
module C_gate2 ( in1, in2, out );
input  in1, in2;
output out;
    adfull_1 U3 ( .co(out), .a(in1), .b(in2), .ci(out) );
endmodule


module mutex ( r1, r2, g1, g2 );
input  r1, r2;
output g1, g2;
    wire gr2, gr1;
    nand2_1 mg2 ( .x(gr2), .a(r2), .b(gr1) );
    nand2_1 U1 ( .x(gr1), .a(r1), .b(gr2) );
    nor3_1 U2 ( .x(g2), .a(gr2), .b(gr2), .c(gr2) );
    nor3_1 U3 ( .x(g1), .a(gr1), .b(gr1), .c(gr1) );
endmodule


module mymux4 ( mux_sel, out, in );
input  [1:0] mux_sel;
input  [0:3] in;
output out;
    mux4_1 U4 ( .x(out), .d0(in[0]), .d1(in[1]), .d2(in[2]), .d3(in[3]), .sl0(
        mux_sel[0]), .sl1(mux_sel[1]) );
endmodule


module sram_latency ( in, out, mux_sel );
input  [1:0] mux_sel;
input  in;
output out;
    wire n1, n2, net1, net2, net3, net4, net5, net6, net7, net8, net9, net10, 
        net11, net12, net13, net14, net15, net16, net17, net18, net19, net20, 
        net21, net22, net23, net24;
    buf_1 U1 ( .x(n1), .a(in) );
    buf_4 U2 ( .x(n2), .a(n1) );
    and2_1 and1 ( .x(net1), .a(n2), .b(n1) );
    and2_1 and2 ( .x(net2), .a(n2), .b(net1) );
    and2_1 and3 ( .x(net3), .a(n2), .b(net2) );
    and2_1 and4 ( .x(net4), .a(n2), .b(net3) );
    and2_1 and5 ( .x(net5), .a(n2), .b(net4) );
    and2_1 and6 ( .x(net6), .a(n2), .b(net5) );
    and2_1 and7 ( .x(net7), .a(n2), .b(net6) );
    and2_1 and8 ( .x(net8), .a(n2), .b(net7) );
    and2_1 and9 ( .x(net9), .a(n2), .b(net8) );
    and2_1 and10 ( .x(net10), .a(n2), .b(net9) );
    and2_1 and11 ( .x(net11), .a(n2), .b(net10) );
    and2_1 and12 ( .x(net12), .a(n2), .b(net11) );
    and2_1 and13 ( .x(net13), .a(n2), .b(net12) );
    and2_1 and14 ( .x(net14), .a(n2), .b(net13) );
    and2_1 and15 ( .x(net15), .a(n2), .b(net14) );
    and2_1 and16 ( .x(net16), .a(n2), .b(net15) );
    and2_1 and17 ( .x(net17), .a(n2), .b(net16) );
    and2_1 and18 ( .x(net18), .a(n2), .b(net17) );
    and2_1 and19 ( .x(net19), .a(n2), .b(net18) );
    and2_1 and20 ( .x(net20), .a(n2), .b(net19) );
    and2_1 and21 ( .x(net21), .a(n2), .b(net20) );
    and2_1 and22 ( .x(net22), .a(n2), .b(net21) );
    and2_1 and23 ( .x(net23), .a(n2), .b(net22) );
    and2_1 and24 ( .x(net24), .a(n2), .b(net23) );
    mymux4 mux ( .mux_sel(mux_sel), .out(out), .in({net3, net6, net12, net24})
         );
endmodule


module delay_shifter ( reset, enable, shift_clk, scan_in, par_out );
output [10:0] par_out;
input  reset, enable, shift_clk, scan_in;
    wire n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12;
    mux2_2 U2 ( .x(n2), .d0(par_out[0]), .sl(enable), .d1(scan_in) );
    mux2_2 U3 ( .x(n3), .d0(par_out[1]), .sl(enable), .d1(par_out[0]) );
    mux2_2 U4 ( .x(n4), .d0(par_out[2]), .sl(enable), .d1(par_out[1]) );
    mux2_2 U5 ( .x(n5), .d0(par_out[3]), .sl(enable), .d1(par_out[2]) );
    mux2_2 U6 ( .x(n6), .d0(par_out[4]), .sl(enable), .d1(par_out[3]) );
    mux2_2 U7 ( .x(n7), .d0(par_out[5]), .sl(enable), .d1(par_out[4]) );
    mux2_2 U8 ( .x(n8), .d0(par_out[6]), .sl(enable), .d1(par_out[5]) );
    mux2_2 U9 ( .x(n9), .d0(par_out[7]), .sl(enable), .d1(par_out[6]) );
    mux2_2 U10 ( .x(n10), .d0(par_out[8]), .sl(enable), .d1(par_out[7]) );
    mux2_2 U11 ( .x(n11), .d0(par_out[9]), .sl(enable), .d1(par_out[8]) );
    inv_2 U12 ( .x(n1), .a(reset) );
    mux2_2 U13 ( .x(n12), .d0(par_out[10]), .sl(enable), .d1(par_out[9]) );
    dffpr_1 par_out_reg_0 ( .q(par_out[0]), .rb(n1), .d(n2), .ck(shift_clk) );
    dffpr_1 par_out_reg_1 ( .q(par_out[1]), .rb(n1), .d(n3), .ck(shift_clk) );
    dffpr_1 par_out_reg_2 ( .q(par_out[2]), .rb(n1), .d(n4), .ck(shift_clk) );
    dffpr_1 par_out_reg_3 ( .q(par_out[3]), .rb(n1), .d(n5), .ck(shift_clk) );
    dffpr_1 par_out_reg_4 ( .q(par_out[4]), .rb(n1), .d(n6), .ck(shift_clk) );
    dffpr_1 par_out_reg_5 ( .q(par_out[5]), .rb(n1), .d(n7), .ck(shift_clk) );
    dffpr_1 par_out_reg_6 ( .q(par_out[6]), .rb(n1), .d(n8), .ck(shift_clk) );
    dffpr_1 par_out_reg_7 ( .q(par_out[7]), .rb(n1), .d(n9), .ck(shift_clk) );
    dffpr_1 par_out_reg_8 ( .q(par_out[8]), .rb(n1), .d(n10), .ck(shift_clk)
         );
    dffpr_1 par_out_reg_9 ( .q(par_out[9]), .rb(n1), .d(n11), .ck(shift_clk)
         );
    dffpr_1 par_out_reg_10 ( .q(par_out[10]), .rb(n1), .d(n12), .ck(shift_clk)
         );
endmodule


module matched_delay32__0_85__1__1_38__1_77 ( in, out, mux_sel );
input  [1:0] mux_sel;
input  in;
output out;
    wire n1, n2, n3, net1, net2, net3, net4, net5, net6, net7, net8, net9, 
        net10, net11, net12, net13, net14, net15, net16, net17, net18, net19, 
        net20;
    buf_1 U1 ( .x(n1), .a(in) );
    buf_4 U2 ( .x(n2), .a(n1) );
    buf_16 U3 ( .x(n3), .a(n2) );
    and2_1 and1 ( .x(net1), .a(n3), .b(n3) );
    and2_1 and2 ( .x(net2), .a(n3), .b(net1) );
    and2_1 and3 ( .x(net3), .a(n3), .b(net2) );
    and2_1 and4 ( .x(net4), .a(n3), .b(net3) );
    and2_1 and5 ( .x(net5), .a(n3), .b(net4) );
    and2_1 and6 ( .x(net6), .a(n3), .b(net5) );
    and2_1 and7 ( .x(net7), .a(n3), .b(net6) );
    and2_1 and8 ( .x(net8), .a(n3), .b(net7) );
    and2_1 and9 ( .x(net9), .a(n3), .b(net8) );
    and2_1 and10 ( .x(net10), .a(n3), .b(net9) );
    and2_1 and11 ( .x(net11), .a(n3), .b(net10) );
    and2_1 and12 ( .x(net12), .a(n3), .b(net11) );
    and2_1 and13 ( .x(net13), .a(n3), .b(net12) );
    and2_1 and14 ( .x(net14), .a(n3), .b(net13) );
    and2_1 and15 ( .x(net15), .a(n3), .b(net14) );
    and2_1 and16 ( .x(net16), .a(n3), .b(net15) );
    and2_1 and17 ( .x(net17), .a(n3), .b(net16) );
    and2_1 and18 ( .x(net18), .a(n3), .b(net17) );
    and2_1 and19 ( .x(net19), .a(n3), .b(net18) );
    and2_1 and20 ( .x(net20), .a(n3), .b(net19) );
    mymux4 mux ( .mux_sel(mux_sel), .out(out), .in({net3, net5, net10, net20})
         );
endmodule


module lc_semi_dec_master ( rst, ri, ai, ro, ao, l );
input  rst, ri, ao;
output ai, ro, l;
    wire lint, aoi1, nri, nrst, nro;
    inv_1 linvg ( .x(l), .a(ai) );
    inv_1 linvi ( .x(lint), .a(ai) );
    aoi23_1 maingate ( .x(ai), .a(aoi1), .b(nri), .c(nri), .d(ro), .e(ao) );
    inv_1 resetinv ( .x(nrst), .a(rst) );
    nand2_1 resetnand ( .x(aoi1), .a(nrst), .b(ai) );
    inv_1 riinv ( .x(nri), .a(ri) );
    aoi21_1 rogate ( .x(ro), .a(nro), .b(ao), .c(lint) );
    inv_1 roint ( .x(nro), .a(ro) );
endmodule


module lc_semi_dec_slave ( rst, ri, ai, ro, ao, l );
input  rst, ri, ao;
output ai, ro, l;
    wire lint, aoi1, nri, nro;
    inv_1 linvg ( .x(l), .a(ai) );
    inv_1 linvi ( .x(lint), .a(ai) );
    aoi23_1 maingate ( .x(ai), .a(aoi1), .b(nri), .c(nri), .d(ro), .e(ao) );
    nor2_1 resetnor ( .x(aoi1), .a(rst), .b(ai) );
    inv_1 riinv ( .x(nri), .a(ri) );
    aoi221_1 rogate ( .x(ro), .a(nro), .b(ao), .c(lint), .d(1'b1), .e(rst) );
    inv_1 roint ( .x(nro), .a(ro) );
endmodule


module controller_d32__0_85__1__1_38__1_77_r1_a2 ( reset, en1, en2, ri1, ai, 
    ro, ao1, ao2, delay_mux_sel );
input  [1:0] delay_mux_sel;
input  reset, ri1, ao1, ao2;
output en1, en2, ai, ro;
    wire ao_synchr, ri_synchr_delayed, rx, ax;
    C_gate2 cgate_ackouts ( .in1(ao1), .in2(ao2), .out(ao_synchr) );
    matched_delay32__0_85__1__1_38__1_77 delay ( .in(ri1), .out(
        ri_synchr_delayed), .mux_sel(delay_mux_sel) );
    lc_semi_dec_master master ( .rst(reset), .ri(ri_synchr_delayed), .ai(ai), 
        .ro(rx), .ao(ax), .l(en1) );
    lc_semi_dec_slave slave ( .rst(reset), .ri(rx), .ai(ax), .ro(ro), .ao(
        ao_synchr), .l(en2) );
endmodule


module matched_delay31__0_85__1__1_47__1_93 ( in, out, mux_sel );
input  [1:0] mux_sel;
input  in;
output out;
    wire n1, n2, n3, net1, net2, net3, net4, net5, net6, net7, net8, net9, 
        net10, net11, net12, net13, net14, net15, net16, net17, net18, net19, 
        net20;
    buf_1 U1 ( .x(n1), .a(in) );
    buf_4 U2 ( .x(n2), .a(n1) );
    buf_16 U3 ( .x(n3), .a(n2) );
    and2_1 and1 ( .x(net1), .a(n3), .b(n3) );
    and2_1 and2 ( .x(net2), .a(n3), .b(net1) );
    and2_1 and3 ( .x(net3), .a(n3), .b(net2) );
    and2_1 and4 ( .x(net4), .a(n3), .b(net3) );
    and2_1 and5 ( .x(net5), .a(n3), .b(net4) );
    and2_1 and6 ( .x(net6), .a(n3), .b(net5) );
    and2_1 and7 ( .x(net7), .a(n3), .b(net6) );
    and2_1 and8 ( .x(net8), .a(n3), .b(net7) );
    and2_1 and9 ( .x(net9), .a(n3), .b(net8) );
    and2_1 and10 ( .x(net10), .a(n3), .b(net9) );
    and2_1 and11 ( .x(net11), .a(n3), .b(net10) );
    and2_1 and12 ( .x(net12), .a(n3), .b(net11) );
    and2_1 and13 ( .x(net13), .a(n3), .b(net12) );
    and2_1 and14 ( .x(net14), .a(n3), .b(net13) );
    and2_1 and15 ( .x(net15), .a(n3), .b(net14) );
    and2_1 and16 ( .x(net16), .a(n3), .b(net15) );
    and2_1 and17 ( .x(net17), .a(n3), .b(net16) );
    and2_1 and18 ( .x(net18), .a(n3), .b(net17) );
    and2_1 and19 ( .x(net19), .a(n3), .b(net18) );
    and2_1 and20 ( .x(net20), .a(n3), .b(net19) );
    mymux4 mux ( .mux_sel(mux_sel), .out(out), .in({net3, net5, net10, net20})
         );
endmodule


module controller_d31__0_85__1__1_47__1_93_r2_a2 ( reset, en1, en2, ri1, ri2, 
    ai, ro, ao1, ao2, delay_mux_sel );
input  [1:0] delay_mux_sel;
input  reset, ri1, ri2, ao1, ao2;
output en1, en2, ai, ro;
    wire ao_synchr, ri_synchr, ri_synchr_delayed, rx, ax;
    C_gate2 cgate_ackouts ( .in1(ao1), .in2(ao2), .out(ao_synchr) );
    C_gate2 cgate_reqins ( .in1(ri1), .in2(ri2), .out(ri_synchr) );
    matched_delay31__0_85__1__1_47__1_93 delay ( .in(ri_synchr), .out(
        ri_synchr_delayed), .mux_sel(delay_mux_sel) );
    lc_semi_dec_master master ( .rst(reset), .ri(ri_synchr_delayed), .ai(ai), 
        .ro(rx), .ao(ax), .l(en1) );
    lc_semi_dec_slave slave ( .rst(reset), .ri(rx), .ai(ax), .ro(ro), .ao(
        ao_synchr), .l(en2) );
endmodule


module matched_delay28__0_85__1__1_48__1_95 ( in, out, mux_sel );
input  [1:0] mux_sel;
input  in;
output out;
    wire n1, n2, n3, net1, net2, net3, net4, net5, net6, net7, net8, net9, 
        net10, net11, net12, net13, net14, net15, net16, net17, net18, net19, 
        net20;
    buf_1 U1 ( .x(n1), .a(in) );
    buf_4 U2 ( .x(n2), .a(n1) );
    buf_16 U3 ( .x(n3), .a(n2) );
    and2_1 and1 ( .x(net1), .a(n3), .b(n3) );
    and2_1 and2 ( .x(net2), .a(n3), .b(net1) );
    and2_1 and3 ( .x(net3), .a(n3), .b(net2) );
    and2_1 and4 ( .x(net4), .a(n3), .b(net3) );
    and2_1 and5 ( .x(net5), .a(n3), .b(net4) );
    and2_1 and6 ( .x(net6), .a(n3), .b(net5) );
    and2_1 and7 ( .x(net7), .a(n3), .b(net6) );
    and2_1 and8 ( .x(net8), .a(n3), .b(net7) );
    and2_1 and9 ( .x(net9), .a(n3), .b(net8) );
    and2_1 and10 ( .x(net10), .a(n3), .b(net9) );
    and2_1 and11 ( .x(net11), .a(n3), .b(net10) );
    and2_1 and12 ( .x(net12), .a(n3), .b(net11) );
    and2_1 and13 ( .x(net13), .a(n3), .b(net12) );
    and2_1 and14 ( .x(net14), .a(n3), .b(net13) );
    and2_1 and15 ( .x(net15), .a(n3), .b(net14) );
    and2_1 and16 ( .x(net16), .a(n3), .b(net15) );
    and2_1 and17 ( .x(net17), .a(n3), .b(net16) );
    and2_1 and18 ( .x(net18), .a(n3), .b(net17) );
    and2_1 and19 ( .x(net19), .a(n3), .b(net18) );
    and2_1 and20 ( .x(net20), .a(n3), .b(net19) );
    mymux4 mux ( .mux_sel(mux_sel), .out(out), .in({net3, net5, net10, net20})
         );
endmodule


module controller_d28__0_85__1__1_48__1_95_r2_a2 ( reset, en1, en2, ri1, ri2, 
    ai, ro, ao1, ao2, delay_mux_sel );
input  [1:0] delay_mux_sel;
input  reset, ri1, ri2, ao1, ao2;
output en1, en2, ai, ro;
    wire ao_synchr, ri_synchr, ri_synchr_delayed, rx, ax;
    C_gate2 cgate_ackouts ( .in1(ao1), .in2(ao2), .out(ao_synchr) );
    C_gate2 cgate_reqins ( .in1(ri1), .in2(ri2), .out(ri_synchr) );
    matched_delay28__0_85__1__1_48__1_95 delay ( .in(ri_synchr), .out(
        ri_synchr_delayed), .mux_sel(delay_mux_sel) );
    lc_semi_dec_master master ( .rst(reset), .ri(ri_synchr_delayed), .ai(ai), 
        .ro(rx), .ao(ax), .l(en1) );
    lc_semi_dec_slave slave ( .rst(reset), .ri(rx), .ai(ax), .ro(ro), .ao(
        ao_synchr), .l(en2) );
endmodule


module matched_delay6__0_85__1__1_18__1_36 ( in, out, mux_sel );
input  [1:0] mux_sel;
input  in;
output out;
    wire n1, n2, net1, net2, net3, net4, net5, net6;
    buf_1 U1 ( .x(n1), .a(in) );
    buf_4 U2 ( .x(n2), .a(n1) );
    and2_1 and1 ( .x(net1), .a(n2), .b(n2) );
    and2_1 and2 ( .x(net2), .a(n2), .b(net1) );
    and2_1 and3 ( .x(net3), .a(n2), .b(net2) );
    and2_1 and4 ( .x(net4), .a(n2), .b(net3) );
    and2_1 and5 ( .x(net5), .a(n2), .b(net4) );
    and2_1 and6 ( .x(net6), .a(n2), .b(net5) );
    mymux4 mux ( .mux_sel(mux_sel), .out(out), .in({net1, net2, net4, net6})
         );
endmodule


module controller_d6__0_85__1__1_18__1_36_r2_a1 ( reset, en1, en2, ri1, ri2, 
    ai, ro, ao1, delay_mux_sel );
input  [1:0] delay_mux_sel;
input  reset, ri1, ri2, ao1;
output en1, en2, ai, ro;
    wire ri_synchr, ri_synchr_delayed, rx, ax;
    C_gate2 cgate_reqins ( .in1(ri1), .in2(ri2), .out(ri_synchr) );
    matched_delay6__0_85__1__1_18__1_36 delay ( .in(ri_synchr), .out(
        ri_synchr_delayed), .mux_sel(delay_mux_sel) );
    lc_semi_dec_master master ( .rst(reset), .ri(ri_synchr_delayed), .ai(ai), 
        .ro(rx), .ao(ax), .l(en1) );
    lc_semi_dec_slave slave ( .rst(reset), .ri(rx), .ai(ax), .ro(ro), .ao(ao1), 
        .l(en2) );
endmodule


module smlatnr_2 ( q, qb, d, sdi, se, g, rb, glob_g, sync_sel );
input  d, sdi, se, g, rb, glob_g, sync_sel;
output q, qb;
    wire data, enable;
    latnr_2 latch ( .q(q), .qb(qb), .rb(rb), .d(data), .g(enable) );
    mux2_1 mux_scan ( .x(data), .d0(d), .sl(se), .d1(sdi) );
    mux2_1 mux_sync ( .x(enable), .d0(glob_g), .sl(sync_sel), .d1(g) );
endmodule


module mlatnr_8 ( q, qb, d, g, rb, glob_g, sync_sel );
input  d, g, rb, glob_g, sync_sel;
output q, qb;
    wire enable;
    latnr_8 latch ( .q(q), .qb(qb), .rb(rb), .d(d), .g(enable) );
    mux2_1 mux_sync ( .x(enable), .d0(glob_g), .sl(sync_sel), .d1(g) );
endmodule


module smlatnr_1 ( q, qb, d, sdi, se, g, rb, glob_g, sync_sel );
input  d, sdi, se, g, rb, glob_g, sync_sel;
output q, qb;
    wire data, enable;
    latnr_1 latch ( .q(q), .qb(qb), .rb(rb), .d(data), .g(enable) );
    mux2_1 mux_scan ( .x(data), .d0(d), .sl(se), .d1(sdi) );
    mux2_1 mux_sync ( .x(enable), .d0(glob_g), .sl(sync_sel), .d1(g) );
endmodule


module mlatnr_4 ( q, qb, d, g, rb, glob_g, sync_sel );
input  d, g, rb, glob_g, sync_sel;
output q, qb;
    wire enable;
    latnr_4 latch ( .q(q), .qb(qb), .rb(rb), .d(d), .g(enable) );
    mux2_1 mux_sync ( .x(enable), .d0(glob_g), .sl(sync_sel), .d1(g) );
endmodule


module mlatnr_2 ( q, qb, d, g, rb, glob_g, sync_sel );
input  d, g, rb, glob_g, sync_sel;
output q, qb;
    wire enable;
    latnr_2 latch ( .q(q), .qb(qb), .rb(rb), .d(d), .g(enable) );
    mux2_1 mux_sync ( .x(enable), .d0(glob_g), .sl(sync_sel), .d1(g) );
endmodule


module mlatnr_1 ( q, qb, d, g, rb, glob_g, sync_sel );
input  d, g, rb, glob_g, sync_sel;
output q, qb;
    wire enable;
    latnr_1 latch ( .q(q), .qb(qb), .rb(rb), .d(d), .g(enable) );
    mux2_1 mux_sync ( .x(enable), .d0(glob_g), .sl(sync_sel), .d1(g) );
endmodule


module EX_DW01_add_32_5_test_1 ( A, B, CI, SUM, CO );
input  [31:0] A;
input  [31:0] B;
output [31:0] SUM;
input  CI;
output CO;
    wire n167, n181, n367, n313, n365, n322, n224, n225, n250, n321, n311, 
        n174, n173, n96, n251, n94, n95, n111, n330, n138, n202, n331, n332, 
        n136, n243, n200, n135, n199, n131, n129, n132, n133, n197, n198, n170, 
        n193, n341, n109, n161, n347, n121, n348, n159, n233, n314, n107, n300, 
        n190, n342, n343, n355, n266, n234, n294, n272, n295, n296, n108, n110, 
        n273, n232, n353, n360, n354, n242, n363, n267, n235, n93, n83, n116, 
        n119, n211, n117, n118, n182, n307, n122, n124, n263, n177, n100, n371, 
        n178, n104, n101, n102, n204, n140, n176, n97, n325, n310, n98, n99, 
        n287, n275, n186, n195, n134, n206, n146, n103, n323, n179, n324, n217, 
        n216, n172, n127, n196, n171, n184, n183, n175, n230, n229, n63, n364, 
        n201, n306, n151, n160, n75, n191, n192, n189, n188, n64, n52, n209, 
        n210, n58, n219, n220, n221, n222, n223, n51, n165, n80, n166, n279, 
        n260, n112, n53, n162, n164, n227, n284, n329, n56, n55, n54, n150, 
        n315, n356, n254, n153, n154, n212, n147, n148, n215, n244, n264, n265, 
        n157, n259, n369, n358, n208, n362, n149, n316, n285, n168, n163, n252, 
        n57, n256, n194, n84, n214, n257, n276, n336, n339, n338, n337, n340, 
        n59, n278, n60, n289, n213, n357, n247, n128, n239, n76, n79, n78, n77, 
        n62, n180, n268, n269, n346, n152, n286, n308, n82, n87, n86, n85, n65, 
        n255, n352, n89, n326, n309, n185, n361, n66, n344, n67, n68, n298, 
        n297, n71, n69, n70, n125, n207, n72, n270, n73, n271, n305, n74, n350, 
        n302, n301, n303, n304, n237, n236, n156, n126, n317, n123, n345, n351, 
        n142, n145, n327, n226, n169, n359, n253, n88, n238, n115, n92, n114, 
        n187, n245, n374, n248, n113, n241, n203, n274, n280, n281, n120, n158, 
        n282, n290, n144, n292, n261, n262, n293, n299, n218, n320, n319, n349, 
        n141, n291, n335, n90, n283, n91, n333, n258, n288, n105, n277, n370, 
        n205, n372, n143, n373, n61, n81, n249, n334, n375, n106, n240, n318, 
        n312, n50, n49, n328, n155, n231, n366, n137, n139, n130, n228, n368;
    exnor2_5 U10 ( .x(SUM[30]), .a(n167), .b(n181) );
    inv_2 U100 ( .x(n367), .a(n313) );
    nand2_0 U101 ( .x(n365), .a(A[0]), .b(B[0]) );
    oai22_1 U102 ( .x(n322), .a(n224), .b(n225), .c(n250), .d(n321) );
    inv_2 U103 ( .x(n250), .a(n311) );
    inv_2 U104 ( .x(n321), .a(n174) );
    inv_2 U107 ( .x(n173), .a(n322) );
    inv_2 U108 ( .x(n96), .a(n251) );
    nor2i_1 U109 ( .x(n94), .a(n95), .b(n96) );
    nor2_2 U11 ( .x(n111), .a(A[15]), .b(B[15]) );
    inv_2 U110 ( .x(n330), .a(n138) );
    nand2i_2 U111 ( .x(n202), .a(n330), .b(n331) );
    inv_2 U112 ( .x(n332), .a(n202) );
    inv_0 U113 ( .x(n136), .a(n243) );
    oai21_1 U114 ( .x(n200), .a(n136), .b(n332), .c(n135) );
    exnor2_1 U115 ( .x(SUM[16]), .a(n199), .b(n131) );
    inv_5 U116 ( .x(n199), .a(n129) );
    nor2i_0 U117 ( .x(n131), .a(n132), .b(n133) );
    exor2_1 U118 ( .x(SUM[17]), .a(n197), .b(n198) );
    nor2_0 U12 ( .x(n170), .a(A[4]), .b(B[4]) );
    nand2i_2 U120 ( .x(n193), .a(n341), .b(n109) );
    inv_2 U121 ( .x(n161), .a(n109) );
    nand2i_0 U122 ( .x(n347), .a(n121), .b(n161) );
    nand2_0 U123 ( .x(n348), .a(A[22]), .b(B[22]) );
    inv_2 U124 ( .x(n341), .a(n159) );
    inv_0 U125 ( .x(n233), .a(B[21]) );
    nand2i_2 U126 ( .x(n314), .a(A[22]), .b(n107) );
    nand2i_2 U127 ( .x(n300), .a(n121), .b(n159) );
    nand2i_2 U128 ( .x(n190), .a(n342), .b(n343) );
    inv_2 U129 ( .x(n355), .a(n266) );
    or3i_2 U130 ( .x(n266), .a(n159), .b(n234), .c(n121) );
    aoi21_1 U131 ( .x(n294), .a(n272), .b(n295), .c(n296) );
    oai31_1 U132 ( .x(n272), .a(n108), .b(n121), .c(n110), .d(n273) );
    nand2i_0 U133 ( .x(n295), .a(B[24]), .b(n232) );
    inv_2 U134 ( .x(n296), .a(n343) );
    inv_2 U135 ( .x(n353), .a(n272) );
    inv_2 U136 ( .x(n234), .a(B[23]) );
    nand2i_2 U137 ( .x(n360), .a(n342), .b(n354) );
    inv_2 U138 ( .x(n342), .a(n295) );
    inv_2 U139 ( .x(n232), .a(A[24]) );
    inv_1 U14 ( .x(n242), .a(n363) );
    inv_2 U140 ( .x(n354), .a(n267) );
    or3i_2 U141 ( .x(n267), .a(n159), .b(n235), .c(n121) );
    inv_2 U142 ( .x(n235), .a(A[23]) );
    inv_2 U143 ( .x(n93), .a(n83) );
    nand2_2 U144 ( .x(n116), .a(A[25]), .b(B[25]) );
    inv_2 U145 ( .x(n119), .a(n211) );
    nor2i_1 U146 ( .x(n117), .a(n118), .b(n119) );
    inv_2 U147 ( .x(n182), .a(n307) );
    exnor2_1 U148 ( .x(SUM[3]), .a(n182), .b(n117) );
    exor2_1 U149 ( .x(SUM[2]), .a(n122), .b(n124) );
    inv_0 U15 ( .x(n263), .a(B[15]) );
    exor2_1 U150 ( .x(SUM[6]), .a(n177), .b(n100) );
    oai21_1 U151 ( .x(n177), .a(n371), .b(n178), .c(n104) );
    nor2i_1 U152 ( .x(n100), .a(n101), .b(n102) );
    exor2_1 U153 ( .x(SUM[12]), .a(n204), .b(n140) );
    exor2_1 U154 ( .x(SUM[7]), .a(n176), .b(n97) );
    oai21_1 U155 ( .x(n176), .a(n102), .b(n325), .c(n101) );
    inv_0 U156 ( .x(n102), .a(n310) );
    inv_2 U157 ( .x(n325), .a(n177) );
    nor2i_1 U158 ( .x(n97), .a(n98), .b(n99) );
    inv_2 U159 ( .x(n99), .a(n287) );
    nand2i_2 U16 ( .x(n275), .a(n138), .b(n243) );
    exor2_1 U160 ( .x(n186), .a(B[27]), .b(A[27]) );
    exor2_1 U162 ( .x(n195), .a(A[20]), .b(B[20]) );
    exor2_1 U163 ( .x(SUM[14]), .a(n202), .b(n134) );
    exor2_1 U164 ( .x(SUM[10]), .a(n206), .b(n146) );
    nor2i_0 U165 ( .x(n103), .a(n104), .b(n371) );
    inv_2 U166 ( .x(n323), .a(n179) );
    aoai211_1 U167 ( .x(n324), .a(n217), .b(n216), .c(n323), .d(n172) );
    inv_2 U168 ( .x(n178), .a(n324) );
    exnor2_1 U169 ( .x(SUM[5]), .a(n178), .b(n103) );
    exnor2_1 U170 ( .x(SUM[19]), .a(n127), .b(n196) );
    exor2_1 U171 ( .x(SUM[4]), .a(n179), .b(n171) );
    exor2_1 U172 ( .x(n184), .a(A[28]), .b(B[28]) );
    exnor2_1 U173 ( .x(SUM[28]), .a(n183), .b(n184) );
    exnor2_1 U174 ( .x(SUM[8]), .a(n174), .b(n175) );
    inv_2 U175 ( .x(n230), .a(B[27]) );
    inv_2 U176 ( .x(n229), .a(A[27]) );
    inv_0 U177 ( .x(n63), .a(n364) );
    exnor2_1 U178 ( .x(SUM[9]), .a(n173), .b(n94) );
    exor2_1 U179 ( .x(SUM[15]), .a(n200), .b(n201) );
    inv_2 U18 ( .x(n306), .a(n151) );
    inv_2 U180 ( .x(n160), .a(n75) );
    exnor2_1 U181 ( .x(SUM[21]), .a(n160), .b(n193) );
    exor2_1 U182 ( .x(SUM[23]), .a(n191), .b(n192) );
    oai211_1 U183 ( .x(n191), .a(n75), .b(n300), .c(n348), .d(n347) );
    exor2_1 U184 ( .x(n192), .a(A[23]), .b(B[23]) );
    exnor2_1 U185 ( .x(SUM[24]), .a(n189), .b(n190) );
    exor2_1 U186 ( .x(n188), .a(B[25]), .b(A[25]) );
    exnor2_1 U187 ( .x(SUM[25]), .a(n93), .b(n188) );
    exnor2_1 U188 ( .x(SUM[29]), .a(n64), .b(n52) );
    inv_2 U189 ( .x(n209), .a(B[1]) );
    inv_2 U19 ( .x(n210), .a(n58) );
    nand4_2 U190 ( .x(n219), .a(n220), .b(n221), .c(n222), .d(n223) );
    ao21_3 U191 ( .x(n51), .a(n165), .b(n80), .c(n166) );
    nand2i_3 U192 ( .x(n279), .a(B[18]), .b(n260) );
    exnor2_1 U193 ( .x(n52), .a(B[29]), .b(A[29]) );
    nor2_1 U194 ( .x(n112), .a(A[17]), .b(B[17]) );
    oai21_1 U195 ( .x(n197), .a(n199), .b(n133), .c(n132) );
    ao21_3 U197 ( .x(n53), .a(n80), .b(n162), .c(n164) );
    nand2i_0 U198 ( .x(n162), .a(B[29]), .b(n227) );
    nand3i_1 U20 ( .x(n223), .a(n284), .b(n310), .c(n287) );
    ao21_4 U200 ( .x(n329), .a(n56), .b(n55), .c(n54) );
    inv_3 U201 ( .x(n55), .a(n219) );
    nand3_1 U202 ( .x(n56), .a(n150), .b(n315), .c(n306) );
    inv_4 U203 ( .x(n356), .a(n254) );
    and3i_4 U204 ( .x(n153), .a(n151), .b(n154), .c(n315) );
    nand3_5 U205 ( .x(n151), .a(n210), .b(n211), .c(n212) );
    nor2i_1 U206 ( .x(n146), .a(n147), .b(n148) );
    inv_2 U208 ( .x(n215), .a(B[6]) );
    nand2i_2 U209 ( .x(n244), .a(A[13]), .b(n264) );
    nand2_0 U21 ( .x(n98), .a(A[7]), .b(B[7]) );
    nand2i_2 U210 ( .x(n243), .a(B[14]), .b(n265) );
    nand2i_2 U211 ( .x(n363), .a(A[15]), .b(n263) );
    nor2_1 U213 ( .x(n157), .a(n111), .b(n135) );
    inv_1 U214 ( .x(n259), .a(A[17]) );
    nand2_0 U215 ( .x(n369), .a(B[1]), .b(A[1]) );
    nand2_0 U216 ( .x(n358), .a(B[1]), .b(A[1]) );
    inv_2 U217 ( .x(n208), .a(A[1]) );
    nand2_1 U218 ( .x(n362), .a(B[1]), .b(A[1]) );
    nor2_2 U219 ( .x(n149), .a(B[1]), .b(A[1]) );
    nand4_1 U22 ( .x(n221), .a(n287), .b(n310), .c(n316), .d(n285) );
    aoi21_3 U220 ( .x(n167), .a(n168), .b(n163), .c(n166) );
    nand2_1 U221 ( .x(n252), .a(n57), .b(n256) );
    inv_1 U222 ( .x(n256), .a(A[10]) );
    exnor2_1 U223 ( .x(SUM[20]), .a(n194), .b(n195) );
    nand2_0 U224 ( .x(n172), .a(B[4]), .b(A[4]) );
    inv_12 U225 ( .x(n216), .a(A[4]) );
    or2_2 U226 ( .x(n147), .a(n256), .b(n84) );
    inv_2 U227 ( .x(n214), .a(B[5]) );
    nand2_5 U228 ( .x(n58), .a(n310), .b(n287) );
    nand2i_2 U23 ( .x(n316), .a(A[5]), .b(n214) );
    inv_1 U230 ( .x(n257), .a(A[11]) );
    exor2_1 U231 ( .x(n201), .a(A[15]), .b(B[15]) );
    aoi21_1 U232 ( .x(n276), .a(A[15]), .b(B[15]), .c(n157) );
    nand4_3 U233 ( .x(n336), .a(n339), .b(n338), .c(n337), .d(n340) );
    inv_0 U234 ( .x(n59), .a(n278) );
    inv_2 U235 ( .x(n60), .a(n59) );
    nand2_0 U236 ( .x(n289), .a(A[8]), .b(B[8]) );
    inv_0 U237 ( .x(n225), .a(A[8]) );
    inv_7 U238 ( .x(n213), .a(A[7]) );
    oai211_3 U239 ( .x(n339), .a(n219), .b(n153), .c(n357), .d(n356) );
    inv_10 U240 ( .x(n357), .a(n247) );
    inv_2 U242 ( .x(n194), .a(n336) );
    nor2i_0 U243 ( .x(n128), .a(n279), .b(n239) );
    oaoi211_2 U244 ( .x(n76), .a(n79), .b(n78), .c(n336), .d(n77) );
    aoai211_1 U245 ( .x(n189), .a(n267), .b(n266), .c(n75), .d(n353) );
    inv_2 U246 ( .x(n62), .a(n180) );
    exor2_1 U247 ( .x(n180), .a(B[31]), .b(A[31]) );
    aoai211_1 U248 ( .x(n64), .a(n268), .b(n269), .c(n63), .d(n346) );
    nand4i_1 U249 ( .x(n220), .a(n152), .b(n310), .c(n287), .d(n286) );
    nor2_1 U25 ( .x(n286), .a(n170), .b(n118) );
    nand2_1 U250 ( .x(n308), .a(B[17]), .b(A[17]) );
    exor2_1 U251 ( .x(SUM[27]), .a(n82), .b(n186) );
    ao221_4 U252 ( .x(n80), .a(n364), .b(n87), .c(n364), .d(n86), .e(n85) );
    inv_0 U253 ( .x(n65), .a(n255) );
    nand2i_2 U254 ( .x(n352), .a(n95), .b(n89) );
    nand3i_1 U255 ( .x(n326), .a(n289), .b(n251), .c(n89) );
    inv_0 U256 ( .x(n148), .a(n89) );
    nand2_1 U257 ( .x(n309), .a(A[16]), .b(B[16]) );
    mx4_4 U258 ( .x(n185), .d0(B[26]), .sl0(A[26]), .d1(n361), .sl1(n66), .d2(
        n344), .sl2(n67), .d3(n361), .sl3(n68) );
    inv_2 U259 ( .x(n66), .a(n298) );
    inv_2 U260 ( .x(n67), .a(n116) );
    inv_2 U261 ( .x(n68), .a(n297) );
    oaoi211_1 U262 ( .x(n71), .a(n69), .b(n260), .c(n278), .d(n70) );
    inv_7 U263 ( .x(n260), .a(A[18]) );
    nand2_4 U264 ( .x(n125), .a(B[2]), .b(A[2]) );
    ao21_2 U265 ( .x(n278), .a(n308), .b(n309), .c(n112) );
    nand2i_6 U266 ( .x(n315), .a(B[2]), .b(n207) );
    nand2_0 U268 ( .x(n104), .a(B[5]), .b(A[5]) );
    nand2_0 U269 ( .x(n284), .a(B[5]), .b(A[5]) );
    inv_2 U27 ( .x(n54), .a(n356) );
    nor2_0 U270 ( .x(n152), .a(A[5]), .b(B[5]) );
    inv_2 U271 ( .x(n72), .a(n270) );
    inv_2 U272 ( .x(n73), .a(n271) );
    inv_0 U273 ( .x(n270), .a(B[30]) );
    inv_2 U274 ( .x(n271), .a(A[30]) );
    nand2_2 U275 ( .x(n305), .a(n306), .b(n307) );
    buf_3 U276 ( .x(n74), .a(n215) );
    inv_2 U279 ( .x(n77), .a(n350) );
    aoi21_1 U28 ( .x(n302), .a(n301), .b(n303), .c(n304) );
    inv_2 U280 ( .x(n78), .a(n237) );
    inv_2 U281 ( .x(n79), .a(n236) );
    nand2_0 U282 ( .x(n350), .a(A[20]), .b(B[20]) );
    inv_0 U283 ( .x(n237), .a(A[20]) );
    inv_0 U284 ( .x(n236), .a(B[20]) );
    nor2_0 U285 ( .x(n156), .a(B[1]), .b(A[1]) );
    nor2i_0 U286 ( .x(n124), .a(n125), .b(n126) );
    inv_2 U287 ( .x(n317), .a(n125) );
    oai211_1 U288 ( .x(n150), .a(n156), .b(n123), .c(n125), .d(n358) );
    aoai211_5 U289 ( .x(n364), .a(n229), .b(n230), .c(n345), .d(n351) );
    nor2_0 U29 ( .x(n301), .a(n142), .b(n145) );
    nand2_0 U290 ( .x(n343), .a(A[24]), .b(B[24]) );
    exor2_1 U291 ( .x(n198), .a(B[17]), .b(A[17]) );
    inv_0 U292 ( .x(n327), .a(n219) );
    ao21_1 U293 ( .x(n175), .a(A[8]), .b(B[8]), .c(n250) );
    inv_0 U294 ( .x(n82), .a(n345) );
    inv_3 U295 ( .x(n226), .a(B[9]) );
    nand2_2 U296 ( .x(n95), .a(B[9]), .b(A[9]) );
    ao221_4 U297 ( .x(n163), .a(n364), .b(n87), .c(n364), .d(n86), .e(n85) );
    nor2_0 U298 ( .x(n169), .a(A[4]), .b(B[4]) );
    aoai211_1 U299 ( .x(n83), .a(n360), .b(n359), .c(n75), .d(n294) );
    inv_0 U30 ( .x(n145), .a(n253) );
    inv_0 U300 ( .x(n84), .a(B[10]) );
    inv_2 U301 ( .x(n85), .a(n346) );
    inv_2 U302 ( .x(n86), .a(n269) );
    inv_2 U303 ( .x(n87), .a(n268) );
    inv_0 U304 ( .x(n183), .a(n364) );
    nand2_0 U305 ( .x(n346), .a(B[28]), .b(A[28]) );
    inv_0 U306 ( .x(n269), .a(B[28]) );
    inv_0 U307 ( .x(n268), .a(A[28]) );
    nand2_2 U308 ( .x(n109), .a(B[21]), .b(A[21]) );
    nand2_0 U309 ( .x(n132), .a(A[16]), .b(B[16]) );
    inv_0 U31 ( .x(n264), .a(B[13]) );
    and2_2 U310 ( .x(n88), .a(A[6]), .b(B[6]) );
    inv_0 U311 ( .x(n101), .a(n88) );
    nand2_1 U312 ( .x(n138), .a(B[13]), .b(A[13]) );
    inv_4 U313 ( .x(n238), .a(B[12]) );
    nor3i_5 U314 ( .x(n115), .a(n116), .b(n92), .c(n114) );
    exnor2_5 U315 ( .x(SUM[26]), .a(n115), .b(n187) );
    inv_6 U316 ( .x(n207), .a(A[2]) );
    nand2i_4 U317 ( .x(n245), .a(n70), .b(n374) );
    or3i_5 U318 ( .x(n247), .a(n248), .b(n113), .c(n241) );
    nand2i_4 U319 ( .x(n254), .a(n142), .b(n255) );
    nand2_3 U32 ( .x(n203), .a(n302), .b(n329) );
    inv_6 U320 ( .x(n265), .a(A[14]) );
    oai21_4 U321 ( .x(n274), .a(n242), .b(n275), .c(n276) );
    exnor2_3 U322 ( .x(n280), .a(n281), .b(n260) );
    mux2i_3 U323 ( .x(SUM[22]), .d0(n120), .sl(n158), .d1(n282) );
    nor2i_5 U324 ( .x(n285), .a(B[4]), .b(n216) );
    nand2_2 U325 ( .x(n290), .a(n144), .b(n147) );
    oai21_4 U326 ( .x(n292), .a(n261), .b(n262), .c(n293) );
    nand2_2 U327 ( .x(n164), .a(n299), .b(n271) );
    exor2_3 U328 ( .x(n181), .a(B[30]), .b(n73) );
    exor2_3 U329 ( .x(n187), .a(A[26]), .b(B[26]) );
    nand2_1 U33 ( .x(n331), .a(n203), .b(n244) );
    nand2i_4 U330 ( .x(n211), .a(B[3]), .b(n218) );
    nand3i_3 U331 ( .x(n307), .a(n317), .b(n320), .c(n319) );
    inv_5 U334 ( .x(n345), .a(n185) );
    oai21_4 U335 ( .x(n206), .a(n173), .b(n96), .c(n95) );
    inv_5 U336 ( .x(n349), .a(n206) );
    nand2i_4 U337 ( .x(n340), .a(n141), .b(n357) );
    nand3i_3 U338 ( .x(n338), .a(n291), .b(n303), .c(n357) );
    nand2i_4 U339 ( .x(n359), .a(n342), .b(n355) );
    nand3_1 U34 ( .x(n241), .a(n363), .b(n243), .c(n244) );
    aoai211_4 U340 ( .x(n337), .a(n248), .b(n274), .c(n292), .d(n335) );
    mux2i_3 U341 ( .x(n90), .d0(n283), .sl(B[18]), .d1(n280) );
    nand2_3 U342 ( .x(SUM[18]), .a(n90), .b(n91) );
    nand2i_6 U344 ( .x(n159), .a(A[21]), .b(n233) );
    nor2i_5 U345 ( .x(n92), .a(B[25]), .b(n93) );
    nor2i_5 U346 ( .x(n114), .a(A[25]), .b(n93) );
    nand2i_6 U347 ( .x(n251), .a(A[9]), .b(n226) );
    nand2i_5 U348 ( .x(n333), .a(n241), .b(n203) );
    inv_10 U349 ( .x(n217), .a(B[4]) );
    inv_2 U35 ( .x(n258), .a(A[16]) );
    nand2i_6 U350 ( .x(n310), .a(A[6]), .b(n74) );
    nand2i_6 U351 ( .x(n287), .a(B[7]), .b(n213) );
    aoi21_4 U352 ( .x(n222), .a(n88), .b(n287), .c(n288) );
    inv_6 U353 ( .x(n248), .a(n245) );
    nand2i_4 U354 ( .x(n291), .a(n142), .b(n253) );
    aoi21_4 U355 ( .x(n212), .a(n217), .b(n216), .c(n105) );
    inv_16 U356 ( .x(n262), .a(A[19]) );
    nor2_8 U357 ( .x(n113), .a(A[19]), .b(B[19]) );
    nor2i_1 U358 ( .x(n283), .a(A[18]), .b(n277) );
    oai21_3 U359 ( .x(n277), .a(n199), .b(n239), .c(n60) );
    nand2_2 U36 ( .x(n273), .a(A[23]), .b(B[23]) );
    inv_0 U360 ( .x(n370), .a(n105) );
    inv_2 U361 ( .x(n371), .a(n370) );
    inv_3 U362 ( .x(n105), .a(n316) );
    exnor2_1 U363 ( .x(SUM[11]), .a(n205), .b(n372) );
    inv_2 U364 ( .x(n372), .a(n143) );
    oai21_2 U365 ( .x(n205), .a(n148), .b(n349), .c(n147) );
    nor2i_0 U366 ( .x(n143), .a(n144), .b(n373) );
    oai211_1 U367 ( .x(n154), .a(n149), .b(n123), .c(n125), .d(n362) );
    nand2_3 U368 ( .x(n123), .a(B[0]), .b(A[0]) );
    oaoi211_2 U369 ( .x(n75), .a(n79), .b(n78), .c(n61), .d(n77) );
    nor2_1 U37 ( .x(n110), .a(A[23]), .b(B[23]) );
    inv_4 U370 ( .x(n61), .a(n194) );
    nand2_1 U371 ( .x(n174), .a(n81), .b(n305) );
    inv_2 U372 ( .x(n81), .a(n219) );
    inv_0 U373 ( .x(n373), .a(n253) );
    nand2i_3 U374 ( .x(n253), .a(B[11]), .b(n257) );
    inv_4 U375 ( .x(n255), .a(n249) );
    nand4i_3 U376 ( .x(n249), .a(n250), .b(n251), .c(n89), .d(n253) );
    buf_6 U377 ( .x(n89), .a(n252) );
    nor2i_3 U378 ( .x(n374), .a(n334), .b(n375) );
    inv_0 U379 ( .x(n239), .a(n374) );
    nor2i_1 U38 ( .x(n108), .a(n109), .b(n106) );
    inv_5 U380 ( .x(n375), .a(n240) );
    inv_0 U381 ( .x(n133), .a(n334) );
    nand2i_2 U382 ( .x(n240), .a(B[17]), .b(n259) );
    nand2i_2 U383 ( .x(n334), .a(B[16]), .b(n258) );
    aoai211_3 U384 ( .x(n361), .a(n360), .b(n359), .c(n76), .d(n294) );
    nor2i_1 U39 ( .x(n106), .a(A[22]), .b(n107) );
    inv_2 U40 ( .x(n107), .a(B[22]) );
    nand3i_1 U41 ( .x(n319), .a(n149), .b(n315), .c(n318) );
    or3i_2 U42 ( .x(n320), .a(n315), .b(n209), .c(n208) );
    inv_2 U43 ( .x(n126), .a(n315) );
    aoi21_1 U44 ( .x(n122), .a(n123), .b(n369), .c(n367) );
    nand2i_2 U45 ( .x(n313), .a(B[1]), .b(n208) );
    inv_2 U46 ( .x(n318), .a(n123) );
    nand2i_2 U47 ( .x(n312), .a(A[12]), .b(n238) );
    inv_2 U48 ( .x(n142), .a(n312) );
    nand2_0 U49 ( .x(n141), .a(A[12]), .b(B[12]) );
    exnor2_3 U5 ( .x(SUM[31]), .a(n50), .b(n49) );
    nor2i_1 U50 ( .x(n140), .a(n141), .b(n142) );
    nand2i_2 U51 ( .x(n328), .a(n373), .b(n303) );
    aoai211_1 U53 ( .x(n204), .a(n327), .b(n305), .c(n65), .d(n328) );
    inv_2 U54 ( .x(n288), .a(n98) );
    nand2i_2 U55 ( .x(n297), .a(n155), .b(B[25]) );
    nand2i_2 U56 ( .x(n298), .a(n155), .b(A[25]) );
    nand2i_2 U57 ( .x(n344), .a(B[26]), .b(n231) );
    inv_2 U58 ( .x(n231), .a(A[26]) );
    inv_2 U59 ( .x(n155), .a(n344) );
    inv_2 U6 ( .x(n49), .a(n62) );
    nor2i_1 U60 ( .x(SUM[0]), .a(n365), .b(n366) );
    nor2_1 U61 ( .x(n366), .a(B[0]), .b(A[0]) );
    nand2_1 U62 ( .x(n144), .a(A[11]), .b(B[11]) );
    inv_2 U64 ( .x(n304), .a(n141) );
    nand2i_2 U65 ( .x(n335), .a(B[19]), .b(n262) );
    inv_2 U66 ( .x(n261), .a(B[19]) );
    nand3i_2 U67 ( .x(n303), .a(n290), .b(n352), .c(n326) );
    nand2_1 U68 ( .x(n135), .a(A[14]), .b(B[14]) );
    nor2i_1 U69 ( .x(n134), .a(n135), .b(n136) );
    aoi22_1 U7 ( .x(n50), .a(n51), .b(n73), .c(n53), .d(n72) );
    exor2_1 U70 ( .x(SUM[13]), .a(n203), .b(n137) );
    nor2i_1 U71 ( .x(n137), .a(n138), .b(n139) );
    inv_2 U72 ( .x(n139), .a(n244) );
    inv_1 U73 ( .x(n57), .a(B[10]) );
    aoi21_1 U74 ( .x(n158), .a(n159), .b(n160), .c(n161) );
    exnor2_1 U75 ( .x(n282), .a(A[22]), .b(B[22]) );
    aoi21_1 U76 ( .x(n120), .a(A[22]), .b(B[22]), .c(n121) );
    inv_3 U77 ( .x(n121), .a(n314) );
    exor2_1 U78 ( .x(n196), .a(A[19]), .b(B[19]) );
    inv_2 U79 ( .x(n70), .a(n279) );
    nand2i_2 U8 ( .x(n311), .a(A[8]), .b(n224) );
    inv_0 U80 ( .x(n69), .a(B[18]) );
    inv_2 U81 ( .x(n293), .a(n71) );
    inv_0 U82 ( .x(n130), .a(n293) );
    nand2i_3 U83 ( .x(n129), .a(n274), .b(n333) );
    aoi21_1 U84 ( .x(n127), .a(n128), .b(n129), .c(n130) );
    nor2i_1 U85 ( .x(n171), .a(n172), .b(n169) );
    oai21_1 U86 ( .x(n179), .a(n119), .b(n182), .c(n118) );
    inv_0 U87 ( .x(n218), .a(A[3]) );
    nand2_1 U88 ( .x(n118), .a(A[3]), .b(B[3]) );
    nand2i_0 U89 ( .x(n91), .a(n279), .b(n277) );
    inv_3 U9 ( .x(n224), .a(B[8]) );
    inv_2 U90 ( .x(n281), .a(n277) );
    inv_2 U91 ( .x(n228), .a(B[29]) );
    nand2i_2 U92 ( .x(n168), .a(A[29]), .b(n228) );
    nand2_2 U93 ( .x(n351), .a(B[27]), .b(A[27]) );
    nand2i_2 U94 ( .x(n165), .a(B[29]), .b(n227) );
    inv_2 U95 ( .x(n227), .a(A[29]) );
    inv_2 U96 ( .x(n166), .a(n299) );
    nand2_2 U97 ( .x(n299), .a(B[29]), .b(A[29]) );
    exnor2_1 U98 ( .x(SUM[1]), .a(n368), .b(n365) );
    nor2i_1 U99 ( .x(n368), .a(n369), .b(n367) );
endmodule


module EX_DW01_add_32_6_test_1 ( A, B, CI, SUM, CO );
input  [31:0] A;
input  [31:0] B;
output [31:0] SUM;
input  CI;
output CO;
    wire n350, n89, n239, n241, n240, n336, n147, n367, n84, n366, n54, n140, 
        n139, n200, n56, n255, n331, n204, n298, n342, n190, n384, n153, n154, 
        n155, n79, n275, n361, n260, n363, n196, n227, n132, n226, n225, n82, 
        n278, n371, n370, n145, n198, n50, n164, n223, n224, n379, n288, n364, 
        n365, n326, n222, n220, n188, n283, n282, n289, n51, n141, n230, n146, 
        n181, n382, n148, n302, n236, n166, n167, n168, n131, n129, n115, n118, 
        n237, n169, n238, n103, n344, n170, n171, n229, n157, n160, n165, n372, 
        n161, n162, n158, n235, n378, n318, n307, n163, n386, n172, n144, n195, 
        n299, n211, n123, n85, n348, n212, n86, n124, n125, n149, n231, n107, 
        n126, n143, n142, n110, n111, n300, n296, n295, n292, n206, n214, n216, 
        n209, n210, n61, n351, n305, n215, n62, n286, n287, n208, n112, n353, 
        n252, n253, n313, n352, n346, n113, n114, n159, n156, n234, n100, n99, 
        n265, n310, n77, n221, n201, n301, n52, n347, n249, n128, n315, n312, 
        n93, n246, n55, n58, n81, n245, n57, n228, n83, n106, n381, n380, n325, 
        n327, n192, n174, n373, n60, n59, n262, n261, n75, n243, n244, n53, 
        n120, n134, n135, n242, n349, n273, n175, n185, n355, n268, n78, n274, 
        n314, n284, n285, n63, n369, n217, n329, n64, n105, n330, n183, n193, 
        n66, n65, n194, n173, n279, n67, n68, n280, n95, n176, n177, n178, 
        n319, n320, n97, n69, n306, n71, n70, n328, n186, n290, n270, n291, 
        n339, n316, n189, n119, n116, n121, n72, n130, n73, n74, n179, n76, 
        n213, n203, n199, n80, n375, n266, n98, n138, n356, n383, n256, n257, 
        n368, n374, n308, n309, n324, n377, n271, n376, n127, n109, n218, n88, 
        n362, n137, n264, n340, n94, n136, n187, n90, n250, n104, n205, n281, 
        n91, n311, n357, n258, n96, n294, n293, n49, n191, n122, n303, n101, 
        n385, n102, n259, n233, n108, n333, n254, n202, n334, n182, n184, n219, 
        n197, n232, n263, n269, n276, n277, n297, n304, n322, n321, n323, n317, 
        n92, n354, n180, n345, n247, n133, n335, n337, n358, n359, n338, n207, 
        n87, n267, n343, n248, n251, n332, n117, n272, n150, n151, n152, n341;
    ao211_2 U10 ( .x(n350), .a(n89), .b(n239), .c(n241), .d(n240) );
    inv_2 U100 ( .x(n336), .a(n147) );
    nand2_1 U101 ( .x(n147), .a(B[2]), .b(A[2]) );
    nand3_3 U102 ( .x(n367), .a(n84), .b(n366), .c(n54) );
    inv_2 U103 ( .x(n140), .a(B[26]) );
    nor2i_1 U104 ( .x(n139), .a(A[26]), .b(n140) );
    nand2i_2 U105 ( .x(n200), .a(n56), .b(n255) );
    nand2_2 U106 ( .x(n331), .a(n56), .b(A[29]) );
    inv_2 U107 ( .x(n255), .a(A[29]) );
    nand2i_2 U108 ( .x(n204), .a(n56), .b(n255) );
    oai21_1 U109 ( .x(n298), .a(A[1]), .b(B[1]), .c(n342) );
    inv_0 U11 ( .x(n190), .a(n350) );
    exor2_1 U110 ( .x(SUM[1]), .a(n298), .b(n384) );
    nor2i_1 U111 ( .x(n153), .a(n154), .b(n155) );
    inv_2 U112 ( .x(n79), .a(n275) );
    inv_2 U113 ( .x(n155), .a(n361) );
    inv_0 U114 ( .x(n260), .a(B[21]) );
    inv_2 U115 ( .x(n363), .a(n196) );
    nand2i_2 U116 ( .x(n227), .a(n363), .b(n132) );
    exor2_1 U117 ( .x(n226), .a(A[23]), .b(B[23]) );
    oai211_1 U118 ( .x(n225), .a(n82), .b(n278), .c(n371), .d(n370) );
    nand2i_2 U119 ( .x(n370), .a(n145), .b(n198) );
    buf_1 U12 ( .x(n50), .a(n164) );
    inv_2 U120 ( .x(n198), .a(n132) );
    exnor2_1 U121 ( .x(SUM[24]), .a(n223), .b(n224) );
    inv_0 U122 ( .x(n379), .a(n288) );
    nand2i_2 U123 ( .x(n224), .a(n364), .b(n365) );
    inv_2 U124 ( .x(n364), .a(n326) );
    exor2_1 U125 ( .x(n222), .a(n54), .b(A[25]) );
    exor2_1 U126 ( .x(n220), .a(A[26]), .b(B[26]) );
    nand2_2 U127 ( .x(n188), .a(A[25]), .b(n54) );
    inv_2 U128 ( .x(n283), .a(A[25]) );
    inv_2 U129 ( .x(n282), .a(n54) );
    nand2_0 U13 ( .x(n289), .a(A[23]), .b(B[23]) );
    exnor2_1 U130 ( .x(SUM[3]), .a(n51), .b(n141) );
    exor2_1 U131 ( .x(SUM[2]), .a(n230), .b(n146) );
    oai21_1 U132 ( .x(n230), .a(n384), .b(n181), .c(n342) );
    inv_7 U133 ( .x(n181), .a(n382) );
    nor2i_1 U134 ( .x(n146), .a(n147), .b(n148) );
    inv_2 U135 ( .x(n148), .a(n302) );
    exor2_1 U136 ( .x(SUM[12]), .a(n236), .b(n166) );
    nor2i_1 U138 ( .x(n166), .a(n167), .b(n168) );
    nor2i_1 U14 ( .x(n131), .a(n132), .b(n129) );
    exnor2_1 U140 ( .x(SUM[7]), .a(n115), .b(n118) );
    exor2_1 U141 ( .x(SUM[11]), .a(n237), .b(n169) );
    ao21_2 U142 ( .x(n237), .a(n238), .b(n103), .c(n344) );
    nor2i_1 U143 ( .x(n169), .a(n170), .b(n171) );
    exor2_1 U144 ( .x(n229), .a(A[20]), .b(B[20]) );
    exor2_1 U145 ( .x(SUM[14]), .a(n157), .b(n160) );
    oai21_1 U146 ( .x(n157), .a(n165), .b(n372), .c(n50) );
    nor2i_1 U147 ( .x(n160), .a(n161), .b(n162) );
    inv_0 U148 ( .x(n162), .a(n158) );
    inv_2 U149 ( .x(n372), .a(n235) );
    nand2i_2 U15 ( .x(n378), .a(n318), .b(n307) );
    nor2i_1 U150 ( .x(n163), .a(n50), .b(n165) );
    inv_2 U151 ( .x(n168), .a(n275) );
    oai21_1 U152 ( .x(n235), .a(n386), .b(n168), .c(n167) );
    exor2_1 U153 ( .x(SUM[13]), .a(n235), .b(n163) );
    exor2_1 U154 ( .x(SUM[10]), .a(n238), .b(n172) );
    mux2i_1 U155 ( .x(SUM[22]), .d0(n144), .sl(n195), .d1(n299) );
    exor2_1 U156 ( .x(SUM[5]), .a(n211), .b(n123) );
    aoi21_1 U157 ( .x(n85), .a(n348), .b(n212), .c(n86) );
    nor2i_1 U158 ( .x(n123), .a(n124), .b(n125) );
    exnor2_1 U159 ( .x(SUM[19]), .a(n149), .b(n231) );
    inv_6 U16 ( .x(n107), .a(A[6]) );
    exor2_1 U160 ( .x(SUM[4]), .a(n212), .b(n126) );
    oai21_1 U161 ( .x(n212), .a(n143), .b(n51), .c(n142) );
    nand2_2 U162 ( .x(SUM[18]), .a(n110), .b(n111) );
    mux2i_1 U163 ( .x(n110), .d0(n300), .sl(B[18]), .d1(n296) );
    nand2i_2 U164 ( .x(n111), .a(n295), .b(n292) );
    exnor2_3 U165 ( .x(SUM[30]), .a(n206), .b(n214) );
    exor2_1 U166 ( .x(n216), .a(A[28]), .b(B[28]) );
    exnor2_1 U167 ( .x(SUM[8]), .a(n209), .b(n210) );
    oai211_1 U168 ( .x(n209), .a(n51), .b(n61), .c(n351), .d(n305) );
    exor2_1 U169 ( .x(n215), .a(n56), .b(A[29]) );
    inv_0 U17 ( .x(n62), .a(B[2]) );
    inv_2 U170 ( .x(n286), .a(B[30]) );
    inv_2 U171 ( .x(n287), .a(A[30]) );
    exnor2_1 U172 ( .x(SUM[9]), .a(n208), .b(n112) );
    oai22_1 U173 ( .x(n353), .a(n252), .b(n253), .c(n313), .d(n352) );
    inv_5 U174 ( .x(n313), .a(n346) );
    inv_2 U175 ( .x(n352), .a(n209) );
    nor2i_0 U176 ( .x(n112), .a(n113), .b(n114) );
    inv_2 U177 ( .x(n159), .a(n161) );
    aoi21_1 U178 ( .x(n156), .a(n157), .b(n158), .c(n159) );
    exnor2_1 U179 ( .x(SUM[15]), .a(n156), .b(n234) );
    aoai211_1 U18 ( .x(n100), .a(n99), .b(n265), .c(n164), .d(n310) );
    exnor2_1 U180 ( .x(SUM[16]), .a(n77), .b(n153) );
    exor2_1 U181 ( .x(SUM[23]), .a(n225), .b(n226) );
    exnor2_1 U182 ( .x(SUM[25]), .a(n221), .b(n222) );
    exor2_1 U183 ( .x(SUM[29]), .a(n201), .b(n215) );
    oa211_2 U184 ( .x(n51), .a(n384), .b(n301), .c(n350), .d(n147) );
    exnor2_1 U186 ( .x(n52), .a(B[31]), .b(A[31]) );
    inv_2 U187 ( .x(n143), .a(n347) );
    nand2i_2 U188 ( .x(n347), .a(B[3]), .b(n249) );
    inv_2 U189 ( .x(n128), .a(n348) );
    inv_5 U19 ( .x(n315), .a(n312) );
    nand2_2 U190 ( .x(n348), .a(n93), .b(n246) );
    buf_3 U191 ( .x(n54), .a(B[25]) );
    inv_0 U192 ( .x(n55), .a(B[29]) );
    inv_2 U193 ( .x(n56), .a(n55) );
    inv_2 U194 ( .x(n58), .a(n81) );
    inv_6 U195 ( .x(n245), .a(A[5]) );
    aoi21_2 U196 ( .x(n57), .a(n228), .b(n83), .c(n106) );
    aoai211_3 U197 ( .x(n84), .a(n381), .b(n380), .c(n57), .d(n325) );
    aoi21_2 U198 ( .x(n325), .a(n288), .b(n326), .c(n327) );
    and3i_1 U20 ( .x(n192), .a(n174), .b(A[9]), .c(B[9]) );
    inv_2 U200 ( .x(n106), .a(n373) );
    nand2_4 U201 ( .x(n60), .a(n59), .b(n262) );
    inv_4 U202 ( .x(n59), .a(B[17]) );
    inv_7 U203 ( .x(n262), .a(A[17]) );
    inv_5 U204 ( .x(n261), .a(A[16]) );
    inv_1 U205 ( .x(n75), .a(B[10]) );
    nand2_2 U207 ( .x(n142), .a(A[3]), .b(B[3]) );
    nand3_1 U208 ( .x(n61), .a(n243), .b(n244), .c(n347) );
    nor2_3 U209 ( .x(n243), .a(n53), .b(n120) );
    nor2i_0 U21 ( .x(n134), .a(B[18]), .b(n135) );
    nand3_2 U210 ( .x(n242), .a(n243), .b(n244), .c(n347) );
    nand2i_3 U211 ( .x(n349), .a(B[5]), .b(n245) );
    oa22_4 U212 ( .x(n77), .a(n273), .b(n175), .c(n386), .d(n185) );
    nand2i_3 U213 ( .x(n355), .a(A[15]), .b(n268) );
    and4i_4 U214 ( .x(n78), .a(n79), .b(n355), .c(n274), .d(n158) );
    inv_2 U215 ( .x(n273), .a(n355) );
    ao21_6 U216 ( .x(n314), .a(n62), .b(n239), .c(n315) );
    aoai211_3 U217 ( .x(n201), .a(n284), .b(n285), .c(n63), .d(n369) );
    nand3i_5 U218 ( .x(n217), .a(n139), .b(n367), .c(n329) );
    aoai211_3 U219 ( .x(n64), .a(n381), .b(n380), .c(n105), .d(n325) );
    inv_8 U22 ( .x(n135), .a(A[18]) );
    aoai211_1 U220 ( .x(n330), .a(n381), .b(n380), .c(n58), .d(n325) );
    and3i_3 U221 ( .x(n183), .a(n193), .b(n66), .c(n65) );
    inv_2 U222 ( .x(n65), .a(n192) );
    or3_5 U223 ( .x(n66), .a(n174), .b(n114), .c(n194) );
    nand2_2 U224 ( .x(n193), .a(n170), .b(n173) );
    inv_2 U225 ( .x(n279), .a(n67) );
    inv_2 U226 ( .x(n68), .a(B[23]) );
    inv_0 U227 ( .x(n280), .a(n278) );
    ao31_6 U228 ( .x(n95), .a(n176), .b(n161), .c(n177), .d(n178) );
    nor2i_3 U229 ( .x(n319), .a(A[4]), .b(n320) );
    inv_5 U23 ( .x(n97), .a(B[16]) );
    inv_5 U230 ( .x(n93), .a(A[4]) );
    buf_1 U231 ( .x(n69), .a(n228) );
    nand2i_2 U233 ( .x(n306), .a(B[5]), .b(n245) );
    ao21_4 U234 ( .x(n238), .a(n353), .b(n71), .c(n70) );
    inv_2 U235 ( .x(n70), .a(n113) );
    inv_0 U236 ( .x(n71), .a(n114) );
    inv_0 U237 ( .x(n208), .a(n353) );
    aoi21_3 U238 ( .x(n329), .a(n64), .b(n328), .c(n186) );
    inv_5 U239 ( .x(n268), .a(B[15]) );
    nand2i_0 U24 ( .x(n290), .a(n270), .b(n291) );
    exor2_1 U240 ( .x(n234), .a(A[15]), .b(B[15]) );
    nand2_0 U241 ( .x(n339), .a(A[15]), .b(B[15]) );
    nand2_1 U242 ( .x(n310), .a(A[15]), .b(B[15]) );
    nor3_5 U243 ( .x(n316), .a(n189), .b(n314), .c(n242) );
    nand2_1 U244 ( .x(n119), .a(A[7]), .b(B[7]) );
    exor2_1 U245 ( .x(SUM[6]), .a(n116), .b(n121) );
    inv_0 U246 ( .x(n72), .a(n130) );
    or2_2 U247 ( .x(n365), .a(n73), .b(n74) );
    inv_1 U248 ( .x(n74), .a(B[24]) );
    and2_2 U249 ( .x(n179), .a(n75), .b(n76) );
    inv_3 U25 ( .x(n270), .a(n60) );
    inv_4 U250 ( .x(n241), .a(B[1]) );
    oai22_2 U251 ( .x(n213), .a(n203), .b(n287), .c(n199), .d(n286) );
    inv_6 U252 ( .x(n185), .a(n78) );
    and3_1 U253 ( .x(n175), .a(n80), .b(n176), .c(n375) );
    and2_1 U254 ( .x(n80), .a(n339), .b(n161) );
    nand2i_2 U255 ( .x(n275), .a(B[12]), .b(n266) );
    inv_1 U256 ( .x(n98), .a(B[17]) );
    inv_2 U257 ( .x(n82), .a(n81) );
    inv_2 U258 ( .x(n83), .a(n138) );
    nand4i_1 U259 ( .x(n381), .a(n145), .b(n196), .c(A[23]), .d(n326) );
    nand2_2 U26 ( .x(n291), .a(n97), .b(n261) );
    inv_14 U260 ( .x(n99), .a(B[14]) );
    exor2_1 U261 ( .x(SUM[20]), .a(n69), .b(n229) );
    nand3_4 U262 ( .x(n176), .a(n274), .b(n158), .c(n356) );
    nand2i_0 U263 ( .x(n375), .a(n164), .b(n158) );
    nand2i_4 U264 ( .x(n161), .a(n265), .b(B[14]) );
    aoai211_5 U265 ( .x(n383), .a(n256), .b(n257), .c(n368), .d(n374) );
    inv_10 U266 ( .x(n368), .a(n217) );
    inv_16 U267 ( .x(n265), .a(A[14]) );
    aoi31_1 U268 ( .x(n305), .a(n306), .b(n307), .c(n308), .d(n309) );
    nand4i_5 U269 ( .x(n324), .a(n309), .b(n351), .c(n377), .d(n378) );
    inv_2 U27 ( .x(n271), .a(n291) );
    inv_6 U270 ( .x(n309), .a(n376) );
    inv_0 U271 ( .x(n211), .a(n85) );
    inv_2 U272 ( .x(n86), .a(n127) );
    nand2_0 U273 ( .x(n127), .a(n109), .b(A[4]) );
    exor2_1 U274 ( .x(SUM[27]), .a(n217), .b(n218) );
    aoai211_2 U275 ( .x(n88), .a(n256), .b(n257), .c(n368), .d(n374) );
    inv_10 U276 ( .x(n240), .a(A[1]) );
    ao23_6 U277 ( .x(n362), .a(n137), .b(n264), .c(n95), .d(n340), .e(n94) );
    inv_2 U278 ( .x(n94), .a(n136) );
    inv_0 U279 ( .x(n264), .a(A[19]) );
    nor2_1 U28 ( .x(n186), .a(n187), .b(n188) );
    inv_2 U280 ( .x(n90), .a(B[7]) );
    inv_6 U281 ( .x(n250), .a(B[6]) );
    aoi21_3 U282 ( .x(n203), .a(n204), .b(n104), .c(n205) );
    inv_2 U283 ( .x(n205), .a(n331) );
    inv_0 U284 ( .x(n281), .a(n91) );
    nand2i_2 U286 ( .x(n178), .a(n273), .b(n311) );
    nand2i_6 U287 ( .x(n302), .a(B[2]), .b(n239) );
    aoai211_1 U288 ( .x(n223), .a(n281), .b(n279), .c(n82), .d(n379) );
    nand2i_2 U289 ( .x(n357), .a(B[10]), .b(n76) );
    nand2i_2 U29 ( .x(n366), .a(B[26]), .b(n258) );
    nor2i_0 U290 ( .x(n136), .a(A[19]), .b(n137) );
    nand2_0 U291 ( .x(n124), .a(B[5]), .b(A[5]) );
    nand2_0 U292 ( .x(n318), .a(B[5]), .b(A[5]) );
    aoi211_1 U293 ( .x(n96), .a(n262), .b(n98), .c(n261), .d(n97) );
    inv_0 U294 ( .x(n294), .a(n96) );
    nand2_1 U295 ( .x(n293), .a(B[17]), .b(A[17]) );
    nor2_5 U296 ( .x(n189), .a(n49), .b(n191) );
    inv_3 U297 ( .x(n177), .a(n100) );
    nor2i_0 U298 ( .x(n121), .a(n122), .b(n53) );
    nor2_2 U299 ( .x(n303), .a(n53), .b(n120) );
    inv_2 U30 ( .x(n258), .a(A[26]) );
    inv_0 U300 ( .x(n101), .a(n53) );
    nor2_0 U301 ( .x(n385), .a(B[0]), .b(A[0]) );
    inv_0 U302 ( .x(n102), .a(n357) );
    inv_2 U303 ( .x(n103), .a(n102) );
    oai21_3 U304 ( .x(n191), .a(n384), .b(n181), .c(n147) );
    nor2i_0 U305 ( .x(n126), .a(n127), .b(n128) );
    nand2i_2 U306 ( .x(n326), .a(B[24]), .b(n259) );
    exor2_1 U307 ( .x(n233), .a(B[17]), .b(A[17]) );
    ao221_4 U308 ( .x(n104), .a(n383), .b(A[28]), .c(n383), .d(B[28]), .e(n108
        ) );
    nand2_2 U309 ( .x(n194), .a(A[8]), .b(B[8]) );
    inv_2 U31 ( .x(n187), .a(n366) );
    ao21_1 U310 ( .x(n210), .a(A[8]), .b(B[8]), .c(n313) );
    inv_0 U311 ( .x(n252), .a(B[8]) );
    nand2_0 U312 ( .x(n373), .a(A[20]), .b(B[20]) );
    nand2_0 U313 ( .x(n333), .a(A[9]), .b(B[9]) );
    inv_3 U314 ( .x(n254), .a(B[9]) );
    nand2_0 U315 ( .x(n113), .a(B[9]), .b(A[9]) );
    exnor2_1 U316 ( .x(SUM[28]), .a(n63), .b(n216) );
    aoi21_2 U317 ( .x(n199), .a(n200), .b(n104), .c(n202) );
    exnor2_3 U318 ( .x(SUM[31]), .a(n213), .b(n52) );
    inv_2 U319 ( .x(n108), .a(n369) );
    nand2_2 U32 ( .x(n374), .a(B[27]), .b(A[27]) );
    nand2_0 U320 ( .x(n369), .a(B[28]), .b(A[28]) );
    inv_0 U321 ( .x(n285), .a(B[28]) );
    inv_0 U322 ( .x(n284), .a(A[28]) );
    inv_0 U323 ( .x(n109), .a(n246) );
    nand2_2 U324 ( .x(n132), .a(B[21]), .b(A[21]) );
    nand2i_0 U325 ( .x(n361), .a(B[16]), .b(n261) );
    nand2_0 U326 ( .x(n154), .a(A[16]), .b(B[16]) );
    nor2i_0 U327 ( .x(n172), .a(n173), .b(n174) );
    oai211_1 U328 ( .x(n334), .a(n174), .b(n333), .c(n170), .d(n173) );
    inv_0 U329 ( .x(n344), .a(n173) );
    inv_0 U33 ( .x(n165), .a(n274) );
    nand2_2 U330 ( .x(n167), .a(A[12]), .b(B[12]) );
    nand2_0 U331 ( .x(n173), .a(A[10]), .b(B[10]) );
    nor3_4 U332 ( .x(n182), .a(n183), .b(n184), .c(n185) );
    exor2_3 U333 ( .x(SUM[26]), .a(n219), .b(n220) );
    exnor2_3 U334 ( .x(SUM[21]), .a(n197), .b(n227) );
    exor2_3 U335 ( .x(SUM[17]), .a(n232), .b(n233) );
    inv_6 U336 ( .x(n263), .a(B[18]) );
    inv_6 U337 ( .x(n266), .a(A[12]) );
    ao211_5 U338 ( .x(n269), .a(n135), .b(n263), .c(n270), .d(n271) );
    or3i_5 U339 ( .x(n276), .a(n277), .b(n179), .c(n114) );
    nand2_6 U34 ( .x(n158), .a(n99), .b(n265) );
    nand2i_4 U340 ( .x(n295), .a(B[18]), .b(n135) );
    exnor2_3 U341 ( .x(n296), .a(n297), .b(n135) );
    nand2i_4 U342 ( .x(n301), .a(n181), .b(n302) );
    nor2_5 U343 ( .x(n304), .a(n125), .b(n142) );
    nor2_5 U344 ( .x(n277), .a(n171), .b(n313) );
    nor3_4 U346 ( .x(n322), .a(n321), .b(n185), .c(n276) );
    aoi22_3 U347 ( .x(n323), .a(n316), .b(n317), .c(n324), .d(n322) );
    nand2_2 U348 ( .x(n202), .a(n331), .b(n287) );
    nand2i_4 U349 ( .x(n346), .a(B[8]), .b(n253) );
    nor2_0 U35 ( .x(n138), .a(A[20]), .b(B[20]) );
    oai221_3 U350 ( .x(n219), .a(n221), .b(n282), .c(n221), .d(n283), .e(n188)
         );
    nand2_2 U351 ( .x(n371), .a(A[22]), .b(n72) );
    oai21_4 U352 ( .x(n232), .a(n77), .b(n155), .c(n154) );
    nand2_8 U353 ( .x(n384), .a(A[0]), .b(B[0]) );
    nand3i_5 U354 ( .x(n228), .a(n182), .b(n362), .c(n323) );
    inv_6 U355 ( .x(n221), .a(n330) );
    inv_7 U356 ( .x(n174), .a(n357) );
    nand2i_6 U358 ( .x(n196), .a(A[21]), .b(n260) );
    nand3_4 U359 ( .x(n351), .a(n303), .b(n348), .c(n304) );
    nor2i_1 U36 ( .x(n91), .a(n280), .b(n92) );
    nand2i_6 U360 ( .x(n354), .a(A[9]), .b(n254) );
    nor2_6 U361 ( .x(n180), .a(n384), .b(n181) );
    nand2i_6 U363 ( .x(n345), .a(A[22]), .b(n130) );
    nor2i_5 U364 ( .x(n328), .a(A[25]), .b(n187) );
    inv_10 U365 ( .x(n256), .a(A[27]) );
    inv_8 U366 ( .x(n257), .a(B[27]) );
    inv_6 U367 ( .x(n307), .a(n247) );
    nand3_5 U368 ( .x(n377), .a(n307), .b(B[4]), .c(n319) );
    nand2i_6 U369 ( .x(n312), .a(A[19]), .b(n137) );
    nand2i_2 U37 ( .x(n278), .a(n145), .b(n196) );
    nor2_8 U371 ( .x(n133), .a(A[23]), .b(B[23]) );
    nand2i_6 U372 ( .x(n382), .a(B[1]), .b(n240) );
    nor2i_8 U373 ( .x(n129), .a(A[22]), .b(n130) );
    oa211_4 U374 ( .x(n386), .a(n335), .b(n337), .c(n358), .d(n359) );
    inv_0 U375 ( .x(n236), .a(n386) );
    nand2i_1 U376 ( .x(n337), .a(n276), .b(n338) );
    oai31_1 U377 ( .x(n335), .a(n190), .b(n336), .c(n180), .d(n302) );
    inv_5 U378 ( .x(n63), .a(n88) );
    aoi21_3 U379 ( .x(n206), .a(n207), .b(n201), .c(n205) );
    inv_2 U38 ( .x(n92), .a(A[23]) );
    nand3i_2 U380 ( .x(n184), .a(n171), .b(n312), .c(n311) );
    nand2i_2 U381 ( .x(n321), .a(n315), .b(n311) );
    and3i_4 U382 ( .x(n317), .a(n185), .b(n87), .c(n311) );
    inv_7 U383 ( .x(n311), .a(n269) );
    inv_4 U384 ( .x(n267), .a(B[13]) );
    aoi21_5 U385 ( .x(n105), .a(n228), .b(n83), .c(n106) );
    inv_2 U39 ( .x(n73), .a(A[24]) );
    inv_2 U40 ( .x(n327), .a(n365) );
    oai31_1 U41 ( .x(n288), .a(n131), .b(n145), .c(n133), .d(n289) );
    nand2_3 U42 ( .x(n380), .a(n67), .b(n326) );
    nor2_3 U43 ( .x(n67), .a(n278), .b(n68) );
    inv_5 U44 ( .x(n130), .a(B[22]) );
    inv_2 U45 ( .x(n259), .a(A[24]) );
    nor2i_1 U46 ( .x(n141), .a(n142), .b(n143) );
    nand2_0 U47 ( .x(n342), .a(B[1]), .b(A[1]) );
    or2_3 U48 ( .x(n122), .a(n107), .b(n250) );
    inv_4 U49 ( .x(n171), .a(n343) );
    nand2i_2 U5 ( .x(n248), .a(B[7]), .b(n251) );
    inv_5 U50 ( .x(n114), .a(n354) );
    nor2_0 U51 ( .x(n332), .a(n114), .b(n194) );
    aoai211_1 U52 ( .x(n359), .a(n332), .b(n103), .c(n334), .d(n343) );
    nand2i_2 U53 ( .x(n358), .a(n276), .b(n324) );
    inv_5 U54 ( .x(n239), .a(A[2]) );
    inv_1 U55 ( .x(n89), .a(B[2]) );
    nor2i_1 U57 ( .x(n118), .a(n119), .b(n120) );
    aoi21_1 U58 ( .x(n115), .a(n116), .b(n101), .c(n117) );
    oai21_1 U59 ( .x(n116), .a(n125), .b(n85), .c(n124) );
    ao22_3 U6 ( .x(n247), .a(n107), .b(n250), .c(n90), .d(n251) );
    inv_4 U60 ( .x(n125), .a(n349) );
    and2_3 U61 ( .x(n53), .a(n107), .b(n250) );
    inv_0 U62 ( .x(n117), .a(n122) );
    exor2_1 U63 ( .x(n218), .a(B[27]), .b(A[27]) );
    nor2i_1 U64 ( .x(SUM[0]), .a(n384), .b(n385) );
    inv_2 U65 ( .x(n272), .a(B[11]) );
    nand2i_3 U66 ( .x(n343), .a(A[11]), .b(n272) );
    nand2_0 U67 ( .x(n170), .a(A[11]), .b(B[11]) );
    inv_4 U68 ( .x(n87), .a(n276) );
    inv_2 U69 ( .x(n137), .a(B[19]) );
    inv_3 U7 ( .x(n251), .a(A[7]) );
    nand2i_3 U70 ( .x(n274), .a(A[13]), .b(n267) );
    nand2i_2 U71 ( .x(n164), .a(n267), .b(A[13]) );
    inv_2 U72 ( .x(n356), .a(n167) );
    inv_4 U73 ( .x(n253), .a(A[8]) );
    inv_2 U74 ( .x(n81), .a(n105) );
    inv_1 U75 ( .x(n197), .a(n58) );
    aoi21_1 U76 ( .x(n195), .a(n196), .b(n197), .c(n198) );
    exnor2_1 U77 ( .x(n299), .a(A[22]), .b(n72) );
    aoi21_1 U78 ( .x(n144), .a(A[22]), .b(n72), .c(n145) );
    inv_5 U79 ( .x(n145), .a(n345) );
    inv_4 U8 ( .x(n76), .a(A[10]) );
    exor2_1 U80 ( .x(n231), .a(A[19]), .b(B[19]) );
    aoi21_1 U81 ( .x(n149), .a(n150), .b(n151), .c(n152) );
    nor2i_1 U82 ( .x(n150), .a(n295), .b(n290) );
    inv_0 U83 ( .x(n151), .a(n77) );
    inv_0 U84 ( .x(n152), .a(n340) );
    oai31_1 U85 ( .x(n340), .a(n134), .b(n96), .c(n341), .d(n295) );
    inv_2 U86 ( .x(n341), .a(n293) );
    inv_2 U87 ( .x(n246), .a(B[4]) );
    nor2i_0 U88 ( .x(n300), .a(A[18]), .b(n292) );
    oai211_1 U89 ( .x(n292), .a(n77), .b(n290), .c(n293), .d(n294) );
    inv_2 U9 ( .x(n49), .a(n350) );
    inv_2 U90 ( .x(n297), .a(n292) );
    exor2_1 U91 ( .x(n214), .a(B[30]), .b(A[30]) );
    nand2i_2 U92 ( .x(n207), .a(A[29]), .b(n55) );
    inv_2 U93 ( .x(n320), .a(n306) );
    ao21_3 U94 ( .x(n376), .a(n119), .b(n122), .c(n120) );
    nand2_2 U95 ( .x(n308), .a(n127), .b(n124) );
    inv_5 U96 ( .x(n120), .a(n248) );
    aoi21_2 U97 ( .x(n244), .a(n93), .b(n246), .c(n125) );
    inv_0 U98 ( .x(n249), .a(A[3]) );
    inv_2 U99 ( .x(n338), .a(n61) );
endmodule


module EX_DW01_add_32_4_test_1 ( A, B, CI, SUM, CO );
input  [31:0] A;
input  [31:0] B;
output [31:0] SUM;
input  CI;
output CO;
    wire n336, n110, n150, n285, n148, n182, n328, n329, n222, n261, n98, n100, 
        n262, n342, n224, n255, n225, n256, n58, n60, n181, n361, n281, n279, 
        n280, n344, n349, n343, n350, n180, n104, n105, n83, n103, n264, n127, 
        n232, n84, n174, n106, n107, n108, n111, n113, n168, n91, n50, n67, 
        n311, n196, n129, n167, n254, n88, n89, n90, n273, n178, n71, n197, 
        n132, n137, n338, n136, n133, n134, n242, n187, n194, n123, n102, n316, 
        n317, n124, n125, n318, n128, n233, n126, n195, n198, n135, n164, n87, 
        n86, n144, n146, n112, n114, n351, n99, n147, n149, n270, n109, n95, 
        n302, n93, n94, n310, n208, n207, n309, n163, n169, n245, n116, n188, 
        n170, n162, n203, n293, n161, n82, n267, n265, n173, n176, n54, n70, 
        n219, n175, n165, n166, n260, n357, n354, n85, n308, n214, n215, n240, 
        n307, n295, n241, n192, n193, n191, n120, n189, n190, n327, n185, n141, 
        n202, n204, n183, n184, n74, n73, n51, n52, n145, n53, n57, n252, n244, 
        n239, n122, n121, n62, n160, n228, n229, n320, n345, n206, n253, n186, 
        n337, n75, n322, n77, n210, n59, n211, n212, n213, n55, n56, n92, n319, 
        n65, n205, n294, n248, n358, n138, n348, n142, n96, n97, n153, n257, 
        n258, n69, n335, n353, n288, n275, n341, n312, n63, n246, n274, n304, 
        n177, n333, n332, n331, n61, n230, n231, n64, n68, n157, n284, n199, 
        n352, n291, n315, n139, n346, n66, n79, n76, n306, n301, n201, n200, 
        n263, n282, n283, n140, n115, n151, n152, n154, n101, n298, n334, n247, 
        n171, n72, n172, n303, n356, n355, n278, n290, n216, n339, n78, n226, 
        n80, n272, n227, n220, n340, n299, n179, n296, n234, n235, n236, n259, 
        n268, n359, n249, n277, n250, n251, n130, n131, n209, n305, n321, n156, 
        n217, n314, n243, n326, n347, n324, n276, n323, n238, n81, n271, n300, 
        n223, n292, n118, n360, n266, n313, n364, n325, n143, n363, n159, n330, 
        n221, n362, n155, n237, n49, n287, n289, n286, n119, n117, n218, n297;
    nand2i_2 U100 ( .x(n336), .a(n110), .b(n150) );
    nand2i_2 U101 ( .x(n285), .a(n110), .b(n148) );
    nand2i_2 U102 ( .x(n182), .a(n328), .b(n329) );
    inv_2 U103 ( .x(n222), .a(A[24]) );
    oai31_2 U104 ( .x(n261), .a(n98), .b(n110), .c(n100), .d(n262) );
    inv_2 U105 ( .x(n342), .a(n261) );
    inv_0 U106 ( .x(n224), .a(B[23]) );
    or3i_2 U107 ( .x(n255), .a(n148), .b(n224), .c(n110) );
    inv_2 U108 ( .x(n225), .a(A[23]) );
    or3i_2 U109 ( .x(n256), .a(n148), .b(n225), .c(n110) );
    inv_2 U11 ( .x(n58), .a(n60) );
    aoai211_1 U110 ( .x(n181), .a(n256), .b(n255), .c(n361), .d(n342) );
    inv_2 U111 ( .x(n281), .a(n329) );
    aoi21_1 U112 ( .x(n279), .a(n261), .b(n280), .c(n281) );
    inv_2 U113 ( .x(n344), .a(n255) );
    nand2i_2 U114 ( .x(n349), .a(n328), .b(n344) );
    inv_2 U115 ( .x(n343), .a(n256) );
    inv_2 U116 ( .x(n328), .a(n280) );
    nand2i_2 U117 ( .x(n350), .a(n328), .b(n343) );
    exor2_1 U118 ( .x(n180), .a(B[25]), .b(A[25]) );
    nor3i_2 U119 ( .x(n104), .a(n105), .b(n83), .c(n103) );
    nand2i_2 U12 ( .x(n264), .a(n127), .b(n232) );
    nand2_2 U120 ( .x(n105), .a(A[25]), .b(B[25]) );
    nor2i_3 U121 ( .x(n83), .a(B[25]), .b(n84) );
    exnor2_1 U122 ( .x(SUM[3]), .a(n174), .b(n106) );
    nor2i_1 U123 ( .x(n106), .a(n107), .b(n108) );
    exor2_1 U124 ( .x(SUM[2]), .a(n111), .b(n113) );
    exor2_1 U125 ( .x(SUM[6]), .a(n168), .b(n91) );
    nor2i_1 U126 ( .x(n91), .a(n50), .b(n67) );
    inv_2 U127 ( .x(n311), .a(n168) );
    exor2_1 U128 ( .x(SUM[12]), .a(n196), .b(n129) );
    oai21_1 U129 ( .x(n167), .a(n67), .b(n311), .c(n50) );
    inv_2 U13 ( .x(n254), .a(A[14]) );
    nor2i_1 U130 ( .x(n88), .a(n89), .b(n90) );
    inv_5 U131 ( .x(n90), .a(n273) );
    exor2_1 U132 ( .x(n178), .a(B[27]), .b(A[27]) );
    exor2_1 U133 ( .x(SUM[27]), .a(n71), .b(n178) );
    exor2_1 U134 ( .x(SUM[11]), .a(n197), .b(n132) );
    oai21_1 U135 ( .x(n197), .a(n137), .b(n338), .c(n136) );
    nor2i_1 U136 ( .x(n132), .a(n133), .b(n134) );
    inv_2 U137 ( .x(n134), .a(n242) );
    exor2_1 U138 ( .x(n187), .a(A[20]), .b(B[20]) );
    exor2_1 U139 ( .x(SUM[14]), .a(n194), .b(n123) );
    nor2_1 U14 ( .x(n102), .a(A[19]), .b(B[19]) );
    nand2i_2 U140 ( .x(n194), .a(n316), .b(n317) );
    nor2i_1 U141 ( .x(n123), .a(n124), .b(n125) );
    inv_2 U142 ( .x(n125), .a(n232) );
    inv_2 U143 ( .x(n318), .a(n194) );
    inv_2 U144 ( .x(n128), .a(n233) );
    nor2i_1 U145 ( .x(n126), .a(n127), .b(n128) );
    exor2_1 U146 ( .x(SUM[13]), .a(n195), .b(n126) );
    exor2_1 U147 ( .x(SUM[10]), .a(n198), .b(n135) );
    oai21_1 U148 ( .x(n198), .a(n164), .b(n87), .c(n86) );
    nor2i_0 U149 ( .x(n135), .a(n136), .b(n137) );
    oai211_1 U15 ( .x(n144), .a(n146), .b(n112), .c(n114), .d(n351) );
    inv_2 U150 ( .x(n338), .a(n198) );
    inv_2 U151 ( .x(n150), .a(n99) );
    aoi21_1 U152 ( .x(n147), .a(n148), .b(n149), .c(n150) );
    exnor2_1 U153 ( .x(n270), .a(A[22]), .b(B[22]) );
    aoi21_1 U154 ( .x(n109), .a(A[22]), .b(B[22]), .c(n110) );
    mux2i_1 U155 ( .x(SUM[22]), .d0(n109), .sl(n147), .d1(n270) );
    inv_2 U156 ( .x(n95), .a(n302) );
    nor2i_1 U157 ( .x(n93), .a(n94), .b(n95) );
    aoai211_1 U158 ( .x(n310), .a(n208), .b(n207), .c(n309), .d(n163) );
    exnor2_1 U159 ( .x(SUM[5]), .a(n169), .b(n93) );
    inv_0 U16 ( .x(n245), .a(A[10]) );
    exnor2_1 U160 ( .x(SUM[19]), .a(n116), .b(n188) );
    exor2_1 U161 ( .x(SUM[4]), .a(n170), .b(n162) );
    oai21_1 U162 ( .x(n170), .a(n108), .b(n174), .c(n107) );
    inv_2 U163 ( .x(n108), .a(n203) );
    inv_2 U164 ( .x(n174), .a(n293) );
    nor2i_1 U165 ( .x(n162), .a(n163), .b(n161) );
    inv_2 U166 ( .x(n309), .a(n170) );
    nand2i_2 U167 ( .x(n82), .a(n267), .b(n265) );
    exor2_1 U168 ( .x(n173), .a(B[30]), .b(A[30]) );
    exor2_1 U169 ( .x(n176), .a(A[28]), .b(B[28]) );
    nand2_2 U17 ( .x(n54), .a(n70), .b(n245) );
    inv_2 U170 ( .x(n219), .a(A[27]) );
    exnor2_1 U171 ( .x(SUM[28]), .a(n175), .b(n176) );
    exnor2_1 U172 ( .x(SUM[8]), .a(n165), .b(n166) );
    inv_2 U173 ( .x(n260), .a(A[30]) );
    exnor2_1 U175 ( .x(SUM[1]), .a(n357), .b(n354) );
    exnor2_1 U176 ( .x(SUM[9]), .a(n164), .b(n85) );
    inv_2 U177 ( .x(n164), .a(n308) );
    oai22_1 U178 ( .x(n308), .a(n214), .b(n215), .c(n240), .d(n307) );
    inv_2 U179 ( .x(n240), .a(n295) );
    inv_1 U18 ( .x(n70), .a(B[10]) );
    inv_2 U180 ( .x(n307), .a(n165) );
    nor2i_1 U181 ( .x(n85), .a(n86), .b(n87) );
    inv_2 U182 ( .x(n87), .a(n241) );
    exor2_1 U183 ( .x(SUM[15]), .a(n192), .b(n193) );
    exnor2_1 U184 ( .x(SUM[16]), .a(n191), .b(n120) );
    exor2_1 U186 ( .x(SUM[17]), .a(n189), .b(n190) );
    inv_2 U187 ( .x(n327), .a(n148) );
    nand2i_2 U188 ( .x(n185), .a(n327), .b(n99) );
    exnor2_1 U189 ( .x(SUM[21]), .a(n149), .b(n185) );
    nand3_3 U19 ( .x(n141), .a(n202), .b(n203), .c(n204) );
    exor2_1 U190 ( .x(SUM[23]), .a(n183), .b(n184) );
    exnor2_1 U191 ( .x(SUM[24]), .a(n181), .b(n182) );
    exnor2_1 U192 ( .x(SUM[25]), .a(n84), .b(n180) );
    inv_2 U193 ( .x(n74), .a(n73) );
    nand2_0 U194 ( .x(n50), .a(A[6]), .b(B[6]) );
    exnor2_1 U195 ( .x(n51), .a(B[29]), .b(A[29]) );
    or2_2 U196 ( .x(n52), .a(n145), .b(n105) );
    oa22_4 U197 ( .x(n53), .a(n57), .b(n252), .c(n124), .d(n58) );
    inv_2 U198 ( .x(n244), .a(n239) );
    oai21_1 U199 ( .x(n189), .a(n191), .b(n122), .c(n121) );
    or2_2 U20 ( .x(n62), .a(n160), .b(n107) );
    nand2i_4 U200 ( .x(n228), .a(n122), .b(n229) );
    inv_5 U201 ( .x(n122), .a(n320) );
    nand2i_0 U202 ( .x(n345), .a(A[5]), .b(n206) );
    nand2i_2 U203 ( .x(n233), .a(A[13]), .b(n253) );
    exnor2_1 U204 ( .x(SUM[20]), .a(n186), .b(n187) );
    oai211_1 U205 ( .x(n183), .a(n361), .b(n285), .c(n337), .d(n336) );
    oaoi211_1 U206 ( .x(n75), .a(B[20]), .b(A[20]), .c(n322), .d(n77) );
    nand2i_2 U207 ( .x(n302), .a(A[5]), .b(n206) );
    nand4_4 U208 ( .x(n210), .a(n59), .b(n211), .c(n212), .d(n213) );
    nor3i_5 U209 ( .x(n55), .a(n56), .b(n92), .c(n90) );
    nand2i_2 U21 ( .x(n319), .a(n65), .b(n195) );
    and2_1 U210 ( .x(n56), .a(B[5]), .b(A[5]) );
    nand2i_3 U211 ( .x(n273), .a(B[7]), .b(n205) );
    or2_8 U212 ( .x(n294), .a(A[6]), .b(B[6]) );
    inv_7 U213 ( .x(n92), .a(n294) );
    inv_1 U214 ( .x(n248), .a(A[17]) );
    nand2_0 U215 ( .x(n358), .a(n74), .b(A[1]) );
    nor2_1 U216 ( .x(n138), .a(n74), .b(A[1]) );
    nand2_2 U217 ( .x(n348), .a(n74), .b(A[1]) );
    nor2_1 U218 ( .x(n142), .a(n74), .b(A[1]) );
    nand2_1 U219 ( .x(n351), .a(B[1]), .b(A[1]) );
    nor2i_0 U22 ( .x(n96), .a(A[22]), .b(n97) );
    aoai211_4 U222 ( .x(n153), .a(n257), .b(n258), .c(n69), .d(n335) );
    inv_6 U223 ( .x(n69), .a(n353) );
    nand3i_2 U224 ( .x(n288), .a(n275), .b(n341), .c(n312) );
    nand2i_2 U225 ( .x(n341), .a(n86), .b(n54) );
    nor2_1 U226 ( .x(n160), .a(A[4]), .b(B[4]) );
    nor2_0 U227 ( .x(n161), .a(A[4]), .b(B[4]) );
    nand2_0 U228 ( .x(n163), .a(B[4]), .b(A[4]) );
    inv_12 U229 ( .x(n207), .a(A[4]) );
    nor2i_1 U23 ( .x(n98), .a(n99), .b(n96) );
    or2_1 U230 ( .x(n63), .a(A[5]), .b(B[5]) );
    inv_2 U231 ( .x(n206), .a(B[5]) );
    exor2_1 U232 ( .x(n193), .a(A[15]), .b(B[15]) );
    inv_2 U233 ( .x(n252), .a(B[15]) );
    inv_2 U234 ( .x(n246), .a(A[11]) );
    nand2_0 U235 ( .x(n274), .a(A[8]), .b(B[8]) );
    inv_0 U236 ( .x(n215), .a(A[8]) );
    inv_7 U237 ( .x(n205), .a(A[7]) );
    nand2_0 U238 ( .x(n89), .a(A[7]), .b(B[7]) );
    inv_0 U239 ( .x(n57), .a(A[15]) );
    inv_0 U24 ( .x(n304), .a(n112) );
    nand4_1 U240 ( .x(n177), .a(n333), .b(n332), .c(n331), .d(n52) );
    aoi23_1 U242 ( .x(n212), .a(A[7]), .b(B[7]), .c(A[6]), .d(B[6]), .e(n273)
         );
    nand2i_4 U243 ( .x(n232), .a(B[14]), .b(n254) );
    or2_2 U244 ( .x(n60), .a(A[15]), .b(B[15]) );
    and4i_5 U245 ( .x(n61), .a(n62), .b(n63), .c(n294), .d(n273) );
    nand3i_3 U246 ( .x(n230), .a(n231), .b(n232), .c(n233) );
    inv_2 U247 ( .x(n64), .a(n68) );
    inv_2 U249 ( .x(n157), .a(n284) );
    inv_2 U25 ( .x(n199), .a(A[2]) );
    nand2i_5 U250 ( .x(n352), .a(A[15]), .b(n252) );
    nand2i_2 U251 ( .x(n165), .a(n210), .b(n291) );
    oai21_1 U252 ( .x(n315), .a(n139), .b(n210), .c(n346) );
    nand3i_0 U253 ( .x(n65), .a(n231), .b(n232), .c(n233) );
    inv_10 U254 ( .x(n231), .a(n352) );
    inv_0 U255 ( .x(n66), .a(n92) );
    inv_2 U256 ( .x(n67), .a(n66) );
    aoai211_3 U257 ( .x(n79), .a(n350), .b(n349), .c(n76), .d(n279) );
    nand2_5 U259 ( .x(n114), .a(B[2]), .b(A[2]) );
    or3i_2 U26 ( .x(n306), .a(n301), .b(n201), .c(n200) );
    oai21_5 U260 ( .x(n263), .a(n231), .b(n264), .c(n53) );
    nand2i_2 U261 ( .x(n333), .a(n282), .b(n79) );
    nand2i_2 U262 ( .x(n332), .a(n283), .b(n79) );
    nor3i_2 U263 ( .x(n139), .a(n140), .b(n115), .c(n141) );
    aoi21_2 U265 ( .x(n151), .a(n152), .b(n153), .c(n154) );
    nor2_1 U266 ( .x(n101), .a(A[17]), .b(B[17]) );
    nand2_1 U267 ( .x(n298), .a(B[17]), .b(A[17]) );
    inv_4 U268 ( .x(n334), .a(n177) );
    inv_0 U269 ( .x(n71), .a(n334) );
    inv_2 U27 ( .x(n201), .a(n74) );
    nand2_1 U270 ( .x(n329), .a(A[24]), .b(B[24]) );
    nand2i_2 U271 ( .x(n320), .a(A[16]), .b(n247) );
    nand2_0 U272 ( .x(n94), .a(B[5]), .b(A[5]) );
    exnor2_3 U273 ( .x(SUM[31]), .a(n171), .b(n72) );
    inv_2 U274 ( .x(n72), .a(n172) );
    exor2_1 U275 ( .x(n172), .a(B[31]), .b(A[31]) );
    nor2i_0 U276 ( .x(n113), .a(n114), .b(n115) );
    inv_1 U277 ( .x(n303), .a(n114) );
    oai211_1 U278 ( .x(n140), .a(n142), .b(n112), .c(n114), .d(n348) );
    nand3i_1 U279 ( .x(n312), .a(n274), .b(n241), .c(n54) );
    aoi21_1 U28 ( .x(n111), .a(n112), .b(n358), .c(n356) );
    inv_0 U280 ( .x(n137), .a(n54) );
    nand4i_1 U281 ( .x(n239), .a(n240), .b(n54), .c(n241), .d(n242) );
    nand2_0 U282 ( .x(n354), .a(A[0]), .b(B[0]) );
    nor2_0 U283 ( .x(n355), .a(B[0]), .b(A[0]) );
    aoai211_2 U284 ( .x(n278), .a(B[18]), .b(A[18]), .c(n290), .d(n267) );
    nand2i_2 U285 ( .x(n280), .a(B[24]), .b(n222) );
    exor2_1 U286 ( .x(n190), .a(B[17]), .b(A[17]) );
    inv_3 U287 ( .x(n214), .a(B[8]) );
    ao21_1 U288 ( .x(n166), .a(A[8]), .b(B[8]), .c(n240) );
    inv_3 U289 ( .x(n216), .a(B[9]) );
    nand2_2 U29 ( .x(n112), .a(B[0]), .b(A[0]) );
    inv_2 U291 ( .x(n77), .a(n339) );
    inv_2 U292 ( .x(n78), .a(n226) );
    nand2_0 U293 ( .x(n339), .a(A[20]), .b(B[20]) );
    inv_0 U294 ( .x(n226), .a(B[20]) );
    inv_0 U295 ( .x(n186), .a(n322) );
    aoai211_1 U296 ( .x(n80), .a(n350), .b(n349), .c(n75), .d(n279) );
    nand4_1 U297 ( .x(n211), .a(n273), .b(n294), .c(n345), .d(n272) );
    nand2_0 U299 ( .x(n335), .a(B[28]), .b(A[28]) );
    inv_0 U30 ( .x(n227), .a(B[12]) );
    inv_0 U300 ( .x(n258), .a(B[28]) );
    inv_0 U301 ( .x(n257), .a(A[28]) );
    aoai211_3 U302 ( .x(n353), .a(n219), .b(n220), .c(n334), .d(n340) );
    nand2_2 U303 ( .x(n99), .a(B[21]), .b(A[21]) );
    nand2_1 U304 ( .x(n299), .a(B[16]), .b(A[16]) );
    nand2_0 U305 ( .x(n121), .a(B[16]), .b(A[16]) );
    exor2_3 U306 ( .x(SUM[7]), .a(n167), .b(n88) );
    exnor2_5 U308 ( .x(SUM[26]), .a(n104), .b(n179) );
    nand2_5 U309 ( .x(n107), .a(A[3]), .b(B[3]) );
    nand2i_0 U31 ( .x(n296), .a(A[12]), .b(n227) );
    nand2i_4 U310 ( .x(n234), .a(n235), .b(n236) );
    inv_6 U311 ( .x(n259), .a(B[30]) );
    exnor2_3 U312 ( .x(n268), .a(n359), .b(n249) );
    nor2_5 U313 ( .x(n202), .a(n92), .b(n90) );
    nor2i_5 U314 ( .x(n272), .a(B[4]), .b(n207) );
    nand2_2 U315 ( .x(n275), .a(n133), .b(n136) );
    oai21_4 U316 ( .x(n277), .a(n250), .b(n251), .c(n278) );
    nand2_2 U317 ( .x(n154), .a(n284), .b(n260) );
    exor2_3 U318 ( .x(n179), .a(A[26]), .b(B[26]) );
    nor2i_1 U32 ( .x(n129), .a(n130), .b(n131) );
    nand2i_4 U320 ( .x(n301), .a(B[2]), .b(n199) );
    nand2i_4 U321 ( .x(n203), .a(B[3]), .b(n209) );
    nand3i_3 U322 ( .x(n305), .a(n138), .b(n301), .c(n304) );
    nand3i_3 U323 ( .x(n293), .a(n303), .b(n306), .c(n305) );
    inv_5 U324 ( .x(n169), .a(n310) );
    oai21_4 U325 ( .x(n168), .a(n95), .b(n169), .c(n94) );
    nand2i_4 U326 ( .x(n242), .a(B[11]), .b(n246) );
    nand2i_4 U327 ( .x(n229), .a(B[17]), .b(n248) );
    nand2i_4 U328 ( .x(n321), .a(B[19]), .b(n251) );
    nand2i_4 U329 ( .x(n156), .a(B[29]), .b(n217) );
    nand2i_2 U33 ( .x(n314), .a(n134), .b(n288) );
    nand2_2 U330 ( .x(n337), .a(A[22]), .b(B[22]) );
    inv_5 U331 ( .x(n346), .a(n243) );
    nand2i_4 U332 ( .x(n326), .a(n130), .b(n347) );
    nand3i_3 U333 ( .x(n324), .a(n276), .b(n288), .c(n347) );
    aoai211_4 U334 ( .x(n323), .a(n238), .b(n263), .c(n277), .d(n321) );
    mux2i_3 U335 ( .x(n81), .d0(n271), .sl(B[18]), .d1(n268) );
    nand2_4 U336 ( .x(SUM[18]), .a(n81), .b(n82) );
    inv_6 U337 ( .x(n84), .a(n80) );
    inv_7 U338 ( .x(n110), .a(n300) );
    nand2i_6 U339 ( .x(n148), .a(A[21]), .b(n223) );
    inv_0 U34 ( .x(n292), .a(n141) );
    nor2i_5 U340 ( .x(n103), .a(A[25]), .b(n84) );
    nand2i_6 U341 ( .x(n241), .a(A[9]), .b(n216) );
    inv_10 U342 ( .x(n220), .a(B[27]) );
    inv_10 U343 ( .x(n208), .a(B[4]) );
    nor2_8 U344 ( .x(n100), .a(A[23]), .b(B[23]) );
    nand2_4 U345 ( .x(n262), .a(A[23]), .b(B[23]) );
    aoi21_4 U346 ( .x(n204), .a(n208), .b(n207), .c(n95) );
    aoi21_3 U347 ( .x(n359), .a(n118), .b(n236), .c(n360) );
    inv_3 U348 ( .x(n265), .a(n359) );
    inv_0 U349 ( .x(n360), .a(n266) );
    aoai211_1 U35 ( .x(n196), .a(n313), .b(n291), .c(n364), .d(n314) );
    inv_0 U350 ( .x(n191), .a(n118) );
    ao21_2 U351 ( .x(n266), .a(n298), .b(n299), .c(n101) );
    inv_5 U352 ( .x(n236), .a(n228) );
    nand2i_2 U353 ( .x(n118), .a(n263), .b(n319) );
    buf_3 U354 ( .x(n361), .a(n75) );
    inv_1 U355 ( .x(n175), .a(n353) );
    exnor2_3 U356 ( .x(SUM[29]), .a(n153), .b(n51) );
    nand4_4 U357 ( .x(n322), .a(n325), .b(n324), .c(n323), .d(n326) );
    oai211_3 U358 ( .x(n325), .a(n143), .b(n210), .c(n347), .d(n346) );
    ao21_3 U359 ( .x(n363), .a(n159), .b(n153), .c(n157) );
    nand2i_2 U36 ( .x(n330), .a(B[26]), .b(n221) );
    exnor2_3 U360 ( .x(SUM[30]), .a(n363), .b(n362) );
    inv_2 U361 ( .x(n362), .a(n173) );
    oai22_2 U362 ( .x(n171), .a(n155), .b(n260), .c(n151), .d(n259) );
    inv_0 U363 ( .x(n364), .a(n244) );
    aoi21_3 U364 ( .x(n155), .a(n156), .b(n153), .c(n157) );
    oaoi211_2 U365 ( .x(n76), .a(n78), .b(A[20]), .c(n322), .d(n77) );
    inv_2 U366 ( .x(n149), .a(n361) );
    inv_2 U37 ( .x(n221), .a(A[26]) );
    nand2_2 U38 ( .x(n331), .a(A[26]), .b(B[26]) );
    nand2i_2 U39 ( .x(n283), .a(n145), .b(A[25]) );
    nand2i_2 U40 ( .x(n282), .a(n145), .b(B[25]) );
    inv_2 U41 ( .x(n145), .a(n330) );
    nor2i_1 U42 ( .x(SUM[0]), .a(n354), .b(n355) );
    nand2_0 U43 ( .x(n133), .a(A[11]), .b(B[11]) );
    inv_5 U44 ( .x(n238), .a(n234) );
    inv_2 U45 ( .x(n251), .a(A[19]) );
    inv_0 U46 ( .x(n250), .a(B[19]) );
    nand2i_2 U47 ( .x(n276), .a(n131), .b(n242) );
    or3i_3 U48 ( .x(n237), .a(n238), .b(n102), .c(n230) );
    inv_5 U49 ( .x(n347), .a(n237) );
    nand2_2 U5 ( .x(n49), .a(n73), .b(n200) );
    nor3i_3 U50 ( .x(n143), .a(n144), .b(n115), .c(n141) );
    nand2_2 U51 ( .x(n195), .a(n287), .b(n315) );
    nand2_2 U52 ( .x(n317), .a(n195), .b(n233) );
    inv_0 U53 ( .x(n253), .a(B[13]) );
    inv_0 U54 ( .x(n316), .a(n127) );
    nand2_0 U55 ( .x(n127), .a(B[13]), .b(A[13]) );
    nand2i_2 U56 ( .x(n243), .a(n131), .b(n244) );
    inv_2 U57 ( .x(n115), .a(n301) );
    nand2_0 U58 ( .x(n130), .a(A[12]), .b(B[12]) );
    inv_2 U59 ( .x(n289), .a(n130) );
    inv_2 U6 ( .x(n146), .a(n49) );
    inv_2 U60 ( .x(n131), .a(n296) );
    nor2_1 U61 ( .x(n286), .a(n131), .b(n134) );
    aoi21_1 U62 ( .x(n287), .a(n286), .b(n288), .c(n289) );
    or2_2 U63 ( .x(n136), .a(n245), .b(n70) );
    inv_4 U64 ( .x(n97), .a(B[22]) );
    nand2i_2 U65 ( .x(n300), .a(A[22]), .b(n97) );
    exor2_1 U66 ( .x(n188), .a(A[19]), .b(B[19]) );
    inv_2 U67 ( .x(n290), .a(n266) );
    inv_0 U68 ( .x(n119), .a(n278) );
    nor2i_0 U69 ( .x(n117), .a(n267), .b(n228) );
    inv_10 U7 ( .x(n200), .a(A[1]) );
    aoi21_1 U70 ( .x(n116), .a(n117), .b(n118), .c(n119) );
    inv_0 U71 ( .x(n209), .a(A[3]) );
    nand2i_2 U72 ( .x(n267), .a(B[18]), .b(n249) );
    inv_7 U73 ( .x(n249), .a(A[18]) );
    inv_2 U74 ( .x(n235), .a(n267) );
    nor2i_1 U75 ( .x(n271), .a(A[18]), .b(n265) );
    nand2i_2 U77 ( .x(n159), .a(A[29]), .b(n218) );
    inv_2 U78 ( .x(n218), .a(B[29]) );
    nand2_2 U79 ( .x(n340), .a(B[27]), .b(A[27]) );
    inv_5 U8 ( .x(n73), .a(B[1]) );
    nand2i_2 U80 ( .x(n295), .a(A[8]), .b(n214) );
    nand2i_2 U81 ( .x(n152), .a(B[29]), .b(n217) );
    nand2_0 U82 ( .x(n284), .a(B[29]), .b(A[29]) );
    inv_2 U83 ( .x(n217), .a(A[29]) );
    nand2i_0 U84 ( .x(n297), .a(n74), .b(n200) );
    inv_2 U85 ( .x(n356), .a(n297) );
    nor2i_1 U86 ( .x(n357), .a(n358), .b(n356) );
    nand2_0 U87 ( .x(n86), .a(B[9]), .b(A[9]) );
    inv_0 U88 ( .x(n313), .a(n210) );
    nand2_2 U89 ( .x(n291), .a(n292), .b(n293) );
    inv_5 U90 ( .x(n213), .a(n55) );
    inv_4 U91 ( .x(n59), .a(n61) );
    inv_0 U92 ( .x(n68), .a(B[14]) );
    nand2i_2 U93 ( .x(n124), .a(n254), .b(n64) );
    oai21_1 U94 ( .x(n192), .a(n125), .b(n318), .c(n124) );
    nor2i_0 U95 ( .x(n120), .a(n121), .b(n122) );
    inv_3 U96 ( .x(n247), .a(B[16]) );
    inv_0 U98 ( .x(n223), .a(B[21]) );
    exor2_1 U99 ( .x(n184), .a(A[23]), .b(B[23]) );
endmodule


module EX_DW01_add_32_3_test_1 ( A, B, CI, SUM, CO );
input  [31:0] A;
input  [31:0] B;
output [31:0] SUM;
input  CI;
output CO;
    wire n327, n326, n294, n144, n145, n369, n146, n199, n85, n337, n115, n111, 
        n225, n162, n163, n164, n265, n340, n77, n127, n78, n91, n209, n165, 
        n169, n218, n354, n223, n353, n224, n161, n55, n160, n156, n159, n61, 
        n257, n256, n310, n166, n172, n190, n122, n187, n188, n189, n297, n141, 
        n323, n140, n200, n114, n118, n336, n64, n267, n261, n325, n58, n219, 
        n148, n66, n81, n149, n370, n73, n341, n71, n289, n285, n125, n288, 
        n201, n116, n139, n324, n331, n204, n158, n234, n105, n287, n126, n49, 
        n104, n298, n295, n296, n304, n203, n194, n279, n191, n192, n193, n196, 
        n197, n205, n135, n244, n368, n365, n195, n106, n335, n107, n108, n272, 
        n154, n151, n220, n142, n95, n215, n216, n212, n266, n69, n260, n211, 
        n346, n186, n147, n124, n155, n286, n207, n74, n80, n174, n320, n271, 
        n56, n299, n301, n332, n268, n292, n305, n167, n243, n117, n54, n53, 
        n50, n311, n312, n51, n52, n59, n60, n363, n362, n62, n314, n338, n258, 
        n255, n293, n306, n175, n70, n221, n157, n228, n303, n112, n232, n300, 
        n233, n57, n302, n309, n322, n177, n84, n246, n247, n349, n356, n98, 
        n97, n217, n96, n222, n308, n88, n227, n68, n230, n313, n343, n342, 
        n179, n182, n181, n237, n329, n86, n63, n290, n291, n339, n241, n242, 
        n273, n274, n67, n75, n173, n226, n121, n119, n307, n137, n138, n283, 
        n183, n150, n184, n185, n330, n238, n270, n269, n72, n282, n284, n176, 
        n264, n65, n348, n76, n79, n236, n344, n358, n210, n319, n345, n263, 
        n262, n153, n347, n90, n99, n132, n93, n92, n133, n134, n208, n231, 
        n152, n82, n83, n317, n316, n130, n87, n315, n249, n214, n239, n235, 
        n180, n109, n110, n170, n89, n202, n94, n253, n355, n254, n245, n100, 
        n101, n350, n102, n278, n103, n277, n248, n113, n321, n198, n371, n251, 
        n328, n352, n276, n131, n240, n360, n361, n250, n252, n275, n120, n229, 
        n123, n281, n333, n178, n366, n364, n136, n259, n171, n168, n367, n143, 
        n351, n318, n213, n357, n280, n128, n129, n359;
    inv_2 U100 ( .x(n327), .a(n326) );
    oai21_1 U101 ( .x(n294), .a(A[2]), .b(B[2]), .c(n326) );
    aoi21_1 U102 ( .x(n144), .a(n145), .b(n369), .c(n146) );
    exnor2_1 U103 ( .x(SUM[2]), .a(n144), .b(n294) );
    oai21_1 U104 ( .x(n199), .a(n85), .b(n337), .c(n115) );
    exor2_1 U105 ( .x(SUM[6]), .a(n199), .b(n111) );
    exor2_1 U106 ( .x(SUM[12]), .a(n225), .b(n162) );
    nor2i_1 U107 ( .x(n162), .a(n163), .b(n164) );
    inv_2 U108 ( .x(n164), .a(n265) );
    inv_4 U109 ( .x(n340), .a(n225) );
    nor2_0 U11 ( .x(n77), .a(n127), .b(n78) );
    exor2_1 U110 ( .x(SUM[27]), .a(n91), .b(n209) );
    exor2_1 U111 ( .x(n209), .a(B[27]), .b(A[27]) );
    exnor2_1 U112 ( .x(SUM[11]), .a(n165), .b(n169) );
    exor2_1 U113 ( .x(n218), .a(A[20]), .b(B[20]) );
    inv_2 U114 ( .x(n354), .a(n223) );
    inv_4 U115 ( .x(n353), .a(n224) );
    inv_5 U116 ( .x(n161), .a(n55) );
    oai21_1 U117 ( .x(n223), .a(n161), .b(n353), .c(n160) );
    exor2_1 U118 ( .x(SUM[14]), .a(n223), .b(n156) );
    exor2_1 U119 ( .x(SUM[13]), .a(n224), .b(n159) );
    aoi21_2 U12 ( .x(n61), .a(n257), .b(n256), .c(n310) );
    exor2_1 U120 ( .x(SUM[10]), .a(n166), .b(n172) );
    inv_2 U121 ( .x(n190), .a(n122) );
    aoi21_1 U122 ( .x(n187), .a(n188), .b(n189), .c(n190) );
    exnor2_1 U123 ( .x(n297), .a(A[22]), .b(B[22]) );
    inv_5 U124 ( .x(n141), .a(n323) );
    aoi21_1 U125 ( .x(n140), .a(A[22]), .b(B[22]), .c(n141) );
    mux2i_1 U126 ( .x(SUM[22]), .d0(n140), .sl(n187), .d1(n297) );
    exor2_1 U127 ( .x(SUM[5]), .a(n200), .b(n114) );
    oai21_1 U128 ( .x(n200), .a(n118), .b(n336), .c(n64) );
    nor2i_0 U129 ( .x(n114), .a(n115), .b(n85) );
    nand2i_3 U13 ( .x(n267), .a(B[14]), .b(n261) );
    inv_0 U130 ( .x(n325), .a(n58) );
    inv_2 U131 ( .x(n337), .a(n200) );
    exor2_1 U132 ( .x(n219), .a(A[19]), .b(B[19]) );
    nor2i_1 U133 ( .x(n148), .a(n66), .b(n81) );
    oai21_1 U134 ( .x(n149), .a(n370), .b(n73), .c(n341) );
    aoi21_1 U135 ( .x(n71), .a(n289), .b(n285), .c(n125) );
    inv_0 U136 ( .x(n288), .a(n149) );
    exor2_1 U137 ( .x(SUM[4]), .a(n201), .b(n116) );
    inv_2 U138 ( .x(n139), .a(n324) );
    inv_2 U139 ( .x(n331), .a(n204) );
    inv_5 U14 ( .x(n158), .a(n267) );
    nor2i_1 U140 ( .x(n116), .a(n64), .b(n118) );
    inv_2 U141 ( .x(n118), .a(n234) );
    inv_2 U142 ( .x(n336), .a(n201) );
    nand2i_2 U143 ( .x(n105), .a(n66), .b(n287) );
    inv_0 U144 ( .x(n66), .a(n310) );
    inv_7 U145 ( .x(n126), .a(A[18]) );
    oai21_1 U146 ( .x(n287), .a(n288), .b(n81), .c(n49) );
    mux2i_1 U147 ( .x(n104), .d0(n298), .sl(B[18]), .d1(n295) );
    nor2i_0 U148 ( .x(n298), .a(A[18]), .b(n287) );
    exnor2_1 U149 ( .x(n295), .a(n296), .b(n126) );
    nor2_2 U15 ( .x(n304), .a(n161), .b(n163) );
    inv_2 U150 ( .x(n296), .a(n287) );
    exor2_1 U151 ( .x(n203), .a(B[30]), .b(A[30]) );
    inv_2 U152 ( .x(n194), .a(n279) );
    aoi21_1 U153 ( .x(n191), .a(n192), .b(n193), .c(n194) );
    exnor2_1 U156 ( .x(SUM[8]), .a(n196), .b(n197) );
    exor2_1 U157 ( .x(n205), .a(B[29]), .b(A[29]) );
    inv_0 U158 ( .x(n135), .a(B[30]) );
    inv_2 U159 ( .x(n244), .a(A[29]) );
    inv_2 U16 ( .x(n261), .a(A[14]) );
    exnor2_1 U160 ( .x(SUM[1]), .a(n368), .b(n365) );
    exnor2_1 U161 ( .x(SUM[9]), .a(n195), .b(n106) );
    inv_2 U162 ( .x(n195), .a(n335) );
    nor2i_1 U163 ( .x(n106), .a(n107), .b(n108) );
    inv_0 U164 ( .x(n108), .a(n272) );
    exor2_1 U165 ( .x(SUM[16]), .a(n149), .b(n154) );
    exnor2_1 U166 ( .x(SUM[17]), .a(n151), .b(n220) );
    exnor2_1 U167 ( .x(SUM[21]), .a(n142), .b(n95) );
    exor2_1 U168 ( .x(SUM[23]), .a(n215), .b(n216) );
    exor2_1 U169 ( .x(n212), .a(B[25]), .b(A[25]) );
    nand2_2 U17 ( .x(n266), .a(n69), .b(n260) );
    exor2_1 U170 ( .x(n211), .a(A[26]), .b(B[26]) );
    inv_2 U171 ( .x(n346), .a(n186) );
    exnor2_1 U172 ( .x(SUM[19]), .a(n147), .b(n219) );
    nand2_2 U173 ( .x(SUM[18]), .a(n104), .b(n105) );
    oa21_1 U174 ( .x(n49), .a(n124), .b(n155), .c(n286) );
    nand2i_4 U175 ( .x(n289), .a(B[18]), .b(n126) );
    inv_4 U176 ( .x(n310), .a(n289) );
    exor2_1 U177 ( .x(n207), .a(A[28]), .b(B[28]) );
    inv_1 U178 ( .x(n74), .a(B[17]) );
    and4i_4 U179 ( .x(n80), .a(n174), .b(n320), .c(n271), .d(n272) );
    inv_4 U18 ( .x(n69), .a(A[13]) );
    oai211_2 U180 ( .x(n56), .a(n58), .b(n299), .c(n301), .d(n332) );
    or3i_4 U181 ( .x(n268), .a(n61), .b(n127), .c(n78) );
    nor2_3 U182 ( .x(n127), .a(A[17]), .b(B[17]) );
    nand4_1 U183 ( .x(n292), .a(n272), .b(n271), .c(n305), .d(n167) );
    nand2i_3 U184 ( .x(n272), .a(A[9]), .b(n243) );
    nand2_2 U185 ( .x(n117), .a(B[4]), .b(A[4]) );
    inv_0 U186 ( .x(n54), .a(n53) );
    nand2_0 U187 ( .x(n50), .a(n61), .b(n77) );
    aoai211_1 U188 ( .x(n311), .a(n54), .b(n256), .c(n71), .d(n312) );
    inv_0 U189 ( .x(n51), .a(n52) );
    inv_7 U190 ( .x(n59), .a(A[5]) );
    aoai211_4 U191 ( .x(n60), .a(n363), .b(n362), .c(n62), .d(n314) );
    nand2_5 U192 ( .x(n338), .a(n52), .b(n258) );
    inv_2 U193 ( .x(n255), .a(A[16]) );
    aoi31_3 U194 ( .x(n293), .a(n167), .b(n271), .c(n306), .d(n175) );
    and2_5 U195 ( .x(n175), .a(n271), .b(n70) );
    oai21_2 U196 ( .x(n221), .a(n158), .b(n354), .c(n157) );
    nor2i_1 U197 ( .x(n156), .a(n157), .b(n158) );
    inv_4 U198 ( .x(n228), .a(B[5]) );
    inv_0 U199 ( .x(n53), .a(n257) );
    nand2_2 U20 ( .x(n303), .a(A[0]), .b(B[0]) );
    nand2_1 U200 ( .x(n112), .a(A[6]), .b(B[6]) );
    nand4i_2 U201 ( .x(n232), .a(n58), .b(n300), .c(n234), .d(n233) );
    and2_3 U202 ( .x(n301), .a(n112), .b(n57) );
    inv_2 U203 ( .x(n57), .a(n302) );
    or3i_4 U204 ( .x(n309), .a(n322), .b(n177), .c(n158) );
    aoai211_5 U206 ( .x(n84), .a(n246), .b(n247), .c(n349), .d(n356) );
    oaoi211_4 U207 ( .x(n62), .a(n98), .b(n97), .c(n217), .d(n96) );
    exor2_1 U208 ( .x(n222), .a(n51), .b(B[15]) );
    nand2_0 U209 ( .x(n308), .a(A[15]), .b(B[15]) );
    aoi22_1 U21 ( .x(n233), .a(n88), .b(n227), .c(n68), .d(n230) );
    inv_2 U210 ( .x(n258), .a(B[15]) );
    nand4i_3 U212 ( .x(n217), .a(n311), .b(n313), .c(n343), .d(n342) );
    nor2_4 U213 ( .x(n313), .a(n179), .b(n182) );
    and4i_4 U214 ( .x(n179), .a(n181), .b(n237), .c(n329), .d(n86) );
    inv_2 U215 ( .x(n68), .a(B[3]) );
    inv_0 U216 ( .x(n63), .a(n117) );
    inv_2 U217 ( .x(n64), .a(n63) );
    nand3i_0 U218 ( .x(n290), .a(n291), .b(n292), .c(n293) );
    inv_2 U219 ( .x(n339), .a(n290) );
    inv_4 U22 ( .x(n88), .a(B[7]) );
    nand2i_0 U220 ( .x(n324), .a(B[3]), .b(n230) );
    nor2i_2 U221 ( .x(n305), .a(A[8]), .b(n241) );
    inv_0 U222 ( .x(n242), .a(A[8]) );
    nand2i_6 U223 ( .x(n181), .a(n273), .b(n274) );
    inv_0 U224 ( .x(n67), .a(n75) );
    aoai211_2 U225 ( .x(n285), .a(n74), .b(n75), .c(n155), .d(n286) );
    inv_2 U226 ( .x(n256), .a(B[19]) );
    inv_2 U227 ( .x(n70), .a(n173) );
    nand2i_5 U228 ( .x(n300), .a(B[6]), .b(n226) );
    exor2_1 U229 ( .x(n220), .a(n67), .b(B[17]) );
    nor2i_1 U23 ( .x(n121), .a(n122), .b(n119) );
    nor2_0 U230 ( .x(n124), .a(B[17]), .b(n67) );
    or3i_4 U231 ( .x(n307), .a(n304), .b(n158), .c(n177) );
    nor2i_0 U232 ( .x(n137), .a(n138), .b(n139) );
    oai21_1 U233 ( .x(n201), .a(n139), .b(n331), .c(n138) );
    nand3_2 U234 ( .x(n283), .a(n307), .b(n309), .c(n308) );
    nor2_3 U235 ( .x(n182), .a(n181), .b(n183) );
    inv_0 U236 ( .x(n150), .a(n71) );
    nor2i_0 U237 ( .x(n172), .a(n173), .b(n174) );
    aoi21_1 U238 ( .x(n147), .a(n148), .b(n149), .c(n150) );
    nor2_1 U239 ( .x(n184), .a(n185), .b(n186) );
    nand2i_0 U24 ( .x(n330), .a(A[2]), .b(n238) );
    oai22_1 U240 ( .x(n335), .a(n241), .b(n242), .c(n270), .d(n370) );
    oai21_3 U241 ( .x(n225), .a(n370), .b(n269), .c(n339) );
    inv_0 U242 ( .x(n72), .a(n273) );
    inv_2 U243 ( .x(n73), .a(n72) );
    or3i_4 U244 ( .x(n282), .a(n284), .b(n176), .c(n283) );
    nand2i_2 U245 ( .x(n284), .a(n264), .b(n65) );
    or3i_2 U247 ( .x(n348), .a(n60), .b(n185), .c(n76) );
    inv_0 U248 ( .x(n76), .a(B[25]) );
    inv_0 U249 ( .x(n341), .a(n282) );
    inv_0 U25 ( .x(n238), .a(B[2]) );
    and2_3 U250 ( .x(n78), .a(n79), .b(n255) );
    inv_2 U251 ( .x(n79), .a(B[16]) );
    inv_4 U252 ( .x(n236), .a(n329) );
    ao21_1 U253 ( .x(n204), .a(n329), .b(n330), .c(n327) );
    oai21_5 U254 ( .x(n329), .a(n146), .b(n303), .c(n369) );
    nand2i_2 U255 ( .x(n363), .a(n344), .b(n358) );
    nand3i_1 U256 ( .x(n210), .a(n346), .b(n319), .c(n345) );
    nand2_4 U258 ( .x(n107), .a(B[9]), .b(A[9]) );
    inv_0 U259 ( .x(n269), .a(n80) );
    nand2_0 U26 ( .x(n326), .a(A[2]), .b(B[2]) );
    inv_0 U260 ( .x(n270), .a(n320) );
    nand2i_4 U261 ( .x(n167), .a(A[10]), .b(n263) );
    nand2i_8 U262 ( .x(n271), .a(A[11]), .b(n262) );
    nor2i_1 U263 ( .x(n154), .a(n155), .b(n78) );
    inv_2 U264 ( .x(n153), .a(n155) );
    inv_2 U265 ( .x(n185), .a(n347) );
    ao21_6 U266 ( .x(n90), .a(A[30]), .b(n99), .c(n132) );
    inv_1 U267 ( .x(n93), .a(n92) );
    aoi21_3 U268 ( .x(n132), .a(n133), .b(n134), .c(n135) );
    inv_7 U269 ( .x(n349), .a(n208) );
    inv_2 U27 ( .x(n231), .a(B[1]) );
    nand2i_0 U270 ( .x(n81), .a(n127), .b(n152) );
    inv_0 U271 ( .x(n82), .a(n217) );
    inv_2 U272 ( .x(n83), .a(n82) );
    inv_0 U274 ( .x(n85), .a(n325) );
    aoi21_2 U275 ( .x(n317), .a(n60), .b(n316), .c(n184) );
    nand3i_3 U276 ( .x(n208), .a(n130), .b(n348), .c(n317) );
    nand2i_4 U277 ( .x(n183), .a(n87), .b(n56) );
    nand2i_2 U278 ( .x(n315), .a(B[24]), .b(n249) );
    exor2_1 U279 ( .x(n214), .a(A[24]), .b(B[24]) );
    nand2_0 U28 ( .x(n145), .a(B[0]), .b(A[0]) );
    exor2_1 U280 ( .x(SUM[20]), .a(n83), .b(n218) );
    nand2i_4 U281 ( .x(n239), .a(n238), .b(n237) );
    nand2i_4 U282 ( .x(n235), .a(n236), .b(n237) );
    inv_5 U283 ( .x(n241), .a(B[8]) );
    ao21_1 U284 ( .x(n197), .a(A[8]), .b(B[8]), .c(n270) );
    inv_2 U286 ( .x(n86), .a(n180) );
    nor2_0 U287 ( .x(n180), .a(A[2]), .b(B[2]) );
    inv_3 U288 ( .x(n243), .a(B[9]) );
    nor2i_0 U289 ( .x(n109), .a(n110), .b(n87) );
    nand2_0 U29 ( .x(n170), .a(A[11]), .b(B[11]) );
    exnor2_5 U290 ( .x(SUM[31]), .a(n90), .b(n89) );
    inv_2 U291 ( .x(n89), .a(n202) );
    exor2_1 U292 ( .x(n202), .a(B[31]), .b(A[31]) );
    nand3i_0 U293 ( .x(n91), .a(n130), .b(n348), .c(n317) );
    inv_0 U294 ( .x(n92), .a(n60) );
    inv_0 U295 ( .x(n94), .a(n62) );
    inv_2 U296 ( .x(n95), .a(n94) );
    inv_0 U297 ( .x(n189), .a(n95) );
    inv_2 U298 ( .x(n98), .a(n253) );
    nand2_0 U299 ( .x(n355), .a(A[20]), .b(B[20]) );
    nand2_2 U30 ( .x(n110), .a(A[7]), .b(B[7]) );
    inv_0 U300 ( .x(n254), .a(A[20]) );
    inv_0 U301 ( .x(n253), .a(B[20]) );
    nand2_2 U302 ( .x(n122), .a(B[21]), .b(A[21]) );
    aoai211_1 U303 ( .x(n99), .a(n244), .b(n245), .c(n100), .d(n279) );
    nand2_1 U304 ( .x(n155), .a(A[16]), .b(B[16]) );
    nand2_0 U306 ( .x(n157), .a(A[14]), .b(B[14]) );
    and3i_1 U307 ( .x(n176), .a(n177), .b(B[14]), .c(A[14]) );
    inv_2 U308 ( .x(n193), .a(n100) );
    inv_2 U309 ( .x(n101), .a(n350) );
    inv_3 U31 ( .x(n227), .a(A[7]) );
    inv_2 U310 ( .x(n102), .a(n278) );
    inv_2 U311 ( .x(n103), .a(n277) );
    nand2_0 U312 ( .x(n350), .a(B[28]), .b(A[28]) );
    inv_0 U313 ( .x(n278), .a(B[28]) );
    inv_0 U314 ( .x(n277), .a(A[28]) );
    nand2_2 U316 ( .x(n163), .a(A[12]), .b(B[12]) );
    exor2_1 U317 ( .x(SUM[25]), .a(n93), .b(n212) );
    nand2_0 U318 ( .x(n319), .a(B[25]), .b(n93) );
    nand2_0 U319 ( .x(n345), .a(A[25]), .b(n93) );
    nand2i_2 U32 ( .x(n347), .a(B[26]), .b(n248) );
    nor2i_0 U320 ( .x(n111), .a(n112), .b(n113) );
    inv_0 U321 ( .x(n321), .a(n112) );
    nand2_1 U322 ( .x(n173), .a(B[10]), .b(A[10]) );
    inv_6 U323 ( .x(n263), .a(B[10]) );
    exor2_3 U324 ( .x(SUM[7]), .a(n198), .b(n109) );
    exnor2_3 U325 ( .x(SUM[30]), .a(n191), .b(n203) );
    exnor2_3 U326 ( .x(SUM[28]), .a(n371), .b(n207) );
    exor2_3 U327 ( .x(SUM[26]), .a(n210), .b(n211) );
    exor2_3 U328 ( .x(SUM[15]), .a(n221), .b(n222) );
    inv_6 U329 ( .x(n251), .a(B[23]) );
    inv_2 U33 ( .x(n248), .a(A[26]) );
    inv_6 U330 ( .x(n134), .a(A[30]) );
    nand3i_3 U331 ( .x(n299), .a(n138), .b(n300), .c(n234) );
    nand2i_4 U332 ( .x(n328), .a(A[1]), .b(n231) );
    inv_5 U333 ( .x(n146), .a(n328) );
    ao211_5 U334 ( .x(n332), .a(n117), .b(n115), .c(n58), .d(n113) );
    ao21_4 U335 ( .x(n198), .a(n199), .b(n300), .c(n321) );
    nand2_2 U336 ( .x(n352), .a(A[22]), .b(B[22]) );
    oai21_4 U337 ( .x(n224), .a(n340), .b(n164), .c(n163) );
    inv_5 U338 ( .x(n358), .a(n276) );
    nand2i_4 U339 ( .x(n342), .a(n50), .b(n282) );
    nor2i_1 U34 ( .x(n130), .a(A[26]), .b(n131) );
    nand3i_5 U340 ( .x(n343), .a(n240), .b(n360), .c(n361) );
    nand2i_6 U341 ( .x(n188), .a(A[21]), .b(n250) );
    or3i_5 U342 ( .x(n276), .a(n188), .b(n252), .c(n141) );
    or3i_5 U343 ( .x(n275), .a(n188), .b(n251), .c(n141) );
    inv_6 U344 ( .x(n113), .a(n300) );
    nand2i_6 U345 ( .x(n323), .a(A[22]), .b(n120) );
    nor2i_5 U346 ( .x(n316), .a(A[25]), .b(n185) );
    inv_10 U347 ( .x(n246), .a(A[27]) );
    inv_10 U348 ( .x(n247), .a(B[27]) );
    nand2_4 U349 ( .x(n356), .a(B[27]), .b(A[27]) );
    inv_2 U35 ( .x(n131), .a(B[26]) );
    nand2i_6 U350 ( .x(n234), .a(A[4]), .b(n229) );
    inv_10 U351 ( .x(n262), .a(B[11]) );
    inv_6 U352 ( .x(n177), .a(n338) );
    inv_14 U353 ( .x(n120), .a(B[22]) );
    nor2_8 U354 ( .x(n123), .a(A[23]), .b(B[23]) );
    nand2_4 U355 ( .x(n281), .a(A[23]), .b(B[23]) );
    inv_10 U356 ( .x(n229), .a(B[4]) );
    nor2i_8 U357 ( .x(n119), .a(A[22]), .b(n120) );
    oa222_4 U358 ( .x(n370), .a(n239), .b(n240), .c(n87), .d(n333), .e(n178), 
        .f(n235) );
    inv_0 U359 ( .x(n196), .a(n370) );
    nor2i_1 U36 ( .x(SUM[0]), .a(n365), .b(n366) );
    inv_3 U360 ( .x(n333), .a(n56) );
    inv_0 U361 ( .x(n240), .a(A[2]) );
    aoi221_4 U362 ( .x(n100), .a(n103), .b(n364), .c(n84), .d(n102), .e(n101)
         );
    aoai211_4 U363 ( .x(n364), .a(n246), .b(n247), .c(n349), .d(n356) );
    inv_5 U364 ( .x(n133), .a(n136) );
    aoai211_4 U365 ( .x(n136), .a(n244), .b(n245), .c(n100), .d(n279) );
    inv_3 U366 ( .x(n361), .a(n181) );
    exnor2_2 U367 ( .x(SUM[29]), .a(n100), .b(n205) );
    inv_2 U368 ( .x(n371), .a(n364) );
    nand4_3 U369 ( .x(n264), .a(n338), .b(n265), .c(n266), .d(n267) );
    nor2_1 U37 ( .x(n366), .a(B[0]), .b(A[0]) );
    nand2i_4 U370 ( .x(n265), .a(B[12]), .b(n259) );
    nand2i_4 U371 ( .x(n273), .a(n264), .b(n80) );
    inv_4 U372 ( .x(n260), .a(B[13]) );
    inv_2 U38 ( .x(n291), .a(n170) );
    inv_2 U39 ( .x(n171), .a(n271) );
    nor2i_1 U40 ( .x(n169), .a(n170), .b(n171) );
    aoi21_1 U41 ( .x(n165), .a(n166), .b(n167), .c(n168) );
    inv_4 U42 ( .x(n274), .a(n268) );
    inv_5 U43 ( .x(n257), .a(A[19]) );
    nand2_0 U44 ( .x(n312), .a(A[19]), .b(B[19]) );
    nor2i_1 U45 ( .x(n159), .a(n160), .b(n161) );
    nand2_1 U46 ( .x(n160), .a(B[13]), .b(A[13]) );
    nand2_2 U47 ( .x(n55), .a(n69), .b(n260) );
    inv_2 U48 ( .x(n322), .a(n160) );
    inv_2 U49 ( .x(n259), .a(A[12]) );
    nand2i_4 U5 ( .x(n320), .a(A[8]), .b(n241) );
    inv_0 U50 ( .x(n168), .a(n173) );
    oai21_1 U51 ( .x(n166), .a(n195), .b(n108), .c(n107) );
    nand2_1 U52 ( .x(n115), .a(B[5]), .b(A[5]) );
    and2_1 U53 ( .x(n125), .a(B[18]), .b(A[18]) );
    inv_5 U54 ( .x(n75), .a(A[17]) );
    inv_2 U55 ( .x(n174), .a(n167) );
    inv_2 U56 ( .x(n230), .a(A[3]) );
    nand2_2 U57 ( .x(n138), .a(A[3]), .b(B[3]) );
    nand2_2 U58 ( .x(n286), .a(A[17]), .b(B[17]) );
    nand2i_2 U59 ( .x(n192), .a(A[29]), .b(n245) );
    inv_5 U6 ( .x(n226), .a(A[6]) );
    and2_6 U60 ( .x(n58), .a(n59), .b(n228) );
    inv_2 U61 ( .x(n302), .a(n110) );
    inv_5 U62 ( .x(n237), .a(n232) );
    nor2_0 U63 ( .x(n178), .a(A[2]), .b(B[2]) );
    and2_1 U64 ( .x(n87), .a(n88), .b(n227) );
    inv_5 U65 ( .x(n360), .a(n239) );
    inv_2 U66 ( .x(n245), .a(B[29]) );
    nand2_2 U68 ( .x(n279), .a(B[29]), .b(A[29]) );
    nand2_0 U69 ( .x(n365), .a(A[0]), .b(B[0]) );
    nand3i_2 U7 ( .x(n65), .a(n291), .b(n292), .c(n293) );
    nor2_1 U70 ( .x(n367), .a(B[1]), .b(A[1]) );
    nand2_2 U71 ( .x(n369), .a(B[1]), .b(A[1]) );
    nor2i_1 U72 ( .x(n368), .a(n369), .b(n367) );
    inv_2 U73 ( .x(n306), .a(n107) );
    inv_2 U75 ( .x(n152), .a(n78) );
    aoi21_1 U76 ( .x(n151), .a(n152), .b(n149), .c(n153) );
    inv_0 U77 ( .x(n250), .a(B[21]) );
    inv_2 U78 ( .x(n143), .a(n188) );
    nor2i_1 U79 ( .x(n142), .a(n122), .b(n143) );
    inv_10 U8 ( .x(n52), .a(A[15]) );
    exor2_1 U80 ( .x(n216), .a(A[23]), .b(B[23]) );
    nand2i_0 U81 ( .x(n351), .a(n141), .b(n190) );
    nand2i_2 U82 ( .x(n318), .a(n141), .b(n188) );
    oai211_1 U83 ( .x(n215), .a(n95), .b(n318), .c(n352), .d(n351) );
    exor2_1 U84 ( .x(SUM[24]), .a(n213), .b(n214) );
    aoai211_1 U85 ( .x(n213), .a(n276), .b(n275), .c(n95), .d(n357) );
    aoi21_1 U86 ( .x(n314), .a(n280), .b(n315), .c(n128) );
    oai31_1 U87 ( .x(n280), .a(n121), .b(n141), .c(n123), .d(n281) );
    nor2i_1 U88 ( .x(n128), .a(A[24]), .b(n129) );
    inv_2 U89 ( .x(n129), .a(B[24]) );
    inv_2 U90 ( .x(n357), .a(n280) );
    inv_2 U91 ( .x(n96), .a(n355) );
    inv_2 U92 ( .x(n97), .a(n254) );
    nand2i_2 U93 ( .x(n362), .a(n344), .b(n359) );
    inv_2 U94 ( .x(n359), .a(n275) );
    inv_2 U95 ( .x(n344), .a(n315) );
    inv_2 U96 ( .x(n249), .a(A[24]) );
    inv_2 U97 ( .x(n252), .a(A[23]) );
    nand2_2 U98 ( .x(n186), .a(A[25]), .b(B[25]) );
    exor2_1 U99 ( .x(SUM[3]), .a(n204), .b(n137) );
endmodule


module EX_DW01_add_32_7_test_1 ( A, B, CI, SUM, CO );
input  [31:0] A;
input  [31:0] B;
output [31:0] SUM;
input  CI;
output CO;
    wire n60, n331, n267, n190, n245, n138, n333, n322, n330, n295, n242, n268, 
        n246, n336, n184, n55, n203, n134, n309, n308, n135, n136, n306, n313, 
        n139, n277, n200, n107, n50, n157, n158, n159, n121, n251, n207, n160, 
        n164, n163, n168, n165, n166, n215, n95, n89, n220, n151, n221, n154, 
        n161, n167, n323, n241, n49, n103, n102, n169, n162, n191, n118, n280, 
        n137, n201, n109, n142, n216, n114, n229, n112, n113, n202, n100, n276, 
        n273, n204, n205, n197, n198, n235, n106, n305, n132, n81, n131, n130, 
        n133, n239, n101, n252, n59, n218, n153, n326, n152, n219, n145, n217, 
        n301, n69, n98, n214, n94, n327, n247, n185, n213, n210, n211, n209, 
        n269, n299, n228, n208, n54, n88, n129, n293, n82, n236, n237, n253, 
        n316, n329, n255, n73, n86, n225, n51, n174, n258, n75, n259, n52, n53, 
        n248, n291, n156, n155, n307, n223, n110, n97, n314, n111, n176, n177, 
        n178, n143, n249, n340, n275, n337, n85, n310, n226, n79, n335, n230, 
        n318, n144, n146, n147, n148, n92, n338, n339, n186, n188, n192, n193, 
        n194, n187, n93, n63, n70, n250, n319, n224, n56, n170, n62, n321, 
        n288, n179, n122, n181, n286, n71, n303, n254, n289, n105, n173, n74, 
        n58, n264, n65, n61, n57, n64, n270, n272, n195, n282, n66, n123, n68, 
        n206, n175, n292, n284, n271, n76, n261, n78, n80, n141, n120, n83, 
        n119, n302, n149, n260, n265, n84, n87, n256, n117, n115, n231, n287, 
        n234, n212, n90, n324, n334, n91, n116, n96, n222, n104, n172, n180, 
        n182, n183, n199, n240, n278, n279, n108, n285, n290, n312, n233, n298, 
        n296, n126, n300, n297, n311, n315, n317, n328, n320, n257, n99, n281, 
        n77, n232, n227, n332, n294, n342, n341, n343, n140, n344, n262, n238, 
        n67, n283, n266, n263, n128, n171, n127, n72, n325, n150, n304, n244, 
        n243, n125, n124;
    inv_2 U10 ( .x(n60), .a(B[14]) );
    inv_2 U100 ( .x(n331), .a(n267) );
    or3i_2 U101 ( .x(n267), .a(n190), .b(n245), .c(n138) );
    inv_2 U102 ( .x(n245), .a(B[23]) );
    nand2i_2 U103 ( .x(n333), .a(n322), .b(n330) );
    inv_2 U104 ( .x(n322), .a(n295) );
    nand2i_0 U105 ( .x(n295), .a(B[24]), .b(n242) );
    inv_2 U106 ( .x(n242), .a(A[24]) );
    inv_2 U107 ( .x(n330), .a(n268) );
    or3i_2 U108 ( .x(n268), .a(n190), .b(n246), .c(n138) );
    inv_2 U109 ( .x(n246), .a(A[23]) );
    nor2_0 U11 ( .x(n336), .a(B[0]), .b(A[0]) );
    nand2_2 U110 ( .x(n184), .a(n55), .b(B[25]) );
    exor2_1 U111 ( .x(SUM[3]), .a(n203), .b(n134) );
    inv_2 U112 ( .x(n309), .a(n308) );
    nor2i_1 U113 ( .x(n134), .a(n135), .b(n136) );
    inv_2 U114 ( .x(n136), .a(n306) );
    inv_2 U115 ( .x(n313), .a(n203) );
    exnor2_1 U116 ( .x(SUM[2]), .a(n139), .b(n277) );
    exor2_1 U117 ( .x(SUM[6]), .a(n200), .b(n107) );
    exnor2_1 U118 ( .x(SUM[12]), .a(n50), .b(n157) );
    nor2i_0 U119 ( .x(n157), .a(n158), .b(n159) );
    nor2_1 U12 ( .x(n121), .a(A[17]), .b(B[17]) );
    inv_0 U120 ( .x(n159), .a(n251) );
    exor2_1 U121 ( .x(n207), .a(B[27]), .b(A[27]) );
    exnor2_1 U122 ( .x(SUM[11]), .a(n160), .b(n164) );
    inv_2 U123 ( .x(n163), .a(n168) );
    nor2i_1 U124 ( .x(n164), .a(n165), .b(n166) );
    exor2_1 U125 ( .x(n215), .a(n95), .b(B[20]) );
    exnor2_1 U126 ( .x(SUM[20]), .a(n89), .b(n215) );
    exor2_1 U127 ( .x(SUM[14]), .a(n220), .b(n151) );
    exor2_1 U128 ( .x(SUM[13]), .a(n221), .b(n154) );
    exor2_1 U129 ( .x(SUM[10]), .a(n161), .b(n167) );
    nand2i_2 U13 ( .x(n323), .a(B[26]), .b(n241) );
    oai21_1 U130 ( .x(n161), .a(n49), .b(n103), .c(n102) );
    nor2i_1 U131 ( .x(n167), .a(n168), .b(n169) );
    inv_0 U132 ( .x(n169), .a(n162) );
    inv_2 U133 ( .x(n191), .a(n118) );
    exnor2_1 U134 ( .x(n280), .a(A[22]), .b(B[22]) );
    aoi21_1 U135 ( .x(n137), .a(A[22]), .b(B[22]), .c(n138) );
    exor2_1 U137 ( .x(SUM[5]), .a(n201), .b(n109) );
    exnor2_1 U138 ( .x(SUM[19]), .a(n142), .b(n216) );
    exor2_1 U139 ( .x(n216), .a(A[19]), .b(B[19]) );
    inv_2 U14 ( .x(n241), .a(A[26]) );
    inv_2 U140 ( .x(n114), .a(n229) );
    nor2i_1 U141 ( .x(n112), .a(n113), .b(n114) );
    exor2_1 U142 ( .x(SUM[4]), .a(n202), .b(n112) );
    nand2i_0 U143 ( .x(n100), .a(n276), .b(n273) );
    exnor2_1 U144 ( .x(SUM[28]), .a(n204), .b(n205) );
    exnor2_1 U145 ( .x(SUM[8]), .a(n197), .b(n198) );
    inv_5 U146 ( .x(n235), .a(A[2]) );
    inv_5 U147 ( .x(n106), .a(n305) );
    inv_0 U149 ( .x(n132), .a(B[30]) );
    and2_3 U15 ( .x(n81), .a(A[0]), .b(B[0]) );
    inv_2 U150 ( .x(n131), .a(A[30]) );
    inv_5 U151 ( .x(n130), .a(n133) );
    inv_2 U152 ( .x(n239), .a(A[29]) );
    nor2i_1 U153 ( .x(n101), .a(n102), .b(n103) );
    exnor2_1 U154 ( .x(SUM[9]), .a(n49), .b(n101) );
    inv_5 U155 ( .x(n252), .a(n59) );
    oai21_1 U156 ( .x(n218), .a(n153), .b(n326), .c(n152) );
    exor2_2 U157 ( .x(SUM[15]), .a(n218), .b(n219) );
    exnor2_1 U158 ( .x(SUM[17]), .a(n145), .b(n217) );
    inv_2 U159 ( .x(n301), .a(n190) );
    nor2i_3 U16 ( .x(n69), .a(n98), .b(A[6]) );
    nand2i_2 U160 ( .x(n214), .a(n301), .b(n118) );
    inv_2 U161 ( .x(n94), .a(n327) );
    inv_1 U162 ( .x(n247), .a(B[20]) );
    exnor2_1 U163 ( .x(SUM[23]), .a(n185), .b(n213) );
    exor2_1 U164 ( .x(n213), .a(A[23]), .b(B[23]) );
    exnor2_1 U165 ( .x(SUM[25]), .a(n210), .b(n211) );
    exor2_1 U166 ( .x(n211), .a(B[25]), .b(n55) );
    exor2_1 U167 ( .x(n209), .a(A[26]), .b(B[26]) );
    inv_2 U168 ( .x(n269), .a(B[25]) );
    inv_5 U169 ( .x(n210), .a(n299) );
    nor2_2 U17 ( .x(n228), .a(n106), .b(n136) );
    oai221_1 U170 ( .x(n208), .a(n210), .b(n269), .c(n210), .d(n54), .e(n184)
         );
    exor2_1 U171 ( .x(SUM[26]), .a(n208), .b(n209) );
    ao21_2 U173 ( .x(n88), .a(n133), .b(A[30]), .c(n129) );
    inv_2 U174 ( .x(n293), .a(n82) );
    oa22_1 U175 ( .x(n49), .a(n236), .b(n237), .c(n253), .d(n316) );
    aoi22_1 U176 ( .x(n50), .a(n329), .b(n255), .c(n197), .d(n73) );
    inv_2 U177 ( .x(n55), .a(n54) );
    inv_2 U178 ( .x(n54), .a(A[25]) );
    inv_1 U179 ( .x(n86), .a(B[19]) );
    nand2i_2 U18 ( .x(n306), .a(B[3]), .b(n225) );
    exnor2_1 U180 ( .x(n51), .a(B[31]), .b(A[31]) );
    inv_2 U181 ( .x(n174), .a(n258) );
    nand2i_2 U182 ( .x(n258), .a(n75), .b(n259) );
    exnor2_1 U183 ( .x(n52), .a(B[30]), .b(A[30]) );
    exnor2_1 U184 ( .x(n53), .a(B[29]), .b(A[29]) );
    exor2_1 U186 ( .x(n205), .a(A[28]), .b(B[28]) );
    inv_2 U187 ( .x(n95), .a(n248) );
    oai211_2 U188 ( .x(n291), .a(n156), .b(n158), .c(n155), .d(n152) );
    nand2_2 U189 ( .x(n158), .a(A[12]), .b(B[12]) );
    inv_2 U19 ( .x(n225), .a(A[3]) );
    nand2i_2 U190 ( .x(n307), .a(A[5]), .b(n223) );
    nand2_1 U191 ( .x(n110), .a(B[5]), .b(A[5]) );
    nor2i_5 U192 ( .x(n97), .a(A[6]), .b(n98) );
    ao211_5 U193 ( .x(n314), .a(n113), .b(n110), .c(n111), .d(n69) );
    nor2_6 U194 ( .x(n176), .a(n177), .b(n178) );
    nor2i_0 U195 ( .x(n143), .a(n276), .b(n249) );
    oai21_1 U196 ( .x(n273), .a(n340), .b(n249), .c(n275) );
    nor2_0 U197 ( .x(n337), .a(n85), .b(A[1]) );
    nand2i_2 U198 ( .x(n310), .a(A[1]), .b(n226) );
    inv_2 U199 ( .x(n79), .a(A[1]) );
    nand2_2 U20 ( .x(n335), .a(A[0]), .b(B[0]) );
    nand2_3 U200 ( .x(n135), .a(A[3]), .b(B[3]) );
    nor2_2 U201 ( .x(n230), .a(n111), .b(n69) );
    oai21_2 U202 ( .x(n200), .a(n111), .b(n318), .c(n110) );
    inv_8 U203 ( .x(n111), .a(n307) );
    aoi21_1 U204 ( .x(n142), .a(n143), .b(n144), .c(n82) );
    aoi21_1 U205 ( .x(n145), .a(n146), .b(n144), .c(n147) );
    exor2_1 U206 ( .x(SUM[16]), .a(n144), .b(n148) );
    exnor2_1 U208 ( .x(SUM[21]), .a(n92), .b(n214) );
    nor2i_1 U21 ( .x(n338), .a(n339), .b(n337) );
    aoi21_1 U210 ( .x(n185), .a(n186), .b(n92), .c(n188) );
    aoi21_1 U211 ( .x(n192), .a(n193), .b(n92), .c(n194) );
    inv_0 U212 ( .x(n187), .a(n93) );
    ao23_3 U214 ( .x(n63), .a(B[15]), .b(A[15]), .c(n291), .d(n252), .e(n70)
         );
    nand4_1 U215 ( .x(n250), .a(n252), .b(n319), .c(n251), .d(n70) );
    nand2_2 U216 ( .x(n113), .a(B[4]), .b(A[4]) );
    nand2i_2 U217 ( .x(n229), .a(A[4]), .b(n224) );
    inv_2 U218 ( .x(n223), .a(B[5]) );
    inv_2 U219 ( .x(n56), .a(n170) );
    inv_2 U22 ( .x(n62), .a(n166) );
    oai222_4 U220 ( .x(n321), .a(n235), .b(n288), .c(n179), .d(n122), .e(n181), 
        .f(n286) );
    exor2_1 U221 ( .x(n219), .a(A[15]), .b(B[15]) );
    inv_5 U222 ( .x(n71), .a(B[15]) );
    and4_5 U223 ( .x(n73), .a(n303), .b(n254), .c(n162), .d(n255) );
    nand2_2 U224 ( .x(n165), .a(A[11]), .b(B[11]) );
    nand2i_2 U225 ( .x(n303), .a(A[8]), .b(n236) );
    inv_0 U226 ( .x(n237), .a(A[8]) );
    ao21_1 U227 ( .x(n198), .a(A[8]), .b(B[8]), .c(n253) );
    nand2_1 U228 ( .x(n289), .a(A[8]), .b(B[8]) );
    nand2_1 U229 ( .x(n105), .a(A[7]), .b(B[7]) );
    inv_5 U23 ( .x(n173), .a(n74) );
    and4i_2 U231 ( .x(n58), .a(n59), .b(n319), .c(n251), .d(n70) );
    nand2i_2 U232 ( .x(n251), .a(B[12]), .b(n264) );
    inv_2 U233 ( .x(n65), .a(A[6]) );
    exnor2_3 U234 ( .x(SUM[30]), .a(n61), .b(n52) );
    oai21_1 U235 ( .x(n61), .a(n57), .b(n64), .c(n270) );
    ao31_6 U236 ( .x(n272), .a(n329), .b(n62), .c(n58), .d(n63) );
    inv_2 U237 ( .x(n64), .a(n195) );
    ao221_3 U238 ( .x(n282), .a(n98), .b(n65), .c(n66), .d(n224), .e(n135) );
    inv_5 U239 ( .x(n224), .a(B[4]) );
    nor2i_1 U24 ( .x(n123), .a(A[19]), .b(n86) );
    inv_10 U240 ( .x(n68), .a(A[13]) );
    inv_0 U241 ( .x(n253), .a(n303) );
    inv_2 U242 ( .x(n166), .a(n255) );
    exor2_1 U243 ( .x(SUM[27]), .a(n206), .b(n207) );
    nand2_5 U246 ( .x(n74), .a(n174), .b(n272) );
    inv_0 U247 ( .x(n175), .a(n272) );
    oai211_4 U248 ( .x(n292), .a(n282), .b(n111), .c(n284), .d(n314) );
    inv_0 U249 ( .x(n276), .a(n75) );
    nand2_2 U25 ( .x(n271), .a(A[23]), .b(B[23]) );
    inv_5 U250 ( .x(n76), .a(B[18]) );
    inv_16 U251 ( .x(n261), .a(A[18]) );
    inv_0 U253 ( .x(n339), .a(n78) );
    inv_6 U254 ( .x(n80), .a(B[1]) );
    inv_0 U255 ( .x(n141), .a(n310) );
    nand2_4 U256 ( .x(n102), .a(A[9]), .b(B[9]) );
    nor2_0 U257 ( .x(n120), .a(B[17]), .b(A[17]) );
    oaoi211_2 U258 ( .x(n82), .a(n83), .b(n261), .c(n275), .d(n75) );
    inv_0 U259 ( .x(n83), .a(B[18]) );
    nor2_1 U26 ( .x(n119), .a(A[23]), .b(B[23]) );
    ao21_3 U260 ( .x(n275), .a(n302), .b(n149), .c(n120) );
    inv_2 U261 ( .x(n260), .a(A[16]) );
    nand2_0 U262 ( .x(n302), .a(A[17]), .b(B[17]) );
    inv_2 U264 ( .x(n265), .a(A[10]) );
    inv_0 U265 ( .x(n84), .a(B[1]) );
    inv_2 U266 ( .x(n85), .a(n84) );
    ao211_5 U267 ( .x(n177), .a(n87), .b(n86), .c(n258), .d(n256) );
    inv_2 U268 ( .x(n87), .a(A[19]) );
    exnor2_3 U269 ( .x(SUM[31]), .a(n88), .b(n51) );
    nor2i_1 U27 ( .x(n117), .a(n118), .b(n115) );
    oa222_1 U270 ( .x(n89), .a(n235), .b(n288), .c(n179), .d(n122), .e(n181), 
        .f(n286) );
    nand2i_5 U271 ( .x(n286), .a(n231), .b(n287) );
    nand2i_4 U272 ( .x(n288), .a(n234), .b(n287) );
    exor2_1 U273 ( .x(n212), .a(A[24]), .b(B[24]) );
    exor2_1 U274 ( .x(n217), .a(A[17]), .b(B[17]) );
    inv_2 U275 ( .x(n90), .a(n324) );
    inv_0 U276 ( .x(n204), .a(n334) );
    nand2_0 U277 ( .x(n324), .a(B[28]), .b(A[28]) );
    inv_2 U278 ( .x(n91), .a(n187) );
    inv_4 U279 ( .x(n92), .a(n91) );
    nor2i_1 U28 ( .x(n115), .a(A[22]), .b(n116) );
    inv_2 U280 ( .x(n96), .a(n247) );
    nand2_0 U281 ( .x(n327), .a(A[20]), .b(B[20]) );
    inv_0 U282 ( .x(n248), .a(A[20]) );
    nand2_3 U283 ( .x(n118), .a(B[21]), .b(A[21]) );
    aoi21_1 U284 ( .x(n160), .a(n161), .b(n162), .c(n163) );
    nand2i_3 U285 ( .x(n162), .a(B[10]), .b(n265) );
    nand2i_2 U286 ( .x(n305), .a(B[7]), .b(n222) );
    nand2_2 U287 ( .x(n168), .a(A[10]), .b(B[10]) );
    nor2i_5 U288 ( .x(n104), .a(n105), .b(n106) );
    nor2_5 U289 ( .x(n172), .a(A[2]), .b(B[2]) );
    inv_2 U29 ( .x(n116), .a(B[22]) );
    nor3_5 U290 ( .x(n179), .a(n176), .b(n173), .c(n180) );
    nor2_5 U291 ( .x(n181), .a(A[2]), .b(B[2]) );
    nor2_5 U292 ( .x(n182), .a(n183), .b(n184) );
    exor2_3 U293 ( .x(SUM[7]), .a(n199), .b(n104) );
    exnor2_3 U294 ( .x(SUM[24]), .a(n192), .b(n212) );
    inv_6 U295 ( .x(n240), .a(B[29]) );
    inv_6 U296 ( .x(n264), .a(A[12]) );
    exnor2_3 U297 ( .x(n278), .a(n279), .b(n261) );
    nor2i_5 U298 ( .x(n284), .a(n108), .b(n285) );
    nand2_2 U299 ( .x(n290), .a(n165), .b(n168) );
    nand2i_2 U30 ( .x(n312), .a(A[2]), .b(n233) );
    nand2i_4 U300 ( .x(n180), .a(n123), .b(n293) );
    aoi21_3 U301 ( .x(n298), .a(n296), .b(n299), .c(n126) );
    aoi21_3 U302 ( .x(n300), .a(n297), .b(n299), .c(n182) );
    nand2_5 U303 ( .x(n308), .a(A[2]), .b(B[2]) );
    ao21_4 U304 ( .x(n203), .a(n311), .b(n312), .c(n309) );
    oai222_4 U305 ( .x(n197), .a(n234), .b(n235), .c(n106), .d(n315), .e(n172), 
        .f(n231) );
    oai21_4 U306 ( .x(n202), .a(n136), .b(n313), .c(n135) );
    inv_5 U307 ( .x(n317), .a(n202) );
    oai21_4 U308 ( .x(n201), .a(n114), .b(n317), .c(n113) );
    inv_5 U309 ( .x(n318), .a(n201) );
    oai21_1 U31 ( .x(n277), .a(A[2]), .b(B[2]), .c(n308) );
    nand2_2 U310 ( .x(n193), .a(n268), .b(n267) );
    nand2_5 U311 ( .x(n270), .a(B[29]), .b(A[29]) );
    nand2i_4 U312 ( .x(n328), .a(n102), .b(n162) );
    nand3i_3 U313 ( .x(n329), .a(n290), .b(n328), .c(n320) );
    inv_5 U314 ( .x(n257), .a(n250) );
    mux2i_3 U315 ( .x(n99), .d0(n281), .sl(B[18]), .d1(n278) );
    nand2_3 U316 ( .x(SUM[18]), .a(n99), .b(n100) );
    aoai211_5 U317 ( .x(n133), .a(n239), .b(n240), .c(n57), .d(n270) );
    aoi21_4 U318 ( .x(n129), .a(n130), .b(n131), .c(n132) );
    nand2i_6 U319 ( .x(n231), .a(n77), .b(n232) );
    inv_5 U32 ( .x(n226), .a(B[1]) );
    nor2_8 U320 ( .x(n122), .a(B[19]), .b(A[19]) );
    nor2i_5 U321 ( .x(n297), .a(n55), .b(n183) );
    nor2i_5 U322 ( .x(n296), .a(B[25]), .b(n183) );
    inv_10 U323 ( .x(n233), .a(B[2]) );
    inv_6 U324 ( .x(n232), .a(n227) );
    inv_10 U325 ( .x(n236), .a(B[8]) );
    nand3_4 U326 ( .x(n227), .a(n228), .b(n229), .c(n230) );
    nand2i_4 U327 ( .x(n178), .a(n106), .b(n292) );
    aoai211_3 U328 ( .x(n299), .a(n333), .b(n332), .c(n93), .d(n294) );
    oaoi211_3 U329 ( .x(n93), .a(n96), .b(n95), .c(n321), .d(n94) );
    nor2_2 U33 ( .x(n78), .a(n80), .b(n79) );
    inv_2 U330 ( .x(n311), .a(n77) );
    aoi21_2 U331 ( .x(n77), .a(n310), .b(n81), .c(n78) );
    aoi21_1 U332 ( .x(n340), .a(n197), .b(n342), .c(n341) );
    inv_2 U333 ( .x(n144), .a(n340) );
    inv_0 U334 ( .x(n341), .a(n175) );
    inv_0 U335 ( .x(n342), .a(n256) );
    inv_0 U336 ( .x(n316), .a(n197) );
    nand2_2 U337 ( .x(n256), .a(n73), .b(n257) );
    exnor2_3 U338 ( .x(SUM[29]), .a(n57), .b(n343) );
    inv_2 U339 ( .x(n343), .a(n53) );
    nand2_0 U34 ( .x(n140), .a(B[0]), .b(A[0]) );
    nand2_1 U340 ( .x(n206), .a(n300), .b(n298) );
    mux2i_3 U341 ( .x(SUM[22]), .d0(n280), .sl(n344), .d1(n137) );
    ao21_3 U342 ( .x(n344), .a(n190), .b(n92), .c(n191) );
    inv_2 U343 ( .x(n262), .a(B[13]) );
    aoi21_1 U35 ( .x(n139), .a(n140), .b(n339), .c(n141) );
    nor2i_1 U36 ( .x(n107), .a(n108), .b(n69) );
    inv_2 U37 ( .x(n108), .a(n97) );
    inv_0 U38 ( .x(n103), .a(n254) );
    inv_2 U39 ( .x(n238), .a(A[9]) );
    inv_2 U40 ( .x(n67), .a(B[9]) );
    nand3i_1 U41 ( .x(n320), .a(n289), .b(n254), .c(n162) );
    inv_2 U42 ( .x(n222), .a(A[7]) );
    inv_2 U43 ( .x(n283), .a(n69) );
    ao21_2 U44 ( .x(n199), .a(n200), .b(n283), .c(n97) );
    nor2i_1 U45 ( .x(SUM[0]), .a(n335), .b(n336) );
    inv_2 U46 ( .x(n266), .a(A[11]) );
    nand2i_2 U47 ( .x(n255), .a(B[11]), .b(n266) );
    nor2i_1 U48 ( .x(n151), .a(n152), .b(n153) );
    nand2_1 U49 ( .x(n152), .a(A[14]), .b(B[14]) );
    oaoi211_4 U5 ( .x(n57), .a(A[28]), .b(B[28]), .c(n334), .d(n90) );
    inv_0 U50 ( .x(n153), .a(n252) );
    and2_5 U51 ( .x(n59), .a(n60), .b(n263) );
    inv_4 U52 ( .x(n263), .a(A[14]) );
    nor2i_0 U53 ( .x(n154), .a(n155), .b(n156) );
    nand2_1 U54 ( .x(n155), .a(B[13]), .b(A[13]) );
    inv_5 U55 ( .x(n156), .a(n319) );
    nor2i_0 U56 ( .x(n109), .a(n110), .b(n111) );
    nand2i_2 U57 ( .x(n249), .a(n121), .b(n146) );
    inv_2 U58 ( .x(n259), .a(n249) );
    and2_3 U59 ( .x(n75), .a(n76), .b(n261) );
    aoai211_3 U6 ( .x(n334), .a(n300), .b(n298), .c(n128), .d(n56) );
    inv_0 U60 ( .x(n279), .a(n273) );
    nor2i_0 U61 ( .x(n281), .a(A[18]), .b(n273) );
    nand2i_2 U62 ( .x(n195), .a(A[29]), .b(n240) );
    nor2i_1 U63 ( .x(n170), .a(B[27]), .b(n171) );
    inv_2 U64 ( .x(n171), .a(A[27]) );
    nor2_1 U65 ( .x(n128), .a(B[27]), .b(A[27]) );
    nor2i_1 U66 ( .x(n126), .a(A[26]), .b(n127) );
    inv_2 U67 ( .x(n127), .a(B[26]) );
    inv_2 U68 ( .x(n183), .a(n323) );
    inv_5 U69 ( .x(n98), .a(B[6]) );
    inv_5 U7 ( .x(n72), .a(A[15]) );
    inv_0 U70 ( .x(n66), .a(A[4]) );
    inv_2 U71 ( .x(n285), .a(n105) );
    inv_2 U72 ( .x(n315), .a(n292) );
    nand2i_5 U74 ( .x(n234), .a(n233), .b(n232) );
    exnor2_1 U75 ( .x(SUM[1]), .a(n338), .b(n335) );
    nand2_2 U76 ( .x(n254), .a(n67), .b(n238) );
    inv_2 U77 ( .x(n326), .a(n220) );
    oai21_1 U78 ( .x(n221), .a(n50), .b(n159), .c(n158) );
    inv_2 U79 ( .x(n325), .a(n221) );
    nand2_5 U8 ( .x(n70), .a(n72), .b(n71) );
    nand2_5 U80 ( .x(n319), .a(n68), .b(n262) );
    oai21_1 U81 ( .x(n220), .a(n156), .b(n325), .c(n155) );
    nor2i_1 U82 ( .x(n148), .a(n149), .b(n150) );
    inv_2 U83 ( .x(n150), .a(n146) );
    nand2_1 U84 ( .x(n149), .a(A[16]), .b(B[16]) );
    inv_2 U85 ( .x(n147), .a(n149) );
    nand2i_2 U86 ( .x(n146), .a(B[16]), .b(n260) );
    inv_5 U87 ( .x(n287), .a(n177) );
    nand2i_2 U88 ( .x(n304), .a(A[22]), .b(n116) );
    inv_0 U89 ( .x(n244), .a(A[22]) );
    oai22_1 U90 ( .x(n188), .a(n116), .b(n244), .c(n138), .d(n118) );
    nor2_1 U91 ( .x(n186), .a(n138), .b(n301) );
    inv_2 U92 ( .x(n138), .a(n304) );
    nand2i_0 U93 ( .x(n190), .a(A[21]), .b(n243) );
    inv_0 U94 ( .x(n243), .a(B[21]) );
    inv_0 U95 ( .x(n125), .a(B[24]) );
    nor2i_1 U96 ( .x(n124), .a(A[24]), .b(n125) );
    oai31_2 U97 ( .x(n194), .a(n117), .b(n138), .c(n119), .d(n271) );
    aoi21_1 U98 ( .x(n294), .a(n194), .b(n295), .c(n124) );
    nand2i_2 U99 ( .x(n332), .a(n322), .b(n331) );
endmodule


module EX_DW01_add_32_1_test_1 ( A, B, CI, SUM, CO );
input  [31:0] A;
input  [31:0] B;
output [31:0] SUM;
input  CI;
output CO;
    wire n253, n199, n200, n201, n89, n90, n91, n92, n132, n137, n133, n134, 
        n82, n249, n218, n184, n94, n143, n262, n263, n250, n278, n270, n101, 
        n217, n198, n135, n181, n152, n227, n223, n254, n255, n229, n237, n215, 
        n203, n248, n142, n228, n195, n119, n121, n75, n98, n157, n158, n144, 
        n145, n159, n129, n54, n247, n153, n154, n155, n156, n140, n139, n50, 
        n160, n161, n194, n112, n85, n100, n188, n108, n70, n103, n95, n93, 
        n151, n226, n120, n245, n49, n71, n164, n66, n51, n60, n177, n59, n234, 
        n122, n202, n252, n56, n55, n124, n235, n77, n83, n73, n258, n169, n57, 
        n128, n189, n264, n216, n58, n221, n53, n267, n146, n147, n260, n207, 
        n130, n162, n214, n186, n251, n180, n61, n179, n149, n150, n138, n78, 
        n63, n279, n213, n62, n65, n136, n72, n99, n64, n206, n67, n238, n76, 
        n52, n74, n68, n224, n265, n69, n87, n275, n204, n81, n80, n79, n231, 
        n230, n182, n185, n192, n268, n269, n211, n209, n243, n131, n261, n205, 
        n172, n208, n105, n106, n107, n109, n110, n111, n113, n114, n115, n116, 
        n117, n118, n123, n125, n126, n127, n171, n170, n174, n175, n168, n183, 
        n190, n196, n197, n219, n210, n176, n220, n222, n225, n187, n236, n232, 
        n212, n163, n266, n277, n276, n102, n233, n166, n97, n167, n191, n193, 
        n148, n240, n272, n241, n242, n274, n246, n244, n178, n141, n239, n273, 
        n271, n256, n257, n165, n173, n259, n86, n88, n104, n84, n96;
    nor3_1 U10 ( .x(n253), .a(n199), .b(n200), .c(n201) );
    nor3i_1 U100 ( .x(n89), .a(n90), .b(n91), .c(n92) );
    nor2i_1 U102 ( .x(n91), .a(n132), .b(n137) );
    nor3i_1 U103 ( .x(n92), .a(n132), .b(n133), .c(n134) );
    exnor2_1 U104 ( .x(SUM[1]), .a(n82), .b(n249) );
    nand2i_2 U105 ( .x(n218), .a(B[9]), .b(n184) );
    nand2_1 U106 ( .x(n94), .a(A[9]), .b(B[9]) );
    nand3_1 U107 ( .x(n143), .a(n262), .b(n263), .c(n250) );
    nand2i_2 U108 ( .x(n262), .a(n278), .b(n270) );
    nand2i_2 U109 ( .x(n263), .a(n101), .b(n217) );
    inv_2 U11 ( .x(n198), .a(A[24]) );
    nor2_1 U110 ( .x(n250), .a(n135), .b(n181) );
    exor2_1 U111 ( .x(n152), .a(A[15]), .b(B[15]) );
    inv_4 U112 ( .x(n227), .a(n223) );
    nand2i_0 U113 ( .x(n254), .a(n255), .b(n227) );
    inv_0 U114 ( .x(n229), .a(n237) );
    nand2i_0 U115 ( .x(n215), .a(A[14]), .b(n203) );
    inv_2 U116 ( .x(n255), .a(n215) );
    exnor2_1 U117 ( .x(SUM[17]), .a(A[17]), .b(n248) );
    oai21_1 U118 ( .x(n248), .a(n142), .b(n228), .c(A[16]) );
    inv_2 U119 ( .x(n195), .a(A[23]) );
    inv_2 U12 ( .x(n201), .a(A[25]) );
    inv_2 U120 ( .x(n119), .a(n199) );
    nor2i_1 U121 ( .x(n121), .a(A[25]), .b(n199) );
    exor2_1 U122 ( .x(SUM[6]), .a(n75), .b(n98) );
    exnor2_1 U123 ( .x(SUM[12]), .a(n157), .b(n158) );
    exnor2_1 U124 ( .x(SUM[7]), .a(n144), .b(n145) );
    exor2_1 U125 ( .x(SUM[11]), .a(n159), .b(n129) );
    buf_1 U126 ( .x(n54), .a(A[20]) );
    exnor2_1 U127 ( .x(SUM[20]), .a(n54), .b(n247) );
    exnor2_1 U128 ( .x(SUM[14]), .a(n153), .b(n154) );
    exnor2_1 U129 ( .x(SUM[13]), .a(n155), .b(n156) );
    nor2i_0 U13 ( .x(n140), .a(n139), .b(n50) );
    exnor2_1 U130 ( .x(SUM[10]), .a(n160), .b(n161) );
    inv_2 U131 ( .x(n194), .a(A[22]) );
    exnor2_1 U132 ( .x(SUM[22]), .a(n112), .b(n194) );
    exnor2_1 U133 ( .x(SUM[5]), .a(n85), .b(n100) );
    inv_0 U134 ( .x(n188), .a(A[19]) );
    exnor2_1 U135 ( .x(SUM[19]), .a(n108), .b(n188) );
    exor2_1 U136 ( .x(SUM[4]), .a(n70), .b(n103) );
    exnor2_1 U137 ( .x(SUM[8]), .a(n89), .b(n95) );
    exor2_1 U138 ( .x(SUM[9]), .a(n143), .b(n93) );
    exor2_1 U139 ( .x(SUM[15]), .a(n151), .b(n152) );
    inv_4 U14 ( .x(n139), .a(n226) );
    inv_2 U140 ( .x(n200), .a(A[26]) );
    exnor2_1 U141 ( .x(SUM[26]), .a(n120), .b(n200) );
    inv_2 U142 ( .x(n245), .a(A[31]) );
    and2_2 U143 ( .x(n49), .a(n71), .b(n164) );
    inv_6 U145 ( .x(n66), .a(n218) );
    oai21_1 U146 ( .x(n51), .a(n60), .b(n177), .c(n59) );
    inv_1 U148 ( .x(n234), .a(A[28]) );
    exnor2_1 U149 ( .x(SUM[28]), .a(n122), .b(n234) );
    inv_0 U15 ( .x(n202), .a(B[15]) );
    nor2i_1 U150 ( .x(n252), .a(n56), .b(n234) );
    inv_2 U151 ( .x(n55), .a(n234) );
    exnor2_1 U152 ( .x(SUM[29]), .a(n124), .b(n235) );
    inv_2 U153 ( .x(n56), .a(n235) );
    inv_2 U154 ( .x(n235), .a(A[29]) );
    aoi21_1 U155 ( .x(n82), .a(n77), .b(A[1]), .c(n83) );
    and2_2 U156 ( .x(n73), .a(B[1]), .b(A[1]) );
    nand2i_2 U157 ( .x(n258), .a(A[1]), .b(n169) );
    inv_2 U158 ( .x(n57), .a(n128) );
    nand4_1 U159 ( .x(n189), .a(A[19]), .b(A[18]), .c(A[16]), .d(A[17]) );
    nand2i_2 U16 ( .x(n264), .a(A[15]), .b(n202) );
    ao21_1 U160 ( .x(n216), .a(n58), .b(n184), .c(n278) );
    inv_0 U161 ( .x(n58), .a(B[9]) );
    inv_2 U162 ( .x(n184), .a(A[9]) );
    nand2i_2 U163 ( .x(n158), .a(n221), .b(n53) );
    inv_2 U164 ( .x(n221), .a(n267) );
    exor2_1 U165 ( .x(SUM[3]), .a(n146), .b(n147) );
    oai21_2 U166 ( .x(n260), .a(A[3]), .b(n146), .c(B[3]) );
    inv_0 U167 ( .x(n207), .a(A[11]) );
    nand2_0 U168 ( .x(n130), .a(A[11]), .b(B[11]) );
    inv_2 U169 ( .x(n162), .a(A[8]) );
    inv_2 U17 ( .x(n214), .a(n264) );
    nand2_1 U170 ( .x(n186), .a(B[7]), .b(A[7]) );
    inv_2 U171 ( .x(n59), .a(n251) );
    inv_0 U172 ( .x(n60), .a(B[4]) );
    inv_0 U173 ( .x(n180), .a(n177) );
    inv_2 U174 ( .x(n251), .a(n101) );
    inv_2 U175 ( .x(n61), .a(n179) );
    exnor2_1 U176 ( .x(SUM[16]), .a(n149), .b(n150) );
    nand2i_6 U177 ( .x(n149), .a(n138), .b(n78) );
    inv_0 U178 ( .x(n179), .a(B[4]) );
    nor2_0 U179 ( .x(n63), .a(n279), .b(n66) );
    nand2i_2 U18 ( .x(n213), .a(n214), .b(n215) );
    nor2_0 U180 ( .x(n62), .a(n278), .b(n66) );
    nor2_3 U181 ( .x(n65), .a(n136), .b(n66) );
    aoi31_3 U182 ( .x(n72), .a(A[0]), .b(n258), .c(B[0]), .d(n73) );
    nand2_1 U183 ( .x(n99), .a(A[6]), .b(B[6]) );
    inv_5 U184 ( .x(n169), .a(B[1]) );
    inv_2 U185 ( .x(n64), .a(n53) );
    nand2i_1 U186 ( .x(n267), .a(B[12]), .b(n206) );
    inv_0 U187 ( .x(n217), .a(n279) );
    inv_2 U188 ( .x(n128), .a(A[30]) );
    inv_2 U189 ( .x(n67), .a(n238) );
    ao21_1 U19 ( .x(n76), .a(n52), .b(n74), .c(n51) );
    inv_2 U190 ( .x(n68), .a(n224) );
    nand2_0 U191 ( .x(n238), .a(B[13]), .b(A[13]) );
    inv_2 U192 ( .x(n224), .a(n265) );
    inv_0 U193 ( .x(n69), .a(n87) );
    inv_2 U194 ( .x(n70), .a(n69) );
    inv_0 U195 ( .x(n71), .a(B[6]) );
    nand2_0 U196 ( .x(n153), .a(n229), .b(n275) );
    oai221_1 U197 ( .x(n151), .a(n255), .b(n229), .c(n50), .d(n254), .e(n204)
         );
    nand2_0 U198 ( .x(n249), .a(A[0]), .b(B[0]) );
    exor2_1 U199 ( .x(SUM[0]), .a(A[0]), .b(B[0]) );
    exor2_1 U200 ( .x(n147), .a(B[3]), .b(A[3]) );
    inv_0 U201 ( .x(n83), .a(n258) );
    inv_0 U202 ( .x(n77), .a(n169) );
    aoi211_5 U203 ( .x(n78), .a(n237), .b(n81), .c(n80), .d(n79) );
    inv_2 U204 ( .x(n79), .a(n231) );
    inv_2 U205 ( .x(n81), .a(n213) );
    nand2_0 U206 ( .x(n231), .a(A[15]), .b(B[15]) );
    nand2i_2 U207 ( .x(n230), .a(n204), .b(n264) );
    aoi21_1 U208 ( .x(n90), .a(n251), .b(n132), .c(n182) );
    oai21_2 U209 ( .x(n182), .a(n185), .b(n99), .c(n186) );
    nand2_1 U21 ( .x(n192), .a(n54), .b(A[21]) );
    aoai211_1 U210 ( .x(n159), .a(n268), .b(n269), .c(n211), .d(n209) );
    nand2i_0 U211 ( .x(n161), .a(n211), .b(n209) );
    oai21_1 U212 ( .x(n243), .a(n131), .b(n209), .c(n130) );
    inv_0 U213 ( .x(n203), .a(B[14]) );
    nand2_0 U214 ( .x(n204), .a(A[14]), .b(B[14]) );
    nor2i_0 U215 ( .x(n98), .a(n99), .b(n49) );
    inv_0 U216 ( .x(n261), .a(n99) );
    nand2i_0 U217 ( .x(n265), .a(A[13]), .b(n205) );
    inv_0 U218 ( .x(n205), .a(B[13]) );
    nand2_0 U219 ( .x(n209), .a(B[10]), .b(A[10]) );
    nand2_1 U22 ( .x(n172), .a(B[2]), .b(A[2]) );
    inv_0 U220 ( .x(n208), .a(B[10]) );
    nor2i_5 U221 ( .x(n93), .a(n94), .b(n66) );
    nor2i_3 U222 ( .x(n105), .a(n106), .b(n107) );
    nor2i_3 U223 ( .x(n108), .a(n109), .b(n107) );
    nor2i_3 U224 ( .x(n110), .a(n111), .b(n107) );
    nor2i_3 U225 ( .x(n112), .a(n113), .b(n107) );
    nor2i_3 U226 ( .x(n114), .a(n115), .b(n107) );
    nor2i_3 U227 ( .x(n116), .a(n117), .b(n107) );
    nor2i_3 U228 ( .x(n118), .a(n119), .b(n107) );
    nor2i_3 U229 ( .x(n120), .a(n121), .b(n107) );
    nor2i_1 U23 ( .x(n106), .a(A[17]), .b(n150) );
    nor2i_3 U230 ( .x(n122), .a(n123), .b(n107) );
    nor2i_3 U231 ( .x(n124), .a(n125), .b(n107) );
    nor2_5 U232 ( .x(n126), .a(n127), .b(n128) );
    aoai211_4 U234 ( .x(n146), .a(n171), .b(n170), .c(n72), .d(n172) );
    nand2_5 U235 ( .x(n174), .a(n74), .b(n175) );
    ao21_4 U236 ( .x(n181), .a(n182), .b(n168), .c(n183) );
    inv_6 U237 ( .x(n190), .a(A[21]) );
    nand2i_4 U238 ( .x(n196), .a(n197), .b(n113) );
    nand2i_4 U239 ( .x(n219), .a(n210), .b(n65) );
    nand2i_2 U24 ( .x(n175), .a(n61), .b(n176) );
    nand2i_4 U240 ( .x(n220), .a(n221), .b(n222) );
    nand2i_4 U241 ( .x(n223), .a(n224), .b(n225) );
    nand2i_4 U242 ( .x(n226), .a(n213), .b(n227) );
    exnor2_5 U243 ( .x(SUM[31]), .a(n126), .b(n245) );
    exnor2_5 U244 ( .x(SUM[25]), .a(n118), .b(n201) );
    exnor2_5 U245 ( .x(SUM[24]), .a(n116), .b(n198) );
    exnor2_5 U246 ( .x(SUM[23]), .a(n114), .b(n195) );
    exnor2_5 U247 ( .x(SUM[21]), .a(n110), .b(n190) );
    exnor2_5 U248 ( .x(SUM[18]), .a(n105), .b(n187) );
    nand2_2 U249 ( .x(n197), .a(A[22]), .b(A[23]) );
    inv_2 U25 ( .x(n176), .a(A[4]) );
    nor2i_5 U250 ( .x(n236), .a(n252), .b(n232) );
    nor2i_5 U251 ( .x(n125), .a(n55), .b(n232) );
    nand2i_4 U252 ( .x(n212), .a(B[11]), .b(n207) );
    inv_5 U253 ( .x(n225), .a(n220) );
    inv_5 U254 ( .x(n117), .a(n196) );
    nor2i_5 U255 ( .x(n138), .a(n139), .b(n50) );
    inv_10 U256 ( .x(n107), .a(n149) );
    inv_10 U257 ( .x(n171), .a(B[2]) );
    inv_16 U258 ( .x(n170), .a(A[2]) );
    nand2i_6 U259 ( .x(n127), .a(n107), .b(n236) );
    inv_2 U26 ( .x(n133), .a(n175) );
    nand2i_6 U261 ( .x(n199), .a(n198), .b(n117) );
    inv_7 U263 ( .x(n163), .a(B[7]) );
    nand2i_5 U264 ( .x(n266), .a(A[10]), .b(n208) );
    oai21_1 U265 ( .x(n75), .a(n277), .b(n134), .c(n276) );
    inv_0 U266 ( .x(n276), .a(n51) );
    inv_2 U267 ( .x(n277), .a(n52) );
    or2_1 U268 ( .x(n52), .a(B[4]), .b(A[4]) );
    nand2i_4 U269 ( .x(n134), .a(n102), .b(n87) );
    nand2i_2 U27 ( .x(n232), .a(n233), .b(n119) );
    or2_6 U270 ( .x(n136), .a(n166), .b(n97) );
    or2_1 U271 ( .x(n279), .a(n166), .b(n97) );
    or2_1 U272 ( .x(n278), .a(n166), .b(n97) );
    inv_0 U273 ( .x(n132), .a(n166) );
    nand2i_2 U274 ( .x(n168), .a(B[8]), .b(n162) );
    inv_3 U275 ( .x(n97), .a(n168) );
    nand2i_3 U276 ( .x(n166), .a(n49), .b(n167) );
    nor2_0 U28 ( .x(n135), .a(n279), .b(n137) );
    nand2i_2 U29 ( .x(n137), .a(n179), .b(n180) );
    nor2i_1 U30 ( .x(n142), .a(n139), .b(n50) );
    aoi21_3 U31 ( .x(n50), .a(n52), .b(n74), .c(n51) );
    nor2i_1 U32 ( .x(n111), .a(n54), .b(n189) );
    nor2i_1 U33 ( .x(n115), .a(A[22]), .b(n191) );
    nand2i_2 U34 ( .x(n191), .a(n192), .b(n193) );
    inv_2 U35 ( .x(n113), .a(n191) );
    exor2_1 U36 ( .x(n148), .a(B[2]), .b(A[2]) );
    exnor2_1 U37 ( .x(SUM[2]), .a(n72), .b(n148) );
    inv_0 U38 ( .x(n164), .a(A[6]) );
    inv_5 U40 ( .x(n74), .a(n134) );
    nand2_0 U41 ( .x(n53), .a(A[12]), .b(B[12]) );
    inv_0 U42 ( .x(n206), .a(A[12]) );
    nand2i_0 U43 ( .x(n157), .a(n240), .b(n272) );
    ao21_3 U44 ( .x(n240), .a(n241), .b(n242), .c(n243) );
    nand2i_2 U45 ( .x(n272), .a(n219), .b(n75) );
    nand2i_2 U46 ( .x(n145), .a(n185), .b(n186) );
    inv_2 U47 ( .x(n185), .a(n167) );
    nand2i_3 U48 ( .x(n167), .a(A[7]), .b(n163) );
    nand2i_2 U49 ( .x(n144), .a(n261), .b(n274) );
    nand3_1 U5 ( .x(n233), .a(A[27]), .b(A[26]), .c(A[25]) );
    nand2i_2 U50 ( .x(n274), .a(n49), .b(n76) );
    inv_4 U51 ( .x(n228), .a(n78) );
    oai21_1 U52 ( .x(n246), .a(n140), .b(n228), .c(n253) );
    exnor2_1 U53 ( .x(SUM[27]), .a(A[27]), .b(n246) );
    inv_2 U54 ( .x(n131), .a(n212) );
    nor2i_1 U55 ( .x(n129), .a(n130), .b(n131) );
    inv_0 U56 ( .x(n268), .a(n242) );
    oai21_2 U57 ( .x(n242), .a(n66), .b(n244), .c(n94) );
    inv_2 U58 ( .x(n244), .a(n181) );
    nand2i_2 U59 ( .x(n269), .a(n216), .b(n75) );
    nand2i_2 U6 ( .x(n177), .a(n176), .b(n178) );
    oai21_1 U60 ( .x(n247), .a(n141), .b(n228), .c(n193) );
    nor2i_0 U61 ( .x(n141), .a(n139), .b(n50) );
    inv_2 U62 ( .x(n80), .a(n230) );
    nand2i_2 U63 ( .x(n154), .a(n255), .b(n204) );
    ao21_3 U64 ( .x(n237), .a(n68), .b(n239), .c(n67) );
    nand2i_0 U65 ( .x(n275), .a(n223), .b(n76) );
    nand2i_2 U66 ( .x(n156), .a(n224), .b(n238) );
    nand2i_2 U67 ( .x(n155), .a(n239), .b(n273) );
    ao21_3 U68 ( .x(n239), .a(n267), .b(n240), .c(n64) );
    nand2i_0 U69 ( .x(n273), .a(n220), .b(n76) );
    inv_0 U7 ( .x(n241), .a(n210) );
    inv_2 U70 ( .x(n211), .a(n266) );
    oai211_1 U71 ( .x(n160), .a(n174), .b(n216), .c(n271), .d(n256) );
    nand2i_2 U72 ( .x(n271), .a(n101), .b(n62) );
    aoi21_1 U73 ( .x(n256), .a(n63), .b(n257), .c(n242) );
    inv_2 U74 ( .x(n257), .a(n137) );
    inv_2 U75 ( .x(n270), .a(n174) );
    inv_2 U76 ( .x(n193), .a(n189) );
    nor2i_1 U77 ( .x(n100), .a(n101), .b(n102) );
    nand2_1 U78 ( .x(n101), .a(A[5]), .b(B[5]) );
    inv_2 U79 ( .x(n102), .a(n178) );
    inv_2 U8 ( .x(n222), .a(n219) );
    nand2i_2 U80 ( .x(n178), .a(B[5]), .b(n165) );
    inv_0 U81 ( .x(n165), .a(A[5]) );
    inv_2 U82 ( .x(n173), .a(A[3]) );
    inv_1 U83 ( .x(n259), .a(n146) );
    nand2i_2 U84 ( .x(n86), .a(n61), .b(n176) );
    aoi21_1 U85 ( .x(n85), .a(n86), .b(n70), .c(n88) );
    inv_0 U86 ( .x(n150), .a(A[16]) );
    and3i_1 U87 ( .x(n109), .a(n150), .b(A[18]), .c(A[17]) );
    oai21_2 U88 ( .x(n87), .a(n259), .b(n173), .c(n260) );
    nor2i_1 U89 ( .x(n103), .a(n104), .b(n84) );
    nand2i_2 U9 ( .x(n210), .a(n211), .b(n212) );
    nand2_2 U90 ( .x(n104), .a(n61), .b(A[4]) );
    nor2_1 U91 ( .x(n84), .a(n61), .b(A[4]) );
    inv_2 U92 ( .x(n88), .a(n104) );
    inv_2 U93 ( .x(n187), .a(A[18]) );
    exnor2_3 U94 ( .x(SUM[30]), .a(n127), .b(n57) );
    inv_2 U95 ( .x(n123), .a(n232) );
    inv_2 U96 ( .x(n183), .a(n96) );
    nand2_0 U98 ( .x(n96), .a(A[8]), .b(B[8]) );
    nor2i_1 U99 ( .x(n95), .a(n96), .b(n97) );
endmodule


module EX_DW01_cmp2_32_3_test_1 ( A, B, LEQ, TC, LT_LE, GE_GT );
input  [31:0] A;
input  [31:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n76, n107, n123, n72, n15, n62, n61, n37, n64, n63, n137, n17, n49, 
        n19, n18, n66, n71, n102, n101, n65, n124, n73, n142, n94, n93, n68, 
        n26, n106, n119, n53, n56, n27, n91, n34, n33, n97, n129, n117, n136, 
        n48, n55, n143, n57, n22, n20, n21, n74, n75, n77, n121, n38, n103, 
        n104, n79, n115, n112, n130, n131, n96, n132, n133, n46, n114, n60, 
        n144, n145, n139, n69, n89, n39, n134, n135, n108, n141, n92, n120, 
        n100, n24, n99, n98, n105, n113, n126, n47, n122, n45, n35, n44, n90, 
        n138, n16, n28, n31, n29, n30, n87, n88, n118, n32, n116, n95, n81, 
        n52, n80, n140, n58, n54, n23, n25, n59, n109, n111, n110, n78, n70, 
        n67, n36, n84, n43, n125, n127, n128, n40, n41, n42, n82, n86, n85, 
        n50, n51, n83;
    nand2i_2 U10 ( .x(n76), .a(n107), .b(n123) );
    inv_2 U100 ( .x(n72), .a(A[28]) );
    oa22_1 U101 ( .x(n15), .a(B[15]), .b(n62), .c(B[16]), .d(n61) );
    oai22_1 U102 ( .x(n37), .a(A[14]), .b(n64), .c(A[15]), .d(n63) );
    nand2i_2 U105 ( .x(n137), .a(A[24]), .b(B[24]) );
    inv_2 U106 ( .x(n17), .a(n49) );
    inv_2 U107 ( .x(n49), .a(A[1]) );
    inv_2 U108 ( .x(n19), .a(n18) );
    inv_2 U109 ( .x(n18), .a(B[30]) );
    inv_2 U110 ( .x(n66), .a(B[19]) );
    nand4_1 U111 ( .x(n71), .a(A[17]), .b(n102), .c(n101), .d(n65) );
    aoi22_1 U112 ( .x(n124), .a(A[30]), .b(n18), .c(A[29]), .d(n73) );
    oai22_1 U114 ( .x(n142), .a(B[6]), .b(n94), .c(B[5]), .d(n93) );
    aoi21_1 U115 ( .x(n68), .a(A[20]), .b(n26), .c(n106) );
    aoi22_1 U116 ( .x(n119), .a(A[13]), .b(n53), .c(A[14]), .d(n64) );
    inv_1 U117 ( .x(n56), .a(B[8]) );
    nor2i_0 U118 ( .x(n27), .a(A[8]), .b(B[8]) );
    inv_0 U119 ( .x(n91), .a(A[11]) );
    nor2i_0 U120 ( .x(n34), .a(B[11]), .b(A[11]) );
    nor2i_0 U121 ( .x(n33), .a(B[3]), .b(A[3]) );
    inv_0 U122 ( .x(n97), .a(A[0]) );
    inv_0 U123 ( .x(n129), .a(B[7]) );
    oai22_1 U124 ( .x(n117), .a(B[7]), .b(n136), .c(n136), .d(n48) );
    inv_0 U125 ( .x(n55), .a(A[9]) );
    oai22_1 U126 ( .x(n143), .a(A[9]), .b(n57), .c(A[8]), .d(n56) );
    inv_0 U127 ( .x(n53), .a(B[13]) );
    and3i_3 U128 ( .x(LT_LE), .a(n22), .b(n20), .c(n21) );
    nand3_3 U129 ( .x(n74), .a(n75), .b(n76), .c(n77) );
    nand2i_3 U13 ( .x(n121), .a(B[27]), .b(A[27]) );
    nand4_1 U130 ( .x(n38), .a(n101), .b(n102), .c(n103), .d(n104) );
    nor3i_5 U131 ( .x(n79), .a(n115), .b(n112), .c(n74) );
    aoi22_3 U132 ( .x(n21), .a(n130), .b(n131), .c(n96), .d(n130) );
    aoi22_3 U133 ( .x(n20), .a(n132), .b(n130), .c(n133), .d(n130) );
    nand4_1 U134 ( .x(n46), .a(A[23]), .b(n114), .c(n137), .d(n60) );
    nand4_1 U135 ( .x(n144), .a(n145), .b(n15), .c(n119), .d(n139) );
    nand2i_5 U136 ( .x(n69), .a(B[22]), .b(A[22]) );
    nand2i_5 U137 ( .x(n107), .a(A[27]), .b(B[27]) );
    inv_0 U138 ( .x(n89), .a(A[29]) );
    nand3i_2 U139 ( .x(n22), .a(n39), .b(n134), .c(n135) );
    nand3_1 U14 ( .x(n75), .a(n121), .b(n108), .c(n123) );
    inv_0 U140 ( .x(n62), .a(A[15]) );
    nand2i_1 U141 ( .x(n141), .a(A[6]), .b(B[6]) );
    inv_0 U142 ( .x(n92), .a(A[23]) );
    nand2i_4 U143 ( .x(n123), .a(B[28]), .b(A[28]) );
    nor2i_2 U144 ( .x(n108), .a(B[26]), .b(A[26]) );
    nor2i_0 U145 ( .x(n120), .a(A[24]), .b(B[24]) );
    nand2i_2 U15 ( .x(n114), .a(A[25]), .b(B[25]) );
    nor2i_1 U16 ( .x(n100), .a(n19), .b(A[30]) );
    nand2i_0 U17 ( .x(n24), .a(A[20]), .b(n99) );
    nand2i_2 U18 ( .x(n98), .a(A[21]), .b(B[21]) );
    nor2i_1 U19 ( .x(n105), .a(A[18]), .b(B[18]) );
    nand2i_2 U20 ( .x(n99), .a(B[21]), .b(A[21]) );
    nand2i_2 U21 ( .x(n104), .a(A[16]), .b(B[16]) );
    nand2i_0 U22 ( .x(n103), .a(A[17]), .b(B[17]) );
    nand2i_2 U23 ( .x(n102), .a(A[18]), .b(B[18]) );
    nand2i_2 U24 ( .x(n101), .a(A[19]), .b(B[19]) );
    nand2i_2 U25 ( .x(n113), .a(A[31]), .b(B[31]) );
    nand2i_2 U26 ( .x(n126), .a(B[31]), .b(A[31]) );
    inv_2 U27 ( .x(n73), .a(B[29]) );
    nand3_1 U28 ( .x(n47), .a(n121), .b(n122), .c(n123) );
    inv_2 U29 ( .x(n60), .a(B[23]) );
    aoi21_1 U30 ( .x(n45), .a(n120), .b(n114), .c(n35) );
    and3i_1 U31 ( .x(n44), .a(n47), .b(n45), .c(n46) );
    inv_0 U32 ( .x(n90), .a(A[12]) );
    oai22_1 U33 ( .x(n138), .a(B[11]), .b(n91), .c(B[12]), .d(n90) );
    nand2_2 U34 ( .x(n139), .a(n16), .b(n138) );
    and3i_1 U35 ( .x(n28), .a(n31), .b(n29), .c(n30) );
    nand2i_0 U36 ( .x(n29), .a(B[3]), .b(A[3]) );
    nand2i_2 U37 ( .x(n30), .a(B[2]), .b(A[2]) );
    nand3_1 U38 ( .x(n31), .a(n87), .b(n97), .c(n88) );
    oai211_1 U39 ( .x(n118), .a(n32), .b(n33), .c(n29), .d(n87) );
    nor2i_0 U40 ( .x(n32), .a(B[2]), .b(A[2]) );
    nand2i_2 U41 ( .x(n87), .a(B[4]), .b(A[4]) );
    inv_2 U42 ( .x(n136), .a(n141) );
    or3i_2 U43 ( .x(n116), .a(n95), .b(n132), .c(n133) );
    and3i_1 U44 ( .x(n95), .a(n96), .b(n49), .c(B[1]) );
    nand2i_0 U45 ( .x(n81), .a(A[10]), .b(B[10]) );
    oa22_1 U46 ( .x(n16), .a(A[13]), .b(n53), .c(A[12]), .d(n52) );
    inv_2 U47 ( .x(n52), .a(B[12]) );
    nand2_2 U48 ( .x(n80), .a(n140), .b(n143) );
    inv_2 U49 ( .x(n140), .a(n58) );
    oai22_1 U50 ( .x(n58), .a(B[9]), .b(n55), .c(B[10]), .d(n54) );
    inv_2 U51 ( .x(n57), .a(B[9]) );
    nand2_2 U52 ( .x(n112), .a(n113), .b(n114) );
    nand2_2 U53 ( .x(n115), .a(n100), .b(n126) );
    inv_0 U54 ( .x(n26), .a(B[20]) );
    nor3_1 U55 ( .x(n23), .a(n24), .b(n25), .c(n26) );
    inv_0 U56 ( .x(n59), .a(B[22]) );
    oai22_1 U57 ( .x(n109), .a(A[22]), .b(n59), .c(n25), .d(n98) );
    inv_2 U58 ( .x(n111), .a(n137) );
    aoi21_1 U59 ( .x(n110), .a(B[23]), .b(n92), .c(n111) );
    nand2i_2 U6 ( .x(n122), .a(B[26]), .b(A[26]) );
    nor3i_1 U60 ( .x(n78), .a(n110), .b(n109), .c(n23) );
    inv_2 U61 ( .x(n25), .a(n69) );
    inv_0 U62 ( .x(n65), .a(B[17]) );
    aoi22_1 U63 ( .x(n70), .a(A[19]), .b(n66), .c(n105), .d(n101) );
    inv_2 U64 ( .x(n106), .a(n99) );
    nand4_1 U65 ( .x(n67), .a(n68), .b(n69), .c(n70), .d(n71) );
    inv_0 U66 ( .x(n63), .a(B[15]) );
    inv_2 U67 ( .x(n64), .a(B[14]) );
    aoi21_1 U68 ( .x(n36), .a(n15), .b(n37), .c(n38) );
    nand2i_2 U69 ( .x(n135), .a(n88), .b(n130) );
    nor2i_1 U7 ( .x(n35), .a(A[25]), .b(B[25]) );
    nand2i_2 U70 ( .x(n88), .a(B[1]), .b(n17) );
    inv_2 U71 ( .x(n84), .a(n43) );
    aoai211_1 U72 ( .x(n134), .a(n84), .b(n144), .c(n125), .d(n127) );
    inv_2 U73 ( .x(n145), .a(n67) );
    oai211_1 U74 ( .x(n125), .a(n44), .b(n74), .c(n124), .d(n126) );
    nor2i_1 U75 ( .x(n127), .a(n115), .b(n128) );
    inv_2 U76 ( .x(n128), .a(n113) );
    aoi211_1 U77 ( .x(n39), .a(n40), .b(n41), .c(n42), .d(n43) );
    nand2_2 U78 ( .x(n40), .a(n142), .b(n117) );
    aoi211_1 U79 ( .x(n41), .a(A[7]), .b(n129), .c(n27), .d(n58) );
    oai211_3 U80 ( .x(n43), .a(n36), .b(n67), .c(n78), .d(n79) );
    inv_5 U81 ( .x(n130), .a(n82) );
    and4i_1 U82 ( .x(n86), .a(n28), .b(n116), .c(n117), .d(n118) );
    nand4i_1 U83 ( .x(n42), .a(n34), .b(n80), .c(n16), .d(n81) );
    inv_2 U84 ( .x(n85), .a(n42) );
    inv_2 U85 ( .x(n50), .a(B[4]) );
    inv_2 U86 ( .x(n51), .a(B[5]) );
    oai22_1 U87 ( .x(n83), .a(A[5]), .b(n51), .c(A[4]), .d(n50) );
    nand4i_1 U88 ( .x(n82), .a(n83), .b(n84), .c(n85), .d(n86) );
    inv_0 U89 ( .x(n54), .a(A[10]) );
    aoi22_1 U9 ( .x(n77), .a(B[29]), .b(n89), .c(B[28]), .d(n72) );
    inv_2 U90 ( .x(n132), .a(n29) );
    inv_2 U91 ( .x(n133), .a(n30) );
    inv_2 U92 ( .x(n131), .a(B[0]) );
    inv_2 U93 ( .x(n96), .a(n87) );
    inv_0 U95 ( .x(n61), .a(A[16]) );
    inv_0 U96 ( .x(n93), .a(A[5]) );
    inv_2 U97 ( .x(n48), .a(A[7]) );
    inv_0 U99 ( .x(n94), .a(A[6]) );
endmodule


module EX_DW01_cmp2_32_0 ( A, B, LEQ, TC, LT_LE, GE_GT );
input  [31:0] A;
input  [31:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n81, n62, n110, n112, n16, n54, n53, n45, n17, n18, n84, n19, n21, 
        n20, n65, n131, n22, n75, n76, n68, n99, n100, n74, n27, n28, n25, n82, 
        n97, n98, n94, n128, n127, n71, n80, n78, n116, n92, n107, n60, n56, 
        n55, n132, n42, n118, n133, n130, n134, n126, n120, n122, n138, n135, 
        n142, n24, n143, n41, n43, n146, n77, n147, n26, n113, n114, n72, n73, 
        n115, n108, n63, n129, n31, n90, n117, n93, n66, n64, n70, n50, n51, 
        n52, n89, n15, n44, n33, n144, n141, n145, n88, n91, n158, n119, n121, 
        n86, n83, n157, n155, n123, n156, n58, n104, n101, n39, n57, n49, n105, 
        n40, n140, n87, n96, n154, n67, n47, n46, n37, n35, n38, n34, n36, 
        n152, n48, n103, n102, n106, n136, n137, n32, n95, n29, n111, n109, 
        n79, n85, n124, n30, n125, n59, n61, n69, n139, n148, n149, n150, n151, 
        n153, n23;
    aoi211_1 U10 ( .x(n81), .a(A[20]), .b(n62), .c(n110), .d(n112) );
    oa22_2 U100 ( .x(n16), .a(A[31]), .b(n54), .c(A[30]), .d(n53) );
    nand2_2 U101 ( .x(n45), .a(n17), .b(B[11]) );
    inv_0 U102 ( .x(n17), .a(A[11]) );
    inv_2 U103 ( .x(n18), .a(n62) );
    inv_2 U104 ( .x(n62), .a(B[20]) );
    inv_2 U105 ( .x(n84), .a(A[3]) );
    inv_2 U106 ( .x(n19), .a(n53) );
    inv_2 U107 ( .x(n53), .a(B[30]) );
    inv_2 U108 ( .x(n21), .a(n20) );
    inv_0 U109 ( .x(n65), .a(B[13]) );
    nand2i_2 U11 ( .x(n131), .a(B[22]), .b(A[22]) );
    inv_0 U110 ( .x(n22), .a(n75) );
    inv_2 U111 ( .x(n76), .a(n68) );
    nand2_2 U112 ( .x(n75), .a(n99), .b(n100) );
    inv_2 U113 ( .x(n74), .a(n45) );
    oai22_1 U114 ( .x(n27), .a(B[5]), .b(n28), .c(B[6]), .d(n25) );
    nand4_1 U115 ( .x(n82), .a(A[17]), .b(n97), .c(n98), .d(n94) );
    nor2i_0 U116 ( .x(n128), .a(B[17]), .b(A[17]) );
    inv_0 U117 ( .x(n28), .a(A[5]) );
    nand2i_0 U118 ( .x(n127), .a(A[5]), .b(B[5]) );
    inv_1 U119 ( .x(n71), .a(B[8]) );
    aoi22_1 U12 ( .x(n80), .a(A[19]), .b(n78), .c(n116), .d(n98) );
    inv_0 U120 ( .x(n92), .a(B[3]) );
    nand2i_0 U121 ( .x(n107), .a(B[24]), .b(A[24]) );
    oai22_1 U122 ( .x(n60), .a(A[25]), .b(n56), .c(A[24]), .d(n55) );
    oai31_1 U123 ( .x(n132), .a(n42), .b(n118), .c(n133), .d(n130) );
    oai222_1 U124 ( .x(n134), .a(n42), .b(n126), .c(n42), .d(n120), .e(n42), 
        .f(n122) );
    oai31_1 U125 ( .x(n138), .a(n42), .b(n127), .c(n27), .d(n135) );
    oai21_1 U126 ( .x(n142), .a(n24), .b(n42), .c(n143) );
    nor2_2 U127 ( .x(n41), .a(n42), .b(n43) );
    oai21_1 U128 ( .x(n146), .a(n42), .b(n77), .c(n147) );
    aoi22_1 U129 ( .x(n24), .a(B[6]), .b(n25), .c(B[7]), .d(n26) );
    inv_2 U13 ( .x(n78), .a(B[19]) );
    nand2i_0 U130 ( .x(n113), .a(B[7]), .b(A[7]) );
    nand2i_0 U131 ( .x(n114), .a(B[8]), .b(A[8]) );
    oai22_1 U132 ( .x(n100), .a(A[9]), .b(n72), .c(A[8]), .d(n71) );
    nand4i_1 U133 ( .x(n73), .a(n74), .b(n75), .c(n76), .d(n77) );
    inv_2 U134 ( .x(n115), .a(n77) );
    nand2i_4 U135 ( .x(n77), .a(A[10]), .b(B[10]) );
    nor2i_0 U136 ( .x(n108), .a(B[21]), .b(A[21]) );
    inv_0 U137 ( .x(n63), .a(A[16]) );
    nand2i_0 U138 ( .x(n129), .a(A[16]), .b(B[16]) );
    inv_0 U139 ( .x(n31), .a(A[14]) );
    nor2i_1 U14 ( .x(n116), .a(A[18]), .b(B[18]) );
    aoi222_1 U140 ( .x(n90), .a(n76), .b(n117), .c(A[13]), .d(n65), .e(A[14]), 
        .f(n93) );
    inv_0 U141 ( .x(n66), .a(A[12]) );
    oai22_1 U142 ( .x(n68), .a(A[13]), .b(n65), .c(A[12]), .d(n64) );
    inv_0 U143 ( .x(n25), .a(A[6]) );
    inv_0 U144 ( .x(n70), .a(A[10]) );
    aoi21_3 U145 ( .x(LT_LE), .a(n50), .b(n51), .c(n52) );
    nor3i_5 U146 ( .x(n89), .a(n15), .b(n44), .c(n33) );
    nand2i_4 U147 ( .x(n144), .a(n142), .b(n141) );
    nor3_4 U148 ( .x(n50), .a(n144), .b(n145), .c(n146) );
    nand4_5 U149 ( .x(n42), .a(n88), .b(n89), .c(n90), .d(n91) );
    nand2i_0 U15 ( .x(n158), .a(B[21]), .b(A[21]) );
    nand3i_5 U150 ( .x(n120), .a(A[0]), .b(n119), .c(n121) );
    oai22_1 U16 ( .x(n86), .a(B[3]), .b(n84), .c(B[4]), .d(n83) );
    nand2i_2 U17 ( .x(n157), .a(B[1]), .b(A[1]) );
    or3i_2 U18 ( .x(n155), .a(n123), .b(n156), .c(A[2]) );
    aoi21_1 U19 ( .x(n58), .a(n104), .b(n101), .c(n39) );
    nor2i_1 U20 ( .x(n104), .a(n21), .b(A[27]) );
    nor2i_1 U21 ( .x(n39), .a(B[28]), .b(A[28]) );
    nand3_1 U22 ( .x(n57), .a(n49), .b(n105), .c(n101) );
    inv_0 U23 ( .x(n20), .a(B[27]) );
    nor2i_1 U24 ( .x(n105), .a(B[26]), .b(A[26]) );
    nor2i_1 U25 ( .x(n40), .a(B[29]), .b(A[29]) );
    nand2i_2 U26 ( .x(n140), .a(A[23]), .b(B[23]) );
    nand2i_2 U27 ( .x(n97), .a(A[18]), .b(B[18]) );
    oai31_2 U28 ( .x(n121), .a(n87), .b(n156), .c(n86), .d(n155) );
    inv_2 U29 ( .x(n96), .a(B[0]) );
    nand3i_1 U30 ( .x(n43), .a(n96), .b(n119), .c(n121) );
    nand2i_2 U31 ( .x(n98), .a(A[19]), .b(B[19]) );
    nand2i_2 U32 ( .x(n91), .a(n113), .b(n154) );
    inv_2 U33 ( .x(n154), .a(n73) );
    inv_2 U34 ( .x(n93), .a(B[14]) );
    inv_0 U35 ( .x(n67), .a(A[11]) );
    oai22_1 U36 ( .x(n117), .a(B[11]), .b(n67), .c(B[12]), .d(n66) );
    nand3_1 U37 ( .x(n33), .a(n80), .b(n81), .c(n82) );
    and3i_1 U38 ( .x(n44), .a(n47), .b(n45), .c(n46) );
    nand2i_2 U39 ( .x(n88), .a(n114), .b(n154) );
    nor2_1 U40 ( .x(n37), .a(n35), .b(n38) );
    nand2i_2 U41 ( .x(n38), .a(B[26]), .b(A[26]) );
    nor2_1 U42 ( .x(n34), .a(n35), .b(n36) );
    nand2i_2 U43 ( .x(n36), .a(B[25]), .b(A[25]) );
    nand2i_2 U44 ( .x(n152), .a(B[31]), .b(A[31]) );
    nand2i_2 U45 ( .x(n101), .a(B[28]), .b(A[28]) );
    nor2_1 U46 ( .x(n48), .a(n35), .b(n49) );
    nand4i_1 U47 ( .x(n35), .a(n40), .b(n57), .c(n58), .d(n16) );
    nand2i_2 U48 ( .x(n49), .a(n21), .b(A[27]) );
    nor2i_1 U49 ( .x(n103), .a(A[29]), .b(B[29]) );
    inv_2 U50 ( .x(n54), .a(B[31]) );
    nor2i_1 U51 ( .x(n102), .a(A[30]), .b(n19) );
    nor2i_1 U52 ( .x(n106), .a(A[23]), .b(B[23]) );
    aoi211_1 U53 ( .x(n135), .a(n128), .b(n136), .c(n137), .d(n32) );
    oai22_1 U54 ( .x(n137), .a(A[22]), .b(n95), .c(n33), .d(n129) );
    inv_0 U55 ( .x(n95), .a(B[22]) );
    nor3i_1 U56 ( .x(n32), .a(n15), .b(n29), .c(n33) );
    aoi22_1 U57 ( .x(n130), .a(n108), .b(n131), .c(n111), .d(n109) );
    nor2i_1 U58 ( .x(n111), .a(n18), .b(n112) );
    inv_2 U59 ( .x(n112), .a(n158) );
    nand2i_2 U6 ( .x(n47), .a(n115), .b(n76) );
    nor2i_1 U60 ( .x(n109), .a(n79), .b(n110) );
    inv_0 U61 ( .x(n79), .a(A[20]) );
    inv_2 U62 ( .x(n110), .a(n131) );
    inv_2 U63 ( .x(n85), .a(A[1]) );
    nand3_1 U64 ( .x(n118), .a(n119), .b(n85), .c(B[1]) );
    oai22_1 U65 ( .x(n124), .a(A[3]), .b(n92), .c(A[2]), .d(n87) );
    inv_2 U66 ( .x(n119), .a(n27) );
    inv_2 U67 ( .x(n83), .a(A[4]) );
    inv_2 U68 ( .x(n123), .a(n86) );
    nand3_1 U69 ( .x(n122), .a(n123), .b(n119), .c(n124) );
    inv_0 U7 ( .x(n30), .a(A[15]) );
    inv_2 U70 ( .x(n156), .a(n157) );
    inv_2 U71 ( .x(n87), .a(B[2]) );
    nand2i_2 U72 ( .x(n125), .a(A[4]), .b(B[4]) );
    nand2i_2 U73 ( .x(n126), .a(n125), .b(n119) );
    nand2i_2 U74 ( .x(n59), .a(n60), .b(n61) );
    inv_2 U75 ( .x(n56), .a(B[25]) );
    inv_2 U76 ( .x(n55), .a(B[24]) );
    inv_2 U77 ( .x(n72), .a(B[9]) );
    inv_0 U78 ( .x(n69), .a(A[9]) );
    oai22_1 U79 ( .x(n46), .a(B[10]), .b(n70), .c(B[9]), .d(n69) );
    aoi22_1 U8 ( .x(n29), .a(B[15]), .b(n30), .c(B[14]), .d(n31) );
    inv_4 U80 ( .x(n99), .a(n46) );
    inv_2 U81 ( .x(n64), .a(B[12]) );
    nor2_1 U82 ( .x(n141), .a(n41), .b(n139) );
    oai21_1 U83 ( .x(n139), .a(n33), .b(n97), .c(n140) );
    inv_0 U84 ( .x(n26), .a(A[7]) );
    nand2i_2 U85 ( .x(n143), .a(n98), .b(n136) );
    inv_2 U86 ( .x(n136), .a(n33) );
    nand4_1 U87 ( .x(n52), .a(n148), .b(n149), .c(n150), .d(n151) );
    aoi222_1 U88 ( .x(n148), .a(n106), .b(n147), .c(n102), .d(n16), .e(n103), 
        .f(n16) );
    nand2i_2 U89 ( .x(n149), .a(n107), .b(n147) );
    inv_2 U9 ( .x(n94), .a(B[17]) );
    aoi21_1 U90 ( .x(n150), .a(n153), .b(n61), .c(n48) );
    inv_2 U91 ( .x(n153), .a(n101) );
    inv_2 U92 ( .x(n61), .a(n35) );
    nor3i_1 U93 ( .x(n151), .a(n152), .b(n34), .c(n37) );
    nor3_1 U94 ( .x(n51), .a(n134), .b(n132), .c(n138) );
    inv_2 U95 ( .x(n133), .a(n121) );
    inv_2 U96 ( .x(n147), .a(n59) );
    inv_5 U97 ( .x(n23), .a(n42) );
    ao222_2 U98 ( .x(n145), .a(n23), .b(n22), .c(n68), .d(n23), .e(n23), .f(
        n74) );
    oa22_1 U99 ( .x(n15), .a(B[15]), .b(n30), .c(B[16]), .d(n63) );
endmodule


module EX_DW01_cmp2_32_5_test_1 ( A, B, LEQ, TC, LT_LE, GE_GT );
input  [31:0] A;
input  [31:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n75, n136, n105, n137, n21, n88, n22, n67, n65, n103, n99, n42, n19, 
        n66, n68, n64, n86, n24, n123, n89, n94, n58, n140, n57, n56, n31, n26, 
        n128, n129, n139, n91, n90, n34, n33, n131, n47, n18, n48, n49, n50, 
        n100, n122, n40, n53, n63, n27, n25, n36, n15, n37, n38, n44, n76, n77, 
        n81, n82, n83, n84, n96, n101, n102, n106, n72, n110, n111, n112, n113, 
        n114, n115, n116, n74, n97, n95, n85, n87, n61, n70, n23, n73, n71, 
        n55, n54, n29, n28, n30, n120, n109, n92, n108, n107, n35, n104, n62, 
        n32, n20, n69, n117, n17, n93, n98, n135, n127, n46, n126, n141, n125, 
        n121, n119, n138, n124, n45, n41, n16, n60, n39, n78, n80, n52, n79, 
        n43, n132, n133, n134, n59, n118, n130, n51;
    nand3_1 U10 ( .x(n75), .a(n136), .b(n105), .c(n137) );
    inv_2 U100 ( .x(n21), .a(n88) );
    inv_2 U101 ( .x(n22), .a(A[28]) );
    aoi22_1 U102 ( .x(n67), .a(A[19]), .b(n65), .c(n103), .d(n99) );
    nand4i_4 U103 ( .x(n42), .a(n19), .b(n66), .c(n67), .d(n68) );
    inv_0 U104 ( .x(n64), .a(B[17]) );
    nand2_0 U105 ( .x(n86), .a(n24), .b(A[3]) );
    oai22_1 U106 ( .x(n123), .a(B[30]), .b(n88), .c(B[29]), .d(n89) );
    inv_0 U107 ( .x(n94), .a(A[6]) );
    inv_0 U108 ( .x(n58), .a(B[20]) );
    oai22_1 U109 ( .x(n140), .a(A[9]), .b(n57), .c(A[8]), .d(n56) );
    nor2i_0 U110 ( .x(n31), .a(A[8]), .b(B[8]) );
    aoi22_1 U111 ( .x(n26), .a(A[0]), .b(n128), .c(n129), .d(n128) );
    nand2i_2 U112 ( .x(n66), .a(B[22]), .b(A[22]) );
    oai22_1 U113 ( .x(n139), .a(B[11]), .b(n91), .c(B[12]), .d(n90) );
    nor2i_0 U114 ( .x(n34), .a(B[11]), .b(A[11]) );
    nor2i_0 U115 ( .x(n33), .a(B[3]), .b(A[3]) );
    inv_0 U116 ( .x(n131), .a(B[0]) );
    aoi221_1 U117 ( .x(n47), .a(n18), .b(n48), .c(A[7]), .d(n49), .e(n50) );
    nand2i_2 U118 ( .x(n100), .a(A[18]), .b(B[18]) );
    inv_0 U119 ( .x(n57), .a(B[9]) );
    inv_2 U12 ( .x(n122), .a(n136) );
    aoi22_1 U120 ( .x(n40), .a(A[13]), .b(n53), .c(A[14]), .d(n63) );
    and3i_3 U121 ( .x(LT_LE), .a(n27), .b(n25), .c(n26) );
    aoi21_3 U122 ( .x(n36), .a(n15), .b(n37), .c(n38) );
    oai211_4 U123 ( .x(n44), .a(n36), .b(n42), .c(n76), .d(n77) );
    nand4i_4 U124 ( .x(n81), .a(n82), .b(n83), .c(n18), .d(n84) );
    nor2i_5 U125 ( .x(n96), .a(B[21]), .b(A[21]) );
    nand4_1 U126 ( .x(n38), .a(n99), .b(n100), .c(n101), .d(n102) );
    nand2i_4 U127 ( .x(n106), .a(A[27]), .b(B[27]) );
    and4i_5 U128 ( .x(n77), .a(n72), .b(n110), .c(n111), .d(n112) );
    nand4_1 U129 ( .x(n82), .a(n113), .b(n114), .c(n115), .d(n116) );
    nand2i_2 U13 ( .x(n74), .a(n106), .b(n137) );
    nand2i_4 U130 ( .x(n97), .a(B[21]), .b(A[21]) );
    nand4_1 U131 ( .x(n113), .a(n95), .b(n85), .c(n86), .d(n87) );
    inv_10 U132 ( .x(n61), .a(A[15]) );
    nand2i_6 U133 ( .x(n136), .a(B[27]), .b(A[27]) );
    inv_3 U134 ( .x(n70), .a(B[28]) );
    nand2i_1 U135 ( .x(n137), .a(B[28]), .b(n23) );
    nor2i_0 U136 ( .x(n105), .a(B[26]), .b(A[26]) );
    nand2i_0 U137 ( .x(n110), .a(A[24]), .b(B[24]) );
    oai22_1 U15 ( .x(n73), .a(A[29]), .b(n71), .c(n23), .d(n70) );
    inv_0 U16 ( .x(n71), .a(B[29]) );
    inv_2 U17 ( .x(n23), .a(n22) );
    inv_2 U18 ( .x(n90), .a(A[12]) );
    inv_2 U19 ( .x(n91), .a(A[11]) );
    inv_2 U20 ( .x(n55), .a(A[9]) );
    inv_2 U21 ( .x(n54), .a(A[10]) );
    nand2i_1 U22 ( .x(n29), .a(n58), .b(n97) );
    nor3_1 U23 ( .x(n28), .a(n29), .b(A[20]), .c(n30) );
    nand2i_2 U24 ( .x(n120), .a(A[25]), .b(B[25]) );
    inv_2 U25 ( .x(n109), .a(n120) );
    inv_2 U26 ( .x(n92), .a(A[23]) );
    aoi21_1 U27 ( .x(n108), .a(B[23]), .b(n92), .c(n109) );
    aoi21_1 U28 ( .x(n107), .a(n96), .b(n66), .c(n35) );
    nor2i_0 U29 ( .x(n35), .a(B[22]), .b(A[22]) );
    nand4_1 U30 ( .x(n68), .a(n100), .b(n64), .c(n99), .d(A[17]) );
    nor2i_1 U31 ( .x(n103), .a(A[18]), .b(B[18]) );
    inv_2 U32 ( .x(n30), .a(n66) );
    inv_2 U33 ( .x(n104), .a(n97) );
    nand2i_0 U34 ( .x(n102), .a(A[16]), .b(B[16]) );
    nand2i_0 U35 ( .x(n101), .a(A[17]), .b(B[17]) );
    nand2i_2 U36 ( .x(n99), .a(A[19]), .b(B[19]) );
    oai22_1 U37 ( .x(n37), .a(A[14]), .b(n63), .c(A[15]), .d(n62) );
    nor2i_0 U38 ( .x(n32), .a(B[2]), .b(A[2]) );
    nor2i_1 U39 ( .x(n95), .a(n20), .b(A[1]) );
    inv_0 U40 ( .x(n69), .a(B[26]) );
    nand2i_0 U41 ( .x(n87), .a(B[2]), .b(A[2]) );
    nand2i_0 U42 ( .x(n117), .a(n20), .b(A[1]) );
    nand2i_2 U43 ( .x(n50), .a(n31), .b(n17) );
    inv_0 U44 ( .x(n93), .a(A[5]) );
    oai22_1 U45 ( .x(n48), .a(B[6]), .b(n94), .c(B[5]), .d(n93) );
    nand2_2 U46 ( .x(n112), .a(n98), .b(n135) );
    nand2i_2 U47 ( .x(n111), .a(A[31]), .b(B[31]) );
    inv_2 U48 ( .x(n127), .a(n111) );
    nand2i_2 U49 ( .x(n46), .a(n127), .b(n112) );
    inv_2 U50 ( .x(n89), .a(A[29]) );
    inv_2 U51 ( .x(n88), .a(A[30]) );
    nand2i_2 U52 ( .x(n135), .a(B[31]), .b(A[31]) );
    inv_2 U53 ( .x(n126), .a(n135) );
    inv_2 U54 ( .x(n141), .a(n137) );
    nand4i_1 U55 ( .x(n125), .a(n141), .b(n121), .c(n119), .d(n138) );
    nand3i_1 U56 ( .x(n72), .a(n73), .b(n74), .c(n75) );
    inv_2 U57 ( .x(n124), .a(n72) );
    aoi211_1 U58 ( .x(n45), .a(n124), .b(n125), .c(n126), .d(n123) );
    nand2_0 U59 ( .x(n41), .a(n16), .b(n139) );
    nor2i_0 U6 ( .x(n98), .a(B[30]), .b(n21) );
    inv_2 U60 ( .x(n60), .a(A[16]) );
    oa22_1 U61 ( .x(n15), .a(B[15]), .b(n61), .c(B[16]), .d(n60) );
    and4i_1 U62 ( .x(n39), .a(n42), .b(n15), .c(n40), .d(n41) );
    inv_2 U63 ( .x(n84), .a(n78) );
    nand2i_0 U64 ( .x(n80), .a(A[10]), .b(B[10]) );
    inv_0 U65 ( .x(n52), .a(B[12]) );
    nand2_2 U66 ( .x(n79), .a(n17), .b(n140) );
    nand4i_1 U67 ( .x(n78), .a(n34), .b(n79), .c(n16), .d(n80) );
    and3i_1 U68 ( .x(n76), .a(n28), .b(n107), .c(n108) );
    inv_5 U69 ( .x(n83), .a(n44) );
    nand4i_1 U7 ( .x(n138), .a(B[23]), .b(n120), .c(A[23]), .d(n110) );
    oai211_1 U70 ( .x(n116), .a(n32), .b(n33), .c(n86), .d(n85) );
    nand2i_0 U71 ( .x(n115), .a(A[4]), .b(B[4]) );
    nand2i_0 U72 ( .x(n114), .a(A[5]), .b(B[5]) );
    nand4i_1 U73 ( .x(n27), .a(n43), .b(n132), .c(n133), .d(n134) );
    oaoi211_1 U74 ( .x(n43), .a(n39), .b(n44), .c(n45), .d(n46) );
    or3i_2 U75 ( .x(n132), .a(n83), .b(n78), .c(n47) );
    nand2i_2 U76 ( .x(n133), .a(n117), .b(n128) );
    inv_5 U77 ( .x(n128), .a(n81) );
    nand2i_2 U78 ( .x(n134), .a(n87), .b(n128) );
    inv_2 U79 ( .x(n129), .a(n85) );
    aoi22_1 U8 ( .x(n119), .a(A[25]), .b(n59), .c(n118), .d(n120) );
    nand2i_2 U80 ( .x(n85), .a(B[4]), .b(A[4]) );
    aoi22_1 U81 ( .x(n25), .a(n130), .b(n128), .c(n128), .d(n131) );
    inv_2 U82 ( .x(n130), .a(n86) );
    inv_0 U83 ( .x(n53), .a(B[13]) );
    inv_2 U84 ( .x(n59), .a(B[25]) );
    inv_2 U85 ( .x(n49), .a(B[7]) );
    inv_0 U86 ( .x(n65), .a(B[19]) );
    inv_0 U87 ( .x(n63), .a(B[14]) );
    inv_0 U88 ( .x(n56), .a(B[8]) );
    inv_0 U89 ( .x(n51), .a(B[6]) );
    aoi21_1 U9 ( .x(n121), .a(A[26]), .b(n69), .c(n122) );
    oa22_3 U91 ( .x(n16), .a(A[13]), .b(n53), .c(A[12]), .d(n52) );
    oa22_1 U92 ( .x(n17), .a(B[9]), .b(n55), .c(B[10]), .d(n54) );
    oa22_1 U93 ( .x(n18), .a(A[6]), .b(n51), .c(A[7]), .d(n49) );
    ao21_3 U94 ( .x(n19), .a(A[20]), .b(n58), .c(n104) );
    inv_2 U95 ( .x(n62), .a(B[15]) );
    nor2i_1 U96 ( .x(n118), .a(A[24]), .b(B[24]) );
    buf_3 U98 ( .x(n20), .a(B[1]) );
    inv_2 U99 ( .x(n24), .a(B[3]) );
endmodule


module EX_DW01_cmp2_32_2 ( A, B, LEQ, TC, LT_LE, GE_GT );
input  [31:0] A;
input  [31:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n18, n48, n68, n129, n95, n125, n34, n100, n24, n39, n38, n17, n76, 
        n72, n71, n108, n67, n42, n66, n117, n93, n118, n41, n43, n90, n119, 
        n121, n92, n91, n89, n73, n105, n106, n107, n22, n140, n131, n97, n40, 
        n96, n55, n59, n56, n57, n58, n47, n74, n75, n86, n87, n88, n32, n98, 
        n99, n16, n132, n133, n15, n61, n135, n136, n134, n137, n120, n122, 
        n35, n94, n31, n25, n126, n127, n26, n27, n30, n142, n29, n23, n141, 
        n80, n79, n84, n116, n49, n46, n50, n83, n115, n112, n54, n113, n70, 
        n114, n103, n109, n111, n110, n77, n124, n123, n53, n44, n52, n102, 
        n62, n63, n64, n101, n85, n128, n130, n28, n33, n36, n45, n37, n19, 
        n20, n21, n81, n139, n82, n104, n51, n60, n69, n65, n78, n138;
    inv_2 U10 ( .x(n18), .a(A[23]) );
    nand2i_2 U100 ( .x(n48), .a(A[24]), .b(B[24]) );
    inv_0 U101 ( .x(n68), .a(B[17]) );
    nor2i_0 U102 ( .x(n129), .a(B[5]), .b(A[5]) );
    inv_0 U103 ( .x(n95), .a(A[0]) );
    nand2i_0 U104 ( .x(n125), .a(B[3]), .b(A[3]) );
    nand2i_0 U105 ( .x(n34), .a(A[3]), .b(B[3]) );
    nand2i_0 U106 ( .x(n100), .a(B[7]), .b(A[7]) );
    nor2i_0 U107 ( .x(n24), .a(A[8]), .b(B[8]) );
    nand2i_0 U108 ( .x(n39), .a(A[8]), .b(B[8]) );
    inv_0 U109 ( .x(n38), .a(B[9]) );
    inv_2 U11 ( .x(n17), .a(A[25]) );
    oai22_1 U110 ( .x(n76), .a(B[22]), .b(n72), .c(B[21]), .d(n71) );
    nor2i_0 U111 ( .x(n108), .a(B[21]), .b(A[21]) );
    oai22_1 U112 ( .x(n67), .a(B[15]), .b(n42), .c(B[16]), .d(n66) );
    aoi22_1 U113 ( .x(n117), .a(B[16]), .b(n66), .c(B[17]), .d(n93) );
    nand2i_0 U114 ( .x(n118), .a(B[14]), .b(A[14]) );
    aoi22_1 U115 ( .x(n41), .a(B[15]), .b(n42), .c(B[14]), .d(n43) );
    inv_0 U116 ( .x(n90), .a(B[13]) );
    nand2i_0 U117 ( .x(n119), .a(B[13]), .b(A[13]) );
    oai22_1 U118 ( .x(n121), .a(B[11]), .b(n92), .c(B[12]), .d(n91) );
    inv_0 U119 ( .x(n89), .a(B[12]) );
    nand3_2 U12 ( .x(n73), .a(n105), .b(n106), .c(n107) );
    nor2i_0 U120 ( .x(n22), .a(A[6]), .b(B[6]) );
    nand2i_0 U121 ( .x(n140), .a(A[6]), .b(B[6]) );
    aoi22_1 U122 ( .x(n131), .a(B[10]), .b(n97), .c(B[11]), .d(n92) );
    oai22_1 U123 ( .x(n40), .a(B[10]), .b(n97), .c(B[9]), .d(n96) );
    and4i_4 U124 ( .x(n55), .a(n59), .b(n56), .c(n57), .d(n58) );
    nand3i_5 U125 ( .x(n47), .a(n73), .b(n74), .c(n75) );
    nand2i_4 U126 ( .x(n86), .a(n87), .b(n88) );
    nand4i_4 U127 ( .x(n32), .a(n24), .b(n98), .c(n99), .d(n100) );
    oai211_4 U128 ( .x(n87), .a(n41), .b(n67), .c(n117), .d(n16) );
    nand2i_4 U129 ( .x(n59), .a(n132), .b(n133) );
    nand2i_2 U13 ( .x(n106), .a(B[26]), .b(A[26]) );
    nand2_2 U130 ( .x(n132), .a(n15), .b(n131) );
    nand4_1 U131 ( .x(n61), .a(n135), .b(n136), .c(n134), .d(n137) );
    nand2i_4 U132 ( .x(n136), .a(n119), .b(n133) );
    nand2i_4 U133 ( .x(n135), .a(n120), .b(n133) );
    nand2i_6 U134 ( .x(n105), .a(B[27]), .b(A[27]) );
    nand2i_2 U14 ( .x(n107), .a(B[28]), .b(A[28]) );
    nand2i_2 U15 ( .x(n122), .a(B[18]), .b(A[18]) );
    inv_2 U16 ( .x(n91), .a(A[12]) );
    inv_2 U17 ( .x(n92), .a(A[11]) );
    nand3_1 U18 ( .x(n35), .a(n125), .b(n94), .c(B[2]) );
    inv_2 U19 ( .x(n94), .a(A[2]) );
    and4i_1 U20 ( .x(n31), .a(n25), .b(n125), .c(n126), .d(n127) );
    nand2i_2 U21 ( .x(n126), .a(B[2]), .b(A[2]) );
    nand2i_0 U22 ( .x(n127), .a(B[4]), .b(A[4]) );
    nor2i_1 U23 ( .x(n25), .a(n26), .b(n27) );
    inv_2 U24 ( .x(n26), .a(B[0]) );
    nand2i_2 U25 ( .x(n30), .a(n95), .b(n142) );
    nand2i_2 U26 ( .x(n142), .a(A[1]), .b(B[1]) );
    inv_2 U27 ( .x(n27), .a(n142) );
    nand2i_2 U28 ( .x(n29), .a(B[1]), .b(A[1]) );
    inv_2 U29 ( .x(n97), .a(A[10]) );
    inv_2 U30 ( .x(n96), .a(A[9]) );
    nor2i_1 U31 ( .x(n23), .a(A[5]), .b(B[5]) );
    oai211_1 U32 ( .x(n98), .a(n22), .b(n23), .c(n140), .d(n141) );
    inv_2 U33 ( .x(n80), .a(B[19]) );
    inv_2 U34 ( .x(n79), .a(B[18]) );
    inv_2 U35 ( .x(n93), .a(A[17]) );
    inv_2 U36 ( .x(n43), .a(A[14]) );
    nor3i_1 U37 ( .x(n84), .a(n116), .b(n49), .c(n46) );
    nor2_0 U38 ( .x(n49), .a(n47), .b(n50) );
    nor2_0 U39 ( .x(n46), .a(n47), .b(n48) );
    aoi21_1 U40 ( .x(n83), .a(n108), .b(n115), .c(n112) );
    inv_2 U41 ( .x(n115), .a(n54) );
    oai33_1 U42 ( .x(n112), .a(n113), .b(A[27]), .c(n70), .d(n113), .e(n114), 
        .f(n103) );
    inv_2 U43 ( .x(n113), .a(n107) );
    inv_2 U44 ( .x(n70), .a(B[27]) );
    nor2i_1 U45 ( .x(n109), .a(B[20]), .b(A[20]) );
    nor2i_1 U46 ( .x(n111), .a(B[23]), .b(A[23]) );
    nor2i_1 U47 ( .x(n110), .a(B[22]), .b(A[22]) );
    inv_0 U48 ( .x(n71), .a(A[21]) );
    inv_0 U49 ( .x(n72), .a(A[22]) );
    nand2i_2 U50 ( .x(n54), .a(n76), .b(n77) );
    nand3_1 U51 ( .x(n124), .a(n16), .b(n68), .c(A[17]) );
    nand2i_2 U52 ( .x(n123), .a(n122), .b(n16) );
    nand3i_1 U53 ( .x(n53), .a(n44), .b(n123), .c(n124) );
    nand2i_2 U54 ( .x(n52), .a(B[20]), .b(A[20]) );
    nand2i_2 U55 ( .x(n137), .a(n118), .b(n133) );
    nor2i_1 U56 ( .x(n102), .a(A[30]), .b(B[30]) );
    inv_2 U57 ( .x(n62), .a(B[30]) );
    inv_2 U58 ( .x(n63), .a(B[31]) );
    oai22_1 U59 ( .x(n64), .a(A[31]), .b(n63), .c(A[30]), .d(n62) );
    nand2i_2 U6 ( .x(n103), .a(A[26]), .b(B[26]) );
    nor2i_1 U60 ( .x(n101), .a(A[29]), .b(B[29]) );
    aoi22_1 U61 ( .x(n134), .a(n101), .b(n85), .c(n102), .d(n85) );
    nand2_2 U62 ( .x(n120), .a(n15), .b(n121) );
    aoi211_1 U63 ( .x(n58), .a(n128), .b(n130), .c(n28), .d(n33) );
    nor2i_1 U64 ( .x(n128), .a(B[4]), .b(A[4]) );
    inv_2 U65 ( .x(n130), .a(n32) );
    inv_2 U66 ( .x(n99), .a(n40) );
    and4i_1 U67 ( .x(n28), .a(n32), .b(n29), .c(n30), .d(n31) );
    aoi211_1 U68 ( .x(n33), .a(n34), .b(n35), .c(n36), .d(n32) );
    inv_2 U69 ( .x(n36), .a(n127) );
    nor2i_2 U7 ( .x(n45), .a(A[25]), .b(B[25]) );
    oaoi211_1 U70 ( .x(n37), .a(A[9]), .b(n38), .c(n39), .d(n40) );
    aoi21_1 U71 ( .x(n57), .a(n129), .b(n130), .c(n37) );
    nand2i_2 U72 ( .x(n56), .a(n19), .b(n130) );
    nor2_1 U73 ( .x(n19), .a(n20), .b(n21) );
    inv_2 U74 ( .x(n20), .a(n140) );
    inv_2 U75 ( .x(n21), .a(n141) );
    inv_4 U76 ( .x(n88), .a(n81) );
    nand2i_2 U77 ( .x(n139), .a(B[31]), .b(A[31]) );
    inv_2 U78 ( .x(n85), .a(n64) );
    nand4_1 U79 ( .x(n81), .a(n82), .b(n83), .c(n84), .d(n85) );
    nor2i_1 U8 ( .x(n104), .a(A[24]), .b(B[24]) );
    nor3i_1 U80 ( .x(n51), .a(n52), .b(n53), .c(n54) );
    inv_2 U81 ( .x(n66), .a(A[16]) );
    inv_0 U82 ( .x(n42), .a(A[15]) );
    nor3i_2 U83 ( .x(LT_LE), .a(n60), .b(n55), .c(n61) );
    inv_5 U84 ( .x(n133), .a(n86) );
    oa22_1 U85 ( .x(n15), .a(A[13]), .b(n90), .c(A[12]), .d(n89) );
    oa22_2 U86 ( .x(n16), .a(A[19]), .b(n80), .c(A[18]), .d(n79) );
    inv_2 U87 ( .x(n69), .a(A[28]) );
    aoi22_1 U88 ( .x(n116), .a(B[28]), .b(n69), .c(n65), .d(B[29]) );
    inv_2 U89 ( .x(n65), .a(A[29]) );
    aoi21_1 U9 ( .x(n75), .a(n104), .b(n50), .c(n45) );
    inv_0 U90 ( .x(n114), .a(n105) );
    nand4i_1 U91 ( .x(n74), .a(n18), .b(n50), .c(n48), .d(n78) );
    inv_5 U92 ( .x(n78), .a(B[23]) );
    inv_7 U93 ( .x(n77), .a(n47) );
    nor2i_1 U94 ( .x(n44), .a(A[19]), .b(B[19]) );
    oai21_1 U95 ( .x(n138), .a(n51), .b(n81), .c(n139) );
    nand2i_0 U96 ( .x(n141), .a(A[7]), .b(B[7]) );
    aoi21_3 U97 ( .x(n60), .a(n133), .b(n67), .c(n138) );
    nand2_5 U98 ( .x(n50), .a(n17), .b(B[25]) );
    aoi222_1 U99 ( .x(n82), .a(n109), .b(n115), .c(n111), .d(n77), .e(n110), 
        .f(n77) );
endmodule


module EX_DW01_cmp2_32_4_test_1 ( A, B, LEQ, TC, LT_LE, GE_GT );
input  [31:0] A;
input  [31:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n116, n59, n115, n117, n27, n16, n47, n17, n18, n84, n23, n24, n25, 
        n97, n61, n120, n85, n119, n131, n26, n28, n21, n141, n55, n54, n29, 
        n19, n147, n44, n94, n135, n87, n86, n76, n91, n40, n49, n118, n64, 
        n77, n43, n42, n37, n56, n32, n53, n52, n111, n50, n20, n31, n33, n34, 
        n98, n99, n101, n74, n106, n67, n110, n92, n140, n35, n128, n129, n82, 
        n72, n145, n108, n107, n109, n68, n69, n70, n66, n144, n132, n148, n79, 
        n80, n81, n39, n71, n73, n38, n65, n100, n134, n123, n133, n113, n41, 
        n45, n46, n51, n75, n137, n30, n130, n96, n114, n63, n62, n142, n143, 
        n60, n22, n105, n104, n103, n88, n102, n57, n58, n124, n122, n121, 
        n112, n136, n15, n146, n126, n125, n89, n90, n139, n36, n138, n95, n93, 
        n48, n83;
    aoi22_1 U10 ( .x(n116), .a(A[25]), .b(n59), .c(n115), .d(n117) );
    inv_2 U101 ( .x(n27), .a(A[20]) );
    inv_2 U102 ( .x(n16), .a(n47) );
    inv_2 U103 ( .x(n47), .a(B[1]) );
    buf_3 U104 ( .x(n17), .a(B[3]) );
    inv_2 U105 ( .x(n18), .a(n84) );
    inv_2 U106 ( .x(n84), .a(A[30]) );
    oai22_1 U107 ( .x(n23), .a(B[17]), .b(n24), .c(B[18]), .d(n25) );
    aoi22_1 U108 ( .x(n97), .a(B[16]), .b(n61), .c(B[17]), .d(n24) );
    oai22_1 U109 ( .x(n120), .a(B[30]), .b(n84), .c(B[29]), .d(n85) );
    inv_2 U11 ( .x(n119), .a(n131) );
    aoi22_1 U110 ( .x(n26), .a(B[20]), .b(n27), .c(B[21]), .d(n28) );
    nor2i_2 U111 ( .x(n21), .a(A[20]), .b(B[20]) );
    oai22_1 U112 ( .x(n141), .a(A[8]), .b(n55), .c(A[9]), .d(n54) );
    nor2i_0 U113 ( .x(n29), .a(A[8]), .b(B[8]) );
    ao222_3 U114 ( .x(n19), .a(A[0]), .b(n147), .c(n147), .d(n44), .e(n94), 
        .f(n147) );
    oai22_1 U115 ( .x(n135), .a(B[11]), .b(n87), .c(B[12]), .d(n86) );
    nand2i_0 U116 ( .x(n76), .a(A[11]), .b(B[11]) );
    nand2i_0 U117 ( .x(n91), .a(A[3]), .b(n17) );
    inv_0 U118 ( .x(n40), .a(A[3]) );
    inv_0 U119 ( .x(n49), .a(B[0]) );
    aoi21_1 U12 ( .x(n118), .a(A[26]), .b(n64), .c(n119) );
    oai22_1 U120 ( .x(n77), .a(A[6]), .b(n43), .c(A[7]), .d(n42) );
    aoi211_1 U121 ( .x(n37), .a(A[7]), .b(n42), .c(n29), .d(n56) );
    nand2i_2 U122 ( .x(n32), .a(A[18]), .b(B[18]) );
    oai22_1 U123 ( .x(n56), .a(B[10]), .b(n53), .c(B[9]), .d(n52) );
    inv_0 U124 ( .x(n54), .a(B[9]) );
    aoi21_1 U125 ( .x(n111), .a(A[13]), .b(n50), .c(n23) );
    nor2_5 U126 ( .x(LT_LE), .a(n19), .b(n20) );
    aoi21_6 U127 ( .x(n31), .a(n32), .b(n33), .c(n34) );
    nor2i_5 U128 ( .x(n98), .a(n99), .b(n34) );
    nand2i_4 U129 ( .x(n101), .a(A[27]), .b(B[27]) );
    nor3i_5 U130 ( .x(n74), .a(n106), .b(n67), .c(n31) );
    nand2i_4 U131 ( .x(n110), .a(n92), .b(n140) );
    nand3i_5 U132 ( .x(n20), .a(n35), .b(n128), .c(n129) );
    nand2i_6 U134 ( .x(n82), .a(B[2]), .b(A[2]) );
    nand2_4 U135 ( .x(n72), .a(n98), .b(n145) );
    nand3i_5 U136 ( .x(n108), .a(n107), .b(n109), .c(n110) );
    nand3i_5 U137 ( .x(n67), .a(n68), .b(n69), .c(n70) );
    nand2i_6 U138 ( .x(n131), .a(B[27]), .b(A[27]) );
    inv_0 U139 ( .x(n66), .a(B[29]) );
    inv_2 U14 ( .x(n144), .a(n132) );
    and4_5 U140 ( .x(n147), .a(n148), .b(n79), .c(n80), .d(n81) );
    inv_3 U141 ( .x(n148), .a(n39) );
    nand4i_2 U142 ( .x(n39), .a(n71), .b(n72), .c(n73), .d(n74) );
    nor2_2 U143 ( .x(n80), .a(n38), .b(n77) );
    nand2i_0 U144 ( .x(n132), .a(B[28]), .b(A[28]) );
    inv_0 U145 ( .x(n65), .a(B[28]) );
    nor2i_0 U146 ( .x(n100), .a(B[26]), .b(A[26]) );
    nand2i_4 U147 ( .x(n134), .a(A[24]), .b(B[24]) );
    nand4i_1 U15 ( .x(n123), .a(n144), .b(n118), .c(n116), .d(n133) );
    nand2i_2 U16 ( .x(n113), .a(B[14]), .b(A[14]) );
    inv_2 U17 ( .x(n86), .a(A[12]) );
    inv_2 U18 ( .x(n87), .a(A[11]) );
    nand2i_0 U19 ( .x(n92), .a(A[2]), .b(B[2]) );
    nand2i_2 U20 ( .x(n109), .a(n91), .b(n140) );
    inv_2 U21 ( .x(n140), .a(n44) );
    inv_2 U22 ( .x(n41), .a(A[4]) );
    inv_2 U23 ( .x(n45), .a(B[4]) );
    oai22_1 U24 ( .x(n107), .a(A[4]), .b(n45), .c(A[5]), .d(n46) );
    inv_0 U25 ( .x(n51), .a(B[12]) );
    nand2_2 U26 ( .x(n75), .a(n137), .b(n141) );
    nor2i_0 U27 ( .x(n30), .a(B[10]), .b(A[10]) );
    nand2i_2 U28 ( .x(n33), .a(A[19]), .b(B[19]) );
    nand3_1 U29 ( .x(n70), .a(n131), .b(n100), .c(n132) );
    nand2i_2 U30 ( .x(n69), .a(n101), .b(n132) );
    oai22_1 U32 ( .x(n68), .a(A[29]), .b(n66), .c(A[28]), .d(n65) );
    nand2i_2 U33 ( .x(n130), .a(B[31]), .b(A[31]) );
    nor2i_1 U34 ( .x(n96), .a(B[30]), .b(n18) );
    inv_0 U35 ( .x(n114), .a(n63) );
    inv_2 U36 ( .x(n61), .a(A[16]) );
    inv_5 U37 ( .x(n62), .a(A[15]) );
    oai22_1 U38 ( .x(n63), .a(B[15]), .b(n62), .c(B[16]), .d(n61) );
    nand2i_2 U39 ( .x(n142), .a(A[14]), .b(B[14]) );
    aoai211_1 U40 ( .x(n145), .a(n143), .b(n142), .c(n63), .d(n97) );
    or3i_2 U41 ( .x(n34), .a(n60), .b(n21), .c(n22) );
    inv_2 U42 ( .x(n25), .a(A[18]) );
    inv_2 U43 ( .x(n24), .a(A[17]) );
    inv_2 U44 ( .x(n99), .a(n23) );
    inv_2 U45 ( .x(n105), .a(n134) );
    nand2i_2 U46 ( .x(n117), .a(A[25]), .b(B[25]) );
    inv_2 U47 ( .x(n104), .a(n117) );
    nor2_1 U48 ( .x(n103), .a(n104), .b(n105) );
    inv_2 U49 ( .x(n88), .a(A[23]) );
    aoi22_1 U50 ( .x(n102), .a(B[23]), .b(n88), .c(B[22]), .d(n57) );
    oai22_1 U51 ( .x(n58), .a(B[21]), .b(n28), .c(B[22]), .d(n57) );
    inv_0 U52 ( .x(n28), .a(A[21]) );
    inv_2 U53 ( .x(n57), .a(A[22]) );
    inv_2 U54 ( .x(n60), .a(n58) );
    inv_0 U55 ( .x(n64), .a(B[26]) );
    inv_2 U56 ( .x(n124), .a(n130) );
    inv_2 U57 ( .x(n122), .a(n67) );
    aoi211_1 U58 ( .x(n121), .a(n122), .b(n123), .c(n124), .d(n120) );
    and4i_1 U59 ( .x(n112), .a(n34), .b(n113), .c(n114), .d(n111) );
    nand2_2 U60 ( .x(n136), .a(n15), .b(n135) );
    aoai211_1 U61 ( .x(n146), .a(n136), .b(n112), .c(n39), .d(n121) );
    nand2i_2 U62 ( .x(n106), .a(A[31]), .b(B[31]) );
    inv_2 U63 ( .x(n126), .a(n106) );
    nand2i_2 U64 ( .x(n125), .a(n126), .b(n73) );
    inv_0 U65 ( .x(n53), .a(A[10]) );
    inv_0 U66 ( .x(n52), .a(A[9]) );
    inv_2 U67 ( .x(n137), .a(n56) );
    inv_0 U68 ( .x(n89), .a(A[5]) );
    inv_0 U69 ( .x(n90), .a(A[6]) );
    nor2i_1 U7 ( .x(n22), .a(A[19]), .b(B[19]) );
    oai22_1 U70 ( .x(n139), .a(B[6]), .b(n90), .c(B[5]), .d(n89) );
    nand2_2 U71 ( .x(n36), .a(n138), .b(n139) );
    aoi21_2 U72 ( .x(n81), .a(n95), .b(n93), .c(n108) );
    nor2_1 U73 ( .x(n95), .a(n44), .b(n47) );
    nor2i_1 U74 ( .x(n93), .a(n48), .b(n94) );
    inv_2 U75 ( .x(n48), .a(A[1]) );
    inv_2 U76 ( .x(n138), .a(n77) );
    nand4i_1 U77 ( .x(n38), .a(n30), .b(n75), .c(n15), .d(n76) );
    nand2i_2 U79 ( .x(n83), .a(n16), .b(A[1]) );
    inv_2 U8 ( .x(n85), .a(A[29]) );
    nand4i_1 U80 ( .x(n79), .a(n49), .b(n140), .c(n83), .d(n82) );
    oai211_1 U82 ( .x(n71), .a(n26), .b(n58), .c(n102), .d(n103) );
    nand2_2 U83 ( .x(n73), .a(n96), .b(n130) );
    nand2i_2 U84 ( .x(n129), .a(n83), .b(n147) );
    nand2i_2 U85 ( .x(n128), .a(n125), .b(n146) );
    aoi211_1 U86 ( .x(n35), .a(n36), .b(n37), .c(n38), .d(n39) );
    inv_2 U87 ( .x(n94), .a(n82) );
    oai22_1 U88 ( .x(n44), .a(B[4]), .b(n41), .c(n17), .d(n40) );
    nand4i_1 U9 ( .x(n133), .a(B[23]), .b(n117), .c(A[23]), .d(n134) );
    inv_0 U90 ( .x(n50), .a(B[13]) );
    inv_0 U91 ( .x(n46), .a(B[5]) );
    inv_2 U92 ( .x(n59), .a(B[25]) );
    inv_2 U93 ( .x(n42), .a(B[7]) );
    inv_0 U94 ( .x(n55), .a(B[8]) );
    inv_0 U95 ( .x(n43), .a(B[6]) );
    oa22_2 U97 ( .x(n15), .a(A[12]), .b(n51), .c(A[13]), .d(n50) );
    nand2i_2 U98 ( .x(n143), .a(A[15]), .b(B[15]) );
    nor2i_1 U99 ( .x(n115), .a(A[24]), .b(B[24]) );
endmodule


module EX_DW01_cmp2_32_1 ( A, B, LEQ, TC, LT_LE, GE_GT );
input  [31:0] A;
input  [31:0] B;
input  LEQ, TC;
output LT_LE, GE_GT;
    wire n18, n85, n84, n81, n103, n109, n112, n87, n86, n88, n32, n106, n102, 
        n66, n67, n65, n60, n57, n56, n97, n27, n37, n35, n98, n71, n72, n25, 
        n104, n43, n111, n64, n33, n58, n93, n94, n95, n78, n63, n45, n46, n47, 
        n48, n49, n50, n51, n80, n79, n125, n135, n30, n105, n128, n108, n127, 
        n124, n121, n76, n26, n114, n70, n59, n17, n139, n140, n15, n34, n28, 
        n24, n36, n22, n23, n19, n61, n68, n101, n100, n89, n107, n31, n118, 
        n122, n123, n119, n55, n96, n75, n38, n39, n40, n16, n110, n130, n131, 
        n129, n83, n82, n134, n133, n54, n77, n42, n44, n113, n20, n29, n117, 
        n62, n115, n116, n73, n74, n69, n99, n91, n137, n138, n136, n90, n41, 
        n52, n53, n126, n132, n21, n92, n120;
    and4_3 U10 ( .x(n18), .a(A[23]), .b(n85), .c(n84), .d(n81) );
    nand2i_0 U100 ( .x(n103), .a(B[5]), .b(A[5]) );
    nand2i_0 U101 ( .x(n109), .a(A[5]), .b(B[5]) );
    oai22_1 U102 ( .x(n112), .a(A[9]), .b(n87), .c(A[8]), .d(n86) );
    inv_0 U103 ( .x(n88), .a(A[0]) );
    inv_0 U104 ( .x(n32), .a(A[3]) );
    nand2i_0 U105 ( .x(n106), .a(B[3]), .b(A[3]) );
    aoi22_1 U106 ( .x(n102), .a(A[7]), .b(n66), .c(A[8]), .d(n86) );
    oai22_1 U107 ( .x(n67), .a(A[7]), .b(n66), .c(A[6]), .d(n65) );
    inv_0 U108 ( .x(n86), .a(B[8]) );
    inv_0 U109 ( .x(n87), .a(B[9]) );
    inv_2 U11 ( .x(n81), .a(B[23]) );
    oai22_1 U110 ( .x(n60), .a(B[21]), .b(n57), .c(B[22]), .d(n56) );
    nand2i_0 U111 ( .x(n97), .a(A[21]), .b(B[21]) );
    inv_0 U112 ( .x(n27), .a(B[16]) );
    nor2i_0 U113 ( .x(n37), .a(B[16]), .b(A[16]) );
    inv_0 U114 ( .x(n35), .a(B[14]) );
    aoi22_1 U115 ( .x(n98), .a(A[13]), .b(n71), .c(A[14]), .d(n35) );
    oai22_1 U116 ( .x(n72), .a(A[13]), .b(n71), .c(A[12]), .d(n25) );
    nand2i_0 U117 ( .x(n104), .a(B[6]), .b(A[6]) );
    inv_0 U118 ( .x(n65), .a(B[6]) );
    aoi221_1 U119 ( .x(n43), .a(n111), .b(n112), .c(B[10]), .d(n64), .e(n33)
         );
    nand3_1 U12 ( .x(n58), .a(n93), .b(n94), .c(n95) );
    oai22_1 U120 ( .x(n78), .a(B[10]), .b(n64), .c(B[9]), .d(n63) );
    nor3i_5 U121 ( .x(n45), .a(n46), .b(n47), .c(n48) );
    aoi21_3 U122 ( .x(LT_LE), .a(n49), .b(n50), .c(n51) );
    or3i_5 U123 ( .x(n48), .a(n80), .b(n78), .c(n79) );
    or3i_4 U124 ( .x(n125), .a(n135), .b(n30), .c(n105) );
    nand2i_4 U125 ( .x(n128), .a(n108), .b(n135) );
    nand2i_4 U126 ( .x(n127), .a(n109), .b(n135) );
    inv_7 U127 ( .x(n135), .a(n48) );
    nand2i_5 U128 ( .x(n124), .a(n121), .b(n125) );
    nand2i_5 U129 ( .x(n76), .a(n26), .b(n114) );
    nand2i_2 U13 ( .x(n94), .a(B[26]), .b(A[26]) );
    inv_6 U130 ( .x(n114), .a(n70) );
    nand2i_5 U131 ( .x(n59), .a(n60), .b(n17) );
    inv_10 U132 ( .x(n57), .a(A[21]) );
    nand2i_2 U14 ( .x(n95), .a(B[28]), .b(A[28]) );
    nor2i_0 U15 ( .x(n33), .a(B[11]), .b(A[11]) );
    inv_0 U16 ( .x(n71), .a(B[13]) );
    nand2i_0 U17 ( .x(n139), .a(B[11]), .b(A[11]) );
    aoai211_1 U18 ( .x(n140), .a(n139), .b(n15), .c(n72), .d(n98) );
    oai22_1 U19 ( .x(n34), .a(A[14]), .b(n35), .c(A[15]), .d(n28) );
    inv_2 U20 ( .x(n24), .a(A[18]) );
    nor2i_1 U21 ( .x(n36), .a(B[17]), .b(A[17]) );
    or3i_2 U22 ( .x(n70), .a(n22), .b(n36), .c(n37) );
    inv_2 U23 ( .x(n28), .a(B[15]) );
    aoi22_1 U24 ( .x(n26), .a(A[16]), .b(n27), .c(A[15]), .d(n28) );
    inv_0 U25 ( .x(n56), .a(A[22]) );
    aoi22_1 U26 ( .x(n22), .a(n24), .b(B[18]), .c(n23), .d(B[19]) );
    inv_2 U27 ( .x(n23), .a(A[19]) );
    inv_2 U28 ( .x(n19), .a(A[20]) );
    inv_2 U29 ( .x(n61), .a(B[20]) );
    inv_0 U30 ( .x(n68), .a(B[19]) );
    nand2i_0 U31 ( .x(n101), .a(B[17]), .b(A[17]) );
    nand2i_2 U32 ( .x(n100), .a(B[18]), .b(A[18]) );
    nand2i_2 U33 ( .x(n89), .a(B[29]), .b(A[29]) );
    nand2_2 U34 ( .x(n105), .a(n106), .b(n107) );
    inv_2 U35 ( .x(n31), .a(A[2]) );
    aoi22_1 U36 ( .x(n30), .a(B[2]), .b(n31), .c(B[3]), .d(n32) );
    nand3i_1 U37 ( .x(n121), .a(n118), .b(n122), .c(n123) );
    inv_2 U38 ( .x(n119), .a(n95) );
    inv_2 U39 ( .x(n55), .a(B[27]) );
    nand2i_0 U40 ( .x(n122), .a(n96), .b(n75) );
    nand2i_0 U41 ( .x(n123), .a(n97), .b(n75) );
    nor2_1 U42 ( .x(n38), .a(n39), .b(n40) );
    nor3_2 U43 ( .x(n17), .a(n58), .b(n18), .c(n16) );
    nand2i_2 U44 ( .x(n40), .a(A[22]), .b(B[22]) );
    nor2i_1 U45 ( .x(n110), .a(B[23]), .b(A[23]) );
    nand2i_2 U46 ( .x(n108), .a(A[4]), .b(B[4]) );
    aoi21_1 U47 ( .x(n130), .a(n131), .b(n17), .c(n129) );
    inv_2 U48 ( .x(n131), .a(n84) );
    nand2i_2 U49 ( .x(n84), .a(A[24]), .b(B[24]) );
    oai22_1 U50 ( .x(n129), .a(A[29]), .b(n83), .c(A[28]), .d(n82) );
    inv_2 U51 ( .x(n83), .a(B[29]) );
    inv_2 U52 ( .x(n82), .a(B[28]) );
    nand2i_2 U53 ( .x(n85), .a(A[25]), .b(B[25]) );
    inv_2 U54 ( .x(n134), .a(n85) );
    aoi21_1 U55 ( .x(n133), .a(n134), .b(n17), .c(n54) );
    nand3i_2 U56 ( .x(n77), .a(n34), .b(n114), .c(n140) );
    nor2i_1 U57 ( .x(n42), .a(n43), .b(n44) );
    nand3i_0 U58 ( .x(n44), .a(n72), .b(n113), .c(n114) );
    inv_2 U59 ( .x(n113), .a(n34) );
    nand2i_2 U6 ( .x(n96), .a(n20), .b(B[20]) );
    oai31_2 U60 ( .x(n47), .a(n88), .b(B[0]), .c(n29), .d(n117) );
    nor2i_1 U61 ( .x(n29), .a(B[1]), .b(A[1]) );
    nand2i_2 U62 ( .x(n117), .a(B[1]), .b(A[1]) );
    aoi211_1 U63 ( .x(n46), .a(A[2]), .b(n62), .c(n115), .d(n116) );
    inv_2 U64 ( .x(n62), .a(B[2]) );
    inv_2 U65 ( .x(n115), .a(n107) );
    nand2i_2 U66 ( .x(n107), .a(B[4]), .b(A[4]) );
    inv_2 U67 ( .x(n116), .a(n106) );
    nand4i_1 U68 ( .x(n73), .a(n74), .b(n75), .c(n76), .d(n77) );
    aoai211_1 U69 ( .x(n74), .a(n100), .b(n101), .c(n69), .d(n99) );
    nand2i_2 U7 ( .x(n91), .a(A[26]), .b(B[26]) );
    inv_5 U70 ( .x(n75), .a(n59) );
    inv_2 U71 ( .x(n80), .a(n73) );
    aoai211_1 U72 ( .x(n79), .a(n103), .b(n104), .c(n67), .d(n102) );
    inv_0 U73 ( .x(n64), .a(A[10]) );
    inv_0 U74 ( .x(n63), .a(A[9]) );
    inv_2 U75 ( .x(n111), .a(n78) );
    nand2i_2 U76 ( .x(n137), .a(B[31]), .b(A[31]) );
    inv_2 U77 ( .x(n138), .a(n54) );
    nand2i_2 U78 ( .x(n136), .a(n89), .b(n138) );
    nand2i_2 U79 ( .x(n90), .a(B[30]), .b(A[30]) );
    nor2i_0 U8 ( .x(n41), .a(A[25]), .b(B[25]) );
    inv_2 U80 ( .x(n52), .a(B[30]) );
    inv_2 U81 ( .x(n53), .a(B[31]) );
    oai22_1 U82 ( .x(n54), .a(A[31]), .b(n53), .c(A[30]), .d(n52) );
    oai211_1 U83 ( .x(n51), .a(n54), .b(n90), .c(n136), .d(n137) );
    and4i_3 U84 ( .x(n50), .a(n124), .b(n127), .c(n128), .d(n126) );
    aoi21_1 U85 ( .x(n126), .a(n110), .b(n17), .c(n38) );
    aoi211_1 U86 ( .x(n49), .a(n135), .b(n67), .c(n45), .d(n132) );
    inv_0 U87 ( .x(n66), .a(B[7]) );
    oai211_1 U88 ( .x(n132), .a(n42), .b(n21), .c(n133), .d(n130) );
    nand2_2 U89 ( .x(n15), .a(n25), .b(A[12]) );
    nor2i_1 U9 ( .x(n92), .a(A[24]), .b(B[24]) );
    ao21_3 U90 ( .x(n16), .a(n92), .b(n85), .c(n41) );
    inv_0 U91 ( .x(n39), .a(n17) );
    oai33_1 U92 ( .x(n118), .a(n119), .b(A[27]), .c(n55), .d(n119), .e(n120), 
        .f(n91) );
    inv_0 U93 ( .x(n120), .a(n93) );
    nand2i_4 U94 ( .x(n93), .a(B[27]), .b(A[27]) );
    inv_2 U95 ( .x(n20), .a(n19) );
    nand4i_1 U96 ( .x(n21), .a(n74), .b(n75), .c(n76), .d(n77) );
    aoi22_1 U97 ( .x(n99), .a(n20), .b(n61), .c(A[19]), .d(n68) );
    inv_2 U98 ( .x(n69), .a(n22) );
    inv_0 U99 ( .x(n25), .a(B[12]) );
endmodule


module EX_DW01_sub_32_2_test_1 ( A, B, CI, DIFF, CO );
input  [31:0] A;
input  [31:0] B;
output [31:0] DIFF;
input  CI;
output CO;
    wire n191, n59, n218, n318, n214, n121, n51, n250, n171, n284, n169, n170, 
        n333, n173, n228, n82, n50, n141, n167, n168, n311, n200, n330, n79, 
        n80, n360, n329, n190, n192, n193, n194, n331, n255, n332, n328, n147, 
        n337, n300, n299, n257, n298, n148, n175, n247, n342, n304, n302, n240, 
        n303, n221, n153, n161, n352, n315, n154, n226, n159, n186, n276, n232, 
        n160, n246, n81, n277, n216, n125, n229, n177, n156, n157, n158, n223, 
        n230, n180, n209, n272, n172, n283, n174, n231, n183, n146, n270, n144, 
        n112, n217, n128, n162, n203, n88, n163, n131, n285, n249, n198, n310, 
        n195, n273, n347, n309, n344, n120, n245, n185, n275, n117, n164, n199, 
        n274, n210, n253, n139, n140, n271, n269, n225, n239, n224, n265, n113, 
        n237, n155, n115, n280, n233, n279, n281, n248, n84, n325, n118, n53, 
        n52, n263, n212, n213, n57, n110, n278, n267, n359, n346, n355, n54, 
        n98, n100, n99, n202, n254, n166, n65, n179, n142, n143, n90, n89, 
        n290, n291, n55, n313, n56, n296, n63, n288, n316, n259, n58, n64, 
        n241, n289, n219, n105, n266, n101, n358, n301, n102, n201, n295, n286, 
        n336, n258, n261, n242, n243, n138, n60, n287, n61, n321, n244, n66, 
        n62, n234, n181, n208, n292, n293, n294, n135, n357, n197, n97, n95, 
        n96, n297, n92, n256, n165, n312, n334, n67, n262, n68, n69, n308, n70, 
        n314, n75, n71, n222, n72, n74, n73, n76, n77, n345, n211, n264, n134, 
        n126, n127, n78, n252, n251, n85, n86, n189, n351, n350, n87, n93, 
        n260, n184, n91, n129, n322, n130, n326, n94, n109, n108, n356, n111, 
        n178, n364, n268, n338, n339, n340, n103, n104, n220, n215, n122, n196, 
        n204, n205, n206, n207, n335, n238, n343, n327, n319, n136, n137, n227, 
        n133, n305, n306, n307, n236, n124, n235, n317, n341, n361, n362, n363, 
        n149, n123, n114, n116, n348, n349, n188, n150, n187, n365, n83, n182, 
        n354, n176, n353, n324, n119, n145, n132, n151, n152, n323, n282, n320;
    inv_2 U10 ( .x(n191), .a(n59) );
    inv_2 U100 ( .x(n218), .a(n318) );
    oai21_1 U101 ( .x(n214), .a(n121), .b(n51), .c(n250) );
    inv_0 U102 ( .x(n171), .a(n284) );
    nor2_1 U103 ( .x(n169), .a(n170), .b(n171) );
    nand2i_2 U104 ( .x(n333), .a(B[14]), .b(A[14]) );
    inv_2 U105 ( .x(n173), .a(n333) );
    oai21_1 U106 ( .x(n228), .a(n82), .b(n50), .c(n141) );
    nor2_1 U107 ( .x(n167), .a(n168), .b(n311) );
    inv_2 U108 ( .x(n168), .a(n200) );
    inv_2 U109 ( .x(n311), .a(n330) );
    nor2_1 U110 ( .x(n79), .a(A[16]), .b(n80) );
    inv_2 U111 ( .x(n360), .a(n329) );
    aoi211_1 U112 ( .x(n190), .a(n191), .b(n192), .c(n193), .d(n194) );
    oai211_2 U113 ( .x(n331), .a(n190), .b(n255), .c(n332), .d(n328) );
    nand2i_2 U114 ( .x(n147), .a(B[21]), .b(A[21]) );
    inv_2 U115 ( .x(n337), .a(n147) );
    nand2i_2 U116 ( .x(n300), .a(B[21]), .b(n299) );
    inv_2 U117 ( .x(n257), .a(A[21]) );
    nand2i_2 U118 ( .x(n298), .a(n257), .b(n299) );
    nor2i_0 U119 ( .x(n148), .a(A[22]), .b(B[22]) );
    inv_5 U12 ( .x(n175), .a(n247) );
    nand2i_2 U120 ( .x(n342), .a(B[25]), .b(A[25]) );
    inv_2 U121 ( .x(n304), .a(n342) );
    inv_2 U122 ( .x(n302), .a(n240) );
    nand2i_2 U123 ( .x(n303), .a(A[25]), .b(B[25]) );
    exor2_1 U124 ( .x(DIFF[3]), .a(n221), .b(n153) );
    oai21_1 U125 ( .x(n221), .a(n161), .b(n352), .c(n315) );
    inv_2 U126 ( .x(n154), .a(B[3]) );
    exor2_1 U127 ( .x(DIFF[2]), .a(n226), .b(n159) );
    aoai211_1 U128 ( .x(n226), .a(B[1]), .b(n186), .c(n276), .d(n232) );
    nor2_1 U129 ( .x(n159), .a(n160), .b(n161) );
    inv_2 U13 ( .x(n246), .a(n81) );
    inv_2 U130 ( .x(n160), .a(n315) );
    inv_2 U131 ( .x(n161), .a(n277) );
    inv_2 U132 ( .x(n352), .a(n226) );
    exor2_1 U133 ( .x(DIFF[6]), .a(n216), .b(n125) );
    exor2_1 U134 ( .x(DIFF[12]), .a(n229), .b(n177) );
    nor2_1 U135 ( .x(n156), .a(n157), .b(n158) );
    exor2_1 U136 ( .x(DIFF[27]), .a(n223), .b(n156) );
    exor2_1 U137 ( .x(DIFF[11]), .a(n230), .b(n180) );
    exnor2_1 U138 ( .x(DIFF[20]), .a(n209), .b(n272) );
    exor2_1 U139 ( .x(DIFF[14]), .a(n228), .b(n172) );
    nor2i_1 U14 ( .x(n283), .a(n284), .b(n173) );
    exnor2_1 U140 ( .x(DIFF[13]), .a(n50), .b(n174) );
    exor2_1 U141 ( .x(DIFF[10]), .a(n231), .b(n183) );
    exnor2_1 U142 ( .x(DIFF[22]), .a(n146), .b(n270) );
    nor3i_1 U143 ( .x(n146), .a(n147), .b(n144), .c(n112) );
    exnor2_1 U144 ( .x(n270), .a(A[22]), .b(B[22]) );
    exor2_1 U145 ( .x(DIFF[5]), .a(n217), .b(n128) );
    exnor2_1 U146 ( .x(DIFF[19]), .a(n162), .b(n203) );
    nor2_0 U147 ( .x(n162), .a(n88), .b(n163) );
    inv_2 U148 ( .x(n163), .a(n328) );
    exnor2_1 U149 ( .x(DIFF[4]), .a(n218), .b(n131) );
    oai21_1 U15 ( .x(n285), .a(n246), .b(n249), .c(n283) );
    inv_2 U150 ( .x(n198), .a(n310) );
    exnor2_1 U151 ( .x(DIFF[18]), .a(n195), .b(n273) );
    inv_2 U152 ( .x(n347), .a(n309) );
    inv_2 U153 ( .x(n157), .a(n344) );
    exnor2_1 U154 ( .x(DIFF[8]), .a(n51), .b(n120) );
    inv_2 U155 ( .x(n121), .a(n245) );
    mux2i_1 U156 ( .x(DIFF[1]), .d0(n185), .sl(n276), .d1(n275) );
    exor2_1 U157 ( .x(DIFF[9]), .a(n214), .b(n117) );
    mux2i_1 U158 ( .x(DIFF[17]), .d0(n164), .sl(n199), .d1(n274) );
    inv_4 U159 ( .x(n210), .a(n253) );
    nor2_1 U16 ( .x(n139), .a(n140), .b(n141) );
    exnor2_1 U160 ( .x(n271), .a(A[21]), .b(B[21]) );
    exnor2_1 U161 ( .x(n269), .a(A[23]), .b(B[23]) );
    nand2_2 U162 ( .x(n225), .a(n303), .b(n342) );
    inv_2 U163 ( .x(n239), .a(A[24]) );
    exnor2_1 U164 ( .x(DIFF[25]), .a(n224), .b(n225) );
    exnor2_1 U165 ( .x(n265), .a(B[26]), .b(A[26]) );
    exnor2_1 U166 ( .x(DIFF[21]), .a(n113), .b(n271) );
    inv_2 U168 ( .x(n237), .a(B[28]) );
    inv_2 U169 ( .x(n155), .a(n115) );
    inv_0 U17 ( .x(n280), .a(n233) );
    oa21_2 U170 ( .x(n51), .a(n218), .b(n279), .c(n281) );
    inv_2 U171 ( .x(n248), .a(n84) );
    nand2i_3 U172 ( .x(n325), .a(B[9]), .b(A[9]) );
    inv_5 U173 ( .x(n118), .a(n325) );
    exnor2_3 U175 ( .x(DIFF[28]), .a(n53), .b(n52) );
    inv_2 U176 ( .x(n52), .a(n263) );
    ao21_3 U177 ( .x(n53), .a(n212), .b(n213), .c(n157) );
    nand2i_2 U179 ( .x(n284), .a(B[15]), .b(A[15]) );
    and4_3 U18 ( .x(n57), .a(n277), .b(n110), .c(n278), .d(n115) );
    exnor2_1 U180 ( .x(n267), .a(A[24]), .b(B[24]) );
    nand2i_2 U181 ( .x(n359), .a(B[24]), .b(n303) );
    nand2i_2 U182 ( .x(n240), .a(B[24]), .b(A[24]) );
    exnor2_1 U183 ( .x(n263), .a(A[28]), .b(B[28]) );
    nand2i_2 U184 ( .x(n346), .a(A[28]), .b(n344) );
    nand2i_0 U185 ( .x(n355), .a(A[28]), .b(B[28]) );
    inv_2 U186 ( .x(n54), .a(n250) );
    nor2i_3 U187 ( .x(n98), .a(n100), .b(n99) );
    inv_2 U188 ( .x(n202), .a(n88) );
    nor2_4 U189 ( .x(n254), .a(n166), .b(n88) );
    inv_5 U19 ( .x(n65), .a(n179) );
    nor2i_1 U190 ( .x(n142), .a(n143), .b(n88) );
    nor2i_3 U191 ( .x(n88), .a(n90), .b(n89) );
    nor2i_3 U192 ( .x(n290), .a(n291), .b(n233) );
    inv_0 U193 ( .x(n82), .a(n247) );
    inv_0 U194 ( .x(n55), .a(n313) );
    inv_2 U195 ( .x(n56), .a(n55) );
    nand3_2 U197 ( .x(n296), .a(n57), .b(n63), .c(n290) );
    or3i_2 U20 ( .x(n288), .a(n316), .b(n160), .c(A[3]) );
    nor2_3 U200 ( .x(n259), .a(n58), .b(n118) );
    nor3i_5 U202 ( .x(n63), .a(n81), .b(n64), .c(n241) );
    or3i_2 U203 ( .x(n289), .a(n63), .b(n233), .c(n155) );
    exor2_1 U204 ( .x(n275), .a(B[1]), .b(A[1]) );
    inv_0 U205 ( .x(n186), .a(A[1]) );
    nand2i_2 U207 ( .x(n278), .a(A[1]), .b(B[1]) );
    aoi21_1 U208 ( .x(n153), .a(A[3]), .b(n154), .c(n155) );
    nand2_8 U209 ( .x(n59), .a(A[16]), .b(n80) );
    exnor2_5 U210 ( .x(DIFF[31]), .a(n219), .b(n105) );
    exnor2_1 U211 ( .x(DIFF[24]), .a(n266), .b(n267) );
    aoai211_3 U212 ( .x(n101), .a(n359), .b(n358), .c(n266), .d(n301) );
    aoai211_4 U213 ( .x(n102), .a(n359), .b(n358), .c(n266), .d(n301) );
    aoi21_2 U214 ( .x(n201), .a(A[20]), .b(n202), .c(n142) );
    oai21_2 U215 ( .x(n295), .a(n286), .b(n289), .c(n296) );
    or3i_3 U216 ( .x(n336), .a(n258), .b(n179), .c(n246) );
    nand2_2 U217 ( .x(n261), .a(n242), .b(n243) );
    inv_3 U218 ( .x(n138), .a(n63) );
    inv_0 U219 ( .x(n60), .a(n241) );
    or3i_3 U22 ( .x(n287), .a(n316), .b(n160), .c(n154) );
    inv_2 U220 ( .x(n61), .a(n60) );
    nand2i_2 U221 ( .x(n321), .a(B[4]), .b(A[4]) );
    nand2i_2 U222 ( .x(n291), .a(A[4]), .b(B[4]) );
    nand4_4 U223 ( .x(n241), .a(n242), .b(n243), .c(n244), .d(n245) );
    inv_10 U224 ( .x(n242), .a(n66) );
    buf_2 U225 ( .x(n62), .a(n234) );
    nand2i_2 U226 ( .x(n181), .a(B[11]), .b(A[11]) );
    inv_0 U227 ( .x(n208), .a(n331) );
    aoi21_3 U229 ( .x(n292), .a(n293), .b(n294), .c(n135) );
    ao211_5 U231 ( .x(n357), .a(n197), .b(n97), .c(n95), .d(n96) );
    inv_3 U232 ( .x(n97), .a(n297) );
    nor2i_1 U233 ( .x(n92), .a(A[5]), .b(B[5]) );
    oai21_1 U234 ( .x(n256), .a(A[17]), .b(n165), .c(n194) );
    aoai211_1 U235 ( .x(n310), .a(A[17]), .b(n165), .c(n311), .d(n312) );
    aoi21_1 U236 ( .x(n164), .a(A[17]), .b(n165), .c(n166) );
    nand2_6 U237 ( .x(n64), .a(n294), .b(n65) );
    inv_7 U238 ( .x(n179), .a(n334) );
    nor2_8 U239 ( .x(n66), .a(A[10]), .b(n67) );
    nand2i_2 U24 ( .x(n115), .a(A[3]), .b(B[3]) );
    exnor2_3 U240 ( .x(DIFF[30]), .a(n262), .b(n68) );
    exnor2_1 U241 ( .x(n68), .a(A[30]), .b(n69) );
    inv_0 U242 ( .x(n69), .a(B[30]) );
    nand2i_2 U244 ( .x(n308), .a(A[30]), .b(n309) );
    buf_1 U245 ( .x(n70), .a(n212) );
    inv_2 U246 ( .x(n165), .a(B[17]) );
    exor2_1 U247 ( .x(n274), .a(A[17]), .b(B[17]) );
    nand2i_0 U248 ( .x(n312), .a(A[17]), .b(B[17]) );
    nand2i_2 U249 ( .x(n329), .a(B[17]), .b(A[17]) );
    nand2i_2 U25 ( .x(n277), .a(A[2]), .b(B[2]) );
    nand2i_2 U250 ( .x(n192), .a(A[17]), .b(B[17]) );
    nor2i_2 U251 ( .x(n193), .a(A[17]), .b(B[17]) );
    nand2i_2 U252 ( .x(n314), .a(A[17]), .b(B[17]) );
    exnor2_3 U253 ( .x(DIFF[29]), .a(n75), .b(n71) );
    inv_2 U254 ( .x(n71), .a(n222) );
    exnor2_1 U255 ( .x(n72), .a(n74), .b(n73) );
    inv_2 U256 ( .x(n222), .a(n72) );
    inv_0 U257 ( .x(n73), .a(B[29]) );
    inv_2 U258 ( .x(n74), .a(A[29]) );
    aoai211_1 U259 ( .x(n75), .a(n70), .b(n76), .c(n77), .d(n355) );
    nand2i_3 U26 ( .x(n315), .a(B[2]), .b(A[2]) );
    inv_2 U260 ( .x(n76), .a(n158) );
    and2_1 U261 ( .x(n77), .a(n346), .b(n345) );
    inv_2 U262 ( .x(n211), .a(n355) );
    inv_2 U263 ( .x(n158), .a(n213) );
    inv_2 U265 ( .x(n264), .a(n102) );
    nand2i_2 U266 ( .x(n309), .a(B[29]), .b(A[29]) );
    exnor2_1 U268 ( .x(n272), .a(A[20]), .b(B[20]) );
    nor2i_0 U269 ( .x(n134), .a(B[20]), .b(A[20]) );
    nor2_1 U27 ( .x(n125), .a(n126), .b(n127) );
    inv_0 U270 ( .x(n143), .a(B[20]) );
    nor2i_2 U271 ( .x(n78), .a(n252), .b(n79) );
    inv_0 U272 ( .x(n251), .a(n78) );
    inv_0 U273 ( .x(n200), .a(n79) );
    inv_2 U274 ( .x(n80), .a(B[16]) );
    nor2_8 U275 ( .x(n81), .a(n84), .b(n175) );
    nor2_8 U276 ( .x(n84), .a(A[14]), .b(n85) );
    inv_0 U277 ( .x(n170), .a(n294) );
    aoai211_1 U278 ( .x(n224), .a(B[24]), .b(n239), .c(n266), .d(n240) );
    nand2i_0 U279 ( .x(n86), .a(n295), .b(n292) );
    nand3i_3 U282 ( .x(n219), .a(n189), .b(n351), .c(n350) );
    inv_0 U283 ( .x(n87), .a(B[30]) );
    ao211_5 U284 ( .x(n93), .a(n197), .b(n97), .c(n96), .d(n95) );
    inv_2 U285 ( .x(n90), .a(A[19]) );
    aoai211_3 U286 ( .x(n258), .a(n259), .b(n260), .c(n261), .d(n181) );
    inv_0 U287 ( .x(n184), .a(n242) );
    inv_2 U288 ( .x(n91), .a(n129) );
    inv_0 U289 ( .x(n129), .a(n322) );
    oai21_1 U29 ( .x(n216), .a(n130), .b(n326), .c(n91) );
    inv_2 U290 ( .x(n322), .a(n92) );
    nand2i_4 U291 ( .x(n299), .a(A[22]), .b(B[22]) );
    inv_8 U292 ( .x(n255), .a(A[18]) );
    ao221_4 U293 ( .x(n94), .a(n102), .b(A[26]), .c(n102), .d(n109), .e(n108)
         );
    inv_2 U294 ( .x(n95), .a(n356) );
    nand2i_0 U295 ( .x(n356), .a(B[20]), .b(A[20]) );
    nand2i_2 U296 ( .x(n297), .a(n134), .b(n210) );
    nand2i_0 U297 ( .x(n111), .a(B[0]), .b(A[0]) );
    exnor2_1 U298 ( .x(n273), .a(A[18]), .b(B[18]) );
    nor2_0 U299 ( .x(n120), .a(n54), .b(n121) );
    nor2_0 U30 ( .x(n177), .a(n178), .b(n179) );
    nand2_2 U300 ( .x(n260), .a(n98), .b(n244) );
    inv_0 U301 ( .x(n250), .a(n98) );
    inv_10 U302 ( .x(n266), .a(n364) );
    nand4i_3 U303 ( .x(n268), .a(n148), .b(n338), .c(n339), .d(n340) );
    inv_0 U304 ( .x(n103), .a(n268) );
    inv_1 U305 ( .x(n104), .a(n103) );
    nand2i_4 U306 ( .x(n338), .a(n298), .b(n93) );
    exor2_1 U307 ( .x(DIFF[23]), .a(n104), .b(n269) );
    inv_2 U308 ( .x(n105), .a(n220) );
    exor2_1 U309 ( .x(n220), .a(A[31]), .b(B[31]) );
    exor2_1 U31 ( .x(DIFF[7]), .a(n215), .b(n122) );
    exor2_1 U310 ( .x(DIFF[16]), .a(n86), .b(n167) );
    aoi21_1 U311 ( .x(n199), .a(n86), .b(n200), .c(n311) );
    aoi21_1 U312 ( .x(n195), .a(n196), .b(n86), .c(n198) );
    aoi22_1 U313 ( .x(n203), .a(n204), .b(n205), .c(n206), .d(n86) );
    aoi21_1 U314 ( .x(n209), .a(n210), .b(n86), .c(n207) );
    inv_0 U315 ( .x(n335), .a(n258) );
    exnor2_1 U316 ( .x(DIFF[26]), .a(n264), .b(n265) );
    oai221_1 U317 ( .x(n223), .a(B[26]), .b(n264), .c(n264), .d(n238), .e(n343
        ) );
    ao221_4 U319 ( .x(n212), .a(n101), .b(A[26]), .c(n101), .d(n109), .e(n108)
         );
    oai21_1 U32 ( .x(n215), .a(n127), .b(n327), .c(n319) );
    inv_2 U320 ( .x(n108), .a(n343) );
    inv_0 U321 ( .x(n109), .a(B[26]) );
    nand2i_0 U322 ( .x(n343), .a(B[26]), .b(A[26]) );
    inv_0 U323 ( .x(n238), .a(A[26]) );
    aoi21_3 U324 ( .x(n135), .a(n136), .b(n137), .c(n138) );
    exor2_3 U325 ( .x(DIFF[15]), .a(n227), .b(n169) );
    nand2_5 U326 ( .x(n253), .a(n254), .b(n78) );
    nand3i_3 U327 ( .x(n286), .a(n133), .b(n287), .c(n288) );
    nor2i_3 U328 ( .x(n305), .a(n306), .b(n211) );
    nor2i_3 U329 ( .x(n307), .a(A[29]), .b(n211) );
    inv_0 U33 ( .x(n127), .a(n236) );
    ao21_4 U330 ( .x(n227), .a(n228), .b(n248), .c(n173) );
    oai21_4 U331 ( .x(n137), .a(n126), .b(n124), .c(n235) );
    nand3i_3 U332 ( .x(n317), .a(n155), .b(n288), .c(n287) );
    nand2i_4 U333 ( .x(n328), .a(B[19]), .b(A[19]) );
    nand2i_4 U334 ( .x(n341), .a(B[23]), .b(A[23]) );
    nand2i_4 U337 ( .x(n339), .a(n300), .b(n357) );
    inv_5 U338 ( .x(n361), .a(n256) );
    oai21_4 U339 ( .x(n332), .a(n311), .b(n360), .c(n361) );
    inv_2 U34 ( .x(n327), .a(n216) );
    nand2i_4 U340 ( .x(n362), .a(n201), .b(n331) );
    nand2i_4 U341 ( .x(n363), .a(n149), .b(n268) );
    nand2_5 U342 ( .x(n364), .a(n363), .b(n341) );
    nand2_4 U344 ( .x(n340), .a(n337), .b(n299) );
    nand2i_6 U345 ( .x(n213), .a(A[27]), .b(B[27]) );
    nand2i_6 U346 ( .x(n249), .a(B[12]), .b(A[12]) );
    nand2i_5 U347 ( .x(n358), .a(n239), .b(n303) );
    aoi21_4 U348 ( .x(n301), .a(n302), .b(n303), .c(n304) );
    nand2i_6 U349 ( .x(n344), .a(B[27]), .b(A[27]) );
    nor2_1 U35 ( .x(n122), .a(n123), .b(n124) );
    nor2i_5 U350 ( .x(n114), .a(n115), .b(n116) );
    nand3i_1 U351 ( .x(n262), .a(n347), .b(n348), .c(n349) );
    nand3i_2 U352 ( .x(n351), .a(n308), .b(n348), .c(n349) );
    aoai211_3 U353 ( .x(n349), .a(n212), .b(n213), .c(n188), .d(n307) );
    or3i_5 U354 ( .x(n293), .a(n336), .b(n139), .c(n285) );
    nand4i_1 U355 ( .x(n350), .a(n87), .b(n349), .c(n348), .d(n309) );
    aoai211_3 U356 ( .x(n348), .a(n213), .b(n94), .c(n150), .d(n305) );
    nand2i_5 U357 ( .x(n316), .a(n232), .b(n277) );
    inv_0 U358 ( .x(n187), .a(n232) );
    nand2i_3 U359 ( .x(n232), .a(B[1]), .b(A[1]) );
    inv_2 U36 ( .x(n123), .a(n235) );
    inv_3 U360 ( .x(n100), .a(B[8]) );
    nand2i_2 U361 ( .x(n245), .a(A[8]), .b(B[8]) );
    inv_3 U362 ( .x(n58), .a(n313) );
    nand2i_3 U363 ( .x(n313), .a(B[10]), .b(A[10]) );
    nand2i_4 U364 ( .x(n197), .a(n295), .b(n292) );
    nand3i_5 U365 ( .x(n233), .a(n365), .b(n235), .c(n236) );
    inv_2 U366 ( .x(n365), .a(n234) );
    nand2i_3 U367 ( .x(n236), .a(A[6]), .b(B[6]) );
    nand2i_2 U368 ( .x(n235), .a(A[7]), .b(B[7]) );
    nand2_0 U369 ( .x(n141), .a(n83), .b(A[13]) );
    nand2_0 U37 ( .x(DIFF[0]), .a(n110), .b(n111) );
    inv_5 U370 ( .x(n83), .a(B[13]) );
    nand2i_2 U371 ( .x(n234), .a(A[5]), .b(B[5]) );
    inv_3 U372 ( .x(n85), .a(B[14]) );
    nand2i_4 U373 ( .x(n294), .a(A[15]), .b(B[15]) );
    nand2i_2 U374 ( .x(n319), .a(B[6]), .b(A[6]) );
    nor2i_0 U375 ( .x(n149), .a(B[23]), .b(A[23]) );
    inv_3 U376 ( .x(n67), .a(B[10]) );
    inv_5 U377 ( .x(n194), .a(B[18]) );
    nand2i_2 U378 ( .x(n252), .a(A[18]), .b(B[18]) );
    inv_0 U38 ( .x(n276), .a(n110) );
    nand2i_2 U39 ( .x(n243), .a(A[11]), .b(B[11]) );
    nor2i_1 U40 ( .x(n180), .a(n181), .b(n182) );
    oai21_1 U41 ( .x(n230), .a(n184), .b(n354), .c(n56) );
    inv_0 U42 ( .x(n89), .a(B[19]) );
    nor2i_1 U43 ( .x(n207), .a(n202), .b(n208) );
    nor2_0 U44 ( .x(n172), .a(n140), .b(n173) );
    inv_2 U45 ( .x(n140), .a(n248) );
    inv_2 U47 ( .x(n176), .a(n141) );
    or2_6 U48 ( .x(n247), .a(A[13]), .b(n83) );
    nor2_1 U49 ( .x(n174), .a(n82), .b(n176) );
    inv_2 U50 ( .x(n178), .a(n249) );
    oai21_1 U51 ( .x(n229), .a(n51), .b(n61), .c(n335) );
    inv_2 U52 ( .x(n353), .a(n229) );
    nand2i_2 U53 ( .x(n334), .a(A[12]), .b(B[12]) );
    oa21_2 U54 ( .x(n50), .a(n179), .b(n353), .c(n249) );
    nor2_1 U55 ( .x(n183), .a(n55), .b(n184) );
    inv_2 U56 ( .x(n354), .a(n231) );
    oai21_1 U57 ( .x(n231), .a(n324), .b(n119), .c(n325) );
    inv_0 U58 ( .x(n113), .a(n93) );
    nor2i_0 U59 ( .x(n112), .a(A[21]), .b(n113) );
    inv_0 U6 ( .x(n182), .a(n243) );
    inv_4 U60 ( .x(n96), .a(n362) );
    inv_2 U61 ( .x(n145), .a(B[21]) );
    nor2i_1 U62 ( .x(n144), .a(n145), .b(n113) );
    inv_2 U63 ( .x(n130), .a(n62) );
    nor2_1 U64 ( .x(n128), .a(n129), .b(n130) );
    oai21_1 U65 ( .x(n217), .a(n218), .b(n133), .c(n321) );
    nand2i_2 U66 ( .x(n318), .a(n114), .b(n317) );
    inv_2 U67 ( .x(n326), .a(n217) );
    inv_2 U68 ( .x(n166), .a(n314) );
    nor2_1 U69 ( .x(n206), .a(n251), .b(n166) );
    nand3_1 U7 ( .x(n116), .a(n277), .b(n110), .c(n278) );
    nand2i_0 U70 ( .x(n205), .a(n194), .b(n310) );
    nand2i_3 U72 ( .x(n330), .a(B[16]), .b(A[16]) );
    aoai211_1 U73 ( .x(n204), .a(n329), .b(n330), .c(n256), .d(n255) );
    nor2_1 U74 ( .x(n131), .a(n132), .b(n133) );
    inv_2 U75 ( .x(n132), .a(n321) );
    inv_2 U76 ( .x(n133), .a(n291) );
    nor2_1 U77 ( .x(n196), .a(n168), .b(n166) );
    nor2_1 U78 ( .x(n188), .a(n151), .b(n152) );
    inv_0 U79 ( .x(n306), .a(B[29]) );
    nand2_2 U8 ( .x(n323), .a(n322), .b(n321) );
    nor2_1 U80 ( .x(n150), .a(n151), .b(n152) );
    nand4_1 U81 ( .x(n136), .a(n62), .b(n235), .c(n323), .d(n236) );
    inv_2 U82 ( .x(n282), .a(n136) );
    inv_2 U83 ( .x(n124), .a(n320) );
    inv_2 U84 ( .x(n126), .a(n319) );
    nor2i_1 U85 ( .x(n281), .a(n137), .b(n282) );
    nand2i_2 U87 ( .x(n279), .a(n133), .b(n280) );
    inv_2 U88 ( .x(n151), .a(n345) );
    inv_2 U89 ( .x(n152), .a(n346) );
    nand2i_0 U9 ( .x(n320), .a(B[7]), .b(A[7]) );
    nand2i_2 U90 ( .x(n345), .a(n237), .b(n344) );
    nor2i_0 U91 ( .x(n189), .a(B[30]), .b(A[30]) );
    nand2i_2 U92 ( .x(n110), .a(A[0]), .b(B[0]) );
    aoi21_1 U93 ( .x(n185), .a(B[1]), .b(n186), .c(n187) );
    nand2i_2 U95 ( .x(n244), .a(A[9]), .b(B[9]) );
    inv_2 U96 ( .x(n119), .a(n244) );
    nor2_1 U97 ( .x(n117), .a(n118), .b(n119) );
    inv_2 U98 ( .x(n324), .a(n214) );
    inv_0 U99 ( .x(n99), .a(A[8]) );
endmodule


module EX_DW01_add_32_2_test_1 ( A, B, CI, SUM, CO );
input  [31:0] A;
input  [31:0] B;
output [31:0] SUM;
input  CI;
output CO;
    wire ___cell__39170_net140238, ___cell__39170_net140310, n224, n203, n216, 
        n205, n223, n180, ___cell__39170_net140214, ___cell__39170_net140460, 
        n202, n104, ___cell__39170_net140251, ___cell__39170_net140286, n98, 
        ___cell__39170_net140285, ___cell__39170_net140357, 
        ___cell__39170_net140264, ___cell__39170_net140355, n175, 
        ___cell__39170_net140279, ___cell__39170_net140209, 
        ___cell__39170_net140484, n233, n134, ___cell__39170_net140210, n121, 
        n184, n49, ___cell__39170_net140316, n245, n247, 
        ___cell__39170_net140273, n144, n120, ___cell__39170_net140502, 
        ___cell__39170_net140193, n145, n146, n168, n150, n166, n167, n70, 
        ___cell__39170_net140246, ___cell__39170_net140199, n135, n194, n141, 
        n142, ___cell__39170_net140307, ___cell__39170_net140504, n232, n177, 
        n56, ___cell__39170_net140284, n58, n240, n241, net150837, n183, 
        ___cell__39170_net140309, ___cell__39170_net140305, n191, n163, n149, 
        n164, n151, n165, n91, n193, n169, ___cell__39170_net140269, 
        ___cell__39170_net140185, ___cell__39170_net140184, 
        ___cell__39170_net140274, ___cell__39170_net140192, n62, 
        ___cell__39170_net140311, ___cell__39170_net140197, n234, n148, n157, 
        n185, n178, n147, ___cell__39170_net140490, ___cell__39170_net140499, 
        ___cell__39170_net140321, ___cell__39170_net140445, 
        ___cell__39170_net140444, ___cell__39170_net140282, n179, n50, 
        net151953, n57, net151951, n93, n95, n94, n231, net156380, 
        ___cell__39170_net140267, n246, n140, ___cell__39170_net140495, n125, 
        ___cell__39170_net140319, n112, ___cell__39170_net140341, 
        ___cell__39170_net140395, ___cell__39170_net140476, 
        ___cell__39170_net140396, n236, n189, net152474, 
        ___cell__39170_net140223, n190, n188, n160, ___cell__39170_net140257, 
        n138, n139, n154, ___cell__39170_net140288, ___cell__39170_net140287, 
        n156, n243, n143, n196, n97, n51, n106, n99, n100, n87, n132, n52, n66, 
        n61, n89, ___cell__39170_net140386, n53, n54, n55, n124, n220, n72, 
        n217, n250, n77, n218, ___cell__39170_net140546, 
        ___cell__39170_net140320, ___cell__39170_net140317, n82, n214, 
        ___cell__39170_net140242, ___cell__39170_net140244, n79, n88, n200, 
        n226, n71, n126, n127, n59, n238, n208, n162, ___cell__39170_net140266, 
        n109, ___cell__39170_net140337, ___cell__39170_net140327, n210, n63, 
        n198, n199, ___cell__39170_net140448, n129, n128, n74, n64, 
        ___cell__39170_net140471, ___cell__39170_net140258, 
        ___cell__39170_net140241, n65, n133, n130, n195, n227, n209, 
        ___cell__39170_net140427, ___cell__39170_net140292, net150142, 
        ___cell__39170_net140561, ___cell__39170_net140560, 
        ___cell__39170_net140455, n171, n131, n69, n68, n67, 
        ___cell__39170_net140514, ___cell__39170_net140513, 
        ___cell__39170_net140259, n172, n173, ___cell__39170_net140249, n122, 
        n155, n212, n211, n215, n114, n73, n153, ___cell__39170_net140451, 
        ___cell__39170_net140256, ___cell__39170_net140218, n197, n80, n81, 
        n83, n96, ___cell__39170_net140401, n237, ___cell__39170_net140566, 
        n152, ___cell__39170_net140452, ___cell__39170_net140525, 
        ___cell__39170_net140268, n85, n86, ___cell__39170_net140397, n113, 
        ___cell__39170_net140392, ___cell__39170_net140412, 
        ___cell__39170_net140398, n60, ___cell__39170_net140236, n207, n90, 
        n108, ___cell__39170_net140276, net150005, ___cell__39170_net140213, 
        net150690, net156215, net151417, n228, ___cell__39170_net140482, 
        ___cell__39170_net140270, ___cell__39170_net140278, 
        ___cell__39170_net140250, ___cell__39170_net140528, 
        ___cell__39170_net140529, n229, ___cell__39170_net140461, 
        ___cell__39170_net140416, ___cell__39170_net140313, net155900, 
        ___cell__39170_net140283, n105, ___cell__39170_net140536, 
        ___cell__39170_net140464, n101, ___cell__39170_net140351, n102, 
        ___cell__39170_net140410, ___cell__39170_net140411, n103, 
        ___cell__39170_net140447, ___cell__39170_net140239, n111, net151032, 
        net151031, net151030, ___cell__39170_net140541, 
        ___cell__39170_net140424, ___cell__39170_net140422, n110, 
        ___cell__39170_net140233, ___cell__39170_net140235, n115, 
        ___cell__39170_net140537, n119, ___cell__39170_net140418, 
        ___cell__39170_net140255, net150555, ___cell__39170_net140277, n174, 
        net152445, n170, n244, n219, n225, n187, n176, n201, n206, n204, 
        net121836, n161, n213, n84, n221, n222, n92, n230, n136, n137, 
        net155899, n76, n181, n248, n182, n239, n249, ___cell__39170_net140231, 
        n192, ___cell__39170_net140485, ___cell__39170_net140232, n78, n75, 
        n251, n252, n107, n158, n159, n123, ___cell__39170_net140463, n116, 
        n117, n118, n242, n235, n186;
    inv_4 U10 ( .x(___cell__39170_net140238), .a(___cell__39170_net140310) );
    nor2i_1 U100 ( .x(n224), .a(n203), .b(n216) );
    inv_0 U101 ( .x(n203), .a(A[21]) );
    inv_0 U102 ( .x(n205), .a(B[20]) );
    exnor2_1 U103 ( .x(n223), .a(n216), .b(n203) );
    exor2_1 U104 ( .x(n180), .a(A[23]), .b(B[23]) );
    inv_2 U105 ( .x(___cell__39170_net140214), .a(___cell__39170_net140460) );
    inv_2 U106 ( .x(n202), .a(A[24]) );
    inv_2 U107 ( .x(n104), .a(A[23]) );
    nand2_2 U108 ( .x(___cell__39170_net140251), .a(B[23]), .b(A[23]) );
    exor2_1 U109 ( .x(___cell__39170_net140286), .a(B[25]), .b(A[25]) );
    inv_5 U11 ( .x(n98), .a(A[2]) );
    exor2_1 U110 ( .x(___cell__39170_net140285), .a(A[26]), .b(B[26]) );
    nand2_2 U111 ( .x(___cell__39170_net140357), .a(B[25]), .b(A[25]) );
    inv_2 U112 ( .x(___cell__39170_net140264), .a(___cell__39170_net140357) );
    inv_2 U113 ( .x(___cell__39170_net140355), .a(A[25]) );
    nand2i_2 U114 ( .x(n175), .a(B[25]), .b(___cell__39170_net140355) );
    exor2_1 U115 ( .x(SUM[3]), .a(___cell__39170_net140279), .b(
        ___cell__39170_net140209) );
    nand3_1 U116 ( .x(___cell__39170_net140279), .a(___cell__39170_net140484), 
        .b(n233), .c(n134) );
    nor2i_1 U117 ( .x(___cell__39170_net140209), .a(___cell__39170_net140210), 
        .b(n121) );
    exnor2_1 U118 ( .x(SUM[2]), .a(n184), .b(n49) );
    nand2i_0 U119 ( .x(n184), .a(___cell__39170_net140238), .b(
        ___cell__39170_net140316) );
    nand2i_4 U12 ( .x(___cell__39170_net140310), .a(B[2]), .b(n98) );
    inv_2 U120 ( .x(n245), .a(n247) );
    exor2_1 U121 ( .x(SUM[6]), .a(___cell__39170_net140273), .b(n144) );
    oai21_1 U122 ( .x(___cell__39170_net140273), .a(n120), .b(
        ___cell__39170_net140502), .c(___cell__39170_net140193) );
    nor2i_0 U123 ( .x(n144), .a(n145), .b(n146) );
    inv_2 U124 ( .x(n168), .a(n150) );
    nor2i_0 U125 ( .x(n166), .a(n167), .b(n168) );
    inv_2 U126 ( .x(n70), .a(___cell__39170_net140246) );
    exor2_1 U127 ( .x(SUM[12]), .a(___cell__39170_net140199), .b(n166) );
    inv_0 U128 ( .x(n135), .a(n194) );
    nor2i_1 U129 ( .x(n141), .a(n142), .b(n135) );
    inv_2 U13 ( .x(___cell__39170_net140307), .a(B[0]) );
    inv_2 U130 ( .x(___cell__39170_net140504), .a(___cell__39170_net140273) );
    inv_0 U131 ( .x(n146), .a(n232) );
    oai21_1 U132 ( .x(n177), .a(n146), .b(___cell__39170_net140504), .c(n145)
         );
    exor2_1 U133 ( .x(SUM[7]), .a(n177), .b(n141) );
    inv_0 U134 ( .x(n56), .a(A[27]) );
    exor2_1 U135 ( .x(___cell__39170_net140284), .a(B[27]), .b(n58) );
    nor2i_1 U136 ( .x(SUM[0]), .a(n240), .b(n241) );
    exor2_1 U139 ( .x(SUM[20]), .a(net150837), .b(n183) );
    or3i_2 U14 ( .x(___cell__39170_net140309), .a(___cell__39170_net140310), 
        .b(___cell__39170_net140305), .c(___cell__39170_net140307) );
    exor2_1 U140 ( .x(SUM[14]), .a(n191), .b(n163) );
    exnor2_1 U141 ( .x(SUM[13]), .a(n149), .b(n164) );
    aoi21_1 U142 ( .x(n149), .a(___cell__39170_net140199), .b(n150), .c(n151)
         );
    inv_2 U143 ( .x(n151), .a(n167) );
    nor2i_0 U144 ( .x(n164), .a(n165), .b(n91) );
    exor2_1 U146 ( .x(SUM[10]), .a(n193), .b(n169) );
    oai21_1 U147 ( .x(n193), .a(___cell__39170_net140269), .b(
        ___cell__39170_net140185), .c(___cell__39170_net140184) );
    exor2_1 U149 ( .x(SUM[5]), .a(___cell__39170_net140274), .b(
        ___cell__39170_net140192) );
    nand2i_1 U15 ( .x(n62), .a(___cell__39170_net140311), .b(
        ___cell__39170_net140310) );
    oai21_1 U150 ( .x(___cell__39170_net140274), .a(___cell__39170_net140197), 
        .b(n234), .c(n148) );
    nor2i_1 U151 ( .x(___cell__39170_net140192), .a(___cell__39170_net140193), 
        .b(n120) );
    inv_2 U152 ( .x(___cell__39170_net140502), .a(___cell__39170_net140274) );
    exnor2_1 U153 ( .x(SUM[19]), .a(n157), .b(n185) );
    exor2_1 U154 ( .x(SUM[4]), .a(n178), .b(n147) );
    nand2i_2 U155 ( .x(n178), .a(___cell__39170_net140490), .b(
        ___cell__39170_net140499) );
    inv_2 U156 ( .x(___cell__39170_net140490), .a(___cell__39170_net140210) );
    nor2i_1 U157 ( .x(n147), .a(n148), .b(___cell__39170_net140197) );
    inv_2 U158 ( .x(___cell__39170_net140197), .a(___cell__39170_net140321) );
    inv_2 U159 ( .x(n234), .a(n178) );
    nor2i_1 U16 ( .x(___cell__39170_net140445), .a(___cell__39170_net140444), 
        .b(n62) );
    exor2_1 U161 ( .x(___cell__39170_net140282), .a(B[28]), .b(A[28]) );
    ao221_1 U162 ( .x(n179), .a(n50), .b(net151953), .c(n50), .d(n57), .e(
        net151951) );
    exor2_1 U163 ( .x(SUM[28]), .a(n179), .b(___cell__39170_net140282) );
    nor2i_1 U164 ( .x(n93), .a(n95), .b(n94) );
    inv_2 U165 ( .x(n94), .a(n231) );
    inv_5 U166 ( .x(net156380), .a(___cell__39170_net140267) );
    exnor2_1 U167 ( .x(SUM[1]), .a(n246), .b(n240) );
    exnor2_1 U168 ( .x(SUM[9]), .a(___cell__39170_net140269), .b(n140) );
    inv_2 U169 ( .x(___cell__39170_net140269), .a(___cell__39170_net140495) );
    inv_4 U17 ( .x(n125), .a(___cell__39170_net140319) );
    oai22_1 U170 ( .x(___cell__39170_net140495), .a(n112), .b(
        ___cell__39170_net140341), .c(___cell__39170_net140395), .d(n93) );
    inv_2 U171 ( .x(n112), .a(B[8]) );
    inv_5 U172 ( .x(___cell__39170_net140341), .a(A[8]) );
    inv_5 U173 ( .x(___cell__39170_net140395), .a(___cell__39170_net140476) );
    nor2i_1 U174 ( .x(n140), .a(___cell__39170_net140184), .b(
        ___cell__39170_net140185) );
    inv_2 U175 ( .x(___cell__39170_net140185), .a(___cell__39170_net140396) );
    inv_2 U176 ( .x(n236), .a(n191) );
    oai21_1 U177 ( .x(n189), .a(net152474), .b(n236), .c(
        ___cell__39170_net140223) );
    exor2_1 U178 ( .x(SUM[15]), .a(n189), .b(n190) );
    exnor2_1 U179 ( .x(SUM[16]), .a(n188), .b(n160) );
    nor2i_3 U18 ( .x(___cell__39170_net140257), .a(___cell__39170_net140444), 
        .b(___cell__39170_net140309) );
    nand2_2 U180 ( .x(SUM[21]), .a(n138), .b(n139) );
    nand2i_2 U181 ( .x(n139), .a(n154), .b(n216) );
    exnor2_1 U182 ( .x(SUM[23]), .a(___cell__39170_net140288), .b(n180) );
    exor2_1 U183 ( .x(SUM[24]), .a(___cell__39170_net140287), .b(n156) );
    or2_2 U184 ( .x(n49), .a(n243), .b(n245) );
    inv_2 U185 ( .x(n143), .a(n194) );
    nand2i_4 U186 ( .x(n194), .a(B[7]), .b(n196) );
    ao21_2 U187 ( .x(n50), .a(n97), .b(n51), .c(n106) );
    or2_2 U188 ( .x(n51), .a(n99), .b(n100) );
    nor2i_4 U189 ( .x(net152474), .a(n87), .b(A[14]) );
    nand2_0 U19 ( .x(n132), .a(A[19]), .b(B[19]) );
    nand2_2 U190 ( .x(n52), .a(n87), .b(n66) );
    nor2i_2 U191 ( .x(n61), .a(n89), .b(A[18]) );
    inv_3 U192 ( .x(___cell__39170_net140386), .a(B[15]) );
    inv_2 U193 ( .x(n53), .a(n54) );
    inv_2 U194 ( .x(n55), .a(n54) );
    inv_0 U195 ( .x(n57), .a(n56) );
    inv_0 U196 ( .x(n58), .a(n56) );
    inv_3 U197 ( .x(n124), .a(A[5]) );
    oai211_2 U198 ( .x(n220), .a(n188), .b(n72), .c(n217), .d(n250) );
    inv_2 U199 ( .x(n77), .a(n218) );
    nand2_2 U20 ( .x(___cell__39170_net140546), .a(A[29]), .b(B[29]) );
    inv_10 U200 ( .x(___cell__39170_net140320), .a(___cell__39170_net140317)
         );
    and3i_4 U201 ( .x(n82), .a(n214), .b(___cell__39170_net140242), .c(n52) );
    and3i_3 U202 ( .x(___cell__39170_net140244), .a(n79), .b(n88), .c(
        ___cell__39170_net140242) );
    nand2i_3 U203 ( .x(___cell__39170_net140242), .a(A[15]), .b(
        ___cell__39170_net140386) );
    or3i_3 U204 ( .x(n200), .a(___cell__39170_net140320), .b(
        ___cell__39170_net140210), .c(n226) );
    nand2_2 U205 ( .x(n71), .a(n126), .b(n127) );
    inv_0 U206 ( .x(n59), .a(n238) );
    nand2i_2 U207 ( .x(n238), .a(B[16]), .b(n208) );
    inv_2 U208 ( .x(n162), .a(n238) );
    nand2_8 U209 ( .x(___cell__39170_net140317), .a(n232), .b(n194) );
    nand2i_2 U21 ( .x(___cell__39170_net140266), .a(A[29]), .b(n109) );
    or3i_3 U211 ( .x(___cell__39170_net140337), .a(___cell__39170_net140320), 
        .b(n124), .c(___cell__39170_net140327) );
    inv_0 U212 ( .x(n210), .a(A[18]) );
    ao21_3 U214 ( .x(n63), .a(n145), .b(n142), .c(n143) );
    nand2_1 U215 ( .x(n142), .a(A[7]), .b(B[7]) );
    nand4_1 U216 ( .x(n198), .a(n199), .b(___cell__39170_net140337), .c(n200), 
        .d(n63) );
    aoai211_1 U217 ( .x(___cell__39170_net140448), .a(n129), .b(n128), .c(n74), 
        .d(n132) );
    inv_2 U218 ( .x(n64), .a(___cell__39170_net140471) );
    nand2_5 U219 ( .x(___cell__39170_net140258), .a(n88), .b(n82) );
    inv_4 U22 ( .x(n196), .a(A[7]) );
    inv_2 U220 ( .x(n66), .a(A[14]) );
    nor2i_0 U222 ( .x(___cell__39170_net140241), .a(___cell__39170_net140242), 
        .b(n79) );
    aoi21_2 U223 ( .x(n79), .a(n65), .b(n133), .c(n130) );
    nand2_0 U224 ( .x(n148), .a(B[4]), .b(A[4]) );
    nand2i_2 U225 ( .x(___cell__39170_net140321), .a(A[4]), .b(n195) );
    nand2_0 U226 ( .x(n227), .a(B[4]), .b(A[4]) );
    inv_0 U227 ( .x(n209), .a(A[17]) );
    inv_6 U228 ( .x(___cell__39170_net140427), .a(___cell__39170_net140292) );
    inv_0 U229 ( .x(___cell__39170_net140327), .a(B[5]) );
    inv_2 U23 ( .x(n87), .a(B[14]) );
    aoai211_3 U230 ( .x(net150142), .a(___cell__39170_net140561), .b(
        ___cell__39170_net140560), .c(___cell__39170_net140427), .d(
        ___cell__39170_net140455) );
    or3i_2 U231 ( .x(n199), .a(___cell__39170_net140320), .b(n171), .c(n227)
         );
    exor2_1 U232 ( .x(n190), .a(A[15]), .b(B[15]) );
    nand2_0 U233 ( .x(n131), .a(A[15]), .b(B[15]) );
    ao211_5 U234 ( .x(___cell__39170_net140199), .a(n70), .b(n69), .c(n68), 
        .d(n67) );
    inv_0 U235 ( .x(n67), .a(___cell__39170_net140514) );
    inv_0 U236 ( .x(n68), .a(___cell__39170_net140513) );
    inv_0 U237 ( .x(n69), .a(___cell__39170_net140259) );
    nor3_4 U238 ( .x(___cell__39170_net140246), .a(n172), .b(n173), .c(
        ___cell__39170_net140249) );
    inv_4 U239 ( .x(n122), .a(n71) );
    inv_0 U24 ( .x(n155), .a(A[22]) );
    inv_0 U240 ( .x(n121), .a(n127) );
    inv_0 U241 ( .x(n120), .a(n126) );
    nand2i_2 U242 ( .x(n126), .a(B[5]), .b(n124) );
    nand2i_0 U243 ( .x(n72), .a(n162), .b(n212) );
    nand2i_4 U244 ( .x(n211), .a(n162), .b(n212) );
    nand2i_2 U245 ( .x(n212), .a(B[17]), .b(n209) );
    inv_6 U246 ( .x(n215), .a(A[11]) );
    nor2i_1 U248 ( .x(n114), .a(A[8]), .b(n112) );
    inv_0 U249 ( .x(n73), .a(___cell__39170_net140311) );
    inv_2 U25 ( .x(n153), .a(B[22]) );
    nor3_2 U250 ( .x(___cell__39170_net140451), .a(___cell__39170_net140448), 
        .b(___cell__39170_net140244), .c(___cell__39170_net140256) );
    inv_0 U251 ( .x(___cell__39170_net140218), .a(n74) );
    inv_4 U252 ( .x(n197), .a(B[6]) );
    inv_2 U253 ( .x(n133), .a(net152474) );
    inv_2 U254 ( .x(n80), .a(___cell__39170_net140445) );
    inv_2 U255 ( .x(n81), .a(n172) );
    exnor2_5 U256 ( .x(SUM[30]), .a(n83), .b(n96) );
    inv_0 U257 ( .x(___cell__39170_net140401), .a(n82) );
    nand2i_2 U258 ( .x(n237), .a(___cell__39170_net140401), .b(
        ___cell__39170_net140199) );
    nand2_5 U259 ( .x(___cell__39170_net140566), .a(n51), .b(n97) );
    aoi21_1 U26 ( .x(n152), .a(n153), .b(n154), .c(n155) );
    nand3_2 U260 ( .x(___cell__39170_net140292), .a(___cell__39170_net140451), 
        .b(___cell__39170_net140452), .c(___cell__39170_net140525) );
    ao21_4 U261 ( .x(n83), .a(___cell__39170_net140267), .b(
        ___cell__39170_net140266), .c(___cell__39170_net140268) );
    inv_2 U263 ( .x(n85), .a(B[13]) );
    inv_10 U264 ( .x(n86), .a(A[6]) );
    nand2i_2 U265 ( .x(___cell__39170_net140397), .a(B[10]), .b(n113) );
    nor2_6 U266 ( .x(n88), .a(___cell__39170_net140392), .b(n211) );
    nand4_1 U268 ( .x(___cell__39170_net140412), .a(___cell__39170_net140398), 
        .b(___cell__39170_net140396), .c(n114), .d(n60) );
    inv_0 U269 ( .x(___cell__39170_net140236), .a(n60) );
    nand2_5 U27 ( .x(n207), .a(A[20]), .b(B[20]) );
    inv_2 U272 ( .x(n90), .a(n89) );
    aoai211_3 U274 ( .x(n108), .a(___cell__39170_net140561), .b(
        ___cell__39170_net140560), .c(___cell__39170_net140427), .d(
        ___cell__39170_net140455) );
    exnor2_3 U275 ( .x(SUM[31]), .a(___cell__39170_net140276), .b(net150005)
         );
    ao21_3 U276 ( .x(___cell__39170_net140525), .a(___cell__39170_net140514), 
        .b(___cell__39170_net140513), .c(___cell__39170_net140258) );
    nor2i_1 U277 ( .x(n156), .a(___cell__39170_net140213), .b(
        ___cell__39170_net140214) );
    inv_2 U278 ( .x(net150690), .a(net156215) );
    buf_2 U279 ( .x(net151417), .a(n97) );
    inv_2 U28 ( .x(n228), .a(n207) );
    inv_2 U280 ( .x(n208), .a(A[16]) );
    inv_2 U281 ( .x(___cell__39170_net140482), .a(___cell__39170_net140309) );
    inv_0 U282 ( .x(___cell__39170_net140270), .a(n93) );
    inv_0 U283 ( .x(n95), .a(n198) );
    nand2_0 U284 ( .x(___cell__39170_net140193), .a(B[5]), .b(A[5]) );
    nor2_0 U285 ( .x(n171), .a(B[5]), .b(A[5]) );
    oai22_1 U286 ( .x(n226), .a(A[4]), .b(B[4]), .c(B[5]), .d(A[5]) );
    inv_2 U287 ( .x(n96), .a(___cell__39170_net140278) );
    nand4i_3 U288 ( .x(n97), .a(___cell__39170_net140250), .b(
        ___cell__39170_net140528), .c(___cell__39170_net140529), .d(
        ___cell__39170_net140213) );
    nand2_1 U289 ( .x(n217), .a(B[17]), .b(A[17]) );
    nand2_2 U29 ( .x(___cell__39170_net140561), .a(n229), .b(B[20]) );
    nand2i_4 U290 ( .x(___cell__39170_net140528), .a(___cell__39170_net140461), 
        .b(n108) );
    exor3_1 U291 ( .x(SUM[29]), .a(A[29]), .b(B[29]), .c(
        ___cell__39170_net140267) );
    aoai211_1 U292 ( .x(___cell__39170_net140287), .a(n104), .b(
        ___cell__39170_net140416), .c(___cell__39170_net140288), .d(
        ___cell__39170_net140251) );
    inv_2 U293 ( .x(___cell__39170_net140416), .a(B[23]) );
    inv_0 U294 ( .x(___cell__39170_net140288), .a(n108) );
    inv_3 U295 ( .x(___cell__39170_net140305), .a(A[0]) );
    nand2i_2 U296 ( .x(___cell__39170_net140313), .a(___cell__39170_net140311), 
        .b(___cell__39170_net140310) );
    nand2_2 U297 ( .x(___cell__39170_net140316), .a(B[2]), .b(A[2]) );
    inv_0 U298 ( .x(net155900), .a(B[1]) );
    nand2i_6 U299 ( .x(___cell__39170_net140283), .a(n106), .b(
        ___cell__39170_net140566) );
    nand2i_2 U30 ( .x(n105), .a(n104), .b(___cell__39170_net140460) );
    nand2i_4 U300 ( .x(___cell__39170_net140536), .a(___cell__39170_net140464), 
        .b(___cell__39170_net140283) );
    oai22_3 U301 ( .x(n106), .a(n101), .b(___cell__39170_net140357), .c(
        ___cell__39170_net140351), .d(n102) );
    nand2i_4 U302 ( .x(___cell__39170_net140529), .a(n105), .b(net150142) );
    inv_0 U303 ( .x(net156215), .a(___cell__39170_net140427) );
    nand3i_3 U304 ( .x(___cell__39170_net140410), .a(___cell__39170_net140411), 
        .b(___cell__39170_net140412), .c(n103) );
    aoi31_1 U305 ( .x(n103), .a(n60), .b(___cell__39170_net140398), .c(
        ___cell__39170_net140447), .d(___cell__39170_net140239) );
    ao221_4 U306 ( .x(___cell__39170_net140276), .a(n111), .b(net151032), .c(
        n111), .d(net151031), .e(net151030) );
    inv_2 U307 ( .x(net151030), .a(___cell__39170_net140541) );
    nand2_0 U308 ( .x(___cell__39170_net140541), .a(A[30]), .b(B[30]) );
    inv_2 U309 ( .x(net151031), .a(___cell__39170_net140424) );
    nand2i_2 U31 ( .x(___cell__39170_net140461), .a(___cell__39170_net140416), 
        .b(___cell__39170_net140460) );
    inv_2 U310 ( .x(___cell__39170_net140424), .a(A[30]) );
    inv_2 U311 ( .x(net151032), .a(___cell__39170_net140422) );
    inv_0 U312 ( .x(___cell__39170_net140422), .a(B[30]) );
    aoai211_4 U313 ( .x(n111), .a(n110), .b(n109), .c(net156380), .d(
        ___cell__39170_net140546) );
    inv_6 U314 ( .x(n109), .a(B[29]) );
    exor2_1 U315 ( .x(___cell__39170_net140278), .a(B[30]), .b(A[30]) );
    nor2_2 U316 ( .x(___cell__39170_net140239), .a(___cell__39170_net140233), 
        .b(___cell__39170_net140235) );
    nand4i_5 U317 ( .x(___cell__39170_net140267), .a(n115), .b(
        ___cell__39170_net140536), .c(___cell__39170_net140537), .d(n119) );
    inv_0 U318 ( .x(___cell__39170_net140418), .a(B[27]) );
    nand2_0 U319 ( .x(___cell__39170_net140255), .a(n57), .b(B[27]) );
    nor2_1 U32 ( .x(___cell__39170_net140250), .a(___cell__39170_net140214), 
        .b(___cell__39170_net140251) );
    inv_0 U320 ( .x(net150555), .a(n125) );
    nand3_4 U321 ( .x(___cell__39170_net140319), .a(___cell__39170_net140320), 
        .b(___cell__39170_net140321), .c(n122) );
    inv_2 U322 ( .x(net151951), .a(___cell__39170_net140255) );
    nand2_2 U323 ( .x(n130), .a(n131), .b(___cell__39170_net140223) );
    inv_10 U324 ( .x(n128), .a(B[19]) );
    inv_2 U325 ( .x(net150005), .a(___cell__39170_net140277) );
    exor2_1 U326 ( .x(___cell__39170_net140277), .a(B[31]), .b(A[31]) );
    aoi21_1 U327 ( .x(n174), .a(n175), .b(net151417), .c(
        ___cell__39170_net140264) );
    exor2_1 U328 ( .x(SUM[25]), .a(net151417), .b(___cell__39170_net140286) );
    nor2_0 U329 ( .x(n134), .a(net152445), .b(n170) );
    and4i_3 U33 ( .x(n170), .a(___cell__39170_net140238), .b(A[0]), .c(B[0]), 
        .d(A[1]) );
    nand2_0 U330 ( .x(n240), .a(A[0]), .b(B[0]) );
    and3i_1 U331 ( .x(n243), .a(n244), .b(B[0]), .c(A[0]) );
    nor2_0 U332 ( .x(n241), .a(B[0]), .b(A[0]) );
    or2_6 U333 ( .x(n172), .a(n170), .b(net152445) );
    nand2_0 U334 ( .x(n219), .a(B[18]), .b(A[18]) );
    nor2i_2 U335 ( .x(n225), .a(A[18]), .b(n220) );
    inv_2 U336 ( .x(net151953), .a(___cell__39170_net140418) );
    exor2_1 U337 ( .x(SUM[27]), .a(n50), .b(___cell__39170_net140284) );
    nand2i_2 U338 ( .x(___cell__39170_net140460), .a(B[24]), .b(n202) );
    nand2_0 U339 ( .x(___cell__39170_net140213), .a(A[24]), .b(B[24]) );
    inv_1 U34 ( .x(___cell__39170_net140311), .a(A[1]) );
    exor2_1 U340 ( .x(n187), .a(B[17]), .b(A[17]) );
    ao21_1 U341 ( .x(n176), .a(A[8]), .b(B[8]), .c(___cell__39170_net140395)
         );
    inv_0 U342 ( .x(net150837), .a(net150690) );
    inv_3 U343 ( .x(n201), .a(B[9]) );
    nand2_3 U344 ( .x(___cell__39170_net140184), .a(B[9]), .b(A[9]) );
    exnor2_1 U345 ( .x(SUM[8]), .a(___cell__39170_net140270), .b(n176) );
    oai22_1 U346 ( .x(n206), .a(B[21]), .b(A[21]), .c(A[22]), .d(B[22]) );
    nand2_4 U347 ( .x(n154), .a(B[21]), .b(A[21]) );
    mux2i_1 U348 ( .x(n138), .d0(n223), .sl(B[21]), .d1(n224) );
    inv_0 U349 ( .x(n204), .a(B[21]) );
    nor2_1 U35 ( .x(n244), .a(net121836), .b(n73) );
    oai211_1 U350 ( .x(n218), .a(A[17]), .b(B[17]), .c(A[16]), .d(B[16]) );
    nand2_0 U351 ( .x(n161), .a(A[16]), .b(B[16]) );
    nor2i_0 U352 ( .x(n169), .a(n64), .b(___cell__39170_net140236) );
    inv_0 U353 ( .x(___cell__39170_net140471), .a(___cell__39170_net140235) );
    inv_3 U355 ( .x(n213), .a(B[12]) );
    nand2_0 U356 ( .x(___cell__39170_net140235), .a(A[10]), .b(B[10]) );
    exnor2_3 U357 ( .x(SUM[26]), .a(n174), .b(___cell__39170_net140285) );
    nand2i_4 U358 ( .x(n214), .a(n168), .b(n84) );
    exnor2_3 U359 ( .x(n221), .a(n222), .b(n210) );
    nand2i_4 U36 ( .x(___cell__39170_net140259), .a(n92), .b(n125) );
    aoi221_4 U360 ( .x(___cell__39170_net140455), .a(n228), .b(n229), .c(B[22]
        ), .d(n230), .e(n152) );
    nand2i_4 U361 ( .x(___cell__39170_net140476), .a(B[8]), .b(
        ___cell__39170_net140341) );
    mux2i_3 U363 ( .x(n136), .d0(n225), .sl(n90), .d1(n221) );
    nand2_3 U364 ( .x(SUM[18]), .a(n136), .b(n137) );
    aoai211_5 U365 ( .x(n216), .a(n205), .b(n54), .c(net150690), .d(n207) );
    nand2i_6 U366 ( .x(___cell__39170_net140398), .a(B[11]), .b(n215) );
    nand2_8 U367 ( .x(___cell__39170_net140560), .a(n229), .b(n53) );
    inv_6 U368 ( .x(n229), .a(n206) );
    inv_10 U369 ( .x(n195), .a(B[4]) );
    inv_2 U37 ( .x(___cell__39170_net140444), .a(net155899) );
    inv_2 U370 ( .x(net121836), .a(net155900) );
    or2_2 U371 ( .x(n137), .a(n76), .b(n222) );
    inv_3 U372 ( .x(n222), .a(n220) );
    exnor2_1 U373 ( .x(SUM[22]), .a(n181), .b(n248) );
    inv_2 U374 ( .x(n248), .a(n182) );
    aoai211_2 U375 ( .x(n181), .a(n204), .b(n203), .c(n239), .d(n154) );
    ao211_4 U376 ( .x(___cell__39170_net140452), .a(n80), .b(n81), .c(
        ___cell__39170_net140258), .d(___cell__39170_net140259) );
    exnor2_3 U377 ( .x(SUM[11]), .a(n249), .b(___cell__39170_net140231) );
    inv_3 U378 ( .x(n249), .a(n192) );
    ao21_2 U379 ( .x(n192), .a(n193), .b(n60), .c(___cell__39170_net140471) );
    inv_2 U38 ( .x(___cell__39170_net140485), .a(___cell__39170_net140313) );
    nor2i_0 U380 ( .x(___cell__39170_net140231), .a(___cell__39170_net140232), 
        .b(___cell__39170_net140233) );
    inv_2 U381 ( .x(n113), .a(A[10]) );
    ao21_3 U382 ( .x(___cell__39170_net140392), .a(n128), .b(n129), .c(n61) );
    inv_4 U383 ( .x(n129), .a(A[19]) );
    nand4i_2 U384 ( .x(n92), .a(___cell__39170_net140395), .b(
        ___cell__39170_net140396), .c(n60), .d(___cell__39170_net140398) );
    buf_8 U385 ( .x(n60), .a(___cell__39170_net140397) );
    nor3i_4 U386 ( .x(___cell__39170_net140256), .a(___cell__39170_net140257), 
        .b(___cell__39170_net140259), .c(___cell__39170_net140258) );
    inv_0 U387 ( .x(n250), .a(n77) );
    oaoi211_2 U388 ( .x(n74), .a(n78), .b(n77), .c(n76), .d(n75) );
    ao21_4 U389 ( .x(n65), .a(n84), .b(n151), .c(n251) );
    nand2_2 U39 ( .x(___cell__39170_net140484), .a(___cell__39170_net140485), 
        .b(___cell__39170_net140444) );
    inv_0 U390 ( .x(n91), .a(n84) );
    inv_0 U391 ( .x(n165), .a(n251) );
    nor2i_1 U392 ( .x(n251), .a(B[13]), .b(n252) );
    nand2i_2 U393 ( .x(n84), .a(A[13]), .b(n85) );
    inv_1 U394 ( .x(n252), .a(A[13]) );
    inv_2 U40 ( .x(___cell__39170_net140249), .a(___cell__39170_net140484) );
    inv_2 U41 ( .x(net155899), .a(B[1]) );
    nand2i_2 U42 ( .x(n233), .a(net155899), .b(___cell__39170_net140482) );
    inv_2 U43 ( .x(n173), .a(n233) );
    inv_2 U44 ( .x(net152445), .a(___cell__39170_net140316) );
    nand2i_5 U45 ( .x(n232), .a(A[6]), .b(n197) );
    or2_5 U46 ( .x(n145), .a(n86), .b(n197) );
    inv_2 U47 ( .x(___cell__39170_net140351), .a(B[26]) );
    inv_2 U48 ( .x(n102), .a(A[26]) );
    nand2i_2 U49 ( .x(n107), .a(B[26]), .b(n102) );
    nor2i_1 U50 ( .x(n99), .a(B[25]), .b(n101) );
    inv_2 U51 ( .x(n101), .a(n107) );
    nor2i_0 U52 ( .x(n100), .a(A[25]), .b(n101) );
    inv_2 U53 ( .x(___cell__39170_net140233), .a(___cell__39170_net140398) );
    inv_2 U54 ( .x(___cell__39170_net140411), .a(___cell__39170_net140232) );
    nand2_0 U55 ( .x(___cell__39170_net140232), .a(A[11]), .b(B[11]) );
    exor2_1 U56 ( .x(n183), .a(n55), .b(B[20]) );
    inv_2 U57 ( .x(n54), .a(A[20]) );
    nor2i_1 U58 ( .x(n163), .a(___cell__39170_net140223), .b(net152474) );
    nand2_1 U59 ( .x(n167), .a(A[12]), .b(B[12]) );
    nand2i_4 U6 ( .x(___cell__39170_net140513), .a(n92), .b(n198) );
    nand2i_5 U60 ( .x(n150), .a(A[12]), .b(n213) );
    exor2_1 U61 ( .x(n182), .a(A[22]), .b(B[22]) );
    exor2_1 U63 ( .x(n185), .a(A[19]), .b(B[19]) );
    aoi21_1 U64 ( .x(n157), .a(n158), .b(n159), .c(___cell__39170_net140218)
         );
    nor2i_1 U65 ( .x(n158), .a(n76), .b(n72) );
    inv_2 U66 ( .x(n76), .a(n61) );
    inv_2 U68 ( .x(n78), .a(n217) );
    inv_2 U69 ( .x(n75), .a(n219) );
    inv_5 U7 ( .x(___cell__39170_net140514), .a(___cell__39170_net140410) );
    nand2_1 U70 ( .x(___cell__39170_net140210), .a(A[3]), .b(B[3]) );
    nand2i_2 U71 ( .x(___cell__39170_net140499), .a(n121), .b(
        ___cell__39170_net140279) );
    nand2i_2 U72 ( .x(n127), .a(B[3]), .b(n123) );
    inv_2 U73 ( .x(n123), .a(A[3]) );
    inv_2 U74 ( .x(n188), .a(n159) );
    nand2i_2 U75 ( .x(n231), .a(net150555), .b(___cell__39170_net140279) );
    nand2_2 U76 ( .x(n119), .a(B[28]), .b(A[28]) );
    nand2i_4 U77 ( .x(___cell__39170_net140537), .a(___cell__39170_net140463), 
        .b(___cell__39170_net140283) );
    nand2i_2 U78 ( .x(___cell__39170_net140463), .a(n116), .b(B[27]) );
    nand2i_2 U79 ( .x(___cell__39170_net140464), .a(n116), .b(n58) );
    inv_7 U8 ( .x(n89), .a(B[18]) );
    inv_2 U80 ( .x(n117), .a(B[28]) );
    nand2i_2 U81 ( .x(n118), .a(A[28]), .b(n117) );
    inv_2 U82 ( .x(n116), .a(n118) );
    nor2_1 U83 ( .x(n115), .a(n116), .b(___cell__39170_net140255) );
    inv_2 U84 ( .x(___cell__39170_net140268), .a(___cell__39170_net140546) );
    inv_2 U85 ( .x(n110), .a(A[29]) );
    nor2_1 U86 ( .x(n242), .a(net121836), .b(n73) );
    nand2_2 U87 ( .x(n247), .a(n73), .b(net121836) );
    nor2i_1 U88 ( .x(n246), .a(n247), .b(n242) );
    nand2i_2 U89 ( .x(___cell__39170_net140396), .a(A[9]), .b(n201) );
    inv_2 U90 ( .x(___cell__39170_net140447), .a(___cell__39170_net140184) );
    nand2i_0 U91 ( .x(n235), .a(n214), .b(___cell__39170_net140199) );
    nand2i_2 U92 ( .x(n191), .a(n65), .b(n235) );
    nand2_1 U93 ( .x(___cell__39170_net140223), .a(A[14]), .b(B[14]) );
    nand2i_2 U94 ( .x(n159), .a(___cell__39170_net140241), .b(n237) );
    nor2i_1 U95 ( .x(n160), .a(n161), .b(n59) );
    exor2_1 U96 ( .x(SUM[17]), .a(n186), .b(n187) );
    oai21_1 U97 ( .x(n186), .a(n188), .b(n59), .c(n161) );
    inv_2 U98 ( .x(n230), .a(n154) );
    inv_2 U99 ( .x(n239), .a(n216) );
endmodule


module EX_DW01_add_32_0_test_1 ( A, B, CI, SUM, CO );
input  [31:0] A;
input  [31:0] B;
output [31:0] SUM;
input  CI;
output CO;
    wire n119, n301, n79, n323, n109, n287, n289, n191, n115, n332, n116, n192, 
        n325, n333, n165, n63, n167, n280, n139, n279, n272, n185, n302, n93, 
        n95, n248, n113, n281, n285, n286, n154, n155, n156, n246, n105, n276, 
        n106, n253, n173, n259, n158, n260, n261, n136, n252, n206, n238, n235, 
        n153, n241, n236, n347, n170, n257, n108, n80, n198, n148, n209, n51, 
        n233, n234, n121, n126, n174, n175, n176, n216, n120, n124, n122, n123, 
        n125, n87, n270, n201, n202, n217, n177, n157, n208, n214, n168, n353, 
        n172, n169, n354, n215, n171, n258, n255, n256, n218, n180, n335, n194, 
        n129, n130, n131, n134, n334, n133, n160, n210, n195, n132, n150, n329, 
        n149, n326, n118, n162, n211, n349, n348, n200, n59, n317, n193, n283, 
        n284, n53, n356, n339, n117, n212, n213, n112, n137, n358, n242, n204, 
        n240, n237, n232, n247, n359, n318, n361, n363, n290, n88, n227, n52, 
        n296, n189, n364, n110, n337, n54, n319, n55, n164, n94, n166, n56, 
        n223, n365, n57, n220, n221, n273, n77, n239, n274, n152, n300, n268, 
        n346, n205, n308, n146, n352, n101, n103, n143, n104, n295, n128, n96, 
        n74, n97, n303, n190, n263, n271, n135, n58, n84, n315, n188, n322, 
        n60, n228, n321, n362, n92, n73, n61, n98, n203, n91, n62, n64, n293, 
        n127, n294, n65, n311, n312, n338, n249, n68, n71, n345, n72, n265, 
        n226, n343, n304, n342, n344, n83, n82, n81, n288, n307, n145, n147, 
        n78, n75, n350, n336, n76, n275, n324, n357, n244, n243, n292, n360, 
        n330, n291, n309, n250, n224, n222, n163, n178, n179, n138, n140, n187, 
        n219, n114, n264, n245, n254, n102, n199, n111, n151, n99, n277, n161, 
        n100, n262, n196, n310, n182, n183, n144, n141, n207, n320, n282, n299, 
        n305, n306, n142, n107, n351, n50, n197, n66, n266, n297, n298, n278, 
        n184, n340, n341, n181, n366, n231, n367, n368, n313, n314, n331, n49, 
        n159, n316, n186, n355, n251, n269, n229, n327, n225, n328, n230, n67, 
        n69, n70, n89, n85, n86;
    inv_2 U10 ( .x(n119), .a(n301) );
    inv_2 U100 ( .x(n79), .a(n323) );
    mux2i_1 U101 ( .x(n109), .d0(n287), .sl(B[1]), .d1(n289) );
    nand2i_2 U102 ( .x(n191), .a(n115), .b(n332) );
    nor2i_0 U103 ( .x(n115), .a(A[8]), .b(n116) );
    nand2_2 U104 ( .x(n332), .a(n192), .b(n325) );
    inv_2 U105 ( .x(n333), .a(n191) );
    nor2i_1 U107 ( .x(n165), .a(n63), .b(n167) );
    inv_2 U108 ( .x(n280), .a(n139) );
    oai21_1 U109 ( .x(n279), .a(n167), .b(n280), .c(n63) );
    nand3_1 U11 ( .x(n272), .a(n185), .b(n301), .c(n302) );
    nand2_4 U110 ( .x(n93), .a(n95), .b(n248) );
    nand2i_2 U111 ( .x(n113), .a(n281), .b(n279) );
    exnor2_1 U112 ( .x(n285), .a(n286), .b(n95) );
    inv_2 U113 ( .x(n286), .a(n279) );
    inv_8 U114 ( .x(n95), .a(B[17]) );
    nor2i_1 U115 ( .x(n154), .a(n155), .b(n156) );
    nand2_2 U116 ( .x(n155), .a(B[21]), .b(A[21]) );
    inv_2 U117 ( .x(n246), .a(B[21]) );
    inv_2 U118 ( .x(n105), .a(n276) );
    inv_2 U119 ( .x(n106), .a(n253) );
    inv_1 U12 ( .x(n173), .a(n259) );
    inv_2 U120 ( .x(n158), .a(n260) );
    nand2i_2 U121 ( .x(n261), .a(n136), .b(n158) );
    inv_2 U122 ( .x(n252), .a(B[19]) );
    exor2_1 U123 ( .x(n206), .a(B[23]), .b(A[23]) );
    inv_0 U124 ( .x(n238), .a(A[24]) );
    inv_2 U125 ( .x(n235), .a(A[26]) );
    inv_2 U127 ( .x(n153), .a(n241) );
    inv_2 U128 ( .x(n236), .a(A[25]) );
    nand2i_2 U129 ( .x(n347), .a(B[25]), .b(n236) );
    inv_0 U13 ( .x(n170), .a(n257) );
    inv_3 U130 ( .x(n108), .a(n80) );
    exor2_1 U131 ( .x(SUM[3]), .a(n198), .b(n148) );
    exnor2_1 U132 ( .x(SUM[2]), .a(n209), .b(n51) );
    nand2i_2 U133 ( .x(n209), .a(n233), .b(n234) );
    exor2_1 U134 ( .x(SUM[6]), .a(n121), .b(n126) );
    nor2i_1 U135 ( .x(n174), .a(n175), .b(n176) );
    exor2_1 U136 ( .x(SUM[12]), .a(n216), .b(n174) );
    exnor2_1 U137 ( .x(SUM[7]), .a(n120), .b(n124) );
    aoi21_1 U138 ( .x(n120), .a(n121), .b(n122), .c(n123) );
    nor2i_1 U139 ( .x(n124), .a(n125), .b(n87) );
    nand2i_0 U14 ( .x(n259), .a(A[13]), .b(n270) );
    exnor2_1 U140 ( .x(SUM[27]), .a(n201), .b(n202) );
    exor2_1 U141 ( .x(SUM[11]), .a(n217), .b(n177) );
    exnor2_1 U142 ( .x(SUM[20]), .a(n157), .b(n208) );
    exor2_1 U143 ( .x(SUM[14]), .a(n214), .b(n168) );
    oai21_1 U144 ( .x(n214), .a(n173), .b(n353), .c(n172) );
    nor2i_1 U145 ( .x(n168), .a(n169), .b(n170) );
    inv_2 U146 ( .x(n354), .a(n214) );
    exor2_1 U147 ( .x(SUM[13]), .a(n215), .b(n171) );
    inv_2 U148 ( .x(n176), .a(n258) );
    nor2i_1 U149 ( .x(n171), .a(n172), .b(n173) );
    nand4i_1 U15 ( .x(n255), .a(n256), .b(n257), .c(n258), .d(n259) );
    inv_2 U150 ( .x(n353), .a(n215) );
    exor2_1 U151 ( .x(SUM[10]), .a(n218), .b(n180) );
    inv_2 U152 ( .x(n335), .a(n194) );
    nor2i_1 U153 ( .x(n129), .a(n130), .b(n131) );
    oai21_1 U154 ( .x(n194), .a(n134), .b(n334), .c(n133) );
    exor2_1 U155 ( .x(SUM[5]), .a(n194), .b(n129) );
    exnor2_1 U156 ( .x(SUM[19]), .a(n160), .b(n210) );
    exor2_1 U157 ( .x(SUM[4]), .a(n195), .b(n132) );
    oai21_1 U158 ( .x(n195), .a(n150), .b(n329), .c(n149) );
    inv_2 U159 ( .x(n150), .a(n326) );
    nand2_1 U16 ( .x(n118), .a(B[9]), .b(A[9]) );
    inv_2 U160 ( .x(n329), .a(n198) );
    nor2i_1 U161 ( .x(n132), .a(n133), .b(n134) );
    inv_2 U162 ( .x(n334), .a(n195) );
    exnor2_1 U163 ( .x(SUM[18]), .a(n162), .b(n211) );
    inv_2 U164 ( .x(n349), .a(n348) );
    exor2_1 U165 ( .x(n200), .a(B[28]), .b(n59) );
    inv_2 U166 ( .x(n317), .a(n325) );
    exnor2_1 U167 ( .x(SUM[8]), .a(n192), .b(n193) );
    exnor2_1 U168 ( .x(SUM[29]), .a(n283), .b(n284) );
    nand2_2 U169 ( .x(SUM[1]), .a(n109), .b(n53) );
    nand3_1 U17 ( .x(n356), .a(n259), .b(n257), .c(n339) );
    exor2_1 U170 ( .x(SUM[9]), .a(n191), .b(n117) );
    exor2_1 U171 ( .x(SUM[15]), .a(n212), .b(n213) );
    exor2_1 U172 ( .x(SUM[16]), .a(n139), .b(n165) );
    nand2_2 U173 ( .x(SUM[17]), .a(n112), .b(n113) );
    exnor2_1 U174 ( .x(SUM[21]), .a(n137), .b(n154) );
    inv_2 U175 ( .x(n358), .a(n242) );
    nand2i_2 U176 ( .x(n204), .a(n240), .b(n237) );
    inv_2 U177 ( .x(n232), .a(B[9]) );
    inv_2 U178 ( .x(n247), .a(B[16]) );
    inv_0 U179 ( .x(n116), .a(B[8]) );
    nand2i_2 U18 ( .x(n359), .a(n172), .b(n257) );
    inv_2 U180 ( .x(n318), .a(B[28]) );
    or2_2 U181 ( .x(n51), .a(n361), .b(n363) );
    inv_2 U182 ( .x(n290), .a(n87) );
    and2_3 U183 ( .x(n87), .a(n88), .b(n227) );
    aoi21_4 U184 ( .x(n52), .a(n296), .b(n302), .c(n189) );
    or2_2 U185 ( .x(n53), .a(n364), .b(n110) );
    inv_2 U186 ( .x(n156), .a(n337) );
    nand2i_2 U187 ( .x(n337), .a(A[21]), .b(n246) );
    nand2_2 U188 ( .x(n54), .a(n348), .b(n319) );
    nand2_2 U189 ( .x(n55), .a(n348), .b(n318) );
    oai22_3 U190 ( .x(n164), .a(n95), .b(n248), .c(n94), .d(n166) );
    ao21_4 U191 ( .x(n56), .a(n363), .b(n223), .c(n365) );
    inv_2 U192 ( .x(n363), .a(n364) );
    and4_3 U193 ( .x(n57), .a(n326), .b(n122), .c(n220), .d(n221) );
    inv_2 U194 ( .x(n273), .a(n77) );
    oa211_2 U195 ( .x(n77), .a(n239), .b(n242), .c(n274), .d(n152) );
    exor2_1 U196 ( .x(n213), .a(B[15]), .b(A[15]) );
    nand2i_2 U197 ( .x(n300), .a(B[15]), .b(n268) );
    nand2i_0 U198 ( .x(n346), .a(B[24]), .b(n238) );
    exor2_1 U199 ( .x(n205), .a(B[24]), .b(A[24]) );
    nor2i_3 U200 ( .x(n308), .a(A[30]), .b(n146) );
    inv_4 U201 ( .x(n146), .a(n352) );
    exnor2_1 U202 ( .x(SUM[23]), .a(n101), .b(n206) );
    aoi21_1 U203 ( .x(n157), .a(n158), .b(n139), .c(n103) );
    oai21_3 U204 ( .x(n143), .a(n156), .b(n104), .c(n155) );
    ao211_5 U205 ( .x(n295), .a(n133), .b(n130), .c(n128), .d(n131) );
    aoai211_4 U206 ( .x(n96), .a(n55), .b(n54), .c(n74), .d(n97) );
    inv_2 U207 ( .x(n59), .a(n319) );
    inv_2 U208 ( .x(n319), .a(A[28]) );
    nor3_2 U209 ( .x(n303), .a(n190), .b(n263), .c(n271) );
    nor2_0 U21 ( .x(n135), .a(A[19]), .b(B[19]) );
    aoi21_3 U210 ( .x(n190), .a(n58), .b(A[0]), .c(n84) );
    nand2i_2 U211 ( .x(n315), .a(n189), .b(n188) );
    ao21_1 U212 ( .x(n201), .a(n108), .b(n322), .c(n273) );
    nand2_0 U213 ( .x(n172), .a(B[13]), .b(A[13]) );
    oai22_2 U214 ( .x(n60), .a(n95), .b(n248), .c(n166), .d(n94) );
    inv_7 U215 ( .x(n94), .a(n93) );
    inv_2 U216 ( .x(n228), .a(A[5]) );
    nand2i_4 U217 ( .x(n321), .a(B[29]), .b(n96) );
    nor2i_0 U218 ( .x(n289), .a(n110), .b(A[1]) );
    nor2_0 U219 ( .x(n362), .a(B[1]), .b(A[1]) );
    inv_3 U22 ( .x(n92), .a(n60) );
    exnor2_1 U220 ( .x(n287), .a(A[1]), .b(n110) );
    nand2_2 U221 ( .x(n364), .a(B[1]), .b(A[1]) );
    inv_2 U222 ( .x(n73), .a(A[3]) );
    exnor2_3 U223 ( .x(SUM[26]), .a(n61), .b(n98) );
    ao21_3 U224 ( .x(n61), .a(n203), .b(n347), .c(n91) );
    inv_0 U225 ( .x(n62), .a(n166) );
    inv_2 U226 ( .x(n63), .a(n62) );
    nand2_4 U227 ( .x(n166), .a(B[16]), .b(A[16]) );
    inv_0 U228 ( .x(n64), .a(n248) );
    inv_6 U229 ( .x(n248), .a(A[17]) );
    nor2i_2 U23 ( .x(n293), .a(n127), .b(n294) );
    nor2_3 U230 ( .x(n65), .a(A[10]), .b(B[10]) );
    aoai211_1 U231 ( .x(n311), .a(A[0]), .b(n58), .c(n84), .d(n312) );
    nand2i_1 U232 ( .x(n338), .a(A[16]), .b(n247) );
    inv_0 U233 ( .x(n167), .a(n338) );
    inv_0 U234 ( .x(n249), .a(A[18]) );
    nand2_2 U235 ( .x(n133), .a(A[4]), .b(B[4]) );
    exnor2_1 U236 ( .x(SUM[25]), .a(n203), .b(n204) );
    inv_2 U237 ( .x(n68), .a(n293) );
    nand2_0 U238 ( .x(n71), .a(B[9]), .b(A[9]) );
    ao211_5 U239 ( .x(n345), .a(n188), .b(n72), .c(n263), .d(n265) );
    nand2_0 U24 ( .x(n125), .a(A[7]), .b(B[7]) );
    inv_0 U240 ( .x(n72), .a(n189) );
    inv_2 U241 ( .x(n188), .a(A[8]) );
    inv_8 U242 ( .x(n226), .a(A[6]) );
    nand4_3 U243 ( .x(n343), .a(n304), .b(n342), .c(n345), .d(n344) );
    oaoi211_2 U245 ( .x(n80), .a(n83), .b(n82), .c(n343), .d(n81) );
    nor2i_0 U246 ( .x(n288), .a(B[17]), .b(n279) );
    nor2i_3 U247 ( .x(n307), .a(n145), .b(n147) );
    oaoi211_3 U248 ( .x(n74), .a(n80), .b(n78), .c(n77), .d(n75) );
    inv_0 U249 ( .x(n350), .a(n74) );
    inv_1 U25 ( .x(n123), .a(n127) );
    inv_2 U250 ( .x(n75), .a(n336) );
    nand2_2 U251 ( .x(n336), .a(n76), .b(n275) );
    inv_0 U252 ( .x(n76), .a(B[27]) );
    nor2i_3 U253 ( .x(n78), .a(n324), .b(n79) );
    inv_2 U254 ( .x(n81), .a(n357) );
    inv_2 U255 ( .x(n82), .a(n244) );
    inv_2 U256 ( .x(n83), .a(n243) );
    inv_0 U257 ( .x(n275), .a(A[27]) );
    nand2i_2 U258 ( .x(n274), .a(n237), .b(n241) );
    nand2_0 U259 ( .x(n152), .a(A[26]), .b(B[26]) );
    nand2i_2 U26 ( .x(n292), .a(n149), .b(n220) );
    nand2_0 U260 ( .x(n242), .a(B[24]), .b(A[24]) );
    nand2i_2 U261 ( .x(n239), .a(n240), .b(n241) );
    nand2_1 U262 ( .x(n324), .a(n360), .b(A[24]) );
    nand2_0 U264 ( .x(n357), .a(B[23]), .b(A[23]) );
    inv_0 U265 ( .x(n244), .a(B[23]) );
    inv_0 U266 ( .x(n243), .a(A[23]) );
    inv_0 U267 ( .x(n330), .a(n84) );
    inv_2 U268 ( .x(n88), .a(B[7]) );
    nand2i_2 U27 ( .x(n291), .a(n128), .b(n221) );
    inv_0 U270 ( .x(n227), .a(A[7]) );
    inv_0 U271 ( .x(n233), .a(n223) );
    inv_2 U272 ( .x(n91), .a(n237) );
    nand2_0 U273 ( .x(n237), .a(A[25]), .b(B[25]) );
    inv_2 U274 ( .x(n240), .a(n347) );
    exnor2_1 U275 ( .x(n284), .a(B[29]), .b(A[29]) );
    exor2_1 U276 ( .x(n208), .a(A[20]), .b(B[20]) );
    nor2_0 U277 ( .x(n136), .a(A[20]), .b(B[20]) );
    nor2i_3 U278 ( .x(n309), .a(n145), .b(n147) );
    oai21_3 U279 ( .x(n250), .a(A[18]), .b(n164), .c(B[18]) );
    nor2i_1 U28 ( .x(n224), .a(n290), .b(n222) );
    aoi21_1 U280 ( .x(n162), .a(n163), .b(n139), .c(n164) );
    nor2i_0 U281 ( .x(n117), .a(n71), .b(n119) );
    oai21_1 U282 ( .x(n218), .a(n333), .b(n119), .c(n71) );
    nor2i_1 U283 ( .x(n177), .a(n178), .b(n179) );
    inv_0 U284 ( .x(n281), .a(n94) );
    exor2_1 U285 ( .x(SUM[24]), .a(n108), .b(n205) );
    ao21_3 U286 ( .x(n203), .a(n346), .b(n108), .c(n358) );
    aoi21_1 U287 ( .x(n137), .a(n138), .b(n139), .c(n140) );
    ao21_1 U288 ( .x(n193), .a(A[8]), .b(B[8]), .c(n317) );
    nor2_0 U289 ( .x(n187), .a(B[8]), .b(A[8]) );
    or3i_2 U29 ( .x(n222), .a(n223), .b(n219), .c(n114) );
    nand2i_2 U290 ( .x(n264), .a(B[22]), .b(n245) );
    nand2i_3 U291 ( .x(n185), .a(B[11]), .b(n254) );
    inv_2 U292 ( .x(n97), .a(n102) );
    exor2_1 U293 ( .x(SUM[28]), .a(n199), .b(n200) );
    nor2_0 U294 ( .x(n111), .a(A[0]), .b(B[0]) );
    and3i_1 U295 ( .x(n361), .a(n362), .b(B[0]), .c(A[0]) );
    nand2_0 U296 ( .x(n110), .a(A[0]), .b(B[0]) );
    mux2i_1 U297 ( .x(n112), .d0(n288), .sl(n64), .d1(n285) );
    exor2_1 U298 ( .x(n211), .a(B[18]), .b(A[18]) );
    inv_2 U299 ( .x(n98), .a(n151) );
    inv_2 U30 ( .x(n360), .a(n239) );
    nor2i_1 U300 ( .x(n151), .a(n152), .b(n153) );
    inv_0 U301 ( .x(n99), .a(n277) );
    oai21_5 U302 ( .x(n161), .a(n92), .b(n249), .c(n250) );
    nand2_5 U303 ( .x(n344), .a(n143), .b(n264) );
    nor2i_3 U304 ( .x(n100), .a(n337), .b(n261) );
    inv_0 U305 ( .x(n262), .a(n100) );
    inv_0 U306 ( .x(n138), .a(n261) );
    inv_0 U307 ( .x(n101), .a(n343) );
    ao221_4 U308 ( .x(n196), .a(n308), .b(n307), .c(n310), .d(n309), .e(n182)
         );
    nor2i_3 U309 ( .x(n310), .a(B[30]), .b(n146) );
    inv_2 U31 ( .x(n183), .a(A[30]) );
    and3i_1 U310 ( .x(n144), .a(n147), .b(n145), .c(n352) );
    exnor2_1 U311 ( .x(SUM[22]), .a(n141), .b(n207) );
    nor2_0 U312 ( .x(n163), .a(n94), .b(n167) );
    nand2i_0 U313 ( .x(n145), .a(B[29]), .b(n320) );
    exnor2_3 U314 ( .x(SUM[30]), .a(n144), .b(n282) );
    aoi22_2 U315 ( .x(n304), .a(n299), .b(n305), .c(n306), .d(n303) );
    nor2i_0 U316 ( .x(n141), .a(n142), .b(n143) );
    exnor2_5 U317 ( .x(SUM[31]), .a(n196), .b(n107) );
    inv_2 U318 ( .x(n102), .a(n351) );
    nand2i_0 U319 ( .x(n351), .a(B[28]), .b(n319) );
    nor2i_1 U32 ( .x(n182), .a(B[30]), .b(n183) );
    buf_1 U320 ( .x(n103), .a(n50) );
    inv_0 U321 ( .x(n140), .a(n104) );
    nand2_0 U322 ( .x(n276), .a(A[20]), .b(B[20]) );
    inv_0 U323 ( .x(n253), .a(B[20]) );
    nand2i_0 U324 ( .x(n199), .a(n349), .b(n350) );
    inv_2 U325 ( .x(n107), .a(n197) );
    exor2_1 U326 ( .x(n197), .a(B[31]), .b(A[31]) );
    aoi21_1 U327 ( .x(n160), .a(n66), .b(n139), .c(n99) );
    inv_0 U328 ( .x(n283), .a(n96) );
    nand2i_4 U329 ( .x(n352), .a(A[29]), .b(n96) );
    inv_5 U33 ( .x(n147), .a(n321) );
    nand3i_5 U330 ( .x(n265), .a(n52), .b(n185), .c(n266) );
    nand2i_4 U331 ( .x(n271), .a(n272), .b(n266) );
    nand2_2 U332 ( .x(n297), .a(n298), .b(n169) );
    nor2i_5 U333 ( .x(n299), .a(n300), .b(n263) );
    nand2i_4 U334 ( .x(n278), .a(n252), .b(n161) );
    nand2i_4 U335 ( .x(n216), .a(n184), .b(n340) );
    inv_5 U336 ( .x(n341), .a(n216) );
    oai21_4 U337 ( .x(n215), .a(n341), .b(n176), .c(n175) );
    oai21_4 U338 ( .x(n212), .a(n170), .b(n354), .c(n169) );
    nand3i_3 U339 ( .x(n305), .a(n297), .b(n359), .c(n356) );
    inv_2 U34 ( .x(n256), .a(n300) );
    inv_5 U340 ( .x(n312), .a(n271) );
    nand2_8 U341 ( .x(n181), .a(B[10]), .b(A[10]) );
    nand2_6 U342 ( .x(n175), .a(B[12]), .b(A[12]) );
    nand2_8 U343 ( .x(n348), .a(A[27]), .b(B[27]) );
    nand2i_6 U345 ( .x(n301), .a(A[9]), .b(n232) );
    inv_6 U347 ( .x(n277), .a(n161) );
    nand2_4 U348 ( .x(n342), .a(A[22]), .b(B[22]) );
    inv_0 U35 ( .x(n268), .a(A[15]) );
    inv_6 U352 ( .x(n266), .a(n255) );
    nor2i_2 U353 ( .x(n296), .a(B[8]), .b(n119) );
    nor2_1 U354 ( .x(n365), .a(n366), .b(n231) );
    inv_0 U355 ( .x(n234), .a(n365) );
    inv_0 U356 ( .x(n366), .a(B[2]) );
    inv_3 U357 ( .x(n231), .a(A[2]) );
    nor2i_3 U358 ( .x(n367), .a(n368), .b(A[14]) );
    inv_4 U359 ( .x(n257), .a(n367) );
    aoi22_1 U36 ( .x(n313), .a(n305), .b(n300), .c(n314), .d(n315) );
    inv_0 U360 ( .x(n368), .a(B[14]) );
    nand2i_4 U361 ( .x(n221), .a(B[5]), .b(n228) );
    nand2_2 U362 ( .x(n130), .a(A[5]), .b(B[5]) );
    nand2_3 U363 ( .x(n169), .a(A[14]), .b(B[14]) );
    nand2_1 U364 ( .x(n298), .a(B[15]), .b(A[15]) );
    nand2i_4 U365 ( .x(n122), .a(B[6]), .b(n226) );
    nand2_2 U366 ( .x(n127), .a(A[6]), .b(B[6]) );
    nand2i_0 U367 ( .x(n241), .a(B[26]), .b(n235) );
    nand2_1 U368 ( .x(n323), .a(n360), .b(B[24]) );
    and2_2 U37 ( .x(n58), .a(n224), .b(n57) );
    inv_2 U38 ( .x(n245), .a(A[22]) );
    inv_2 U39 ( .x(n314), .a(n265) );
    nand2_2 U40 ( .x(n263), .a(n100), .b(n264) );
    oai211_1 U41 ( .x(n189), .a(n65), .b(n118), .c(n178), .d(n181) );
    nand2i_2 U42 ( .x(n306), .a(B[8]), .b(n188) );
    nor2i_0 U43 ( .x(n148), .a(n149), .b(n150) );
    inv_2 U44 ( .x(n219), .a(B[0]) );
    nand2i_2 U45 ( .x(n223), .a(B[2]), .b(n231) );
    nor2i_0 U46 ( .x(n126), .a(n127), .b(n128) );
    inv_5 U48 ( .x(n128), .a(n122) );
    nand2_1 U49 ( .x(n192), .a(n330), .b(n331) );
    inv_0 U5 ( .x(n49), .a(n159) );
    nand3i_1 U50 ( .x(n316), .a(n317), .b(n185), .c(n302) );
    or3i_2 U51 ( .x(n340), .a(n192), .b(n119), .c(n316) );
    inv_2 U52 ( .x(n302), .a(n65) );
    inv_2 U53 ( .x(n186), .a(n315) );
    nor3i_1 U54 ( .x(n184), .a(n185), .b(n186), .c(n52) );
    inv_2 U55 ( .x(n294), .a(n125) );
    oai21_1 U56 ( .x(n121), .a(n131), .b(n335), .c(n130) );
    inv_2 U57 ( .x(n131), .a(n221) );
    nand2_2 U58 ( .x(n202), .a(n336), .b(n348) );
    nand2_2 U59 ( .x(n322), .a(n323), .b(n324) );
    inv_2 U6 ( .x(n50), .a(n49) );
    nor2i_1 U60 ( .x(SUM[0]), .a(n110), .b(n111) );
    inv_2 U61 ( .x(n254), .a(A[11]) );
    inv_2 U62 ( .x(n179), .a(n185) );
    nand2_2 U63 ( .x(n178), .a(A[11]), .b(B[11]) );
    oai21_1 U64 ( .x(n217), .a(n65), .b(n355), .c(n181) );
    inv_0 U65 ( .x(n251), .a(A[19]) );
    nand2i_2 U66 ( .x(n260), .a(n135), .b(n66) );
    inv_0 U67 ( .x(n270), .a(B[13]) );
    nand2i_2 U68 ( .x(n258), .a(A[12]), .b(n269) );
    inv_0 U69 ( .x(n269), .a(B[12]) );
    aoai211_3 U7 ( .x(n159), .a(n277), .b(n252), .c(n251), .d(n278) );
    inv_2 U70 ( .x(n339), .a(n175) );
    nor2i_1 U71 ( .x(n180), .a(n181), .b(n65) );
    inv_2 U72 ( .x(n355), .a(n218) );
    exor2_1 U73 ( .x(n207), .a(A[22]), .b(B[22]) );
    nand2i_1 U74 ( .x(n142), .a(n262), .b(n139) );
    exor2_1 U76 ( .x(n210), .a(A[19]), .b(B[19]) );
    oa211_3 U77 ( .x(n66), .a(A[18]), .b(B[18]), .c(n93), .d(n338) );
    inv_0 U78 ( .x(n134), .a(n220) );
    inv_2 U79 ( .x(n229), .a(A[4]) );
    oaoi211_2 U8 ( .x(n104), .a(A[20]), .b(n106), .c(n159), .d(n105) );
    nand2i_2 U80 ( .x(n220), .a(B[4]), .b(n229) );
    nand2i_2 U81 ( .x(n198), .a(n56), .b(n327) );
    nand2i_2 U82 ( .x(n327), .a(n225), .b(n328) );
    inv_0 U83 ( .x(n328), .a(n222) );
    nand2i_2 U84 ( .x(n326), .a(B[3]), .b(n230) );
    inv_0 U85 ( .x(n230), .a(A[3]) );
    nand2i_2 U86 ( .x(n149), .a(n73), .b(B[3]) );
    oai21_2 U87 ( .x(n139), .a(n187), .b(n311), .c(n313) );
    exnor2_1 U88 ( .x(n282), .a(B[30]), .b(A[30]) );
    inv_2 U89 ( .x(n320), .a(A[29]) );
    nor2_0 U9 ( .x(n114), .a(B[1]), .b(A[1]) );
    nand2i_2 U90 ( .x(n325), .a(B[8]), .b(n188) );
    inv_2 U91 ( .x(n67), .a(n295) );
    inv_2 U92 ( .x(n69), .a(n292) );
    inv_2 U93 ( .x(n70), .a(n291) );
    aoi211_1 U94 ( .x(n89), .a(n70), .b(n69), .c(n68), .d(n67) );
    inv_2 U95 ( .x(n85), .a(n56) );
    inv_2 U96 ( .x(n86), .a(n57) );
    oaoi211_1 U97 ( .x(n84), .a(n86), .b(n85), .c(n89), .d(n87) );
    nand2i_2 U98 ( .x(n331), .a(n225), .b(n58) );
    inv_0 U99 ( .x(n225), .a(A[0]) );
endmodule


module EX_DW01_sub_32_0_test_1 ( A, B, CI, DIFF, CO );
input  [31:0] A;
input  [31:0] B;
output [31:0] DIFF;
input  CI;
output CO;
    wire n298, n175, n186, n111, n116, n313, n85, n206, n74, n187, n112, n113, 
        n204, n194, n195, n329, n328, n272, n327, n61, n249, n285, n282, n283, 
        n314, n130, n178, n179, n242, n81, n332, n147, n296, n247, n126, n148, 
        n157, n158, n71, n89, n160, n324, n237, n228, n164, n52, n201, n159, 
        n284, n161, n227, n166, n84, n165, n79, n286, n127, n141, n51, n125, 
        n128, n142, n143, n244, n188, n117, n211, n311, n304, n303, n189, n104, 
        n118, n305, n156, n224, n205, n149, n91, n274, n150, n151, n246, n190, 
        n180, n309, n100, n152, n291, n223, n236, n101, n256, n153, n94, n260, 
        n129, n131, n269, n185, n108, n307, n121, n109, n110, n240, n193, n58, 
        n192, n184, n105, n231, n106, n107, n239, n230, n312, n154, n155, n96, 
        n275, n221, n144, n145, n146, n273, n270, n271, n215, n140, n216, n138, 
        n139, n316, n214, n136, n219, n137, n251, n191, n132, n50, n217, n54, 
        n56, n53, n297, n57, n254, n212, n317, n60, n133, n281, n93, n259, 
        n261, n262, n99, n92, n95, n122, n170, n245, n229, n119, n243, n277, 
        n225, n290, n82, n59, n326, n77, n62, n55, n287, n292, n73, n330, n97, 
        n333, n63, n90, n64, n65, n66, n67, n252, n68, n182, n183, n69, n70, 
        n174, n218, n72, n76, n80, n234, n293, n257, n295, n75, n315, n294, 
        n98, n320, n253, n266, n78, n267, n172, n173, n120, n167, n168, n169, 
        n200, n83, n222, n299, n86, n87, n88, n102, n103, n123, n124, n135, 
        n171, n258, n196, n197, n238, n241, n263, n264, n265, n268, n276, n310, 
        n210, n306, n318, n323, n202, n325, n203, n220, n322, n255, n334, n279, 
        n181, n331, n300, n335, n235, n336, n233, n226, n319, n308, n208, n301, 
        n289, n134, n177, n250, n213, n302, n280, n209, n278, n248, n176, n321, 
        n198, n199, n207, n114, n115, n162, n163;
    inv_1 U10 ( .x(n298), .a(n175) );
    exor2_1 U100 ( .x(DIFF[7]), .a(n186), .b(n111) );
    oai21_1 U101 ( .x(n186), .a(n116), .b(n313), .c(n85) );
    inv_2 U102 ( .x(n206), .a(n74) );
    inv_2 U103 ( .x(n313), .a(n187) );
    nor2i_1 U104 ( .x(n111), .a(n112), .b(n113) );
    inv_2 U105 ( .x(n113), .a(n204) );
    exnor2_1 U106 ( .x(DIFF[27]), .a(n194), .b(n195) );
    aoai211_1 U107 ( .x(n194), .a(n329), .b(n328), .c(n272), .d(n327) );
    inv_2 U108 ( .x(n272), .a(n61) );
    inv_2 U109 ( .x(n327), .a(n249) );
    nand2_2 U11 ( .x(n285), .a(n282), .b(n283) );
    nand2_2 U110 ( .x(n195), .a(n314), .b(n130) );
    nand2_2 U111 ( .x(DIFF[0]), .a(n178), .b(n179) );
    inv_2 U112 ( .x(n242), .a(n81) );
    exor2_1 U113 ( .x(DIFF[20]), .a(n332), .b(n147) );
    inv_2 U115 ( .x(n296), .a(n247) );
    nor2_1 U116 ( .x(n147), .a(n126), .b(n148) );
    nor2_1 U117 ( .x(n157), .a(n158), .b(n71) );
    oai21_1 U118 ( .x(n89), .a(n160), .b(n324), .c(n237) );
    exor2_1 U119 ( .x(DIFF[14]), .a(n89), .b(n157) );
    nand2i_2 U12 ( .x(n228), .a(n164), .b(n52) );
    exor2_1 U120 ( .x(DIFF[13]), .a(n201), .b(n159) );
    inv_2 U121 ( .x(n164), .a(n284) );
    nor2_1 U122 ( .x(n159), .a(n160), .b(n161) );
    inv_2 U123 ( .x(n160), .a(n227) );
    inv_2 U124 ( .x(n161), .a(n237) );
    inv_2 U125 ( .x(n324), .a(n201) );
    inv_0 U126 ( .x(n166), .a(n84) );
    nor2_0 U127 ( .x(n165), .a(n81), .b(n166) );
    inv_2 U13 ( .x(n79), .a(n286) );
    exnor2_1 U130 ( .x(DIFF[22]), .a(n127), .b(n141) );
    aoi21_1 U131 ( .x(n127), .a(n51), .b(n125), .c(n128) );
    nor2i_1 U132 ( .x(n141), .a(n142), .b(n143) );
    inv_2 U133 ( .x(n143), .a(n244) );
    exor2_1 U134 ( .x(DIFF[5]), .a(n188), .b(n117) );
    oai21_1 U135 ( .x(n188), .a(n211), .b(n311), .c(n304) );
    inv_2 U136 ( .x(n211), .a(n303) );
    inv_5 U137 ( .x(n311), .a(n189) );
    nor2_1 U138 ( .x(n117), .a(n104), .b(n118) );
    inv_2 U139 ( .x(n104), .a(n305) );
    inv_2 U14 ( .x(n156), .a(n224) );
    inv_2 U140 ( .x(n118), .a(n205) );
    mux2i_1 U141 ( .x(DIFF[19]), .d0(n149), .sl(n91), .d1(n274) );
    aoi21_1 U142 ( .x(n149), .a(A[19]), .b(n150), .c(n151) );
    inv_0 U143 ( .x(n150), .a(B[19]) );
    inv_2 U144 ( .x(n151), .a(n246) );
    exor2_1 U145 ( .x(n274), .a(B[19]), .b(A[19]) );
    exnor2_1 U146 ( .x(DIFF[4]), .a(n189), .b(n190) );
    nand2i_4 U147 ( .x(n189), .a(n180), .b(n309) );
    nand2_2 U148 ( .x(n190), .a(n304), .b(n303) );
    exnor2_1 U149 ( .x(DIFF[18]), .a(n100), .b(n152) );
    oai22_1 U15 ( .x(n291), .a(n223), .b(n237), .c(n156), .d(n236) );
    inv_0 U150 ( .x(n101), .a(n256) );
    nor2_1 U151 ( .x(n152), .a(n153), .b(n94) );
    inv_2 U152 ( .x(n94), .a(n260) );
    nor2i_0 U153 ( .x(n129), .a(n130), .b(n131) );
    exnor2_1 U154 ( .x(n269), .a(A[28]), .b(B[28]) );
    exnor2_1 U155 ( .x(DIFF[8]), .a(n185), .b(n108) );
    inv_2 U156 ( .x(n307), .a(n121) );
    nor2_1 U157 ( .x(n108), .a(n109), .b(n110) );
    inv_2 U158 ( .x(n110), .a(n240) );
    exor2_1 U159 ( .x(n193), .a(B[29]), .b(n58) );
    exor2_1 U160 ( .x(DIFF[29]), .a(n192), .b(n193) );
    exor2_1 U161 ( .x(DIFF[9]), .a(n184), .b(n105) );
    inv_2 U162 ( .x(n109), .a(n231) );
    nor2_1 U163 ( .x(n105), .a(n106), .b(n107) );
    inv_2 U164 ( .x(n106), .a(n239) );
    inv_2 U165 ( .x(n107), .a(n230) );
    inv_2 U166 ( .x(n312), .a(n184) );
    nor2i_1 U167 ( .x(n154), .a(n155), .b(n156) );
    exnor2_1 U168 ( .x(DIFF[17]), .a(n96), .b(n275) );
    inv_2 U169 ( .x(n126), .a(n221) );
    nor2i_1 U170 ( .x(n144), .a(n145), .b(n146) );
    exnor2_1 U171 ( .x(DIFF[23]), .a(n272), .b(n273) );
    exor2_1 U172 ( .x(DIFF[24]), .a(n270), .b(n271) );
    inv_2 U173 ( .x(n215), .a(A[23]) );
    inv_2 U174 ( .x(n140), .a(n216) );
    nor2i_1 U175 ( .x(n138), .a(n139), .b(n140) );
    inv_2 U176 ( .x(n316), .a(n214) );
    inv_2 U177 ( .x(n136), .a(n219) );
    inv_2 U178 ( .x(n137), .a(n251) );
    exor2_1 U179 ( .x(DIFF[3]), .a(n191), .b(n132) );
    inv_2 U180 ( .x(n236), .a(n71) );
    and2_1 U181 ( .x(n50), .a(n216), .b(n217) );
    and3_5 U183 ( .x(n54), .a(n204), .b(n205), .c(n206) );
    ao221_1 U184 ( .x(n56), .a(n296), .b(n53), .c(n128), .d(n244), .e(n297) );
    inv_2 U186 ( .x(n57), .a(n254) );
    inv_2 U187 ( .x(n254), .a(A[30]) );
    inv_2 U188 ( .x(n58), .a(n212) );
    inv_10 U189 ( .x(n131), .a(n317) );
    inv_2 U19 ( .x(n84), .a(n60) );
    nand2i_1 U190 ( .x(n133), .a(B[3]), .b(A[3]) );
    nand2i_2 U191 ( .x(n281), .a(A[3]), .b(B[3]) );
    nand3_1 U192 ( .x(n93), .a(n259), .b(n261), .c(n262) );
    nand2i_6 U193 ( .x(n259), .a(B[17]), .b(n99) );
    nand2i_3 U194 ( .x(n303), .a(A[4]), .b(B[4]) );
    aoi211_1 U195 ( .x(n91), .a(n92), .b(n93), .c(n94), .d(n95) );
    inv_2 U196 ( .x(n153), .a(n92) );
    and3i_1 U197 ( .x(n95), .a(n122), .b(n92), .c(n101) );
    nand2_2 U198 ( .x(n170), .a(n92), .b(n246) );
    nand2_2 U199 ( .x(n245), .a(n92), .b(n246) );
    nand4i_1 U20 ( .x(n229), .a(n119), .b(n84), .c(n230), .d(n231) );
    inv_0 U200 ( .x(n243), .a(A[11]) );
    exnor2_1 U201 ( .x(n277), .a(A[11]), .b(B[11]) );
    nand2i_2 U202 ( .x(n240), .a(B[8]), .b(A[8]) );
    nand2i_2 U203 ( .x(n204), .a(A[7]), .b(B[7]) );
    exnor2_1 U204 ( .x(DIFF[28]), .a(n129), .b(n269) );
    or3i_1 U205 ( .x(n286), .a(n227), .b(n225), .c(n223) );
    inv_2 U208 ( .x(n290), .a(n155) );
    nor2i_2 U209 ( .x(n60), .a(n82), .b(n59) );
    nand2i_2 U21 ( .x(n328), .a(n215), .b(n326) );
    inv_0 U210 ( .x(n59), .a(B[10]) );
    inv_2 U211 ( .x(n82), .a(A[10]) );
    ao211_1 U212 ( .x(n61), .a(n77), .b(n62), .c(n56), .d(n55) );
    nand4_3 U213 ( .x(n62), .a(n287), .b(n292), .c(n73), .d(n330) );
    nand4_1 U214 ( .x(n97), .a(n73), .b(n292), .c(n333), .d(n330) );
    inv_2 U215 ( .x(n122), .a(n97) );
    nand2_1 U216 ( .x(n260), .a(n63), .b(A[18]) );
    inv_0 U217 ( .x(n63), .a(B[18]) );
    nand2i_3 U218 ( .x(n90), .a(A[14]), .b(B[14]) );
    nor2i_1 U219 ( .x(n64), .a(n65), .b(n212) );
    nand2i_2 U22 ( .x(n329), .a(B[23]), .b(n326) );
    inv_0 U220 ( .x(n65), .a(B[29]) );
    nor2_1 U221 ( .x(n66), .a(n212), .b(n67) );
    inv_2 U222 ( .x(n67), .a(n252) );
    ao21_6 U223 ( .x(n68), .a(n182), .b(n183), .c(n131) );
    and2_1 U224 ( .x(n69), .a(n65), .b(n252) );
    ao21_6 U225 ( .x(n70), .a(n182), .b(n183), .c(n131) );
    inv_2 U226 ( .x(n212), .a(A[29]) );
    nand2i_0 U227 ( .x(n252), .a(A[28]), .b(B[28]) );
    nand2i_2 U228 ( .x(n261), .a(B[17]), .b(A[17]) );
    nor3i_2 U229 ( .x(n174), .a(A[17]), .b(B[17]), .c(n175) );
    inv_2 U23 ( .x(n326), .a(n218) );
    nor2i_3 U230 ( .x(n71), .a(n72), .b(n76) );
    inv_0 U231 ( .x(n72), .a(B[14]) );
    aoi31_3 U232 ( .x(n73), .a(n80), .b(n234), .c(n293), .d(n79) );
    exnor2_1 U233 ( .x(n275), .a(B[17]), .b(A[17]) );
    nand2i_0 U234 ( .x(n257), .a(A[17]), .b(B[17]) );
    nand2i_2 U235 ( .x(n295), .a(A[17]), .b(B[17]) );
    nand2i_2 U236 ( .x(n305), .a(B[5]), .b(A[5]) );
    nand2i_2 U237 ( .x(n205), .a(A[5]), .b(B[5]) );
    nor2_3 U238 ( .x(n74), .a(A[6]), .b(n75) );
    nand2_2 U239 ( .x(n85), .a(n75), .b(A[6]) );
    nand2_2 U24 ( .x(n218), .a(n50), .b(n219) );
    inv_0 U240 ( .x(n158), .a(n90) );
    inv_0 U241 ( .x(n76), .a(A[14]) );
    nand2i_0 U242 ( .x(n179), .a(B[0]), .b(A[0]) );
    nand2i_2 U243 ( .x(n92), .a(A[18]), .b(B[18]) );
    ao211_5 U244 ( .x(n315), .a(n77), .b(n62), .c(n56), .d(n55) );
    nand4i_1 U245 ( .x(n294), .a(n245), .b(n53), .c(n98), .d(n295) );
    exnor2_1 U246 ( .x(n271), .a(A[24]), .b(B[24]) );
    nand2i_2 U247 ( .x(n217), .a(A[24]), .b(B[24]) );
    nand2i_2 U249 ( .x(n320), .a(B[30]), .b(n253) );
    nand2i_2 U25 ( .x(n247), .a(B[19]), .b(A[19]) );
    exnor2_3 U250 ( .x(DIFF[31]), .a(n266), .b(n78) );
    inv_2 U251 ( .x(n78), .a(n267) );
    exnor2_1 U252 ( .x(n267), .a(A[31]), .b(B[31]) );
    nand2i_2 U253 ( .x(n231), .a(A[8]), .b(B[8]) );
    nand2i_3 U254 ( .x(n239), .a(B[9]), .b(A[9]) );
    aoai211_1 U255 ( .x(n172), .a(n182), .b(n183), .c(n131), .d(n69) );
    aoai211_1 U256 ( .x(n173), .a(n182), .b(n183), .c(n131), .d(n66) );
    aoai211_1 U257 ( .x(n192), .a(n182), .b(n183), .c(n131), .d(n252) );
    or2_6 U258 ( .x(n80), .a(n120), .b(n121) );
    inv_4 U259 ( .x(n293), .a(n228) );
    aoi21_1 U26 ( .x(n167), .a(n168), .b(n169), .c(n170) );
    exnor2_1 U260 ( .x(DIFF[16]), .a(n97), .b(n200) );
    aoi21_1 U262 ( .x(n96), .a(n97), .b(n98), .c(n99) );
    aoi21_1 U263 ( .x(n100), .a(n101), .b(n97), .c(n93) );
    inv_0 U264 ( .x(n116), .a(n206) );
    nor2i_3 U265 ( .x(n81), .a(n83), .b(n82) );
    inv_0 U266 ( .x(n83), .a(B[10]) );
    nand2i_4 U267 ( .x(n222), .a(A[21]), .b(B[21]) );
    nand2i_2 U268 ( .x(n98), .a(A[16]), .b(B[16]) );
    nand2i_2 U269 ( .x(n227), .a(A[13]), .b(B[13]) );
    nor2i_1 U27 ( .x(n168), .a(n261), .b(n299) );
    nand2i_3 U271 ( .x(n284), .a(A[12]), .b(B[12]) );
    nand2i_2 U272 ( .x(n225), .a(B[12]), .b(A[12]) );
    nand2_2 U273 ( .x(DIFF[1]), .a(n86), .b(n87) );
    aoi21_3 U274 ( .x(n88), .a(n89), .b(n90), .c(n71) );
    nor2_5 U275 ( .x(n102), .a(n103), .b(n104) );
    nor2i_5 U276 ( .x(n119), .a(B[11]), .b(A[11]) );
    aoi21_3 U277 ( .x(n123), .a(n124), .b(n332), .c(n126) );
    nor2_5 U278 ( .x(n135), .a(n136), .b(n137) );
    and3i_3 U279 ( .x(n171), .a(n64), .b(n172), .c(n173) );
    inv_0 U28 ( .x(n169), .a(n258) );
    exor2_3 U280 ( .x(DIFF[26]), .a(n196), .b(n135) );
    exor2_3 U281 ( .x(DIFF[25]), .a(n197), .b(n138) );
    exnor2_3 U282 ( .x(DIFF[21]), .a(n123), .b(n144) );
    exnor2_5 U283 ( .x(DIFF[15]), .a(n88), .b(n154) );
    aoai211_4 U285 ( .x(n238), .a(n239), .b(n240), .c(n241), .d(n242) );
    aoai211_4 U286 ( .x(n263), .a(n264), .b(B[11]), .c(n243), .d(n265) );
    exnor2_5 U287 ( .x(DIFF[30]), .a(n171), .b(n268) );
    exor2_3 U288 ( .x(DIFF[11]), .a(n276), .b(n277) );
    aoi21_3 U289 ( .x(n292), .a(n293), .b(n263), .c(n291) );
    nand2_2 U29 ( .x(n258), .a(n259), .b(n260) );
    nand2i_4 U290 ( .x(n304), .a(B[4]), .b(A[4]) );
    oai211_4 U291 ( .x(n310), .a(n311), .b(n210), .c(n307), .d(n306) );
    oai21_4 U292 ( .x(n184), .a(n185), .b(n109), .c(n240) );
    nand2i_4 U293 ( .x(n314), .a(A[27]), .b(B[27]) );
    inv_5 U294 ( .x(n264), .a(n238) );
    aoai211_4 U295 ( .x(n317), .a(n318), .b(n315), .c(n249), .d(n314) );
    inv_5 U296 ( .x(n323), .a(n202) );
    oai21_4 U297 ( .x(n201), .a(n164), .b(n323), .c(n225) );
    inv_5 U298 ( .x(n325), .a(n203) );
    oai21_4 U299 ( .x(n276), .a(n166), .b(n325), .c(n242) );
    nand2i_2 U30 ( .x(n244), .a(A[22]), .b(B[22]) );
    aoai211_4 U300 ( .x(n270), .a(B[23]), .b(n215), .c(n272), .d(n220) );
    exnor2_3 U301 ( .x(n268), .a(n57), .b(B[30]) );
    nand2i_5 U302 ( .x(n202), .a(n263), .b(n322) );
    ao21_4 U303 ( .x(n197), .a(n217), .b(n270), .c(n316) );
    ao21_4 U304 ( .x(n196), .a(n50), .b(n270), .c(n255) );
    inv_6 U305 ( .x(n185), .a(n310) );
    nand2i_5 U306 ( .x(n322), .a(n229), .b(n310) );
    or3i_5 U307 ( .x(n330), .a(n334), .b(n285), .c(n279) );
    nand2i_6 U308 ( .x(n282), .a(A[2]), .b(B[2]) );
    nor2i_5 U309 ( .x(n180), .a(n178), .b(n181) );
    nand2i_0 U31 ( .x(n142), .a(B[22]), .b(A[22]) );
    nand2i_4 U310 ( .x(n265), .a(B[11]), .b(n238) );
    nand2i_6 U311 ( .x(n224), .a(A[15]), .b(B[15]) );
    nand2i_8 U312 ( .x(n246), .a(A[19]), .b(B[19]) );
    nand2i_6 U313 ( .x(n210), .a(n211), .b(n54) );
    nand2i_5 U314 ( .x(n306), .a(n102), .b(n54) );
    nand2_6 U315 ( .x(n223), .a(n224), .b(n90) );
    nand2i_6 U316 ( .x(n175), .a(n170), .b(n53) );
    exnor2_1 U317 ( .x(DIFF[10]), .a(n203), .b(n331) );
    inv_2 U318 ( .x(n331), .a(n165) );
    oai21_2 U319 ( .x(n203), .a(n312), .b(n107), .c(n239) );
    oai21_1 U32 ( .x(n128), .a(n146), .b(n221), .c(n145) );
    or3i_3 U320 ( .x(n332), .a(n300), .b(n296), .c(n167) );
    or3i_3 U321 ( .x(n300), .a(n97), .b(n245), .c(n256) );
    or3i_1 U322 ( .x(n125), .a(n300), .b(n296), .c(n167) );
    and4_5 U323 ( .x(n334), .a(n335), .b(n234), .c(n52), .d(n235) );
    buf_1 U324 ( .x(n333), .a(n287) );
    aoi21_3 U325 ( .x(n287), .a(n334), .b(n336), .c(n290) );
    inv_2 U326 ( .x(n335), .a(n233) );
    inv_6 U327 ( .x(n234), .a(n229) );
    inv_4 U328 ( .x(n235), .a(n210) );
    and2_5 U329 ( .x(n52), .a(n226), .b(n227) );
    inv_0 U33 ( .x(n146), .a(n222) );
    nand2_0 U330 ( .x(n233), .a(n284), .b(n281) );
    and2_6 U331 ( .x(n53), .a(n51), .b(n244) );
    and2_5 U332 ( .x(n51), .a(n124), .b(n222) );
    aoai211_2 U333 ( .x(n266), .a(B[30]), .b(n319), .c(n254), .d(n320) );
    inv_5 U334 ( .x(n319), .a(n253) );
    oai211_1 U335 ( .x(n336), .a(n308), .b(n208), .c(n133), .d(n301) );
    oai211_1 U336 ( .x(n289), .a(n308), .b(n208), .c(n133), .d(n301) );
    nand2i_0 U337 ( .x(n237), .a(B[13]), .b(A[13]) );
    nand2i_0 U34 ( .x(n221), .a(B[20]), .b(A[20]) );
    inv_0 U35 ( .x(n148), .a(n124) );
    nand2i_2 U36 ( .x(n124), .a(A[20]), .b(B[20]) );
    nand2i_2 U38 ( .x(n309), .a(n134), .b(n289) );
    nand3_1 U39 ( .x(n181), .a(n281), .b(n282), .c(n283) );
    inv_4 U4 ( .x(n226), .a(n223) );
    nand2i_5 U40 ( .x(n178), .a(A[0]), .b(B[0]) );
    nand2_2 U41 ( .x(n256), .a(n98), .b(n257) );
    inv_2 U42 ( .x(n299), .a(n262) );
    inv_2 U43 ( .x(n177), .a(A[17]) );
    nand2i_2 U44 ( .x(n262), .a(n177), .b(n99) );
    oai21_1 U45 ( .x(n121), .a(n113), .b(n85), .c(n112) );
    inv_2 U46 ( .x(n75), .a(B[6]) );
    nand2i_0 U47 ( .x(n112), .a(B[7]), .b(A[7]) );
    inv_2 U48 ( .x(n103), .a(n304) );
    inv_4 U49 ( .x(n120), .a(n306) );
    oai211_1 U51 ( .x(n249), .a(n218), .b(n220), .c(n250), .d(n251) );
    nand2_2 U52 ( .x(n318), .a(n329), .b(n328) );
    nand2i_2 U53 ( .x(n183), .a(n213), .b(n130) );
    inv_2 U54 ( .x(n213), .a(B[28]) );
    nand2i_0 U55 ( .x(n130), .a(B[27]), .b(A[27]) );
    nand2i_2 U56 ( .x(n182), .a(A[28]), .b(n130) );
    ao221_4 U57 ( .x(n253), .a(n70), .b(n69), .c(n68), .d(n66), .e(n64) );
    inv_2 U58 ( .x(n279), .a(n178) );
    nand2i_2 U59 ( .x(n208), .a(B[1]), .b(A[1]) );
    nand2_2 U6 ( .x(n241), .a(n84), .b(n230) );
    inv_2 U60 ( .x(n302), .a(n208) );
    nand2_2 U61 ( .x(n87), .a(n302), .b(n178) );
    nor2i_1 U62 ( .x(n280), .a(B[1]), .b(n178) );
    inv_2 U63 ( .x(n209), .a(B[1]) );
    exnor2_1 U64 ( .x(n278), .a(n279), .b(n209) );
    mux2i_1 U65 ( .x(n86), .d0(n278), .sl(A[1]), .d1(n280) );
    nand2i_2 U66 ( .x(n230), .a(A[9]), .b(B[9]) );
    nand2i_0 U67 ( .x(n155), .a(B[15]), .b(A[15]) );
    nand2i_2 U68 ( .x(n248), .a(B[16]), .b(A[16]) );
    nand2_0 U69 ( .x(n200), .a(n248), .b(n98) );
    nand2i_2 U7 ( .x(n283), .a(A[1]), .b(B[1]) );
    inv_2 U70 ( .x(n99), .a(n248) );
    nand2i_0 U71 ( .x(n145), .a(B[21]), .b(A[21]) );
    exnor2_1 U72 ( .x(n273), .a(A[23]), .b(B[23]) );
    inv_2 U73 ( .x(n77), .a(n294) );
    inv_2 U74 ( .x(n297), .a(n142) );
    ao211_2 U75 ( .x(n55), .a(n298), .b(n258), .c(n174), .d(n176) );
    nand2i_2 U76 ( .x(n220), .a(B[23]), .b(A[23]) );
    nand2i_2 U77 ( .x(n251), .a(B[26]), .b(A[26]) );
    nand2i_2 U78 ( .x(n219), .a(A[26]), .b(B[26]) );
    oai21_1 U79 ( .x(n255), .a(n140), .b(n214), .c(n139) );
    nand2_2 U8 ( .x(n250), .a(n255), .b(n219) );
    nand2i_0 U80 ( .x(n214), .a(B[24]), .b(A[24]) );
    nand2i_2 U81 ( .x(n139), .a(B[25]), .b(A[25]) );
    nand2i_2 U82 ( .x(n216), .a(A[25]), .b(B[25]) );
    inv_2 U83 ( .x(n134), .a(n281) );
    nor2i_1 U84 ( .x(n132), .a(n133), .b(n134) );
    nand2i_2 U85 ( .x(n301), .a(B[2]), .b(A[2]) );
    inv_2 U86 ( .x(n308), .a(n282) );
    oai21_1 U87 ( .x(n191), .a(n308), .b(n321), .c(n301) );
    inv_2 U88 ( .x(n321), .a(n198) );
    nand2_2 U89 ( .x(n199), .a(n282), .b(n301) );
    nor3i_1 U9 ( .x(n176), .a(n99), .b(n177), .c(n175) );
    inv_2 U90 ( .x(n207), .a(A[1]) );
    aoai211_1 U91 ( .x(n198), .a(B[1]), .b(n207), .c(n279), .d(n208) );
    exnor2_1 U92 ( .x(DIFF[2]), .a(n198), .b(n199) );
    exor2_1 U93 ( .x(DIFF[6]), .a(n187), .b(n114) );
    ao21_1 U94 ( .x(n187), .a(n188), .b(n205), .c(n104) );
    nor2_1 U95 ( .x(n114), .a(n115), .b(n116) );
    inv_2 U96 ( .x(n115), .a(n85) );
    exor2_1 U97 ( .x(DIFF[12]), .a(n202), .b(n162) );
    nor2_1 U98 ( .x(n162), .a(n163), .b(n164) );
    inv_2 U99 ( .x(n163), .a(n225) );
endmodule


module EX_DW01_sub_32_1_test_1 ( A, B, CI, DIFF, CO );
input  [31:0] A;
input  [31:0] B;
output [31:0] DIFF;
input  CI;
output CO;
    wire n102, n258, n282, n254, n230, n151, n154, n152, n52, n166, n82, n88, 
        n87, n85, n86, n118, n174, n117, n179, n116, n159, n269, n160, n121, 
        n187, n188, n189, n272, n96, n182, n91, n95, n93, n94, n119, n120, 
        n262, n266, n205, n267, n260, n268, n171, n207, n202, n130, n178, n100, 
        n69, n206, n75, n215, n79, n246, n73, n74, n76, n158, n104, n155, n270, 
        n105, n106, n72, n216, n71, n128, n263, n150, n67, n68, n168, n265, 
        n238, n170, n101, n103, n279, n271, n231, n176, n255, n55, n157, n199, 
        n259, n141, n186, n126, n275, n125, n224, n252, n251, n277, n139, n137, 
        n140, n185, n163, n235, n98, n97, n122, n99, n222, n219, n220, n223, 
        n90, n221, n83, n243, n208, n60, n209, n210, n211, n248, n214, n80, 
        n81, n53, n247, n78, n77, n162, n132, n108, n114, n135, n146, n56, 
        n107, n111, n218, n236, n237, n89, n92, n165, n142, n138, n144, n167, 
        n253, n164, n233, n234, n84, n191, n153, n192, n232, n50, n195, n281, 
        n177, n280, n51, n264, n217, n183, n181, n175, n148, n273, n201, n261, 
        n180, n54, n57, n109, n58, n149, n59, n225, n241, n70, n193, n61, n62, 
        n172, n110, n115, n64, n65, n66, n257, n127, n196, n197, n198, n203, 
        n204, n226, n227, n228, n256, n274, n242, n212, n184, n173, n249, n250, 
        n156, n213, n240, n200, n283, n284, n63, n245, n244, n169, n239, n113, 
        n124, n143, n194, n161, n129, n134, n276, n133, n131, n147, n136, n112, 
        n278, n190, n123, n145, n229;
    inv_4 U10 ( .x(n102), .a(n258) );
    nand2i_2 U100 ( .x(n282), .a(n254), .b(n230) );
    and3i_1 U101 ( .x(n151), .a(n154), .b(n152), .c(n52) );
    nand3i_1 U102 ( .x(n166), .a(n151), .b(n258), .c(n282) );
    inv_2 U103 ( .x(n82), .a(n88) );
    inv_0 U104 ( .x(n87), .a(A[22]) );
    aoai211_1 U105 ( .x(DIFF[22]), .a(n85), .b(n86), .c(n87), .d(n88) );
    inv_2 U106 ( .x(n118), .a(n174) );
    inv_2 U107 ( .x(n117), .a(n179) );
    nor2_1 U108 ( .x(n116), .a(n117), .b(n118) );
    ao21_1 U109 ( .x(n159), .a(n269), .b(n160), .c(n121) );
    nand2_2 U11 ( .x(n187), .a(n188), .b(n189) );
    nand2i_2 U110 ( .x(n269), .a(A[4]), .b(B[4]) );
    inv_2 U111 ( .x(n272), .a(n159) );
    nand2i_0 U112 ( .x(n96), .a(n182), .b(n91) );
    inv_0 U113 ( .x(n95), .a(A[19]) );
    aoai211_1 U114 ( .x(DIFF[19]), .a(n93), .b(n94), .c(n95), .d(n96) );
    nor2_1 U115 ( .x(n119), .a(n120), .b(n121) );
    inv_2 U116 ( .x(n121), .a(n262) );
    nand2i_0 U117 ( .x(n262), .a(B[4]), .b(A[4]) );
    inv_2 U118 ( .x(n266), .a(n205) );
    aoai211_1 U119 ( .x(n267), .a(n260), .b(n268), .c(n171), .d(n207) );
    nand2i_2 U12 ( .x(n202), .a(n130), .b(n178) );
    nand4i_1 U120 ( .x(n205), .a(n100), .b(n69), .c(n206), .d(n207) );
    nand2i_3 U121 ( .x(n75), .a(n215), .b(n91) );
    nand2i_2 U122 ( .x(n79), .a(n246), .b(n91) );
    oai211_1 U123 ( .x(DIFF[28]), .a(n73), .b(n74), .c(n75), .d(n76) );
    exor2_1 U124 ( .x(DIFF[8]), .a(n158), .b(n104) );
    nand2_2 U125 ( .x(n158), .a(n155), .b(n270) );
    nor2_0 U126 ( .x(n104), .a(n105), .b(n106) );
    nand2i_3 U127 ( .x(n72), .a(n216), .b(A[29]) );
    nand2_1 U128 ( .x(DIFF[29]), .a(n71), .b(n72) );
    inv_2 U129 ( .x(n128), .a(A[30]) );
    nand2i_2 U13 ( .x(n263), .a(n150), .b(n260) );
    oai21_1 U130 ( .x(DIFF[1]), .a(A[1]), .b(n67), .c(n68) );
    exnor2_1 U131 ( .x(n67), .a(n69), .b(n168) );
    inv_2 U132 ( .x(n168), .a(B[1]) );
    mux2i_1 U133 ( .x(n68), .d0(n260), .sl(n265), .d1(n238) );
    inv_2 U134 ( .x(n260), .a(n170) );
    inv_2 U135 ( .x(n265), .a(n69) );
    nor2_0 U136 ( .x(n101), .a(n102), .b(n103) );
    inv_2 U137 ( .x(n279), .a(n271) );
    inv_2 U138 ( .x(n105), .a(n231) );
    inv_2 U139 ( .x(n152), .a(n176) );
    nor2i_0 U14 ( .x(n150), .a(B[2]), .b(A[2]) );
    nand2_2 U140 ( .x(n255), .a(n55), .b(B[8]) );
    inv_5 U141 ( .x(n106), .a(n255) );
    oai211_1 U142 ( .x(n157), .a(n106), .b(n155), .c(n231), .d(n271) );
    inv_2 U143 ( .x(n199), .a(n259) );
    inv_2 U144 ( .x(n141), .a(n186) );
    inv_2 U145 ( .x(n126), .a(n275) );
    inv_2 U146 ( .x(n125), .a(n224) );
    aoi21_1 U147 ( .x(n252), .a(n125), .b(n189), .c(n126) );
    nand2_2 U148 ( .x(n251), .a(n188), .b(n189) );
    oai21_1 U149 ( .x(n277), .a(n139), .b(n137), .c(n140) );
    nor3_0 U15 ( .x(n185), .a(A[22]), .b(A[20]), .c(A[21]) );
    aoai211_1 U150 ( .x(n163), .a(n186), .b(n277), .c(n251), .d(n252) );
    exor2_1 U151 ( .x(DIFF[16]), .a(n235), .b(n98) );
    inv_2 U152 ( .x(n93), .a(n97) );
    inv_0 U153 ( .x(n122), .a(A[17]) );
    nor2i_1 U154 ( .x(n99), .a(n122), .b(n93) );
    inv_0 U155 ( .x(n98), .a(A[16]) );
    nand4_1 U156 ( .x(n97), .a(n222), .b(n219), .c(n220), .d(n223) );
    aoi31_1 U157 ( .x(DIFF[17]), .a(n97), .b(n98), .c(n91), .d(n99) );
    nand4i_1 U158 ( .x(n90), .a(A[20]), .b(n219), .c(n220), .d(n221) );
    inv_2 U159 ( .x(n83), .a(A[23]) );
    nor2_1 U16 ( .x(n243), .a(A[25]), .b(A[24]) );
    nand4_2 U160 ( .x(n208), .a(n60), .b(n209), .c(n210), .d(n211) );
    nand2i_2 U161 ( .x(n248), .a(A[23]), .b(n214) );
    nand2_2 U162 ( .x(DIFF[25]), .a(n80), .b(n81) );
    oai21_1 U163 ( .x(n81), .a(n53), .b(n247), .c(A[25]) );
    inv_2 U164 ( .x(n78), .a(A[26]) );
    inv_2 U165 ( .x(n77), .a(n80) );
    oai21_1 U166 ( .x(DIFF[26]), .a(n77), .b(n78), .c(n79) );
    exor2_1 U167 ( .x(DIFF[2]), .a(n162), .b(n132) );
    exor2_1 U168 ( .x(DIFF[6]), .a(n108), .b(n114) );
    exnor2_1 U169 ( .x(DIFF[12]), .a(n135), .b(n146) );
    inv_4 U17 ( .x(n56), .a(A[9]) );
    exnor2_1 U170 ( .x(DIFF[7]), .a(n107), .b(n111) );
    exnor2_1 U171 ( .x(DIFF[27]), .a(n73), .b(n218) );
    inv_2 U172 ( .x(n73), .a(n79) );
    inv_0 U173 ( .x(n218), .a(A[27]) );
    exor2_1 U174 ( .x(DIFF[11]), .a(n236), .b(n237) );
    inv_1 U175 ( .x(n89), .a(n182) );
    aoi31_1 U176 ( .x(DIFF[20]), .a(n89), .b(n90), .c(n91), .d(n92) );
    exor2_1 U177 ( .x(DIFF[14]), .a(n165), .b(n142) );
    exnor2_1 U178 ( .x(DIFF[13]), .a(n138), .b(n144) );
    exnor2_1 U179 ( .x(DIFF[10]), .a(n166), .b(n167) );
    nor2_0 U18 ( .x(n253), .a(n106), .b(n103) );
    exor2_1 U180 ( .x(DIFF[5]), .a(n159), .b(n116) );
    exor2_1 U181 ( .x(DIFF[4]), .a(n160), .b(n119) );
    inv_2 U182 ( .x(n94), .a(A[18]) );
    exnor2_1 U183 ( .x(DIFF[18]), .a(n93), .b(n94) );
    exor2_1 U184 ( .x(DIFF[9]), .a(n157), .b(n101) );
    exnor2_1 U185 ( .x(DIFF[15]), .a(n163), .b(n164) );
    inv_2 U186 ( .x(n86), .a(A[21]) );
    exnor2_1 U187 ( .x(DIFF[21]), .a(n85), .b(n86) );
    exnor2_1 U188 ( .x(DIFF[24]), .a(n233), .b(n234) );
    inv_2 U189 ( .x(n233), .a(n84) );
    nand2_3 U19 ( .x(n191), .a(n153), .b(n192) );
    inv_2 U190 ( .x(n234), .a(A[24]) );
    inv_2 U191 ( .x(n232), .a(A[31]) );
    and2_6 U192 ( .x(n50), .a(n195), .b(n140) );
    nand2i_2 U193 ( .x(n281), .a(A[4]), .b(B[4]) );
    inv_2 U194 ( .x(n120), .a(n269) );
    inv_2 U195 ( .x(n177), .a(n280) );
    and2_1 U196 ( .x(n51), .a(n264), .b(n263) );
    inv_0 U197 ( .x(n74), .a(A[28]) );
    nand2_0 U198 ( .x(n76), .a(A[27]), .b(A[28]) );
    inv_2 U199 ( .x(n217), .a(A[29]) );
    nand2_2 U20 ( .x(n230), .a(n155), .b(n231) );
    nand2_8 U200 ( .x(n71), .a(n216), .b(n217) );
    inv_10 U201 ( .x(n216), .a(n75) );
    nor2_0 U202 ( .x(n183), .a(A[18]), .b(A[19]) );
    inv_2 U203 ( .x(n52), .a(n103) );
    inv_0 U204 ( .x(n103), .a(n153) );
    aoi21_5 U205 ( .x(n155), .a(n181), .b(n175), .c(n148) );
    inv_7 U206 ( .x(n273), .a(n201) );
    nand2i_0 U207 ( .x(n261), .a(B[7]), .b(A[7]) );
    nand2i_2 U208 ( .x(n175), .a(A[7]), .b(B[7]) );
    ao21_6 U209 ( .x(n180), .a(n181), .b(n175), .c(n148) );
    inv_2 U21 ( .x(n55), .a(A[8]) );
    inv_2 U210 ( .x(n53), .a(n91) );
    nand2_2 U211 ( .x(n186), .a(n54), .b(A[12]) );
    inv_0 U212 ( .x(n54), .a(B[12]) );
    nand2_4 U213 ( .x(n153), .a(n56), .b(B[9]) );
    inv_0 U214 ( .x(n57), .a(n109) );
    inv_2 U215 ( .x(n58), .a(n57) );
    nand2i_0 U216 ( .x(n174), .a(A[5]), .b(B[5]) );
    nand2i_4 U217 ( .x(n179), .a(B[5]), .b(A[5]) );
    oai211_4 U218 ( .x(n149), .a(n59), .b(A[5]), .c(n58), .d(n175) );
    inv_4 U219 ( .x(n59), .a(B[5]) );
    nand2_0 U22 ( .x(n254), .a(n52), .b(n255) );
    aoai211_3 U220 ( .x(n211), .a(n50), .b(n225), .c(n241), .d(n259) );
    nand2i_2 U221 ( .x(n69), .a(A[0]), .b(B[0]) );
    nand2i_0 U222 ( .x(n70), .a(B[0]), .b(A[0]) );
    inv_2 U223 ( .x(n193), .a(n61) );
    inv_0 U224 ( .x(n62), .a(B[10]) );
    nand2i_4 U225 ( .x(n172), .a(B[3]), .b(A[3]) );
    aoi21_1 U226 ( .x(n107), .a(n108), .b(n58), .c(n110) );
    inv_2 U227 ( .x(n115), .a(n58) );
    nand2i_3 U228 ( .x(n231), .a(B[8]), .b(A[8]) );
    inv_0 U229 ( .x(n64), .a(B[10]) );
    nand2i_0 U23 ( .x(n154), .a(n106), .b(n160) );
    inv_0 U230 ( .x(n65), .a(A[10]) );
    nand2_0 U231 ( .x(n109), .a(n66), .b(B[6]) );
    nand2i_3 U232 ( .x(n189), .a(A[14]), .b(B[14]) );
    nand2i_2 U233 ( .x(n188), .a(A[13]), .b(B[13]) );
    nand2i_4 U234 ( .x(n140), .a(A[12]), .b(B[12]) );
    nand2i_0 U235 ( .x(n257), .a(B[6]), .b(A[6]) );
    oai21_4 U236 ( .x(DIFF[23]), .a(n82), .b(n83), .c(n84) );
    nor2i_5 U237 ( .x(n127), .a(n128), .b(n71) );
    nor3i_5 U238 ( .x(n148), .a(A[4]), .b(B[4]), .c(n149) );
    nand2_5 U239 ( .x(n196), .a(n197), .b(n198) );
    inv_0 U24 ( .x(n264), .a(n171) );
    nand2i_4 U240 ( .x(n201), .a(n202), .b(n203) );
    nand2i_4 U241 ( .x(n204), .a(n149), .b(n203) );
    oai211_3 U242 ( .x(n225), .a(n191), .b(n226), .c(n227), .d(n228) );
    exnor2_5 U243 ( .x(DIFF[31]), .a(n127), .b(n232) );
    exnor2_3 U244 ( .x(DIFF[30]), .a(A[30]), .b(n71) );
    nand4_1 U246 ( .x(n235), .a(n211), .b(n256), .c(n220), .d(n219) );
    inv_5 U247 ( .x(n198), .a(n191) );
    or3i_5 U248 ( .x(n219), .a(n273), .b(n51), .c(n177) );
    or3i_5 U249 ( .x(n220), .a(n274), .b(n177), .c(n205) );
    nand2i_4 U250 ( .x(n242), .a(B[15]), .b(A[15]) );
    nand2_5 U251 ( .x(n256), .a(n203), .b(n180) );
    nand2i_4 U252 ( .x(n80), .a(n212), .b(n91) );
    nand2i_4 U253 ( .x(n88), .a(n184), .b(n91) );
    nand2i_4 U254 ( .x(n84), .a(n248), .b(n91) );
    nand2_2 U255 ( .x(n164), .a(n242), .b(n259) );
    inv_5 U256 ( .x(n274), .a(n204) );
    nand3_3 U257 ( .x(n209), .a(n274), .b(n281), .c(n266) );
    inv_12 U258 ( .x(n91), .a(n208) );
    nand2_8 U259 ( .x(n160), .a(n205), .b(n267) );
    nand2_2 U26 ( .x(n171), .a(n172), .b(n173) );
    nand2i_5 U260 ( .x(n259), .a(A[15]), .b(B[15]) );
    nor3i_5 U261 ( .x(n221), .a(n89), .b(n249), .c(n250) );
    nand3i_5 U262 ( .x(n271), .a(n106), .b(n160), .c(n152) );
    inv_6 U263 ( .x(n203), .a(n156) );
    nand2i_6 U264 ( .x(n206), .a(A[2]), .b(B[2]) );
    nand2i_4 U265 ( .x(n213), .a(A[23]), .b(n243) );
    oai21_5 U266 ( .x(n226), .a(n102), .b(n105), .c(n240) );
    nand3i_5 U267 ( .x(n156), .a(n199), .b(n50), .c(n200) );
    nand2i_5 U268 ( .x(n192), .a(A[11]), .b(B[11]) );
    and2_2 U269 ( .x(n283), .a(n284), .b(A[2]) );
    nand2i_0 U27 ( .x(n268), .a(A[2]), .b(B[2]) );
    inv_2 U270 ( .x(n173), .a(n283) );
    inv_2 U271 ( .x(n284), .a(B[2]) );
    inv_4 U272 ( .x(n240), .a(n63) );
    nor2_3 U273 ( .x(n197), .a(n106), .b(n63) );
    nor2i_3 U274 ( .x(n63), .a(n65), .b(n64) );
    nand2i_2 U28 ( .x(n207), .a(A[3]), .b(B[3]) );
    nor2i_0 U29 ( .x(n100), .a(B[1]), .b(A[1]) );
    nand2i_2 U30 ( .x(n212), .a(n213), .b(n214) );
    inv_2 U31 ( .x(n245), .a(n212) );
    nor2_0 U32 ( .x(n244), .a(A[26]), .b(A[27]) );
    nand3i_1 U33 ( .x(n215), .a(A[28]), .b(n244), .c(n245) );
    nand2i_0 U34 ( .x(n176), .a(n177), .b(n178) );
    nand2_2 U35 ( .x(n270), .a(n152), .b(n160) );
    nor2i_1 U36 ( .x(n238), .a(B[1]), .b(n169) );
    inv_2 U37 ( .x(n178), .a(n149) );
    nor2_1 U38 ( .x(n239), .a(n110), .b(n113) );
    oai21_3 U39 ( .x(n181), .a(n149), .b(n179), .c(n239) );
    nor2_1 U4 ( .x(n124), .a(n125), .b(n126) );
    nor2_1 U40 ( .x(n223), .a(n250), .b(n249) );
    inv_5 U41 ( .x(n250), .a(n211) );
    nor2_0 U42 ( .x(n222), .a(A[16]), .b(A[17]) );
    inv_2 U43 ( .x(n249), .a(n256) );
    nand2i_2 U44 ( .x(n280), .a(A[4]), .b(B[4]) );
    oai221_1 U45 ( .x(n241), .a(n143), .b(n124), .c(n186), .d(n187), .e(n242)
         );
    inv_2 U46 ( .x(n195), .a(n187) );
    or3i_3 U47 ( .x(n210), .a(n273), .b(n120), .c(n51) );
    inv_2 U48 ( .x(n200), .a(n196) );
    or2_2 U49 ( .x(n60), .a(n155), .b(n156) );
    nand2i_2 U5 ( .x(n228), .a(n194), .b(n61) );
    nand3i_0 U50 ( .x(n247), .a(A[23]), .b(n234), .c(n214) );
    nand2i_2 U51 ( .x(n184), .a(n182), .b(n185) );
    nand2i_0 U52 ( .x(n246), .a(A[26]), .b(n245) );
    inv_2 U53 ( .x(n214), .a(n184) );
    exor2_1 U54 ( .x(DIFF[3]), .a(n161), .b(n129) );
    oai21_1 U55 ( .x(n161), .a(n134), .b(n276), .c(n133) );
    nor2_1 U56 ( .x(n129), .a(n130), .b(n131) );
    inv_2 U57 ( .x(n130), .a(n207) );
    inv_0 U58 ( .x(n131), .a(n172) );
    inv_2 U59 ( .x(n134), .a(n206) );
    inv_2 U6 ( .x(n194), .a(A[11]) );
    nand2i_0 U60 ( .x(n133), .a(B[2]), .b(A[2]) );
    nor2i_1 U61 ( .x(n132), .a(n133), .b(n134) );
    aoai211_1 U62 ( .x(n162), .a(B[1]), .b(n169), .c(n265), .d(n170) );
    inv_2 U63 ( .x(n169), .a(A[1]) );
    nand2i_2 U64 ( .x(n170), .a(B[1]), .b(A[1]) );
    inv_2 U65 ( .x(n276), .a(n162) );
    nor2_1 U66 ( .x(n114), .a(n110), .b(n115) );
    nor2_1 U67 ( .x(n146), .a(n141), .b(n147) );
    nand4_1 U68 ( .x(n136), .a(n200), .b(n178), .c(n280), .d(n160) );
    nor2i_1 U69 ( .x(n135), .a(n136), .b(n137) );
    nor2i_0 U7 ( .x(n61), .a(n62), .b(n65) );
    nor2_1 U70 ( .x(n111), .a(n112), .b(n113) );
    inv_2 U71 ( .x(n112), .a(n175) );
    inv_2 U72 ( .x(n113), .a(n261) );
    oai21_1 U73 ( .x(n108), .a(n118), .b(n272), .c(n179) );
    inv_0 U74 ( .x(n66), .a(A[6]) );
    inv_2 U75 ( .x(n110), .a(n257) );
    nand2_2 U76 ( .x(DIFF[0]), .a(n69), .b(n70) );
    exnor2_1 U77 ( .x(n237), .a(B[11]), .b(A[11]) );
    oai21_1 U79 ( .x(n278), .a(n279), .b(n230), .c(n253) );
    inv_0 U8 ( .x(n190), .a(B[11]) );
    nand2i_2 U80 ( .x(n258), .a(B[9]), .b(A[9]) );
    aoai211_1 U81 ( .x(n236), .a(n258), .b(n278), .c(n63), .d(n193) );
    or3i_1 U82 ( .x(n182), .a(n183), .b(A[16]), .c(A[17]) );
    nor2i_1 U83 ( .x(n92), .a(n123), .b(n85) );
    inv_0 U84 ( .x(n123), .a(A[20]) );
    inv_2 U85 ( .x(n85), .a(n90) );
    nor2_1 U86 ( .x(n142), .a(n143), .b(n126) );
    inv_2 U87 ( .x(n143), .a(n189) );
    nand2i_0 U88 ( .x(n275), .a(B[14]), .b(A[14]) );
    nand2i_0 U89 ( .x(n224), .a(B[13]), .b(A[13]) );
    oai21_1 U9 ( .x(n227), .a(n61), .b(A[11]), .c(n190) );
    aoai211_1 U90 ( .x(n165), .a(n186), .b(n277), .c(n145), .d(n224) );
    inv_2 U91 ( .x(n145), .a(n188) );
    nor2_1 U92 ( .x(n144), .a(n145), .b(n125) );
    inv_2 U93 ( .x(n147), .a(n140) );
    inv_2 U94 ( .x(n229), .a(n225) );
    oai21_1 U95 ( .x(n137), .a(n155), .b(n196), .c(n229) );
    inv_2 U96 ( .x(n139), .a(n136) );
    oaoi211_1 U97 ( .x(n138), .a(n139), .b(n137), .c(n140), .d(n141) );
    nand2_2 U99 ( .x(n167), .a(n240), .b(n193) );
endmodule


module EX_test_1_desync ( ALU_result, reg_out_B_EX, mem_write_EX, mem_read_EX, 
    mem_to_reg_EX, reg_write_EX, reset, IR_opcode_field, IR_function_field, 
    reg_out_A, reg_out_B, Imm, reg_dst, reg_write, mem_to_reg, mem_read, 
    mem_write, _byte, word, counter, test_si, test_so, test_se, sync_sel, 
    global_g1, global_g2, Ctrl__Regs_1__en1, Ctrl__Regs_1__en2 );
output [31:0] ALU_result;
output [31:0] reg_out_B_EX;
input  [5:0] IR_opcode_field;
input  [5:0] IR_function_field;
input  [31:0] reg_out_A;
input  [31:0] reg_out_B;
input  [31:0] Imm;
input  [1:0] counter;
input  reset, reg_dst, reg_write, mem_to_reg, mem_read, mem_write, test_si, 
    test_se, sync_sel, global_g1, global_g2, Ctrl__Regs_1__en1, 
    Ctrl__Regs_1__en2;
output mem_write_EX, mem_read_EX, mem_to_reg_EX, reg_write_EX, _byte, word, 
    test_so;
    wire ALU_result_reg_0__m2s, n4049, n4017, n4018, ALU_result_reg_10__m2s, 
        n4059, n4020, ALU_result_reg_11__m2s, n4060, n542, n4021, 
        ALU_result_reg_12__m2s, n4061, n4154, ALU_result_reg_13__m2s, n4062, 
        n543, n4022, ALU_result_reg_14__m2s, n4063, n4153, 
        ALU_result_reg_15__m2s, n4064, n4023, ALU_result_reg_16__m2s, n4065, 
        n4024, ALU_result_reg_17__m2s, n4066, n4025, ALU_result_reg_18__m2s, 
        n4067, n4152, ALU_result_reg_19__m2s, n4068, n4151, 
        ALU_result_reg_1__m2s, n4050, n4019, ALU_result_reg_20__m2s, n4069, 
        n4027, ALU_result_reg_21__m2s, n4070, n4028, ALU_result_reg_22__m2s, 
        n4071, n4029, ALU_result_reg_23__m2s, n4072, n4030, 
        ALU_result_reg_24__m2s, n4073, n4031, ALU_result_reg_25__m2s, n4074, 
        n4032, ALU_result_reg_26__m2s, n4075, n4033, ALU_result_reg_27__m2s, 
        n4076, n4034, ALU_result_reg_28__m2s, n4077, n4035, 
        ALU_result_reg_29__m2s, n4078, n4036, ALU_result_reg_2__m2s, n4051, 
        n4026, ALU_result_reg_30__m2s, n4079, n4038, ALU_result_reg_31__m2s, 
        _ALU_result_reg_31_net106451, n4039, ALU_result_reg_3__m2s, n4052, 
        n4037, ALU_result_reg_4__m2s, n4053, n4040, ALU_result_reg_5__m2s, 
        n4054, n4041, ALU_result_reg_6__m2s, n4055, n4042, 
        ALU_result_reg_7__m2s, n4056, n4043, ALU_result_reg_8__m2s, n4057, 
        n4044, ALU_result_reg_9__m2s, n4058, n4045, n3235, n1577, n1729, n665, 
        n1964, n1070, n1235, n734, n2635, N1754, ___cell__39620_net145150, 
        n2639, n1801, n809, N1655, n2631, n829, n634, n2638, 
        ___cell__39620_net145285, n2645, n1805, n1987, N1820, n1315, n2722, 
        n3236, n1147, n1136, n2644, n1055, n2557, n661, n869, n3648, n844, 
        n1804, N1953, ___cell__39620_net143845, ___cell__39620_net144360, n708, 
        n1236, N1986, n3821, n3460, n1623, n2602, n3820, n1233, 
        ___cell__39620_net143864, n1234, n1322, n1972, n2609, n3418, n4004, 
        n1565, n1807, n3234, n1625, n2806, n2608, n649, n650, n2574, n2604, 
        n1486, n690, n2605, n1063, n646, n2607, n3826, n2620, 
        ___cell__39620_net144707, ___cell__39620_net145617, n811, n606, n1228, 
        N1854, n946, n1230, N1821, n1229, n1077, n1795, N1954, n3239, 
        ___cell__39620_net144201, net152465, n1794, N1887, n2595, n3997, n1226, 
        N1755, ___cell__39620_net143710, n2594, N1722, 
        ___cell__39620_net145190, n1227, n2593, n1793, N1656, n1788, N1955, 
        n1214, N1822, n1213, n565, n1302, n1043, n3524, n4007, n1806, n1653, 
        n497, n676, n2546, N1756, n1212, n2549, n1785, N1657, n2545, n689, 
        n590, n2548, n1060, n1061, n645, n1531, n2566, 
        ___cell__39620_net144517, n2375, n2564, n3811, n2649, n2266, n1091, 
        n1427, n1428, n1429, n3812, n2562, n2584, n688, n3385, n3384, n3444, 
        n3443, n1650, n2001, n1539, n2560, n2475, n1687, n1648, n1690, n2561, 
        n1256, n2477, n3815, n1578, n3684, n3447, n2738, n3232, n3229, n3230, 
        n3813, n1249, n1220, n1221, n1222, n2492, n2572, n1484, n2139, n1483, 
        n2571, n2543, n1626, net149120, n1218, n1781, n530, n1216, n1217, 
        n1219, n2544, n1451, n670, n3228, n3226, n3227, n3782, n2480, n3781, 
        n2479, n3780, n2435, n1711, n2436, n1712, n1443, n1659, n1542, n1540, 
        n1538, n1661, n2474, n1715, n1713, n3225, n3223, n3224, n2476, n3784, 
        n4009, n2286, n507, n1546, n3407, n3408, n2478, n2373, n1194, 
        ___cell__39620_net144302, n1533, n675, n1619, n1519, n1618, 
        ___cell__39620_net144303, n1525, n1523, n1526, n3798, n2779, n3222, 
        n3220, n3221, n1093, n3799, n3797, n1714, n2306, n1150, n2518, n2433, 
        n2270, n2273, n904, n1590, n1522, n1700, n3779, n3778, n3281, n1939, 
        n1951, n3806, n915, n813, n3386, n2568, n1481, n540, n3810, 
        ___cell__39620_net144199, n1116, ___cell__39620_net147732, n2526, 
        n2193, n1482, n2525, n737, n3801, n3315, n855, n882, n825, n2432, 
        n1122, n3739, n536, n3738, n2629, n854, n1330, n2981, n3585, n3783, 
        n3425, n3424, n1559, n1728, n1442, n1444, n1582, n1545, n3762, n3343, 
        n1160, n1568, n1543, n1612, n2677, n1207, n1208, n2506, n1775, n2502, 
        n3280, n2505, ___cell__39620_net147791, n810, n3726, n4125, n1290, 
        n1198, n2423, n2363, n1742, n2837, N310, n571, n3435, n2361, n1186, 
        n2197, n2356, n621, n3757, n2352, n1473, n2353, n3275, n3272, n3273, 
        n2354, n2355, n2357, ___cell__39620_net145524, 
        ___cell__39620_net145444, n2365, n2366, n1647, n1646, n2367, n2364, 
        n2368, n2369, n2370, n1173, n2347, n2345, n2348, n2349, n1182, n2168, 
        n2165, n1743, N1635, n1167, N1833, n3271, n3264, n3265, n3268, n1168, 
        N1999, n1169, n1172, N1966, ___cell__39620_net145508, n1745, N1933, 
        n1171, n3662, n1164, n1165, n1166, n2346, N1701, n1163, n1746, N1800, 
        n2351, n1744, N1866, n2350, n3263, n3261, n3262, n2836, n692, n1733, 
        n917, n2838, n2835, n3705, n1589, n2834, n2360, n1588, n1639, n2825, 
        n502, n2826, n1267, n2827, n2829, n1496, n2828, n1284, n2824, n1064, 
        n815, n2823, n3260, n1518, n3258, n3259, n1436, n1620, n2822, n3760, 
        n2814, N1733, n1271, n1270, n1838, N1634, n2816, n2815, n1839, N1932, 
        n2820, n3999, n1841, N1965, n2819, n1585, n608, n1840, N1832, n2818, 
        n4000, n1275, n1842, n3624, N1998, n1692, N313, n2142, n2141, n1566, 
        n2138, n2134, n2155, n3693, n2156, n2157, n1085, n2106, n1204, n1693, 
        N346, n1508, n644, n1694, N2002, n1696, N1936, n3697, n1699, N1969, 
        n2125, n1698, N1803, n2124, n1697, N1836, n2123, n2122, n2121, n3631, 
        n3559, ___cell__39620_net144331, n2120, N1704, n1111, n1695, N1638, 
        n2119, n2118, n3104, n3078, n3000, n3101, n3075, n2014, n3102, n3109, 
        n2022, n3110, n1389, n3115, n3118, n894, n3057, n3107, n1900, n977, 
        N352, n3961, n3291, n1906, N1975, n3096, n1905, N1842, n3095, n735, 
        n3094, n1095, n1988, n1197, n1397, n3093, n662, n594, n1381, n1386, 
        n1385, n1901, N2008, n1904, N1942, n712, n526, n504, n3020, n1384, 
        n1379, n1380, n1903, N1875, n3092, n3090, N1644, n1378, n1376, n1902, 
        N1743, n3091, n1383, n1675, N347, n2095, n3547, n3548, n3549, n2088, 
        n2089, n2090, n2094, n2091, n2092, n589, n2135, n2096, n2107, n2103, 
        n1681, N1970, n2077, n1680, N1804, n2076, n2074, n1318, n1993, n1992, 
        n2075, n2043, n1099, n1103, n1102, n1677, N2003, n1679, N1937, n1101, 
        n2071, n2068, n1678, N1639, n2072, n2501, ___cell__39620_net144406, 
        n3785, n3352, n658, n2500, n784, n2498, n2499, n1206, n2496, n1761, 
        N334, n2493, n2494, n2491, n2488, n2484, n2400, n539, n2489, n535, 
        n2490, n2481, n2485, n2486, n2487, n3794, n512, n3353, n3422, n1760, 
        n680, n2399, n3419, n3571, n2495, n1191, n681, n1573, n1769, N1857, 
        n2472, n1768, N1824, n2471, n2131, n1570, n1770, N1990, n2470, n2469, 
        n2473, n1196, n1201, n1763, N2023, n1162, n2384, n1764, N1659, n1765, 
        N1725, n3244, ___cell__39620_net143785, n3245, n1438, n3248, n3251, 
        n3253, n3254, n3255, n1110, n922, n1440, n3992, n3991, n1609, n2004, 
        n1937, n1638, n1627, n3290, n3214, N340, n1597, n1445, n3287, n1576, 
        n3288, n3289, n1453, n3131, n1574, n3129, n3130, n3134, n1908, N318, 
        n3133, n3126, n1403, n1907, n3127, n3128, n3132, n3041, n3147, n3117, 
        n3146, n3170, n900, n3137, n1909, N351, ___cell__39620_net144655, 
        n3135, n3139, n3141, n3142, n3143, n3710, n4008, n2024, n3116, n3113, 
        n1915, N1974, n3125, n1914, N1808, n3124, n3123, n1054, n1401, n1910, 
        N2007, n1913, N1941, n4010, n694, n891, n1400, n1396, n3119, N1643, 
        n1395, n1393, n1911, N1742, n3120, n1399, n3121, n2796, n2797, n513, 
        n2800, n702, n570, n2794, n1824, N327, n2184, n3354, n1558, n2788, 
        n2902, n2863, n1266, n1268, n3368, n3365, n1265, n2768, n2767, n1260, 
        n1828, ___cell__39620_net143660, n1827, N1751, N1718, n947, n1261, 
        N1883, n1833, N2016, n1999, n627, n3584, n3448, n659, n1264, n1829, 
        N1950, n1263, n2774, n3856, n1832, N1983, n2777, n1831, N1850, n2776, 
        n1830, N1817, n2775, n3701, n3196, n3046, n3001, n3039, n3040, n3042, 
        n3050, n3012, n3051, n3049, n3008, n1359, n3055, n3964, n3052, n3054, 
        n3047, n1884, N354, n1889, N1844, n3031, n2186, n2187, n1121, n3028, 
        N1811, n1339, n1890, N1977, n3030, n1354, n1885, N2010, n1888, N1944, 
        n1353, n1351, N1745, n3024, n1350, n3025, n3026, n3027, n2989, n1323, 
        n3937, n3936, n3935, n2230, n3079, n3973, n3086, n1892, N353, n3083, 
        n1374, n3067, n1364, n1898, N1976, n3066, n1897, N1810, n3065, n1367, 
        n1893, n2231, n2130, N2009, n1896, N1943, n1366, n1363, N1744, n1894, 
        N1645, n3062, ___cell__39620_net143872, n3061, n3063, 
        ___cell__39620_net144347, ___cell__39620_net144343, n1365, n2011, 
        n2054, n3163, n1917, n1686, n1684, N317, n3162, n3158, n3159, n1572, 
        n3155, n3173, n3174, n1415, n3167, n3168, n2023, n1414, n3164, n1916, 
        n3983, n1918, N350, n3153, n1409, n1922, N1807, n3154, n3150, n4141, 
        n1413, n1412, n1919, N2006, n1921, N1940, n1411, n3149, n1408, n1923, 
        N1973, n3152, n2176, n1584, n2177, n3148, N1642, n1407, n1405, n1920, 
        N1873, n3151, n3998, n2717, n1658, n3830, n2716, n3835, n2704, n1808, 
        N329, n2699, n3849, n2702, n2703, n2709, n2706, n2113, n2070, n583, 
        n1982, n2685, n1616, n3839, n2687, n1815, N1985, n2688, n1814, N1852, 
        n2678, n1240, n2679, n2680, n2681, n1810, N2018, n2684, n1812, N1885, 
        n2683, n944, n2114, n2115, n1246, n2682, n1813, N1952, n1245, n1243, 
        N1819, n1242, ___cell__39620_net144350, n2199, n2196, n2191, n2192, 
        n2194, n2195, n2198, n2188, n664, ___cell__39620_net144326, n2201, 
        n1703, N345, n2200, n2209, n2207, n2202, n2208, n1705, N1637, n2170, 
        n1706, N1703, n2169, n2166, n2167, n1129, n2164, n2069, n636, n1128, 
        n1704, N2001, n1708, N1935, n1127, n1709, N1968, n2175, n2174, N1802, 
        N1835, n1707, N1736, n2173, n2862, n743, n1297, n3706, n1561, n2855, 
        n887, n2856, n2857, n2861, n1498, n2860, n1497, n2858, n2859, n2871, 
        n2872, n842, n2869, n2867, n1844, N326, n1850, N1982, n2848, n3707, 
        ___cell__39620_net144317, n1361, n2845, n2846, n1291, n1848, N1882, 
        n2847, n1296, n2842, n1295, n2849, N1849, n1293, n1849, N1949, n1294, 
        n2243, n2241, n2234, n2211, n2235, n2212, n750, n1142, n940, n938, 
        n2240, n1468, n2239, n1467, n2237, n2238, n2242, n1717, N344, n2244, 
        n1718, N1636, n2221, n2219, n1140, n1725, n783, N2000, n1721, N1934, 
        n1139, n1138, n2222, n2223, n2224, n2225, n1722, N1801, n1723, N1834, 
        n1724, N1967, n3298, n1579, n928, n1720, n1719, N1867, N1735, n2909, 
        n1852, N325, n633, n632, n2905, n2908, n2906, n2907, n2904, n863, n862, 
        n2883, n1307, n2884, n2885, n2886, n1856, N1981, n2880, n865, n1304, 
        N1749, n1319, n2882, N1848, n1305, n1309, N2014, n2308, 
        ___cell__39620_net143784, n2311, n2309, n2310, n3789, n3478, n3745, 
        n1736, n821, n1161, n2328, n3749, n2327, n2331, n703, 
        ___cell__39620_net147270, n2329, n2330, n2332, n2317, n2318, n2319, 
        n2323, ___cell__39620_net143722, n2324, n2320, n2326, n2300, n3741, 
        ___cell__39620_net145472, ___cell__39620_net144555, n706, n710, n709, 
        n707, ___cell__39620_net145470, ___cell__39620_net145450, n798, 
        ___cell__39620_net145451, n3776, n1477, n2441, n2440, n1478, n2438, 
        n2439, n2442, n2443, n2444, n2445, n2402, n1190, n2454, n2453, n2457, 
        n1192, n2452, n615, N1662, n616, n2451, n2455, n2456, n2420, n588, 
        n663, n1757, N1726, n2419, n1188, N1759, n2418, n2421, n1755, N2024, 
        n2417, n1756, N1660, n2416, n3269, n1472, n2415, n2412, n2414, n3727, 
        n2413, n1758, N1958, n2427, n1759, N1825, n2057, n2059, n2027, n2052, 
        n3614, n3613, n2051, n2012, n2049, n1670, N1971, n2042, n2039, n1076, 
        n1669, N1838, n2041, n2040, n1666, N2004, n2038, n2035, N1640, n1075, 
        n1073, n1471, n1667, N1871, n2037, n2036, N1739, n1080, n1668, N1938, 
        n1079, n578, n2395, n2396, n2394, n2393, n3775, n1752, n3740, n2403, 
        n2405, n2407, n2408, n2409, n2401, n1185, n3724, n3723, n2404, n3765, 
        n2391, n816, n3720, n2372, n3767, n3766, n2390, n2185, n2389, n2377, 
        n2378, n2379, n2380, n2381, n2376, n1750, N2025, n2383, N1992, n1181, 
        n791, n782, n3719, n792, n794, ___cell__39620_net145428, n2288, n2289, 
        n1727, N1961, ___cell__39620_net144355, ___cell__39620_net143653, 
        n1726, N2027, n2293, n1153, n2294, n678, n1662, n1087, n1663, n701, 
        n2428, n1529, n2429, n3988, n1424, n3190, n3987, n3192, N1997, n1426, 
        n1517, n1425, n3207, n3209, n3206, n3205, n3180, 
        ___cell__39620_net144175, n3989, n1924, N308, n1437, n3219, n3216, 
        n3215, n1657, n3217, n3218, n941, n3212, n942, N341, n3611, n3610, 
        n2093, n2016, n1594, n1475, N316, n2013, n2007, n3623, n3622, n3620, 
        n3619, n1062, n1532, n2008, n2009, n2026, n2028, n2025, n720, n2021, 
        n2020, n2029, n3266, n1476, n2019, n1598, N349, n2033, n3172, n1615, 
        N1839, n1991, n1986, N1806, n1617, N1972, n1990, n1989, n1089, n713, 
        n927, n1058, n1599, N2005, n1613, N1939, n1057, n1056, n1053, n1984, 
        n1985, n1983, n1600, N1740, n1601, N1872, N1641, n1052, n1050, n498, 
        n3011, n3013, n3003, n3004, ___cell__39620_net143982, n2999, n3002, 
        n2899, n2996, n1876, N355, n3006, n2987, n1881, n2985, n1308, n1340, 
        n1882, N1978, n2986, n3761, n1635, n1344, n1877, N2011, n1880, N1945, 
        n1343, n1879, N1878, n1878, N1746, n2983, n2982, N1647, n1337, n1335, 
        n1868, N356, n2965, n1327, ___cell__39620_net147350, n718, n2970, 
        n1867, N323, n2963, n2962, n2961, n2964, n1871, N1946, n3938, n1873, 
        N2012, n3939, n2954, n2955, n2956, n2957, n2953, n3940, n2950, n3912, 
        n2920, n2918, n3910, n3911, n2921, n2922, n2923, n2924, n1863, N1947, 
        n1865, N2013, n2931, n2932, n2933, n2934, n2947, n1857, N324, n2946, 
        n1858, N357, n2752, n1817, N328, n2749, n2747, n2748, n2745, n1816, 
        n567, n2759, n757, n2803, n3854, n758, n2761, n4001, n2714, n2750, 
        n2760, n2724, n2723, n2725, n2726, n2727, n1821, N1884, n648, n2736, 
        n2732, n2733, n1253, n1818, N1653, n2735, n2734, n2731, n1822, n1823, 
        N1818, n2730, n2728, n1251, n2729, n1252, N2017, n1470, n4144, n2668, 
        n3553, n3552, n2671, n2624, n3825, n3824, n3823, n3822, n2660, n2661, 
        n2663, n2707, n2662, n2664, n2665, n3841, n3840, n2652, n1488, n1149, 
        n509, n2651, n1487, n2650, n3837, n747, n3836, n2628, n2655, n2654, 
        n2656, n2659, n1798, N330, n3842, n1797, n2658, n1313, n3401, n1691, 
        n901, n2657, n1800, N2019, n2642, n1803, N1886, n2641, n1802, N1721, 
        n2640, n1239, n2636, n2647, n2646, n2600, n1237, n3729, n1564, n3591, 
        n2627, n2626, n3816, n2625, n2618, n2623, n1791, N364, n2617, n2611, 
        n1790, N331, n3827, n2615, n2269, n1971, n1177, n2271, n2613, n3828, 
        n2614, n2612, n2610, n2621, n1232, n2598, n2596, n2592, n2597, n1796, 
        N1987, n2589, n1231, n1792, N2020, n2559, n3462, n2265, n2555, n1215, 
        N1988, n2558, n2556, n1784, N2021, n2554, n1787, N1888, n2553, n1786, 
        N1723, n2552, n2550, n3819, n3492, n3493, n2547, n2551, n1454, n1591, 
        n2587, n2586, n2579, n2580, n2573, n2532, n2567, n1223, n1224, n2585, 
        n2264, n2079, n2542, n2541, n2540, n2538, n2537, n1772, n1710, n1447, 
        n2536, n1210, n1211, n1595, n1534, n3805, n3804, n3807, n2529, n3809, 
        n3808, n2524, n2523, n1580, n2527, n2528, n2530, n3420, n2673, n2531, 
        n2263, n2302, n3423, n2534, n2763, n2533, n1520, n1184, n1209, N1956, 
        n1774, N2022, n2511, n1777, N1889, n3734, n3594, n2510, n1776, N1724, 
        n2509, n2507, n3803, n2515, n1779, N1989, n2517, n1780, 
        ___cell__39620_net144312, ___cell__39620_net144166, n805, n1005, N343, 
        n1004, ___cell__39620_net147731, n1006, n1151, n1152, n953, N309, N342, 
        ___cell__39620_net143326, n999, n1000, n1899, N319, n968, n1674, N314, 
        n959, n989, n2497, n1762, N367, n988, n1456, n2259, n1281, n2260, 
        n1036, n1825, N360, n1022, n1021, n2795, n2793, n2792, n1020, n1262, 
        n1883, N321, n971, n1891, N320, n1032, n1938, n965, n3160, n3161, 
        n1809, N362, n1019, n1018, n2705, n2700, n1017, n1247, n1244, n1702, 
        N312, n956, n954, n1126, n1845, N359, n1025, n3861, n1834, n1024, 
        n2868, n2865, n1023, n1716, N311, n1003, n1001, 
        ___cell__39620_net143287, n1002, n1853, N358, n3891, n976, n975, n2896, 
        n2903, n859, n1753, N335, n1007, n1754, N368, n1009, n1665, N315, n997, 
        n996, n1081, n993, n2387, n2382, n1416, n1417, n1418, 
        ___cell__39620_net144062, n991, n1748, N336, n1942, 
        ___cell__39620_net143655, n3211, n948, n3213, n1875, N322, n1030, n972, 
        n1026, n2937, n2940, n1027, n1421, N1864, n978, n807, n806, n1799, 
        N363, n981, n986, n1783, N365, n985, n1782, N332, n984, n1013, n1773, 
        n1420, N366, n733, n4117, n945, ___cell__6067_net21981, N3297, n4116, 
        n1530, n744, n1671, n4146, n3558, n3664, n1664, n830, N144, N70, n653, 
        n496, n3630, n499, n2890, n1602, n3532, n500, n1685, n541, n501, n549, 
        n548, n619, n503, n517, n4140, n803, n726, n725, n575, n576, n577, 
        n1676, ___cell__39620_net144330, n1524, n510, n1651, n890, n3758, 
        n1655, n671, n748, n3716, n3379, n729, n3374, n3335, n2133, n3699, 
        n834, n833, n514, n515, n3009, n3010, n637, n1333, n4005, 
        ___cell__39620_net144170, n518, n2988, n1837, n2268, n910, n519, n1238, 
        n2581, n3788, n943, n520, n1644, n889, n521, n858, n857, n3307, n761, 
        n3019, n880, n822, n3357, n523, n930, n3279, n3554, n3555, n524, n525, 
        n1643, n3366, n3369, n1629, n881, n2866, n3098, n1997, n3036, n3035, 
        n3918, n1767, N1890, n3339, n749, n527, n799, n2925, n2851, n2852, 
        n538, n1874, n1505, n1956, n1955, n1789, n1485, n1688, n1035, n3138, 
        n3136, n1034, n1402, n528, n529, n883, n3302, n531, n532, n1603, n533, 
        n1587, n3690, n1968, n1433, n1944, n2569, n2570, n2449, n1732, n2410, 
        n1682, n1683, n3694, n1349, n3717, n1042, n534, n935, 
        ___cell__39620_net144257, n537, n3433, n3602, n1183, n2385, n2388, 
        n3340, n1649, N1727, n556, N1892, N1760, n562, n1278, n1279, n3318, 
        n2313, N1761, N1728, n613, n3179, n2066, n902, n2067, n1630, n544, 
        n719, n3858, n2782, n2520, n2802, n1556, n2017, n2030, n2034, n868, 
        n2031, n2032, n2910, n2911, n546, n545, n888, n2160, n3350, n779, 
        ___cell__39620_net144029, n780, n774, n775, n3085, n764, n3112, n765, 
        n856, n848, n2232, n2233, n1134, n3692, n3668, n547, n584, n1175, n823, 
        n585, n1014, n1012, n1011, n893, n1569, n1551, n1960, n1958, n600, 
        n601, n4139, n1586, n836, n3391, n897, n899, n898, n1423, n3506, n2812, 
        n1049, n2938, n3895, n3894, n3893, n3892, n3069, n551, 
        ___cell__39620_net144781, n2344, n1047, n1738, n3355, n762, n3416, 
        n2939, n2941, n2942, n508, n3871, n3483, n2743, n2653, n2698, n552, 
        n3283, n1949, n1948, n3450, n797, n652, N1994, n2298, n1596, N371, 
        n3878, n3877, n2887, n2888, n2690, n769, n704, n839, n569, n3108, 
        n3114, n3111, n3484, n3644, n3652, n3470, n3471, n3472, n553, n3426, 
        n618, n3572, n2386, n3070, n2994, n2995, n2798, n2780, n2778, n554, 
        N370, n992, n1749, n840, ___cell__39620_net144345, n3199, n3200, n3321, 
        n3322, n3323, n1521, n3593, ___cell__39620_net145426, N1828, n555, 
        n557, n838, n937, n3362, n1583, n871, n3575, n1973, n1040, n1974, 
        n3608, n3325, n3603, n3311, n3607, n2213, n2214, n2159, n3276, n1730, 
        ___cell__39620_net144329, n923, n3754, n3687, n559, n1283, 
        ___cell__39620_net143997, n860, n3140, n3410, n625, n850, n2713, n1254, 
        n574, n3656, n2675, n3846, n960, n961, n962, n1541, n1448, n3919, 
        n1634, n1631, net151904, n3481, n3465, n969, n970, n558, n1995, n2715, 
        n3327, n763, n1739, n3573, n684, N1891, n3480, n3635, 
        ___cell__39620_net144322, n778, n560, n561, ___cell__39620_net144321, 
        n647, N1661, n2247, n3702, n563, n564, n2210, n3479, n3653, n1016, 
        n2616, n884, n623, n2753, n2754, n2755, n2756, n845, n2622, n846, 
        net150405, n2841, n875, n831, ___cell__39620_net143596, n788, n790, 
        n3945, n566, n3081, n660, n3074, n3080, n3077, n3171, n3358, n3313, 
        n1994, n1996, n1067, n568, ___cell__39620_net144173, n643, n3946, 
        n2927, n934, n987, n1105, n1555, n2228, n1391, n2226, n2126, n1066, 
        n3853, n3852, n2737, n2053, n1083, n2085, n3947, n2854, n892, n3928, 
        n1632, n572, n3691, n824, n1562, n1969, n3434, n2111, n3601, n3598, 
        n771, n573, n772, n607, n1980, n1979, n1978, n776, 
        ___cell__39620_net145078, ___cell__39620_net145077, n2003, n1065, 
        n3665, n2044, n3458, n3742, n3456, n579, n2056, n2424, N1991, n1189, 
        n1751, n1084, n878, n1331, n1976, n3446, n3445, n1654, n3414, n3545, 
        n3145, n3144, n2278, n2279, n2280, n925, n2303, n2603, n580, n581, 
        n3667, n3666, n3669, n1506, net151622, n609, n2691, n903, n3531, n2843, 
        n2840, n2844, n1847, n3486, n3654, n1450, n3862, n3165, n3166, n3169, 
        n3476, n3577, n751, n3576, n2064, n3518, n3198, n3449, 
        ___cell__39620_net143597, n657, N1894, n3475, n582, n1981, 
        ___cell__39620_net144328, n3914, n3303, n3795, n3770, n2708, net150620, 
        n3533, n3485, n979, n2751, n3579, n2179, n3678, n3915, n3033, n2336, 
        n2337, n2178, n886, n1100, n1094, n2073, n587, n895, n1656, n3746, 
        n2314, n2312, n1552, n1547, n1548, n1550, n1549, n3310, n3387, n913, 
        n851, n2181, n3324, n2619, n592, n3996, n591, n2583, n3916, n4127, 
        n593, n1332, n3954, n3953, n3952, n2512, n2513, n595, n3525, n2637, 
        n2590, n3523, n2218, n3181, n3187, n2813, n2811, n2343, n2217, n2215, 
        n3917, ___cell__39620_net144374, n3034, n1352, n3064, n597, n1660, 
        n598, n603, n4015, n2149, n2152, n2151, n2147, n2150, n3582, n604, 
        n3600, n3599, n738, n980, n982, n3539, n2216, n1419, n1345, n879, 
        n3921, n622, n1962, n656, n1961, n736, n936, n1086, n679, n610, n1605, 
        n1606, n2274, n3721, n2276, n3722, n2599, n3927, N1855, n3639, n2721, 
        n3855, n611, net156363, n612, n614, N1651, n2839, n617, net149627, 
        n3929, n3764, ___cell__39620_net143595, ___cell__39620_net145427, 
        ___cell__39620_net145418, ___cell__39620_net145425, n3516, n2514, 
        n2516, n620, n1452, n3294, n1037, n1038, n3477, n2227, n3451, n3233, 
        ___cell__39620_net145421, ___cell__39620_net145419, net150643, n3509, 
        n1607, n624, n3510, n3511, n3922, n3646, ___cell__39620_net147278, 
        n2807, n843, n1033, n3082, n3677, n3314, n739, n626, n3923, n629, n905, 
        n3122, n1398, n3029, n841, n2334, n3753, ___cell__39620_net143962, 
        n1334, n3924, n2783, n2116, ___cell__39620_net143658, n2112, n2801, 
        n2582, n2182, n2183, n1622, net149167, n801, n1614, n3925, n2784, n641, 
        n642, n1502, n2928, n2929, n2930, n1528, n777, n631, n651, n896, n789, 
        N1729, n1503, n1954, n1953, n1952, n3902, n654, n3903, n655, n516, 
        n766, n1701, n1633, n1324, n3421, n4006, n1689, n966, n967, n957, n958, 
        n3071, n1642, n3596, n828, n819, n1861, N1748, n3378, n826, 
        ___cell__39620_net144324, net151578, n2874, n752, n2850, n1159, n3382, 
        n4012, n3763, n666, n667, n1624, n3981, n668, n818, n1637, n669, n3007, 
        n3015, n773, n3638, n3948, n2299, N1861, n3191, N1831, N1964, n3628, 
        n3395, n3626, ___cell__39620_net143693, ___cell__39620_net143983, 
        n1866, n3818, n1072, n672, n673, n1289, n674, n677, 
        ___cell__39620_net144344, n3884, n3658, n3497, n3645, n2710, n3536, 
        n3535, n2006, ___cell__39620_net144605, n832, n3542, n3627, n921, 
        n3417, n2975, n1967, n3021, n3022, n3920, n685, n3306, n1557, n1039, 
        n686, n1133, n1120, n2790, n1493, n691, n3304, n3305, n3647, n3885, 
        n1940, n2002, n693, n3464, net149107, n696, n698, n697, n699, n727, 
        n3886, n700, n3612, n3499, N1663, n705, n808, n3904, n2719, n802, n800, 
        n3618, n3759, n3906, n2153, n2146, n2158, n2154, n3963, n3415, n711, 
        n908, n907, n714, n715, n635, n3905, n717, n3452, n723, n722, n721, 
        n724, n847, n3059, n3817, n728, n3317, n3504, n1178, n3328, n3329, 
        n3411, n3412, n963, n964, n1410, n3301, n1563, n926, n1636, n2891, 
        n2892, ___cell__39620_net144356, n804, n1257, n1560, n2810, n3336, 
        n812, n3334, n3337, n3338, n2236, n768, n3296, n874, n3467, n3312, 
        n2431, n3930, n2045, n2991, n740, n741, n742, n1449, n3860, n1608, 
        n2912, n640, n1501, ___cell__39620_net143954, n745, n2341, n2992, 
        n1998, n2000, n746, n3546, n3442, n2189, n912, n2190, n1130, n3604, 
        n3491, n2161, n1465, n2143, n2773, n1491, n628, N333, n3629, n2765, 
        n3859, n1672, n1673, n3528, n3551, n753, n754, n2277, n914, n1082, 
        n2281, n3375, n3592, n4134, n1459, n2283, n755, n756, n760, n759, 
        n2789, n2785, n2296, n1592, N338, N3304, n1250, n827, n767, n2669, 
        n2666, ___cell__39620_net143767, n770, N69, n3373, n793, n785, n787, 
        n786, N1762, ___cell__39620_net145429, n796, n3377, 
        ___cell__39620_net147296, n795, ___cell__39620_net145037, net151497, 
        ___cell__39620_net144309, ___cell__39620_net144200, net149616, n1535, 
        n3346, n3394, n3396, n3345, n3347, n3348, n814, n3319, n3320, n870, 
        n817, n2127, n2128, n1108, n1109, n3496, n2297, net149122, n820, n3881, 
        n4003, ___cell__39620_net144572, n2316, n2315, n3597, n3247, n3237, 
        n3238, n3241, n3256, n909, n1513, net149628, n3640, n885, n1179, n2148, 
        n1117, n1474, ___cell__39620_net143720, n2711, net151577, n1446, n1527, 
        n3274, n1628, n3461, n3257, n2588, n1104, n852, n1092, n1119, n3494, 
        n1088, n695, n1461, n1462, n861, n835, n3637, n506, n3495, n3588, 
        n3589, n1835, n1851, n1500, n2805, n3490, n4147, n1457, n2873, n4129, 
        ___cell__39620_net143694, ___cell__39620_net143836, n1460, n3488, 
        n3308, n3309, n3566, n3501, n3487, n3463, n3466, n3543, n3469, n3498, 
        n3390, n995, net150830, n2080, n1641, n2018, n4136, n1051, n1458, n924, 
        n2258, n998, n3578, n1604, n1158, n853, N369, n3473, n3563, n3404, 
        n3540, n2333, N337, n2083, n3383, n994, n2325, n2936, n2901, n2295, 
        n864, n2290, n2291, n866, n3786, n867, n3787, n3616, n2117, n2632, 
        n3838, n872, n2676, n2634, n2267, n877, n876, n919, n3556, n3969, n931, 
        n2606, n3737, n3792, n1404, n3053, n3056, n2799, n1269, n3014, n1347, 
        n2978, n1328, n2697, n3848, n2254, n1145, n2105, n1107, n2063, n1118, 
        n1652, n687, n1492, n2720, ___cell__39620_net144765, 
        ___cell__39620_net146131, n1504, n1507, n3023, n916, n3564, n3500, 
        n3405, n3474, n1571, n1510, n920, n1509, n3060, n1375, n1511, n682, 
        n1377, n3530, ___cell__39620_net143735, n1463, n1406, n1516, n1610, 
        n949, n950, n951, n952, n955, n683, n3202, n973, n983, n1015, n1028, 
        n1029, n1031, n1068, n1069, n1097, n1098, n1135, n1141, n1170, n1180, 
        N1959, n1187, n1193, n2565, n1195, N1957, n1202, n1199, n1200, N1984, 
        N2015, n1306, n1338, n1355, n1368, n1434, ___cell__39620_net144340, 
        n4137, n1621, N1870, N1893, n1740, n1741, N1658, n1778, N1823, N1856, 
        n1820, N1752, n4080, n4047, n1941, n4048, n4046, N3024, n1943, N3029, 
        n1945, n1946, n1947, N1392, N1402, N1407, n1957, n1963, n1965, n1966, 
        n1575, n1581, n1975, n1977, n1059, n2010, n2015, n2284, n2060, n2061, 
        n2058, n2062, n2078, n1090, n2097, n2100, n2101, n2102, n2098, n2110, 
        n1112, n2144, n2145, n2162, n2163, n2171, n522, n2180, n2205, n2203, 
        n2204, n2220, n1137, n2229, n2245, n2248, n2249, n2250, n2251, n2252, 
        n2246, n2253, n2255, n2256, n2257, n2301, n2342, n2358, n2359, n2362, 
        n2437, n2446, n2447, n2448, net149121, net156024, n2450, n1008, n2459, 
        n2463, n2464, n2466, n2467, n2468, n1203, n2504, n2503, n2519, n2262, 
        n2522, n2521, n2535, n2539, n2577, n2575, n2578, n1225, n2591, n2601, 
        n2643, n2648, n2674, n1241, n2686, n2695, n2696, n2692, n2701, n2712, 
        n2740, n2741, n2742, n2746, n1143, n2757, n2758, n2772, n2769, n2770, 
        n2771, n2791, n1836, n1277, n2817, n1273, n1276, n2821, n2830, n2831, 
        n2832, n2833, n2893, n2897, n2898, n2460, n1317, n2917, n2919, n2914, 
        n2943, n2944, n2945, n2958, n2966, n2967, n2968, n2969, n2971, n2972, 
        n2973, n2974, n2976, n2977, n2979, n2458, n1342, n2984, n3005, n3018, 
        n3016, n3017, n3045, n3037, n3044, n3048, n3076, n1372, n3084, n3105, 
        n3099, n3106, n3185, n3186, n3182, n1422, n3193, n3194, n3203, n3204, 
        n3208, n3210, n3595, n1514, n1495, n1499, n1490, n1494, n1479, n1469, 
        n3246, n3242, n1435, n1441, n1489, n1480, n1466, n1464, n3282, n3284, 
        n3292, n3293, n3316, n3326, n639, n638, n3351, n3332, n3333, n3344, 
        n3370, n3371, n3409, n3406, n1157, n3454, n3457, n3341, n3459, n3468, 
        n1045, n1156, n3482, n3537, n1123, n3538, n3541, n3544, n3278, n3557, 
        n3560, n3561, n3562, n3489, n3570, n3574, n3605, n3389, n3615, n3657, 
        n3682, n3683, n2065, n3695, n3696, n3681, n3703, n3704, n3176, n3436, 
        n3689, n3711, n2371, n3712, n3802, n3713, n3714, n3715, n3430, n2282, 
        n3718, n3367, n2285, n2275, n3625, n3392, n3750, n3751, n3752, n3755, 
        n1176, n2338, n3769, n2430, n3773, n3777, n3796, n3800, n2508, n3814, 
        n3636, n2670, n3829, n2667, n3843, n3403, n3844, n2689, n3851, n2739, 
        n3521, n3864, n2876, n3897, n3901, n3900, n3899, n3898, n3944, n630, 
        n3965, n3068, n3438, n3514, n1390, n3974, n3976, n3975, n3977, n3984, 
        n3175, n3985, n3195, n3990, n1950, n3993, n3994, n3995, n2104, n3380, 
        n3529, n3534, n3522, n3515, N3014, N361, n1455, n1439, n3270, n2881, 
        n2879, n2465, n4002, n2808, n2206, n3058, n1970, n1912, n1387, n3100, 
        n1593, n1369, n3072, n3073, n1356, n3038, n2949, n2951, n2948, n2952, 
        N1734, n1288, n3868, n3870, n3869, n1855, n1854, n1310, n2894, n2895, 
        n1300, n2576, n1205, n2422, n1124, n2172, n2099, n1106, n1285, n3197, 
        n3431, n3432, n1536, n1041, n3634, n3633, n3632, n1048, n3661, n3660, 
        n3659, n3590, n1348, n3960, n3959, n3958, n849, n3972, n3971, n3439, 
        n2980, n2339, n3756, n3957, n3032, n3413, n3970, n1321, n3934, n3933, 
        n3932, n3774, n1314, n3909, n3908, n3907, n511, n2340, n3962, n1312, 
        n1301, n3883, n3882, n1286, n3867, n3866, n3865, n1316, n3850, n2718, 
        n3889, n3876, n2889, n596, n3342, n3875, n3437, n1431, n2781, n1258, 
        n1255, N1700, n1298, n3834, n3833, n3832, n3831, N1853, n1272, N1865, 
        n3427, n3428, n3429, n4130, N1757, N1858, n3735, n3507, n3508, n3440, 
        n3441, n3709, n3672, n3671, n3670, n1044, n3643, n3642, n3641, n1071, 
        n3675, n3674, n3673, n1096, N1738, N1837, n1274, N1799, n3583, n3177, 
        n1553, n1430, n1432, n1640, n3349, n4011, n2766, n1360, n3967, n3966, 
        n3651, n3649, n1392, n4142, n3512, n2137, n3698, n3621, n3617, n3655, 
        n2108, n1329, n3790, n2109, n3744, n1299, n3880, n2136, n3879, n2998, 
        n1287, n2960, n3896, n2926, n2935, n3887, n2140, n1114, n3913, n3857, 
        n2915, n2630, n3526, n3872, n3845, n3565, n1282, n2804, n3863, n3400, 
        n1259, n2744, n2633, n1115, n3772, n1645, n1771, n3743, n2411, n1554, 
        n3731, n3730, n2397, n2322, n2292, n2081, n3685, n2084, n3680, n2048, 
        n3580, n3183, n3184, n1174, n2335, n3980, n3979, n3356, n3505, n3567, 
        n3568, n3361, n3297, n3363, n3364, n3372, n3300, n3725, n3888, n3376, 
        n3295, n3569, n4013, n1113, N1869, n1248, n1148, n3453, n3791, n2305, 
        n3402, n1146, N1737, n3398, n3399, n3733, n2261, n3103, n1512, n3503, 
        n3517, n1388, n1382, N1809, n4119, n4118, n3089, n3088, n4122, n4121, 
        n4120, n3331, n4124, n3388, n4123, n730, n3873, N1710, n2050, n2046, 
        n2875, n732, n731, N348, n2055, n4126, n3890, n1567, n3686, n3393, 
        N1650, n1303, n2878, N1716, n2082, n4128, n3502, n3097, n3299, n2853, 
        n2563, n3359, n3360, n1010, n2425, n4131, n4132, n550, n911, n4133, 
        n3397, n990, n3679, n933, n932, n2426, ___cell__39620_net143598, N1859, 
        n2392, N1705, N1826, n929, N1654, n2809, n1731, n4135, net149617, 
        n2087, n4138, N1720, n3688, n2086, N1827, N1860, n918, n4014, n4016, 
        n602, n605, n3968, n837, n3231, n974, n4143, n4145, n4224, n1959, 
        n4156, n4158, n4160, n4162, n4164, n4166, n4168, n4170, n4172, n4174, 
        n4176, n4178, n4180, n4182, n3793, n4184, n4186, n4188, n4190, n4192, 
        n4194, n4196, n4198, n4200, n4202, n2483, n4203, n4204, n4206, n4208, 
        n4210, n4212, n4214, n4216, n4218, n4220, n2482, n4222, n505, n2461, 
        n1766, N1758, n2462, n1933, N1797, n1936, N1830, n3252, n1930, N1731, 
        n1929, N1698, n3249, n3250, n1934, N1996, n1932, N1930, n1935, N1963, 
        N1632, n3240, n3243, n1544, n3286, n3285, n3277, n1537, N307, n3982, 
        n716, N1841, n1394, N1709, N1874, n1515, n2787, n2786, n1826, N1652, 
        n2764, n3043, n1357, n1358, n1887, N1877, n1886, N1646, N1712, n1373, 
        n3267, n1370, n1371, N1843, n1895, N1876, n1362, N1711, n3157, n3156, 
        n3513, n3978, N1840, N1741, N1708, n3847, n2694, n2693, n1811, N1753, 
        n1131, n1132, n3708, n2132, n2129, n1125, N1868, n2672, n3874, n1843, 
        n2870, n3519, n3520, n1292, N1816, n1846, N1717, N1750, n3606, n1144, 
        n3700, N1702, n586, n1311, n3381, N1948, N1815, n2877, N1881, n1734, 
        N1993, n2307, n1735, N1960, n1737, N2026, n599, n3747, n3748, n2321, 
        n3771, n2434, n873, n2047, n3676, n1078, N1805, n1074, N1706, n2398, 
        n3768, n2304, n2406, n1747, n2287, ___cell__39620_net144307, n495, 
        n3728, n3736, n2272, n3732, n1154, n1155, n2005, n1927, N1931, n1928, 
        N1798, n3986, n1926, N1732, n3189, n3188, N1699, n1925, N1633, n3178, 
        n3201, n3663, n3586, n3587, n3581, n3650, n1046, n1280, N1707, n3956, 
        n3931, n3926, n2990, n3943, n3949, n3950, n3951, n2993, n3942, n3955, 
        n2997, n1346, N1845, n1341, N1812, n1336, N1713, n1326, n2959, n3941, 
        n939, n1870, N1879, N1648, n1325, ___cell__39620_net146132, N1714, 
        n1869, N1747, N1979, N1846, n1872, N1813, net149106, n2913, n2916, 
        n1860, N1715, n1859, N1649, n1862, N1880, N1847, N1980, n1864, N1814, 
        n2762, net156025, n1320, n3609, n2864, n3527, n3550, n1819, N1719, 
        N1851, n1931, N1863, N1951, byte_reg__m2s, mem_read_EX_reg__m2s, 
        mem_to_reg_EX_reg__m2s, n4201, mem_write_EX_reg__m2s, 
        reg_out_B_EX_reg_0__m2s, n4213, reg_out_B_EX_reg_10__m2s, n4209, n4183, 
        reg_out_B_EX_reg_11__m2s, n4215, reg_out_B_EX_reg_12__m2s, n4181, 
        reg_out_B_EX_reg_13__m2s, n4217, reg_out_B_EX_reg_14__m2s, n4179, 
        reg_out_B_EX_reg_15__m2s, n4159, reg_out_B_EX_reg_16__m2s, n4177, 
        reg_out_B_EX_reg_17__m2s, n4223, reg_out_B_EX_reg_18__m2s, n4211, 
        reg_out_B_EX_reg_19__m2s, n4175, reg_out_B_EX_reg_1__m2s, n4161, 
        reg_out_B_EX_reg_20__m2s, n4219, reg_out_B_EX_reg_21__m2s, n4163, 
        reg_out_B_EX_reg_22__m2s, n4205, reg_out_B_EX_reg_23__m2s, n4173, 
        reg_out_B_EX_reg_24__m2s, n4157, reg_out_B_EX_reg_25__m2s, n4171, 
        reg_out_B_EX_reg_26__m2s, n4207, reg_out_B_EX_reg_27__m2s, n4169, 
        reg_out_B_EX_reg_28__m2s, n4167, reg_out_B_EX_reg_29__m2s, n4221, 
        reg_out_B_EX_reg_2__m2s, n4197, reg_out_B_EX_reg_30__m2s, n4165, 
        reg_out_B_EX_reg_31__m2s, n4150, reg_out_B_EX_reg_3__m2s, n4195, 
        reg_out_B_EX_reg_4__m2s, n4193, reg_out_B_EX_reg_5__m2s, n4191, 
        reg_out_B_EX_reg_6__m2s, n4189, reg_out_B_EX_reg_7__m2s, n4187, 
        reg_out_B_EX_reg_8__m2s, n4185, reg_out_B_EX_reg_9__m2s, 
        reg_write_EX_reg__m2s, n4199, word_reg__m2s;
    assign word = test_so;
    smlatnr_2 ALU_result_reg_0__master ( .q(ALU_result_reg_0__m2s), .d(n4049), 
        .sdi(test_si), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4017), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_8 ALU_result_reg_0__slave ( .q(ALU_result[0]), .qb(n4018), .d(
        ALU_result_reg_0__m2s), .g(Ctrl__Regs_1__en2), .rb(n4017), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 ALU_result_reg_10__master ( .q(ALU_result_reg_10__m2s), .d(n4059
        ), .sdi(ALU_result[9]), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4017
        ), .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_4 ALU_result_reg_10__slave ( .q(ALU_result[10]), .qb(n4020), .d(
        ALU_result_reg_10__m2s), .g(Ctrl__Regs_1__en2), .rb(n4017), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_2 ALU_result_reg_11__master ( .q(ALU_result_reg_11__m2s), .d(n4060
        ), .sdi(ALU_result[10]), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n542
        ), .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_8 ALU_result_reg_11__slave ( .q(ALU_result[11]), .qb(n4021), .d(
        ALU_result_reg_11__m2s), .g(Ctrl__Regs_1__en2), .rb(n542), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 ALU_result_reg_12__master ( .q(ALU_result_reg_12__m2s), .d(n4061
        ), .sdi(ALU_result[11]), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n542
        ), .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_4 ALU_result_reg_12__slave ( .q(ALU_result[12]), .qb(n4154), .d(
        ALU_result_reg_12__m2s), .g(Ctrl__Regs_1__en2), .rb(n542), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 ALU_result_reg_13__master ( .q(ALU_result_reg_13__m2s), .d(n4062
        ), .sdi(n4154), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n543), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_4 ALU_result_reg_13__slave ( .q(ALU_result[13]), .qb(n4022), .d(
        ALU_result_reg_13__m2s), .g(Ctrl__Regs_1__en2), .rb(n543), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 ALU_result_reg_14__master ( .q(ALU_result_reg_14__m2s), .d(n4063
        ), .sdi(ALU_result[13]), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n543
        ), .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_4 ALU_result_reg_14__slave ( .q(ALU_result[14]), .qb(n4153), .d(
        ALU_result_reg_14__m2s), .g(Ctrl__Regs_1__en2), .rb(n543), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 ALU_result_reg_15__master ( .q(ALU_result_reg_15__m2s), .d(n4064
        ), .sdi(n4153), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n543), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 ALU_result_reg_15__slave ( .q(ALU_result[15]), .qb(n4023), .d(
        ALU_result_reg_15__m2s), .g(Ctrl__Regs_1__en2), .rb(n543), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 ALU_result_reg_16__master ( .q(ALU_result_reg_16__m2s), .d(n4065
        ), .sdi(ALU_result[15]), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n543
        ), .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 ALU_result_reg_16__slave ( .q(ALU_result[16]), .qb(n4024), .d(
        ALU_result_reg_16__m2s), .g(Ctrl__Regs_1__en2), .rb(n543), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 ALU_result_reg_17__master ( .q(ALU_result_reg_17__m2s), .d(n4066
        ), .sdi(ALU_result[16]), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(
        n4017), .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 ALU_result_reg_17__slave ( .q(ALU_result[17]), .qb(n4025), .d(
        ALU_result_reg_17__m2s), .g(Ctrl__Regs_1__en2), .rb(n4017), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 ALU_result_reg_18__master ( .q(ALU_result_reg_18__m2s), .d(n4067
        ), .sdi(ALU_result[17]), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n543
        ), .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_4 ALU_result_reg_18__slave ( .q(ALU_result[18]), .qb(n4152), .d(
        ALU_result_reg_18__m2s), .g(Ctrl__Regs_1__en2), .rb(n543), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 ALU_result_reg_19__master ( .q(ALU_result_reg_19__m2s), .d(n4068
        ), .sdi(n4152), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n543), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_4 ALU_result_reg_19__slave ( .q(ALU_result[19]), .qb(n4151), .d(
        ALU_result_reg_19__m2s), .g(Ctrl__Regs_1__en2), .rb(n543), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 ALU_result_reg_1__master ( .q(ALU_result_reg_1__m2s), .d(n4050), 
        .sdi(ALU_result[0]), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4017), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 ALU_result_reg_1__slave ( .q(ALU_result[1]), .qb(n4019), .d(
        ALU_result_reg_1__m2s), .g(Ctrl__Regs_1__en2), .rb(n4017), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_2 ALU_result_reg_20__master ( .q(ALU_result_reg_20__m2s), .d(n4069
        ), .sdi(n4151), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n542), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_8 ALU_result_reg_20__slave ( .q(ALU_result[20]), .qb(n4027), .d(
        ALU_result_reg_20__m2s), .g(Ctrl__Regs_1__en2), .rb(n542), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 ALU_result_reg_21__master ( .q(ALU_result_reg_21__m2s), .d(n4070
        ), .sdi(ALU_result[20]), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n542
        ), .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 ALU_result_reg_21__slave ( .q(ALU_result[21]), .qb(n4028), .d(
        ALU_result_reg_21__m2s), .g(Ctrl__Regs_1__en2), .rb(n542), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 ALU_result_reg_22__master ( .q(ALU_result_reg_22__m2s), .d(n4071
        ), .sdi(ALU_result[21]), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(
        n4017), .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_4 ALU_result_reg_22__slave ( .q(ALU_result[22]), .qb(n4029), .d(
        ALU_result_reg_22__m2s), .g(Ctrl__Regs_1__en2), .rb(n4017), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 ALU_result_reg_23__master ( .q(ALU_result_reg_23__m2s), .d(n4072
        ), .sdi(ALU_result[22]), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n543
        ), .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 ALU_result_reg_23__slave ( .q(ALU_result[23]), .qb(n4030), .d(
        ALU_result_reg_23__m2s), .g(Ctrl__Regs_1__en2), .rb(n543), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 ALU_result_reg_24__master ( .q(ALU_result_reg_24__m2s), .d(n4073
        ), .sdi(ALU_result[23]), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n542
        ), .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 ALU_result_reg_24__slave ( .q(ALU_result[24]), .qb(n4031), .d(
        ALU_result_reg_24__m2s), .g(Ctrl__Regs_1__en2), .rb(n542), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 ALU_result_reg_25__master ( .q(ALU_result_reg_25__m2s), .d(n4074
        ), .sdi(ALU_result[24]), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n543
        ), .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 ALU_result_reg_25__slave ( .q(ALU_result[25]), .qb(n4032), .d(
        ALU_result_reg_25__m2s), .g(Ctrl__Regs_1__en2), .rb(n543), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 ALU_result_reg_26__master ( .q(ALU_result_reg_26__m2s), .d(n4075
        ), .sdi(ALU_result[25]), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n542
        ), .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 ALU_result_reg_26__slave ( .q(ALU_result[26]), .qb(n4033), .d(
        ALU_result_reg_26__m2s), .g(Ctrl__Regs_1__en2), .rb(n542), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 ALU_result_reg_27__master ( .q(ALU_result_reg_27__m2s), .d(n4076
        ), .sdi(ALU_result[26]), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n542
        ), .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_4 ALU_result_reg_27__slave ( .q(ALU_result[27]), .qb(n4034), .d(
        ALU_result_reg_27__m2s), .g(Ctrl__Regs_1__en2), .rb(n542), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 ALU_result_reg_28__master ( .q(ALU_result_reg_28__m2s), .d(n4077
        ), .sdi(ALU_result[27]), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n542
        ), .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_4 ALU_result_reg_28__slave ( .q(ALU_result[28]), .qb(n4035), .d(
        ALU_result_reg_28__m2s), .g(Ctrl__Regs_1__en2), .rb(n542), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_2 ALU_result_reg_29__master ( .q(ALU_result_reg_29__m2s), .d(n4078
        ), .sdi(ALU_result[28]), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n543
        ), .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_8 ALU_result_reg_29__slave ( .q(ALU_result[29]), .qb(n4036), .d(
        ALU_result_reg_29__m2s), .g(Ctrl__Regs_1__en2), .rb(n543), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 ALU_result_reg_2__master ( .q(ALU_result_reg_2__m2s), .d(n4051), 
        .sdi(ALU_result[1]), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4017), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 ALU_result_reg_2__slave ( .q(ALU_result[2]), .qb(n4026), .d(
        ALU_result_reg_2__m2s), .g(Ctrl__Regs_1__en2), .rb(n4017), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_2 ALU_result_reg_30__master ( .q(ALU_result_reg_30__m2s), .d(n4079
        ), .sdi(ALU_result[29]), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(
        n4017), .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_8 ALU_result_reg_30__slave ( .q(ALU_result[30]), .qb(n4038), .d(
        ALU_result_reg_30__m2s), .g(Ctrl__Regs_1__en2), .rb(n4017), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_2 ALU_result_reg_31__master ( .q(ALU_result_reg_31__m2s), .d(
        _ALU_result_reg_31_net106451), .sdi(ALU_result[30]), .se(test_se), .g(
        Ctrl__Regs_1__en1), .rb(n4017), .glob_g(global_g1), .sync_sel(sync_sel
        ) );
    mlatnr_8 ALU_result_reg_31__slave ( .q(ALU_result[31]), .qb(n4039), .d(
        ALU_result_reg_31__m2s), .g(Ctrl__Regs_1__en2), .rb(n4017), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 ALU_result_reg_3__master ( .q(ALU_result_reg_3__m2s), .d(n4052), 
        .sdi(ALU_result[2]), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4017), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 ALU_result_reg_3__slave ( .q(ALU_result[3]), .qb(n4037), .d(
        ALU_result_reg_3__m2s), .g(Ctrl__Regs_1__en2), .rb(n4017), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 ALU_result_reg_4__master ( .q(ALU_result_reg_4__m2s), .d(n4053), 
        .sdi(ALU_result[3]), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4017), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 ALU_result_reg_4__slave ( .q(ALU_result[4]), .qb(n4040), .d(
        ALU_result_reg_4__m2s), .g(Ctrl__Regs_1__en2), .rb(n4017), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 ALU_result_reg_5__master ( .q(ALU_result_reg_5__m2s), .d(n4054), 
        .sdi(ALU_result[4]), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4017), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_4 ALU_result_reg_5__slave ( .q(ALU_result[5]), .qb(n4041), .d(
        ALU_result_reg_5__m2s), .g(Ctrl__Regs_1__en2), .rb(n4017), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 ALU_result_reg_6__master ( .q(ALU_result_reg_6__m2s), .d(n4055), 
        .sdi(ALU_result[5]), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n543), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 ALU_result_reg_6__slave ( .q(ALU_result[6]), .qb(n4042), .d(
        ALU_result_reg_6__m2s), .g(Ctrl__Regs_1__en2), .rb(n543), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 ALU_result_reg_7__master ( .q(ALU_result_reg_7__m2s), .d(n4056), 
        .sdi(ALU_result[6]), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n542), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_4 ALU_result_reg_7__slave ( .q(ALU_result[7]), .qb(n4043), .d(
        ALU_result_reg_7__m2s), .g(Ctrl__Regs_1__en2), .rb(n542), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 ALU_result_reg_8__master ( .q(ALU_result_reg_8__m2s), .d(n4057), 
        .sdi(ALU_result[7]), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n543), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_1 ALU_result_reg_8__slave ( .q(ALU_result[8]), .qb(n4044), .d(
        ALU_result_reg_8__m2s), .g(Ctrl__Regs_1__en2), .rb(n543), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 ALU_result_reg_9__master ( .q(ALU_result_reg_9__m2s), .d(n4058), 
        .sdi(ALU_result[8]), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n543), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 ALU_result_reg_9__slave ( .q(ALU_result[9]), .qb(n4045), .d(
        ALU_result_reg_9__m2s), .g(Ctrl__Regs_1__en2), .rb(n543), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    oai21_1 U100 ( .x(n3235), .a(n1577), .b(n1729), .c(n665) );
    inv_2 U1000 ( .x(n1964), .a(n1070) );
    nor2i_0 U1001 ( .x(n1235), .a(Imm[7]), .b(n734) );
    aoi21_1 U1002 ( .x(n2635), .a(N1754), .b(___cell__39620_net145150), .c(
        n1235) );
    nand2i_2 U1003 ( .x(n2639), .a(n1801), .b(n809) );
    inv_2 U1004 ( .x(n1801), .a(N1655) );
    nand2_2 U1005 ( .x(n2631), .a(n829), .b(n634) );
    nand2i_2 U1006 ( .x(n2638), .a(n2631), .b(___cell__39620_net145285) );
    nand2i_2 U1007 ( .x(n2645), .a(n1805), .b(n1987) );
    inv_2 U1008 ( .x(n1805), .a(N1820) );
    inv_5 U1009 ( .x(n1315), .a(n2722) );
    ao21_1 U101 ( .x(n3236), .a(n1147), .b(n1136), .c(n3235) );
    nand2i_2 U1010 ( .x(n2644), .a(n1055), .b(n2557) );
    inv_2 U1011 ( .x(n661), .a(n869) );
    inv_5 U1012 ( .x(n3648), .a(n844) );
    inv_2 U1013 ( .x(n1804), .a(N1953) );
    nand2i_2 U1014 ( .x(___cell__39620_net143845), .a(___cell__39620_net144360
        ), .b(n708) );
    nor2i_1 U1015 ( .x(n1236), .a(N1986), .b(___cell__39620_net143845) );
    oai211_2 U1016 ( .x(n3821), .a(n3460), .b(n1623), .c(n2602), .d(n3820) );
    nor2i_3 U1017 ( .x(n1233), .a(___cell__39620_net143864), .b(n1234) );
    inv_8 U1018 ( .x(n1322), .a(n1972) );
    oai221_4 U1019 ( .x(n2609), .a(n3418), .b(n4004), .c(n1322), .d(n1565), 
        .e(n1807) );
    nand2i_2 U102 ( .x(n3234), .a(n1625), .b(n2806) );
    aoi22_1 U1020 ( .x(n2608), .a(n649), .b(n2609), .c(n650), .d(n2574) );
    oai21_1 U1021 ( .x(n2604), .a(n1486), .b(n690), .c(n2605) );
    inv_2 U1022 ( .x(n1063), .a(n646) );
    inv_2 U1023 ( .x(n2607), .a(n3826) );
    nand2i_0 U1024 ( .x(n2620), .a(___cell__39620_net144707), .b(
        ___cell__39620_net145617) );
    inv_8 U1025 ( .x(n811), .a(n606) );
    nor2i_1 U1026 ( .x(n1228), .a(N1854), .b(n946) );
    inv_2 U1027 ( .x(n1230), .a(N1821) );
    nor2_1 U1028 ( .x(n1229), .a(n1077), .b(n1230) );
    inv_2 U1029 ( .x(n1795), .a(N1954) );
    mux2i_1 U103 ( .x(n3239), .d0(___cell__39620_net144201), .sl(net152465), 
        .d1(___cell__39620_net145285) );
    inv_2 U1030 ( .x(n1794), .a(N1887) );
    nand2i_2 U1031 ( .x(n2595), .a(n1794), .b(n3997) );
    nor2i_1 U1032 ( .x(n1226), .a(N1755), .b(___cell__39620_net143710) );
    aoi211_1 U1033 ( .x(n2594), .a(N1722), .b(___cell__39620_net145190), .c(
        n1227), .d(n1226) );
    nand2i_2 U1034 ( .x(n2593), .a(n1793), .b(n809) );
    inv_2 U1035 ( .x(n1793), .a(N1656) );
    inv_2 U1036 ( .x(n1788), .a(N1955) );
    inv_2 U1037 ( .x(n1214), .a(N1822) );
    nor2_1 U1038 ( .x(n1213), .a(n1077), .b(n1214) );
    oai221_3 U1039 ( .x(n565), .a(n1302), .b(n1043), .c(n3524), .d(n4007), .e(
        n1806) );
    nand2i_2 U104 ( .x(n1653), .a(n497), .b(n676) );
    aoi21_1 U1040 ( .x(n2546), .a(N1756), .b(___cell__39620_net145150), .c(
        n1212) );
    nand2i_2 U1041 ( .x(n2549), .a(n1785), .b(n809) );
    inv_2 U1042 ( .x(n1785), .a(N1657) );
    nand2_2 U1043 ( .x(n2545), .a(n689), .b(n590) );
    nand2i_2 U1044 ( .x(n2548), .a(n2545), .b(___cell__39620_net145285) );
    nor2_1 U1045 ( .x(n1060), .a(n1061), .b(n645) );
    nand2i_2 U1046 ( .x(n1531), .a(IR_function_field[1]), .b(IR_function_field
        [0]) );
    aoi21_1 U1047 ( .x(n2566), .a(___cell__39620_net144517), .b(n2375), .c(
        n2564) );
    nand2i_2 U1048 ( .x(n3811), .a(n1625), .b(n2649) );
    inv_5 U1049 ( .x(n2266), .a(n1091) );
    nor2_1 U105 ( .x(n1427), .a(n1428), .b(n1429) );
    nand3_1 U1050 ( .x(n3812), .a(n2562), .b(n3811), .c(n2566) );
    nand2i_2 U1051 ( .x(n2584), .a(n688), .b(___cell__39620_net145617) );
    inv_8 U1052 ( .x(n3385), .a(n3384) );
    inv_2 U1053 ( .x(n3444), .a(n3443) );
    nor2i_1 U1054 ( .x(n1650), .a(n2001), .b(n1539) );
    oai22_1 U1055 ( .x(n2560), .a(n2475), .b(n1687), .c(n1648), .d(n1690) );
    aoi21_1 U1056 ( .x(n2561), .a(n1256), .b(n2477), .c(n2560) );
    nand2i_2 U1057 ( .x(n3815), .a(n1578), .b(n3684) );
    inv_5 U1058 ( .x(n1578), .a(reg_out_A[24]) );
    inv_2 U1059 ( .x(n3447), .a(n2738) );
    nor2_1 U106 ( .x(n3232), .a(n3229), .b(n3230) );
    nand2_2 U1060 ( .x(n3813), .a(n1249), .b(n2738) );
    nor2i_1 U1061 ( .x(n1220), .a(n1221), .b(n1222) );
    inv_2 U1062 ( .x(n1222), .a(n2492) );
    nand2i_2 U1063 ( .x(n2572), .a(n1484), .b(n2139) );
    exnor2_1 U1064 ( .x(n1483), .a(n590), .b(n689) );
    oai21_1 U1065 ( .x(n2571), .a(n1483), .b(n690), .c(n2572) );
    nor2_0 U1066 ( .x(n2543), .a(n1626), .b(net149120) );
    nand2i_2 U1067 ( .x(n1218), .a(n1781), .b(n530) );
    aoi21_1 U1068 ( .x(n1216), .a(n1217), .b(n1218), .c(n1219) );
    nor2i_1 U1069 ( .x(n2544), .a(n1451), .b(n670) );
    nor2_1 U107 ( .x(n3228), .a(n3226), .b(n3227) );
    nand4_1 U1070 ( .x(n3782), .a(n2480), .b(n3781), .c(n2479), .d(n3780) );
    inv_2 U1071 ( .x(n2435), .a(n1711) );
    inv_2 U1072 ( .x(n2436), .a(n1712) );
    nand2i_2 U1073 ( .x(n3780), .a(n1623), .b(n2649) );
    nand2i_2 U1074 ( .x(n1443), .a(n1659), .b(n1542) );
    inv_2 U1075 ( .x(n1542), .a(n1539) );
    nand2i_2 U1076 ( .x(n1539), .a(IR_function_field[5]), .b(n1540) );
    inv_2 U1077 ( .x(n1540), .a(n1538) );
    inv_2 U1078 ( .x(n1661), .a(n1443) );
    oai22_1 U1079 ( .x(n2474), .a(n1648), .b(n1715), .c(n2475), .d(n1713) );
    nor2_1 U108 ( .x(n3225), .a(n3223), .b(n3224) );
    aoi21_1 U1080 ( .x(n2476), .a(n1249), .b(n2477), .c(n2474) );
    nand2i_2 U1081 ( .x(n3784), .a(n4009), .b(n2286) );
    oai211_2 U1082 ( .x(n2286), .a(n507), .b(n1546), .c(n3407), .d(n3408) );
    aoi21_1 U1083 ( .x(n2478), .a(n1256), .b(n2373), .c(n1194) );
    nand2i_2 U1084 ( .x(___cell__39620_net144302), .a(n1533), .b(n675) );
    nor2i_0 U1085 ( .x(n1619), .a(IR_opcode_field[0]), .b(n1519) );
    nand2_2 U1086 ( .x(n1618), .a(n1619), .b(___cell__39620_net144303) );
    inv_2 U1087 ( .x(n1061), .a(n1531) );
    nand2i_2 U1088 ( .x(n1525), .a(n1523), .b(n1526) );
    nand2_2 U1089 ( .x(n3798), .a(n1249), .b(n2779) );
    nor2_1 U109 ( .x(n3222), .a(n3220), .b(n3221) );
    inv_2 U1090 ( .x(n3684), .a(n1093) );
    nand2i_2 U1091 ( .x(n3799), .a(n1219), .b(n3684) );
    nand2_2 U1092 ( .x(n3797), .a(n1714), .b(n2306) );
    inv_2 U1093 ( .x(n1150), .a(n1687) );
    aoi222_1 U1094 ( .x(n2518), .a(n1256), .b(n2433), .c(n1150), .d(n2270), 
        .e(n2273), .f(n904) );
    nand2i_2 U1095 ( .x(n1590), .a(IR_function_field[2]), .b(n1526) );
    inv_2 U1096 ( .x(n1526), .a(n1522) );
    or3i_1 U1097 ( .x(n1522), .a(IR_function_field[5]), .b(IR_function_field
        [4]), .c(IR_function_field[3]) );
    inv_8 U1098 ( .x(n1217), .a(n1700) );
    inv_5 U1099 ( .x(n3779), .a(n3778) );
    nor2_1 U110 ( .x(n3281), .a(n1939), .b(n1951) );
    nand2i_2 U1100 ( .x(n3806), .a(n670), .b(n3778) );
    inv_14 U1101 ( .x(n915), .a(n813) );
    inv_2 U1102 ( .x(n3386), .a(n2568) );
    exnor2_1 U1103 ( .x(n1481), .a(n540), .b(Imm[26]) );
    inv_2 U1104 ( .x(n3810), .a(n1481) );
    inv_2 U1105 ( .x(___cell__39620_net144201), .a(___cell__39620_net144199)
         );
    nand2_2 U1106 ( .x(n1116), .a(___cell__39620_net147732), .b(
        ___cell__39620_net144201) );
    nand2_2 U1107 ( .x(n2526), .a(n2193), .b(n3810) );
    exnor2_1 U1108 ( .x(n1482), .a(n540), .b(reg_out_B[26]) );
    nand2i_2 U1109 ( .x(n2525), .a(n1482), .b(n2139) );
    inv_5 U111 ( .x(n1093), .a(n737) );
    nand2_2 U1110 ( .x(n3801), .a(n3315), .b(n855) );
    inv_10 U1111 ( .x(n882), .a(n825) );
    inv_2 U1112 ( .x(n2432), .a(n1122) );
    oai21_1 U1113 ( .x(n3739), .a(n536), .b(n3738), .c(n1807) );
    inv_2 U1114 ( .x(n3738), .a(n2629) );
    inv_2 U1115 ( .x(n854), .a(n1807) );
    inv_2 U1116 ( .x(n1330), .a(n1565) );
    nand2i_4 U1117 ( .x(n2981), .a(n3585), .b(n3783) );
    nand2i_2 U1118 ( .x(n3425), .a(n1565), .b(n2981) );
    nand2i_0 U1119 ( .x(n3424), .a(n1559), .b(n1728) );
    nor2i_1 U112 ( .x(n1442), .a(n1443), .b(n1444) );
    nand2i_2 U1120 ( .x(n1582), .a(n1451), .b(n1545) );
    nand2_2 U1121 ( .x(n3762), .a(n3343), .b(n855) );
    nand2i_2 U1124 ( .x(n1160), .a(n1568), .b(n1543) );
    nor2i_1 U1125 ( .x(n1612), .a(IR_opcode_field[0]), .b(IR_opcode_field[1])
         );
    inv_8 U1126 ( .x(n1302), .a(n2677) );
    nor2_1 U1127 ( .x(n1207), .a(n734), .b(n1208) );
    nand2i_3 U1128 ( .x(n2506), .a(n1775), .b(n809) );
    nand2_0 U1129 ( .x(n2502), .a(Imm[26]), .b(n540) );
    oai21_1 U113 ( .x(n3280), .a(n1442), .b(n1093), .c(n3281) );
    nand2i_2 U1130 ( .x(n2505), .a(n2502), .b(___cell__39620_net147791) );
    nand2i_2 U1131 ( .x(___cell__39620_net144360), .a(n675), .b(n810) );
    oai21_3 U1132 ( .x(n3726), .a(n4125), .b(n1290), .c(n1806) );
    inv_8 U1133 ( .x(n1198), .a(n2423) );
    nand2i_2 U1134 ( .x(n2363), .a(n1742), .b(n2837) );
    inv_2 U1135 ( .x(n1742), .a(N310) );
    inv_2 U1136 ( .x(n571), .a(n3435) );
    nand2i_1 U1137 ( .x(n2361), .a(n1186), .b(n2197) );
    nand2i_2 U1138 ( .x(n2356), .a(n621), .b(n3757) );
    oai21_1 U1139 ( .x(n2352), .a(n1473), .b(n690), .c(n2353) );
    nor2_1 U114 ( .x(n3275), .a(n3272), .b(n3273) );
    nand4i_1 U1140 ( .x(n2354), .a(n2352), .b(n2355), .c(n2356), .d(n2357) );
    inv_2 U1141 ( .x(___cell__39620_net145524), .a(___cell__39620_net145444)
         );
    oai221_1 U1142 ( .x(n2365), .a(n2366), .b(n1647), .c(
        ___cell__39620_net145524), .d(n1646), .e(n2367) );
    nand4i_1 U1143 ( .x(n2364), .a(n2365), .b(n2368), .c(n2369), .d(n2370) );
    nand4_1 U1144 ( .x(n1173), .a(n2347), .b(n2345), .c(n2348), .d(n2349) );
    nand2i_2 U1145 ( .x(n2347), .a(n1182), .b(n2168) );
    nand2i_2 U1146 ( .x(n2348), .a(n1055), .b(n2165) );
    nand2i_2 U1147 ( .x(n2349), .a(n1743), .b(n809) );
    inv_2 U1148 ( .x(n1743), .a(N1635) );
    nor2i_1 U1149 ( .x(n1167), .a(N1833), .b(n946) );
    and3i_1 U115 ( .x(n3271), .a(n3264), .b(n3265), .c(n3268) );
    nor2i_1 U1150 ( .x(n1168), .a(N1999), .b(n1169) );
    aoi211_1 U1151 ( .x(n1172), .a(N1966), .b(___cell__39620_net145508), .c(
        n1168), .d(n1167) );
    inv_2 U1152 ( .x(n1745), .a(N1933) );
    nand2i_2 U1153 ( .x(n1171), .a(n1745), .b(n3662) );
    nor2i_2 U1154 ( .x(n1164), .a(n1165), .b(n1166) );
    aoi21_1 U1155 ( .x(n2346), .a(N1701), .b(___cell__39620_net145190), .c(
        n1163) );
    inv_2 U1156 ( .x(n1746), .a(N1800) );
    nand2i_2 U1157 ( .x(n2351), .a(n1746), .b(n1987) );
    inv_2 U1158 ( .x(n1744), .a(N1866) );
    nand2i_2 U1159 ( .x(n2350), .a(n1744), .b(n3997) );
    nor2_1 U116 ( .x(n3263), .a(n3261), .b(n3262) );
    aoi221_1 U1160 ( .x(n2836), .a(n692), .b(n1733), .c(n917), .d(
        ___cell__39620_net145444), .e(n2838) );
    nand2i_2 U1161 ( .x(n2835), .a(n1647), .b(n3705) );
    inv_2 U1162 ( .x(n1589), .a(n1582) );
    oai211_2 U1163 ( .x(n2834), .a(n2360), .b(n1588), .c(n2835), .d(n2836) );
    inv_5 U1164 ( .x(n1428), .a(n1639) );
    ao22_2 U1165 ( .x(n2825), .a(n502), .b(n2826), .c(n1267), .d(n2827) );
    inv_2 U1166 ( .x(n2829), .a(n1496) );
    aoi21_1 U1167 ( .x(n2828), .a(n2139), .b(n2829), .c(n1284) );
    aoai211_1 U1168 ( .x(n2824), .a(n692), .b(n530), .c(n1064), .d(n815) );
    nand2i_2 U1169 ( .x(n2823), .a(n670), .b(n3757) );
    nor3i_1 U117 ( .x(n3260), .a(n1518), .b(n3258), .c(n3259) );
    inv_2 U1170 ( .x(n1436), .a(n1620) );
    inv_2 U1171 ( .x(n2822), .a(n3760) );
    aoi211_1 U1172 ( .x(n2814), .a(N1733), .b(___cell__39620_net145150), .c(
        n1271), .d(n1270) );
    inv_2 U1173 ( .x(n1838), .a(N1634) );
    nand2i_2 U1174 ( .x(n2816), .a(n1838), .b(n809) );
    nand2i_2 U1175 ( .x(n2815), .a(n1182), .b(n2165) );
    inv_2 U1176 ( .x(n1839), .a(N1932) );
    nand2i_2 U1177 ( .x(n2820), .a(n1839), .b(n3999) );
    inv_2 U1178 ( .x(n1841), .a(N1965) );
    nand2i_2 U1179 ( .x(n2819), .a(n1841), .b(___cell__39620_net145508) );
    inv_5 U118 ( .x(n1585), .a(n608) );
    inv_2 U1180 ( .x(n1840), .a(N1832) );
    nand2i_2 U1181 ( .x(n2818), .a(n1840), .b(n4000) );
    nand2i_2 U1182 ( .x(n1275), .a(n1842), .b(n3624) );
    inv_2 U1183 ( .x(n1842), .a(N1998) );
    inv_2 U1184 ( .x(n1692), .a(N313) );
    inv_2 U1185 ( .x(n2142), .a(n2197) );
    oai211_1 U1186 ( .x(n2141), .a(n2142), .b(n1566), .c(n2138), .d(n2134) );
    nand2i_2 U1187 ( .x(n2155), .a(n621), .b(n3693) );
    aoi22_1 U1188 ( .x(n2156), .a(n2157), .b(n1085), .c(n2106), .d(n1204) );
    inv_2 U1189 ( .x(n1693), .a(N346) );
    exnor2_1 U119 ( .x(n1508), .a(reg_out_B[14]), .b(n644) );
    inv_2 U1190 ( .x(n1694), .a(N2002) );
    inv_2 U1191 ( .x(n1696), .a(N1936) );
    nand2i_2 U1192 ( .x(n3697), .a(n1696), .b(n3999) );
    inv_2 U1193 ( .x(n1699), .a(N1969) );
    nand2i_2 U1194 ( .x(n2125), .a(n1699), .b(___cell__39620_net145508) );
    inv_2 U1195 ( .x(n1698), .a(N1803) );
    nand2i_2 U1196 ( .x(n2124), .a(n1698), .b(n1987) );
    inv_2 U1197 ( .x(n1697), .a(N1836) );
    nand2i_2 U1198 ( .x(n2123), .a(n1697), .b(n4000) );
    and4i_1 U1199 ( .x(n2122), .a(n2121), .b(n2123), .c(n2124), .d(n2125) );
    nand2_2 U120 ( .x(n3631), .a(n3559), .b(___cell__39620_net144331) );
    aoi21_1 U1200 ( .x(n2120), .a(N1704), .b(___cell__39620_net145190), .c(
        n1111) );
    inv_2 U1201 ( .x(n1695), .a(N1638) );
    nand2i_2 U1202 ( .x(n2119), .a(n1695), .b(n809) );
    nand2i_2 U1203 ( .x(n2118), .a(n1166), .b(n2168) );
    aoi22_1 U1204 ( .x(n3104), .a(n650), .b(n3078), .c(n1221), .d(n3000) );
    aoi221_1 U1205 ( .x(n3101), .a(n1204), .b(n3075), .c(n649), .d(n2014), .e(
        n3102) );
    aoi21_1 U1206 ( .x(n3109), .a(n2022), .b(n3110), .c(n1389) );
    aoi222_1 U1207 ( .x(n3115), .a(n3118), .b(___cell__39620_net143864), .c(
        n894), .d(n1700), .e(ALU_result[12]), .f(n3057) );
    nand2i_2 U1208 ( .x(n3107), .a(n1900), .b(n977) );
    inv_2 U1209 ( .x(n1900), .a(N352) );
    nand2i_2 U121 ( .x(n3961), .a(n1625), .b(n3291) );
    inv_2 U1210 ( .x(n1906), .a(N1975) );
    nand2i_2 U1211 ( .x(n3096), .a(n1906), .b(___cell__39620_net145508) );
    inv_2 U1212 ( .x(n1905), .a(N1842) );
    nand2i_2 U1213 ( .x(n3095), .a(n1905), .b(n735) );
    aoi22_1 U1214 ( .x(n3094), .a(n1095), .b(n1988), .c(n1197), .d(n1397) );
    aoi21_1 U1215 ( .x(n3093), .a(n662), .b(n594), .c(n1381) );
    nand4_1 U1216 ( .x(n1386), .a(n3093), .b(n3094), .c(n3095), .d(n3096) );
    nand2i_2 U1217 ( .x(n1385), .a(n1901), .b(n3624) );
    inv_2 U1218 ( .x(n1901), .a(N2008) );
    inv_2 U1219 ( .x(n1904), .a(N1942) );
    ao22_2 U122 ( .x(n712), .a(n526), .b(n1256), .c(n504), .d(n3020) );
    nand2i_2 U1220 ( .x(n1384), .a(n1904), .b(n3999) );
    nor2i_3 U1221 ( .x(n1379), .a(n1380), .b(n1055) );
    inv_2 U1222 ( .x(n1903), .a(N1875) );
    nand2i_2 U1223 ( .x(n3092), .a(n1903), .b(n3997) );
    aoi211_1 U1224 ( .x(n3090), .a(N1644), .b(n809), .c(n1378), .d(n1376) );
    inv_2 U1225 ( .x(n1902), .a(N1743) );
    nand2i_2 U1226 ( .x(n3091), .a(n1902), .b(___cell__39620_net145150) );
    and4i_1 U1227 ( .x(n1383), .a(n1379), .b(n3091), .c(n3090), .d(n3092) );
    inv_2 U1228 ( .x(n1675), .a(N347) );
    nand2i_2 U1229 ( .x(n2095), .a(n1675), .b(n977) );
    nand2_2 U123 ( .x(n3547), .a(n3548), .b(n3549) );
    aoi22_1 U1231 ( .x(n2088), .a(n649), .b(n2089), .c(n650), .d(n2090) );
    nand4_1 U1232 ( .x(n2094), .a(n2091), .b(n2088), .c(n2092), .d(n2095) );
    inv_2 U1233 ( .x(n589), .a(n2135) );
    aoi221_3 U1234 ( .x(n2096), .a(n2106), .b(___cell__39620_net143864), .c(
        n2107), .d(n1204), .e(n2103) );
    inv_2 U1235 ( .x(n1681), .a(N1970) );
    nand2i_2 U1236 ( .x(n2077), .a(n1681), .b(___cell__39620_net145508) );
    inv_2 U1237 ( .x(n1680), .a(N1804) );
    nand2i_2 U1238 ( .x(n2076), .a(n1680), .b(n1987) );
    aoi22_1 U1239 ( .x(n2074), .a(n1318), .b(n1993), .c(n662), .d(n1992) );
    inv_5 U124 ( .x(n2273), .a(n1690) );
    aoi21_1 U1240 ( .x(n2075), .a(n1197), .b(n2043), .c(n1099) );
    nand4_1 U1241 ( .x(n1103), .a(n2075), .b(n2074), .c(n2076), .d(n2077) );
    nand2i_2 U1242 ( .x(n1102), .a(n1677), .b(n3624) );
    inv_2 U1243 ( .x(n1677), .a(N2003) );
    inv_2 U1244 ( .x(n1679), .a(N1937) );
    nand2i_2 U1245 ( .x(n1101), .a(n1679), .b(n3662) );
    nand2i_2 U1246 ( .x(n2071), .a(n2068), .b(___cell__39620_net145285) );
    inv_2 U1247 ( .x(n1678), .a(N1639) );
    nand2i_2 U1248 ( .x(n2072), .a(n1678), .b(n809) );
    nand2i_2 U1249 ( .x(n2501), .a(___cell__39620_net144406), .b(n3785) );
    inv_4 U125 ( .x(n3352), .a(n658) );
    nand2i_2 U1250 ( .x(n2500), .a(n784), .b(n3782) );
    aoi21_1 U1251 ( .x(n2498), .a(n1085), .b(n2499), .c(n1206) );
    nand2i_2 U1253 ( .x(n2496), .a(n1761), .b(n2837) );
    inv_2 U1254 ( .x(n1761), .a(N334) );
    and4i_3 U1255 ( .x(n2493), .a(n2494), .b(n2491), .c(n2488), .d(n2484) );
    aoi22_1 U1256 ( .x(n2491), .a(n650), .b(n2492), .c(n1221), .d(n2400) );
    aoi22_1 U1257 ( .x(n2488), .a(n539), .b(n2489), .c(n535), .d(n2490) );
    and4i_3 U1258 ( .x(n2484), .a(n2481), .b(n2485), .c(n2486), .d(n2487) );
    inv_2 U1259 ( .x(n2494), .a(n3794) );
    and2_5 U126 ( .x(n512), .a(n3352), .b(n3353) );
    nand2i_2 U1260 ( .x(n3794), .a(n1566), .b(n3422) );
    inv_5 U1261 ( .x(n1760), .a(reg_out_B[27]) );
    inv_5 U1262 ( .x(n680), .a(Imm[27]) );
    oai21_2 U1263 ( .x(n2399), .a(n3419), .b(n1565), .c(n3571) );
    aoi222_1 U1264 ( .x(n2495), .a(n1191), .b(n2399), .c(n681), .d(
        ___cell__39620_net145617), .e(reg_out_B[27]), .f(n1064) );
    inv_8 U1265 ( .x(n1573), .a(reg_out_A[26]) );
    inv_2 U1266 ( .x(n1769), .a(N1857) );
    nand2i_2 U1267 ( .x(n2472), .a(n1769), .b(n735) );
    inv_2 U1268 ( .x(n1768), .a(N1824) );
    nand2i_2 U1269 ( .x(n2471), .a(n1768), .b(n1987) );
    oai22_1 U127 ( .x(n2131), .a(n512), .b(n1687), .c(n1570), .d(n1690) );
    inv_2 U1270 ( .x(n1770), .a(N1990) );
    nand2i_2 U1271 ( .x(n2470), .a(n1770), .b(___cell__39620_net145508) );
    aoi21_1 U1272 ( .x(n2469), .a(n1095), .b(n2473), .c(n1196) );
    nand2i_2 U1273 ( .x(n1201), .a(n1763), .b(n3624) );
    inv_2 U1274 ( .x(n1763), .a(N2023) );
    inv_2 U1275 ( .x(n1162), .a(n2384) );
    inv_2 U1276 ( .x(n1764), .a(N1659) );
    inv_2 U1277 ( .x(n1765), .a(N1725) );
    aoi21_1 U1278 ( .x(n3244), .a(___cell__39620_net143785), .b(n3245), .c(
        n1438) );
    and4i_3 U1279 ( .x(n3248), .a(n3251), .b(n3253), .c(n3254), .d(n3255) );
    nor2i_0 U128 ( .x(n1110), .a(n922), .b(n1093) );
    ao21_3 U1280 ( .x(n1440), .a(n3992), .b(n3991), .c(n1609) );
    inv_2 U1281 ( .x(n2004), .a(n1937) );
    inv_2 U1282 ( .x(n1638), .a(n1627) );
    aoi221_1 U1283 ( .x(n3290), .a(n1638), .b(n3214), .c(N340), .d(n1597), .e(
        n1445) );
    aoi221_3 U1284 ( .x(n3287), .a(n1576), .b(n3288), .c(n1589), .d(n3289), 
        .e(n1453) );
    nand2i_2 U1285 ( .x(n3131), .a(n1574), .b(n2014) );
    oai21_1 U1287 ( .x(n3129), .a(n3130), .b(n1566), .c(n3131) );
    nand2i_2 U1288 ( .x(n3134), .a(n1908), .b(n2837) );
    inv_2 U1289 ( .x(n1908), .a(N318) );
    nand2i_2 U1290 ( .x(n3133), .a(n1588), .b(n3078) );
    oai211_1 U1291 ( .x(n3126), .a(n1403), .b(n1907), .c(n3127), .d(n3128) );
    aoi21_1 U1292 ( .x(n3132), .a(n1221), .b(n3041), .c(n3126) );
    nand2_1 U1293 ( .x(n3147), .a(n1085), .b(n3117) );
    nand2_2 U1294 ( .x(n3146), .a(n3170), .b(___cell__39620_net143864) );
    inv_5 U1295 ( .x(n900), .a(reg_out_A[11]) );
    nand2i_2 U1296 ( .x(n3137), .a(n1909), .b(n977) );
    inv_2 U1297 ( .x(n1909), .a(N351) );
    inv_14 U1298 ( .x(___cell__39620_net144655), .a(Imm[11]) );
    and4i_3 U1299 ( .x(n3135), .a(n3139), .b(n3141), .c(n3142), .d(n3143) );
    nand2i_2 U130 ( .x(n3710), .a(n4008), .b(n2806) );
    nand2_2 U1300 ( .x(n3141), .a(n2024), .b(n3116) );
    nand2_2 U1301 ( .x(n3142), .a(n2022), .b(n3113) );
    inv_2 U1302 ( .x(n1915), .a(N1974) );
    nand2i_2 U1303 ( .x(n3125), .a(n1915), .b(___cell__39620_net145508) );
    inv_2 U1304 ( .x(n1914), .a(N1808) );
    nand2i_2 U1305 ( .x(n3124), .a(n1914), .b(n1987) );
    aoi22_1 U1306 ( .x(n3123), .a(n1095), .b(n1054), .c(n1197), .d(n1988) );
    nand2i_2 U1307 ( .x(n1401), .a(n1910), .b(n3624) );
    inv_2 U1308 ( .x(n1910), .a(N2007) );
    inv_2 U1309 ( .x(n1913), .a(N1941) );
    nand2i_2 U131 ( .x(n4010), .a(n694), .b(n891) );
    nand2i_2 U1310 ( .x(n1400), .a(n1913), .b(n3662) );
    nor2i_3 U1311 ( .x(n1396), .a(n1397), .b(n1055) );
    aoi211_1 U1312 ( .x(n3119), .a(N1643), .b(n809), .c(n1395), .d(n1393) );
    inv_2 U1313 ( .x(n1911), .a(N1742) );
    nand2i_2 U1314 ( .x(n3120), .a(n1911), .b(___cell__39620_net145150) );
    and4i_3 U1315 ( .x(n1399), .a(n1396), .b(n3120), .c(n3121), .d(n3119) );
    aoi22_1 U1316 ( .x(n2796), .a(n2797), .b(n2022), .c(n513), .d(n2024) );
    nand2i_2 U1317 ( .x(n2800), .a(n702), .b(n570) );
    nand2i_2 U1318 ( .x(n2794), .a(n1824), .b(n2837) );
    inv_2 U1319 ( .x(n1824), .a(N327) );
    nand2_4 U132 ( .x(n2184), .a(n3354), .b(n1558) );
    ao22_3 U1320 ( .x(n2788), .a(n2902), .b(n649), .c(n2863), .d(n650) );
    nor2i_2 U1321 ( .x(n1266), .a(n1267), .b(n1268) );
    inv_5 U1322 ( .x(n3368), .a(n3365) );
    or3i_2 U1323 ( .x(n1265), .a(n2768), .b(n2767), .c(n1260) );
    oai22_1 U1324 ( .x(n2767), .a(___cell__39620_net143710), .b(n1828), .c(
        ___cell__39620_net143660), .d(n1827) );
    inv_2 U1325 ( .x(n1828), .a(N1751) );
    inv_2 U1326 ( .x(n1827), .a(N1718) );
    nor2_1 U1327 ( .x(n1260), .a(n947), .b(n1261) );
    inv_2 U1328 ( .x(n1261), .a(N1883) );
    inv_2 U1329 ( .x(n1833), .a(N2016) );
    ao22_4 U133 ( .x(n1999), .a(n627), .b(n3584), .c(n3448), .d(n659) );
    nand2i_2 U1330 ( .x(n1264), .a(n1833), .b(n3624) );
    inv_2 U1331 ( .x(n1829), .a(N1950) );
    nand2i_2 U1332 ( .x(n1263), .a(n1829), .b(n3662) );
    inv_8 U1333 ( .x(n2774), .a(n3856) );
    inv_2 U1334 ( .x(n1832), .a(N1983) );
    nand2i_2 U1335 ( .x(n2777), .a(n1832), .b(___cell__39620_net145508) );
    inv_2 U1336 ( .x(n1831), .a(N1850) );
    nand2i_2 U1337 ( .x(n2776), .a(n1831), .b(n4000) );
    inv_2 U1338 ( .x(n1830), .a(N1817) );
    nand2i_2 U1339 ( .x(n2775), .a(n1830), .b(n1987) );
    nand2i_2 U134 ( .x(n3701), .a(n4009), .b(n3196) );
    nand2i_2 U1340 ( .x(n3046), .a(n1588), .b(n3001) );
    aoi221_2 U1341 ( .x(n3039), .a(___cell__39620_net143864), .b(n3040), .c(
        n649), .d(n3041), .e(n3042) );
    aoi22_1 U1342 ( .x(n3050), .a(n2024), .b(n3012), .c(n1267), .d(n3051) );
    aoi21_1 U1343 ( .x(n3049), .a(n2022), .b(n3008), .c(n1359) );
    inv_2 U1344 ( .x(n3055), .a(n3964) );
    aoi21_1 U1345 ( .x(n3052), .a(n502), .b(n3054), .c(n3055) );
    nand2i_2 U1346 ( .x(n3047), .a(n1884), .b(n977) );
    inv_2 U1347 ( .x(n1884), .a(N354) );
    inv_2 U1348 ( .x(n1889), .a(N1844) );
    nand2i_2 U1349 ( .x(n3031), .a(n1889), .b(n4000) );
    aoi21_1 U135 ( .x(n2186), .a(n1249), .b(n2187), .c(n1121) );
    aoi22_1 U1350 ( .x(n3028), .a(N1811), .b(n1987), .c(n662), .d(n1339) );
    inv_2 U1351 ( .x(n1890), .a(N1977) );
    nand2i_2 U1352 ( .x(n3030), .a(n1890), .b(___cell__39620_net145508) );
    nand2i_2 U1353 ( .x(n1354), .a(n1885), .b(n3624) );
    inv_2 U1354 ( .x(n1885), .a(N2010) );
    inv_2 U1355 ( .x(n1888), .a(N1944) );
    nand2i_2 U1356 ( .x(n1353), .a(n1888), .b(n3999) );
    nor2i_1 U1357 ( .x(n1351), .a(N1745), .b(___cell__39620_net143710) );
    nand4i_1 U1358 ( .x(n3024), .a(n1350), .b(n3025), .c(n3026), .d(n3027) );
    nand4i_3 U1359 ( .x(n2989), .a(n1323), .b(n3937), .c(n3936), .d(n3935) );
    oai22_1 U136 ( .x(n2230), .a(n1570), .b(n1715), .c(n512), .d(n1713) );
    inv_2 U1360 ( .x(n3079), .a(n3973) );
    nand2i_2 U1361 ( .x(n3086), .a(n1892), .b(n977) );
    inv_2 U1362 ( .x(n1892), .a(N353) );
    ao21_3 U1363 ( .x(n3083), .a(n2022), .b(n3051), .c(n1374) );
    aoi21_1 U1364 ( .x(n3067), .a(n1197), .b(n1380), .c(n1364) );
    inv_2 U1365 ( .x(n1898), .a(N1976) );
    nand2i_2 U1366 ( .x(n3066), .a(n1898), .b(___cell__39620_net145508) );
    inv_2 U1367 ( .x(n1897), .a(N1810) );
    nand2i_2 U1368 ( .x(n3065), .a(n1897), .b(n1987) );
    nand2i_2 U1369 ( .x(n1367), .a(n1893), .b(n3624) );
    aoi21_1 U137 ( .x(n2231), .a(n1256), .b(n2130), .c(n2230) );
    inv_2 U1370 ( .x(n1893), .a(N2009) );
    inv_2 U1371 ( .x(n1896), .a(N1943) );
    nand2i_2 U1372 ( .x(n1366), .a(n1896), .b(n3662) );
    nor2i_1 U1373 ( .x(n1363), .a(N1744), .b(___cell__39620_net143710) );
    inv_2 U1374 ( .x(n1894), .a(N1645) );
    oai211_1 U1375 ( .x(n3062), .a(___cell__39620_net143872), .b(n1894), .c(
        n3061), .d(n3063) );
    inv_2 U1376 ( .x(___cell__39620_net144347), .a(___cell__39620_net144343)
         );
    aoi211_1 U1377 ( .x(n1365), .a(n1318), .b(n594), .c(n3062), .d(n1363) );
    inv_5 U1378 ( .x(n2011), .a(n2054) );
    nand2i_2 U1379 ( .x(n3163), .a(n1917), .b(n2837) );
    inv_8 U138 ( .x(n1686), .a(n1684) );
    inv_2 U1380 ( .x(n1917), .a(N317) );
    nand2i_2 U1381 ( .x(n3162), .a(n1588), .b(n2014) );
    aoai211_1 U1382 ( .x(n3158), .a(n1217), .b(n3159), .c(n1572), .d(n3155) );
    aoi21_1 U1383 ( .x(n3173), .a(n3174), .b(n1085), .c(n1415) );
    aoi221_1 U1384 ( .x(n3167), .a(n2022), .b(n3168), .c(n1267), .d(n2023), 
        .e(n1414) );
    nand2i_2 U1385 ( .x(n3164), .a(n1916), .b(n1064) );
    nand2i_2 U1386 ( .x(n3983), .a(n1918), .b(n977) );
    inv_2 U1387 ( .x(n1918), .a(N350) );
    aoi21_1 U1388 ( .x(n3153), .a(n1197), .b(n1054), .c(n1409) );
    inv_2 U1389 ( .x(n1922), .a(N1807) );
    nand2_2 U139 ( .x(n1712), .a(n1686), .b(___cell__39620_net144517) );
    nand2i_2 U1390 ( .x(n3154), .a(n1922), .b(n1987) );
    aoi22_1 U1391 ( .x(n3150), .a(n662), .b(n4141), .c(n1095), .d(n1992) );
    nand3_1 U1392 ( .x(n1413), .a(n3150), .b(n3154), .c(n3153) );
    nand2i_2 U1393 ( .x(n1412), .a(n1919), .b(n3624) );
    inv_2 U1394 ( .x(n1919), .a(N2006) );
    inv_2 U1395 ( .x(n1921), .a(N1940) );
    nand2i_2 U1396 ( .x(n1411), .a(n1921), .b(n3999) );
    ao21_3 U1397 ( .x(n3149), .a(n1318), .b(n1988), .c(n1408) );
    inv_2 U1398 ( .x(n1923), .a(N1973) );
    nand2i_2 U1399 ( .x(n3152), .a(n1923), .b(___cell__39620_net145508) );
    oai22_1 U140 ( .x(n2176), .a(n1584), .b(n1712), .c(n2177), .d(n1711) );
    aoi211_1 U1400 ( .x(n3148), .a(N1642), .b(n809), .c(n1407), .d(n1405) );
    inv_2 U1401 ( .x(n1920), .a(N1873) );
    nand2i_2 U1402 ( .x(n3151), .a(n1920), .b(n3998) );
    nand2i_2 U1403 ( .x(n2717), .a(n1658), .b(n3830) );
    nand2_2 U1404 ( .x(n2716), .a(n1085), .b(n3835) );
    nand2i_2 U1405 ( .x(n2704), .a(n1808), .b(n2837) );
    inv_2 U1406 ( .x(n1808), .a(N329) );
    inv_2 U1407 ( .x(n2699), .a(n3849) );
    nand2i_2 U1408 ( .x(n2702), .a(n1186), .b(n2574) );
    nor2i_3 U1409 ( .x(n2703), .a(n2709), .b(n2706) );
    aoi21_1 U141 ( .x(n2113), .a(n2070), .b(n583), .c(n1982) );
    nand2i_2 U1410 ( .x(n2685), .a(n1616), .b(n3839) );
    nand2i_2 U1411 ( .x(n2687), .a(n1815), .b(___cell__39620_net145508) );
    inv_2 U1412 ( .x(n1815), .a(N1985) );
    nand2i_2 U1413 ( .x(n2688), .a(n1814), .b(n735) );
    inv_2 U1414 ( .x(n1814), .a(N1852) );
    nand4i_1 U1415 ( .x(n2678), .a(n1240), .b(n2679), .c(n2680), .d(n2681) );
    inv_2 U1416 ( .x(n1810), .a(N2018) );
    nand2i_2 U1417 ( .x(n2684), .a(n1810), .b(n3624) );
    inv_2 U1418 ( .x(n1812), .a(N1885) );
    nand2i_2 U1419 ( .x(n2683), .a(n1812), .b(n944) );
    nand2_2 U142 ( .x(n2114), .a(n2115), .b(n2113) );
    and4i_3 U1420 ( .x(n1246), .a(n2678), .b(n2682), .c(n2683), .d(n2684) );
    inv_2 U1421 ( .x(n1813), .a(N1952) );
    nand2i_2 U1422 ( .x(n1245), .a(n1813), .b(n3999) );
    inv_2 U1423 ( .x(n1243), .a(N1819) );
    nor2_1 U1424 ( .x(n1242), .a(n1077), .b(n1243) );
    inv_2 U1425 ( .x(___cell__39620_net143785), .a(___cell__39620_net144350)
         );
    nand2i_2 U1426 ( .x(n2199), .a(n1588), .b(n2089) );
    aoi22_1 U1427 ( .x(n2196), .a(n650), .b(n2197), .c(n1221), .d(n2090) );
    aoi222_2 U1428 ( .x(n2191), .a(n649), .b(n2192), .c(n2193), .d(n2194), .e(
        n2139), .f(n2195) );
    nand4_1 U1429 ( .x(n2198), .a(n2191), .b(n2188), .c(n2196), .d(n2199) );
    inv_2 U143 ( .x(n664), .a(___cell__39620_net144326) );
    nand2i_2 U1430 ( .x(n2201), .a(n1703), .b(n977) );
    inv_2 U1431 ( .x(n1703), .a(N345) );
    and4i_3 U1432 ( .x(n2200), .a(n2209), .b(n2207), .c(n2202), .d(n2208) );
    nand2i_2 U1433 ( .x(n2207), .a(n670), .b(n3693) );
    inv_2 U1434 ( .x(n1705), .a(N1637) );
    nand2i_2 U1435 ( .x(n2170), .a(n1705), .b(n809) );
    inv_2 U1436 ( .x(n1706), .a(N1703) );
    nand2i_2 U1437 ( .x(n2169), .a(n1706), .b(___cell__39620_net145190) );
    aoi22_1 U1438 ( .x(n2166), .a(n1318), .b(n2167), .c(n1197), .d(n2168) );
    nand4_1 U1439 ( .x(n1129), .a(n2166), .b(n2164), .c(n2169), .d(n2170) );
    aoi21_1 U144 ( .x(n2069), .a(n2070), .b(n636), .c(n1982) );
    nand2i_2 U1440 ( .x(n1128), .a(n1704), .b(n3624) );
    inv_2 U1441 ( .x(n1704), .a(N2001) );
    inv_2 U1442 ( .x(n1708), .a(N1935) );
    nand2i_2 U1443 ( .x(n1127), .a(n1708), .b(n3662) );
    inv_2 U1444 ( .x(n1709), .a(N1968) );
    nand2i_2 U1445 ( .x(n2175), .a(n1709), .b(___cell__39620_net145508) );
    aoi22_1 U1446 ( .x(n2174), .a(N1802), .b(n1987), .c(N1835), .d(n4000) );
    inv_2 U1447 ( .x(n1707), .a(N1736) );
    nand2i_2 U1448 ( .x(n2173), .a(n1707), .b(___cell__39620_net145150) );
    aoi221_1 U1449 ( .x(n2862), .a(n1191), .b(n2863), .c(n1221), .d(n743), .e(
        n1297) );
    nand2i_0 U145 ( .x(n3706), .a(n1561), .b(n2070) );
    aoi22_1 U1450 ( .x(n2855), .a(n887), .b(n2856), .c(n502), .d(n2857) );
    inv_2 U1451 ( .x(n2861), .a(n1498) );
    inv_2 U1452 ( .x(n2860), .a(n1497) );
    aoi222_1 U1453 ( .x(n2858), .a(n649), .b(n2859), .c(n2193), .d(n2860), .e(
        n2139), .f(n2861) );
    aoi221_1 U1454 ( .x(n2871), .a(n2872), .b(n2022), .c(n842), .d(n2024), .e(
        n2869) );
    nand2i_2 U1456 ( .x(n2867), .a(n1844), .b(n2837) );
    inv_2 U1457 ( .x(n1844), .a(N326) );
    inv_2 U1458 ( .x(n1850), .a(N1982) );
    nand2i_2 U1459 ( .x(n2848), .a(n1850), .b(___cell__39620_net145508) );
    nand2i_2 U146 ( .x(n3707), .a(___cell__39620_net144317), .b(n1361) );
    aoi21_1 U1460 ( .x(n2845), .a(n1095), .b(n2846), .c(n1291) );
    inv_2 U1461 ( .x(n1848), .a(N1882) );
    nand2i_2 U1462 ( .x(n2847), .a(n1848), .b(n3998) );
    nand4_1 U1463 ( .x(n1296), .a(n2842), .b(n2847), .c(n2845), .d(n2848) );
    aoi221_1 U1464 ( .x(n1295), .a(n1197), .b(n2849), .c(N1849), .d(n735), .e(
        n1293) );
    inv_2 U1465 ( .x(n1849), .a(N1949) );
    nand2i_2 U1466 ( .x(n1294), .a(n1849), .b(n3999) );
    nand2i_2 U1467 ( .x(n2243), .a(n1574), .b(n2192) );
    aoi22_1 U1468 ( .x(n2241), .a(n1191), .b(n2197), .c(n1221), .d(n2089) );
    aoi221_1 U1469 ( .x(n2234), .a(n2211), .b(n2235), .c(n2212), .d(n750), .e(
        n1142) );
    inv_14 U147 ( .x(n940), .a(n938) );
    inv_2 U1470 ( .x(n2240), .a(n1468) );
    inv_2 U1471 ( .x(n2239), .a(n1467) );
    aoi222_1 U1472 ( .x(n2237), .a(n649), .b(n2238), .c(n2193), .d(n2239), .e(
        n2139), .f(n2240) );
    nand4_1 U1473 ( .x(n2242), .a(n2237), .b(n2234), .c(n2241), .d(n2243) );
    inv_2 U1474 ( .x(n1717), .a(N344) );
    nand2i_2 U1475 ( .x(n2244), .a(n1717), .b(n977) );
    inv_2 U1476 ( .x(n1718), .a(N1636) );
    nand2i_2 U1477 ( .x(n2221), .a(n1718), .b(n809) );
    aoi22_2 U1478 ( .x(n2219), .a(n1197), .b(n2165), .c(n662), .d(n2167) );
    nand2i_2 U1479 ( .x(n1140), .a(n1725), .b(n3624) );
    inv_5 U148 ( .x(n783), .a(Imm[0]) );
    inv_2 U1480 ( .x(n1725), .a(N2000) );
    inv_2 U1481 ( .x(n1721), .a(N1934) );
    nand2i_2 U1482 ( .x(n1139), .a(n1721), .b(n3999) );
    and4i_1 U1483 ( .x(n1138), .a(n2222), .b(n2223), .c(n2224), .d(n2225) );
    nand2i_2 U1484 ( .x(n2223), .a(n1722), .b(n1987) );
    inv_2 U1485 ( .x(n1722), .a(N1801) );
    nand2i_2 U1486 ( .x(n2224), .a(n1723), .b(n735) );
    inv_2 U1487 ( .x(n1723), .a(N1834) );
    nand2i_2 U1488 ( .x(n2225), .a(n1724), .b(___cell__39620_net145508) );
    inv_2 U1489 ( .x(n1724), .a(N1967) );
    nand2i_2 U149 ( .x(n3298), .a(n1579), .b(n928) );
    oai22_1 U1490 ( .x(n2222), .a(n947), .b(n1720), .c(
        ___cell__39620_net143710), .d(n1719) );
    inv_2 U1491 ( .x(n1720), .a(N1867) );
    inv_2 U1492 ( .x(n1719), .a(N1735) );
    nand2i_2 U1493 ( .x(n2909), .a(n1852), .b(n2837) );
    inv_2 U1494 ( .x(n1852), .a(N325) );
    inv_5 U1495 ( .x(n633), .a(n632) );
    and3i_2 U1496 ( .x(n2905), .a(n2908), .b(n2906), .c(n2907) );
    nand2i_2 U1499 ( .x(n2904), .a(n1574), .b(n2859) );
    inv_10 U150 ( .x(n863), .a(n862) );
    and4i_2 U1500 ( .x(n2883), .a(n1307), .b(n2884), .c(n2885), .d(n2886) );
    nand2i_2 U1501 ( .x(n2884), .a(n1856), .b(___cell__39620_net145508) );
    inv_2 U1502 ( .x(n1856), .a(N1981) );
    oai22_2 U1503 ( .x(n2880), .a(n2774), .b(n1182), .c(n865), .d(n1055) );
    nor2i_3 U1504 ( .x(n1304), .a(N1749), .b(___cell__39620_net143710) );
    inv_2 U1505 ( .x(n1319), .a(n2846) );
    aoi221_1 U1506 ( .x(n2882), .a(n1197), .b(n2846), .c(N1848), .d(n4000), 
        .e(n1305) );
    nor2i_1 U1507 ( .x(n1309), .a(N2014), .b(n1169) );
    and4i_4 U1508 ( .x(n2308), .a(___cell__39620_net143784), .b(n2311), .c(
        n2309), .d(n2310) );
    nand2_2 U151 ( .x(n3789), .a(n3478), .b(___cell__39620_net144331) );
    nand2i_4 U1510 ( .x(n3745), .a(n1736), .b(n944) );
    inv_2 U1511 ( .x(n821), .a(n1161) );
    inv_2 U1512 ( .x(n2328), .a(n3749) );
    aoi21_1 U1513 ( .x(n2327), .a(n1191), .b(n1728), .c(n2328) );
    nand2i_2 U1514 ( .x(n2331), .a(n703), .b(___cell__39620_net147270) );
    nand4i_1 U1515 ( .x(n2329), .a(n2330), .b(n2331), .c(n2332), .d(n2327) );
    aoi22_1 U1516 ( .x(n2317), .a(n535), .b(n2318), .c(
        ___cell__39620_net143864), .d(n2319) );
    aoi21_1 U1517 ( .x(n2323), .a(___cell__39620_net143722), .b(n2324), .c(
        n2320) );
    nand2i_2 U1518 ( .x(n2326), .a(n2300), .b(n3741) );
    inv_2 U1519 ( .x(___cell__39620_net145472), .a(___cell__39620_net144555)
         );
    aoi22_1 U152 ( .x(n706), .a(n710), .b(n709), .c(n708), .d(n707) );
    aoi22_1 U1520 ( .x(___cell__39620_net145470), .a(___cell__39620_net145450), 
        .b(n798), .c(___cell__39620_net145451), .d(___cell__39620_net145472)
         );
    inv_2 U1521 ( .x(n3776), .a(n1477) );
    nand2_2 U1522 ( .x(n2441), .a(n2193), .b(n3776) );
    nand2i_2 U1523 ( .x(n2440), .a(n1478), .b(n2139) );
    oai211_2 U1524 ( .x(n2438), .a(n2439), .b(n1658), .c(n2440), .d(n2441) );
    nand3i_2 U1525 ( .x(n2442), .a(n2443), .b(n2444), .c(n2445) );
    aoi21_1 U1526 ( .x(n2444), .a(n1221), .b(n2402), .c(n1190) );
    aoi22_1 U1527 ( .x(n2454), .a(reg_out_B[28]), .b(n1064), .c(Imm[28]), .d(
        ___cell__39620_net145617) );
    aoi21_1 U1528 ( .x(n2453), .a(n2457), .b(___cell__39620_net143864), .c(
        n1192) );
    nand2i_2 U1529 ( .x(n2452), .a(___cell__39620_net144406), .b(n2499) );
    nand2_5 U153 ( .x(n615), .a(N1662), .b(n616) );
    aoi22_1 U1530 ( .x(n2451), .a(n2022), .b(n2455), .c(n2024), .d(n2456) );
    nand2i_2 U1531 ( .x(n2420), .a(n588), .b(n663) );
    inv_2 U1532 ( .x(n1757), .a(N1726) );
    nand2i_2 U1533 ( .x(n2419), .a(n1757), .b(___cell__39620_net145190) );
    nor2i_1 U1534 ( .x(n1188), .a(N1759), .b(___cell__39620_net143710) );
    nand4i_1 U1535 ( .x(n2418), .a(n1188), .b(n2419), .c(n2420), .d(n2421) );
    inv_2 U1536 ( .x(n1755), .a(N2024) );
    nand2i_2 U1537 ( .x(n2417), .a(n1755), .b(n3624) );
    inv_2 U1538 ( .x(n1756), .a(N1660) );
    nand2i_2 U1539 ( .x(n2416), .a(n1756), .b(n809) );
    inv_2 U154 ( .x(n3269), .a(n1472) );
    nand2i_2 U1540 ( .x(n2415), .a(n2412), .b(___cell__39620_net145285) );
    nand2i_2 U1541 ( .x(n2414), .a(n1182), .b(n3727) );
    nand4_1 U1542 ( .x(n2413), .a(n2414), .b(n2415), .c(n2416), .d(n2417) );
    inv_2 U1543 ( .x(n1758), .a(N1958) );
    nand2i_4 U1544 ( .x(n2427), .a(n1758), .b(n3662) );
    inv_2 U1545 ( .x(n1759), .a(N1825) );
    aoi22_1 U1547 ( .x(n2057), .a(n1267), .b(n2059), .c(n2024), .d(n2027) );
    nand2i_1 U1548 ( .x(n2052), .a(n1566), .b(n2090) );
    inv_5 U1549 ( .x(n3614), .a(n3613) );
    exnor2_1 U155 ( .x(n1472), .a(reg_out_A[30]), .b(reg_out_B[30]) );
    oai211_1 U1550 ( .x(n2051), .a(n2012), .b(n1574), .c(n2052), .d(n2049) );
    inv_2 U1551 ( .x(n1670), .a(N1971) );
    nand2i_2 U1552 ( .x(n2042), .a(n1670), .b(___cell__39620_net145508) );
    aoi21_2 U1553 ( .x(n2039), .a(n662), .b(n1054), .c(n1076) );
    inv_2 U1554 ( .x(n1669), .a(N1838) );
    nand2i_2 U1555 ( .x(n2041), .a(n1669), .b(n735) );
    aoi22_1 U1556 ( .x(n2040), .a(n1197), .b(n1993), .c(n1095), .d(n2043) );
    inv_2 U1557 ( .x(n1666), .a(N2004) );
    nand2i_2 U1558 ( .x(n2038), .a(n1666), .b(n3624) );
    aoi211_1 U1559 ( .x(n2035), .a(N1640), .b(n809), .c(n1075), .d(n1073) );
    exnor2_1 U156 ( .x(n1471), .a(reg_out_A[30]), .b(Imm[30]) );
    inv_2 U1560 ( .x(n1667), .a(N1871) );
    nand2i_2 U1561 ( .x(n2037), .a(n1667), .b(n944) );
    aoi22_1 U1562 ( .x(n2036), .a(N1739), .b(___cell__39620_net145150), .c(
        n1318), .d(n1992) );
    nand4_1 U1563 ( .x(n1080), .a(n2036), .b(n2037), .c(n2035), .d(n2038) );
    inv_2 U1564 ( .x(n1668), .a(N1938) );
    nand2i_2 U1565 ( .x(n1079), .a(n1668), .b(n3999) );
    inv_2 U1566 ( .x(n2400), .a(n578) );
    aoi221_1 U1567 ( .x(n2395), .a(n649), .b(n2399), .c(n650), .d(n2400), .e(
        n2396) );
    nand2i_2 U1568 ( .x(n2394), .a(n702), .b(n2324) );
    inv_2 U1569 ( .x(n2393), .a(n2319) );
    nand2i_2 U157 ( .x(n3775), .a(n1752), .b(n1063) );
    inv_2 U1571 ( .x(n3740), .a(n2402) );
    nand4i_1 U1572 ( .x(n2403), .a(n2405), .b(n2407), .c(n2408), .d(n2409) );
    aoi211_1 U1573 ( .x(n2401), .a(n1191), .b(n2402), .c(n2403), .d(n1185) );
    inv_7 U1574 ( .x(n3724), .a(n3723) );
    nand2i_2 U1576 ( .x(n2404), .a(n784), .b(n3765) );
    oai21_2 U1577 ( .x(n2391), .a(n816), .b(n3720), .c(n2372) );
    inv_2 U1578 ( .x(n3767), .a(n3766) );
    nand2i_2 U1579 ( .x(n2390), .a(n3767), .b(n1217) );
    inv_2 U158 ( .x(n2185), .a(n1715) );
    aoi22_1 U1580 ( .x(n2389), .a(n539), .b(n2390), .c(
        ___cell__39620_net143722), .d(n2391) );
    nand4_1 U1581 ( .x(n2377), .a(n2378), .b(n2379), .c(n2380), .d(n2381) );
    nand2i_2 U1582 ( .x(n2378), .a(n1055), .b(n3727) );
    nand2i_2 U1583 ( .x(n2379), .a(n2376), .b(___cell__39620_net147791) );
    nand2i_2 U1584 ( .x(n2381), .a(n1750), .b(n3624) );
    inv_2 U1585 ( .x(n1750), .a(N2025) );
    aoi221_1 U1587 ( .x(n2383), .a(n1197), .b(n2384), .c(N1992), .d(
        ___cell__39620_net145508), .e(n1181) );
    aoi21_1 U1588 ( .x(n791), .a(n535), .b(___cell__39620_net145444), .c(n782)
         );
    inv_7 U1589 ( .x(n3720), .a(n3719) );
    inv_2 U1590 ( .x(n792), .a(___cell__39620_net147270) );
    inv_2 U1591 ( .x(n798), .a(n794) );
    nand2_2 U1592 ( .x(___cell__39620_net145428), .a(n2288), .b(n2289) );
    inv_2 U1593 ( .x(n1727), .a(N1961) );
    inv_2 U1594 ( .x(___cell__39620_net144355), .a(___cell__39620_net143653)
         );
    inv_5 U1595 ( .x(___cell__39620_net143872), .a(n809) );
    inv_4 U1596 ( .x(n1726), .a(N2027) );
    oai21_1 U1597 ( .x(n2293), .a(n1153), .b(n1658), .c(n2294) );
    inv_2 U1598 ( .x(n678), .a(n1662) );
    nand3_3 U1599 ( .x(n1087), .a(n678), .b(n1663), .c(n701) );
    oai22_1 U160 ( .x(n2428), .a(n1529), .b(n1715), .c(n2429), .d(n1713) );
    nand4i_1 U1600 ( .x(n3988), .a(n1424), .b(n3190), .c(n3987), .d(n3192) );
    nor2i_1 U1601 ( .x(n1424), .a(N1997), .b(n1169) );
    nand2i_2 U1602 ( .x(n3987), .a(___cell__39620_net144343), .b(n3245) );
    inv_2 U1603 ( .x(n1426), .a(n1517) );
    nor2i_1 U1604 ( .x(n1425), .a(n1426), .b(n690) );
    ao21_2 U1605 ( .x(n3207), .a(n2024), .b(n2826), .c(n1425) );
    nand2i_2 U1606 ( .x(n3209), .a(n1518), .b(n2139) );
    nand2i_3 U1607 ( .x(n3206), .a(n1626), .b(n2827) );
    aoai211_1 U1608 ( .x(n3205), .a(n917), .b(n530), .c(n1064), .d(n816) );
    nand2i_0 U1609 ( .x(n3180), .a(___cell__39620_net144175), .b(n1545) );
    inv_5 U161 ( .x(n938), .a(reg_out_A[2]) );
    nand2i_2 U1610 ( .x(n3989), .a(n1924), .b(n2837) );
    inv_2 U1611 ( .x(n1924), .a(N308) );
    inv_5 U1612 ( .x(n1437), .a(n3219) );
    inv_5 U1613 ( .x(n3216), .a(n1733) );
    oai211_1 U1614 ( .x(n3215), .a(n3216), .b(n1657), .c(n3217), .d(n3218) );
    inv_5 U1615 ( .x(n941), .a(reg_out_A[0]) );
    aoi222_1 U1616 ( .x(n3212), .a(n502), .b(n3214), .c(n942), .d(
        ___cell__39620_net145444), .e(N341), .f(n977) );
    inv_5 U1617 ( .x(n3611), .a(n3610) );
    inv_5 U1618 ( .x(n2012), .a(n2093) );
    nand2i_2 U1619 ( .x(n2016), .a(n1594), .b(n2837) );
    exnor2_1 U162 ( .x(n1475), .a(reg_out_A[29]), .b(Imm[29]) );
    inv_2 U1620 ( .x(n1594), .a(N316) );
    aoi21_1 U1622 ( .x(n2013), .a(n1221), .b(n2014), .c(n2007) );
    inv_2 U1623 ( .x(n3623), .a(n3622) );
    inv_5 U1624 ( .x(n3620), .a(n3619) );
    oai211_1 U1625 ( .x(n2007), .a(n1062), .b(n1532), .c(n2008), .d(n2009) );
    aoi22_1 U1626 ( .x(n2026), .a(n502), .b(n2027), .c(
        ___cell__39620_net143722), .d(n2028) );
    inv_2 U1627 ( .x(n2025), .a(n720) );
    aoi22_1 U1628 ( .x(n2021), .a(n2022), .b(n2023), .c(n2024), .d(n2025) );
    nand3_1 U1629 ( .x(n2020), .a(n2021), .b(n2029), .c(n2026) );
    inv_2 U163 ( .x(n3266), .a(n1476) );
    nand2i_2 U1630 ( .x(n2019), .a(n1598), .b(n977) );
    inv_2 U1631 ( .x(n1598), .a(N349) );
    nand2i_2 U1633 ( .x(n2033), .a(n1658), .b(n3172) );
    inv_2 U1634 ( .x(n1615), .a(N1839) );
    nand2i_2 U1635 ( .x(n1991), .a(n1615), .b(n4000) );
    aoi22_1 U1636 ( .x(n1986), .a(N1806), .b(n1987), .c(n662), .d(n1988) );
    inv_2 U1637 ( .x(n1617), .a(N1972) );
    nand2i_2 U1638 ( .x(n1990), .a(n1617), .b(___cell__39620_net145508) );
    aoi22_1 U1639 ( .x(n1989), .a(n1197), .b(n1992), .c(n1095), .d(n1993) );
    nand2_5 U164 ( .x(n1089), .a(n713), .b(n927) );
    nand2i_2 U1640 ( .x(n1058), .a(n1599), .b(n3624) );
    inv_2 U1641 ( .x(n1599), .a(N2005) );
    inv_2 U1642 ( .x(n1613), .a(N1939) );
    nand2i_2 U1643 ( .x(n1057), .a(n1613), .b(n3662) );
    and4i_3 U1644 ( .x(n1056), .a(n1053), .b(n1984), .c(n1985), .d(n1983) );
    nand2i_2 U1645 ( .x(n1984), .a(n1600), .b(___cell__39620_net145150) );
    inv_2 U1646 ( .x(n1600), .a(N1740) );
    nand2i_2 U1647 ( .x(n1985), .a(n1601), .b(n3998) );
    inv_2 U1648 ( .x(n1601), .a(N1872) );
    aoi211_1 U1649 ( .x(n1983), .a(N1641), .b(n809), .c(n1052), .d(n1050) );
    nand2i_1 U165 ( .x(___cell__39620_net144555), .a(n498), .b(n1728) );
    aoi22_1 U1650 ( .x(n3011), .a(n502), .b(n3012), .c(
        ___cell__39620_net143722), .d(n3013) );
    aoi21_1 U1651 ( .x(n3003), .a(n1191), .b(n3004), .c(
        ___cell__39620_net143982) );
    aoi22_1 U1652 ( .x(n2999), .a(n649), .b(n3000), .c(n650), .d(n3001) );
    aoi21_1 U1653 ( .x(n3002), .a(n1221), .b(n2899), .c(n2996) );
    inv_2 U1654 ( .x(n1876), .a(N355) );
    nand2i_2 U1655 ( .x(n3006), .a(n1876), .b(n977) );
    nand2i_4 U1656 ( .x(n2987), .a(n1881), .b(n735) );
    aoi21_1 U1657 ( .x(n2985), .a(n662), .b(n1308), .c(n1340) );
    inv_4 U1658 ( .x(n1882), .a(N1978) );
    nand2i_4 U1659 ( .x(n2986), .a(n1882), .b(___cell__39620_net145508) );
    nand2i_2 U166 ( .x(n3761), .a(n1635), .b(___cell__39620_net145472) );
    nand2i_2 U1660 ( .x(n1344), .a(n1877), .b(n3624) );
    inv_2 U1661 ( .x(n1877), .a(N2011) );
    inv_2 U1662 ( .x(n1880), .a(N1945) );
    nand2i_2 U1663 ( .x(n1343), .a(n1880), .b(n3662) );
    inv_2 U1664 ( .x(n1879), .a(N1878) );
    inv_2 U1665 ( .x(n1878), .a(N1746) );
    nand2i_2 U1666 ( .x(n2983), .a(n1878), .b(___cell__39620_net145150) );
    aoi211_1 U1667 ( .x(n2982), .a(N1647), .b(n809), .c(n1337), .d(n1335) );
    inv_2 U1668 ( .x(n1868), .a(N356) );
    aoi21_1 U1669 ( .x(n2965), .a(n1191), .b(n2899), .c(n1327) );
    nand2i_2 U167 ( .x(___cell__39620_net147350), .a(n718), .b(n798) );
    nand2i_2 U1670 ( .x(n2970), .a(n1867), .b(n2837) );
    inv_2 U1671 ( .x(n1867), .a(N323) );
    nand2i_2 U1672 ( .x(n2963), .a(n1574), .b(n3004) );
    and3i_1 U1673 ( .x(n2962), .a(n2961), .b(n2963), .c(n2964) );
    inv_2 U1674 ( .x(n1871), .a(N1946) );
    nand2i_2 U1675 ( .x(n3938), .a(n1871), .b(n3662) );
    inv_2 U1676 ( .x(n1873), .a(N2012) );
    nand2i_2 U1677 ( .x(n3939), .a(n1873), .b(n3624) );
    nand4_1 U1678 ( .x(n2954), .a(n2955), .b(n2956), .c(n2957), .d(n2953) );
    nand4i_1 U1679 ( .x(n3940), .a(n2954), .b(n2950), .c(n3939), .d(n3938) );
    or2_1 U168 ( .x(n498), .a(reg_out_B[4]), .b(reg_out_B[3]) );
    nand4i_1 U1680 ( .x(n3912), .a(n2920), .b(n2918), .c(n3910), .d(n3911) );
    nand4_1 U1681 ( .x(n2920), .a(n2921), .b(n2922), .c(n2923), .d(n2924) );
    nand2i_2 U1682 ( .x(n3910), .a(n1863), .b(n3999) );
    inv_2 U1683 ( .x(n1863), .a(N1947) );
    nand2i_2 U1684 ( .x(n3911), .a(n1865), .b(n3624) );
    inv_2 U1685 ( .x(n1865), .a(N2013) );
    nand3i_1 U1686 ( .x(n2931), .a(n2932), .b(n2933), .c(n2934) );
    nand2i_2 U1687 ( .x(n2947), .a(n1857), .b(n2837) );
    inv_2 U1688 ( .x(n1857), .a(N324) );
    nand2i_2 U1689 ( .x(n2946), .a(n1858), .b(n977) );
    inv_5 U169 ( .x(___cell__39620_net144707), .a(Imm[24]) );
    inv_2 U1690 ( .x(n1858), .a(N357) );
    nand2i_2 U1691 ( .x(n2752), .a(n1817), .b(n2837) );
    inv_2 U1692 ( .x(n1817), .a(N328) );
    nor3i_2 U1693 ( .x(n2749), .a(n2747), .b(n2748), .c(n2745) );
    inv_2 U1694 ( .x(n1816), .a(n567) );
    ao22_3 U1695 ( .x(n2759), .a(n757), .b(n2803), .c(n3854), .d(n758) );
    nand2i_2 U1696 ( .x(n2761), .a(n4001), .b(n2714) );
    and3i_3 U1697 ( .x(n2750), .a(n2759), .b(n2760), .c(n2761) );
    nand4i_2 U1698 ( .x(n2724), .a(n2723), .b(n2725), .c(n2726), .d(n2727) );
    inv_2 U1699 ( .x(n1821), .a(N1884) );
    inv_5 U170 ( .x(n648), .a(Imm[29]) );
    nand2i_2 U1700 ( .x(n2736), .a(n1821), .b(n3997) );
    aoi21_1 U1701 ( .x(n2732), .a(n1197), .b(n2733), .c(n1253) );
    inv_2 U1702 ( .x(n1818), .a(N1653) );
    nand2i_2 U1703 ( .x(n2735), .a(n1818), .b(n809) );
    and4i_3 U1704 ( .x(n2734), .a(n2724), .b(n2735), .c(n2732), .d(n2736) );
    nand2i_4 U1705 ( .x(n2731), .a(n1822), .b(n3662) );
    inv_2 U1706 ( .x(n1823), .a(N1818) );
    nand2i_2 U1707 ( .x(n2730), .a(n1823), .b(n1987) );
    nand4i_1 U1708 ( .x(n2728), .a(n1251), .b(n2729), .c(n2730), .d(n2731) );
    nor2i_1 U1709 ( .x(n1252), .a(N2017), .b(n1169) );
    exnor2_1 U171 ( .x(n1470), .a(reg_out_A[31]), .b(n4144) );
    inv_2 U1710 ( .x(n2668), .a(n3835) );
    inv_5 U1711 ( .x(n3553), .a(n3552) );
    nand2i_2 U1712 ( .x(n2671), .a(n4030), .b(n3057) );
    nand4_1 U1713 ( .x(n2624), .a(n3825), .b(n3824), .c(n3823), .d(n3822) );
    aoi22_1 U1714 ( .x(n2660), .a(n829), .b(___cell__39620_net145617), .c(
        n2661), .d(n2024) );
    nand2_2 U1715 ( .x(n2663), .a(n2707), .b(n502) );
    nand4_1 U1716 ( .x(n2662), .a(n2663), .b(n2664), .c(n2660), .d(n2665) );
    buf_10 U1717 ( .x(n636), .a(reg_out_A[23]) );
    inv_2 U1718 ( .x(n3841), .a(n3840) );
    inv_2 U1719 ( .x(n2652), .a(n1488) );
    nor2i_1 U172 ( .x(n1149), .a(n1150), .b(n509) );
    inv_2 U1720 ( .x(n2651), .a(n1487) );
    aoi22_1 U1721 ( .x(n2650), .a(n2139), .b(n2651), .c(n2193), .d(n2652) );
    oai211_3 U1722 ( .x(n3837), .a(n747), .b(n1565), .c(n3836), .d(n2628) );
    inv_5 U1723 ( .x(n2655), .a(n3837) );
    oai211_1 U1724 ( .x(n2654), .a(n2655), .b(n1566), .c(n2650), .d(n2656) );
    nand2i_2 U1725 ( .x(n2659), .a(n1798), .b(n2837) );
    inv_2 U1726 ( .x(n1798), .a(N330) );
    nand2i_2 U1727 ( .x(n3842), .a(n1797), .b(n1064) );
    inv_2 U1728 ( .x(n2658), .a(n3842) );
    oai221_4 U1729 ( .x(n2574), .a(n3419), .b(n1070), .c(n1313), .d(n1565), 
        .e(n1807) );
    nand2_1 U173 ( .x(n3401), .a(n1691), .b(n901) );
    aoi21_1 U1730 ( .x(n2657), .a(n1191), .b(n2574), .c(n2658) );
    inv_2 U1731 ( .x(n1800), .a(N2019) );
    nand2i_2 U1732 ( .x(n2642), .a(n1800), .b(n3624) );
    inv_2 U1733 ( .x(n1803), .a(N1886) );
    nand2i_2 U1734 ( .x(n2641), .a(n1803), .b(n3998) );
    inv_2 U1735 ( .x(n1802), .a(N1721) );
    nand2i_2 U1736 ( .x(n2640), .a(n1802), .b(___cell__39620_net145190) );
    and4i_1 U1737 ( .x(n1239), .a(n2636), .b(n2640), .c(n2641), .d(n2642) );
    nand2i_2 U1738 ( .x(n2647), .a(n1804), .b(n3999) );
    aoi211_1 U1739 ( .x(n2646), .a(n1197), .b(n2600), .c(n1237), .d(n1236) );
    nand2i_3 U174 ( .x(n3729), .a(n1564), .b(n3591) );
    nand2i_2 U1740 ( .x(n2627), .a(n1658), .b(n3812) );
    nand2_2 U1741 ( .x(n2626), .a(n1085), .b(n3816) );
    nand2i_2 U1742 ( .x(n2625), .a(n4031), .b(n3057) );
    nand4_1 U1743 ( .x(n2618), .a(n2625), .b(n2626), .c(n2623), .d(n2627) );
    inv_2 U1744 ( .x(n1791), .a(N364) );
    nand2i_2 U1745 ( .x(n2617), .a(n1791), .b(n977) );
    inv_5 U1746 ( .x(n2611), .a(n3422) );
    inv_2 U1747 ( .x(n1790), .a(N331) );
    nand2i_2 U1748 ( .x(n3827), .a(n1790), .b(n2837) );
    inv_2 U1749 ( .x(n2615), .a(n3827) );
    aoi22_1 U175 ( .x(n2269), .a(n1971), .b(n2270), .c(n1177), .d(n2271) );
    inv_2 U1750 ( .x(n2613), .a(n3828) );
    nor3i_2 U1751 ( .x(n2614), .a(n2612), .b(n2615), .c(n2610) );
    nand2_2 U1752 ( .x(n2621), .a(n2661), .b(n502) );
    and4i_3 U1753 ( .x(n1232), .a(n2598), .b(n2596), .c(n2592), .d(n2597) );
    nand2i_2 U1754 ( .x(n2596), .a(n1796), .b(___cell__39620_net145508) );
    inv_2 U1755 ( .x(n1796), .a(N1987) );
    and4i_3 U1756 ( .x(n2592), .a(n2589), .b(n2593), .c(n2594), .d(n2595) );
    nand2i_2 U1757 ( .x(n1231), .a(n1792), .b(n3624) );
    inv_2 U1758 ( .x(n1792), .a(N2020) );
    nand2i_2 U1759 ( .x(n2559), .a(n1788), .b(n3999) );
    inv_3 U176 ( .x(n3462), .a(n2265) );
    aoi221_1 U1760 ( .x(n2555), .a(n1318), .b(n2473), .c(n662), .d(n2423), .e(
        n1213) );
    nor2i_3 U1761 ( .x(n1215), .a(N1988), .b(___cell__39620_net143845) );
    nand4i_1 U1762 ( .x(n2558), .a(n1215), .b(n2555), .c(n2556), .d(n2559) );
    inv_2 U1763 ( .x(n1784), .a(N2021) );
    nand2i_2 U1764 ( .x(n2554), .a(n1784), .b(n3624) );
    inv_2 U1765 ( .x(n1787), .a(N1888) );
    nand2i_2 U1766 ( .x(n2553), .a(n1787), .b(n944) );
    inv_2 U1767 ( .x(n1786), .a(N1723) );
    nand2i_2 U1768 ( .x(n2552), .a(n1786), .b(___cell__39620_net145190) );
    inv_2 U1769 ( .x(n2550), .a(n3819) );
    nand2i_2 U177 ( .x(n2265), .a(n3492), .b(n3493) );
    and4i_1 U1770 ( .x(n2547), .a(n2550), .b(n2548), .c(n2549), .d(n2546) );
    nand4_1 U1771 ( .x(n2551), .a(n2547), .b(n2552), .c(n2553), .d(n2554) );
    nand2i_2 U1772 ( .x(n1454), .a(n1060), .b(n1591) );
    nand2i_2 U1773 ( .x(n2587), .a(n784), .b(n3812) );
    inv_2 U1774 ( .x(n2586), .a(n3816) );
    oai211_2 U1775 ( .x(n2579), .a(n2586), .b(___cell__39620_net144406), .c(
        n2580), .d(n2587) );
    aoi22_1 U1776 ( .x(n2573), .a(n649), .b(n2574), .c(n650), .d(n2532) );
    aoi21_1 U1777 ( .x(n2567), .a(n2544), .b(n2568), .c(n1216) );
    nor2i_3 U1778 ( .x(n1223), .a(n1204), .b(n1224) );
    nand2i_2 U1779 ( .x(n2585), .a(n4032), .b(n3057) );
    aoi22_1 U178 ( .x(n2264), .a(n2079), .b(n2265), .c(n2266), .d(n608) );
    nand2i_2 U1780 ( .x(n2542), .a(n4001), .b(n3782) );
    nand2i_2 U1781 ( .x(n2541), .a(n4033), .b(n3057) );
    inv_2 U1782 ( .x(n2540), .a(n3785) );
    oai211_1 U1783 ( .x(n2538), .a(n2540), .b(n702), .c(n2541), .d(n2542) );
    nand2i_2 U1784 ( .x(n2537), .a(n1772), .b(n2837) );
    inv_2 U1785 ( .x(n1710), .a(n1447) );
    aoi22_1 U1786 ( .x(n2536), .a(reg_out_B[26]), .b(n1064), .c(Imm[26]), .d(
        ___cell__39620_net145617) );
    nor2i_3 U1787 ( .x(n1210), .a(___cell__39620_net143722), .b(n1211) );
    inv_2 U1788 ( .x(n1591), .a(n1590) );
    nand2i_2 U1789 ( .x(n1595), .a(n1534), .b(n1591) );
    inv_2 U1790 ( .x(n1597), .a(n1595) );
    inv_2 U1791 ( .x(n3805), .a(n3804) );
    inv_2 U1792 ( .x(n3807), .a(n3806) );
    aoai211_1 U1793 ( .x(n2529), .a(n502), .b(n2568), .c(n3807), .d(n1451) );
    inv_4 U1794 ( .x(n3809), .a(n3808) );
    inv_2 U1795 ( .x(n2524), .a(n2489) );
    oai211_1 U1796 ( .x(n2523), .a(n2524), .b(n1580), .c(n2525), .d(n2526) );
    nand4i_3 U1797 ( .x(n2527), .a(n2523), .b(n2528), .c(n2529), .d(n2530) );
    inv_2 U1798 ( .x(n3420), .a(n2673) );
    aoi22_1 U1799 ( .x(n2531), .a(n539), .b(n2490), .c(n649), .d(n2532) );
    nand2i_2 U180 ( .x(n2263), .a(n1625), .b(n2302) );
    inv_2 U1800 ( .x(n3423), .a(n3739) );
    nand2i_2 U1801 ( .x(n2534), .a(n1574), .b(n3422) );
    inv_8 U1802 ( .x(n3418), .a(n2763) );
    aoi22_1 U1803 ( .x(n2533), .a(n1221), .b(n2399), .c(n1191), .d(n2492) );
    inv_8 U1804 ( .x(n1520), .a(n1519) );
    nand3_1 U1805 ( .x(n1184), .a(n1520), .b(n810), .c(n1612) );
    nor2i_1 U1806 ( .x(n1209), .a(N1956), .b(n1184) );
    inv_2 U1807 ( .x(n1774), .a(N2022) );
    nand2i_2 U1808 ( .x(n2511), .a(n1774), .b(n3624) );
    inv_2 U1809 ( .x(n1777), .a(N1889) );
    nand2i_2 U181 ( .x(n3734), .a(n1564), .b(n3594) );
    nand2i_2 U1810 ( .x(n2510), .a(n1777), .b(n3998) );
    inv_4 U1811 ( .x(n1776), .a(N1724) );
    nand2i_3 U1812 ( .x(n2509), .a(n1776), .b(___cell__39620_net145190) );
    inv_2 U1813 ( .x(n2507), .a(n3803) );
    nand2i_2 U1814 ( .x(n2515), .a(n1616), .b(n2473) );
    inv_2 U1815 ( .x(n1779), .a(N1989) );
    nand2i_2 U1816 ( .x(n2517), .a(n1780), .b(n4000) );
    nor2i_1 U1817 ( .x(___cell__39620_net144312), .a(___cell__39620_net144166), 
        .b(n805) );
    aoi211_1 U1818 ( .x(n1005), .a(n977), .b(N343), .c(n2364), .d(n2354) );
    oai211_1 U1819 ( .x(n4052), .a(n1004), .b(___cell__39620_net147731), .c(
        n1005), .d(n1006) );
    nor2i_3 U182 ( .x(n1151), .a(n1147), .b(n1152) );
    aoi221_1 U1820 ( .x(n953), .a(N309), .b(n2837), .c(N342), .d(n977), .e(
        n2834) );
    ao21_2 U1821 ( .x(n4055), .a(___cell__39620_net143326), .b(n999), .c(n1000
        ) );
    inv_2 U1822 ( .x(n1899), .a(N319) );
    nand2i_2 U1823 ( .x(n968), .a(n1899), .b(n2837) );
    inv_2 U1824 ( .x(n1674), .a(N314) );
    nand2i_2 U1825 ( .x(n959), .a(n1674), .b(n2837) );
    and4i_3 U1826 ( .x(n989), .a(n2497), .b(n2495), .c(n2493), .d(n2496) );
    inv_2 U1827 ( .x(n1762), .a(N367) );
    nand2i_2 U1828 ( .x(n988), .a(n1762), .b(n977) );
    nand2i_2 U1829 ( .x(n1456), .a(n4018), .b(n3057) );
    oai21_1 U183 ( .x(n2259), .a(n1529), .b(n1281), .c(n2260) );
    and4i_1 U1830 ( .x(n1036), .a(n3129), .b(n3132), .c(n3133), .d(n3134) );
    inv_2 U1831 ( .x(n1825), .a(N360) );
    nand2i_2 U1832 ( .x(n1022), .a(n1825), .b(n977) );
    and4i_3 U1833 ( .x(n1021), .a(n2795), .b(n2793), .c(n2792), .d(n2794) );
    and4i_2 U1834 ( .x(n1020), .a(n1265), .b(n1262), .c(n1263), .d(n1264) );
    inv_2 U1836 ( .x(n1883), .a(N321) );
    nand2i_2 U1837 ( .x(n971), .a(n1883), .b(n2837) );
    inv_2 U1838 ( .x(n1891), .a(N320) );
    nand2i_2 U1839 ( .x(n1032), .a(n1891), .b(n2837) );
    nor2_0 U184 ( .x(n1938), .a(IR_function_field[4]), .b(IR_function_field[1]
        ) );
    and4i_1 U1840 ( .x(n965), .a(n3160), .b(n3161), .c(n3162), .d(n3163) );
    inv_2 U1841 ( .x(n1809), .a(N362) );
    nand2i_2 U1842 ( .x(n1019), .a(n1809), .b(n977) );
    and4i_3 U1843 ( .x(n1018), .a(n2705), .b(n2703), .c(n2700), .d(n2704) );
    and4i_2 U1844 ( .x(n1017), .a(n1247), .b(n1244), .c(n1245), .d(n1246) );
    inv_2 U1845 ( .x(n1702), .a(N312) );
    nand2i_2 U1846 ( .x(n956), .a(n1702), .b(n2837) );
    and4i_2 U1847 ( .x(n954), .a(n1129), .b(n1126), .c(n1127), .d(n1128) );
    inv_2 U1848 ( .x(n1845), .a(N359) );
    nand2i_2 U1849 ( .x(n1025), .a(n1845), .b(n977) );
    inv_4 U185 ( .x(n3861), .a(n1834) );
    nor3i_2 U1850 ( .x(n1024), .a(n2867), .b(n2868), .c(n2865) );
    and3i_2 U1851 ( .x(n1023), .a(n1296), .b(n1294), .c(n1295) );
    inv_2 U1852 ( .x(n1716), .a(N311) );
    nand2i_2 U1853 ( .x(n1003), .a(n1716), .b(n2837) );
    oai211_1 U1854 ( .x(n4053), .a(n1001), .b(___cell__39620_net143287), .c(
        n1002), .d(n1003) );
    inv_2 U1855 ( .x(n1853), .a(N358) );
    nand2i_2 U1856 ( .x(n3891), .a(n1853), .b(n977) );
    inv_2 U1857 ( .x(n976), .a(n3891) );
    nand4_1 U1858 ( .x(n975), .a(n2905), .b(n2896), .c(n2903), .d(n2909) );
    inv_2 U1860 ( .x(n859), .a(n2329) );
    inv_2 U1861 ( .x(n1753), .a(N335) );
    nand2i_2 U1862 ( .x(n1007), .a(n1753), .b(n2837) );
    inv_2 U1863 ( .x(n1754), .a(N368) );
    nand2i_4 U1864 ( .x(n1009), .a(n1754), .b(n977) );
    inv_2 U1866 ( .x(n1665), .a(N315) );
    nand2i_2 U1867 ( .x(n997), .a(n1665), .b(n2837) );
    nor3i_1 U1868 ( .x(n996), .a(n1079), .b(n1080), .c(n1081) );
    oai31_2 U1869 ( .x(n993), .a(n2387), .b(n2377), .c(n2382), .d(
        ___cell__39620_net147732) );
    oaoi211_1 U187 ( .x(n1416), .a(n1417), .b(n1418), .c(n665), .d(
        ___cell__39620_net144062) );
    nand2i_2 U1870 ( .x(n991), .a(n1748), .b(n2837) );
    inv_2 U1871 ( .x(n1748), .a(N336) );
    nand3i_1 U1872 ( .x(n1942), .a(IR_opcode_field[0]), .b(n1533), .c(
        ___cell__39620_net143655) );
    inv_2 U1873 ( .x(n3211), .a(n3989) );
    nand3i_1 U1874 ( .x(n948), .a(n3211), .b(n3212), .c(n3213) );
    inv_2 U1875 ( .x(n1875), .a(N322) );
    nand2i_2 U1876 ( .x(n1030), .a(n1875), .b(n2837) );
    nand2i_2 U1877 ( .x(n972), .a(___cell__39620_net143287), .b(n3940) );
    and4i_4 U1878 ( .x(n1026), .a(n2937), .b(n2940), .c(n2946), .d(n2947) );
    nand2i_2 U1879 ( .x(n1027), .a(___cell__39620_net147731), .b(n3912) );
    inv_2 U188 ( .x(n1421), .a(N1864) );
    or3i_2 U1880 ( .x(n978), .a(n2734), .b(n1252), .c(n2728) );
    inv_8 U1881 ( .x(n807), .a(n806) );
    inv_2 U1882 ( .x(n1799), .a(N363) );
    nand2i_2 U1883 ( .x(n981), .a(n1799), .b(n977) );
    oai21_1 U1884 ( .x(n986), .a(n2551), .b(n2558), .c(
        ___cell__39620_net143326) );
    inv_2 U1885 ( .x(n1783), .a(N365) );
    nand2i_2 U1886 ( .x(n985), .a(n1783), .b(n977) );
    inv_2 U1887 ( .x(n1782), .a(N332) );
    nand2i_2 U1888 ( .x(n984), .a(n1782), .b(n2837) );
    nand2i_2 U1889 ( .x(n1013), .a(n1773), .b(n977) );
    nor2_1 U189 ( .x(n1420), .a(n947), .b(n1421) );
    inv_2 U1890 ( .x(n1773), .a(N366) );
    inv_2 U1891 ( .x(n1533), .a(n733) );
    aoi21_1 U1892 ( .x(n4117), .a(n3997), .b(n945), .c(___cell__6067_net21981)
         );
    nor2i_1 U1893 ( .x(N3297), .a(n4144), .b(n4116) );
    inv_2 U1894 ( .x(n1530), .a(IR_function_field[0]) );
    inv_5 U1895 ( .x(n744), .a(Imm[22]) );
    inv_2 U1896 ( .x(n1781), .a(reg_out_B[25]) );
    inv_2 U1897 ( .x(n1671), .a(n4146) );
    inv_2 U1899 ( .x(n1797), .a(reg_out_B[23]) );
    inv_2 U190 ( .x(n3558), .a(n3664) );
    inv_2 U1900 ( .x(n1523), .a(IR_function_field[2]) );
    inv_0 U1901 ( .x(n1664), .a(reg_out_B[8]) );
    inv_5 U1902 ( .x(n830), .a(Imm[23]) );
    inv_2 U1903 ( .x(n1752), .a(reg_out_B[28]) );
    inv_2 U1905 ( .x(N144), .a(Imm[31]) );
    inv_2 U1906 ( .x(N70), .a(reg_out_B[31]) );
    inv_8 U1907 ( .x(n653), .a(reg_out_B[12]) );
    or2_2 U1908 ( .x(n496), .a(reg_out_B[0]), .b(IR_function_field[0]) );
    or2_2 U1909 ( .x(n497), .a(IR_opcode_field[1]), .b(net152465) );
    nand2_2 U191 ( .x(n3559), .a(n665), .b(n3630) );
    aoi21_6 U1910 ( .x(n499), .a(n2890), .b(n1602), .c(n3532) );
    aoi21_4 U1911 ( .x(n500), .a(n1685), .b(n541), .c(n3558) );
    and2_3 U1912 ( .x(n501), .a(n549), .b(n548) );
    and2_8 U1913 ( .x(n502), .a(n619), .b(n1444) );
    inv_16 U1914 ( .x(n650), .a(n1574) );
    oa21_2 U1915 ( .x(n503), .a(net149120), .b(n517), .c(n4140) );
    inv_2 U1916 ( .x(n805), .a(n810) );
    and2_6 U1917 ( .x(n810), .a(n803), .b(IR_opcode_field[3]) );
    and2_8 U1918 ( .x(n504), .a(n726), .b(n725) );
    oaoi211_4 U1919 ( .x(n578), .a(n3585), .b(n575), .c(n576), .d(n577) );
    nand2i_2 U192 ( .x(n1418), .a(n1676), .b(___cell__39620_net144330) );
    inv_16 U1920 ( .x(n855), .a(reg_out_B[4]) );
    inv_2 U1921 ( .x(n675), .a(IR_opcode_field[1]) );
    or2_4 U1922 ( .x(n1524), .a(IR_function_field[1]), .b(IR_function_field[0]
        ) );
    oa22_4 U1923 ( .x(n510), .a(n1580), .b(n1651), .c(n1578), .d(n890) );
    inv_2 U1924 ( .x(n1584), .a(n634) );
    buf_12 U1925 ( .x(n583), .a(reg_out_A[22]) );
    inv_2 U1926 ( .x(n3532), .a(n3758) );
    nand2i_2 U1927 ( .x(n3758), .a(n1655), .b(n811) );
    inv_2 U1928 ( .x(n671), .a(n891) );
    inv_12 U1929 ( .x(n748), .a(reg_out_A[20]) );
    nand2i_2 U193 ( .x(n3716), .a(n748), .b(n2070) );
    mux2_4 U1930 ( .x(n513), .d0(n3379), .sl(n729), .d1(n3374) );
    inv_5 U1931 ( .x(n3335), .a(n2133) );
    nand2i_2 U1932 ( .x(n3699), .a(n1693), .b(n977) );
    inv_14 U1933 ( .x(n834), .a(n833) );
    and2_1 U1934 ( .x(n514), .a(n675), .b(net152465) );
    aoi222_1 U1935 ( .x(n515), .a(n1267), .b(n3008), .c(n2022), .d(n3009), .e(
        n2024), .f(n3010) );
    or2_6 U1936 ( .x(n1043), .a(n637), .b(Imm[3]) );
    inv_2 U1937 ( .x(n1333), .a(n4005) );
    nand2i_8 U1938 ( .x(___cell__39620_net144170), .a(IR_opcode_field[0]), .b(
        n1520) );
    ao22_3 U1939 ( .x(n518), .a(n1095), .b(n2988), .c(n1197), .d(n2989) );
    nand2_2 U194 ( .x(n1837), .a(n2268), .b(n910) );
    ao21_4 U1940 ( .x(n519), .a(n1238), .b(n1239), .c(___cell__39620_net143287
        ) );
    mux2i_1 U1941 ( .x(n2581), .d0(n3444), .sl(net149120), .d1(n3788) );
    inv_16 U1942 ( .x(n943), .a(n941) );
    oa22_4 U1943 ( .x(n520), .a(n1644), .b(n889), .c(n1646), .d(n1651) );
    ao22_6 U1944 ( .x(n521), .a(n858), .b(n3584), .c(n2184), .d(n857) );
    inv_2 U1945 ( .x(n3307), .a(n761) );
    inv_14 U1946 ( .x(n862), .a(reg_out_A[17]) );
    oai22_5 U1947 ( .x(n3019), .a(n1529), .b(n880), .c(n822), .d(n1657) );
    inv_7 U1948 ( .x(n3357), .a(n3019) );
    inv_0 U1949 ( .x(n523), .a(n930) );
    nand2_2 U195 ( .x(n3279), .a(n3554), .b(n3555) );
    inv_2 U1950 ( .x(n524), .a(n523) );
    oai22_1 U1951 ( .x(n525), .a(n880), .b(n1648), .c(n822), .d(n1647) );
    inv_14 U1952 ( .x(n880), .a(n1643) );
    inv_10 U1953 ( .x(n3366), .a(n3369) );
    oai22_6 U1954 ( .x(n3369), .a(n1580), .b(n1629), .c(n748), .d(n881) );
    nand4_1 U1955 ( .x(n2865), .a(n2858), .b(n2866), .c(n2855), .d(n2862) );
    aoi22_2 U1956 ( .x(n3098), .a(n1256), .b(n1997), .c(n1249), .d(n3036) );
    aoi22_2 U1957 ( .x(n3035), .a(n1714), .b(n1997), .c(n1256), .d(n3036) );
    nand2i_2 U1958 ( .x(n3918), .a(n4009), .b(n1997) );
    inv_2 U1959 ( .x(n1767), .a(N1890) );
    nand2_2 U196 ( .x(n3339), .a(n1691), .b(n749) );
    inv_2 U1960 ( .x(n526), .a(n3357) );
    inv_1 U1961 ( .x(n527), .a(n799) );
    aoi22_3 U1962 ( .x(n2925), .a(n1714), .b(n2851), .c(n1256), .d(n2852) );
    inv_5 U1963 ( .x(n538), .a(n1580) );
    inv_0 U1964 ( .x(n1874), .a(reg_out_B[15]) );
    exnor2_1 U1965 ( .x(n1505), .a(reg_out_B[15]), .b(n608) );
    nand2i_2 U1966 ( .x(n1956), .a(reg_out_B[15]), .b(n1955) );
    inv_0 U1967 ( .x(n1789), .a(reg_out_B[24]) );
    exnor2_1 U1968 ( .x(n1485), .a(n541), .b(reg_out_B[24]) );
    inv_8 U197 ( .x(n1691), .a(n1688) );
    and4i_2 U1970 ( .x(n1035), .a(n3138), .b(n3135), .c(n3136), .d(n3137) );
    and4i_3 U1971 ( .x(n1034), .a(n1402), .b(n1399), .c(n1400), .d(n1401) );
    inv_14 U1972 ( .x(n689), .a(n688) );
    aoi22_4 U1973 ( .x(n528), .a(reg_out_A[29]), .b(n529), .c(reg_out_A[21]), 
        .d(n883) );
    inv_5 U1974 ( .x(n3302), .a(n528) );
    inv_12 U1975 ( .x(n530), .a(n646) );
    and2_8 U1976 ( .x(n531), .a(n532), .b(___cell__39620_net144317) );
    inv_6 U1977 ( .x(n532), .a(n1603) );
    inv_12 U1979 ( .x(n533), .a(n1587) );
    nand2i_2 U198 ( .x(n3690), .a(n1546), .b(n1968) );
    oai21_3 U1980 ( .x(n3992), .a(n1433), .b(n1944), .c(n810) );
    inv_16 U1981 ( .x(n536), .a(n1546) );
    aoi221_1 U1982 ( .x(n2569), .a(n2543), .b(n2570), .c(n538), .d(n2490), .e(
        n2571) );
    oai21_1 U1983 ( .x(n2449), .a(n1732), .b(n2410), .c(n538) );
    nand2_0 U1984 ( .x(n2412), .a(Imm[28]), .b(n538) );
    nand2i_2 U1985 ( .x(n1711), .a(___cell__39620_net144317), .b(
        ___cell__39620_net144517) );
    nand2i_2 U1986 ( .x(n1682), .a(___cell__39620_net144317), .b(n1683) );
    nand2i_2 U1987 ( .x(n3694), .a(___cell__39620_net144317), .b(n1349) );
    nand2i_2 U1988 ( .x(n3717), .a(___cell__39620_net144317), .b(n1042) );
    inv_2 U1989 ( .x(n534), .a(___cell__39620_net144317) );
    inv_4 U199 ( .x(n935), .a(reg_out_A[6]) );
    inv_2 U1991 ( .x(n535), .a(___cell__39620_net144257) );
    inv_2 U1992 ( .x(___cell__39620_net144257), .a(reg_out_A[30]) );
    inv_5 U1993 ( .x(n1546), .a(reg_out_B[3]) );
    inv_2 U1994 ( .x(n537), .a(n1587) );
    inv_8 U1995 ( .x(n1580), .a(reg_out_A[28]) );
    inv_5 U1996 ( .x(n539), .a(n1564) );
    inv_5 U1997 ( .x(n1564), .a(reg_out_A[29]) );
    inv_10 U1998 ( .x(n3433), .a(n3602) );
    nand4i_2 U1999 ( .x(n2387), .a(n1183), .b(n2385), .c(n2383), .d(n2388) );
    nand2i_4 U200 ( .x(n3340), .a(n1649), .b(n883) );
    mx4_4 U2000 ( .x(n2382), .d0(N1727), .sl0(___cell__39620_net145190), .d1(
        n556), .sl1(n663), .d2(N1892), .sl2(n3998), .d3(N1760), .sl3(n562) );
    nor2i_1 U2001 ( .x(n1278), .a(n1177), .b(n1279) );
    inv_2 U2002 ( .x(n1279), .a(n3318) );
    inv_16 U2003 ( .x(n590), .a(n1219) );
    inv_5 U2004 ( .x(n540), .a(n1573) );
    inv_5 U2005 ( .x(n541), .a(n1578) );
    inv_2 U2006 ( .x(n543), .a(reset) );
    inv_2 U2007 ( .x(n542), .a(reset) );
    inv_2 U2008 ( .x(n4017), .a(reset) );
    aoi221_3 U2009 ( .x(n2313), .a(N1761), .b(___cell__39620_net145150), .c(
        N1728), .d(___cell__39620_net145190), .e(n613) );
    aoai211_1 U201 ( .x(n3179), .a(n2066), .b(n902), .c(n2067), .d(n504) );
    nand2_8 U2010 ( .x(n825), .a(n1630), .b(n1546) );
    oai211_1 U2011 ( .x(n544), .a(n3460), .b(n719), .c(n3858), .d(n2782) );
    nand2i_6 U2012 ( .x(n3858), .a(___cell__39620_net144062), .b(n2520) );
    oai211_3 U2013 ( .x(n2802), .a(n3460), .b(n719), .c(n3858), .d(n2782) );
    inv_10 U2014 ( .x(n1630), .a(n1556) );
    and3i_3 U2015 ( .x(n2017), .a(n2030), .b(n2033), .c(n2034) );
    oai211_4 U2016 ( .x(n2030), .a(n868), .b(n702), .c(n2031), .d(n2032) );
    aoi22_1 U2017 ( .x(n2906), .a(___cell__39620_net143722), .b(n2910), .c(
        ___cell__39620_net143864), .d(n2911) );
    inv_2 U2018 ( .x(n546), .a(n545) );
    inv_14 U2019 ( .x(n889), .a(n888) );
    inv_2 U202 ( .x(n2160), .a(n3350) );
    nand2_2 U2020 ( .x(n779), .a(___cell__39620_net144029), .b(n780) );
    inv_10 U2021 ( .x(___cell__39620_net144029), .a(Imm[12]) );
    or3i_5 U2023 ( .x(n774), .a(n775), .b(Imm[7]), .c(Imm[30]) );
    ao22_6 U2024 ( .x(n3085), .a(n764), .b(n3112), .c(n3054), .d(n765) );
    mux2i_3 U2025 ( .x(n842), .d0(n856), .sl(n848), .d1(n3368) );
    aoi21_1 U2026 ( .x(n2232), .a(n1249), .b(n2233), .c(n1134) );
    nand2_1 U2027 ( .x(n3692), .a(n1256), .b(n2233) );
    nand2_1 U2028 ( .x(n3668), .a(n1714), .b(n2233) );
    buf_3 U2029 ( .x(n547), .a(n584) );
    inv_5 U203 ( .x(n1175), .a(n823) );
    and2_3 U2030 ( .x(n584), .a(n585), .b(n644) );
    nand4_1 U2031 ( .x(n4075), .a(n1014), .b(n1012), .c(n1013), .d(n1011) );
    inv_2 U2032 ( .x(n548), .a(n1577) );
    inv_5 U2033 ( .x(n1577), .a(n893) );
    inv_2 U2034 ( .x(n549), .a(n1603) );
    inv_5 U2035 ( .x(n1569), .a(n910) );
    and4i_5 U2036 ( .x(n1551), .a(n1960), .b(n1958), .c(n600), .d(n601) );
    inv_2 U2037 ( .x(n600), .a(n4139) );
    oai22_5 U2039 ( .x(n2520), .a(n1586), .b(n836), .c(n3391), .d(n4125) );
    nor2_1 U204 ( .x(n897), .a(n899), .b(n898) );
    oai211_3 U2040 ( .x(n1423), .a(n3506), .b(n1602), .c(n665), .d(n2812) );
    aoi21_3 U2041 ( .x(n2812), .a(n1147), .b(n1049), .c(n1834) );
    nand4_4 U2042 ( .x(n2938), .a(n3895), .b(n3894), .c(n3893), .d(n3892) );
    nand2i_6 U2043 ( .x(n3895), .a(n719), .b(n3069) );
    inv_5 U2044 ( .x(n551), .a(___cell__39620_net144781) );
    inv_5 U2045 ( .x(___cell__39620_net144781), .a(Imm[20]) );
    aoi21_3 U2046 ( .x(n2344), .a(n1147), .b(n1047), .c(n1738) );
    inv_16 U2047 ( .x(n3355), .a(n521) );
    inv_5 U2048 ( .x(n762), .a(n3416) );
    nor3_5 U2049 ( .x(n2940), .a(n2939), .b(n2941), .c(n2942) );
    oa22_3 U205 ( .x(n508), .a(n880), .b(n1648), .c(n822), .d(n1647) );
    nand2i_1 U2050 ( .x(n3871), .a(n4010), .b(n3483) );
    nand2i_3 U2051 ( .x(n3893), .a(n1623), .b(n3483) );
    aoi21_2 U2052 ( .x(n2747), .a(n1221), .b(n2609), .c(n2743) );
    aoi22_1 U2053 ( .x(n2653), .a(n1221), .b(n2532), .c(n650), .d(n2609) );
    aoi21_1 U2054 ( .x(n2698), .a(n1191), .b(n2609), .c(n2699) );
    nand3_0 U2055 ( .x(n552), .a(n810), .b(___cell__39620_net144166), .c(
        ___cell__39620_net143655) );
    inv_2 U2056 ( .x(n3998), .a(n552) );
    inv_2 U2057 ( .x(___cell__39620_net144166), .a(IR_opcode_field[0]) );
    mux2i_3 U2058 ( .x(n3283), .d0(n1949), .sl(IR_function_field[2]), .d1(
        n1948) );
    inv_2 U206 ( .x(n3450), .a(n897) );
    nand4i_2 U2060 ( .x(n797), .a(___cell__39620_net147731), .b(n652), .c(n708
        ), .d(N1994) );
    nand2i_4 U2061 ( .x(n2298), .a(n1596), .b(N371) );
    nand3_2 U2062 ( .x(n2910), .a(n3878), .b(n3877), .c(n2887) );
    aoi22_2 U2063 ( .x(n2887), .a(n1249), .b(n2888), .c(n1714), .d(n2690) );
    inv_6 U2064 ( .x(n769), .a(n704) );
    inv_14 U2065 ( .x(n839), .a(n569) );
    nand4_1 U2066 ( .x(n3108), .a(n3115), .b(n3114), .c(n3109), .d(n3111) );
    nand2i_8 U2067 ( .x(n3484), .a(n1584), .b(n928) );
    nand2_0 U2068 ( .x(n3644), .a(___cell__39620_net144330), .b(n533) );
    nand2_0 U2069 ( .x(n3652), .a(___cell__39620_net144330), .b(reg_out_A[30])
         );
    nand2i_3 U207 ( .x(n3470), .a(n3471), .b(n3472) );
    oa21_6 U2070 ( .x(n553), .a(n3426), .b(n618), .c(n3572) );
    inv_10 U2071 ( .x(n2386), .a(n553) );
    aoi22_4 U2072 ( .x(n3070), .a(n1256), .b(n2994), .c(n1249), .d(n2995) );
    nand2_8 U2074 ( .x(n2798), .a(n2780), .b(n2778) );
    nor2i_1 U2075 ( .x(n554), .a(N370), .b(n1596) );
    nand2i_1 U2076 ( .x(n3825), .a(n1635), .b(n2433) );
    or2_5 U2077 ( .x(n992), .a(n1749), .b(n1596) );
    nand2i_8 U2078 ( .x(n1596), .a(___cell__39620_net144175), .b(n1597) );
    oai211_3 U2079 ( .x(n3219), .a(n840), .b(___cell__39620_net144345), .c(
        n3199), .d(n3200) );
    nand2i_3 U208 ( .x(n3321), .a(n3322), .b(n3323) );
    nand3i_1 U2080 ( .x(n1937), .a(n1521), .b(IR_function_field[3]), .c(n1938)
         );
    mux2i_1 U2081 ( .x(n3593), .d0(n1531), .sl(IR_function_field[3]), .d1(
        IR_function_field[4]) );
    or3i_3 U2082 ( .x(___cell__39620_net145426), .a(N1828), .b(
        ___cell__39620_net147731), .c(n1077) );
    inv_2 U2084 ( .x(n556), .a(n555) );
    inv_2 U2085 ( .x(n557), .a(n627) );
    buf_16 U2086 ( .x(n838), .a(n937) );
    nand2i_2 U2087 ( .x(n3362), .a(n1583), .b(n928) );
    aoi22_1 U2088 ( .x(n3111), .a(n2024), .b(n3112), .c(n1267), .d(n3113) );
    inv_10 U209 ( .x(n871), .a(n3575) );
    nand2_5 U2090 ( .x(n1973), .a(n1040), .b(n1974) );
    nand2_5 U2091 ( .x(n3343), .a(n1040), .b(n3608) );
    nand2_5 U2092 ( .x(n3325), .a(n1040), .b(n3603) );
    nand2_5 U2093 ( .x(n3311), .a(n1040), .b(n3607) );
    nor2i_3 U2094 ( .x(n2213), .a(n1040), .b(n2214) );
    nor2i_3 U2095 ( .x(n2159), .a(n1040), .b(n2160) );
    oai21_1 U2096 ( .x(n3276), .a(n1577), .b(n1730), .c(n1040) );
    nand2i_8 U2097 ( .x(n1603), .a(___cell__39620_net144329), .b(
        ___cell__39620_net144331) );
    inv_10 U2098 ( .x(n923), .a(n1603) );
    nand2i_4 U2099 ( .x(n3754), .a(n1602), .b(n3687) );
    oai22_1 U210 ( .x(n559), .a(n1569), .b(n871), .c(n4125), .d(n1283) );
    inv_16 U2100 ( .x(___cell__39620_net143997), .a(Imm[14]) );
    inv_2 U2101 ( .x(n3174), .a(n860) );
    oai22_2 U2102 ( .x(n3139), .a(___cell__39620_net144406), .b(n860), .c(
        n3140), .d(n621) );
    mux2i_3 U2103 ( .x(n860), .d0(n3410), .sl(n625), .d1(n850) );
    aoi21_2 U2104 ( .x(n2760), .a(n1085), .b(n2713), .c(n1254) );
    oai211_2 U2105 ( .x(n574), .a(n3656), .b(n1043), .c(n2675), .d(n3846) );
    oai211_3 U2106 ( .x(n4058), .a(n960), .b(___cell__39620_net143287), .c(
        n961), .d(n962) );
    and3i_3 U2107 ( .x(n1545), .a(n1541), .b(IR_function_field[0]), .c(n1448)
         );
    nand2i_2 U2108 ( .x(n3919), .a(n1634), .b(n3369) );
    nand2_6 U2109 ( .x(n1631), .a(n1630), .b(n1546) );
    ao211_4 U211 ( .x(n1042), .a(net151904), .b(n3481), .c(n3465), .d(n1982)
         );
    oai211_2 U2110 ( .x(n4063), .a(n969), .b(___cell__39620_net147731), .c(
        n970), .d(n971) );
    oai22_1 U2111 ( .x(n558), .a(n1569), .b(n871), .c(n4125), .d(n1283) );
    oai22_2 U2112 ( .x(n1995), .a(n1569), .b(n871), .c(n4125), .d(n1283) );
    nand2i_3 U2113 ( .x(n2715), .a(n4029), .b(n3057) );
    ao22_5 U2114 ( .x(n2187), .a(n3327), .b(n763), .c(n887), .d(n3584) );
    inv_2 U2115 ( .x(n1583), .a(n887) );
    exnor2_1 U2116 ( .x(n1498), .a(n887), .b(reg_out_B[19]) );
    nand2_2 U2117 ( .x(n1739), .a(n3573), .b(n887) );
    exnor2_1 U2118 ( .x(n1497), .a(n887), .b(n684) );
    nand2i_2 U2119 ( .x(n2421), .a(n947), .b(N1891) );
    nand2_2 U212 ( .x(n3480), .a(n665), .b(n3635) );
    and4i_4 U2120 ( .x(___cell__39620_net144322), .a(n778), .b(n560), .c(n561), 
        .d(___cell__39620_net144707) );
    inv_2 U2121 ( .x(n560), .a(Imm[31]) );
    inv_2 U2122 ( .x(n561), .a(Imm[19]) );
    inv_2 U2123 ( .x(n562), .a(___cell__39620_net143710) );
    and3i_4 U2124 ( .x(___cell__39620_net144321), .a(n774), .b(n648), .c(n647)
         );
    inv_5 U2125 ( .x(n647), .a(Imm[28]) );
    nand2_1 U2126 ( .x(n2380), .a(n809), .b(N1661) );
    ao221_4 U2127 ( .x(n2209), .a(n2247), .b(n1267), .c(n3702), .d(n563), .e(
        n564) );
    inv_2 U2128 ( .x(n563), .a(n621) );
    inv_2 U2129 ( .x(n564), .a(n2210) );
    nand2_2 U213 ( .x(n3479), .a(n665), .b(n3653) );
    and4i_3 U2130 ( .x(n1016), .a(n2618), .b(n2616), .c(n2614), .d(n2617) );
    inv_10 U2131 ( .x(n884), .a(n623) );
    oai211_4 U2132 ( .x(n2753), .a(n670), .b(n2754), .c(n2755), .d(n2756) );
    nand2_2 U2133 ( .x(n2665), .a(n845), .b(n2022) );
    nand2_2 U2134 ( .x(n2622), .a(n845), .b(n1267) );
    mux2i_3 U2135 ( .x(n845), .d0(n846), .sl(net150405), .d1(n510) );
    oai22_6 U2136 ( .x(n2841), .a(n875), .b(n1182), .c(n2774), .d(n1055) );
    inv_5 U2138 ( .x(n831), .a(n830) );
    nor2_4 U2139 ( .x(___cell__39620_net143596), .a(n788), .b(n790) );
    nand2i_2 U214 ( .x(n3945), .a(n4010), .b(n3547) );
    buf_3 U2140 ( .x(n567), .a(n4139) );
    buf_3 U2141 ( .x(n566), .a(n4139) );
    nand4_3 U2142 ( .x(n3081), .a(n660), .b(n3074), .c(n3080), .d(n3077) );
    mux2i_2 U2143 ( .x(n3171), .d0(n3358), .sl(n816), .d1(n3313) );
    aoi22_3 U2144 ( .x(n1994), .a(n559), .b(n1683), .c(
        ___cell__39620_net144517), .d(n1996) );
    inv_7 U2145 ( .x(n1067), .a(n1996) );
    inv_0 U2146 ( .x(n568), .a(n806) );
    nand2i_8 U2147 ( .x(n806), .a(___cell__39620_net144173), .b(n708) );
    nor2_1 U2148 ( .x(n1206), .a(n1087), .b(n4034) );
    inv_14 U2149 ( .x(n644), .a(n643) );
    nand2i_2 U215 ( .x(n3946), .a(n718), .b(n2927) );
    inv_4 U2150 ( .x(n643), .a(n934) );
    oai211_3 U2151 ( .x(n4076), .a(n987), .b(___cell__39620_net143287), .c(
        n988), .d(n989) );
    aoi21_1 U2152 ( .x(n2092), .a(n1191), .b(n2093), .c(n1105) );
    nand2_8 U2153 ( .x(n569), .a(n1555), .b(n855) );
    aoi21_2 U2154 ( .x(n2228), .a(n1391), .b(n558), .c(n2226) );
    aoi22_2 U2155 ( .x(n2126), .a(n1391), .b(n1996), .c(n1066), .d(n1995) );
    nand3_1 U2156 ( .x(n570), .a(n3853), .b(n3852), .c(n2737) );
    aoi21_2 U2157 ( .x(n2053), .a(n1191), .b(n2054), .c(n1083) );
    aoi21_1 U2158 ( .x(n2091), .a(n1221), .b(n2054), .c(n2085) );
    inv_10 U2159 ( .x(n1417), .a(reg_out_A[17]) );
    nand2i_2 U216 ( .x(n3947), .a(___cell__39620_net144062), .b(n2854) );
    inv_10 U2160 ( .x(n892), .a(reg_out_A[16]) );
    nand2i_1 U2161 ( .x(n3928), .a(n1632), .b(n3019) );
    ao221_5 U2162 ( .x(n2197), .a(n3602), .b(n572), .c(n3691), .d(n824), .e(
        n571) );
    inv_0 U2163 ( .x(n572), .a(n1562) );
    nand2i_4 U2164 ( .x(n3435), .a(n4004), .b(n1969) );
    nand2_4 U2165 ( .x(n1562), .a(n815), .b(reg_out_B[3]) );
    inv_5 U2166 ( .x(n3434), .a(n3691) );
    nand2i_6 U2167 ( .x(n3691), .a(n2111), .b(n3690) );
    nand2i_3 U2168 ( .x(n3602), .a(n3601), .b(n3598) );
    nand4_5 U2169 ( .x(n771), .a(n573), .b(___cell__39620_net144322), .c(n772), 
        .d(___cell__39620_net144321) );
    and4_5 U2170 ( .x(n573), .a(n607), .b(n1980), .c(n1979), .d(n1978) );
    and3i_4 U2171 ( .x(n772), .a(n776), .b(___cell__39620_net145078), .c(
        ___cell__39620_net145077) );
    nor2i_1 U2172 ( .x(n2003), .a(IR_function_field[5]), .b(IR_function_field
        [2]) );
    inv_2 U2173 ( .x(n1521), .a(IR_function_field[5]) );
    nand3i_3 U2174 ( .x(n2059), .a(n1065), .b(n3665), .c(n2044) );
    oai211_2 U2175 ( .x(n4071), .a(n1017), .b(___cell__39620_net147731), .c(
        n1018), .d(n1019) );
    inv_6 U2176 ( .x(n875), .a(n574) );
    inv_10 U2177 ( .x(n3460), .a(n3458) );
    inv_5 U2178 ( .x(n575), .a(n3742) );
    inv_2 U2179 ( .x(n576), .a(n1565) );
    nand2i_4 U218 ( .x(n3456), .a(n1584), .b(n3575) );
    inv_2 U2180 ( .x(n577), .a(n3571) );
    inv_16 U2181 ( .x(n3585), .a(n1558) );
    inv_5 U2183 ( .x(n579), .a(n2056) );
    aoi221_3 U2185 ( .x(n2424), .a(n1197), .b(n2386), .c(N1991), .d(
        ___cell__39620_net145508), .e(n1189) );
    nand2i_4 U2186 ( .x(n2388), .a(n1751), .b(n4000) );
    nand2i_2 U2187 ( .x(n2408), .a(n4036), .b(n3057) );
    nor2i_3 U2188 ( .x(n1084), .a(n1085), .b(n878) );
    inv_2 U2189 ( .x(n2028), .a(n878) );
    inv_5 U219 ( .x(n1331), .a(n1976) );
    inv_10 U2190 ( .x(n3446), .a(n3445) );
    oai22_6 U2191 ( .x(n3445), .a(n889), .b(n1655), .c(n1651), .d(n1654) );
    mux2i_2 U2192 ( .x(n878), .d0(n3414), .sl(reg_out_B[1]), .d1(n3545) );
    nand4_1 U2193 ( .x(n3138), .a(n3145), .b(n3144), .c(n3146), .d(n3147) );
    aoi222_3 U2194 ( .x(n2278), .a(n1066), .b(n2279), .c(n2266), .d(n644), .e(
        n2079), .f(n2280) );
    inv_10 U2195 ( .x(n925), .a(n923) );
    aoi22_4 U2196 ( .x(n2602), .a(n1683), .b(n2303), .c(
        ___cell__39620_net144517), .d(n2603) );
    and4i_3 U2198 ( .x(n580), .a(n581), .b(n3668), .c(n3667), .d(n3666) );
    inv_2 U2199 ( .x(n3669), .a(n580) );
    exnor2_1 U220 ( .x(n1506), .a(net151622), .b(n609) );
    and2_5 U2200 ( .x(n581), .a(n504), .b(n2130) );
    aoi22_4 U2201 ( .x(n2691), .a(n1683), .b(n2603), .c(
        ___cell__39620_net144517), .d(n2520) );
    inv_10 U2202 ( .x(n903), .a(reg_out_A[9]) );
    nand2_2 U2203 ( .x(n3145), .a(n3118), .b(n1204) );
    mux2i_5 U2204 ( .x(n3118), .d0(n499), .sl(n694), .d1(n3531) );
    and4i_3 U2205 ( .x(n2842), .a(n2841), .b(n2843), .c(n2840), .d(n2844) );
    nand2i_2 U2206 ( .x(n2843), .a(n1847), .b(___cell__39620_net145150) );
    inv_6 U2207 ( .x(n3486), .a(n3654) );
    inv_6 U2208 ( .x(n1450), .a(n3862) );
    nand4i_2 U2209 ( .x(n3165), .a(n3166), .b(n3167), .c(n3173), .d(n3169) );
    inv_5 U221 ( .x(n3476), .a(n3577) );
    inv_8 U2210 ( .x(n751), .a(n3576) );
    mux2i_5 U2211 ( .x(n2064), .d0(n520), .sl(net150405), .d1(n3518) );
    nand2i_2 U2212 ( .x(n3198), .a(n1687), .b(n3448) );
    nand2_2 U2213 ( .x(n3448), .a(n3449), .b(n3450) );
    nand3_5 U2215 ( .x(___cell__39620_net143597), .a(___cell__39620_net143326), 
        .b(n657), .c(N1894) );
    oai22_6 U2216 ( .x(n2994), .a(n1219), .b(n822), .c(n557), .d(n881) );
    nand2_5 U2217 ( .x(n3475), .a(n582), .b(n1981) );
    inv_7 U2218 ( .x(n582), .a(n3476) );
    aoi21_2 U2219 ( .x(n1981), .a(net151904), .b(___cell__39620_net144328), 
        .c(n1982) );
    nand2i_2 U222 ( .x(n3914), .a(n1623), .b(n3303) );
    nand2i_2 U2220 ( .x(n3795), .a(n4010), .b(n2603) );
    nand2i_2 U2221 ( .x(n3770), .a(n1623), .b(n2603) );
    mux2_6 U2222 ( .x(n2708), .d0(n3443), .sl(net150620), .d1(n3533) );
    oai22_2 U2223 ( .x(n3443), .a(n1564), .b(n1651), .c(n1219), .d(n889) );
    oai22_5 U2224 ( .x(n3533), .a(n1587), .b(n1651), .c(n891), .d(n3485) );
    nand4_2 U2225 ( .x(n979), .a(n2750), .b(n2751), .c(n2749), .d(n2752) );
    inv_1 U2226 ( .x(n585), .a(n1603) );
    nand2i_3 U2228 ( .x(n3579), .a(n4008), .b(n2179) );
    nand2i_2 U2229 ( .x(n3678), .a(n719), .b(n2179) );
    nand2i_2 U223 ( .x(n3915), .a(n1625), .b(n3033) );
    aoi22_1 U2230 ( .x(n2336), .a(n1391), .b(n2179), .c(
        ___cell__39620_net144517), .d(n2337) );
    aoi21_2 U2231 ( .x(n2178), .a(n1066), .b(n2179), .c(n2176) );
    inv_7 U2232 ( .x(n886), .a(reg_out_A[19]) );
    and4i_4 U2233 ( .x(n1100), .a(n1094), .b(n2073), .c(n2072), .d(n2071) );
    inv_0 U2235 ( .x(n587), .a(___cell__39620_net144029) );
    inv_2 U2236 ( .x(n588), .a(n587) );
    oa22_1 U2237 ( .x(n895), .a(n889), .b(n1656), .c(n1651), .d(n1657) );
    nand4_3 U2238 ( .x(n3746), .a(n2314), .b(n3745), .c(n2312), .d(n2308) );
    inv_10 U2239 ( .x(n1552), .a(n1547) );
    nand4i_4 U2240 ( .x(n1547), .a(n1548), .b(n1551), .c(n1550), .d(n1549) );
    oai21_5 U2241 ( .x(n2433), .a(n536), .b(n3310), .c(n3387) );
    inv_10 U2242 ( .x(n913), .a(reg_out_A[8]) );
    inv_1 U2243 ( .x(n851), .a(reg_out_A[7]) );
    oai22_6 U2244 ( .x(n2181), .a(n1583), .b(n871), .c(n4125), .d(n3324) );
    ao221_4 U2246 ( .x(n2619), .a(n592), .b(n3996), .c(n2022), .d(n2581), .e(
        n591) );
    inv_2 U2247 ( .x(n591), .a(n2620) );
    inv_0 U2248 ( .x(n592), .a(n670) );
    inv_6 U2249 ( .x(n2583), .a(n3996) );
    nand2i_2 U225 ( .x(n3916), .a(___cell__39620_net144062), .b(n4127) );
    mux2i_6 U2250 ( .x(n3996), .d0(n3385), .sl(n816), .d1(n3779) );
    or2_8 U2251 ( .x(n3576), .a(n4140), .b(n593) );
    inv_0 U2252 ( .x(n593), .a(net151904) );
    nand4i_5 U2254 ( .x(n594), .a(n1332), .b(n3954), .c(n3953), .d(n3952) );
    oai221_5 U2255 ( .x(n2512), .a(n1198), .b(n1055), .c(n553), .d(n1182), .e(
        n2513) );
    mux2i_3 U2256 ( .x(n2106), .d0(n520), .sl(n595), .d1(n3525) );
    inv_2 U2257 ( .x(n595), .a(net150620) );
    inv_5 U2258 ( .x(n3525), .a(n2235) );
    nand2i_2 U2259 ( .x(n2637), .a(n1182), .b(n565) );
    nand2i_2 U2260 ( .x(n2590), .a(n1055), .b(n3523) );
    nand2i_2 U2261 ( .x(n3819), .a(n1616), .b(n565) );
    nand2i_2 U2262 ( .x(n3803), .a(n1166), .b(n565) );
    oai21_5 U2263 ( .x(n1738), .a(n890), .b(n1654), .c(n1739) );
    aoi221_1 U2264 ( .x(n3190), .a(n662), .b(n2218), .c(n3181), .d(
        ___cell__39620_net145285), .e(n3187) );
    aoi22_1 U2265 ( .x(n2813), .a(n2811), .b(___cell__39620_net145285), .c(
        n1318), .d(n2218) );
    aoi22_1 U2266 ( .x(n2345), .a(n2343), .b(___cell__39620_net147791), .c(
        n1197), .d(n2218) );
    aoi22_1 U2267 ( .x(n2217), .a(n2215), .b(___cell__39620_net145285), .c(
        n1095), .d(n2218) );
    inv_12 U2268 ( .x(n890), .a(n888) );
    nand2i_2 U227 ( .x(n3917), .a(___cell__39620_net144374), .b(n3034) );
    aoi211_1 U2270 ( .x(n1352), .a(n1318), .b(n2989), .c(n3024), .d(n1351) );
    aoi22_1 U2271 ( .x(n3064), .a(n662), .b(n2989), .c(n1095), .d(n4141) );
    nand2i_4 U2272 ( .x(n2956), .a(n1166), .b(n2989) );
    inv_2 U2273 ( .x(n597), .a(n1660) );
    inv_2 U2274 ( .x(n598), .a(n4001) );
    oai211_2 U2275 ( .x(n4068), .a(___cell__39620_net147731), .b(n1023), .c(
        n1024), .d(n1025) );
    buf_16 U2276 ( .x(n603), .a(n4015) );
    nand4_1 U2277 ( .x(n2149), .a(n2152), .b(n2151), .c(n2147), .d(n2150) );
    nand2_8 U2278 ( .x(n3582), .a(n604), .b(n2181) );
    inv_2 U2279 ( .x(n604), .a(___cell__39620_net144374) );
    oai22_5 U228 ( .x(n1997), .a(n1577), .b(n881), .c(n1578), .d(n822) );
    inv_12 U2280 ( .x(n3600), .a(n3599) );
    nand2i_4 U2281 ( .x(n606), .a(n738), .b(n531) );
    inv_5 U2282 ( .x(n738), .a(Imm[2]) );
    nand4_1 U2284 ( .x(n4072), .a(n519), .b(n980), .c(n981), .d(n982) );
    inv_5 U2285 ( .x(n607), .a(Imm[26]) );
    nand4_3 U2286 ( .x(n3539), .a(n3717), .b(n3716), .c(n2216), .d(n1419) );
    nand4i_2 U2287 ( .x(n1345), .a(n518), .b(n2986), .c(n2985), .d(n2987) );
    inv_5 U2289 ( .x(n879), .a(reg_out_B[1]) );
    nand2i_2 U229 ( .x(n3921), .a(n1635), .b(n3036) );
    and2_2 U2290 ( .x(n622), .a(reg_out_A[9]), .b(n923) );
    and4_5 U2291 ( .x(n1550), .a(n1962), .b(n656), .c(n1961), .d(n1760) );
    inv_5 U2292 ( .x(n1961), .a(n736) );
    inv_2 U2294 ( .x(n936), .a(n935) );
    or2_6 U2295 ( .x(n1519), .a(IR_opcode_field[4]), .b(IR_opcode_field[5]) );
    nor2_1 U2296 ( .x(n1086), .a(n679), .b(n4044) );
    nand2i_8 U2297 ( .x(n610), .a(n1605), .b(n1606) );
    nand4i_5 U2298 ( .x(n3723), .a(n2274), .b(n3721), .c(n2276), .d(n3722) );
    aoi221_1 U2299 ( .x(n2599), .a(n1095), .b(n2600), .c(n1197), .d(n2557), 
        .e(n1228) );
    nand2i_2 U230 ( .x(n3927), .a(n1634), .b(n2888) );
    aoi21_1 U2300 ( .x(n1244), .a(n662), .b(n2557), .c(n1242) );
    aoi22_1 U2301 ( .x(n2556), .a(N1855), .b(n4000), .c(n1095), .d(n2557) );
    oai211_4 U2302 ( .x(n3856), .a(n3639), .b(n4005), .c(n2721), .d(n3855) );
    inv_0 U2303 ( .x(n611), .a(net156363) );
    inv_0 U2304 ( .x(n612), .a(n663) );
    or2_2 U2305 ( .x(n614), .a(n611), .b(n612) );
    inv_0 U2306 ( .x(n616), .a(n706) );
    aoi222_1 U2307 ( .x(n2840), .a(N1651), .b(n809), .c(n2839), .d(
        ___cell__39620_net147791), .e(n663), .f(n534) );
    nor2i_3 U2308 ( .x(n617), .a(net149627), .b(n779) );
    inv_4 U2309 ( .x(n776), .a(n617) );
    nand2i_2 U231 ( .x(n3929), .a(n1635), .b(n3020) );
    inv_12 U2310 ( .x(net149627), .a(Imm[8]) );
    inv_2 U2311 ( .x(n618), .a(n1333) );
    inv_10 U2312 ( .x(n3426), .a(n3764) );
    and4i_5 U2313 ( .x(___cell__39620_net143595), .a(___cell__39620_net145427), 
        .b(___cell__39620_net145418), .c(___cell__39620_net145426), .d(
        ___cell__39620_net145425) );
    inv_10 U2314 ( .x(n3518), .a(n3516) );
    nand4i_5 U2315 ( .x(n2514), .a(n2512), .b(n2515), .c(n2516), .d(n2517) );
    and2_8 U2316 ( .x(n619), .a(n620), .b(n807) );
    inv_16 U2317 ( .x(___cell__39620_net144175), .a(n619) );
    nand2_8 U2318 ( .x(n621), .a(n619), .b(n1444) );
    inv_10 U2319 ( .x(n1444), .a(n1452) );
    inv_5 U232 ( .x(n3294), .a(n3291) );
    nand2_6 U2320 ( .x(___cell__6067_net21981), .a(n1037), .b(n1038) );
    nand2_2 U2321 ( .x(n3477), .a(n665), .b(n3652) );
    nand2_2 U2322 ( .x(n3478), .a(n665), .b(n3644) );
    inv_5 U2323 ( .x(n1038), .a(counter[0]) );
    oai22_1 U2324 ( .x(n2226), .a(n1570), .b(n1712), .c(n2227), .d(n1711) );
    oai22_6 U2325 ( .x(n3451), .a(n1570), .b(n836), .c(n4125), .d(n2227) );
    oai22_1 U2327 ( .x(n3233), .a(n1577), .b(n1091), .c(n500), .d(n1682) );
    and4i_4 U2328 ( .x(___cell__39620_net145418), .a(n769), .b(
        ___cell__39620_net145421), .c(___cell__39620_net145419), .d(net150643)
         );
    oai221_4 U2329 ( .x(n623), .a(n3509), .b(n1607), .c(n624), .d(n3510), .e(
        n3511) );
    nand2i_2 U233 ( .x(n3922), .a(n1623), .b(n3291) );
    inv_2 U2330 ( .x(n624), .a(n671) );
    inv_4 U2331 ( .x(n3509), .a(n3646) );
    nand2i_1 U2332 ( .x(n3828), .a(n1789), .b(n1064) );
    nand2i_2 U2333 ( .x(n3826), .a(n1789), .b(n1063) );
    oai21_5 U2334 ( .x(___cell__39620_net147278), .a(n3724), .b(
        ___cell__39620_net144345), .c(n2278) );
    oa22_5 U2335 ( .x(n2807), .a(n843), .b(n512), .c(n1175), .d(n1570) );
    and3i_3 U2336 ( .x(n1033), .a(n3081), .b(n3082), .c(n3086) );
    mux2i_5 U2337 ( .x(n3677), .d0(n3313), .sl(n625), .d1(n3314) );
    inv_2 U2338 ( .x(n625), .a(n739) );
    inv_0 U2339 ( .x(n626), .a(n4140) );
    nand2i_2 U234 ( .x(n3923), .a(n4010), .b(n2890) );
    nand2i_0 U2340 ( .x(n3136), .a(___cell__39620_net144655), .b(
        ___cell__39620_net145617) );
    inv_0 U2341 ( .x(n627), .a(n1417) );
    inv_0 U2342 ( .x(n629), .a(n905) );
    oai211_1 U2344 ( .x(n4060), .a(n1034), .b(___cell__39620_net147731), .c(
        n1035), .d(n1036) );
    aoi21_1 U2345 ( .x(n3122), .a(n662), .b(n1380), .c(n1398) );
    aoi22_1 U2346 ( .x(n3029), .a(n1095), .b(n1380), .c(n1197), .d(n594) );
    and4i_5 U2347 ( .x(n840), .a(n841), .b(n2334), .c(n3758), .d(n3753) );
    inv_16 U2348 ( .x(___cell__39620_net143962), .a(Imm[16]) );
    inv_10 U2349 ( .x(n1334), .a(n3475) );
    nand2i_2 U235 ( .x(n3924), .a(n718), .b(n2783) );
    oai22_2 U2350 ( .x(n2116), .a(n884), .b(n1616), .c(
        ___cell__39620_net143658), .d(n2112) );
    nor2i_3 U2351 ( .x(n1094), .a(n1095), .b(n884) );
    aoi22_1 U2352 ( .x(n2801), .a(n544), .b(___cell__39620_net143864), .c(
        n1204), .d(n2803) );
    aoi221_1 U2353 ( .x(n2580), .a(n2581), .b(n1267), .c(reg_out_B[25]), .d(
        n1064), .e(n2582) );
    aoi222_2 U2354 ( .x(n2182), .a(n1256), .b(n1999), .c(n2183), .d(n2184), 
        .e(n2185), .f(n636) );
    inv_14 U2355 ( .x(n1256), .a(n1634) );
    nand2_5 U2356 ( .x(n1622), .a(n923), .b(net149167) );
    inv_1 U2357 ( .x(n632), .a(Imm[18]) );
    nor2_0 U2358 ( .x(n801), .a(IR_opcode_field[2]), .b(IR_opcode_field[4]) );
    nand2i_0 U2359 ( .x(n1614), .a(IR_opcode_field[4]), .b(IR_opcode_field[5])
         );
    nand2i_2 U236 ( .x(n3925), .a(n4008), .b(n2784) );
    buf_10 U2360 ( .x(n634), .a(reg_out_A[23]) );
    inv_0 U2361 ( .x(n641), .a(Imm[6]) );
    inv_2 U2362 ( .x(n642), .a(n641) );
    exnor2_1 U2363 ( .x(n1502), .a(reg_out_B[17]), .b(n902) );
    aoi22_1 U2364 ( .x(n2928), .a(reg_out_B[17]), .b(n2929), .c(n2024), .d(
        n2930) );
    nand3i_4 U2365 ( .x(n646), .a(___cell__39620_net144175), .b(n1528), .c(
        n645) );
    inv_2 U2366 ( .x(n645), .a(n1524) );
    nor2_8 U2367 ( .x(n777), .a(Imm[20]), .b(n631) );
    nor2i_3 U2368 ( .x(n651), .a(n896), .b(n1573) );
    or3i_3 U2369 ( .x(n789), .a(N1729), .b(___cell__39620_net147731), .c(
        ___cell__39620_net143660) );
    exnor2_1 U237 ( .x(n1503), .a(reg_out_B[16]), .b(n893) );
    inv_2 U2370 ( .x(n652), .a(___cell__39620_net144360) );
    nand4_1 U2371 ( .x(n1548), .a(n1954), .b(n653), .c(n1953), .d(n1952) );
    ao221_4 U2372 ( .x(n2939), .a(n3902), .b(n654), .c(n3903), .d(n655), .e(
        n516) );
    inv_0 U2373 ( .x(n654), .a(n621) );
    inv_2 U2374 ( .x(n655), .a(___cell__39620_net144406) );
    inv_2 U2375 ( .x(n656), .a(reg_out_B[31]) );
    nand2i_8 U2376 ( .x(n1700), .a(n766), .b(n1701) );
    nand2_8 U2377 ( .x(n1633), .a(n896), .b(reg_out_B[4]) );
    oai221_5 U2378 ( .x(n2600), .a(n1324), .b(n4005), .c(n3421), .d(n4006), 
        .e(n1806) );
    inv_2 U2379 ( .x(n657), .a(n947) );
    inv_14 U238 ( .x(n631), .a(___cell__39620_net143962) );
    nand2i_6 U2380 ( .x(n1688), .a(reg_out_B[3]), .b(n1689) );
    and2_8 U2381 ( .x(n658), .a(n1689), .b(reg_out_A[30]) );
    oai211_2 U2382 ( .x(n4061), .a(___cell__39620_net143287), .b(n966), .c(
        n967), .d(n968) );
    inv_0 U2383 ( .x(n659), .a(reg_out_B[3]) );
    oai211_2 U2384 ( .x(n4056), .a(___cell__39620_net143287), .b(n957), .c(
        n958), .d(n959) );
    inv_6 U2385 ( .x(n660), .a(n3071) );
    nand2i_8 U2386 ( .x(n1642), .a(reg_out_B[2]), .b(n882) );
    oai211_2 U2387 ( .x(n1968), .a(n855), .b(n3596), .c(n1040), .d(n3353) );
    inv_16 U2388 ( .x(n815), .a(n828) );
    ao31_4 U2389 ( .x(n2402), .a(n2629), .b(n763), .c(n828), .d(n819) );
    inv_2 U239 ( .x(n1861), .a(N1748) );
    ao22_1 U2390 ( .x(n3378), .a(n828), .b(n3307), .c(n826), .d(n813) );
    nand2_2 U2391 ( .x(n1419), .a(n664), .b(___cell__39620_net144328) );
    nand2_8 U2392 ( .x(n665), .a(n664), .b(___cell__39620_net144328) );
    inv_16 U2393 ( .x(___cell__39620_net144328), .a(___cell__39620_net144324)
         );
    inv_2 U2394 ( .x(___cell__39620_net144326), .a(net151578) );
    oai221_2 U2395 ( .x(n2874), .a(n752), .b(n1635), .c(n3447), .d(n4009), .e(
        n2850) );
    inv_14 U2396 ( .x(n1728), .a(n1159) );
    oai22_2 U2397 ( .x(n3382), .a(n1580), .b(n915), .c(n1578), .d(n1642) );
    oa22_2 U2398 ( .x(n761), .a(n1570), .b(n1631), .c(___cell__39620_net144257
        ), .d(n4012) );
    inv_3 U2399 ( .x(n833), .a(reg_out_A[4]) );
    nand2i_5 U240 ( .x(n3764), .a(n751), .b(n3763) );
    nor2i_3 U2400 ( .x(n666), .a(n667), .b(___cell__39620_net144329) );
    inv_4 U2401 ( .x(n1624), .a(n666) );
    inv_0 U2402 ( .x(n667), .a(___cell__39620_net144331) );
    ao22_3 U2403 ( .x(n3166), .a(n3981), .b(n668), .c(n766), .d(n818) );
    inv_2 U2404 ( .x(n668), .a(n670) );
    nand2_2 U2405 ( .x(n1637), .a(n669), .b(n1638) );
    inv_1 U2406 ( .x(n669), .a(___cell__39620_net144175) );
    nand2_5 U2407 ( .x(n670), .a(n669), .b(n1638) );
    nand3_2 U2408 ( .x(n3007), .a(n3011), .b(n515), .c(n3015) );
    nand2i_8 U2409 ( .x(___cell__39620_net144329), .a(Imm[5]), .b(n773) );
    inv_4 U241 ( .x(n3639), .a(n3638) );
    nand2i_2 U2410 ( .x(n3948), .a(n1632), .b(n525) );
    nand3_4 U2411 ( .x(n2299), .a(N1861), .b(n4000), .c(
        ___cell__39620_net147732) );
    aoi22_1 U2412 ( .x(n3191), .a(N1831), .b(n4000), .c(N1964), .d(
        ___cell__39620_net145508) );
    or2_8 U2413 ( .x(n3628), .a(n3395), .b(n610) );
    inv_3 U2414 ( .x(n3395), .a(n3626) );
    nor2_0 U2415 ( .x(___cell__39620_net143982), .a(___cell__39620_net143693), 
        .b(___cell__39620_net143983) );
    nor2_3 U2418 ( .x(n1962), .a(reg_out_B[16]), .b(reg_out_B[17]) );
    inv_0 U2419 ( .x(n1866), .a(reg_out_B[16]) );
    nand2i_4 U242 ( .x(n2722), .a(n751), .b(n3818) );
    or2_8 U2420 ( .x(n3511), .a(n1072), .b(n672) );
    and2_8 U2421 ( .x(n673), .a(net149167), .b(n891) );
    nand2i_2 U2422 ( .x(n1072), .a(net149167), .b(n891) );
    inv_16 U2423 ( .x(n1289), .a(n1607) );
    oai21_6 U2424 ( .x(n2384), .a(n3524), .b(n4005), .c(n3572) );
    nand2i_2 U2425 ( .x(n3572), .a(n4140), .b(n1043) );
    and3i_4 U2426 ( .x(n674), .a(___cell__39620_net147731), .b(n676), .c(n514)
         );
    inv_12 U2427 ( .x(n784), .a(n674) );
    and2_8 U2428 ( .x(n676), .a(n677), .b(___cell__39620_net144344) );
    inv_0 U2429 ( .x(n677), .a(IR_opcode_field[0]) );
    nand2i_2 U243 ( .x(n3884), .a(n4005), .b(n3658) );
    or2_8 U2430 ( .x(n3646), .a(n3497), .b(n610) );
    inv_3 U2431 ( .x(n3497), .a(n3645) );
    inv_16 U2432 ( .x(n942), .a(n941) );
    mux2i_3 U2433 ( .x(n2710), .d0(n3536), .sl(net149120), .d1(n510) );
    inv_10 U2434 ( .x(n3536), .a(n3535) );
    nor2i_3 U2435 ( .x(n1663), .a(n2006), .b(n1543) );
    oai22_3 U2436 ( .x(n2570), .a(n1573), .b(n890), .c(
        ___cell__39620_net144257), .d(n1651) );
    inv_16 U2437 ( .x(n1651), .a(n811) );
    inv_0 U2438 ( .x(___cell__39620_net144605), .a(Imm[29]) );
    buf_16 U2439 ( .x(n832), .a(reg_out_A[1]) );
    nand2i_6 U244 ( .x(n3658), .a(n3542), .b(n3627) );
    buf_16 U2440 ( .x(n921), .a(n937) );
    inv_14 U2441 ( .x(n681), .a(n680) );
    aoi22_2 U2442 ( .x(n3114), .a(n502), .b(n3116), .c(n3117), .d(
        ___cell__39620_net143722) );
    mux2i_2 U2443 ( .x(n3117), .d0(n3417), .sl(n816), .d1(n3358) );
    nand2i_2 U2444 ( .x(n2975), .a(n621), .b(n3010) );
    aoi22_2 U2445 ( .x(n1967), .a(n1964), .b(n1968), .c(n1330), .d(n1969) );
    aoi22_2 U2446 ( .x(n3021), .a(n1971), .b(n3022), .c(n1330), .d(n1968) );
    nand4_1 U2447 ( .x(n3010), .a(n3921), .b(n3920), .c(n3919), .d(n3918) );
    exnor2_1 U2448 ( .x(n1476), .a(reg_out_A[29]), .b(reg_out_B[29]) );
    inv_10 U2449 ( .x(n747), .a(n685) );
    inv_5 U245 ( .x(n3306), .a(n3303) );
    nand2i_8 U2450 ( .x(n1557), .a(n1039), .b(n1558) );
    buf_12 U2451 ( .x(n686), .a(reg_out_A[22]) );
    nor2i_3 U2452 ( .x(n1134), .a(n838), .b(n1122) );
    nor2i_3 U2453 ( .x(n1133), .a(n838), .b(n1120) );
    aoai211_1 U2454 ( .x(n2790), .a(n749), .b(n530), .c(n1064), .d(reg_out_B
        [20]) );
    exnor2_1 U2455 ( .x(n1493), .a(reg_out_B[20]), .b(n749) );
    inv_16 U2456 ( .x(n691), .a(n940) );
    inv_16 U2457 ( .x(n692), .a(n691) );
    nand2_6 U2458 ( .x(n3303), .a(n3304), .b(n3305) );
    nand2_2 U2459 ( .x(n3647), .a(n923), .b(n634) );
    nand2i_2 U246 ( .x(n3885), .a(n1625), .b(n3303) );
    or3i_2 U2461 ( .x(n1940), .a(n2002), .b(n693), .c(n1521) );
    inv_0 U2462 ( .x(n693), .a(IR_function_field[4]) );
    ao22_6 U2463 ( .x(n1996), .a(reg_out_A[20]), .b(n3575), .c(n3464), .d(n799
        ) );
    buf_16 U2464 ( .x(n694), .a(net149107) );
    nand2_8 U2465 ( .x(n696), .a(n713), .b(n928) );
    ao211_5 U2466 ( .x(n2857), .a(n3374), .b(n625), .c(n698), .d(n697) );
    and2_2 U2467 ( .x(n698), .a(n699), .b(n2995) );
    inv_2 U2468 ( .x(n699), .a(n727) );
    inv_16 U2469 ( .x(n816), .a(n879) );
    nand2i_2 U247 ( .x(n3886), .a(___cell__39620_net144062), .b(n3034) );
    inv_0 U2470 ( .x(n700), .a(n702) );
    nand2_8 U2471 ( .x(n703), .a(n701), .b(n1661) );
    nand2i_5 U2472 ( .x(n3613), .a(n3612), .b(n3598) );
    nand2i_2 U2473 ( .x(n3499), .a(n1647), .b(n1689) );
    oa22_2 U2474 ( .x(n856), .a(n815), .b(n761), .c(n1573), .d(n915) );
    inv_16 U2475 ( .x(n901), .a(n900) );
    or3i_4 U2476 ( .x(n704), .a(N1663), .b(n705), .c(___cell__39620_net143872)
         );
    inv_0 U2477 ( .x(n705), .a(___cell__39620_net147732) );
    inv_16 U2478 ( .x(n809), .a(n706) );
    inv_2 U2479 ( .x(n707), .a(n808) );
    nand2i_2 U248 ( .x(n3904), .a(n1562), .b(n2719) );
    inv_0 U2480 ( .x(n710), .a(IR_opcode_field[3]) );
    aoi21_1 U2481 ( .x(n802), .a(IR_opcode_field[0]), .b(
        ___cell__39620_net143655), .c(n800) );
    nand2i_0 U2482 ( .x(n808), .a(IR_opcode_field[1]), .b(n810) );
    inv_2 U2483 ( .x(n726), .a(n816) );
    inv_5 U2484 ( .x(n1451), .a(n816) );
    nand2i_6 U2485 ( .x(n3619), .a(n3618), .b(n3598) );
    inv_2 U2486 ( .x(n841), .a(n3759) );
    nand2i_2 U2487 ( .x(n3906), .a(n4004), .b(n3610) );
    nand4_1 U2488 ( .x(n1000), .a(n3699), .b(n2153), .c(n2146), .d(n2158) );
    nand2i_2 U2489 ( .x(n2158), .a(n1692), .b(n2837) );
    inv_5 U249 ( .x(n1971), .a(n1562) );
    and4i_2 U2490 ( .x(n2153), .a(n2149), .b(n2154), .c(n2155), .d(n2156) );
    oai22_6 U2491 ( .x(n3384), .a(n1564), .b(n915), .c(n1219), .d(n1642) );
    inv_10 U2492 ( .x(n902), .a(n862) );
    ao21_4 U2493 ( .x(n3963), .a(n3415), .b(n711), .c(n712) );
    inv_0 U2494 ( .x(n711), .a(n1451) );
    inv_16 U2495 ( .x(n908), .a(n907) );
    inv_16 U2496 ( .x(n907), .a(reg_out_A[10]) );
    inv_16 U2497 ( .x(n3598), .a(n1557) );
    inv_4 U2498 ( .x(n714), .a(n1067) );
    inv_2 U2499 ( .x(n715), .a(___cell__39620_net144374) );
    buf_1 U25 ( .x(n635), .a(reg_out_A[23]) );
    nand2i_2 U250 ( .x(n3905), .a(n1565), .b(n3613) );
    nand2i_8 U2500 ( .x(___cell__39620_net144062), .a(n891), .b(n717) );
    or2_4 U2501 ( .x(___cell__39620_net144374), .a(n637), .b(n717) );
    or2_4 U2502 ( .x(n719), .a(n637), .b(n717) );
    or2_4 U2503 ( .x(n718), .a(n637), .b(n717) );
    inv_5 U2504 ( .x(n3452), .a(n3451) );
    aoi221_5 U2505 ( .x(n720), .a(n2133), .b(n723), .c(n722), .d(n721), .e(
        n724) );
    inv_2 U2506 ( .x(n721), .a(n727) );
    inv_2 U2507 ( .x(n723), .a(n1635) );
    ao22_3 U2508 ( .x(n724), .a(n1249), .b(n1997), .c(n1256), .d(n847) );
    nand2_1 U2509 ( .x(n727), .a(n726), .b(n725) );
    nand2i_4 U251 ( .x(n3059), .a(n3585), .b(n3817) );
    nor2i_3 U2510 ( .x(n728), .a(n725), .b(n726) );
    inv_10 U2511 ( .x(n1635), .a(n728) );
    inv_5 U2512 ( .x(n3317), .a(n2233) );
    oai22_4 U2513 ( .x(n2130), .a(n3504), .b(n536), .c(n1577), .d(n1629) );
    inv_2 U2514 ( .x(n1178), .a(n3327) );
    inv_16 U2515 ( .x(n887), .a(n886) );
    nand2_1 U2516 ( .x(n3327), .a(n3328), .b(n3329) );
    oai21_5 U2517 ( .x(n3410), .a(n3411), .b(n815), .c(n3412) );
    oai211_2 U2518 ( .x(n4059), .a(n963), .b(___cell__39620_net147731), .c(
        n964), .d(n965) );
    and4i_2 U2519 ( .x(n963), .a(n1413), .b(n1410), .c(n1411), .d(n1412) );
    nand2i_2 U252 ( .x(n3301), .a(n1563), .b(n926) );
    inv_2 U2520 ( .x(n729), .a(n816) );
    oai221_2 U2522 ( .x(n3903), .a(n752), .b(n1636), .c(n3411), .d(n1632), .e(
        n2925) );
    aoi22_2 U2523 ( .x(n2891), .a(n910), .b(n2892), .c(n2024), .d(n2857) );
    and2_8 U2524 ( .x(n735), .a(___cell__39620_net144356), .b(
        ___cell__39620_net143655) );
    inv_14 U2525 ( .x(n946), .a(n735) );
    inv_4 U2526 ( .x(___cell__39620_net143655), .a(n804) );
    nor2_1 U2527 ( .x(___cell__39620_net144356), .a(n805), .b(
        ___cell__39620_net144166) );
    oai22_6 U2528 ( .x(n2888), .a(n1586), .b(n881), .c(n822), .d(n1654) );
    inv_10 U2529 ( .x(n773), .a(n771) );
    inv_5 U2530 ( .x(n1257), .a(n2690) );
    oai211_2 U2531 ( .x(n3289), .a(n3434), .b(n1560), .c(n1040), .d(n2810) );
    ao22_6 U2532 ( .x(n2133), .a(n3336), .b(n812), .c(reg_out_A[20]), .d(n3584
        ) );
    inv_3 U2533 ( .x(n3334), .a(n3336) );
    nand2_2 U2534 ( .x(n3336), .a(n3337), .b(n3338) );
    nor2_8 U2535 ( .x(n813), .a(n1560), .b(n825) );
    oai22_3 U2536 ( .x(n3545), .a(n915), .b(n1646), .c(n1642), .d(n1644) );
    oai22_3 U2537 ( .x(n2236), .a(n1642), .b(n1649), .c(n915), .d(n1647) );
    nor2i_8 U2538 ( .x(n737), .a(n768), .b(n825) );
    inv_16 U2539 ( .x(n883), .a(n825) );
    nand2i_2 U254 ( .x(n3296), .a(n1654), .b(n874) );
    or2_4 U2540 ( .x(n4009), .a(n816), .b(n815) );
    nand2i_8 U2541 ( .x(n1558), .a(n855), .b(n1728) );
    inv_10 U2542 ( .x(n1283), .a(n3467) );
    inv_0 U2543 ( .x(n739), .a(n816) );
    inv_12 U2544 ( .x(n3313), .a(n3312) );
    oai22_5 U2545 ( .x(n2995), .a(n1587), .b(n822), .c(n1583), .d(n881) );
    aoi22_1 U2546 ( .x(n2431), .a(n2432), .b(n590), .c(n1249), .d(n2433) );
    nand2i_2 U2547 ( .x(n3930), .a(n4009), .b(n2690) );
    aoi22_2 U2548 ( .x(n2044), .a(n1683), .b(n2045), .c(
        ___cell__39620_net144517), .d(n1995) );
    oai22_4 U2549 ( .x(n2045), .a(n1577), .b(n871), .c(n500), .d(n4125) );
    nand2i_2 U255 ( .x(n3892), .a(n4008), .b(n2991) );
    aoai211_5 U2550 ( .x(n740), .a(n3862), .b(n741), .c(n742), .d(n1444) );
    inv_5 U2551 ( .x(n1449), .a(n740) );
    inv_2 U2552 ( .x(n741), .a(n1451) );
    nand4i_2 U2553 ( .x(n3862), .a(n1278), .b(n3860), .c(n2807), .d(n3412) );
    nand2i_1 U2554 ( .x(n3759), .a(n1608), .b(n3321) );
    nand2_0 U2555 ( .x(n2912), .a(n640), .b(n902) );
    exnor2_1 U2556 ( .x(n1501), .a(n902), .b(n640) );
    inv_0 U2557 ( .x(___cell__39620_net143954), .a(n640) );
    inv_16 U2558 ( .x(n745), .a(n744) );
    nand2i_2 U2559 ( .x(n2341), .a(n1632), .b(n1999) );
    nand2i_2 U256 ( .x(n3894), .a(n4010), .b(n2992) );
    aoi22_1 U2560 ( .x(n1998), .a(n1999), .b(n504), .c(n1256), .d(n2000) );
    mux2_4 U2561 ( .x(n746), .d0(n3546), .sl(n816), .d1(n3442) );
    aoi221_1 U2562 ( .x(n2188), .a(n2189), .b(___cell__39620_net144345), .c(
        n912), .d(n2190), .e(n1130) );
    inv_2 U2563 ( .x(n3604), .a(n3491) );
    nor2i_0 U2564 ( .x(n2161), .a(net151578), .b(n1656) );
    exnor2_1 U2565 ( .x(n1465), .a(n912), .b(net151578) );
    inv_16 U2566 ( .x(n749), .a(n748) );
    nor2_3 U2567 ( .x(n2146), .a(n2143), .b(n2141) );
    buf_5 U2568 ( .x(n750), .a(n2236) );
    and4i_3 U2569 ( .x(n1262), .a(n2773), .b(n2775), .c(n2776), .d(n2777) );
    exnor2_1 U257 ( .x(n1491), .a(n628), .b(n566) );
    or2_8 U2570 ( .x(n1281), .a(n1684), .b(n671) );
    nand2i_3 U2571 ( .x(n1684), .a(net149167), .b(n1685) );
    inv_4 U2572 ( .x(n1772), .a(N333) );
    oai22_2 U2574 ( .x(n2773), .a(n2774), .b(n1616), .c(n865), .d(n1166) );
    oa211_5 U2575 ( .x(n865), .a(n3629), .b(n1043), .c(n2765), .d(n3859) );
    nand2i_1 U2576 ( .x(n3603), .a(n1587), .b(n896) );
    nand2i_1 U2577 ( .x(n3607), .a(n1219), .b(n896) );
    nand2i_2 U2578 ( .x(n3608), .a(n1564), .b(n896) );
    nand2i_2 U2579 ( .x(n1672), .a(n1673), .b(n896) );
    nand2i_2 U258 ( .x(n3528), .a(n891), .b(n2992) );
    nand2i_3 U2580 ( .x(n3596), .a(___cell__39620_net144257), .b(n896) );
    oa21_6 U2581 ( .x(n752), .a(n2475), .b(reg_out_B[3]), .c(n3551) );
    nand2i_4 U2582 ( .x(n3551), .a(n1648), .b(n3584) );
    inv_16 U2583 ( .x(n753), .a(___cell__39620_net144655) );
    and2_8 U2584 ( .x(n754), .a(n839), .b(reg_out_B[3]) );
    inv_16 U2585 ( .x(n1629), .a(n754) );
    aoi22_1 U2586 ( .x(n2479), .a(n2435), .b(n2277), .c(n2436), .d(n914) );
    aoi21_1 U2587 ( .x(n1082), .a(n914), .b(n530), .c(n1064) );
    aoi22_1 U2588 ( .x(n2281), .a(n2268), .b(n894), .c(n823), .d(n914) );
    inv_2 U2589 ( .x(n1648), .a(n914) );
    nand2i_5 U259 ( .x(n3375), .a(n1219), .b(n3592) );
    aoi22_1 U2590 ( .x(n2562), .a(n2266), .b(n914), .c(n1391), .d(n4134) );
    exnor2_1 U2591 ( .x(n1459), .a(reg_out_B[8]), .b(n914) );
    inv_16 U2592 ( .x(n2475), .a(n2283) );
    inv_0 U2593 ( .x(n755), .a(n703) );
    inv_2 U2594 ( .x(n756), .a(n1658) );
    inv_12 U2595 ( .x(n1249), .a(n1632) );
    inv_0 U2596 ( .x(n757), .a(n784) );
    inv_0 U2597 ( .x(n758), .a(___cell__39620_net144406) );
    and3i_1 U2598 ( .x(n760), .a(reg_out_B[4]), .b(n759), .c(n1552) );
    inv_0 U2599 ( .x(n899), .a(n760) );
    inv_8 U26 ( .x(n1654), .a(reg_out_A[3]) );
    inv_8 U260 ( .x(n529), .a(n1629) );
    inv_3 U2600 ( .x(n1570), .a(n583) );
    oai211_3 U2601 ( .x(n2789), .a(n2655), .b(n1186), .c(n2785), .d(n2790) );
    ao21_4 U2602 ( .x(n3415), .a(n2888), .b(n828), .c(n762) );
    inv_0 U2604 ( .x(n763), .a(reg_out_B[3]) );
    inv_0 U2605 ( .x(n764), .a(n621) );
    inv_2 U2606 ( .x(n765), .a(n670) );
    nand2i_4 U2607 ( .x(n2296), .a(n1592), .b(N338) );
    inv_16 U2608 ( .x(N3304), .a(___cell__6067_net21981) );
    and3i_4 U2609 ( .x(n964), .a(n3165), .b(n3983), .c(n3164) );
    inv_5 U261 ( .x(n1250), .a(n2851) );
    ao222_4 U2610 ( .x(n2930), .a(reg_out_B[1]), .b(n3365), .c(n827), .d(n767), 
        .e(n3036), .f(n768) );
    inv_2 U2611 ( .x(n767), .a(n1634) );
    inv_2 U2612 ( .x(n768), .a(n4009) );
    nor3_3 U2613 ( .x(n982), .a(n2662), .b(n2669), .c(n2666) );
    inv_2 U2614 ( .x(net150643), .a(___cell__39620_net143767) );
    nor2_0 U2615 ( .x(___cell__39620_net143767), .a(n4140), .b(n770) );
    inv_16 U2616 ( .x(___cell__39620_net147732), .a(___cell__39620_net147731)
         );
    nand2i_6 U2618 ( .x(___cell__39620_net144324), .a(N69), .b(n773) );
    nor2_1 U2619 ( .x(___cell__39620_net145077), .a(Imm[14]), .b(Imm[11]) );
    nand2i_2 U262 ( .x(n3373), .a(n1644), .b(n874) );
    nand2i_4 U2620 ( .x(n778), .a(Imm[17]), .b(n777) );
    oai221_4 U2621 ( .x(n790), .a(n792), .b(___cell__39620_net144406), .c(n793
        ), .d(n784), .e(n791) );
    inv_6 U2622 ( .x(n793), .a(___cell__39620_net147278) );
    oai211_3 U2623 ( .x(n788), .a(n503), .b(n785), .c(n787), .d(n789) );
    aoi23_4 U2624 ( .x(n787), .a(n786), .b(___cell__39620_net147732), .c(N1762
        ), .d(___cell__39620_net143326), .e(___cell__39620_net145150) );
    nor2i_5 U2625 ( .x(n786), .a(net151622), .b(n734) );
    inv_16 U2626 ( .x(___cell__39620_net145150), .a(___cell__39620_net143710)
         );
    nand2i_4 U2627 ( .x(n785), .a(___cell__39620_net144343), .b(
        ___cell__39620_net143326) );
    nor2i_5 U2628 ( .x(___cell__39620_net143784), .a(___cell__39620_net143785), 
        .b(n503) );
    nand4i_4 U2629 ( .x(___cell__39620_net145427), .a(___cell__39620_net145428
        ), .b(___cell__39620_net145429), .c(n796), .d(n797) );
    nand2i_2 U263 ( .x(n3377), .a(n1655), .b(n874) );
    inv_16 U2630 ( .x(___cell__39620_net145508), .a(___cell__39620_net143845)
         );
    nand3i_5 U2631 ( .x(n796), .a(___cell__39620_net144062), .b(
        ___cell__39620_net147296), .c(n798) );
    nand2i_6 U2632 ( .x(n794), .a(n4140), .b(n795) );
    inv_16 U2633 ( .x(net151904), .a(___cell__39620_net144331) );
    inv_16 U2634 ( .x(___cell__39620_net144331), .a(Imm[4]) );
    inv_10 U2635 ( .x(n803), .a(IR_opcode_field[2]) );
    and2_5 U2636 ( .x(___cell__39620_net145037), .a(n803), .b(net151497) );
    nand2i_8 U2637 ( .x(___cell__39620_net143710), .a(n803), .b(
        ___cell__39620_net144309) );
    and3i_1 U2638 ( .x(n800), .a(___cell__39620_net143653), .b(n801), .c(
        IR_opcode_field[5]) );
    or3i_1 U2639 ( .x(n804), .a(IR_opcode_field[5]), .b(IR_opcode_field[4]), 
        .c(IR_opcode_field[1]) );
    oai22_5 U264 ( .x(n2690), .a(n1585), .b(n881), .c(n1629), .d(n1655) );
    nand2i_8 U2640 ( .x(___cell__39620_net147731), .a(n807), .b(N3304) );
    nand2i_8 U2641 ( .x(___cell__39620_net143287), .a(n568), .b(N3304) );
    nand2i_6 U2642 ( .x(___cell__39620_net144199), .a(___cell__39620_net144200
        ), .b(n708) );
    nand2_8 U2643 ( .x(___cell__39620_net143658), .a(___cell__39620_net144303), 
        .b(n708) );
    buf_2 U2644 ( .x(n926), .a(n531) );
    inv_16 U2645 ( .x(n1602), .a(Imm[2]) );
    inv_2 U2646 ( .x(net149616), .a(Imm[9]) );
    nand2i_0 U2647 ( .x(n1535), .a(IR_function_field[0]), .b(IR_function_field
        [1]) );
    inv_2 U2648 ( .x(n1534), .a(IR_function_field[1]) );
    ao22_6 U2649 ( .x(n2000), .a(n3346), .b(n812), .c(n628), .d(n3584) );
    nand2i_3 U265 ( .x(n3394), .a(n3395), .b(n3396) );
    inv_0 U2650 ( .x(n812), .a(reg_out_B[3]) );
    inv_4 U2651 ( .x(n3345), .a(n3346) );
    nand2_2 U2652 ( .x(n3346), .a(n3347), .b(n3348) );
    inv_3 U2653 ( .x(n1560), .a(n815) );
    inv_2 U2654 ( .x(n814), .a(n1569) );
    nand2_2 U2655 ( .x(n3318), .a(n3319), .b(n3320) );
    mux2_4 U2656 ( .x(n870), .d0(n3446), .sl(n694), .d1(n589) );
    and2_3 U2657 ( .x(n1978), .a(n817), .b(n905) );
    aoi211_1 U2658 ( .x(n2127), .a(n2079), .b(n2128), .c(n1108), .d(n1109) );
    inv_5 U266 ( .x(n3391), .a(n3496) );
    inv_2 U2660 ( .x(n818), .a(n817) );
    nand2i_0 U2661 ( .x(n2297), .a(n4039), .b(n3057) );
    oai21_3 U2662 ( .x(n3760), .a(net149122), .b(n840), .c(n2336) );
    inv_0 U2663 ( .x(n819), .a(n1159) );
    inv_2 U2664 ( .x(n820), .a(n819) );
    nand2i_2 U2665 ( .x(n3881), .a(n4003), .b(n3599) );
    oai22_1 U2666 ( .x(n2330), .a(n1087), .b(n4038), .c(
        ___cell__39620_net143693), .d(___cell__39620_net144572) );
    and4_5 U2667 ( .x(n2314), .a(n2313), .b(n2316), .c(n2315), .d(n821) );
    nand2i_0 U2668 ( .x(n2315), .a(n4140), .b(n1318) );
    nand2i_3 U2669 ( .x(n3599), .a(n3597), .b(n3598) );
    buf_16 U2670 ( .x(n822), .a(n4012) );
    nor2_3 U2671 ( .x(n823), .a(n1688), .b(n824) );
    inv_0 U2672 ( .x(n824), .a(n815) );
    nand3_5 U2673 ( .x(n3702), .a(n2186), .b(n3701), .c(n2182) );
    buf_16 U2675 ( .x(net149120), .a(net149107) );
    oai21_1 U2677 ( .x(n3247), .a(n3237), .b(n3238), .c(n943) );
    oai21_1 U2678 ( .x(n3241), .a(n943), .b(___cell__39620_net144199), .c(
        n1618) );
    nor3_0 U2679 ( .x(n3256), .a(n1521), .b(IR_function_field[2]), .c(
        IR_function_field[4]) );
    inv_2 U2680 ( .x(n826), .a(n1573) );
    inv_10 U2681 ( .x(n829), .a(n830) );
    inv_6 U2682 ( .x(n909), .a(reg_out_A[18]) );
    exnor2_1 U2684 ( .x(n1513), .a(reg_out_B[11]), .b(n901) );
    inv_0 U2685 ( .x(n1907), .a(reg_out_B[11]) );
    inv_10 U2686 ( .x(net149628), .a(net149627) );
    nand2i_1 U2687 ( .x(n3640), .a(n1603), .b(n902) );
    aoi21_1 U2688 ( .x(n2369), .a(n885), .b(n1733), .c(n1179) );
    aoi21_1 U2689 ( .x(n2147), .a(n885), .b(n2148), .c(n1117) );
    inv_16 U269 ( .x(n874), .a(n1622) );
    aoai211_1 U2690 ( .x(n2357), .a(n885), .b(n530), .c(n1064), .d(n536) );
    exnor2_1 U2691 ( .x(n1473), .a(net149167), .b(n885) );
    exnor2_1 U2692 ( .x(n1474), .a(reg_out_B[3]), .b(n885) );
    inv_0 U2693 ( .x(___cell__39620_net143720), .a(Imm[7]) );
    inv_0 U2694 ( .x(___cell__39620_net144572), .a(Imm[30]) );
    aoi22_2 U2695 ( .x(n2709), .a(n2710), .b(n1267), .c(n2711), .d(n502) );
    inv_2 U2696 ( .x(net151577), .a(Imm[5]) );
    mux2i_1 U2697 ( .x(n1951), .d0(n1446), .sl(reg_out_B[0]), .d1(n1527) );
    exnor2_1 U2698 ( .x(n3274), .a(reg_out_B[0]), .b(n942) );
    nand2i_0 U2699 ( .x(n1628), .a(IR_function_field[0]), .b(reg_out_B[0]) );
    inv_8 U27 ( .x(___cell__39620_net143983), .a(Imm[15]) );
    nand2i_2 U270 ( .x(n3461), .a(n1563), .b(n874) );
    nand2_0 U2700 ( .x(n1568), .a(reg_out_B[0]), .b(IR_function_field[0]) );
    nor2i_0 U2701 ( .x(n2001), .a(reg_out_B[0]), .b(n1524) );
    nand2i_0 U2702 ( .x(n1659), .a(reg_out_B[0]), .b(n645) );
    nand2_0 U2703 ( .x(n3257), .a(IR_function_field[3]), .b(IR_function_field
        [1]) );
    or3i_2 U2704 ( .x(n1538), .a(IR_function_field[2]), .b(IR_function_field
        [4]), .c(IR_function_field[3]) );
    nand2_0 U2705 ( .x(n2588), .a(Imm[24]), .b(n541) );
    exnor2_1 U2706 ( .x(n1486), .a(n541), .b(Imm[24]) );
    aoi21_1 U2707 ( .x(n1104), .a(n852), .b(n530), .c(n1064) );
    nor2i_3 U2708 ( .x(n1092), .a(n852), .b(n1093) );
    nor2i_3 U2709 ( .x(n1119), .a(n852), .b(n1120) );
    nand2i_2 U271 ( .x(n3494), .a(n1654), .b(n1689) );
    nor2i_3 U2710 ( .x(n1088), .a(n852), .b(n695) );
    nor2i_3 U2711 ( .x(n1121), .a(n852), .b(n1122) );
    exnor2_1 U2712 ( .x(n1461), .a(n4146), .b(n852) );
    inv_2 U2713 ( .x(n1655), .a(reg_out_A[7]) );
    exnor2_1 U2714 ( .x(n1462), .a(Imm[7]), .b(n852) );
    nand2_0 U2715 ( .x(n2068), .a(n852), .b(Imm[7]) );
    ao21_6 U2716 ( .x(n3741), .a(n861), .b(n835), .c(n1728) );
    nand2i_2 U2717 ( .x(n3645), .a(n925), .b(n887) );
    nand2i_2 U2718 ( .x(n3637), .a(n925), .b(n628) );
    nand2i_2 U2719 ( .x(n3654), .a(n925), .b(n686) );
    and2_3 U272 ( .x(n506), .a(n3494), .b(n3495) );
    nand2i_2 U2720 ( .x(n3588), .a(n925), .b(n894) );
    nand2i_2 U2721 ( .x(n3626), .a(n925), .b(n749) );
    nand2i_2 U2722 ( .x(n3664), .a(n925), .b(n914) );
    nand2i_4 U2723 ( .x(n3577), .a(n925), .b(n609) );
    nand2i_2 U2724 ( .x(n3589), .a(n925), .b(n908) );
    oai21_2 U2725 ( .x(n1834), .a(n1646), .b(n890), .c(n1835) );
    aoi22_1 U2726 ( .x(n2907), .a(reg_out_B[18]), .b(n1064), .c(n633), .d(
        ___cell__39620_net145617) );
    inv_0 U2727 ( .x(n1851), .a(reg_out_B[18]) );
    exnor2_1 U2728 ( .x(n1500), .a(n910), .b(reg_out_B[18]) );
    aoi22_1 U2729 ( .x(n2805), .a(___cell__39620_net144517), .b(n2806), .c(
        n1391), .d(n2045) );
    and2_3 U273 ( .x(n509), .a(n3490), .b(n3491) );
    aoi21_1 U2731 ( .x(n3213), .a(n3219), .b(n1267), .c(n3215) );
    inv_0 U2732 ( .x(n1532), .a(n4147) );
    exnor2_1 U2733 ( .x(n1457), .a(n4147), .b(n904) );
    aoi22_1 U2734 ( .x(n2873), .a(___cell__39620_net143722), .b(n2874), .c(
        ___cell__39620_net143864), .d(n4129) );
    inv_0 U2736 ( .x(___cell__39620_net143694), .a(net149628) );
    nor2i_0 U2737 ( .x(n1227), .a(net149628), .b(___cell__39620_net143836) );
    exnor2_1 U2738 ( .x(n1460), .a(net149628), .b(n914) );
    nand2i_2 U2739 ( .x(n3488), .a(n1219), .b(n1685) );
    nand2_2 U274 ( .x(n2271), .a(n3308), .b(n3309) );
    nand2i_2 U2740 ( .x(n3566), .a(n1657), .b(n1685) );
    nand2i_2 U2741 ( .x(n3501), .a(n1647), .b(n1685) );
    nand2i_2 U2742 ( .x(n3487), .a(n1644), .b(n1685) );
    nand2i_2 U2743 ( .x(n3463), .a(___cell__39620_net144257), .b(n1685) );
    nand2i_1 U2744 ( .x(n3323), .a(n1587), .b(n1685) );
    nand2i_1 U2745 ( .x(n3472), .a(n1564), .b(n1685) );
    nand2i_1 U2746 ( .x(n3466), .a(n1580), .b(n1685) );
    nand2i_1 U2747 ( .x(n3543), .a(n1646), .b(n1685) );
    nand2i_2 U2748 ( .x(n3493), .a(n1655), .b(n1685) );
    nand2i_1 U2749 ( .x(n3469), .a(n1573), .b(n1685) );
    nand2i_2 U275 ( .x(n3387), .a(n1563), .b(n3584) );
    nand2i_1 U2750 ( .x(n3498), .a(n1654), .b(n1685) );
    nand2i_2 U2751 ( .x(n3396), .a(n1649), .b(n1685) );
    nand2i_2 U2752 ( .x(n3390), .a(n1656), .b(n1685) );
    nand2i_2 U2753 ( .x(n2729), .a(n1166), .b(n3856) );
    nand2i_4 U2754 ( .x(n995), .a(___cell__39620_net143287), .b(n3746) );
    inv_0 U2755 ( .x(net150830), .a(net149167) );
    inv_2 U2756 ( .x(n2177), .a(n2080) );
    nand2i_2 U2757 ( .x(n2355), .a(n1641), .b(n3760) );
    nand2_0 U2758 ( .x(n2018), .a(___cell__39620_net145617), .b(n4136) );
    nor2i_0 U2759 ( .x(n1212), .a(n4136), .b(___cell__39620_net143836) );
    inv_6 U276 ( .x(n3485), .a(n3483) );
    nor2i_0 U2760 ( .x(n1051), .a(n4136), .b(n1529) );
    exnor2_1 U2761 ( .x(n1458), .a(n904), .b(n4136) );
    inv_2 U2762 ( .x(n924), .a(n923) );
    oai22_2 U2763 ( .x(n2235), .a(n1649), .b(n889), .c(n1647), .d(n1651) );
    nand3i_0 U2764 ( .x(___cell__39620_net145419), .a(n2258), .b(
        ___cell__39620_net147791), .c(___cell__39620_net143326) );
    inv_0 U2765 ( .x(net150620), .a(net149120) );
    inv_16 U2766 ( .x(n893), .a(n892) );
    oai211_2 U2767 ( .x(n4057), .a(n996), .b(___cell__39620_net147731), .c(
        n998), .d(n997) );
    nand2_1 U2768 ( .x(n3578), .a(n923), .b(n524) );
    inv_5 U2769 ( .x(n843), .a(n1971) );
    oai21_5 U277 ( .x(n3483), .a(net151904), .b(n1806), .c(n3484) );
    inv_4 U2770 ( .x(n2754), .a(n2711) );
    nor2i_8 U2771 ( .x(n844), .a(n3647), .b(n610) );
    nand2i_8 U2772 ( .x(n1604), .a(n1605), .b(n1606) );
    inv_0 U2773 ( .x(net150405), .a(net149122) );
    inv_4 U2774 ( .x(n846), .a(n2570) );
    oai22_2 U2775 ( .x(n847), .a(n1570), .b(n1629), .c(n512), .d(n536) );
    inv_16 U2776 ( .x(n3627), .a(n1604) );
    nand2i_2 U2777 ( .x(n3667), .a(n1632), .b(n847) );
    inv_0 U2778 ( .x(n848), .a(n816) );
    nor2_0 U2779 ( .x(n1158), .a(n820), .b(n1160) );
    aoi22_2 U278 ( .x(n853), .a(n858), .b(n883), .c(n855), .d(n854) );
    nor2_1 U2780 ( .x(n1185), .a(n820), .b(n1186) );
    inv_5 U2781 ( .x(n1749), .a(N369) );
    nand2i_2 U2782 ( .x(n3554), .a(n1578), .b(n1689) );
    nand2i_2 U2783 ( .x(n3473), .a(n1644), .b(n1689) );
    nand2i_1 U2784 ( .x(n3347), .a(n1564), .b(n1689) );
    nand2i_1 U2785 ( .x(n3337), .a(n1580), .b(n1689) );
    nand2i_2 U2786 ( .x(n3563), .a(n1657), .b(n1689) );
    nand2i_1 U2787 ( .x(n3404), .a(n1649), .b(n1689) );
    nand2i_1 U2788 ( .x(n3540), .a(n1646), .b(n1689) );
    nand2i_1 U2789 ( .x(n3328), .a(n1587), .b(n1689) );
    inv_10 U279 ( .x(n2067), .a(n1040) );
    nand2i_1 U2790 ( .x(n3319), .a(n1573), .b(n1689) );
    nand2i_2 U2791 ( .x(n3308), .a(n1656), .b(n1689) );
    nand2i_1 U2792 ( .x(n3490), .a(n1655), .b(n1689) );
    nand2_2 U2793 ( .x(n2333), .a(N337), .b(n2837) );
    inv_0 U2794 ( .x(n857), .a(reg_out_B[3]) );
    inv_2 U2795 ( .x(n858), .a(n1584) );
    inv_4 U2796 ( .x(n2083), .a(n2184) );
    inv_2 U2797 ( .x(n3383), .a(n3382) );
    and3i_3 U2798 ( .x(n994), .a(n2325), .b(n2333), .c(n859) );
    inv_0 U2799 ( .x(n861), .a(n816) );
    inv_8 U28 ( .x(net151622), .a(___cell__39620_net143983) );
    nor2i_3 U280 ( .x(n1039), .a(n855), .b(n1040) );
    aoi222_1 U2800 ( .x(n2936), .a(n1191), .b(n2859), .c(n650), .d(n2899), .e(
        n1221), .f(n2902) );
    aoi22_1 U2801 ( .x(n2901), .a(n1221), .b(n2863), .c(n1191), .d(n2902) );
    or3i_5 U2802 ( .x(n2295), .a(n2296), .b(n2293), .c(n864) );
    ao21_3 U2803 ( .x(n864), .a(n1085), .b(n2290), .c(n2291) );
    inv_12 U2804 ( .x(n3629), .a(n3628) );
    oai21_1 U2805 ( .x(n866), .a(n1587), .b(n889), .c(n3786) );
    oai21_1 U2806 ( .x(n867), .a(n1587), .b(n546), .c(n3786) );
    inv_2 U2807 ( .x(n3788), .a(n3787) );
    mux2_4 U2808 ( .x(n868), .d0(n3358), .sl(n816), .d1(n3313) );
    nand2i_2 U2809 ( .x(n3920), .a(n1632), .b(n827) );
    nand2i_0 U281 ( .x(n3616), .a(n1578), .b(n896) );
    and4i_2 U2810 ( .x(n2117), .a(n2116), .b(n2118), .c(n2119), .d(n2120) );
    oa211_5 U2811 ( .x(n869), .a(n844), .b(n4005), .c(n2632), .d(n3838) );
    inv_5 U2812 ( .x(n2107), .a(n870) );
    inv_14 U2813 ( .x(n872), .a(n874) );
    aoi221_1 U2814 ( .x(n2793), .a(n842), .b(n502), .c(
        ___cell__39620_net143722), .d(n2798), .e(n1266) );
    aoi21_3 U2815 ( .x(n2675), .a(n2676), .b(n2677), .c(n2634) );
    oa22_4 U2816 ( .x(n2267), .a(n1730), .b(n877), .c(n1175), .d(n876) );
    inv_0 U2817 ( .x(n876), .a(n904) );
    inv_0 U2818 ( .x(n877), .a(n919) );
    nand2i_3 U2819 ( .x(n1730), .a(n1565), .b(n1689) );
    nand2_2 U282 ( .x(n3556), .a(n1040), .b(n3616) );
    inv_16 U2820 ( .x(n881), .a(n1643) );
    nand2i_2 U2821 ( .x(n3969), .a(n1634), .b(n525) );
    buf_1 U2822 ( .x(n919), .a(n931) );
    oaoi211_1 U2823 ( .x(n2606), .a(n2607), .b(n1700), .c(n541), .d(n2604) );
    oai21_1 U2824 ( .x(n2288), .a(n3737), .b(n1700), .c(reg_out_A[31]) );
    oai21_1 U2825 ( .x(n2486), .a(n3792), .b(n1700), .c(n537) );
    aoi21_1 U2826 ( .x(n3144), .a(n901), .b(n1700), .c(n1404) );
    aoi222_1 U2827 ( .x(n3053), .a(n1204), .b(n3056), .c(n644), .d(n1700), .e(
        ALU_result[14]), .f(n3057) );
    aoi21_1 U2828 ( .x(n2799), .a(n749), .b(n1700), .c(n1269) );
    oai21_1 U2829 ( .x(n2656), .a(n3841), .b(n1700), .c(n636) );
    inv_2 U283 ( .x(n3492), .a(n3647) );
    oai21_1 U2830 ( .x(n2530), .a(n3805), .b(n1700), .c(n540) );
    aoi21_1 U2831 ( .x(n3014), .a(n609), .b(n1700), .c(n1347) );
    aoi21_1 U2832 ( .x(n2978), .a(n893), .b(n1700), .c(n1328) );
    oai21_1 U2833 ( .x(n2697), .a(n3848), .b(n1700), .c(n686) );
    aoi21_1 U2834 ( .x(n2254), .a(n834), .b(n1700), .c(n1145) );
    aoi21_1 U2835 ( .x(n2105), .a(n852), .b(n1700), .c(n1107) );
    nand2i_1 U2836 ( .x(n2032), .a(n1529), .b(n1700) );
    aoi21_1 U2837 ( .x(n2063), .a(n914), .b(n1700), .c(n1086) );
    aoi21_1 U2838 ( .x(n2154), .a(n838), .b(n1700), .c(n1118) );
    inv_16 U2839 ( .x(n888), .a(n1652) );
    buf_3 U284 ( .x(n687), .a(reg_out_A[22]) );
    inv_16 U2840 ( .x(n891), .a(n1602) );
    buf_16 U2841 ( .x(n922), .a(n937) );
    exnor2_1 U2842 ( .x(n1492), .a(n628), .b(Imm[21]) );
    nand2_0 U2843 ( .x(n2720), .a(Imm[21]), .b(n628) );
    inv_0 U2844 ( .x(___cell__39620_net144765), .a(Imm[21]) );
    inv_16 U2845 ( .x(n894), .a(n1579) );
    nand2i_4 U2846 ( .x(n1652), .a(n891), .b(n531) );
    nand2_0 U2847 ( .x(___cell__39620_net146131), .a(n631), .b(n893) );
    exnor2_1 U2848 ( .x(n1504), .a(n893), .b(n631) );
    inv_0 U2849 ( .x(n898), .a(n904) );
    nand2i_2 U285 ( .x(n2605), .a(n1485), .b(n2139) );
    exnor2_1 U2850 ( .x(n1507), .a(net156363), .b(n644) );
    nand2_0 U2851 ( .x(n3023), .a(net156363), .b(n644) );
    inv_14 U2852 ( .x(n917), .a(n916) );
    inv_16 U2853 ( .x(n904), .a(n903) );
    nand2i_2 U2854 ( .x(n3354), .a(n1585), .b(n839) );
    nand2i_2 U2855 ( .x(n3555), .a(n1648), .b(n839) );
    nand2i_2 U2856 ( .x(n3564), .a(n862), .b(n839) );
    nand2i_2 U2857 ( .x(n3309), .a(n1561), .b(n839) );
    nand2i_2 U2858 ( .x(n3348), .a(n1563), .b(n839) );
    nand2i_2 U2859 ( .x(n3500), .a(n1577), .b(n839) );
    oai221_1 U286 ( .x(n3523), .a(n1302), .b(n1043), .c(n3524), .d(n4007), .e(
        n1806) );
    nand2i_2 U2860 ( .x(n3405), .a(n748), .b(n839) );
    nand2i_2 U2861 ( .x(n3338), .a(n1579), .b(n839) );
    nand2i_2 U2862 ( .x(n3474), .a(n1570), .b(n839) );
    nand2i_2 U2863 ( .x(n3353), .a(n1571), .b(n839) );
    nand2i_2 U2864 ( .x(n3320), .a(n1572), .b(n839) );
    nand2i_2 U2865 ( .x(n3329), .a(n1586), .b(n839) );
    nand2i_2 U2866 ( .x(n3495), .a(n1583), .b(n839) );
    nand2i_2 U2867 ( .x(n3491), .a(n1584), .b(n839) );
    inv_16 U2868 ( .x(n910), .a(n909) );
    exnor2_1 U2869 ( .x(n1510), .a(reg_out_B[13]), .b(n919) );
    and2_3 U287 ( .x(n733), .a(IR_opcode_field[3]), .b(IR_opcode_field[2]) );
    nand2_1 U2870 ( .x(n2260), .a(n3573), .b(n919) );
    inv_2 U2871 ( .x(n1563), .a(n930) );
    buf_1 U2872 ( .x(n920), .a(n937) );
    inv_16 U2873 ( .x(n914), .a(n913) );
    inv_0 U2874 ( .x(n945), .a(reg_dst) );
    aoai211_3 U2875 ( .x(n4116), .a(n946), .b(n947), .c(reg_dst), .d(N3304) );
    exnor2_1 U2876 ( .x(n1509), .a(n629), .b(n919) );
    nor2i_0 U2877 ( .x(n3060), .a(n629), .b(n1563) );
    inv_0 U2878 ( .x(n1375), .a(n629) );
    exnor2_1 U2879 ( .x(n1511), .a(n682), .b(n894) );
    nand3_0 U288 ( .x(___cell__39620_net143836), .a(n733), .b(n1520), .c(
        ___cell__39620_net144355) );
    nor2i_0 U2880 ( .x(n1377), .a(n682), .b(n1579) );
    inv_6 U2881 ( .x(n916), .a(n4015) );
    inv_2 U2882 ( .x(n1037), .a(counter[1]) );
    inv_10 U2883 ( .x(n937), .a(n935) );
    mux2i_5 U2884 ( .x(n3172), .d0(n3531), .sl(net149120), .d1(n3446) );
    inv_10 U2885 ( .x(n3531), .a(n3530) );
    nand2_0 U2886 ( .x(n2112), .a(n838), .b(n642) );
    inv_0 U2887 ( .x(___cell__39620_net143735), .a(n642) );
    exnor2_1 U2888 ( .x(n1463), .a(n642), .b(n922) );
    inv_0 U2889 ( .x(n1208), .a(n818) );
    inv_5 U289 ( .x(n2079), .a(n1682) );
    nor2i_0 U2890 ( .x(n1406), .a(n818), .b(n1572) );
    exnor2_1 U2891 ( .x(n1516), .a(n818), .b(n908) );
    nand2i_0 U2892 ( .x(n1610), .a(IR_opcode_field[3]), .b(IR_opcode_field[2])
         );
    oai21_1 U2895 ( .x(n3238), .a(n1166), .b(n546), .c(n3239) );
    oai21_1 U2896 ( .x(n3787), .a(n1587), .b(n889), .c(n3786) );
    nand3i_3 U2897 ( .x(n4050), .a(n948), .b(n949), .c(n950) );
    oai211_4 U2898 ( .x(n4051), .a(n951), .b(___cell__39620_net147731), .c(
        n952), .d(n953) );
    oai211_3 U2899 ( .x(n4054), .a(n954), .b(___cell__39620_net147731), .c(
        n955), .d(n956) );
    inv_8 U29 ( .x(n684), .a(n683) );
    inv_4 U290 ( .x(n3202), .a(n695) );
    nand2_2 U2900 ( .x(n4065), .a(n972), .b(n973) );
    nand4_1 U2901 ( .x(n4074), .a(n983), .b(n984), .c(n985), .d(n986) );
    nand3i_3 U2902 ( .x(n4079), .a(n554), .b(n994), .c(n995) );
    nand2i_4 U2903 ( .x(n4073), .a(n1015), .b(n1016) );
    nand2_2 U2904 ( .x(n4066), .a(n1026), .b(n1027) );
    oai211_4 U2905 ( .x(n4064), .a(n1028), .b(___cell__39620_net143287), .c(
        n1029), .d(n1030) );
    oai211_3 U2906 ( .x(n4062), .a(n1031), .b(___cell__39620_net143287), .c(
        n1032), .d(n1033) );
    nor2i_5 U2907 ( .x(n1053), .a(n1054), .b(n1055) );
    nor2i_5 U2908 ( .x(n1068), .a(n1069), .b(n4004) );
    nor2_6 U2909 ( .x(n1097), .a(n947), .b(n1098) );
    and4i_4 U2910 ( .x(n957), .a(n1103), .b(n1100), .c(n1101), .d(n1102) );
    nor2i_5 U2911 ( .x(n1108), .a(n922), .b(n1089) );
    nor2i_5 U2912 ( .x(n1135), .a(n1136), .b(n4007) );
    and4i_4 U2913 ( .x(n1001), .a(n1141), .b(n1138), .c(n1139), .d(n1140) );
    and4i_4 U2914 ( .x(n1004), .a(n1173), .b(n1170), .c(n1171), .d(n1172) );
    nor2_6 U2915 ( .x(n1180), .a(n679), .b(n4037) );
    nor2i_5 U2916 ( .x(n1183), .a(N1959), .b(n1184) );
    nor2i_5 U2917 ( .x(n1187), .a(n590), .b(n1120) );
    nor2i_5 U2918 ( .x(n1193), .a(n541), .b(n1120) );
    nor2i_5 U2919 ( .x(n1194), .a(n541), .b(n1122) );
    oai22_1 U292 ( .x(n2564), .a(n1578), .b(n695), .c(n2565), .d(n1682) );
    nor2i_5 U2920 ( .x(n1195), .a(N1957), .b(n1184) );
    and4i_4 U2921 ( .x(n987), .a(n1202), .b(n1199), .c(n1200), .d(n1201) );
    aoi21_3 U2922 ( .x(n1015), .a(n1231), .b(n1232), .c(
        ___cell__39620_net147731) );
    nor2i_5 U2923 ( .x(n1251), .a(N1984), .b(___cell__39620_net143845) );
    nor2i_5 U2924 ( .x(n1293), .a(N2015), .b(n1169) );
    nor2_6 U2925 ( .x(n1305), .a(n947), .b(n1306) );
    nor2i_5 U2926 ( .x(n1307), .a(n1308), .b(n1166) );
    nor2i_5 U2927 ( .x(n1338), .a(n1339), .b(n1055) );
    and4i_4 U2928 ( .x(n969), .a(n1355), .b(n1352), .c(n1353), .d(n1354) );
    and4i_4 U2929 ( .x(n1031), .a(n1368), .b(n1365), .c(n1366), .d(n1367) );
    nand2i_5 U293 ( .x(n4012), .a(n1556), .b(reg_out_B[3]) );
    and4i_4 U2930 ( .x(n966), .a(n1386), .b(n1383), .c(n1384), .d(n1385) );
    nor2i_5 U2931 ( .x(n1433), .a(n1434), .b(___cell__39620_net143653) );
    nand2i_4 U2932 ( .x(n1541), .a(n1534), .b(n1542) );
    nand2i_4 U2933 ( .x(n1070), .a(reg_out_B[3]), .b(n815) );
    inv_6 U2935 ( .x(n1572), .a(n908) );
    nand3i_5 U2936 ( .x(n1169), .a(___cell__39620_net143653), .b(n810), .c(
        n1520) );
    nand2i_4 U2937 ( .x(___cell__39620_net144340), .a(n1610), .b(n4137) );
    or3i_5 U2938 ( .x(___cell__39620_net144343), .a(___cell__39620_net144344), 
        .b(net152465), .c(___cell__39620_net143653) );
    nand2i_4 U2939 ( .x(n1620), .a(n1621), .b(n676) );
    exnor2_1 U294 ( .x(n1484), .a(n590), .b(reg_out_B[25]) );
    nand2i_4 U2940 ( .x(n1627), .a(n1628), .b(n1543) );
    or2_8 U2942 ( .x(n1636), .a(n816), .b(n815) );
    inv_6 U2943 ( .x(n1098), .a(N1870) );
    inv_6 U2944 ( .x(n1736), .a(N1893) );
    oai21_5 U2945 ( .x(n1740), .a(n1642), .b(n1654), .c(n1741) );
    inv_6 U2946 ( .x(n1775), .a(N1658) );
    inv_6 U2947 ( .x(n1778), .a(N1823) );
    inv_6 U2948 ( .x(n1780), .a(N1856) );
    inv_6 U2949 ( .x(n1820), .a(N1752) );
    nand2_2 U295 ( .x(n2283), .a(n3499), .b(n3500) );
    oai21_4 U2950 ( .x(n1939), .a(n1531), .b(n1940), .c(n1447) );
    mux2i_3 U2951 ( .x(n4080), .d0(n4047), .sl(N3304), .d1(n1941) );
    mux2i_3 U2952 ( .x(n4048), .d0(n4046), .sl(N3304), .d1(n1942) );
    inv_6 U2953 ( .x(n1434), .a(N3024) );
    mux2i_3 U2954 ( .x(n1943), .d0(N3024), .sl(IR_opcode_field[0]), .d1(N3029)
         );
    mux2i_3 U2955 ( .x(n1944), .d0(n1945), .sl(IR_opcode_field[1]), .d1(n1946)
         );
    inv_6 U2956 ( .x(n1947), .a(N1392) );
    mux2i_3 U2957 ( .x(n1948), .d0(N1402), .sl(IR_function_field[0]), .d1(
        N1407) );
    nand2i_4 U2958 ( .x(___cell__39620_net144173), .a(IR_opcode_field[1]), .b(
        ___cell__39620_net145037) );
    nor2_5 U2959 ( .x(n1549), .a(n1956), .b(n1957) );
    inv_2 U296 ( .x(n2183), .a(n1713) );
    aoi22_3 U2960 ( .x(n1963), .a(n1964), .b(n1965), .c(n1330), .d(n1966) );
    nor2i_5 U2961 ( .x(n1575), .a(n1451), .b(___cell__39620_net144175) );
    nor2_6 U2962 ( .x(n1581), .a(___cell__39620_net144175), .b(n1451) );
    aoi22_3 U2963 ( .x(n1975), .a(n1964), .b(n1976), .c(n1330), .d(n1977) );
    nand4_1 U2964 ( .x(n1059), .a(n1989), .b(n1990), .c(n1986), .d(n1991) );
    oai22_3 U2965 ( .x(n2010), .a(n2011), .b(n1574), .c(n2012), .d(n1566) );
    and4i_4 U2966 ( .x(n962), .a(n2010), .b(n2013), .c(n2015), .d(n2016) );
    and4i_4 U2967 ( .x(n961), .a(n2020), .b(n2017), .c(n2018), .d(n2019) );
    nand4_1 U2968 ( .x(n1081), .a(n2040), .b(n2041), .c(n2039), .d(n2042) );
    nand2_2 U297 ( .x(n2284), .a(n3404), .b(n3405) );
    oai211_4 U2970 ( .x(n2056), .a(n580), .b(n621), .c(n2060), .d(n2061) );
    aoi211_5 U2971 ( .x(n2058), .a(n1204), .b(n2064), .c(n1084), .d(n2062) );
    nand2i_4 U2972 ( .x(n1676), .a(net149167), .b(net151904) );
    aoi211_4 U2973 ( .x(n2078), .a(n2079), .b(n2080), .c(n1088), .d(n1090) );
    nand4_1 U2974 ( .x(n2097), .a(n2100), .b(n2101), .c(n2102), .d(n2098) );
    oai21_5 U2975 ( .x(n2111), .a(n881), .b(n1644), .c(n2110) );
    ao221_4 U2976 ( .x(n2121), .a(n662), .b(n1993), .c(n1318), .d(n2043), .e(
        n1112) );
    oai211_3 U2977 ( .x(n2143), .a(n2012), .b(n1186), .c(n2144), .d(n2145) );
    nor2i_5 U2978 ( .x(n2162), .a(n2163), .b(n1982) );
    and4i_4 U2979 ( .x(n1126), .a(n2171), .b(n2173), .c(n2174), .d(n2175) );
    and2_3 U298 ( .x(n507), .a(n3540), .b(n522) );
    aoi21_3 U2980 ( .x(n2180), .a(n1391), .b(n2181), .c(n1119) );
    and3i_3 U2981 ( .x(n955), .a(n2198), .b(n2200), .c(n2201) );
    and3i_3 U2982 ( .x(n2202), .a(n2205), .b(n2203), .c(n2204) );
    aoi21_3 U2983 ( .x(n2220), .a(n1318), .b(n2168), .c(n1137) );
    nand4_1 U2984 ( .x(n1141), .a(n2219), .b(n2217), .c(n2221), .d(n2220) );
    aoi21_3 U2985 ( .x(n2229), .a(n1066), .b(n2045), .c(n1133) );
    and3i_3 U2986 ( .x(n1002), .a(n2242), .b(n2244), .c(n2245) );
    nand4_1 U2987 ( .x(n2248), .a(n2249), .b(n2250), .c(n2251), .d(n2252) );
    nor2i_3 U2988 ( .x(n2245), .a(n2246), .b(n2253) );
    nand4_1 U2989 ( .x(n2253), .a(n2255), .b(n2256), .c(n2254), .d(n2257) );
    inv_14 U299 ( .x(n1689), .a(n1633) );
    nor2i_5 U2990 ( .x(___cell__39620_net145450), .a(n1683), .b(n1626) );
    aoi22_3 U2991 ( .x(n2301), .a(___cell__39620_net144517), .b(n2302), .c(
        n1391), .d(n2303) );
    nand4_1 U2992 ( .x(n2325), .a(___cell__39620_net145470), .b(n2326), .c(
        n2323), .d(n2317) );
    aoi21_3 U2993 ( .x(n2342), .a(n1177), .b(n1977), .c(n2067) );
    and4i_5 U2994 ( .x(n1170), .a(n1164), .b(n2350), .c(n2351), .d(n2346) );
    oai22_3 U2995 ( .x(n2358), .a(n2359), .b(n1588), .c(n2360), .d(n1574) );
    and4i_4 U2996 ( .x(n1006), .a(n2358), .b(n2361), .c(n2362), .d(n2363) );
    aoi21_3 U2998 ( .x(n2437), .a(n1066), .b(n2303), .c(n1187) );
    nand4_1 U2999 ( .x(n2443), .a(n2446), .b(n2447), .c(n2448), .d(n2449) );
    buf_10 U3 ( .x(net149121), .a(net149107) );
    inv_2 U30 ( .x(net156024), .a(Imm[17]) );
    nand4_1 U3000 ( .x(n2450), .a(n2453), .b(n2452), .c(n2451), .d(n2454) );
    nor3_4 U3001 ( .x(n1008), .a(n2450), .b(n2442), .c(n2438) );
    nand2_5 U3002 ( .x(n2459), .a(n1267), .b(___cell__39620_net144345) );
    oai221_3 U3003 ( .x(n2463), .a(___cell__39620_net143872), .b(n1764), .c(
        ___cell__39620_net143660), .d(n1765), .e(n2464) );
    oai211_3 U3004 ( .x(n2466), .a(n553), .b(n1055), .c(n2467), .d(n2468) );
    nand4_1 U3005 ( .x(n1202), .a(n2469), .b(n2470), .c(n2471), .d(n2472) );
    aoi21_3 U3006 ( .x(n2480), .a(n1066), .b(n2375), .c(n1193) );
    nand4i_4 U3007 ( .x(n2497), .a(n1203), .b(n2498), .c(n2500), .d(n2501) );
    and4i_4 U3008 ( .x(n2504), .a(n2507), .b(n2505), .c(n2506), .d(n2503) );
    aoi22_3 U3009 ( .x(n2519), .a(n2079), .b(n2262), .c(n1391), .d(n2520) );
    inv_5 U301 ( .x(n1219), .a(reg_out_A[25]) );
    aoi21_3 U3010 ( .x(n2522), .a(___cell__39620_net144517), .b(n2303), .c(
        n2521) );
    and4i_4 U3011 ( .x(n1012), .a(n2527), .b(n2533), .c(n2534), .d(n2531) );
    and4i_4 U3012 ( .x(n1011), .a(n2538), .b(n2535), .c(n2536), .d(n2537) );
    nor2i_5 U3013 ( .x(n2535), .a(n2539), .b(n1210) );
    and4i_4 U3014 ( .x(n2577), .a(n2575), .b(n2567), .c(n2569), .d(n2573) );
    and3i_3 U3015 ( .x(n983), .a(n2579), .b(n2578), .c(n2577) );
    nor3i_5 U3016 ( .x(n2578), .a(n2585), .b(n1223), .c(n1225) );
    nand2_5 U3017 ( .x(n2589), .a(n2590), .b(n2591) );
    nand3i_3 U3018 ( .x(n2598), .a(n1229), .b(n2601), .c(n2599) );
    oai211_3 U3019 ( .x(n2610), .a(n2611), .b(n1186), .c(n2606), .d(n2608) );
    nand2_6 U302 ( .x(n1091), .a(n1686), .b(n1683) );
    aoi21_3 U3020 ( .x(n2612), .a(n1191), .b(n2532), .c(n2613) );
    and3i_3 U3021 ( .x(n2616), .a(n2619), .b(n2621), .c(n2622) );
    aoi21_3 U3022 ( .x(n2623), .a(___cell__39620_net143722), .b(n2624), .c(
        n1233) );
    nand4_1 U3023 ( .x(n2636), .a(n2637), .b(n2638), .c(n2639), .d(n2635) );
    oai211_3 U3024 ( .x(n2643), .a(n869), .b(n1166), .c(n2644), .d(n2645) );
    and3i_4 U3025 ( .x(n1238), .a(n2643), .b(n2646), .c(n2647) );
    aoi22_4 U3026 ( .x(n2648), .a(n1683), .b(n2375), .c(
        ___cell__39620_net144517), .d(n2649) );
    aoi21_6 U3027 ( .x(n2682), .a(n2674), .b(___cell__39620_net147791), .c(
        n1241) );
    nand4_1 U3028 ( .x(n1247), .a(n2685), .b(n2686), .c(n2687), .d(n2688) );
    oai211_3 U3029 ( .x(n2695), .a(n2696), .b(n1566), .c(n2692), .d(n2697) );
    oai22_1 U303 ( .x(n2521), .a(n1529), .b(n1091), .c(n1219), .d(n695) );
    and4i_4 U3030 ( .x(n2700), .a(n2695), .b(n2701), .c(n2702), .d(n2698) );
    nand4_1 U3031 ( .x(n2705), .a(n2715), .b(n2716), .c(n2717), .d(n2712) );
    aoi22_4 U3032 ( .x(n2740), .a(n2139), .b(n2741), .c(n2193), .d(n2742) );
    oai22_3 U3033 ( .x(n2745), .a(n2696), .b(n1574), .c(n2746), .d(n1566) );
    oai22_3 U3034 ( .x(n2748), .a(n1143), .b(n1816), .c(n2655), .d(n1588) );
    and3i_3 U3035 ( .x(n2751), .a(n2753), .b(n2757), .c(n2758) );
    and4i_4 U3036 ( .x(n2768), .a(n2772), .b(n2769), .c(n2770), .d(n2771) );
    oai22_3 U3037 ( .x(n2791), .a(___cell__39620_net143693), .b(
        ___cell__39620_net144781), .c(n2696), .d(n1588) );
    nor3_4 U3038 ( .x(n2792), .a(n2791), .b(n2788), .c(n2789) );
    nand4_1 U3039 ( .x(n2795), .a(n2799), .b(n2800), .c(n2801), .d(n2796) );
    inv_5 U304 ( .x(n1528), .a(n1525) );
    aoi21_6 U3040 ( .x(n2810), .a(n1177), .b(n1969), .c(n1836) );
    nand4_1 U3041 ( .x(n1277), .a(n2813), .b(n2815), .c(n2816), .d(n2814) );
    aoi221_4 U3042 ( .x(n2817), .a(n1095), .b(n1423), .c(n1197), .d(n1165), 
        .e(n1273) );
    nand4_3 U3043 ( .x(n1276), .a(n2817), .b(n2818), .c(n2819), .d(n2820) );
    oai211_4 U3044 ( .x(n2821), .a(n2822), .b(n1626), .c(n2823), .d(n2824) );
    nand4_3 U3045 ( .x(n2830), .a(n2831), .b(n2832), .c(n2828), .d(n2833) );
    nor3_4 U3046 ( .x(n952), .a(n2821), .b(n2830), .c(n2825) );
    and3i_3 U3048 ( .x(n2896), .a(n2893), .b(n2891), .c(n2897) );
    and3i_3 U3049 ( .x(n2903), .a(n2898), .b(n2901), .c(n2904) );
    nand2i_0 U305 ( .x(n2460), .a(reg_out_B[4]), .b(n1964) );
    and4i_4 U3050 ( .x(n2918), .a(n1317), .b(n2917), .c(n2919), .d(n2914) );
    nand3i_3 U3051 ( .x(n2937), .a(n2931), .b(n2928), .c(n2936) );
    oai22_3 U3052 ( .x(n2942), .a(n2943), .b(n1658), .c(n2944), .d(n784) );
    ao21_4 U3053 ( .x(n2941), .a(n1085), .b(n2910), .c(n2945) );
    ao21_4 U3054 ( .x(n2961), .a(n1221), .b(n2859), .c(n2958) );
    nand4_1 U3055 ( .x(n2966), .a(n2967), .b(n2968), .c(n2965), .d(n2969) );
    and3i_3 U3056 ( .x(n973), .a(n2966), .b(n2962), .c(n2970) );
    nand2_5 U3057 ( .x(n2971), .a(n2972), .b(n2973) );
    and4i_4 U3058 ( .x(n2968), .a(n2971), .b(n2974), .c(n2975), .d(n2976) );
    and3i_4 U3059 ( .x(n2967), .a(n2977), .b(n2978), .c(n2979) );
    nor2i_3 U306 ( .x(n2458), .a(___cell__39620_net144331), .b(n1072) );
    and4i_5 U3060 ( .x(n1342), .a(n1338), .b(n2982), .c(n2983), .d(n2984) );
    nand3_3 U3061 ( .x(n3005), .a(n3002), .b(n2999), .c(n3003) );
    and4i_4 U3062 ( .x(n3015), .a(n3018), .b(n3016), .c(n3017), .d(n3014) );
    nand4_1 U3063 ( .x(n1355), .a(n3029), .b(n3030), .c(n3028), .d(n3031) );
    nand4i_4 U3064 ( .x(n3045), .a(n3037), .b(n3039), .c(n3044), .d(n3046) );
    nand4_1 U3065 ( .x(n3048), .a(n3052), .b(n3053), .c(n3049), .d(n3050) );
    nand4_1 U3066 ( .x(n1368), .a(n3064), .b(n3065), .c(n3066), .d(n3067) );
    aoi221_4 U3067 ( .x(n3074), .a(___cell__39620_net143864), .b(n3075), .c(
        ___cell__39620_net143722), .d(n3076), .e(n1372) );
    aoi221_4 U3068 ( .x(n3077), .a(n650), .b(n3041), .c(n649), .d(n3078), .e(
        n3079) );
    nor3_4 U3069 ( .x(n3082), .a(n3083), .b(n3084), .c(n3085) );
    nand2i_2 U307 ( .x(___cell__39620_net144200), .a(n1533), .b(
        IR_opcode_field[1]) );
    nand4i_4 U3071 ( .x(n3105), .a(n3099), .b(n3101), .c(n3104), .d(n3106) );
    nand4_1 U3072 ( .x(n1402), .a(n3123), .b(n3124), .c(n3122), .d(n3125) );
    and4i_4 U3073 ( .x(n1410), .a(n3149), .b(n3151), .c(n3148), .d(n3152) );
    oai22_3 U3074 ( .x(n3160), .a(n3130), .b(n1574), .c(n2011), .d(n1566) );
    ao21_4 U3075 ( .x(n3185), .a(n1066), .b(n3186), .c(n3182) );
    and4i_5 U3076 ( .x(n3192), .a(n1422), .b(n3193), .c(n3194), .d(n3191) );
    oai211_3 U3077 ( .x(n3203), .a(n3204), .b(n3180), .c(n3205), .d(n3206) );
    oai211_3 U3078 ( .x(n3208), .a(n2360), .b(n1186), .c(n3209), .d(n3210) );
    nor3_4 U3079 ( .x(n949), .a(n3203), .b(n3208), .c(n3207) );
    nand2_2 U308 ( .x(n3315), .a(n1040), .b(n3595) );
    nand4_1 U3080 ( .x(n3220), .a(n1514), .b(n1511), .c(n1516), .d(n1517) );
    nand4_1 U3081 ( .x(n3223), .a(n1497), .b(n1495), .c(n1501), .d(n1499) );
    nand4_1 U3082 ( .x(n3224), .a(n1490), .b(n1488), .c(n1494), .d(n1492) );
    nand4_1 U3083 ( .x(n3226), .a(n1481), .b(n1479), .c(n1486), .d(n1483) );
    nand4_1 U3084 ( .x(n3227), .a(n1473), .b(n1471), .c(n1477), .d(n1475) );
    nand4_1 U3085 ( .x(n3229), .a(n1465), .b(n1463), .c(n1469), .d(n1467) );
    nor3i_5 U3086 ( .x(n3246), .a(n3247), .b(n3242), .c(n1435) );
    nand3_3 U3087 ( .x(n1441), .a(n3246), .b(n3244), .c(n3248) );
    nand4_1 U3088 ( .x(n3261), .a(n1498), .b(n1496), .c(n1502), .d(n1500) );
    nand4_1 U3089 ( .x(n3262), .a(n1489), .b(n1487), .c(n1493), .d(n1491) );
    inv_2 U309 ( .x(n3595), .a(n651) );
    nand4_1 U3090 ( .x(n3264), .a(n1482), .b(n1480), .c(n1485), .d(n1484) );
    nand4_1 U3091 ( .x(n3272), .a(n1466), .b(n1464), .c(n1470), .d(n1468) );
    nand4_1 U3092 ( .x(n3273), .a(n1461), .b(n1459), .c(n3274), .d(n1457) );
    aoi211_4 U3093 ( .x(n3282), .a(n3283), .b(n2004), .c(n1449), .d(n3284) );
    nand2_5 U3094 ( .x(n3291), .a(n3292), .b(n3293) );
    ao211_5 U3095 ( .x(n1966), .a(reg_out_B[4]), .b(n3311), .c(n897), .d(n2067
        ) );
    oai22_5 U3096 ( .x(n3312), .a(n915), .b(n1654), .c(n1642), .d(n1655) );
    ao211_5 U3097 ( .x(n1969), .a(reg_out_B[4]), .b(n3315), .c(n3316), .d(
        n2067) );
    inv_5 U3098 ( .x(n3324), .a(n3321) );
    ao211_5 U3099 ( .x(n1977), .a(reg_out_B[4]), .b(n3325), .c(n3326), .d(
        n2067) );
    inv_2 U31 ( .x(n639), .a(n638) );
    nand2_2 U310 ( .x(n3351), .a(n1040), .b(n3596) );
    ao211_5 U3100 ( .x(n1069), .a(reg_out_B[4]), .b(n3332), .c(n3333), .d(
        n2067) );
    ao211_5 U3101 ( .x(n1965), .a(reg_out_B[4]), .b(n3343), .c(n3344), .d(
        n2067) );
    nand2i_4 U3102 ( .x(n1976), .a(n1973), .b(n3354) );
    nand2_5 U3103 ( .x(n2992), .a(n3370), .b(n3371) );
    oai22_5 U3104 ( .x(n2568), .a(n1573), .b(n1642), .c(
        ___cell__39620_net144257), .d(n915) );
    oai22_3 U3105 ( .x(n2306), .a(n509), .b(n536), .c(n1585), .d(n1629) );
    oai22_3 U3106 ( .x(n2373), .a(n3409), .b(n536), .c(n1571), .d(n1629) );
    oai211_4 U3107 ( .x(n3422), .a(n3423), .b(n1560), .c(n3424), .d(n3425) );
    oai22_3 U3108 ( .x(n2738), .a(n507), .b(reg_out_B[3]), .c(n1572), .d(n822)
         );
    oai22_3 U3109 ( .x(n2477), .a(n3406), .b(n536), .c(n1579), .d(n1629) );
    nand2i_2 U311 ( .x(n1157), .a(N69), .b(n1552) );
    oai22_5 U3111 ( .x(n2375), .a(n1571), .b(n871), .c(n3454), .d(n4125) );
    oai22_5 U3112 ( .x(n3457), .a(n1561), .b(n872), .c(net149167), .d(n3341)
         );
    oai22_3 U3113 ( .x(n3458), .a(n1529), .b(n872), .c(n3459), .d(n4125) );
    nand2i_4 U3114 ( .x(n3464), .a(n3465), .b(n3466) );
    nand2i_4 U3115 ( .x(n3467), .a(n3468), .b(n3469) );
    ao211_5 U3116 ( .x(n1349), .a(net151904), .b(n3477), .c(n547), .d(n1982)
         );
    ao211_5 U3117 ( .x(n1047), .a(net151904), .b(n3478), .c(n3322), .d(n1982)
         );
    ao211_5 U3118 ( .x(n1049), .a(net151904), .b(n3479), .c(n3468), .d(n1982)
         );
    ao211_5 U3119 ( .x(n1045), .a(net151904), .b(n3480), .c(n622), .d(n1982)
         );
    nor2i_0 U312 ( .x(n1156), .a(n855), .b(n1157) );
    ao211_5 U3120 ( .x(n1361), .a(net151904), .b(n3482), .c(n3471), .d(n1982)
         );
    nand2i_4 U3121 ( .x(n3496), .a(n3497), .b(n3498) );
    oai221_3 U3122 ( .x(n2167), .a(n3509), .b(n1607), .c(n891), .d(n3510), .e(
        n3511) );
    ao221_5 U3123 ( .x(n2165), .a(n1289), .b(n3537), .c(n3186), .d(n1602), .e(
        n1123) );
    ao221_5 U3124 ( .x(n2218), .a(n1289), .b(n3538), .c(n3539), .d(n1602), .e(
        n1135) );
    nand2i_4 U3125 ( .x(n3541), .a(n3542), .b(n3543) );
    oai22_5 U3126 ( .x(n3544), .a(n1572), .b(n880), .c(n822), .d(n1646) );
    ao211_5 U3127 ( .x(n3278), .a(reg_out_B[4]), .b(n3556), .c(n2067), .d(
        n3557) );
    ao211_5 U3128 ( .x(n1136), .a(net151904), .b(n3559), .c(n1982), .d(n3558)
         );
    nand2_5 U3129 ( .x(n3560), .a(n3561), .b(n3562) );
    nand2_2 U313 ( .x(n3783), .a(n3325), .b(n855) );
    oai22_5 U3130 ( .x(n2179), .a(n557), .b(n836), .c(n3489), .d(n4125) );
    nand2i_4 U3131 ( .x(n3570), .a(n1562), .b(n1728) );
    inv_5 U3132 ( .x(n3322), .a(n3574) );
    inv_5 U3133 ( .x(n3471), .a(n3578) );
    inv_5 U3134 ( .x(n3465), .a(n3588) );
    inv_5 U3135 ( .x(n3468), .a(n3589) );
    inv_5 U3136 ( .x(n3605), .a(n3495) );
    nand2i_4 U3138 ( .x(n1606), .a(net151904), .b(n1982) );
    inv_5 U3139 ( .x(n3389), .a(n3637) );
    nand2_2 U314 ( .x(n3332), .a(n1040), .b(n3615) );
    inv_5 U3140 ( .x(n3542), .a(n3657) );
    nand2i_4 U3142 ( .x(n3682), .a(n1655), .b(n883) );
    oai211_3 U3143 ( .x(n3683), .a(n1331), .b(n1546), .c(n2065), .d(n3682) );
    nand2_2 U3144 ( .x(n2100), .a(n2024), .b(n3669) );
    nand2i_4 U3146 ( .x(n3695), .a(n2114), .b(n3694) );
    nand4_1 U3147 ( .x(n999), .a(n2117), .b(n2122), .c(n3697), .d(n3696) );
    nand2i_4 U3148 ( .x(n2151), .a(n1626), .b(n3681) );
    nand2i_0 U315 ( .x(n3615), .a(n1580), .b(n896) );
    nand2i_4 U3150 ( .x(n3703), .a(n1561), .b(n2066) );
    nand2i_4 U3151 ( .x(n3704), .a(n1546), .b(n1965) );
    nand3_3 U3152 ( .x(n3176), .a(n3704), .b(n3703), .c(n2159) );
    inv_5 U3153 ( .x(n3436), .a(n3176) );
    oai22_5 U3154 ( .x(n3705), .a(n1660), .b(n1122), .c(n4001), .d(n1120) );
    nand3_3 U3155 ( .x(n3186), .a(n3707), .b(n3706), .c(n2162) );
    nand2i_4 U3156 ( .x(n2208), .a(n1626), .b(n3689) );
    nand3_3 U3157 ( .x(n3711), .a(n2229), .b(n3710), .c(n2228) );
    nand3_3 U3159 ( .x(n2371), .a(n2232), .b(n3712), .c(n2231) );
    nand2_2 U316 ( .x(n3802), .a(n3479), .b(___cell__39620_net144331) );
    nand2i_4 U3160 ( .x(n3713), .a(n748), .b(n2066) );
    nand2i_4 U3161 ( .x(n3714), .a(n1546), .b(n1069) );
    nand3_3 U3162 ( .x(n3715), .a(n3714), .b(n3713), .c(n2213) );
    inv_5 U3163 ( .x(n3430), .a(n3715) );
    nand2i_4 U3164 ( .x(n2250), .a(n1654), .b(___cell__39620_net145444) );
    nand4_3 U3166 ( .x(n3719), .a(n2282), .b(n3718), .c(n2281), .d(n3367) );
    oai21_4 U3167 ( .x(___cell__39620_net147270), .a(n3720), .b(n1451), .c(
        n2285) );
    nand2_5 U3168 ( .x(n2275), .a(n3573), .b(n894) );
    or3i_4 U3169 ( .x(___cell__39620_net145421), .a(___cell__39620_net147732), 
        .b(n1169), .c(n1726) );
    nand2_2 U317 ( .x(n3481), .a(n665), .b(n3625) );
    or3i_4 U3170 ( .x(___cell__39620_net145425), .a(___cell__39620_net143326), 
        .b(n1184), .c(n1727) );
    nand2_5 U3171 ( .x(n3392), .a(n1686), .b(n901) );
    aoai211_4 U3172 ( .x(___cell__39620_net145429), .a(n1545), .b(n3741), .c(
        n1158), .d(n619) );
    inv_5 U3173 ( .x(n3750), .a(n1740) );
    nand2i_4 U3174 ( .x(n3751), .a(n1560), .b(n3683) );
    nand3i_5 U3175 ( .x(n3752), .a(n1740), .b(n3751), .c(n2342) );
    nand4i_4 U3176 ( .x(n3755), .a(n1176), .b(n3750), .c(n2338), .d(n3416) );
    nand2i_4 U3177 ( .x(n2367), .a(n1657), .b(n3705) );
    inv_5 U3178 ( .x(n2439), .a(n3765) );
    nand3_3 U3179 ( .x(n2499), .a(n2431), .b(n3769), .c(n2430) );
    nand2_2 U318 ( .x(n3773), .a(n3481), .b(___cell__39620_net144331) );
    nand2i_4 U3180 ( .x(n3777), .a(n2460), .b(n1728) );
    nand2i_4 U3181 ( .x(n3781), .a(n4008), .b(n2279) );
    nand3_3 U3182 ( .x(n3785), .a(n2478), .b(n3784), .c(n2476) );
    nand3_3 U3183 ( .x(n3796), .a(n2519), .b(n3795), .c(n2522) );
    inv_5 U3184 ( .x(n1224), .a(n3796) );
    nand4_1 U3185 ( .x(n3800), .a(n2518), .b(n3797), .c(n3799), .d(n3798) );
    inv_5 U3186 ( .x(n1211), .a(n3800) );
    nand2i_4 U3187 ( .x(n3808), .a(n1626), .b(n867) );
    oai31_2 U3188 ( .x(n1014), .a(n2514), .b(n2508), .c(n1209), .d(
        ___cell__39620_net147732) );
    nand4_1 U3189 ( .x(n3816), .a(n3814), .b(n3813), .c(n3815), .d(n2561) );
    nand2_2 U319 ( .x(n3482), .a(n665), .b(n3636) );
    inv_5 U3190 ( .x(n2670), .a(n2624) );
    oai211_3 U3191 ( .x(n3830), .a(n3553), .b(n1623), .c(n3829), .d(n2648) );
    inv_5 U3192 ( .x(n2667), .a(n3830) );
    oai211_3 U3193 ( .x(n2714), .a(n3460), .b(n4010), .c(n3843), .d(n2691) );
    oai211_3 U3194 ( .x(n2713), .a(n3403), .b(n1635), .c(n3844), .d(n2689) );
    nand2i_4 U3195 ( .x(n2701), .a(n1574), .b(n3837) );
    oai211_3 U3196 ( .x(n2803), .a(n3553), .b(n1625), .c(n3851), .d(n2739) );
    nand2i_4 U3197 ( .x(n3521), .a(n891), .b(n3033) );
    nand2_5 U3198 ( .x(n2827), .a(n2805), .b(n3864) );
    nand2i_4 U3199 ( .x(n2831), .a(n1186), .b(n2192) );
    inv_5 U32 ( .x(n683), .a(Imm[19]) );
    nand2_2 U320 ( .x(n3763), .a(n3482), .b(___cell__39620_net144331) );
    nand2i_4 U3201 ( .x(n2876), .a(n1658), .b(n2802) );
    inv_5 U3203 ( .x(n2944), .a(n3897) );
    nand4_3 U3204 ( .x(n3902), .a(n3901), .b(n3900), .c(n3899), .d(n3898) );
    nand2i_4 U3205 ( .x(n2973), .a(n1626), .b(n2938) );
    nand2i_4 U3207 ( .x(n3944), .a(n1623), .b(n3560) );
    oai211_3 U3208 ( .x(n3110), .a(n630), .b(n718), .c(n3965), .d(n3068) );
    nand2i_2 U321 ( .x(n3438), .a(n1562), .b(n3613) );
    nand2i_4 U3210 ( .x(n3514), .a(n891), .b(n3547) );
    nand4i_4 U3211 ( .x(n3168), .a(n1390), .b(n3974), .c(n3976), .d(n3975) );
    nand2i_4 U3212 ( .x(n3977), .a(n1632), .b(n2994) );
    nand2_5 U3214 ( .x(n3288), .a(n3984), .b(n3175) );
    inv_5 U3215 ( .x(n3204), .a(n3288) );
    nand2_5 U3216 ( .x(n3214), .a(n3985), .b(n3195) );
    nand2i_4 U3217 ( .x(n3210), .a(n1574), .b(n3289) );
    nand4_1 U3218 ( .x(n3990), .a(n3232), .b(n3228), .c(n3225), .d(n3222) );
    nand2i_4 U3219 ( .x(n3991), .a(n1943), .b(___cell__39620_net144303) );
    inv_5 U322 ( .x(n2268), .a(n1730) );
    nand4_1 U3220 ( .x(n1950), .a(n3275), .b(n3271), .c(n3263), .d(n3260) );
    nand3i_3 U3221 ( .x(n3993), .a(n3257), .b(n3256), .c(n3994) );
    nand4_3 U3222 ( .x(n3995), .a(n3287), .b(n3290), .c(n3993), .d(n3282) );
    nand3i_3 U3223 ( .x(n1941), .a(___cell__39620_net144166), .b(n1533), .c(
        ___cell__39620_net143655) );
    inv_5 U3224 ( .x(n2104), .a(n3677) );
    mux2i_3 U3225 ( .x(n2661), .d0(n3383), .sl(n816), .d1(n3386) );
    mux2i_3 U3226 ( .x(n2707), .d0(n3380), .sl(n816), .d1(n3385) );
    mux2i_3 U3227 ( .x(n2797), .d0(n3529), .sl(net149122), .d1(n3534) );
    mux2i_3 U3228 ( .x(n2872), .d0(n3522), .sl(net149122), .d1(n3536) );
    mux2i_3 U3229 ( .x(n3170), .d0(n3515), .sl(net149122), .d1(n3518) );
    nand2_2 U323 ( .x(n1741), .a(n2268), .b(n887) );
    nand2i_4 U3230 ( .x(n1946), .a(IR_opcode_field[0]), .b(N3014) );
    ao221_5 U3232 ( .x(n4070), .a(N361), .b(n977), .c(___cell__39620_net147732
        ), .d(n978), .e(n979) );
    nand2_8 U3233 ( .x(n947), .a(___cell__39620_net144312), .b(
        ___cell__39620_net143655) );
    inv_8 U3234 ( .x(n944), .a(n947) );
    inv_10 U3235 ( .x(n3997), .a(n947) );
    nand2i_5 U3236 ( .x(n1455), .a(___cell__39620_net144175), .b(n3995) );
    nor2i_5 U3237 ( .x(n1439), .a(n1440), .b(n1441) );
    nand2i_5 U3238 ( .x(n950), .a(___cell__39620_net143287), .b(n3988) );
    nor3i_5 U3239 ( .x(n967), .a(n3107), .b(n3108), .c(n3105) );
    nand2i_2 U324 ( .x(n2353), .a(n1474), .b(n2139) );
    nor3i_5 U3240 ( .x(n970), .a(n3047), .b(n3048), .c(n3045) );
    and4i_5 U3241 ( .x(n1028), .a(n1345), .b(n1342), .c(n1343), .d(n1344) );
    nor3i_5 U3242 ( .x(n1029), .a(n3006), .b(n3005), .c(n3007) );
    nor3i_5 U3243 ( .x(n951), .a(n1275), .b(n1276), .c(n1277) );
    inv_16 U3244 ( .x(n977), .a(n1596) );
    and4i_5 U3245 ( .x(n980), .a(n2654), .b(n2653), .c(n2657), .d(n2659) );
    nor3i_5 U3246 ( .x(n958), .a(n2096), .b(n2094), .c(n2097) );
    and4i_5 U3247 ( .x(n960), .a(n1059), .b(n1056), .c(n1057), .d(n1058) );
    inv_16 U3248 ( .x(n3057), .a(n1087) );
    aoi21_4 U3249 ( .x(n3161), .a(n1221), .b(n3078), .c(n3158) );
    inv_2 U325 ( .x(n3270), .a(n1474) );
    inv_16 U3250 ( .x(n2837), .a(n1592) );
    nor3i_5 U3251 ( .x(n2881), .a(n2879), .b(n1304), .c(n2880) );
    oai221_5 U3252 ( .x(n2669), .a(n2670), .b(n703), .c(n1234), .d(n4001), .e(
        n2671) );
    oai22_4 U3253 ( .x(n2666), .a(n2667), .b(n784), .c(n2668), .d(
        ___cell__39620_net144406) );
    nand4_2 U3254 ( .x(n2508), .a(n2504), .b(n2509), .c(n2510), .d(n2511) );
    nor3i_5 U3255 ( .x(n1199), .a(n2465), .b(n2463), .c(n2466) );
    aoi21_4 U3256 ( .x(n1200), .a(n662), .b(n2384), .c(n1195) );
    nand2i_5 U3257 ( .x(n2362), .a(n1566), .b(n3752) );
    nand2i_5 U3258 ( .x(n3696), .a(n1694), .b(n3624) );
    oai22_6 U3259 ( .x(___cell__39620_net145444), .a(n784), .b(n696), .c(
        ___cell__39620_net144406), .d(n1093) );
    nor2i_1 U326 ( .x(n1179), .a(n534), .b(n4002) );
    inv_16 U3260 ( .x(n1267), .a(n1641) );
    inv_7 U3261 ( .x(n2360), .a(n2238) );
    nand2_8 U3262 ( .x(n1186), .a(n1581), .b(n1576) );
    inv_16 U3263 ( .x(n2024), .a(n670) );
    oai21_6 U3264 ( .x(n2826), .a(n816), .b(n1450), .c(n2808) );
    inv_10 U3265 ( .x(n3662), .a(n1184) );
    inv_10 U3266 ( .x(n3999), .a(n1184) );
    inv_16 U3267 ( .x(n3624), .a(n1169) );
    inv_16 U3268 ( .x(n1064), .a(n1143) );
    aoi222_4 U3269 ( .x(n3169), .a(n3170), .b(n1204), .c(n3171), .d(
        ___cell__39620_net143722), .e(n3172), .f(___cell__39620_net143864) );
    inv_4 U327 ( .x(n2206), .a(n3705) );
    inv_16 U3270 ( .x(n1221), .a(n1186) );
    oai221_5 U3271 ( .x(n3078), .a(n3614), .b(n4003), .c(n3611), .d(n1559), 
        .e(n3058) );
    nand2i_8 U3272 ( .x(n1588), .a(___cell__39620_net144175), .b(n1589) );
    oai221_5 U3273 ( .x(n2014), .a(n3623), .b(n4004), .c(n3620), .d(n1559), 
        .e(n1970) );
    nand2_8 U3274 ( .x(n1574), .a(n1575), .b(n1576) );
    nand2i_5 U3276 ( .x(n3121), .a(n1912), .b(n944) );
    oai221_5 U3277 ( .x(n3041), .a(n3433), .b(n1070), .c(n3600), .d(n1559), 
        .e(n3021) );
    nand2i_5 U3278 ( .x(n3099), .a(n1387), .b(n3100) );
    nand2i_5 U3279 ( .x(n3106), .a(n1588), .b(n3041) );
    nor2i_0 U328 ( .x(n2343), .a(n534), .b(n1654) );
    nand2i_5 U3280 ( .x(n1592), .a(___cell__39620_net144175), .b(n1593) );
    inv_16 U3281 ( .x(n1318), .a(n1055) );
    nand3i_5 U3282 ( .x(n3071), .a(n1369), .b(n3072), .c(n3073) );
    aoi22_4 U3283 ( .x(n3080), .a(n1221), .b(n3001), .c(n1191), .d(n3000) );
    nand2i_5 U3284 ( .x(n3037), .a(n1356), .b(n3038) );
    aoi22_4 U3285 ( .x(n3044), .a(n650), .b(n3000), .c(n1221), .d(n3004) );
    nand2i_5 U3286 ( .x(n2984), .a(n1879), .b(n3997) );
    and4i_5 U3287 ( .x(n2950), .a(n2949), .b(n2951), .c(n2948), .d(n2952) );
    nand2i_5 U3288 ( .x(n2964), .a(n1566), .b(n3001) );
    nand2i_6 U3289 ( .x(n2969), .a(n1868), .b(n977) );
    nor2i_1 U329 ( .x(n1163), .a(N1734), .b(___cell__39620_net143710) );
    inv_16 U3290 ( .x(n1197), .a(n1616) );
    nand4i_5 U3291 ( .x(n2846), .a(n1288), .b(n3868), .c(n3870), .d(n3869) );
    inv_16 U3292 ( .x(n4000), .a(n946) );
    nand2i_5 U3293 ( .x(n2885), .a(n1855), .b(n1987) );
    nand2i_5 U3294 ( .x(n2886), .a(n1854), .b(n3662) );
    nand3i_5 U3295 ( .x(n2893), .a(n1310), .b(n2894), .c(n2895) );
    oai211_5 U3296 ( .x(n2849), .a(n3629), .b(n1043), .c(n2765), .d(n3859) );
    nand2_8 U3297 ( .x(n1626), .a(n1436), .b(___cell__39620_net147732) );
    nand2i_6 U3298 ( .x(n2832), .a(n1574), .b(n3752) );
    nand2i_5 U3299 ( .x(n2833), .a(n1566), .b(n3289) );
    inv_2 U330 ( .x(n4002), .a(n766) );
    inv_16 U3300 ( .x(___cell__39620_net143722), .a(___cell__39620_net144406)
         );
    nand2_5 U3301 ( .x(n2757), .a(n513), .b(n502) );
    nand2_5 U3302 ( .x(n2758), .a(n2797), .b(n1267) );
    oai221_5 U3303 ( .x(n2557), .a(n1315), .b(n1043), .c(n3426), .d(n1072), 
        .e(n1806) );
    nand2i_5 U3304 ( .x(n2686), .a(n1166), .b(n2733) );
    ao222_5 U3305 ( .x(n2706), .a(n2707), .b(n2024), .c(n745), .d(
        ___cell__39620_net145617), .e(n2708), .f(n2022) );
    oai221_5 U3306 ( .x(n2532), .a(n3420), .b(n4003), .c(n1300), .d(n1565), 
        .e(n1807) );
    inv_16 U3307 ( .x(n1191), .a(n1588) );
    nand2_5 U3308 ( .x(n2664), .a(n2708), .b(n1267) );
    inv_6 U3309 ( .x(n1234), .a(n3821) );
    nand2_8 U3310 ( .x(n1658), .a(n1429), .b(___cell__39620_net147732) );
    nand2_8 U3311 ( .x(n4001), .a(n1429), .b(___cell__39620_net147732) );
    nand2i_8 U3312 ( .x(___cell__39620_net144406), .a(___cell__39620_net144175
        ), .b(n1650) );
    nand2i_5 U3313 ( .x(n2597), .a(n1795), .b(n3662) );
    nor2i_5 U3314 ( .x(n1225), .a(n1085), .b(n1211) );
    nand2i_5 U3315 ( .x(n2575), .a(n1220), .b(n2576) );
    nand2i_4 U3316 ( .x(n2539), .a(n784), .b(n3796) );
    oai22_6 U3317 ( .x(n2490), .a(n1637), .b(n1122), .c(n1626), .d(n1120) );
    aoai211_5 U3318 ( .x(n2528), .a(n1267), .b(n2570), .c(n3809), .d(
        ___cell__39620_net144345) );
    nand2i_5 U3319 ( .x(n2516), .a(n1779), .b(___cell__39620_net145508) );
    oai22_1 U332 ( .x(n2838), .a(n679), .b(n4026), .c(n1602), .d(n4002) );
    nand2i_5 U3320 ( .x(n2465), .a(n1767), .b(n3997) );
    nor2i_5 U3321 ( .x(n1203), .a(n1204), .b(n1205) );
    nand2i_5 U3322 ( .x(n2445), .a(n703), .b(n2391) );
    aoi22_4 U3323 ( .x(n2422), .a(n1318), .b(n2384), .c(n1095), .d(n2423) );
    aoi21_6 U3325 ( .x(n2368), .a(n2024), .b(n2371), .c(n1180) );
    nand2i_6 U3326 ( .x(n2370), .a(n1626), .b(n3711) );
    inv_6 U3327 ( .x(n2359), .a(n2192) );
    nand2i_6 U3328 ( .x(n2332), .a(n1658), .b(___cell__39620_net147278) );
    nand3i_5 U3329 ( .x(n1077), .a(n1614), .b(n810), .c(
        ___cell__39620_net144355) );
    exnor2_1 U333 ( .x(n1496), .a(n815), .b(n692) );
    aoi21_4 U3330 ( .x(n2246), .a(n2022), .b(n2247), .c(n2248) );
    nand2i_5 U3331 ( .x(n2171), .a(n1124), .b(n2172) );
    aoi22_4 U3332 ( .x(n2164), .a(n2161), .b(___cell__39620_net147791), .c(
        n1095), .d(n2165) );
    inv_16 U3333 ( .x(___cell__39620_net143864), .a(n784) );
    inv_16 U3334 ( .x(n1204), .a(n4001) );
    oai21_5 U3335 ( .x(n2103), .a(n703), .b(n2104), .c(n2105) );
    nand2i_4 U3336 ( .x(n2101), .a(n1626), .b(n2059) );
    aoi21_5 U3337 ( .x(n2098), .a(n502), .b(n2099), .c(n1106) );
    nand2i_4 U3338 ( .x(n2034), .a(n784), .b(n2064) );
    nor2i_1 U334 ( .x(n1284), .a(n1285), .b(n690) );
    aoi21_5 U3340 ( .x(n3195), .a(n1256), .b(n3196), .c(n3197) );
    nand2_8 U3341 ( .x(n1641), .a(n1428), .b(___cell__39620_net143326) );
    inv_16 U3342 ( .x(___cell__39620_net144345), .a(net149122) );
    inv_16 U3343 ( .x(n1657), .a(n917) );
    oai211_5 U3344 ( .x(n2238), .a(n3430), .b(n815), .c(n3431), .d(n3432) );
    inv_16 U3345 ( .x(n2139), .a(n1536) );
    inv_12 U3346 ( .x(___cell__39620_net147791), .a(___cell__39620_net143658)
         );
    and2_8 U3347 ( .x(n1422), .a(n1197), .b(n1423) );
    nand4i_5 U3348 ( .x(n1988), .a(n1041), .b(n3634), .c(n3633), .d(n3632) );
    inv_16 U3349 ( .x(n1095), .a(n1166) );
    inv_2 U335 ( .x(n1285), .a(n1495) );
    nand4i_5 U3350 ( .x(n1992), .a(n1048), .b(n3661), .c(n3660), .d(n3659) );
    inv_16 U3351 ( .x(n1987), .a(n1077) );
    nand2i_8 U3352 ( .x(n1143), .a(___cell__39620_net144175), .b(n1710) );
    nand2i_8 U3353 ( .x(___cell__39620_net143693), .a(n1618), .b(
        ___cell__39620_net143326) );
    oai211_4 U3354 ( .x(n2023), .a(n3452), .b(n1625), .c(n3590), .d(n1994) );
    inv_16 U3355 ( .x(n1085), .a(n703) );
    nand2i_5 U3356 ( .x(n4003), .a(reg_out_B[3]), .b(n815) );
    nand2i_4 U3357 ( .x(n4004), .a(reg_out_B[3]), .b(n815) );
    nand2i_8 U3358 ( .x(n1559), .a(n815), .b(reg_out_B[3]) );
    aoi22_4 U3359 ( .x(n3058), .a(n1971), .b(n3059), .c(n1330), .d(n1965) );
    exnor2_1 U336 ( .x(n1495), .a(n891), .b(n692) );
    aoi22_4 U3360 ( .x(n1970), .a(n1971), .b(n1972), .c(n1330), .d(n1069) );
    oai221_4 U3361 ( .x(n2054), .a(n3433), .b(n1559), .c(n3600), .d(n1562), 
        .e(n1967) );
    nand2i_8 U3362 ( .x(n1055), .a(___cell__39620_net144345), .b(
        ___cell__39620_net144347) );
    nand4i_5 U3363 ( .x(n1380), .a(n1348), .b(n3960), .c(n3959), .d(n3958) );
    oai221_4 U3365 ( .x(n3112), .a(n3355), .b(n1635), .c(n849), .d(n727), .e(
        n3070) );
    nand2i_5 U3366 ( .x(n3100), .a(n702), .b(n3076) );
    oai211_5 U3367 ( .x(n3075), .a(n3515), .b(___cell__39620_net144345), .c(
        n3972), .d(n3971) );
    oai221_5 U3368 ( .x(n3000), .a(n3439), .b(n4003), .c(n747), .d(n1559), .e(
        n2980) );
    nor2i_5 U3369 ( .x(n1332), .a(n1333), .b(n1334) );
    nand2i_2 U337 ( .x(n3757), .a(n2339), .b(n3756) );
    nand2i_5 U3370 ( .x(n3953), .a(n4007), .b(n3646) );
    oai211_4 U3371 ( .x(n3051), .a(n3452), .b(n4008), .c(n3957), .d(n3032) );
    nand2i_5 U3372 ( .x(n3072), .a(n702), .b(n3963) );
    nand2i_6 U3373 ( .x(n3073), .a(n4001), .b(n3040) );
    oai211_4 U3374 ( .x(n3076), .a(n3413), .b(n1451), .c(n3970), .d(n3969) );
    nand4i_5 U3375 ( .x(n3001), .a(n1321), .b(n3934), .c(n3933), .d(n3932) );
    nand2i_5 U3376 ( .x(n3936), .a(n1072), .b(n3628) );
    nand2i_6 U3377 ( .x(n3935), .a(n1607), .b(n3774) );
    nand4i_5 U3378 ( .x(n1339), .a(n1314), .b(n3909), .c(n3908), .d(n3907) );
    oai221_4 U3379 ( .x(n3054), .a(n3366), .b(n1632), .c(n511), .d(n1636), .e(
        n3035) );
    nand2_2 U338 ( .x(n2339), .a(n2340), .b(n2341) );
    nand2i_5 U3380 ( .x(n3038), .a(___cell__39620_net144406), .b(n3963) );
    oai211_5 U3381 ( .x(n3040), .a(n499), .b(___cell__39620_net144345), .c(
        n3961), .d(n3962) );
    nand4i_5 U3382 ( .x(n3004), .a(n1312), .b(n3906), .c(n3905), .d(n3904) );
    nand4i_5 U3383 ( .x(n1308), .a(n1301), .b(n3884), .c(n3883), .d(n3882) );
    ao22_6 U3385 ( .x(n2949), .a(n662), .b(n2846), .c(n1318), .d(n1308) );
    nand4i_5 U3386 ( .x(n2859), .a(n1286), .b(n3867), .c(n3866), .d(n3865) );
    aoi21_5 U3387 ( .x(n2917), .a(n662), .b(n2849), .c(n1316) );
    nor2i_5 U3388 ( .x(n1317), .a(n1318), .b(n1319) );
    nand2_8 U3389 ( .x(___cell__39620_net143653), .a(IR_opcode_field[1]), .b(
        IR_opcode_field[0]) );
    inv_4 U339 ( .x(n3341), .a(n3470) );
    nand2i_6 U3390 ( .x(n1616), .a(net149122), .b(___cell__39620_net143785) );
    nor2i_5 U3391 ( .x(n1288), .a(n1289), .b(n1290) );
    nand2i_5 U3392 ( .x(n3868), .a(n4006), .b(n3648) );
    nand2i_6 U3393 ( .x(n3870), .a(n4005), .b(n3646) );
    nand2i_8 U3394 ( .x(n1182), .a(___cell__39620_net144345), .b(
        ___cell__39620_net143785) );
    nand2i_6 U3395 ( .x(n1166), .a(net149120), .b(___cell__39620_net144347) );
    oai211_5 U3396 ( .x(n2863), .a(n3611), .b(n1565), .c(n3850), .d(n2718) );
    nand2i_6 U3397 ( .x(n2892), .a(n3889), .b(n1217) );
    oai211_5 U3399 ( .x(n2911), .a(n3460), .b(n4008), .c(n3876), .d(n2889) );
    inv_2 U34 ( .x(n596), .a(n886) );
    oai211_1 U340 ( .x(n2337), .a(n3341), .b(___cell__39620_net144317), .c(
        n3342), .d(n2163) );
    or2_8 U3400 ( .x(n4005), .a(n891), .b(net149167) );
    inv_16 U3401 ( .x(n2193), .a(n1116) );
    nand2i_6 U3402 ( .x(n2856), .a(n3875), .b(n1217) );
    oai211_5 U3403 ( .x(n2192), .a(n3436), .b(n815), .c(n3437), .d(n3438) );
    nand2i_6 U3404 ( .x(n3864), .a(net149120), .b(n1431) );
    nand2i_5 U3406 ( .x(n2769), .a(n1055), .b(n2733) );
    aoi21_5 U3407 ( .x(n2780), .a(n1714), .b(n2781), .c(n1258) );
    aoi21_4 U3408 ( .x(n2778), .a(n504), .b(n2779), .c(n1255) );
    inv_10 U3409 ( .x(n2746), .a(n2863) );
    nor2i_1 U341 ( .x(n1270), .a(N1700), .b(___cell__39620_net143660) );
    inv_10 U3410 ( .x(n1298), .a(n2902) );
    oai22_6 U3411 ( .x(n2723), .a(___cell__39620_net143710), .b(n1820), .c(
        ___cell__39620_net143658), .d(n2720) );
    nand2_5 U3412 ( .x(n2756), .a(n2710), .b(n2022) );
    nand2i_4 U3413 ( .x(n4006), .a(net149167), .b(n891) );
    nand2i_4 U3414 ( .x(n4007), .a(net149167), .b(n891) );
    nand2i_8 U3415 ( .x(n1806), .a(n4140), .b(net149167) );
    nand4_3 U3417 ( .x(n3835), .a(n3834), .b(n3833), .c(n3832), .d(n3831) );
    nor2i_8 U3418 ( .x(n1237), .a(N1853), .b(n946) );
    nand2_8 U3419 ( .x(n1807), .a(n1728), .b(reg_out_B[3]) );
    inv_2 U342 ( .x(n1272), .a(N1865) );
    inv_7 U3420 ( .x(n1429), .a(n1653) );
    nand2i_5 U3421 ( .x(n2601), .a(n1182), .b(n2473) );
    nand2i_5 U3422 ( .x(n2576), .a(n1588), .b(n3422) );
    oai21_5 U3423 ( .x(n2582), .a(n621), .b(n2583), .c(n2584) );
    oai211_5 U3424 ( .x(n2473), .a(n3427), .b(n1602), .c(n3428), .d(n3429) );
    oai21_6 U3425 ( .x(n2423), .a(n3421), .b(n4005), .c(n3572) );
    nand2_8 U3426 ( .x(n3571), .a(n1728), .b(n1565) );
    nand2i_8 U3427 ( .x(n1122), .a(n1635), .b(n883) );
    nand2i_8 U3428 ( .x(n1120), .a(n718), .b(n4130) );
    aoi21_6 U3429 ( .x(n2503), .a(N1757), .b(___cell__39620_net145150), .c(
        n1207) );
    nor2_1 U343 ( .x(n1271), .a(n947), .b(n1272) );
    nand2i_6 U3430 ( .x(n2513), .a(n1778), .b(n1987) );
    nor2i_8 U3431 ( .x(n1196), .a(n1197), .b(n1198) );
    nand2i_5 U3433 ( .x(n2446), .a(n1566), .b(n2492) );
    nor2i_8 U3434 ( .x(n1189), .a(N1858), .b(n946) );
    oai21_6 U3436 ( .x(n2319), .a(n694), .b(n3735), .c(n2301) );
    oai211_4 U3437 ( .x(n2168), .a(n891), .b(n3506), .c(n3507), .d(n3508) );
    inv_16 U3438 ( .x(n1646), .a(n692) );
    or2_8 U3439 ( .x(n4008), .a(n637), .b(net149120) );
    nor2i_1 U344 ( .x(n2811), .a(n891), .b(n1646) );
    nand2i_5 U3440 ( .x(n2256), .a(n670), .b(n3702) );
    oai211_5 U3441 ( .x(n2089), .a(n3439), .b(n1562), .c(n3440), .d(n3441) );
    nand2i_5 U3442 ( .x(n2172), .a(n1182), .b(n2043) );
    nand2i_6 U3443 ( .x(n2190), .a(n3709), .b(n1217) );
    nand4i_5 U3444 ( .x(n2090), .a(n1068), .b(n3672), .c(n3671), .d(n3670) );
    nand4i_5 U3445 ( .x(n1993), .a(n1044), .b(n3643), .c(n3642), .d(n3641) );
    nand4i_5 U3446 ( .x(n2043), .a(n1071), .b(n3675), .c(n3674), .d(n3673) );
    nand2i_5 U3447 ( .x(n2145), .a(n1588), .b(n2090) );
    nor2i_8 U3448 ( .x(n1096), .a(N1738), .b(___cell__39620_net143710) );
    nor2i_8 U3449 ( .x(n1099), .a(N1837), .b(n946) );
    inv_2 U345 ( .x(n1274), .a(N1799) );
    oai221_4 U3450 ( .x(n2093), .a(n3614), .b(n1559), .c(n3611), .d(n1562), 
        .e(n1963) );
    nand2_8 U3451 ( .x(n2060), .a(n3677), .b(___cell__39620_net143722) );
    nand2i_6 U3452 ( .x(n2061), .a(n1626), .b(n3583) );
    oai21_5 U3453 ( .x(n2062), .a(n784), .b(n870), .c(n2063) );
    nand2i_6 U3454 ( .x(n2009), .a(n1457), .b(n2139) );
    aoi21_5 U3455 ( .x(n3175), .a(n1256), .b(n3176), .c(n3177) );
    nand2i_8 U3456 ( .x(n1040), .a(n759), .b(n1553) );
    nand2i_6 U3457 ( .x(n1446), .a(n1535), .b(n1528) );
    aoi21_6 U3458 ( .x(n1430), .a(n694), .b(n1431), .c(n1432) );
    nand2i_6 U3459 ( .x(n1639), .a(n1640), .b(n676) );
    nor2_1 U346 ( .x(n1273), .a(n1077), .b(n1274) );
    oai211_5 U3460 ( .x(n3196), .a(n3345), .b(n1546), .c(n3349), .d(n3350) );
    inv_16 U3461 ( .x(n1643), .a(n4011) );
    inv_16 U3462 ( .x(n1066), .a(n4010) );
    inv_16 U3463 ( .x(n1714), .a(n1635) );
    nand2i_6 U3465 ( .x(n3538), .a(n501), .b(n3627) );
    nor2i_6 U3466 ( .x(n1041), .a(n1042), .b(n1043) );
    nand2i_5 U3467 ( .x(n3634), .a(n1608), .b(n3628) );
    nand2i_5 U3468 ( .x(n3633), .a(n4007), .b(n3538) );
    nand2i_6 U3469 ( .x(n3632), .a(n1607), .b(n2766) );
    nand3_4 U347 ( .x(n1165), .a(n3754), .b(n665), .c(n2344) );
    nor2i_6 U3470 ( .x(n1360), .a(n1361), .b(n4005) );
    nand2i_5 U3471 ( .x(n3967), .a(n4007), .b(n3537) );
    nand2i_6 U3472 ( .x(n3966), .a(n1607), .b(n2722) );
    nand2i_5 U3473 ( .x(n3651), .a(n1608), .b(n3646) );
    nand2i_6 U3474 ( .x(n3649), .a(n1607), .b(n3648) );
    nor2i_5 U3475 ( .x(n1390), .a(n1391), .b(n1392) );
    nand2i_5 U3476 ( .x(n3974), .a(n4010), .b(n4142) );
    nand2i_6 U3477 ( .x(n3976), .a(n4008), .b(n2181) );
    nand2i_6 U3478 ( .x(n1625), .a(n694), .b(n891) );
    inv_6 U3479 ( .x(n3515), .a(n3512) );
    nand2i_2 U348 ( .x(n2137), .a(n1064), .b(n3698) );
    nand2i_6 U3480 ( .x(n3622), .a(n3621), .b(n3598) );
    nand2i_6 U3481 ( .x(n1972), .a(n3585), .b(n3617) );
    nor2i_6 U3482 ( .x(n1348), .a(n1349), .b(n1043) );
    nand2i_5 U3483 ( .x(n3960), .a(n1608), .b(n3655) );
    nand2i_5 U3484 ( .x(n3959), .a(n4007), .b(n3658) );
    nand2i_6 U3485 ( .x(n3958), .a(n1607), .b(n2677) );
    nand2i_5 U3486 ( .x(n1701), .a(___cell__39620_net144175), .b(n1939) );
    nand2i_6 U3487 ( .x(n3022), .a(n3585), .b(n3801) );
    aoi22_4 U3488 ( .x(n3068), .a(n1066), .b(n2991), .c(n1391), .d(n3069) );
    nand2i_6 U3489 ( .x(n3972), .a(n4008), .b(n2927) );
    nor2i_1 U349 ( .x(n2108), .a(n1451), .b(___cell__39620_net144406) );
    nand2i_5 U3490 ( .x(n3971), .a(n4010), .b(n3560) );
    aoi21_5 U3491 ( .x(n2980), .a(n1971), .b(n2981), .c(n1329) );
    nand2i_6 U3492 ( .x(n1608), .a(n891), .b(net149167) );
    nand2i_6 U3493 ( .x(n3790), .a(n751), .b(n3789) );
    nor2i_5 U3494 ( .x(n1321), .a(n1177), .b(n1322) );
    nand2i_5 U3495 ( .x(n3934), .a(n1070), .b(n3619) );
    nand2i_6 U3496 ( .x(n3932), .a(n1562), .b(n2763) );
    inv_16 U3497 ( .x(n1147), .a(n1608) );
    nand2i_6 U3498 ( .x(n3774), .a(n751), .b(n3773) );
    nor2i_8 U3499 ( .x(n1314), .a(n1147), .b(n1315) );
    inv_5 U35 ( .x(n640), .a(n638) );
    nor2_1 U350 ( .x(n2109), .a(n784), .b(n694) );
    nand2i_6 U3500 ( .x(n3909), .a(n4005), .b(n3537) );
    nand2i_5 U3501 ( .x(n3908), .a(n4006), .b(n3638) );
    nand2i_6 U3502 ( .x(n3907), .a(n1607), .b(n3764) );
    nand2i_6 U3503 ( .x(n3962), .a(n4008), .b(n2783) );
    nor2i_5 U3504 ( .x(n1312), .a(n1177), .b(n1313) );
    nor2i_5 U3505 ( .x(n1301), .a(n1147), .b(n1302) );
    nand2i_5 U3506 ( .x(n3883), .a(n1072), .b(n3655) );
    nand2i_6 U3507 ( .x(n3882), .a(n1607), .b(n3744) );
    nor2i_5 U3508 ( .x(n1299), .a(n1177), .b(n1300) );
    nand2i_6 U3509 ( .x(n3880), .a(n1565), .b(n3602) );
    aoi222_1 U351 ( .x(n2134), .a(n2109), .b(n2135), .c(n2108), .d(n2136), .e(
        reg_out_B[6]), .f(n2137) );
    nand2i_6 U3510 ( .x(n3879), .a(n1562), .b(n2673) );
    nand2i_6 U3511 ( .x(n2998), .a(n1505), .b(n2139) );
    nor2i_5 U3512 ( .x(n1286), .a(n1177), .b(n1287) );
    nand2i_5 U3513 ( .x(n3867), .a(n1070), .b(n685) );
    nand2i_6 U3514 ( .x(n2960), .a(n1503), .b(n2139) );
    oai211_4 U3515 ( .x(n3897), .a(n3553), .b(n4008), .c(n3896), .d(n2926) );
    nand2i_5 U3516 ( .x(n2972), .a(n670), .b(n3902) );
    nand2i_5 U3517 ( .x(n3877), .a(n1634), .b(n3020) );
    nand2i_6 U3518 ( .x(n2935), .a(n1502), .b(n2139) );
    oai211_5 U3519 ( .x(n3887), .a(n3522), .b(___cell__39620_net144345), .c(
        n3886), .d(n3885) );
    aoi21_1 U352 ( .x(n2138), .a(n2139), .b(n2140), .c(n1114) );
    nand2i_6 U3520 ( .x(n3913), .a(n1417), .b(n530) );
    nand2i_5 U3521 ( .x(n3857), .a(n4004), .b(n1972) );
    nand2i_5 U3522 ( .x(n2915), .a(n1861), .b(___cell__39620_net145150) );
    aoi21_5 U3523 ( .x(n2718), .a(n1177), .b(n2719), .c(n2630) );
    inv_6 U3525 ( .x(n3529), .a(n3526) );
    nand2i_6 U3526 ( .x(n3872), .a(n4008), .b(n3069) );
    aoi22_4 U3527 ( .x(n2889), .a(n1391), .b(n2890), .c(n1066), .d(n2783) );
    nand2i_6 U3528 ( .x(n2766), .a(n751), .b(n3631) );
    nand2_8 U3529 ( .x(n1623), .a(n694), .b(n891) );
    inv_2 U353 ( .x(n2140), .a(n1464) );
    nand2i_5 U3530 ( .x(n3845), .a(n1070), .b(n3022) );
    nand2i_6 U3531 ( .x(n3537), .a(n3565), .b(n3627) );
    nand2i_6 U3532 ( .x(n3756), .a(n816), .b(n3755) );
    nand2i_5 U3533 ( .x(n3437), .a(n1070), .b(n1966) );
    inv_16 U3534 ( .x(___cell__39620_net144517), .a(___cell__39620_net144374)
         );
    inv_16 U3536 ( .x(n1391), .a(n1623) );
    nand4i_5 U3537 ( .x(n1431), .a(n1282), .b(n3861), .c(n2804), .d(n3863) );
    oai21_5 U3538 ( .x(n3365), .a(n3366), .b(n815), .c(n3367) );
    oai21_6 U3539 ( .x(n2781), .a(n2429), .b(n536), .c(n3400) );
    exnor2_1 U354 ( .x(n1464), .a(reg_out_B[6]), .b(n922) );
    nor2i_5 U3540 ( .x(n1258), .a(n1249), .b(n1259) );
    nor2i_8 U3541 ( .x(n1255), .a(n1256), .b(n1257) );
    aoi22_4 U3542 ( .x(n2782), .a(n1391), .b(n2783), .c(n1066), .d(n2784) );
    aoi21_4 U3544 ( .x(n2721), .a(n2676), .b(n2722), .c(n2634) );
    nand2i_5 U3545 ( .x(n3855), .a(n1608), .b(n3764) );
    nand2i_5 U3546 ( .x(n3846), .a(n1608), .b(n3744) );
    nand2i_6 U3547 ( .x(n2744), .a(n1816), .b(n530) );
    aoi21_4 U3548 ( .x(n2632), .a(n1147), .b(n2633), .c(n2634) );
    nand2i_5 U3549 ( .x(n3838), .a(n4007), .b(n3790) );
    nor2i_1 U355 ( .x(n1114), .a(n1115), .b(n690) );
    nand2_4 U3550 ( .x(n3834), .a(n504), .b(n2373) );
    nand2i_6 U3552 ( .x(n2673), .a(n3585), .b(n3742) );
    nand2i_6 U3553 ( .x(n2763), .a(n3585), .b(n3772) );
    nand2i_6 U3554 ( .x(n2719), .a(n3585), .b(n3762) );
    nand2i_6 U3555 ( .x(n3840), .a(n1797), .b(n530) );
    nand2i_5 U3556 ( .x(n2591), .a(n2588), .b(___cell__39620_net147791) );
    nand2_3 U3557 ( .x(n3814), .a(n1714), .b(n2373) );
    nand2i_8 U3558 ( .x(n1645), .a(n1560), .b(n883) );
    nand2i_6 U3559 ( .x(n3428), .a(n4140), .b(n1147) );
    inv_2 U356 ( .x(n1115), .a(n1463) );
    nand2i_6 U3560 ( .x(n3429), .a(n1043), .b(n3790) );
    nand2i_6 U3561 ( .x(n3804), .a(n1771), .b(n530) );
    nand2i_6 U3562 ( .x(n3744), .a(n751), .b(n3743) );
    oai21_6 U3563 ( .x(n3778), .a(n1587), .b(n1642), .c(n3777) );
    nand2i_6 U3564 ( .x(n2410), .a(n2411), .b(n1217) );
    inv_10 U3565 ( .x(n1555), .a(n1554) );
    inv_6 U3566 ( .x(n3731), .a(n3730) );
    nand2i_6 U3567 ( .x(n2397), .a(n1476), .b(n2139) );
    nand2i_6 U3568 ( .x(n3508), .a(n1607), .b(n3658) );
    oai22_6 U3569 ( .x(n2148), .a(n784), .b(n1120), .c(
        ___cell__39620_net144406), .d(n1122) );
    nand2i_2 U357 ( .x(n2144), .a(n1574), .b(n2089) );
    inv_16 U3570 ( .x(n1177), .a(n1559) );
    inv_16 U3571 ( .x(n1683), .a(n4008) );
    nand2i_6 U3572 ( .x(n2322), .a(n1472), .b(n2139) );
    nand2i_6 U3573 ( .x(n2292), .a(n1470), .b(n2139) );
    nand2i_6 U3574 ( .x(n3441), .a(n815), .b(n3683) );
    inv_16 U3575 ( .x(n1656), .a(n912) );
    nand2i_6 U3576 ( .x(n3672), .a(n1562), .b(n3619) );
    nor2i_8 U3577 ( .x(n1044), .a(n1045), .b(n4005) );
    nand2i_5 U3578 ( .x(n3643), .a(n1608), .b(n3537) );
    nand2i_5 U3579 ( .x(n3642), .a(n1072), .b(n1361) );
    nand3_2 U358 ( .x(n2099), .a(n2081), .b(n3685), .c(n2084) );
    nand2i_6 U3580 ( .x(n3641), .a(n1607), .b(n3638) );
    nand2i_6 U3581 ( .x(n3674), .a(n1607), .b(n3628) );
    oai22_6 U3582 ( .x(n2136), .a(n1642), .b(n1656), .c(n915), .d(n1657) );
    nor2i_5 U3583 ( .x(n1065), .a(n1066), .b(n1067) );
    nand2i_5 U3584 ( .x(n3680), .a(n4010), .b(n2181) );
    nand2i_6 U3585 ( .x(n2048), .a(n1459), .b(n2139) );
    inv_16 U3586 ( .x(n1529), .a(n904) );
    nand2i_6 U3587 ( .x(n3580), .a(n1623), .b(n4142) );
    inv_7 U3588 ( .x(n1553), .a(n1157) );
    oai21_6 U3589 ( .x(n1836), .a(n1642), .b(n1646), .c(n1837) );
    nand2i_2 U359 ( .x(n2150), .a(n670), .b(n2099) );
    inv_16 U3590 ( .x(n3591), .a(n1642) );
    nand2i_5 U3591 ( .x(n1432), .a(n3233), .b(n3234) );
    nand3i_5 U3592 ( .x(n3182), .a(n1416), .b(n3183), .c(n3184) );
    nor2i_5 U3593 ( .x(n1176), .a(n1177), .b(n1178) );
    aoi21_5 U3594 ( .x(n2338), .a(n1971), .b(n2184), .c(n1174) );
    nand2i_6 U3595 ( .x(n3416), .a(n1655), .b(n3592) );
    nand2_8 U3596 ( .x(n3349), .a(n1691), .b(n628) );
    nand2i_6 U3597 ( .x(n3350), .a(n1656), .b(n883) );
    nand2_8 U3598 ( .x(n1690), .a(n1691), .b(n504) );
    buf_16 U3599 ( .x(n4011), .a(n1631) );
    inv_8 U36 ( .x(net156363), .a(___cell__39620_net143997) );
    nor2_1 U360 ( .x(n1117), .a(n4002), .b(___cell__39620_net143735) );
    aoi22_4 U3600 ( .x(n2334), .a(n1289), .b(n2080), .c(n2335), .d(n636) );
    nand2_8 U3601 ( .x(n3342), .a(n1686), .b(n628) );
    nand2i_6 U3603 ( .x(n3412), .a(n1644), .b(n3592) );
    nand2i_8 U3604 ( .x(n3638), .a(n3389), .b(n3627) );
    nand2i_8 U3605 ( .x(n3655), .a(n3486), .b(n3627) );
    nand2_3 U3606 ( .x(n3980), .a(n504), .b(n2187) );
    nand2_3 U3607 ( .x(n3979), .a(n1714), .b(n2000) );
    oai22_6 U3608 ( .x(n3356), .a(n915), .b(n1656), .c(n3357), .d(n815) );
    oai22_6 U3609 ( .x(n3530), .a(n891), .b(n3294), .c(n1651), .d(n1656) );
    inv_2 U361 ( .x(n3505), .a(n2045) );
    nand2_8 U3610 ( .x(n3817), .a(n3311), .b(n855) );
    nand2_8 U3611 ( .x(n3617), .a(n3556), .b(n855) );
    inv_16 U3612 ( .x(n1586), .a(n901) );
    nand2i_6 U3613 ( .x(n2677), .a(n751), .b(n3802) );
    oai22_6 U3614 ( .x(n3036), .a(n1573), .b(n1629), .c(n1569), .d(n825) );
    nand2_8 U3615 ( .x(n2991), .a(n3567), .b(n3568) );
    nand2_8 U3616 ( .x(n3069), .a(n3361), .b(n3362) );
    nand2_8 U3617 ( .x(n2927), .a(n3297), .b(n3298) );
    nor2i_5 U3618 ( .x(n1329), .a(n1330), .b(n1331) );
    inv_10 U3619 ( .x(n1605), .a(n3576) );
    mux2i_1 U362 ( .x(n2157), .d0(n3546), .sl(n816), .d1(n3442) );
    nand2_6 U3620 ( .x(n3033), .a(n3363), .b(n3364) );
    oai22_6 U3621 ( .x(n2852), .a(n1629), .b(n1649), .c(n1579), .d(n881) );
    nand2_8 U3622 ( .x(n2854), .a(n3372), .b(n3373) );
    inv_16 U3623 ( .x(n1571), .a(n644) );
    nand2_8 U3624 ( .x(n2783), .a(n3300), .b(n3301) );
    oai22_6 U3625 ( .x(n2851), .a(n1571), .b(n881), .c(n1629), .d(n1644) );
    inv_7 U3626 ( .x(n1287), .a(n2981) );
    nand2i_5 U3627 ( .x(n2629), .a(n1156), .b(n1558) );
    aoi22_6 U3628 ( .x(n2926), .a(n1066), .b(n2927), .c(
        ___cell__39620_net144517), .d(n2854) );
    nand2i_5 U3629 ( .x(n3901), .a(n1635), .b(n2995) );
    nor2_1 U363 ( .x(n1118), .a(n1087), .b(n4042) );
    oai22_6 U3630 ( .x(n3020), .a(n1629), .b(n1656), .c(n1563), .d(n881) );
    nand2i_6 U3631 ( .x(n2633), .a(n1605), .b(n3725) );
    nand2i_6 U3632 ( .x(n3888), .a(n1851), .b(n530) );
    nand2_8 U3633 ( .x(n2784), .a(n3376), .b(n3377) );
    nand2_6 U3634 ( .x(n2890), .a(n3295), .b(n3296) );
    nand2i_6 U3635 ( .x(n3569), .a(n4140), .b(n1289) );
    oai22_6 U3636 ( .x(n3535), .a(n891), .b(n3306), .c(n1573), .d(n1651) );
    buf_16 U3639 ( .x(n4013), .a(n1622) );
    inv_2 U364 ( .x(n1113), .a(N1869) );
    nor2i_5 U3640 ( .x(n1282), .a(n1147), .b(n1283) );
    nand2i_6 U3641 ( .x(n3863), .a(n1644), .b(n811) );
    nand2i_6 U3642 ( .x(n3367), .a(n1578), .b(n3592) );
    nand2i_6 U3643 ( .x(n3400), .a(n1529), .b(n3584) );
    nor2i_5 U3644 ( .x(n1248), .a(n1249), .b(n1250) );
    oai21_6 U3645 ( .x(n2649), .a(n4125), .b(n1148), .c(n3453) );
    nand2_8 U3646 ( .x(n3742), .a(n3351), .b(n855) );
    nand2_8 U3647 ( .x(n3772), .a(n3332), .b(n855) );
    nand2i_6 U3648 ( .x(n2262), .a(n3565), .b(n3566) );
    nand2i_6 U3649 ( .x(n2277), .a(n501), .b(n3501) );
    nor2_1 U365 ( .x(n1112), .a(n947), .b(n1113) );
    nand2i_6 U3650 ( .x(n3791), .a(n1760), .b(n1063) );
    nand2i_6 U3651 ( .x(n3786), .a(n4140), .b(n2458) );
    oai211_5 U3652 ( .x(n2305), .a(n506), .b(n1546), .c(n3401), .d(n3402) );
    nand2i_6 U3653 ( .x(n3718), .a(n1580), .b(n3591) );
    nand2_8 U3654 ( .x(n3407), .a(n1691), .b(n908) );
    nand2i_6 U3655 ( .x(n3408), .a(n1573), .b(n883) );
    nand2i_6 U3656 ( .x(n3721), .a(n1578), .b(n811) );
    aoi21_4 U3657 ( .x(n2276), .a(n1289), .b(n2277), .c(n1146) );
    nand2i_6 U3658 ( .x(n3722), .a(n1580), .b(n3594) );
    nor2i_1 U366 ( .x(n1111), .a(N1737), .b(___cell__39620_net143710) );
    nand2_8 U3660 ( .x(n3398), .a(n1686), .b(n908) );
    nand2i_6 U3661 ( .x(n3399), .a(n1573), .b(n928) );
    aoi21_6 U3662 ( .x(n2065), .a(n2066), .b(n634), .c(n2067) );
    nand2i_6 U3663 ( .x(n3733), .a(n1219), .b(n811) );
    aoi21_4 U3664 ( .x(n2261), .a(n1289), .b(n2262), .c(n1151) );
    nor2i_8 U3665 ( .x(n1109), .a(n686), .b(n1091) );
    inv_16 U3666 ( .x(n1644), .a(n922) );
    nand2i_6 U3667 ( .x(n2080), .a(n1605), .b(n3577) );
    nor2i_8 U3668 ( .x(n1090), .a(n634), .b(n1091) );
    nand2i_8 U3669 ( .x(n1687), .a(n1546), .b(n504) );
    nand2i_2 U367 ( .x(n3103), .a(n1512), .b(n2139) );
    nand2i_6 U3670 ( .x(n3183), .a(n1682), .b(n1045) );
    nand2i_6 U3671 ( .x(n3184), .a(n1657), .b(n3202) );
    nor2i_8 U3672 ( .x(n1174), .a(n634), .b(n1175) );
    inv_16 U3673 ( .x(n3592), .a(n1645) );
    inv_14 U3674 ( .x(n1685), .a(n1624) );
    inv_8 U3675 ( .x(n2070), .a(n1418) );
    inv_16 U3676 ( .x(n1982), .a(n1419) );
    inv_10 U3677 ( .x(n2227), .a(n2128) );
    nand2i_6 U3679 ( .x(n3503), .a(n1577), .b(n927) );
    nand2_2 U368 ( .x(n690), .a(___cell__39620_net147732), .b(
        ___cell__39620_net144201) );
    inv_6 U3680 ( .x(n3517), .a(n3560) );
    nand2i_5 U3683 ( .x(n3567), .a(n1219), .b(n874) );
    nand2i_5 U3685 ( .x(n3361), .a(n1587), .b(n874) );
    nand2i_5 U3686 ( .x(n3297), .a(n1649), .b(n874) );
    nand2i_5 U3687 ( .x(n3363), .a(n1580), .b(n874) );
    nand2i_6 U3689 ( .x(n3372), .a(n1571), .b(n928) );
    oai21_1 U369 ( .x(n3102), .a(n1511), .b(n690), .c(n3103) );
    nand2i_6 U3690 ( .x(n3548), .a(n1572), .b(n927) );
    nand2i_5 U3691 ( .x(n3549), .a(n1646), .b(n874) );
    nand2i_6 U3692 ( .x(n3292), .a(n1529), .b(n928) );
    nand2i_6 U3693 ( .x(n3304), .a(n1570), .b(n928) );
    nand2_8 U3694 ( .x(n3725), .a(___cell__39620_net144328), .b(
        ___cell__39620_net144331) );
    nand2i_6 U3695 ( .x(n3376), .a(n1585), .b(n928) );
    inv_6 U3698 ( .x(n1148), .a(n3394) );
    nand2i_5 U3699 ( .x(n3453), .a(n1579), .b(n874) );
    inv_12 U37 ( .x(n609), .a(n1585) );
    nand2i_0 U370 ( .x(n1388), .a(n1579), .b(n530) );
    nand2_8 U3700 ( .x(n1715), .a(n1691), .b(n1714) );
    nand2i_6 U3701 ( .x(n1713), .a(n1546), .b(n1714) );
    nand2i_6 U3702 ( .x(n3402), .a(n1587), .b(n883) );
    nor2i_5 U3704 ( .x(n1146), .a(n1147), .b(n1148) );
    aoi21_6 U3705 ( .x(n2110), .a(n2066), .b(n686), .c(n2067) );
    inv_10 U3706 ( .x(n2066), .a(n1672) );
    nand2i_6 U3707 ( .x(n1974), .a(n855), .b(n1553) );
    inv_6 U3708 ( .x(n2214), .a(n3340) );
    nand2_8 U3709 ( .x(n1556), .a(n1555), .b(n855) );
    aoi21_1 U371 ( .x(n1387), .a(n1143), .b(n1388), .c(n653) );
    nand2i_6 U3710 ( .x(n3657), .a(n924), .b(n910) );
    nand2i_5 U3711 ( .x(n3574), .a(n924), .b(n901) );
    inv_16 U3712 ( .x(n3575), .a(n4013) );
    nand2i_6 U3713 ( .x(n2115), .a(n1644), .b(n928) );
    nor2_1 U372 ( .x(n1389), .a(n4002), .b(n588) );
    inv_2 U373 ( .x(n1382), .a(N1809) );
    nor2_1 U374 ( .x(n1381), .a(n1077), .b(n1382) );
    inv_12 U375 ( .x(n1579), .a(reg_out_A[12]) );
    ao211_5 U3750 ( .x(n3084), .a(n3110), .b(n1267), .c(n4119), .d(n4118) );
    inv_0 U3751 ( .x(n4118), .a(n3089) );
    inv_2 U3752 ( .x(n4119), .a(n3088) );
    nand2i_1 U3753 ( .x(n3088), .a(n4022), .b(n3057) );
    ao211_5 U3754 ( .x(n2806), .a(n3464), .b(n4122), .c(n4121), .d(n4120) );
    inv_2 U3755 ( .x(n4120), .a(n2216) );
    inv_4 U3756 ( .x(n4121), .a(n3331) );
    inv_0 U3757 ( .x(n4122), .a(___cell__39620_net144317) );
    nand2i_5 U3758 ( .x(n2216), .a(n1649), .b(n4130) );
    nand2_1 U3759 ( .x(n3331), .a(n1686), .b(n749) );
    nor2i_1 U376 ( .x(n1376), .a(n1377), .b(___cell__39620_net143658) );
    ao21_6 U3760 ( .x(n2603), .a(n4124), .b(n3388), .c(n4123) );
    inv_2 U3761 ( .x(n4123), .a(n3461) );
    inv_3 U3762 ( .x(n4124), .a(n4125) );
    inv_14 U3763 ( .x(n4125), .a(___cell__39620_net144317) );
    inv_4 U3764 ( .x(n1152), .a(n3388) );
    nand2i_6 U3765 ( .x(n3388), .a(n3389), .b(n3390) );
    nand3_2 U3766 ( .x(n2868), .a(n730), .b(n2873), .c(n2871) );
    inv_3 U3767 ( .x(___cell__39620_net144317), .a(Imm[3]) );
    inv_12 U3768 ( .x(net149167), .a(n799) );
    nand2i_2 U3769 ( .x(n2897), .a(n1626), .b(n3873) );
    nor2i_1 U377 ( .x(n1378), .a(N1710), .b(___cell__39620_net143660) );
    nand2i_1 U3770 ( .x(n2866), .a(n1641), .b(n3873) );
    oai211_3 U3771 ( .x(n3873), .a(n3529), .b(___cell__39620_net144345), .c(
        n3871), .d(n3872) );
    inv_5 U3772 ( .x(n3130), .a(n2050) );
    aoi21_1 U3773 ( .x(n2049), .a(n1221), .b(n2050), .c(n2046) );
    nand2i_0 U3774 ( .x(n2015), .a(n1588), .b(n2050) );
    oai221_4 U3775 ( .x(n2050), .a(n3439), .b(n1559), .c(n747), .d(n1562), .e(
        n1975) );
    ao222_4 U3776 ( .x(n2908), .a(n2874), .b(n755), .c(n2875), .d(n756), .e(
        ALU_result[18]), .f(n3057) );
    aoi211_2 U3777 ( .x(n730), .a(n2798), .b(n1085), .c(n732), .d(n731) );
    inv_6 U3778 ( .x(n731), .a(n2876) );
    aoi211_1 U3779 ( .x(n998), .a(n977), .b(N348), .c(n2051), .d(n2055) );
    inv_5 U378 ( .x(n3546), .a(n3545) );
    nand2i_3 U3780 ( .x(n3300), .a(n1656), .b(n874) );
    oai21_2 U3781 ( .x(n2898), .a(n1566), .b(n4126), .c(n3890) );
    inv_5 U3782 ( .x(n4126), .a(n2899) );
    nand4i_4 U3783 ( .x(n2899), .a(n1299), .b(n3881), .c(n3880), .d(n3879) );
    inv_16 U3784 ( .x(n649), .a(n1566) );
    nand2i_0 U3785 ( .x(n3890), .a(n1500), .b(n2139) );
    nand2i_5 U3786 ( .x(n1566), .a(___cell__39620_net144175), .b(n1567) );
    nand2_3 U3787 ( .x(n695), .a(n713), .b(n4130) );
    nand2i_2 U3788 ( .x(n2163), .a(n1656), .b(n4130) );
    nand2i_2 U3789 ( .x(n3568), .a(n862), .b(n4130) );
    nor2i_3 U379 ( .x(n1106), .a(___cell__39620_net143722), .b(n746) );
    nand2i_2 U3790 ( .x(n3562), .a(n1648), .b(n4130) );
    nand2i_2 U3791 ( .x(n3364), .a(n748), .b(n4130) );
    nand2i_2 U3792 ( .x(n3686), .a(n1655), .b(n4130) );
    nand2i_2 U3793 ( .x(n3295), .a(n1586), .b(n4130) );
    nand2i_1 U3794 ( .x(n3393), .a(n1587), .b(n4130) );
    oai22_2 U3795 ( .x(n2189), .a(n895), .b(n4001), .c(n3525), .d(n784) );
    aoi211_2 U3796 ( .x(n2879), .a(N1650), .b(n809), .c(n1303), .d(n2878) );
    nor2i_5 U3797 ( .x(n1303), .a(N1716), .b(___cell__39620_net143660) );
    aoi22_2 U3798 ( .x(n2712), .a(n2713), .b(___cell__39620_net143722), .c(
        ___cell__39620_net143864), .d(n2714) );
    inv_3 U3799 ( .x(n1205), .a(n2457) );
    nand4_1 U38 ( .x(n3221), .a(n1506), .b(n1504), .c(n1509), .d(n1507) );
    aoi21_1 U380 ( .x(n2084), .a(n1249), .b(n2000), .c(n2082) );
    nand2_1 U3800 ( .x(n4128), .a(n3502), .b(n3503) );
    nand2_2 U3801 ( .x(n4127), .a(n3502), .b(n3503) );
    nand2i_3 U3802 ( .x(n3502), .a(n1578), .b(n874) );
    nand2_1 U3803 ( .x(n3097), .a(n3502), .b(n3503) );
    oai221_1 U3804 ( .x(n4129), .a(n3553), .b(___cell__39620_net144374), .c(
        n3299), .d(n1623), .e(n2853) );
    aoi22_2 U3805 ( .x(n2853), .a(n1066), .b(n2854), .c(n1683), .d(n2563) );
    buf_14 U3806 ( .x(n4130), .a(n531) );
    buf_8 U3807 ( .x(n927), .a(n531) );
    buf_14 U3808 ( .x(n928), .a(n531) );
    nand2_5 U3809 ( .x(n3034), .a(n3359), .b(n3360) );
    nand2_1 U381 ( .x(n3685), .a(n1256), .b(n2187) );
    nand2i_4 U3810 ( .x(n3360), .a(n1569), .b(n928) );
    nand2i_4 U3811 ( .x(n3359), .a(n1573), .b(n874) );
    oai31_2 U3812 ( .x(n1010), .a(n2425), .b(n2413), .c(n2418), .d(
        ___cell__39620_net143326) );
    ao21_6 U3813 ( .x(n3765), .a(n4131), .b(n3723), .c(n4132) );
    inv_0 U3814 ( .x(n4131), .a(net149122) );
    ao22_3 U3815 ( .x(n4132), .a(___cell__39620_net144517), .b(n2279), .c(
        n1391), .d(n2375) );
    buf_16 U3816 ( .x(net149122), .a(net149107) );
    oai211_3 U3817 ( .x(n2302), .a(n550), .b(___cell__39620_net144317), .c(
        n3392), .d(n3393) );
    inv_4 U3818 ( .x(n550), .a(n3496) );
    oai221_2 U3819 ( .x(n3116), .a(n511), .b(n1635), .c(n3335), .d(n4009), .e(
        n3098) );
    aoi21_1 U382 ( .x(n2081), .a(n1714), .b(n1999), .c(n1092) );
    oa22_5 U3820 ( .x(n511), .a(n1570), .b(n1629), .c(n512), .d(n536) );
    inv_7 U3821 ( .x(n912), .a(n911) );
    oai22_1 U3822 ( .x(n4133), .a(n1572), .b(n836), .c(n3397), .d(n4125) );
    oai22_1 U3823 ( .x(n4134), .a(n1572), .b(n836), .c(n3397), .d(n4125) );
    oai22_1 U3824 ( .x(n2563), .a(n1572), .b(n836), .c(n3397), .d(n4125) );
    inv_10 U3825 ( .x(n3397), .a(n3541) );
    nand4_2 U3826 ( .x(n4078), .a(n993), .b(n992), .c(n991), .d(n990) );
    nand4_1 U3827 ( .x(n4077), .a(n1010), .b(n1008), .c(n1009), .d(n1007) );
    aoi22_1 U3828 ( .x(n2739), .a(n1683), .b(n2649), .c(
        ___cell__39620_net144517), .d(n4134) );
    nand2i_1 U3829 ( .x(n3829), .a(n1625), .b(n4133) );
    nand2i_2 U383 ( .x(n3679), .a(n1623), .b(n3457) );
    inv_6 U3830 ( .x(n933), .a(n932) );
    inv_10 U3831 ( .x(n934), .a(n932) );
    inv_7 U3832 ( .x(n932), .a(reg_out_A[14]) );
    nand4_2 U3833 ( .x(n2055), .a(n2058), .b(n2057), .c(n579), .d(n2053) );
    nand4_2 U3834 ( .x(n2425), .a(n2422), .b(n2426), .c(n2427), .d(n2424) );
    nand4_3 U3835 ( .x(_ALU_result_reg_31_net106451), .a(
        ___cell__39620_net143598), .b(___cell__39620_net143595), .c(
        ___cell__39620_net143597), .d(___cell__39620_net143596) );
    and4i_5 U3836 ( .x(___cell__39620_net143598), .a(n2295), .b(n2299), .c(
        n2298), .d(n2297) );
    nand2i_4 U3837 ( .x(n2426), .a(n1759), .b(n1987) );
    inv_3 U3838 ( .x(n1751), .a(N1859) );
    and4i_3 U3839 ( .x(n990), .a(n2392), .b(n2389), .c(n2404), .d(n2401) );
    nand4_1 U384 ( .x(n3681), .a(n3679), .b(n3678), .c(n3680), .d(n2078) );
    oai211_2 U3840 ( .x(n2392), .a(n2393), .b(n4001), .c(n2394), .d(n2395) );
    aoi211_2 U3841 ( .x(n2073), .a(N1705), .b(___cell__39620_net145190), .c(
        n1097), .d(n1096) );
    aoi22_3 U3842 ( .x(n2385), .a(N1826), .b(n1987), .c(n1095), .d(n2386) );
    inv_14 U3843 ( .x(n637), .a(n738) );
    inv_7 U3844 ( .x(n2429), .a(n2270) );
    nand2_5 U3845 ( .x(n2270), .a(n3563), .b(n3564) );
    inv_4 U3846 ( .x(n931), .a(n929) );
    inv_10 U3847 ( .x(n930), .a(n929) );
    inv_6 U3848 ( .x(n929), .a(reg_out_A[13]) );
    nor2i_2 U3849 ( .x(n1240), .a(N1654), .b(___cell__39620_net143872) );
    nor2_1 U385 ( .x(n1105), .a(___cell__39620_net143693), .b(
        ___cell__39620_net143720) );
    aoai211_4 U3850 ( .x(n4049), .a(___cell__39620_net143287), .b(n1455), .c(
        n1439), .d(n1456) );
    nand2_4 U3851 ( .x(n613), .a(n615), .b(n614) );
    nand2i_2 U3852 ( .x(n3712), .a(n727), .b(n2809) );
    oai211_3 U3853 ( .x(n2809), .a(n3334), .b(n1546), .c(n3339), .d(n3340) );
    nor2_2 U3854 ( .x(n1953), .a(reg_out_B[8]), .b(reg_out_B[9]) );
    nand2i_4 U3855 ( .x(n736), .a(reg_out_B[29]), .b(n1731) );
    inv_0 U3856 ( .x(n4135), .a(net149617) );
    inv_2 U3857 ( .x(n4136), .a(n4135) );
    inv_6 U3858 ( .x(net149617), .a(net149616) );
    nand3_4 U3859 ( .x(n679), .a(n678), .b(n1663), .c(n701) );
    nand2i_2 U386 ( .x(n2087), .a(n1461), .b(n2139) );
    inv_6 U3860 ( .x(n701), .a(___cell__39620_net144175) );
    buf_2 U3861 ( .x(n4015), .a(reg_out_A[1]) );
    and2_1 U3862 ( .x(n4137), .a(n4138), .b(IR_opcode_field[4]) );
    inv_2 U3863 ( .x(n1609), .a(n4137) );
    inv_0 U3864 ( .x(n4138), .a(IR_opcode_field[5]) );
    buf_8 U3865 ( .x(net149107), .a(Imm[1]) );
    inv_10 U3866 ( .x(n896), .a(n1554) );
    nand2i_8 U3867 ( .x(n1554), .a(reg_out_B[5]), .b(n1552) );
    and2_5 U3868 ( .x(n1241), .a(N1720), .b(___cell__39620_net145190) );
    nand2i_4 U3869 ( .x(___cell__39620_net143660), .a(IR_opcode_field[2]), .b(
        ___cell__39620_net144309) );
    inv_2 U387 ( .x(n3688), .a(n1462) );
    inv_16 U3870 ( .x(___cell__39620_net145190), .a(___cell__39620_net143660)
         );
    nand2i_2 U3871 ( .x(n2152), .a(n1641), .b(n3689) );
    nand2i_2 U3872 ( .x(n2257), .a(n1641), .b(n3711) );
    nand2i_4 U3873 ( .x(n2895), .a(n1641), .b(n3887) );
    nand2i_2 U3874 ( .x(n2407), .a(n1641), .b(n2455) );
    nand2i_2 U3875 ( .x(n2976), .a(n1641), .b(n3009) );
    nand2i_1 U3876 ( .x(n2029), .a(n1641), .b(n3583) );
    nand2i_2 U3877 ( .x(n2102), .a(n1641), .b(n3681) );
    oai22_2 U3878 ( .x(n2489), .a(n621), .b(n1122), .c(n1641), .d(n1120) );
    nand2i_2 U3879 ( .x(n3143), .a(n1641), .b(n3168) );
    nand2_2 U388 ( .x(n2086), .a(n2193), .b(n3688) );
    inv_3 U3880 ( .x(n905), .a(Imm[13]) );
    inv_2 U3881 ( .x(n555), .a(Imm[13]) );
    aoi22_3 U3882 ( .x(n2312), .a(N1827), .b(n1987), .c(N1860), .d(n4000) );
    nand2_2 U3883 ( .x(n1632), .a(n816), .b(reg_out_B[2]) );
    or2_6 U3884 ( .x(n1565), .a(reg_out_B[2]), .b(reg_out_B[3]) );
    nand2_1 U3885 ( .x(n1634), .a(n879), .b(reg_out_B[2]) );
    inv_7 U3886 ( .x(n828), .a(reg_out_B[2]) );
    buf_10 U3887 ( .x(n608), .a(reg_out_A[15]) );
    buf_4 U3888 ( .x(n4139), .a(reg_out_B[21]) );
    buf_8 U3889 ( .x(n918), .a(n931) );
    oai211_1 U389 ( .x(n2085), .a(n1104), .b(n1671), .c(n2086), .d(n2087) );
    buf_6 U3890 ( .x(n4014), .a(reg_out_A[15]) );
    buf_5 U3891 ( .x(n4016), .a(reg_out_A[15]) );
    buf_4 U3892 ( .x(n602), .a(reg_out_A[15]) );
    nand2_8 U3893 ( .x(n4140), .a(___cell__39620_net144330), .b(reg_out_A[31])
         );
    inv_10 U3894 ( .x(n817), .a(Imm[10]) );
    or3i_5 U3895 ( .x(n1957), .a(n605), .b(reg_out_B[20]), .c(reg_out_B[18])
         );
    nand4i_1 U3896 ( .x(n4141), .a(n1360), .b(n3968), .c(n3967), .d(n3966) );
    oai211_2 U3897 ( .x(n4069), .a(n1020), .b(___cell__39620_net143287), .c(
        n1021), .d(n1022) );
    ao21_4 U3898 ( .x(n4142), .a(net150830), .b(n2080), .c(n837) );
    inv_5 U3899 ( .x(n837), .a(n3456) );
    exnor2_1 U39 ( .x(n3231), .a(net152465), .b(n942) );
    nor2_1 U390 ( .x(n1107), .a(n1087), .b(n4043) );
    ao211_2 U3900 ( .x(n4067), .a(___cell__39620_net143326), .b(n974), .c(n975
        ), .d(n976) );
    nand4i_2 U3901 ( .x(n974), .a(n1309), .b(n2882), .c(n2881), .d(n2883) );
    inv_16 U3902 ( .x(N69), .a(reg_out_A[31]) );
    nand2_8 U3903 ( .x(n1159), .a(n896), .b(reg_out_A[31]) );
    inv_0 U3904 ( .x(n4143), .a(reg_out_B[31]) );
    inv_2 U3905 ( .x(n4144), .a(n4143) );
    nor2_2 U3906 ( .x(n1955), .a(reg_out_B[13]), .b(reg_out_B[14]) );
    inv_6 U3907 ( .x(n4145), .a(reg_out_B[7]) );
    inv_10 U3908 ( .x(n4146), .a(n4145) );
    inv_5 U3909 ( .x(n759), .a(reg_out_B[5]) );
    oai22_2 U391 ( .x(n2135), .a(n890), .b(n1656), .c(n1651), .d(n1657) );
    buf_1 U3910 ( .x(n4147), .a(reg_out_B[9]) );
    buf_16 U3911 ( .x(mem_to_reg_EX), .a(n4224) );
    nor2_1 U3912 ( .x(n1952), .a(reg_out_B[6]), .b(n4146) );
    nor2_2 U3913 ( .x(n1958), .a(reg_out_B[23]), .b(reg_out_B[24]) );
    nor2_3 U3914 ( .x(n1959), .a(reg_out_B[25]), .b(reg_out_B[26]) );
    nor2_1 U3915 ( .x(n1954), .a(reg_out_B[10]), .b(reg_out_B[11]) );
    nor2i_0 U3916 ( .x(n4156), .a(reg_out_B[24]), .b(n4116) );
    and2_1 U3917 ( .x(n4158), .a(reg_out_B[15]), .b(n4117) );
    nor2i_0 U3918 ( .x(n4160), .a(n816), .b(___cell__6067_net21981) );
    nor2i_0 U3919 ( .x(n4162), .a(n566), .b(n4116) );
    inv_5 U392 ( .x(n852), .a(n851) );
    nor2i_0 U3920 ( .x(n4164), .a(reg_out_B[30]), .b(n4116) );
    nor2i_0 U3921 ( .x(n4166), .a(reg_out_B[28]), .b(n4116) );
    nor2i_0 U3922 ( .x(n4168), .a(reg_out_B[27]), .b(n4116) );
    nor2i_0 U3923 ( .x(n4170), .a(reg_out_B[25]), .b(n4116) );
    nor2i_0 U3924 ( .x(n4172), .a(reg_out_B[23]), .b(n4116) );
    nor2i_0 U3925 ( .x(n4174), .a(reg_out_B[19]), .b(n4116) );
    nor2i_0 U3926 ( .x(n4176), .a(reg_out_B[16]), .b(n4116) );
    and2_1 U3927 ( .x(n4178), .a(reg_out_B[14]), .b(n4117) );
    and2_1 U3928 ( .x(n4180), .a(reg_out_B[12]), .b(n4117) );
    and2_1 U3929 ( .x(n4182), .a(reg_out_B[10]), .b(n4117) );
    inv_2 U393 ( .x(n3793), .a(n1479) );
    and2_1 U3930 ( .x(n4184), .a(reg_out_B[8]), .b(n4117) );
    nor2i_0 U3931 ( .x(n4186), .a(n4146), .b(___cell__6067_net21981) );
    nor2i_0 U3932 ( .x(n4188), .a(reg_out_B[6]), .b(___cell__6067_net21981) );
    nor2i_0 U3933 ( .x(n4190), .a(reg_out_B[5]), .b(___cell__6067_net21981) );
    nor2i_0 U3934 ( .x(n4192), .a(reg_out_B[4]), .b(___cell__6067_net21981) );
    nor2i_0 U3935 ( .x(n4194), .a(n536), .b(___cell__6067_net21981) );
    nor2i_0 U3936 ( .x(n4196), .a(n815), .b(___cell__6067_net21981) );
    and2_1 U3937 ( .x(n4198), .a(reg_write), .b(N3304) );
    and2_1 U3938 ( .x(n4200), .a(mem_to_reg), .b(N3304) );
    and2_1 U3939 ( .x(n4202), .a(mem_read), .b(N3304) );
    nand2_2 U394 ( .x(n2483), .a(n2193), .b(n3793) );
    and2_1 U3940 ( .x(n4203), .a(mem_write), .b(N3304) );
    nor2i_0 U3941 ( .x(n4204), .a(reg_out_B[22]), .b(n4116) );
    nor2i_0 U3942 ( .x(n4206), .a(reg_out_B[26]), .b(n4116) );
    and2_1 U3943 ( .x(n4208), .a(n4147), .b(n4117) );
    nor2i_0 U3944 ( .x(n4210), .a(reg_out_B[18]), .b(n4116) );
    nor2i_0 U3945 ( .x(n4212), .a(reg_out_B[0]), .b(___cell__6067_net21981) );
    and2_1 U3946 ( .x(n4214), .a(reg_out_B[11]), .b(n4117) );
    and2_1 U3947 ( .x(n4216), .a(reg_out_B[13]), .b(n4117) );
    nor2i_0 U3948 ( .x(n4218), .a(reg_out_B[20]), .b(n4116) );
    nor2i_0 U3949 ( .x(n4220), .a(reg_out_B[29]), .b(n4116) );
    nand2i_2 U395 ( .x(n2482), .a(n1480), .b(n2139) );
    nor2i_0 U3950 ( .x(n4222), .a(reg_out_B[17]), .b(n4116) );
    oa22_2 U396 ( .x(n505), .a(n1637), .b(n1093), .c(n1626), .d(n1089) );
    oai211_1 U397 ( .x(n2481), .a(n505), .b(n1580), .c(n2482), .d(n2483) );
    nand2i_3 U398 ( .x(n2487), .a(n2459), .b(n866) );
    inv_2 U399 ( .x(n3792), .a(n3791) );
    nand4_1 U40 ( .x(n3230), .a(n3231), .b(n1458), .c(n1462), .d(n1460) );
    nand2i_2 U400 ( .x(n2461), .a(n816), .b(n502) );
    nand2i_2 U401 ( .x(n2485), .a(n2461), .b(n3778) );
    nand2_2 U402 ( .x(n3743), .a(n3477), .b(___cell__39620_net144331) );
    inv_2 U403 ( .x(n1766), .a(N1758) );
    nand2i_2 U404 ( .x(n2468), .a(n1766), .b(___cell__39620_net145150) );
    nand2i_0 U405 ( .x(n2467), .a(___cell__39620_net144655), .b(n663) );
    nand2_2 U406 ( .x(n2462), .a(n681), .b(n537) );
    nand2i_2 U407 ( .x(n2464), .a(n2462), .b(___cell__39620_net145285) );
    inv_2 U408 ( .x(n1933), .a(N1797) );
    inv_2 U409 ( .x(n1936), .a(N1830) );
    inv_2 U41 ( .x(n2194), .a(n1465) );
    oai22_1 U410 ( .x(n3252), .a(n946), .b(n1936), .c(n1077), .d(n1933) );
    inv_2 U411 ( .x(n1930), .a(N1731) );
    inv_2 U412 ( .x(n1929), .a(N1698) );
    oai221_1 U413 ( .x(n3249), .a(___cell__39620_net143660), .b(n1929), .c(
        ___cell__39620_net143710), .d(n1930), .e(n3250) );
    ao211_3 U414 ( .x(n3251), .a(n1318), .b(n1423), .c(n3249), .d(n3252) );
    nand2i_2 U415 ( .x(n3255), .a(n1934), .b(n3624) );
    inv_2 U416 ( .x(n1934), .a(N1996) );
    inv_2 U417 ( .x(n1932), .a(N1930) );
    nand2i_2 U418 ( .x(n3254), .a(n1932), .b(n3662) );
    nand2i_2 U419 ( .x(n3253), .a(n1935), .b(___cell__39620_net145508) );
    inv_5 U42 ( .x(net152465), .a(n783) );
    inv_2 U420 ( .x(n1935), .a(N1963) );
    nor2i_1 U421 ( .x(n1438), .a(N1632), .b(___cell__39620_net143872) );
    nor2i_3 U422 ( .x(n1435), .a(n1436), .b(n1437) );
    aoi21_1 U423 ( .x(n3240), .a(net152465), .b(n3241), .c(n701) );
    aoai211_1 U424 ( .x(n3243), .a(n891), .b(n3539), .c(n3236), .d(n1095) );
    oai211_2 U425 ( .x(n3242), .a(n1430), .b(n1639), .c(n3243), .d(n3240) );
    oai21_1 U426 ( .x(n3237), .a(n1427), .b(n1089), .c(n1618) );
    inv_1 U427 ( .x(n545), .a(n889) );
    exnor2_1 U428 ( .x(n1945), .a(n3990), .b(___cell__39620_net144166) );
    ao222_2 U429 ( .x(n742), .a(n1256), .b(n2809), .c(n2273), .d(n893), .e(
        n1150), .f(n3279) );
    nand2i_0 U43 ( .x(n1527), .a(n1524), .b(n1528) );
    inv_5 U430 ( .x(n3860), .a(n1836) );
    inv_2 U431 ( .x(n1567), .a(n1544) );
    aoai211_1 U432 ( .x(n3286), .a(n3591), .b(n1567), .c(n3280), .d(n942) );
    nand2i_2 U433 ( .x(n1544), .a(n816), .b(n1545) );
    nand2i_2 U434 ( .x(n3285), .a(n1560), .b(n3715) );
    aoi21_1 U435 ( .x(n3277), .a(n1177), .b(n3278), .c(n3276) );
    aoai211_1 U436 ( .x(n3284), .a(n3277), .b(n3285), .c(n1544), .d(n3286) );
    exnor2_1 U437 ( .x(n1949), .a(n1950), .b(n1530) );
    mux2i_2 U438 ( .x(n3994), .d0(n1947), .sl(IR_function_field[0]), .d1(N1402
        ) );
    oaoi211_1 U439 ( .x(n1445), .a(n942), .b(n1446), .c(n1447), .d(n1448) );
    nand4_1 U44 ( .x(n3259), .a(n1505), .b(n1503), .c(n1510), .d(n1508) );
    nand2i_2 U440 ( .x(n1447), .a(n1531), .b(n1528) );
    inv_1 U441 ( .x(n1448), .a(reg_out_B[0]) );
    inv_2 U442 ( .x(n1537), .a(n1446) );
    nor2i_1 U443 ( .x(n1453), .a(N307), .b(n1454) );
    inv_2 U444 ( .x(n1593), .a(n1454) );
    nand2i_2 U445 ( .x(n3128), .a(n1513), .b(n2139) );
    exnor2_1 U446 ( .x(n1514), .a(n753), .b(n901) );
    inv_2 U447 ( .x(n3982), .a(n1514) );
    nand2_2 U448 ( .x(n3127), .a(n2193), .b(n3982) );
    aoi21_1 U449 ( .x(n1403), .a(n901), .b(n530), .c(n1064) );
    inv_0 U45 ( .x(n1916), .a(reg_out_B[10]) );
    inv_4 U450 ( .x(n1300), .a(n3022) );
    inv_3 U451 ( .x(n3417), .a(n3415) );
    nor2_0 U452 ( .x(n1404), .a(n1087), .b(n4021) );
    ao22_2 U453 ( .x(n716), .a(n1391), .b(n3034), .c(n1066), .d(n3097) );
    ao221_4 U454 ( .x(n3113), .a(n3451), .b(n715), .c(n714), .d(n713), .e(n716
        ) );
    nor2i_1 U455 ( .x(n1398), .a(N1841), .b(n946) );
    nor2i_0 U456 ( .x(n1394), .a(n753), .b(n1586) );
    nor2i_0 U457 ( .x(n1393), .a(n1394), .b(___cell__39620_net143658) );
    nor2i_3 U458 ( .x(n1395), .a(N1709), .b(___cell__39620_net143660) );
    inv_2 U459 ( .x(n1912), .a(N1874) );
    nand3_1 U46 ( .x(n3258), .a(n1513), .b(n1512), .c(n1515) );
    inv_5 U460 ( .x(n3459), .a(n2262) );
    nor2_1 U461 ( .x(n1269), .a(n679), .b(n4027) );
    exnor2_1 U462 ( .x(n1494), .a(n749), .b(n551) );
    inv_2 U463 ( .x(n2787), .a(n1494) );
    inv_2 U464 ( .x(n2786), .a(n1493) );
    aoi22_1 U465 ( .x(n2785), .a(n2139), .b(n2786), .c(n2193), .d(n2787) );
    inv_2 U466 ( .x(n1259), .a(n3020) );
    ao22_2 U467 ( .x(n2772), .a(n661), .b(n662), .c(net151904), .d(n663) );
    inv_2 U468 ( .x(n1826), .a(N1652) );
    nand2i_2 U469 ( .x(n2771), .a(n1826), .b(n809) );
    inv_0 U47 ( .x(n1771), .a(reg_out_B[26]) );
    nand2_2 U470 ( .x(n2764), .a(n551), .b(n749) );
    nand2i_2 U471 ( .x(n2770), .a(n2764), .b(___cell__39620_net147791) );
    inv_5 U472 ( .x(n3656), .a(n3655) );
    nand2i_2 U473 ( .x(n3043), .a(n1508), .b(n2139) );
    oai21_1 U474 ( .x(n3042), .a(n1507), .b(n690), .c(n3043) );
    nand2i_2 U475 ( .x(n1357), .a(n1571), .b(n530) );
    aoi21_1 U476 ( .x(n1356), .a(n1143), .b(n1357), .c(n1358) );
    nor2_1 U477 ( .x(n1359), .a(n4002), .b(___cell__39620_net143997) );
    nand2i_2 U478 ( .x(n3964), .a(n703), .b(n3013) );
    nor2_1 U48 ( .x(n3268), .a(n3269), .b(n3270) );
    inv_2 U480 ( .x(n1887), .a(N1877) );
    nand2i_2 U481 ( .x(n3027), .a(n1887), .b(n944) );
    nand2i_2 U482 ( .x(n3026), .a(n3023), .b(___cell__39620_net147791) );
    nand2i_2 U483 ( .x(n3025), .a(n1886), .b(n809) );
    inv_2 U484 ( .x(n1886), .a(N1646) );
    nor2i_1 U485 ( .x(n1350), .a(N1712), .b(___cell__39620_net143660) );
    nand2i_2 U486 ( .x(n3937), .a(n1043), .b(n3538) );
    nor2i_3 U487 ( .x(n1323), .a(n1147), .b(n1324) );
    nand2i_2 U488 ( .x(n3973), .a(n1510), .b(n2139) );
    inv_2 U489 ( .x(n1373), .a(n1509) );
    nor2_1 U49 ( .x(n3265), .a(n3266), .b(n3267) );
    nor2i_1 U490 ( .x(n1372), .a(n1373), .b(n690) );
    nand2i_2 U491 ( .x(n3970), .a(n727), .b(n2852) );
    nand2_2 U493 ( .x(n702), .a(n701), .b(n1661) );
    nand2i_2 U494 ( .x(n1370), .a(n1563), .b(n530) );
    aoi21_1 U495 ( .x(n1369), .a(n1143), .b(n1370), .c(n1371) );
    oa22_2 U499 ( .x(n849), .a(n3345), .b(n536), .c(n1561), .d(n1629) );
    inv_2 U50 ( .x(n2195), .a(n1466) );
    nand2i_2 U500 ( .x(n3965), .a(___cell__39620_net144062), .b(n3457) );
    aoi21_4 U501 ( .x(n630), .a(net150830), .b(n2080), .c(n837) );
    nand2i_0 U502 ( .x(n3089), .a(n1563), .b(n1700) );
    nor2_1 U504 ( .x(n1374), .a(___cell__39620_net143693), .b(n1375) );
    aoi22_1 U505 ( .x(n3032), .a(n1391), .b(n3033), .c(n1066), .d(n3034) );
    nand2i_2 U506 ( .x(n3957), .a(___cell__39620_net144374), .b(n4128) );
    inv_0 U507 ( .x(n1371), .a(reg_out_B[13]) );
    nor2i_1 U508 ( .x(n1364), .a(N1843), .b(n946) );
    inv_2 U509 ( .x(n1895), .a(N1876) );
    inv_8 U51 ( .x(n682), .a(___cell__39620_net144029) );
    nand2i_2 U510 ( .x(n3063), .a(n1895), .b(n3998) );
    nor2i_1 U511 ( .x(n1362), .a(N1711), .b(___cell__39620_net143660) );
    inv_14 U512 ( .x(n708), .a(___cell__39620_net144170) );
    inv_2 U513 ( .x(___cell__39620_net145285), .a(___cell__39620_net143658) );
    aoi21_1 U515 ( .x(n3061), .a(n3060), .b(___cell__39620_net145285), .c(
        n1362) );
    inv_2 U516 ( .x(n3157), .a(n1516) );
    exnor2_1 U517 ( .x(n1515), .a(n908), .b(reg_out_B[10]) );
    inv_2 U518 ( .x(n3156), .a(n1515) );
    aoi22_1 U519 ( .x(n3155), .a(n2139), .b(n3156), .c(n2193), .d(n3157) );
    nand2i_2 U520 ( .x(n3159), .a(n1916), .b(n530) );
    inv_5 U521 ( .x(n1313), .a(n3059) );
    inv_8 U522 ( .x(n3358), .a(n3356) );
    oai22_3 U523 ( .x(n3516), .a(n1649), .b(n1651), .c(n3517), .d(n891) );
    inv_2 U524 ( .x(n3513), .a(n3863) );
    nand2i_2 U525 ( .x(n3512), .a(n3513), .b(n3514) );
    inv_5 U526 ( .x(n3413), .a(n3410) );
    oai22_1 U527 ( .x(n850), .a(n915), .b(n1649), .c(n508), .d(n815) );
    inv_5 U528 ( .x(n3411), .a(n3544) );
    nor2_1 U529 ( .x(n1415), .a(n1087), .b(n4020) );
    nor2_5 U53 ( .x(n775), .a(Imm[18]), .b(Imm[21]) );
    nor2i_2 U530 ( .x(n1414), .a(n502), .b(n720) );
    nand2i_2 U531 ( .x(n3975), .a(n719), .b(n3457) );
    inv_2 U532 ( .x(n1392), .a(n2991) );
    nand4_1 U533 ( .x(n3981), .a(n3980), .b(n3979), .c(n3978), .d(n3977) );
    nand2i_2 U534 ( .x(n3978), .a(n1634), .b(n521) );
    inv_2 U535 ( .x(n3140), .a(n3981) );
    nor2i_1 U536 ( .x(n1409), .a(N1840), .b(n946) );
    nand2i_2 U537 ( .x(n3968), .a(n1608), .b(n3638) );
    nand4i_1 U538 ( .x(n1397), .a(n1360), .b(n3968), .c(n3967), .d(n3966) );
    nor2i_1 U539 ( .x(n1408), .a(N1741), .b(___cell__39620_net143710) );
    inv_3 U54 ( .x(n780), .a(Imm[6]) );
    nor2i_1 U540 ( .x(n1405), .a(n1406), .b(___cell__39620_net143658) );
    nor2i_1 U541 ( .x(n1407), .a(N1708), .b(___cell__39620_net143660) );
    inv_2 U542 ( .x(n3848), .a(n3847) );
    nand2i_2 U543 ( .x(n3847), .a(n601), .b(n530) );
    exnor2_1 U544 ( .x(n1490), .a(n583), .b(n745) );
    inv_2 U545 ( .x(n2694), .a(n1490) );
    exnor2_1 U546 ( .x(n1489), .a(n583), .b(reg_out_B[22]) );
    inv_2 U547 ( .x(n2693), .a(n1489) );
    aoi22_1 U548 ( .x(n2692), .a(n2139), .b(n2693), .c(n2193), .d(n2694) );
    nand2i_2 U549 ( .x(n3849), .a(n601), .b(n1064) );
    nor2_1 U55 ( .x(___cell__39620_net145078), .a(Imm[9]), .b(Imm[15]) );
    nand2i_2 U550 ( .x(n2681), .a(___cell__39620_net143735), .b(n663) );
    inv_2 U551 ( .x(n663), .a(n734) );
    inv_2 U552 ( .x(n1811), .a(N1753) );
    nand2i_2 U553 ( .x(n2680), .a(n1811), .b(___cell__39620_net145150) );
    inv_5 U554 ( .x(n3421), .a(n3774) );
    inv_5 U555 ( .x(n1324), .a(n2766) );
    nand2i_2 U556 ( .x(n2679), .a(n1055), .b(n2600) );
    nor2i_0 U558 ( .x(n2674), .a(n745), .b(n1570) );
    nand2_2 U559 ( .x(n3818), .a(n3480), .b(___cell__39620_net144331) );
    nor2_0 U56 ( .x(n1979), .a(Imm[22]), .b(Imm[23]) );
    aoi21_1 U560 ( .x(n1130), .a(n1131), .b(n1132), .c(n816) );
    nand2i_2 U561 ( .x(n1131), .a(n702), .b(n2136) );
    nand2i_2 U562 ( .x(n1132), .a(___cell__39620_net144406), .b(n750) );
    nand2i_2 U563 ( .x(n3708), .a(n759), .b(n530) );
    inv_2 U564 ( .x(n3709), .a(n3708) );
    exnor2_1 U565 ( .x(n1466), .a(n912), .b(reg_out_B[5]) );
    nand2i_2 U566 ( .x(n2210), .a(n4041), .b(n3057) );
    oai211_2 U567 ( .x(n3689), .a(n3505), .b(n718), .c(n2126), .d(n2127) );
    oai22_1 U568 ( .x(n2205), .a(___cell__39620_net144326), .b(n4002), .c(
        n2206), .d(n1654) );
    inv_2 U569 ( .x(n2366), .a(n2148) );
    nor2_1 U57 ( .x(n1980), .a(Imm[25]), .b(Imm[27]) );
    nand2i_2 U570 ( .x(n2204), .a(n1646), .b(n2148) );
    nand2i_2 U571 ( .x(n2203), .a(n759), .b(n1064) );
    aoi21_1 U572 ( .x(n2132), .a(n1249), .b(n2133), .c(n2131) );
    aoi21_1 U573 ( .x(n2129), .a(n1714), .b(n2130), .c(n1110) );
    nand3_1 U574 ( .x(n3693), .a(n2129), .b(n3692), .c(n2132) );
    inv_5 U575 ( .x(net151578), .a(net151577) );
    inv_2 U576 ( .x(n1125), .a(N1868) );
    nor2_1 U577 ( .x(n1124), .a(n947), .b(n1125) );
    nor2i_3 U578 ( .x(n1297), .a(n650), .b(n1298) );
    inv_2 U579 ( .x(n2630), .a(n3570) );
    inv_2 U58 ( .x(n688), .a(Imm[25]) );
    oai211_1 U580 ( .x(n743), .a(n3600), .b(n1565), .c(n3845), .d(n2672) );
    nand2i_2 U581 ( .x(n3874), .a(n1843), .b(n530) );
    inv_2 U582 ( .x(n3875), .a(n3874) );
    nand2i_2 U583 ( .x(n2870), .a(n1843), .b(n1064) );
    oai21_1 U584 ( .x(n2869), .a(___cell__39620_net143693), .b(n683), .c(n2870
        ) );
    inv_4 U585 ( .x(n1268), .a(n2872) );
    nand2i_2 U586 ( .x(n3519), .a(n3520), .b(n3521) );
    and2_1 U588 ( .x(n732), .a(ALU_result[19]), .b(n3057) );
    inv_2 U589 ( .x(n1292), .a(N1816) );
    nand2i_3 U59 ( .x(n1729), .a(n1043), .b(n1685) );
    nor2_1 U590 ( .x(n1291), .a(n1077), .b(n1292) );
    inv_2 U592 ( .x(n1846), .a(N1717) );
    nand2i_2 U593 ( .x(n2844), .a(n1846), .b(___cell__39620_net145190) );
    nor2i_0 U594 ( .x(n2839), .a(n684), .b(n1583) );
    inv_2 U595 ( .x(n1847), .a(N1750) );
    nand2i_2 U596 ( .x(n3440), .a(n4003), .b(n1977) );
    nand2i_3 U597 ( .x(n3606), .a(n3605), .b(n3598) );
    inv_5 U598 ( .x(n3442), .a(n2236) );
    nand2i_0 U599 ( .x(n1144), .a(n1649), .b(n530) );
    inv_2 U60 ( .x(n3573), .a(n1729) );
    aoi21_1 U600 ( .x(n1142), .a(n1143), .b(n1144), .c(n855) );
    nor2i_1 U601 ( .x(n2212), .a(n1085), .b(n816) );
    nor2i_1 U602 ( .x(n2211), .a(___cell__39620_net144345), .b(n1658) );
    exnor2_1 U603 ( .x(n1468), .a(reg_out_B[4]), .b(n834) );
    exnor2_1 U604 ( .x(n1467), .a(n834), .b(net151904) );
    nor2_1 U605 ( .x(n1145), .a(n679), .b(n4040) );
    nand2i_2 U606 ( .x(n2255), .a(n621), .b(n2371) );
    nand2i_2 U607 ( .x(n2252), .a(n1646), .b(n3705) );
    nand2i_2 U608 ( .x(n2251), .a(n1657), .b(n2148) );
    inv_5 U609 ( .x(___cell__39620_net145617), .a(___cell__39620_net143693) );
    nand2_2 U61 ( .x(n1835), .a(n3573), .b(n910) );
    nand2_0 U610 ( .x(n2249), .a(___cell__39620_net145617), .b(net151904) );
    nand3_2 U611 ( .x(n2247), .a(n2180), .b(n3700), .c(n2178) );
    nand2i_2 U612 ( .x(n3700), .a(___cell__39620_net144062), .b(n2337) );
    nor2i_1 U613 ( .x(n1137), .a(N1702), .b(___cell__39620_net143660) );
    nand2i_2 U614 ( .x(n3507), .a(n4006), .b(n1049) );
    nor2i_0 U615 ( .x(n2215), .a(net151904), .b(n1649) );
    inv_5 U616 ( .x(n1649), .a(n834) );
    inv_2 U617 ( .x(n672), .a(n1047) );
    oai211_2 U618 ( .x(n3687), .a(n1334), .b(___cell__39620_net144317), .c(
        n2069), .d(n3686) );
    inv_5 U619 ( .x(n3510), .a(n3687) );
    nand2_0 U62 ( .x(n3630), .a(___cell__39620_net144330), .b(n541) );
    nor2i_1 U620 ( .x(n1123), .a(n1045), .b(n4006) );
    inv_12 U621 ( .x(n1607), .a(n673) );
    inv_8 U622 ( .x(n885), .a(n1654) );
    inv_12 U623 ( .x(n586), .a(n1417) );
    inv_2 U625 ( .x(n3299), .a(n2927) );
    ao22_1 U626 ( .x(n3552), .a(reg_out_A[8]), .b(n3575), .c(n2277), .d(n799)
         );
    oai221_2 U627 ( .x(n2875), .a(n3553), .b(___cell__39620_net144374), .c(
        n3299), .d(n1623), .e(n2853) );
    aoi23_1 U628 ( .x(n2850), .a(n1249), .b(n2852), .c(n879), .d(n2851), .e(
        reg_out_B[2]) );
    inv_5 U629 ( .x(n3522), .a(n3519) );
    nand2i_2 U63 ( .x(n1673), .a(reg_out_B[3]), .b(reg_out_B[4]) );
    nand2i_2 U630 ( .x(n2894), .a(n621), .b(n2930) );
    exnor2_1 U631 ( .x(n1499), .a(n910), .b(n633) );
    inv_2 U632 ( .x(n1311), .a(n1499) );
    nor2i_1 U633 ( .x(n1310), .a(n1311), .b(n690) );
    oai21_1 U636 ( .x(n3374), .a(n815), .b(n528), .c(n3375) );
    and2_1 U637 ( .x(n697), .a(n767), .b(n3381) );
    inv_4 U638 ( .x(n3381), .a(n853) );
    inv_2 U639 ( .x(n3889), .a(n3888) );
    nand2i_1 U64 ( .x(n3449), .a(n1219), .b(n1689) );
    inv_2 U640 ( .x(n1854), .a(N1948) );
    inv_2 U641 ( .x(n1855), .a(N1815) );
    nand2i_2 U642 ( .x(n3859), .a(n1608), .b(n3774) );
    inv_2 U643 ( .x(n2634), .a(n3569) );
    aoi21_2 U644 ( .x(n2765), .a(n2676), .b(n2766), .c(n2634) );
    nand2_2 U645 ( .x(n2877), .a(n633), .b(n910) );
    oai22_1 U646 ( .x(n2878), .a(n1602), .b(n734), .c(___cell__39620_net143658
        ), .d(n2877) );
    inv_4 U648 ( .x(n1306), .a(N1881) );
    nand2i_2 U649 ( .x(n3869), .a(n1608), .b(n3790) );
    nand2_0 U65 ( .x(n3635), .a(___cell__39620_net144330), .b(n590) );
    nand2i_4 U650 ( .x(n2310), .a(n1734), .b(___cell__39620_net145508) );
    inv_4 U651 ( .x(n1734), .a(N1993) );
    nand2_2 U652 ( .x(n2307), .a(Imm[30]), .b(n535) );
    nand2i_2 U653 ( .x(n2309), .a(n2307), .b(___cell__39620_net147791) );
    inv_2 U654 ( .x(n1735), .a(N1960) );
    nand2i_2 U655 ( .x(n2311), .a(n1735), .b(n3999) );
    nor2i_1 U656 ( .x(n1161), .a(n1095), .b(n1162) );
    inv_8 U657 ( .x(n3524), .a(n3744) );
    nand2i_2 U658 ( .x(n2316), .a(n1737), .b(n3624) );
    inv_2 U659 ( .x(n1737), .a(N2026) );
    nand2_0 U66 ( .x(n3653), .a(___cell__39620_net144330), .b(n540) );
    nand2i_0 U661 ( .x(n3749), .a(n1731), .b(n1064) );
    inv_10 U662 ( .x(n1731), .a(reg_out_B[30]) );
    ao221_4 U663 ( .x(n1733), .a(n737), .b(n597), .c(n598), .d(n599), .e(n1700
        ) );
    nand2i_0 U664 ( .x(n3747), .a(n1731), .b(n530) );
    nand3i_1 U665 ( .x(n2318), .a(n1732), .b(n3747), .c(n3216) );
    inv_2 U666 ( .x(n3748), .a(n1471) );
    nand2_2 U667 ( .x(n2321), .a(n2193), .b(n3748) );
    oai211_1 U668 ( .x(n2320), .a(n578), .b(n1566), .c(n2321), .d(n2322) );
    nand2i_0 U669 ( .x(n2300), .a(___cell__39620_net144175), .b(n1576) );
    inv_10 U67 ( .x(___cell__39620_net144330), .a(___cell__39620_net144329) );
    inv_5 U670 ( .x(n1576), .a(n1160) );
    inv_2 U671 ( .x(n725), .a(n815) );
    nor2i_1 U672 ( .x(___cell__39620_net145451), .a(n504), .b(n670) );
    inv_12 U673 ( .x(n1587), .a(reg_out_A[27]) );
    exnor2_1 U674 ( .x(n1477), .a(reg_out_A[28]), .b(Imm[28]) );
    exnor2_1 U675 ( .x(n1478), .a(reg_out_A[28]), .b(reg_out_B[28]) );
    inv_2 U676 ( .x(n3267), .a(n1478) );
    nor2i_5 U677 ( .x(n1190), .a(n1191), .b(n578) );
    inv_2 U678 ( .x(n2411), .a(n3775) );
    oai22_1 U679 ( .x(n1732), .a(n621), .b(n1093), .c(n1641), .d(n1089) );
    inv_2 U68 ( .x(n1647), .a(n942) );
    nand2i_2 U680 ( .x(n2448), .a(___cell__39620_net144257), .b(n2489) );
    inv_5 U681 ( .x(n3419), .a(n2719) );
    nand2i_2 U682 ( .x(n2447), .a(n1574), .b(n2399) );
    oai21_3 U683 ( .x(n2492), .a(n3418), .b(n1565), .c(n3571) );
    nor2_1 U684 ( .x(n1192), .a(n679), .b(n4035) );
    nand4_1 U685 ( .x(n2457), .a(n2437), .b(n3771), .c(n2434), .d(n3770) );
    nand2i_2 U686 ( .x(n3771), .a(___cell__39620_net144062), .b(n2302) );
    aoi22_1 U687 ( .x(n2434), .a(n2435), .b(n2262), .c(n2436), .d(n904) );
    aoi21_1 U688 ( .x(n2430), .a(n1256), .b(n2306), .c(n2428) );
    nand2i_2 U689 ( .x(n3769), .a(n1636), .b(n2305) );
    nand2i_2 U69 ( .x(n3561), .a(n1647), .b(n873) );
    nor2_1 U690 ( .x(n1083), .a(n4002), .b(___cell__39620_net143694) );
    nand2_2 U691 ( .x(n3665), .a(n1391), .b(n3451) );
    inv_5 U692 ( .x(n2022), .a(n1626) );
    inv_5 U693 ( .x(n3314), .a(n2136) );
    nand2_2 U694 ( .x(n3666), .a(n1256), .b(n2133) );
    oai211_1 U695 ( .x(n2046), .a(n1082), .b(n1664), .c(n2047), .d(n2048) );
    nand2_2 U696 ( .x(n2047), .a(n2193), .b(n3676) );
    inv_2 U697 ( .x(n3676), .a(n1460) );
    nand2i_2 U698 ( .x(n3670), .a(n1565), .b(n3278) );
    nand2i_2 U699 ( .x(n3671), .a(n1559), .b(n3622) );
    nand2i_2 U70 ( .x(n3293), .a(n1657), .b(n873) );
    inv_2 U700 ( .x(n1078), .a(N1805) );
    nor2_1 U701 ( .x(n1076), .a(n1077), .b(n1078) );
    nand2i_2 U702 ( .x(n3673), .a(n4005), .b(n1136) );
    nand2i_2 U703 ( .x(n3675), .a(n1608), .b(n3538) );
    nor2i_2 U704 ( .x(n1071), .a(n1042), .b(n1072) );
    inv_5 U705 ( .x(___cell__39620_net144303), .a(___cell__39620_net144302) );
    nor2i_0 U706 ( .x(n1074), .a(n914), .b(___cell__39620_net143694) );
    nor2i_1 U707 ( .x(n1073), .a(n1074), .b(___cell__39620_net143658) );
    nor2i_0 U708 ( .x(n1075), .a(N1706), .b(___cell__39620_net143660) );
    oai211_1 U709 ( .x(n2396), .a(n505), .b(___cell__39620_net144257), .c(
        n2397), .d(n2398) );
    inv_5 U71 ( .x(n873), .a(n1622) );
    nand2_2 U710 ( .x(n2398), .a(n2193), .b(n3768) );
    inv_2 U711 ( .x(n3768), .a(n1475) );
    aoi22_1 U712 ( .x(n2304), .a(n1714), .b(n2305), .c(n1249), .d(n2306) );
    oai21_1 U713 ( .x(n2324), .a(n816), .b(n3731), .c(n2304) );
    oai22_5 U714 ( .x(n2303), .a(n1585), .b(n836), .c(n3462), .d(n4125) );
    oai21_2 U715 ( .x(n2456), .a(n1564), .b(n1093), .c(n3761) );
    nand2i_2 U716 ( .x(n2409), .a(n621), .b(n2456) );
    oai21_1 U717 ( .x(n2455), .a(n1564), .b(n695), .c(___cell__39620_net147350
        ) );
    nand2i_2 U718 ( .x(n2406), .a(n1747), .b(n1064) );
    oai21_1 U719 ( .x(n2405), .a(n4002), .b(___cell__39620_net144605), .c(
        n2406) );
    nand2i_2 U72 ( .x(n3305), .a(___cell__39620_net144257), .b(n873) );
    inv_2 U720 ( .x(n717), .a(net149122) );
    inv_2 U722 ( .x(n3409), .a(n2287) );
    aoi22_1 U723 ( .x(n2372), .a(n1714), .b(n2286), .c(n1249), .d(n2373) );
    nand2i_2 U724 ( .x(n3766), .a(n1747), .b(n530) );
    inv_0 U725 ( .x(n1747), .a(reg_out_B[29]) );
    inv_2 U726 ( .x(net151497), .a(IR_opcode_field[3]) );
    inv_2 U727 ( .x(___cell__39620_net144309), .a(___cell__39620_net144307) );
    or2_1 U728 ( .x(n495), .a(IR_opcode_field[0]), .b(IR_opcode_field[3]) );
    nand2i_2 U729 ( .x(___cell__39620_net144307), .a(n495), .b(
        ___cell__39620_net143655) );
    nand2i_2 U73 ( .x(n3371), .a(n1561), .b(n926) );
    nand2_0 U730 ( .x(n2376), .a(Imm[29]), .b(n539) );
    inv_5 U731 ( .x(n1290), .a(n2633) );
    inv_5 U732 ( .x(n3427), .a(n3726) );
    oai21_1 U733 ( .x(n3727), .a(n891), .b(n3427), .c(n4140) );
    inv_12 U734 ( .x(n662), .a(n1182) );
    nor2_0 U735 ( .x(n1181), .a(n4140), .b(n1182) );
    nor2i_1 U736 ( .x(n782), .a(Imm[31]), .b(___cell__39620_net143693) );
    inv_2 U737 ( .x(n3520), .a(n3721) );
    inv_4 U738 ( .x(n3594), .a(n890) );
    oai21_1 U739 ( .x(n2274), .a(n1648), .b(n1281), .c(n2275) );
    nand2i_2 U74 ( .x(n3370), .a(n1564), .b(n874) );
    nand2i_4 U740 ( .x(n2280), .a(n3486), .b(n3487) );
    oai211_3 U741 ( .x(n2279), .a(n3397), .b(___cell__39620_net144317), .c(
        n3398), .d(n3399) );
    aoi22_1 U742 ( .x(n2282), .a(n1971), .b(n2283), .c(n1177), .d(n2284) );
    nand2_2 U743 ( .x(n2287), .a(n3473), .b(n3474) );
    aoi222_1 U744 ( .x(n2285), .a(n1256), .b(n2286), .c(n1150), .d(n2287), .e(
        n2273), .f(n644) );
    nand3_1 U745 ( .x(n734), .a(n733), .b(n1520), .c(___cell__39620_net144355)
         );
    aoi21_1 U746 ( .x(n517), .a(n671), .b(n3726), .c(n626) );
    nor2_0 U747 ( .x(n795), .a(net151904), .b(net149167) );
    inv_8 U748 ( .x(___cell__39620_net143326), .a(___cell__39620_net147731) );
    nand2_0 U749 ( .x(___cell__39620_net147296), .a(n1658), .b(n1641) );
    nor2_0 U75 ( .x(n2002), .a(IR_function_field[2]), .b(IR_function_field[3])
         );
    inv_2 U750 ( .x(n835), .a(n3740) );
    nand2i_2 U751 ( .x(n3728), .a(n1085), .b(n621) );
    nand3i_1 U752 ( .x(n2289), .a(n1636), .b(n3728), .c(
        ___cell__39620_net145472) );
    nand2i_2 U753 ( .x(n3736), .a(N70), .b(n530) );
    inv_2 U754 ( .x(n3737), .a(n3736) );
    inv_5 U755 ( .x(___cell__39620_net144344), .a(___cell__39620_net144340) );
    or3i_1 U756 ( .x(___cell__39620_net144350), .a(___cell__39620_net144344), 
        .b(n783), .c(___cell__39620_net143653) );
    nand2i_2 U757 ( .x(n770), .a(___cell__39620_net144350), .b(
        ___cell__39620_net147732) );
    nand2_2 U758 ( .x(n2258), .a(reg_out_A[31]), .b(Imm[31]) );
    exnor2_1 U759 ( .x(n1469), .a(reg_out_A[31]), .b(Imm[31]) );
    oai21_1 U760 ( .x(n2291), .a(n1469), .b(n690), .c(n2292) );
    aoi21_1 U761 ( .x(n2272), .a(n2273), .b(n609), .c(n1149) );
    nand2i_2 U762 ( .x(n3732), .a(n1634), .b(n2305) );
    nand4_1 U763 ( .x(n3730), .a(n2269), .b(n3729), .c(n2267), .d(n3375) );
    oai211_1 U764 ( .x(n2290), .a(n3731), .b(n1451), .c(n3732), .d(n2272) );
    nand2i_2 U765 ( .x(n2294), .a(N70), .b(n1064) );
    inv_4 U766 ( .x(n3735), .a(n1154) );
    nand2_2 U767 ( .x(n1155), .a(n2263), .b(n2264) );
    nand4i_1 U768 ( .x(n1154), .a(n2259), .b(n3733), .c(n2261), .d(n3734) );
    aoi21_1 U769 ( .x(n1153), .a(net149120), .b(n1154), .c(n1155) );
    nand2i_2 U77 ( .x(n1960), .a(reg_out_B[28]), .b(n1959) );
    nand3i_1 U770 ( .x(n1662), .a(n2004), .b(n1590), .c(n2005) );
    nand2_2 U771 ( .x(n2005), .a(n2003), .b(n3593) );
    aoi22_1 U772 ( .x(n2006), .a(n1526), .b(n1534), .c(n1540), .d(n1530) );
    inv_5 U773 ( .x(n3506), .a(n3695) );
    inv_2 U774 ( .x(n1927), .a(N1931) );
    nand2i_2 U775 ( .x(n3194), .a(n1927), .b(n3999) );
    nand2i_2 U776 ( .x(n3193), .a(n1928), .b(n1987) );
    inv_2 U777 ( .x(n1928), .a(N1798) );
    nand2i_3 U778 ( .x(n3986), .a(___cell__39620_net144345), .b(n1165) );
    nand2i_4 U779 ( .x(n3245), .a(n3185), .b(n3986) );
    inv_5 U78 ( .x(n601), .a(reg_out_B[22]) );
    inv_2 U780 ( .x(n1926), .a(N1732) );
    nand2i_2 U781 ( .x(n3189), .a(n1926), .b(___cell__39620_net145150) );
    aoi21_1 U782 ( .x(n3188), .a(N1699), .b(___cell__39620_net145190), .c(
        n1420) );
    inv_2 U783 ( .x(n1925), .a(N1633) );
    oai211_1 U784 ( .x(n3187), .a(___cell__39620_net143872), .b(n1925), .c(
        n3188), .d(n3189) );
    nor2i_1 U785 ( .x(n3181), .a(n694), .b(n1657) );
    exnor2_1 U786 ( .x(n1517), .a(n917), .b(net149122) );
    inv_2 U787 ( .x(n3504), .a(n3279) );
    aoi22_1 U788 ( .x(n2808), .a(n1714), .b(n2809), .c(n1249), .d(n2130) );
    exnor2_1 U789 ( .x(n1518), .a(n816), .b(n917) );
    nand2i_2 U790 ( .x(n3432), .a(n1562), .b(n3622) );
    inv_2 U791 ( .x(n3557), .a(n3555) );
    nand2i_2 U792 ( .x(n3431), .a(n4003), .b(n3278) );
    oai221_1 U793 ( .x(n3177), .a(n3178), .b(n1687), .c(n1657), .d(n1093), .e(
        n3179) );
    nand2i_3 U794 ( .x(n3984), .a(n1451), .b(n3752) );
    nand2_2 U795 ( .x(n1660), .a(n701), .b(n1661) );
    nand2_0 U796 ( .x(n3218), .a(___cell__39620_net145617), .b(net149122) );
    nand2i_2 U797 ( .x(n3217), .a(n4019), .b(n3057) );
    nand2i_2 U798 ( .x(n1640), .a(net152465), .b(IR_opcode_field[1]) );
    aoi22_1 U799 ( .x(n3200), .a(n2079), .b(n3201), .c(n3202), .d(n917) );
    nand2i_2 U800 ( .x(n3201), .a(n622), .b(n3488) );
    inv_2 U801 ( .x(n3489), .a(n3201) );
    aoi22_1 U802 ( .x(n3199), .a(n2266), .b(n902), .c(n1066), .d(n2337) );
    inv_4 U803 ( .x(n3753), .a(n1738) );
    inv_2 U804 ( .x(n2335), .a(n1281) );
    inv_2 U805 ( .x(n599), .a(n696) );
    oai221_1 U806 ( .x(n3197), .a(n1417), .b(n1690), .c(n1657), .d(n1093), .e(
        n3198) );
    nand2i_2 U807 ( .x(n3985), .a(n1451), .b(n3755) );
    inv_2 U808 ( .x(n1543), .a(n1541) );
    nand2i_2 U809 ( .x(n1452), .a(n496), .b(n1543) );
    inv_8 U81 ( .x(n628), .a(n1561) );
    inv_2 U810 ( .x(n3612), .a(n3564) );
    inv_2 U811 ( .x(n3178), .a(n1966) );
    inv_2 U812 ( .x(n3344), .a(n3348) );
    or2_1 U813 ( .x(n522), .a(n569), .b(n1569) );
    inv_2 U814 ( .x(n3601), .a(n522) );
    inv_2 U815 ( .x(n3316), .a(n3320) );
    inv_2 U816 ( .x(n3326), .a(n3329) );
    inv_2 U817 ( .x(n3663), .a(n1458) );
    nand2_2 U818 ( .x(n2008), .a(n2193), .b(n3663) );
    aoi21_1 U819 ( .x(n1062), .a(n904), .b(n530), .c(n1064) );
    nand2_0 U82 ( .x(n3625), .a(___cell__39620_net144330), .b(reg_out_A[28])
         );
    inv_2 U820 ( .x(n3621), .a(n3500) );
    inv_2 U821 ( .x(n3333), .a(n3338) );
    oai22_1 U822 ( .x(n3414), .a(n915), .b(n1649), .c(n508), .d(n815) );
    nand2i_2 U823 ( .x(n3586), .a(n1632), .b(n521) );
    nand2_1 U824 ( .x(n3587), .a(n1714), .b(n2187) );
    nand3_1 U825 ( .x(n2027), .a(n3587), .b(n3586), .c(n1998) );
    nand4_3 U826 ( .x(n3583), .a(n3582), .b(n3580), .c(n3579), .d(n3581) );
    nand2i_2 U827 ( .x(n3581), .a(n1625), .b(n3457) );
    ao22_5 U828 ( .x(n2233), .a(n3318), .b(n857), .c(n814), .d(n3584) );
    inv_5 U829 ( .x(n722), .a(n3317) );
    nand2_0 U83 ( .x(n3636), .a(___cell__39620_net144330), .b(reg_out_A[29])
         );
    nand2i_2 U830 ( .x(n3590), .a(n1623), .b(n4127) );
    nand2i_2 U831 ( .x(n2031), .a(n4045), .b(n3057) );
    nand2i_2 U833 ( .x(n3659), .a(n1607), .b(n3655) );
    nand2i_2 U834 ( .x(n3660), .a(n4007), .b(n1349) );
    nand2i_2 U835 ( .x(n3661), .a(n1608), .b(n3658) );
    nor2i_3 U836 ( .x(n1048), .a(n1049), .b(n4005) );
    nand2i_2 U837 ( .x(n3650), .a(n4006), .b(n3475) );
    nor2i_3 U838 ( .x(n1046), .a(n1047), .b(n1043) );
    nand4i_2 U839 ( .x(n1054), .a(n1046), .b(n3651), .c(n3650), .d(n3649) );
    nor2i_1 U84 ( .x(n1280), .a(n583), .b(n1281) );
    nor2i_1 U840 ( .x(n1050), .a(n1051), .b(___cell__39620_net143658) );
    nor2i_1 U841 ( .x(n1052), .a(N1707), .b(___cell__39620_net143660) );
    inv_2 U842 ( .x(n3018), .a(n3956) );
    nand2i_2 U843 ( .x(n3956), .a(n703), .b(n3931) );
    nor2_1 U844 ( .x(n1347), .a(n679), .b(n4023) );
    nand4_1 U845 ( .x(n3056), .a(n3947), .b(n3946), .c(n3945), .d(n3944) );
    nand2i_2 U846 ( .x(n3017), .a(n784), .b(n3056) );
    nand2i_2 U847 ( .x(n3016), .a(n1658), .b(n3926) );
    inv_2 U848 ( .x(n713), .a(___cell__39620_net144062) );
    nand2i_4 U85 ( .x(n2128), .a(n547), .b(n3463) );
    aoi22_1 U850 ( .x(n2990), .a(___cell__39620_net144517), .b(n2991), .c(
        n1391), .d(n2992) );
    nand2i_2 U851 ( .x(n3943), .a(n1625), .b(n3069) );
    oai211_1 U852 ( .x(n3008), .a(n630), .b(___cell__39620_net144062), .c(
        n3943), .d(n2990) );
    nand2i_2 U853 ( .x(n3949), .a(n1634), .b(n3544) );
    nand2i_2 U854 ( .x(n3950), .a(n727), .b(n2851) );
    nand2i_2 U855 ( .x(n3951), .a(n1635), .b(n2852) );
    nand4_1 U856 ( .x(n3013), .a(n3951), .b(n3950), .c(n3949), .d(n3948) );
    aoi22_2 U857 ( .x(n2993), .a(n1714), .b(n2994), .c(n1256), .d(n2995) );
    nand2i_2 U858 ( .x(n3942), .a(n1632), .b(n3302) );
    inv_12 U859 ( .x(n3584), .a(n822) );
    aoi21_1 U86 ( .x(n2804), .a(n1289), .b(n2128), .c(n1280) );
    oai211_1 U860 ( .x(n3012), .a(n3355), .b(n1636), .c(n3942), .d(n2993) );
    inv_5 U861 ( .x(n3439), .a(n3606) );
    inv_2 U862 ( .x(n3955), .a(n1506) );
    nand2_2 U863 ( .x(n2997), .a(n2193), .b(n3955) );
    aoi21_1 U864 ( .x(n1346), .a(n609), .b(n530), .c(n1064) );
    oai211_1 U865 ( .x(n2996), .a(n1346), .b(n1874), .c(n2997), .d(n2998) );
    inv_0 U866 ( .x(n1358), .a(reg_out_B[14]) );
    inv_2 U867 ( .x(n1881), .a(N1845) );
    inv_2 U868 ( .x(n1341), .a(N1812) );
    nor2_1 U869 ( .x(n1340), .a(n1077), .b(n1341) );
    nand2i_2 U87 ( .x(n2340), .a(n1635), .b(n3196) );
    nand2i_2 U870 ( .x(n3952), .a(n1607), .b(n3790) );
    nand2i_3 U871 ( .x(n3954), .a(n1608), .b(n3648) );
    nand4i_1 U872 ( .x(n2988), .a(n1332), .b(n3954), .c(n3953), .d(n3952) );
    nor2i_1 U873 ( .x(n1336), .a(net151622), .b(n1585) );
    nor2i_1 U874 ( .x(n1335), .a(n1336), .b(___cell__39620_net143658) );
    nor2i_1 U875 ( .x(n1337), .a(N1713), .b(___cell__39620_net143660) );
    and4i_2 U876 ( .x(n766), .a(n568), .b(N3304), .c(___cell__39620_net144303), 
        .d(n1619) );
    nor2_0 U877 ( .x(n1327), .a(n4002), .b(___cell__39620_net143962) );
    nand4_1 U878 ( .x(n3009), .a(n3917), .b(n3916), .c(n3915), .d(n3914) );
    nand4_1 U879 ( .x(n3931), .a(n3930), .b(n3929), .c(n3928), .d(n3927) );
    nand2i_2 U880 ( .x(n2974), .a(___cell__39620_net144406), .b(n3931) );
    nand4_1 U881 ( .x(n3926), .a(n3925), .b(n3924), .c(n3923), .d(n3922) );
    ao22_3 U882 ( .x(n2977), .a(n3903), .b(n700), .c(n3926), .d(n757) );
    nand2i_2 U883 ( .x(n2979), .a(n4001), .b(n3897) );
    nor2_1 U884 ( .x(n1328), .a(n679), .b(n4024) );
    oai211_1 U885 ( .x(n2958), .a(n1326), .b(n1866), .c(n2959), .d(n2960) );
    aoi21_1 U886 ( .x(n1326), .a(n893), .b(n530), .c(n1064) );
    nand2_2 U887 ( .x(n2959), .a(n2193), .b(n3941) );
    inv_2 U888 ( .x(n3941), .a(n1504) );
    nand2i_2 U889 ( .x(n3933), .a(n1565), .b(n3622) );
    inv_8 U89 ( .x(n939), .a(n938) );
    inv_2 U890 ( .x(n1870), .a(N1879) );
    nand2i_2 U891 ( .x(n2952), .a(n1870), .b(n3998) );
    aoi211_1 U892 ( .x(n2948), .a(N1648), .b(n809), .c(n1325), .d(
        ___cell__39620_net146132) );
    nor2i_1 U893 ( .x(n1325), .a(N1714), .b(___cell__39620_net143660) );
    oai22_1 U894 ( .x(___cell__39620_net146132), .a(n783), .b(n734), .c(
        ___cell__39620_net143658), .d(___cell__39620_net146131) );
    inv_2 U895 ( .x(n1869), .a(N1747) );
    nand2i_2 U896 ( .x(n2951), .a(n1869), .b(___cell__39620_net145150) );
    aoi22_1 U897 ( .x(n2953), .a(N1979), .b(___cell__39620_net145508), .c(
        N1846), .d(n4000) );
    nand2i_2 U898 ( .x(n2957), .a(n1872), .b(n1987) );
    inv_2 U899 ( .x(n1872), .a(N1813) );
    buf_2 U90 ( .x(net149106), .a(Imm[1]) );
    nand2i_2 U900 ( .x(n2955), .a(n1616), .b(n1339) );
    and3i_1 U901 ( .x(n2914), .a(n2913), .b(n2915), .c(n2916) );
    nand2i_2 U902 ( .x(n2916), .a(n1860), .b(___cell__39620_net145190) );
    inv_2 U903 ( .x(n1860), .a(N1715) );
    oai22_1 U904 ( .x(n2913), .a(___cell__39620_net143872), .b(n1859), .c(
        ___cell__39620_net143658), .d(n2912) );
    inv_2 U905 ( .x(n1859), .a(N1649) );
    inv_2 U906 ( .x(n1862), .a(N1880) );
    nand2i_2 U907 ( .x(n2919), .a(n1862), .b(n944) );
    nor2i_1 U908 ( .x(n1316), .a(n694), .b(n734) );
    aoi22_1 U909 ( .x(n2924), .a(N1847), .b(n4000), .c(N1980), .d(
        ___cell__39620_net145508) );
    nand2i_2 U91 ( .x(n3698), .a(n1644), .b(n530) );
    nand2i_2 U910 ( .x(n2923), .a(n1864), .b(n1987) );
    inv_2 U911 ( .x(n1864), .a(N1814) );
    nand2i_2 U912 ( .x(n2922), .a(n1166), .b(n1339) );
    nand2i_2 U913 ( .x(n2921), .a(n1616), .b(n1308) );
    aoi21_2 U914 ( .x(n2762), .a(n1177), .b(n2763), .c(n2630) );
    inv_2 U915 ( .x(n3618), .a(n3405) );
    oai211_3 U916 ( .x(n2902), .a(n3620), .b(n1565), .c(n3857), .d(n2762) );
    nand2i_2 U917 ( .x(n3865), .a(n1562), .b(n2629) );
    nand2i_2 U918 ( .x(n3866), .a(n1565), .b(n3606) );
    inv_1 U919 ( .x(n827), .a(n761) );
    inv_2 U92 ( .x(n911), .a(reg_out_A[5]) );
    nand2i_2 U920 ( .x(n2929), .a(n1064), .b(n3913) );
    nand2i_2 U921 ( .x(n2934), .a(n1626), .b(n3887) );
    nand2i_2 U922 ( .x(n2933), .a(n1566), .b(n3004) );
    inv_1 U923 ( .x(net156025), .a(net156024) );
    inv_2 U924 ( .x(n638), .a(net156025) );
    oai21_1 U925 ( .x(n2932), .a(n1501), .b(n690), .c(n2935) );
    nand2i_2 U926 ( .x(n3896), .a(n1623), .b(n3547) );
    inv_5 U927 ( .x(n2943), .a(n2911) );
    nand2i_2 U928 ( .x(n3876), .a(n719), .b(n2784) );
    oai22_1 U929 ( .x(n2945), .a(n1087), .b(n4025), .c(n1217), .d(n1417) );
    exnor2_1 U93 ( .x(n1512), .a(reg_out_B[12]), .b(n894) );
    nand2i_2 U930 ( .x(n3878), .a(n1636), .b(n2781) );
    ao21_2 U931 ( .x(n516), .a(n1267), .b(n2938), .c(n1320) );
    nor2_1 U932 ( .x(n1320), .a(___cell__39620_net143693), .b(
        ___cell__39620_net143954) );
    nand2i_2 U933 ( .x(n3898), .a(n727), .b(n2994) );
    nand2i_2 U934 ( .x(n3899), .a(n1634), .b(n3302) );
    nand2i_2 U935 ( .x(n3900), .a(n1632), .b(n3381) );
    nand2i_2 U936 ( .x(n3850), .a(n4003), .b(n3059) );
    inv_2 U937 ( .x(n3609), .a(n3309) );
    nand2i_4 U938 ( .x(n3610), .a(n3609), .b(n3598) );
    inv_6 U939 ( .x(n2696), .a(n2864) );
    oai22_1 U94 ( .x(n2082), .a(n2083), .b(n1687), .c(n1584), .d(n1690) );
    aoi21_2 U940 ( .x(n2672), .a(n1177), .b(n2673), .c(n2630) );
    inv_2 U941 ( .x(n3597), .a(n3474) );
    oai211_3 U942 ( .x(n2864), .a(n3600), .b(n1565), .c(n3845), .d(n2672) );
    aoai211_1 U943 ( .x(n2743), .a(n1217), .b(n2744), .c(n1561), .d(n2740) );
    inv_2 U944 ( .x(n2741), .a(n1491) );
    inv_2 U945 ( .x(n2742), .a(n1492) );
    mux2_2 U946 ( .x(n2711), .d0(n3378), .sl(n816), .d1(n3382) );
    nand2i_2 U947 ( .x(n2755), .a(___cell__39620_net144765), .b(
        ___cell__39620_net145617) );
    inv_2 U948 ( .x(n3527), .a(n3733) );
    nand2i_2 U949 ( .x(n3526), .a(n3527), .b(n3528) );
    exnor2_1 U95 ( .x(n1479), .a(n533), .b(n681) );
    oai22_1 U950 ( .x(n3379), .a(n1587), .b(n915), .c(n853), .d(n815) );
    aoi21_1 U951 ( .x(n2737), .a(n1714), .b(n2738), .c(n1248) );
    nand2i_2 U952 ( .x(n3852), .a(n1634), .b(n3550) );
    nand2_1 U953 ( .x(n3853), .a(n504), .b(n2477) );
    nand3_1 U954 ( .x(n3854), .a(n3853), .b(n3852), .c(n2737) );
    nand2i_2 U955 ( .x(n3851), .a(n1623), .b(n2854) );
    inv_5 U956 ( .x(n799), .a(Imm[3]) );
    nand2i_2 U957 ( .x(n3843), .a(n1623), .b(n2784) );
    nor2_1 U958 ( .x(n1254), .a(n1087), .b(n4028) );
    aoi22_1 U959 ( .x(n2689), .a(n2690), .b(n1249), .c(n504), .d(n2433) );
    exnor2_1 U96 ( .x(n1480), .a(n533), .b(reg_out_B[27]) );
    nand2i_2 U960 ( .x(n3844), .a(n1634), .b(n2781) );
    oai22_2 U961 ( .x(n2779), .a(n506), .b(n536), .c(n1586), .d(n1629) );
    aoi22_1 U962 ( .x(n2727), .a(n663), .b(Imm[5]), .c(n662), .d(n2600) );
    inv_2 U963 ( .x(n1819), .a(N1719) );
    nand2i_2 U964 ( .x(n2726), .a(n1819), .b(___cell__39620_net145190) );
    oai211_1 U965 ( .x(n3839), .a(n844), .b(n4005), .c(n2632), .d(n3838) );
    nand2i_2 U966 ( .x(n2725), .a(n1055), .b(n3839) );
    nor2i_1 U967 ( .x(n1253), .a(N1851), .b(n946) );
    oai211_3 U968 ( .x(n2733), .a(n3656), .b(n1043), .c(n3846), .d(n2675) );
    inv_2 U969 ( .x(n709), .a(n802) );
    inv_2 U97 ( .x(n1931), .a(N1863) );
    inv_4 U970 ( .x(n1822), .a(N1951) );
    inv_2 U971 ( .x(n2676), .a(n4006) );
    inv_0 U972 ( .x(n1843), .a(reg_out_B[19]) );
    inv_2 U973 ( .x(n605), .a(reg_out_B[19]) );
    inv_5 U974 ( .x(n3550), .a(n752) );
    nand2i_2 U975 ( .x(n3831), .a(n1632), .b(n3550) );
    inv_2 U976 ( .x(n3406), .a(n2284) );
    nand2_2 U977 ( .x(n3832), .a(n1714), .b(n2477) );
    nand2_2 U978 ( .x(n3833), .a(n1256), .b(n2738) );
    inv_2 U979 ( .x(n2565), .a(n2277) );
    nand2i_2 U98 ( .x(n3250), .a(n1931), .b(n3997) );
    inv_5 U980 ( .x(n3454), .a(n2280) );
    inv_2 U981 ( .x(n3565), .a(n3640) );
    nand2i_4 U982 ( .x(n3820), .a(n4010), .b(n2520) );
    inv_16 U984 ( .x(n836), .a(n3575) );
    inv_2 U985 ( .x(n3403), .a(n2779) );
    nand2_2 U986 ( .x(n3822), .a(n1256), .b(n2779) );
    nand2_2 U987 ( .x(n3823), .a(n504), .b(n2306) );
    nand2i_2 U988 ( .x(n3824), .a(n1632), .b(n2781) );
    inv_2 U989 ( .x(n3310), .a(n2271) );
    nand2_0 U99 ( .x(n1621), .a(net152465), .b(IR_opcode_field[1]) );
    inv_2 U990 ( .x(n3534), .a(n3533) );
    inv_2 U991 ( .x(n3380), .a(n3379) );
    inv_8 U992 ( .x(n1561), .a(reg_out_A[21]) );
    exnor2_1 U993 ( .x(n1488), .a(n636), .b(n829) );
    exnor2_1 U994 ( .x(n1487), .a(n636), .b(reg_out_B[23]) );
    inv_2 U995 ( .x(n620), .a(___cell__6067_net21981) );
    nand2i_2 U996 ( .x(n1536), .a(___cell__39620_net144175), .b(n1537) );
    nand2i_5 U997 ( .x(n685), .a(n3604), .b(n3598) );
    aoi21_1 U998 ( .x(n2628), .a(n1177), .b(n2629), .c(n2630) );
    nand2i_2 U999 ( .x(n3836), .a(n4004), .b(n2981) );
    EX_DW01_add_32_5_test_1 add_271 ( .A({reg_out_A[31], reg_out_A[30], 
        reg_out_A[29], reg_out_A[28], n537, reg_out_A[26], n590, reg_out_A[24], 
        n634, n686, reg_out_A[21], n749, reg_out_A[19], reg_out_A[18], 
        reg_out_A[17], reg_out_A[16], n4016, n934, n930, reg_out_A[12], 
        reg_out_A[11], reg_out_A[10], reg_out_A[9], reg_out_A[8], reg_out_A[7], 
        n922, reg_out_A[5], reg_out_A[4], reg_out_A[3], n940, n832, n942}), 
        .B({Imm[31], Imm[30], Imm[29], Imm[28], n681, Imm[26], n689, Imm[24], 
        n829, n745, Imm[21], Imm[20], n684, Imm[18], Imm[17], Imm[16], Imm[15], 
        Imm[14], Imm[13], n682, n753, Imm[10], Imm[9], Imm[8], Imm[7], Imm[6], 
        Imm[5], Imm[4], Imm[3], Imm[2], net149122, Imm[0]}), .CI(1'b0), .SUM({
        N1729, N1728, N1727, N1726, N1725, N1724, N1723, N1722, N1721, N1720, 
        N1719, N1718, N1717, N1716, N1715, N1714, N1713, N1712, N1711, N1710, 
        N1709, N1708, N1707, N1706, N1705, N1704, N1703, N1702, N1701, N1700, 
        N1699, N1698}) );
    EX_DW01_add_32_6_test_1 add_277 ( .A({reg_out_A[31], reg_out_A[30], n539, 
        reg_out_A[28], n533, reg_out_A[26], n590, reg_out_A[24], n634, n583, 
        reg_out_A[21], n749, reg_out_A[19], reg_out_A[18], reg_out_A[17], 
        reg_out_A[16], n4014, n934, n930, reg_out_A[12], reg_out_A[11], 
        reg_out_A[10], reg_out_A[9], reg_out_A[8], reg_out_A[7], n921, 
        reg_out_A[5], reg_out_A[4], reg_out_A[3], n939, n832, n943}), .B({
        Imm[31], Imm[30], Imm[29], Imm[28], n681, Imm[26], n689, Imm[24], n831, 
        n745, Imm[21], Imm[20], Imm[19], Imm[18], Imm[17], Imm[16], Imm[15], 
        Imm[14], Imm[13], Imm[12], Imm[11], Imm[10], Imm[9], Imm[8], Imm[7], 
        Imm[6], Imm[5], Imm[4], Imm[3], Imm[2], net149121, Imm[0]}), .CI(1'b0), 
        .SUM({N1762, N1761, N1760, N1759, N1758, N1757, N1756, N1755, N1754, 
        N1753, N1752, N1751, N1750, N1749, N1748, N1747, N1746, N1745, N1744, 
        N1743, N1742, N1741, N1740, N1739, N1738, N1737, N1736, N1735, N1734, 
        N1733, N1732, N1731}) );
    EX_DW01_add_32_4_test_1 add_289 ( .A({reg_out_A[31], reg_out_A[30], 
        reg_out_A[29], reg_out_A[28], n537, reg_out_A[26], n590, reg_out_A[24], 
        n636, n583, reg_out_A[21], reg_out_A[20], reg_out_A[19], reg_out_A[18], 
        reg_out_A[17], reg_out_A[16], n608, n934, n930, reg_out_A[12], 
        reg_out_A[11], reg_out_A[10], reg_out_A[9], reg_out_A[8], reg_out_A[7], 
        n922, reg_out_A[5], reg_out_A[4], reg_out_A[3], n940, n832, n943}), 
        .B({Imm[31], Imm[30], Imm[29], Imm[28], n681, Imm[26], n689, Imm[24], 
        n831, n745, Imm[21], Imm[20], Imm[19], Imm[18], Imm[17], Imm[16], 
        Imm[15], Imm[14], Imm[13], Imm[12], Imm[11], Imm[10], Imm[9], Imm[8], 
        Imm[7], Imm[6], Imm[5], Imm[4], Imm[3], Imm[2], net149121, Imm[0]}), 
        .CI(1'b0), .SUM({N1828, N1827, N1826, N1825, N1824, N1823, N1822, 
        N1821, N1820, N1819, N1818, N1817, N1816, N1815, N1814, N1813, N1812, 
        N1811, N1810, N1809, N1808, N1807, N1806, N1805, N1804, N1803, N1802, 
        N1801, N1800, N1799, N1798, N1797}) );
    EX_DW01_add_32_3_test_1 add_295 ( .A({reg_out_A[31], n535, n539, n538, 
        n533, reg_out_A[26], n590, reg_out_A[24], n636, n687, reg_out_A[21], 
        reg_out_A[20], reg_out_A[19], reg_out_A[18], n863, reg_out_A[16], 
        n4014, n933, n930, reg_out_A[12], reg_out_A[11], reg_out_A[10], 
        reg_out_A[9], reg_out_A[8], reg_out_A[7], n936, reg_out_A[5], 
        reg_out_A[4], reg_out_A[3], n940, n603, n942}), .B({Imm[31], Imm[30], 
        Imm[29], Imm[28], n681, Imm[26], n689, Imm[24], n831, n745, Imm[21], 
        Imm[20], Imm[19], Imm[18], Imm[17], Imm[16], Imm[15], Imm[14], Imm[13], 
        Imm[12], Imm[11], Imm[10], Imm[9], Imm[8], Imm[7], Imm[6], Imm[5], 
        Imm[4], Imm[3], Imm[2], net149106, Imm[0]}), .CI(1'b0), .SUM({N1861, 
        N1860, N1859, N1858, N1857, N1856, N1855, N1854, N1853, N1852, N1851, 
        N1850, N1849, N1848, N1847, N1846, N1845, N1844, N1843, N1842, N1841, 
        N1840, N1839, N1838, N1837, N1836, N1835, N1834, N1833, N1832, N1831, 
        N1830}) );
    EX_DW01_add_32_7_test_1 add_301 ( .A({reg_out_A[31], reg_out_A[30], n539, 
        n538, n533, n540, n590, reg_out_A[24], n636, n686, reg_out_A[21], n749, 
        reg_out_A[19], reg_out_A[18], reg_out_A[17], reg_out_A[16], n602, n933, 
        n930, reg_out_A[12], reg_out_A[11], reg_out_A[10], reg_out_A[9], 
        reg_out_A[8], reg_out_A[7], n838, reg_out_A[5], reg_out_A[4], 
        reg_out_A[3], n692, n603, n942}), .B({Imm[31], Imm[30], Imm[29], 
        Imm[28], n681, Imm[26], n689, Imm[24], n829, n745, Imm[21], n551, 
        Imm[19], Imm[18], Imm[17], Imm[16], Imm[15], Imm[14], Imm[13], Imm[12], 
        Imm[11], Imm[10], Imm[9], Imm[8], Imm[7], Imm[6], Imm[5], Imm[4], 
        Imm[3], n637, net149120, Imm[0]}), .CI(1'b0), .SUM({N1894, N1893, 
        N1892, N1891, N1890, N1889, N1888, N1887, N1886, N1885, N1884, N1883, 
        N1882, N1881, N1880, N1879, N1878, N1877, N1876, N1875, N1874, N1873, 
        N1872, N1871, N1870, N1869, N1868, N1867, N1866, N1865, N1864, N1863})
         );
    EX_DW01_add_32_1_test_1 add_310 ( .A({reg_out_A[31], reg_out_A[30], 
        reg_out_A[29], n538, n537, n540, n590, n541, n634, n686, n628, n749, 
        n887, n910, n902, n893, n609, n934, n930, n894, reg_out_A[11], n908, 
        n904, reg_out_A[8], reg_out_A[7], n921, n912, n834, n885, n940, n832, 
        n943}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, net151622, net156363, n556, n682, 
        n753, Imm[10], net149617, Imm[8], Imm[7], Imm[6], net151578, net151904, 
        net149167, n637, net149122, Imm[0]}), .CI(1'b0), .SUM({N1961, N1960, 
        N1959, N1958, N1957, N1956, N1955, N1954, N1953, N1952, N1951, N1950, 
        N1949, N1948, N1947, N1946, N1945, N1944, N1943, N1942, N1941, N1940, 
        N1939, N1938, N1937, N1936, N1935, N1934, N1933, N1932, N1931, N1930})
         );
    smlatnr_1 byte_reg__master ( .q(byte_reg__m2s), .d(n4048), .sdi(ALU_result
        [31]), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n542), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 byte_reg__slave ( .q(_byte), .qb(n4046), .d(byte_reg__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n542), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    EX_DW01_cmp2_32_3_test_1 gte_246 ( .A({N70, reg_out_B[30], reg_out_B[29], 
        reg_out_B[28], reg_out_B[27], reg_out_B[26], reg_out_B[25], 
        reg_out_B[24], reg_out_B[23], reg_out_B[22], n566, reg_out_B[20], 
        reg_out_B[19], reg_out_B[18], reg_out_B[17], reg_out_B[16], 
        reg_out_B[15], reg_out_B[14], reg_out_B[13], reg_out_B[12], 
        reg_out_B[11], reg_out_B[10], reg_out_B[9], reg_out_B[8], n4146, 
        reg_out_B[6], reg_out_B[5], reg_out_B[4], reg_out_B[3], n815, n816, 
        reg_out_B[0]}), .B({N69, reg_out_A[30], reg_out_A[29], reg_out_A[28], 
        n533, reg_out_A[26], reg_out_A[25], reg_out_A[24], n634, n583, 
        reg_out_A[21], n749, n887, n910, n902, n893, n4016, n644, n930, n894, 
        n901, n908, n904, n914, n852, n838, n912, n834, reg_out_A[3], n692, 
        n917, n942}), .LEQ(1'b1), .TC(1'b0), .LT_LE(N1407) );
    EX_DW01_cmp2_32_0 gte_348 ( .A({N144, Imm[30], Imm[29], Imm[28], n681, 
        Imm[26], n689, Imm[24], n829, n745, Imm[21], n551, n684, n633, n640, 
        n631, net151622, net156363, n556, n682, n753, Imm[10], net149617, 
        net149628, Imm[7], n642, net151578, net151904, n527, n891, n694, 
        net152465}), .B({N69, reg_out_A[30], reg_out_A[29], reg_out_A[28], 
        n533, reg_out_A[26], n590, n541, n636, n583, reg_out_A[21], n749, n887, 
        n910, n902, n893, n608, n644, n930, n894, n901, n908, n904, n914, n852, 
        n838, n912, n834, n885, n692, n917, n942}), .LEQ(1'b1), .TC(1'b0), 
        .LT_LE(N3029) );
    EX_DW01_cmp2_32_5_test_1 lt_240 ( .A({N69, reg_out_A[30], reg_out_A[29], 
        reg_out_A[28], n533, reg_out_A[26], reg_out_A[25], reg_out_A[24], n634, 
        n686, n628, n749, n887, n910, n902, n893, n609, n644, n919, n894, n901, 
        n908, n904, n914, n852, n838, n912, n834, reg_out_A[3], n692, n917, 
        n943}), .B({N70, reg_out_B[30], reg_out_B[29], reg_out_B[28], 
        reg_out_B[27], reg_out_B[26], reg_out_B[25], reg_out_B[24], 
        reg_out_B[23], reg_out_B[22], n566, reg_out_B[20], reg_out_B[19], 
        reg_out_B[18], reg_out_B[17], reg_out_B[16], reg_out_B[15], 
        reg_out_B[14], reg_out_B[13], reg_out_B[12], reg_out_B[11], 
        reg_out_B[10], reg_out_B[9], reg_out_B[8], n4146, reg_out_B[6], 
        reg_out_B[5], reg_out_B[4], reg_out_B[3], n815, n816, reg_out_B[0]}), 
        .LEQ(1'b0), .TC(1'b0), .LT_LE(N1392) );
    EX_DW01_cmp2_32_2 lt_342 ( .A({N69, reg_out_A[30], reg_out_A[29], 
        reg_out_A[28], n533, reg_out_A[26], reg_out_A[25], reg_out_A[24], n635, 
        n583, reg_out_A[21], n749, n887, n910, n902, n893, n602, n644, n919, 
        n894, n901, n908, n904, n914, reg_out_A[7], n920, n912, n834, 
        reg_out_A[3], n692, n917, n943}), .B({N144, Imm[30], Imm[29], Imm[28], 
        n681, Imm[26], n689, Imm[24], n831, n745, Imm[21], n551, n684, n633, 
        n640, n631, net151622, net156363, n629, n682, n753, n818, net149617, 
        net149628, Imm[7], Imm[6], net151578, net151904, Imm[3], n891, 
        net149120, net152465}), .LEQ(1'b0), .TC(1'b0), .LT_LE(N3014) );
    EX_DW01_cmp2_32_4_test_1 lte_242 ( .A({N69, reg_out_A[30], reg_out_A[29], 
        reg_out_A[28], n533, reg_out_A[26], reg_out_A[25], reg_out_A[24], n636, 
        n686, reg_out_A[21], n749, n596, n910, n902, n893, n609, n644, n524, 
        n894, n901, n908, n904, n914, n852, n922, n912, n834, reg_out_A[3], 
        n692, n917, n943}), .B({N70, reg_out_B[30], reg_out_B[29], 
        reg_out_B[28], reg_out_B[27], reg_out_B[26], reg_out_B[25], 
        reg_out_B[24], reg_out_B[23], reg_out_B[22], n566, reg_out_B[20], 
        reg_out_B[19], reg_out_B[18], reg_out_B[17], reg_out_B[16], 
        reg_out_B[15], reg_out_B[14], reg_out_B[13], reg_out_B[12], 
        reg_out_B[11], reg_out_B[10], reg_out_B[9], reg_out_B[8], n4146, 
        reg_out_B[6], reg_out_B[5], reg_out_B[4], reg_out_B[3], n815, n816, 
        reg_out_B[0]}), .LEQ(1'b1), .TC(1'b0), .LT_LE(N1402) );
    EX_DW01_cmp2_32_1 lte_344 ( .A({N69, reg_out_A[30], reg_out_A[29], 
        reg_out_A[28], n533, reg_out_A[26], reg_out_A[25], reg_out_A[24], n634, 
        n686, n628, n749, n887, n910, n902, n893, n609, n644, n524, n894, n901, 
        n908, n904, n914, n852, n922, n912, n834, n885, n692, n917, n943}), 
        .B({N144, Imm[30], Imm[29], Imm[28], n681, Imm[26], n689, Imm[24], 
        n829, n745, Imm[21], n551, n684, n633, n639, n631, net151622, Imm[14], 
        Imm[13], Imm[12], n753, n818, net149617, net149628, Imm[7], n642, 
        net151578, net151904, Imm[3], n891, net149120, net152465}), .LEQ(1'b1), 
        .TC(1'b0), .LT_LE(N3024) );
    smlatnr_1 mem_read_EX_reg__master ( .q(mem_read_EX_reg__m2s), .d(n4202), 
        .sdi(_byte), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n542), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_1 mem_read_EX_reg__slave ( .q(mem_read_EX), .d(mem_read_EX_reg__m2s
        ), .g(Ctrl__Regs_1__en2), .rb(n542), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 mem_to_reg_EX_reg__master ( .q(mem_to_reg_EX_reg__m2s), .d(n4200
        ), .sdi(mem_read_EX), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n543), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_4 mem_to_reg_EX_reg__slave ( .q(n4224), .qb(n4201), .d(
        mem_to_reg_EX_reg__m2s), .g(Ctrl__Regs_1__en2), .rb(n543), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 mem_write_EX_reg__master ( .q(mem_write_EX_reg__m2s), .d(n4203), 
        .sdi(n4201), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n543), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_1 mem_write_EX_reg__slave ( .q(mem_write_EX), .d(
        mem_write_EX_reg__m2s), .g(Ctrl__Regs_1__en2), .rb(n543), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    EX_DW01_sub_32_2_test_1 r1860_0 ( .A({reg_out_A[31], reg_out_A[30], n539, 
        n538, n537, n540, n590, n541, n634, n583, n628, reg_out_A[20], 
        reg_out_A[19], reg_out_A[18], n586, n893, n608, n934, n918, 
        reg_out_A[12], reg_out_A[11], n908, reg_out_A[9], reg_out_A[8], 
        reg_out_A[7], n838, reg_out_A[5], reg_out_A[4], reg_out_A[3], n939, 
        n832, n943}), .B({n4144, reg_out_B[30], reg_out_B[29], reg_out_B[28], 
        reg_out_B[27], reg_out_B[26], reg_out_B[25], reg_out_B[24], 
        reg_out_B[23], reg_out_B[22], n567, reg_out_B[20], reg_out_B[19], 
        reg_out_B[18], reg_out_B[17], reg_out_B[16], reg_out_B[15], 
        reg_out_B[14], reg_out_B[13], reg_out_B[12], reg_out_B[11], 
        reg_out_B[10], reg_out_B[9], reg_out_B[8], n4146, reg_out_B[6], 
        reg_out_B[5], reg_out_B[4], reg_out_B[3], reg_out_B[2], reg_out_B[1], 
        reg_out_B[0]}), .CI(1'b0), .DIFF({N371, N370, N369, N368, N367, N366, 
        N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, 
        N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, 
        N341, N340}) );
    EX_DW01_add_32_2_test_1 r1865_0 ( .A({reg_out_A[31], reg_out_A[30], n539, 
        reg_out_A[28], reg_out_A[27], reg_out_A[26], reg_out_A[25], 
        reg_out_A[24], n634, n687, reg_out_A[21], n749, reg_out_A[19], 
        reg_out_A[18], reg_out_A[17], reg_out_A[16], n4016, n934, n918, 
        reg_out_A[12], reg_out_A[11], reg_out_A[10], reg_out_A[9], 
        reg_out_A[8], reg_out_A[7], n921, reg_out_A[5], reg_out_A[4], 
        reg_out_A[3], n939, n832, n943}), .B({Imm[31], Imm[30], Imm[29], 
        Imm[28], n681, Imm[26], n689, Imm[24], n829, n745, Imm[21], n551, 
        Imm[19], Imm[18], Imm[17], Imm[16], Imm[15], Imm[14], Imm[13], Imm[12], 
        Imm[11], Imm[10], Imm[9], Imm[8], Imm[7], Imm[6], Imm[5], Imm[4], 
        Imm[3], Imm[2], net149106, Imm[0]}), .CI(1'b0), .SUM({N1663, N1662, 
        N1661, N1660, N1659, N1658, N1657, N1656, N1655, N1654, N1653, N1652, 
        N1651, N1650, N1649, N1648, N1647, N1646, N1645, N1644, N1643, N1642, 
        N1641, N1640, N1639, N1638, N1637, N1636, N1635, N1634, N1633, N1632})
         );
    EX_DW01_add_32_0_test_1 r247_0 ( .A({reg_out_A[31], n535, reg_out_A[29], 
        reg_out_A[28], n533, reg_out_A[26], reg_out_A[25], reg_out_A[24], n634, 
        n583, reg_out_A[21], reg_out_A[20], reg_out_A[19], reg_out_A[18], 
        reg_out_A[17], reg_out_A[16], n608, n644, n930, n894, n901, n908, n904, 
        n914, reg_out_A[7], n922, reg_out_A[5], reg_out_A[4], reg_out_A[3], 
        n940, n832, n942}), .B({n4144, reg_out_B[30], reg_out_B[29], 
        reg_out_B[28], reg_out_B[27], reg_out_B[26], reg_out_B[25], 
        reg_out_B[24], reg_out_B[23], reg_out_B[22], n567, reg_out_B[20], 
        reg_out_B[19], reg_out_B[18], reg_out_B[17], reg_out_B[16], 
        reg_out_B[15], reg_out_B[14], reg_out_B[13], reg_out_B[12], 
        reg_out_B[11], reg_out_B[10], reg_out_B[9], reg_out_B[8], n4146, 
        reg_out_B[6], reg_out_B[5], reg_out_B[4], reg_out_B[3], reg_out_B[2], 
        reg_out_B[1], reg_out_B[0]}), .CI(1'b0), .SUM({N338, N337, N336, N335, 
        N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, 
        N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, 
        N310, N309, N308, N307}) );
    smlatnr_1 reg_out_B_EX_reg_0__master ( .q(reg_out_B_EX_reg_0__m2s), .d(
        n4212), .sdi(mem_write_EX), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(
        n4017), .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_1 reg_out_B_EX_reg_0__slave ( .q(reg_out_B_EX[0]), .qb(n4213), .d(
        reg_out_B_EX_reg_0__m2s), .g(Ctrl__Regs_1__en2), .rb(n4017), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_EX_reg_10__master ( .q(reg_out_B_EX_reg_10__m2s), .d(
        n4182), .sdi(n4209), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n543), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_1 reg_out_B_EX_reg_10__slave ( .q(reg_out_B_EX[10]), .qb(n4183), 
        .d(reg_out_B_EX_reg_10__m2s), .g(Ctrl__Regs_1__en2), .rb(n543), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_EX_reg_11__master ( .q(reg_out_B_EX_reg_11__m2s), .d(
        n4214), .sdi(n4183), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4017), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_1 reg_out_B_EX_reg_11__slave ( .q(reg_out_B_EX[11]), .qb(n4215), 
        .d(reg_out_B_EX_reg_11__m2s), .g(Ctrl__Regs_1__en2), .rb(n4017), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_EX_reg_12__master ( .q(reg_out_B_EX_reg_12__m2s), .d(
        n4180), .sdi(n4215), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4017), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_1 reg_out_B_EX_reg_12__slave ( .q(reg_out_B_EX[12]), .qb(n4181), 
        .d(reg_out_B_EX_reg_12__m2s), .g(Ctrl__Regs_1__en2), .rb(n4017), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_EX_reg_13__master ( .q(reg_out_B_EX_reg_13__m2s), .d(
        n4216), .sdi(n4181), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n543), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_1 reg_out_B_EX_reg_13__slave ( .q(reg_out_B_EX[13]), .qb(n4217), 
        .d(reg_out_B_EX_reg_13__m2s), .g(Ctrl__Regs_1__en2), .rb(n543), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_EX_reg_14__master ( .q(reg_out_B_EX_reg_14__m2s), .d(
        n4178), .sdi(n4217), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4017), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_1 reg_out_B_EX_reg_14__slave ( .q(reg_out_B_EX[14]), .qb(n4179), 
        .d(reg_out_B_EX_reg_14__m2s), .g(Ctrl__Regs_1__en2), .rb(n4017), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_EX_reg_15__master ( .q(reg_out_B_EX_reg_15__m2s), .d(
        n4158), .sdi(n4179), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4017), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_1 reg_out_B_EX_reg_15__slave ( .q(reg_out_B_EX[15]), .qb(n4159), 
        .d(reg_out_B_EX_reg_15__m2s), .g(Ctrl__Regs_1__en2), .rb(n4017), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_EX_reg_16__master ( .q(reg_out_B_EX_reg_16__m2s), .d(
        n4176), .sdi(n4159), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4017), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_1 reg_out_B_EX_reg_16__slave ( .q(reg_out_B_EX[16]), .qb(n4177), 
        .d(reg_out_B_EX_reg_16__m2s), .g(Ctrl__Regs_1__en2), .rb(n4017), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_EX_reg_17__master ( .q(reg_out_B_EX_reg_17__m2s), .d(
        n4222), .sdi(n4177), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n543), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_1 reg_out_B_EX_reg_17__slave ( .q(reg_out_B_EX[17]), .qb(n4223), 
        .d(reg_out_B_EX_reg_17__m2s), .g(Ctrl__Regs_1__en2), .rb(n543), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_EX_reg_18__master ( .q(reg_out_B_EX_reg_18__m2s), .d(
        n4210), .sdi(n4223), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n542), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_1 reg_out_B_EX_reg_18__slave ( .q(reg_out_B_EX[18]), .qb(n4211), 
        .d(reg_out_B_EX_reg_18__m2s), .g(Ctrl__Regs_1__en2), .rb(n542), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_EX_reg_19__master ( .q(reg_out_B_EX_reg_19__m2s), .d(
        n4174), .sdi(n4211), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n543), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_1 reg_out_B_EX_reg_19__slave ( .q(reg_out_B_EX[19]), .qb(n4175), 
        .d(reg_out_B_EX_reg_19__m2s), .g(Ctrl__Regs_1__en2), .rb(n543), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_EX_reg_1__master ( .q(reg_out_B_EX_reg_1__m2s), .d(
        n4160), .sdi(n4213), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n542), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_1 reg_out_B_EX_reg_1__slave ( .q(reg_out_B_EX[1]), .qb(n4161), .d(
        reg_out_B_EX_reg_1__m2s), .g(Ctrl__Regs_1__en2), .rb(n542), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_EX_reg_20__master ( .q(reg_out_B_EX_reg_20__m2s), .d(
        n4218), .sdi(n4175), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n543), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_1 reg_out_B_EX_reg_20__slave ( .q(reg_out_B_EX[20]), .qb(n4219), 
        .d(reg_out_B_EX_reg_20__m2s), .g(Ctrl__Regs_1__en2), .rb(n543), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_EX_reg_21__master ( .q(reg_out_B_EX_reg_21__m2s), .d(
        n4162), .sdi(n4219), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n542), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_1 reg_out_B_EX_reg_21__slave ( .q(reg_out_B_EX[21]), .qb(n4163), 
        .d(reg_out_B_EX_reg_21__m2s), .g(Ctrl__Regs_1__en2), .rb(n542), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_EX_reg_22__master ( .q(reg_out_B_EX_reg_22__m2s), .d(
        n4204), .sdi(n4163), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n542), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_1 reg_out_B_EX_reg_22__slave ( .q(reg_out_B_EX[22]), .qb(n4205), 
        .d(reg_out_B_EX_reg_22__m2s), .g(Ctrl__Regs_1__en2), .rb(n542), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_EX_reg_23__master ( .q(reg_out_B_EX_reg_23__m2s), .d(
        n4172), .sdi(n4205), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n543), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_1 reg_out_B_EX_reg_23__slave ( .q(reg_out_B_EX[23]), .qb(n4173), 
        .d(reg_out_B_EX_reg_23__m2s), .g(Ctrl__Regs_1__en2), .rb(n543), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_EX_reg_24__master ( .q(reg_out_B_EX_reg_24__m2s), .d(
        n4156), .sdi(n4173), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4017), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_1 reg_out_B_EX_reg_24__slave ( .q(reg_out_B_EX[24]), .qb(n4157), 
        .d(reg_out_B_EX_reg_24__m2s), .g(Ctrl__Regs_1__en2), .rb(n4017), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_EX_reg_25__master ( .q(reg_out_B_EX_reg_25__m2s), .d(
        n4170), .sdi(n4157), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4017), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_1 reg_out_B_EX_reg_25__slave ( .q(reg_out_B_EX[25]), .qb(n4171), 
        .d(reg_out_B_EX_reg_25__m2s), .g(Ctrl__Regs_1__en2), .rb(n4017), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_EX_reg_26__master ( .q(reg_out_B_EX_reg_26__m2s), .d(
        n4206), .sdi(n4171), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n542), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_1 reg_out_B_EX_reg_26__slave ( .q(reg_out_B_EX[26]), .qb(n4207), 
        .d(reg_out_B_EX_reg_26__m2s), .g(Ctrl__Regs_1__en2), .rb(n542), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_EX_reg_27__master ( .q(reg_out_B_EX_reg_27__m2s), .d(
        n4168), .sdi(n4207), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n542), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_1 reg_out_B_EX_reg_27__slave ( .q(reg_out_B_EX[27]), .qb(n4169), 
        .d(reg_out_B_EX_reg_27__m2s), .g(Ctrl__Regs_1__en2), .rb(n542), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_EX_reg_28__master ( .q(reg_out_B_EX_reg_28__m2s), .d(
        n4166), .sdi(n4169), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n542), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_1 reg_out_B_EX_reg_28__slave ( .q(reg_out_B_EX[28]), .qb(n4167), 
        .d(reg_out_B_EX_reg_28__m2s), .g(Ctrl__Regs_1__en2), .rb(n542), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_EX_reg_29__master ( .q(reg_out_B_EX_reg_29__m2s), .d(
        n4220), .sdi(n4167), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n542), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_1 reg_out_B_EX_reg_29__slave ( .q(reg_out_B_EX[29]), .qb(n4221), 
        .d(reg_out_B_EX_reg_29__m2s), .g(Ctrl__Regs_1__en2), .rb(n542), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_EX_reg_2__master ( .q(reg_out_B_EX_reg_2__m2s), .d(
        n4196), .sdi(n4161), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n543), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_1 reg_out_B_EX_reg_2__slave ( .q(reg_out_B_EX[2]), .qb(n4197), .d(
        reg_out_B_EX_reg_2__m2s), .g(Ctrl__Regs_1__en2), .rb(n543), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_EX_reg_30__master ( .q(reg_out_B_EX_reg_30__m2s), .d(
        n4164), .sdi(n4221), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n542), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_1 reg_out_B_EX_reg_30__slave ( .q(reg_out_B_EX[30]), .qb(n4165), 
        .d(reg_out_B_EX_reg_30__m2s), .g(Ctrl__Regs_1__en2), .rb(n542), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_EX_reg_31__master ( .q(reg_out_B_EX_reg_31__m2s), .d(
        N3297), .sdi(n4165), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4017), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 reg_out_B_EX_reg_31__slave ( .q(reg_out_B_EX[31]), .qb(n4150), 
        .d(reg_out_B_EX_reg_31__m2s), .g(Ctrl__Regs_1__en2), .rb(n4017), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_EX_reg_3__master ( .q(reg_out_B_EX_reg_3__m2s), .d(
        n4194), .sdi(n4197), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n542), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_1 reg_out_B_EX_reg_3__slave ( .q(reg_out_B_EX[3]), .qb(n4195), .d(
        reg_out_B_EX_reg_3__m2s), .g(Ctrl__Regs_1__en2), .rb(n542), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_EX_reg_4__master ( .q(reg_out_B_EX_reg_4__m2s), .d(
        n4192), .sdi(n4195), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n542), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_1 reg_out_B_EX_reg_4__slave ( .q(reg_out_B_EX[4]), .qb(n4193), .d(
        reg_out_B_EX_reg_4__m2s), .g(Ctrl__Regs_1__en2), .rb(n542), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_EX_reg_5__master ( .q(reg_out_B_EX_reg_5__m2s), .d(
        n4190), .sdi(n4193), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n543), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_1 reg_out_B_EX_reg_5__slave ( .q(reg_out_B_EX[5]), .qb(n4191), .d(
        reg_out_B_EX_reg_5__m2s), .g(Ctrl__Regs_1__en2), .rb(n543), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_EX_reg_6__master ( .q(reg_out_B_EX_reg_6__m2s), .d(
        n4188), .sdi(n4191), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4017), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_1 reg_out_B_EX_reg_6__slave ( .q(reg_out_B_EX[6]), .qb(n4189), .d(
        reg_out_B_EX_reg_6__m2s), .g(Ctrl__Regs_1__en2), .rb(n4017), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_EX_reg_7__master ( .q(reg_out_B_EX_reg_7__m2s), .d(
        n4186), .sdi(n4189), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4017), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_1 reg_out_B_EX_reg_7__slave ( .q(reg_out_B_EX[7]), .qb(n4187), .d(
        reg_out_B_EX_reg_7__m2s), .g(Ctrl__Regs_1__en2), .rb(n4017), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_EX_reg_8__master ( .q(reg_out_B_EX_reg_8__m2s), .d(
        n4184), .sdi(n4187), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n543), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_1 reg_out_B_EX_reg_8__slave ( .q(reg_out_B_EX[8]), .qb(n4185), .d(
        reg_out_B_EX_reg_8__m2s), .g(Ctrl__Regs_1__en2), .rb(n543), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_EX_reg_9__master ( .q(reg_out_B_EX_reg_9__m2s), .d(
        n4208), .sdi(n4185), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n543), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_1 reg_out_B_EX_reg_9__slave ( .q(reg_out_B_EX[9]), .qb(n4209), .d(
        reg_out_B_EX_reg_9__m2s), .g(Ctrl__Regs_1__en2), .rb(n543), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_write_EX_reg__master ( .q(reg_write_EX_reg__m2s), .d(n4198), 
        .sdi(n4150), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4017), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_1 reg_write_EX_reg__slave ( .q(reg_write_EX), .qb(n4199), .d(
        reg_write_EX_reg__m2s), .g(Ctrl__Regs_1__en2), .rb(n4017), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    EX_DW01_sub_32_0_test_1 sub_312 ( .A({reg_out_A[31], reg_out_A[30], 
        reg_out_A[29], reg_out_A[28], n533, reg_out_A[26], reg_out_A[25], 
        reg_out_A[24], n636, n686, reg_out_A[21], reg_out_A[20], reg_out_A[19], 
        reg_out_A[18], n902, n893, n602, n934, n930, reg_out_A[12], 
        reg_out_A[11], reg_out_A[10], reg_out_A[9], reg_out_A[8], reg_out_A[7], 
        n922, reg_out_A[5], reg_out_A[4], reg_out_A[3], n940, n917, n943}), 
        .B({Imm[31], Imm[30], Imm[29], Imm[28], n681, Imm[26], n689, Imm[24], 
        n829, n745, Imm[21], Imm[20], n684, Imm[18], n640, n631, net151622, 
        net156363, Imm[13], Imm[12], n753, Imm[10], Imm[9], Imm[8], Imm[7], 
        Imm[6], Imm[5], Imm[4], Imm[3], n637, n694, net152465}), .CI(1'b0), 
        .DIFF({N1994, N1993, N1992, N1991, N1990, N1989, N1988, N1987, N1986, 
        N1985, N1984, N1983, N1982, N1981, N1980, N1979, N1978, N1977, N1976, 
        N1975, N1974, N1973, N1972, N1971, N1970, N1969, N1968, N1967, N1966, 
        N1965, N1964, N1963}) );
    EX_DW01_sub_32_1_test_1 sub_314 ( .A({reg_out_A[31], reg_out_A[30], 
        reg_out_A[29], n538, n533, n540, n590, n541, n636, n583, n628, n749, 
        n887, n910, n902, n893, n608, n934, n930, reg_out_A[12], n901, 
        reg_out_A[10], n904, n914, reg_out_A[7], n921, n912, n834, n885, n692, 
        n917, n943}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, net151622, net156363, 
        Imm[13], Imm[12], n753, Imm[10], net149617, net149628, Imm[7], Imm[6], 
        net151578, net151904, Imm[3], n637, net149120, net152465}), .CI(1'b0), 
        .DIFF({N2027, N2026, N2025, N2024, N2023, N2022, N2021, N2020, N2019, 
        N2018, N2017, N2016, N2015, N2014, N2013, N2012, N2011, N2010, N2009, 
        N2008, N2007, N2006, N2005, N2004, N2003, N2002, N2001, N2000, N1999, 
        N1998, N1997, N1996}) );
    smlatnr_1 word_reg__master ( .q(word_reg__m2s), .d(n4080), .sdi(n4199), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n542), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 word_reg__slave ( .q(test_so), .qb(n4047), .d(word_reg__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n542), .glob_g(global_g2), .sync_sel(sync_sel)
         );
endmodule


module DLX_sync_MUX_OP_32_5_32_2_test_1 ( D0_31, D0_30, D0_29, D0_28, D0_27, 
    D0_26, D0_25, D0_24, D0_23, D0_22, D0_21, D0_20, D0_19, D0_18, D0_17, 
    D0_16, D0_15, D0_14, D0_13, D0_12, D0_11, D0_10, D0_9, D0_8, D0_7, D0_6, 
    D0_5, D0_4, D0_3, D0_2, D0_1, D0_0, D1_31, D1_30, D1_29, D1_28, D1_27, 
    D1_26, D1_25, D1_24, D1_23, D1_22, D1_21, D1_20, D1_19, D1_18, D1_17, 
    D1_16, D1_15, D1_14, D1_13, D1_12, D1_11, D1_10, D1_9, D1_8, D1_7, D1_6, 
    D1_5, D1_4, D1_3, D1_2, D1_1, D1_0, D2_31, D2_30, D2_29, D2_28, D2_27, 
    D2_26, D2_25, D2_24, D2_23, D2_22, D2_21, D2_20, D2_19, D2_18, D2_17, 
    D2_16, D2_15, D2_14, D2_13, D2_12, D2_11, D2_10, D2_9, D2_8, D2_7, D2_6, 
    D2_5, D2_4, D2_3, D2_2, D2_1, D2_0, D3_31, D3_30, D3_29, D3_28, D3_27, 
    D3_26, D3_25, D3_24, D3_23, D3_22, D3_21, D3_20, D3_19, D3_18, D3_17, 
    D3_16, D3_15, D3_14, D3_13, D3_12, D3_11, D3_10, D3_9, D3_8, D3_7, D3_6, 
    D3_5, D3_4, D3_3, D3_2, D3_1, D3_0, D4_31, D4_30, D4_29, D4_28, D4_27, 
    D4_26, D4_25, D4_24, D4_23, D4_22, D4_21, D4_20, D4_19, D4_18, D4_17, 
    D4_16, D4_15, D4_14, D4_13, D4_12, D4_11, D4_10, D4_9, D4_8, D4_7, D4_6, 
    D4_5, D4_4, D4_3, D4_2, D4_1, D4_0, D5_31, D5_30, D5_29, D5_28, D5_27, 
    D5_26, D5_25, D5_24, D5_23, D5_22, D5_21, D5_20, D5_19, D5_18, D5_17, 
    D5_16, D5_15, D5_14, D5_13, D5_12, D5_11, D5_10, D5_9, D5_8, D5_7, D5_6, 
    D5_5, D5_4, D5_3, D5_2, D5_1, D5_0, D6_31, D6_30, D6_29, D6_28, D6_27, 
    D6_26, D6_25, D6_24, D6_23, D6_22, D6_21, D6_20, D6_19, D6_18, D6_17, 
    D6_16, D6_15, D6_14, D6_13, D6_12, D6_11, D6_10, D6_9, D6_8, D6_7, D6_6, 
    D6_5, D6_4, D6_3, D6_2, D6_1, D6_0, D7_31, D7_30, D7_29, D7_28, D7_27, 
    D7_26, D7_25, D7_24, D7_23, D7_22, D7_21, D7_20, D7_19, D7_18, D7_17, 
    D7_16, D7_15, D7_14, D7_13, D7_12, D7_11, D7_10, D7_9, D7_8, D7_7, D7_6, 
    D7_5, D7_4, D7_3, D7_2, D7_1, D7_0, D8_31, D8_30, D8_29, D8_28, D8_27, 
    D8_26, D8_25, D8_24, D8_23, D8_22, D8_21, D8_20, D8_19, D8_18, D8_17, 
    D8_16, D8_15, D8_14, D8_13, D8_12, D8_11, D8_10, D8_9, D8_8, D8_7, D8_6, 
    D8_5, D8_4, D8_3, D8_2, D8_1, D8_0, D9_31, D9_30, D9_29, D9_28, D9_27, 
    D9_26, D9_25, D9_24, D9_23, D9_22, D9_21, D9_20, D9_19, D9_18, D9_17, 
    D9_16, D9_15, D9_14, D9_13, D9_12, D9_11, D9_10, D9_9, D9_8, D9_7, D9_6, 
    D9_5, D9_4, D9_3, D9_2, D9_1, D9_0, D10_31, D10_30, D10_29, D10_28, D10_27, 
    D10_26, D10_25, D10_24, D10_23, D10_22, D10_21, D10_20, D10_19, D10_18, 
    D10_17, D10_16, D10_15, D10_14, D10_13, D10_12, D10_11, D10_10, D10_9, 
    D10_8, D10_7, D10_6, D10_5, D10_4, D10_3, D10_2, D10_1, D10_0, D11_31, 
    D11_30, D11_29, D11_28, D11_27, D11_26, D11_25, D11_24, D11_23, D11_22, 
    D11_21, D11_20, D11_19, D11_18, D11_17, D11_16, D11_15, D11_14, D11_13, 
    D11_12, D11_11, D11_10, D11_9, D11_8, D11_7, D11_6, D11_5, D11_4, D11_3, 
    D11_2, D11_1, D11_0, D12_31, D12_30, D12_29, D12_28, D12_27, D12_26, 
    D12_25, D12_24, D12_23, D12_22, D12_21, D12_20, D12_19, D12_18, D12_17, 
    D12_16, D12_15, D12_14, D12_13, D12_12, D12_11, D12_10, D12_9, D12_8, 
    D12_7, D12_6, D12_5, D12_4, D12_3, D12_2, D12_1, D12_0, D13_31, D13_30, 
    D13_29, D13_28, D13_27, D13_26, D13_25, D13_24, D13_23, D13_22, D13_21, 
    D13_20, D13_19, D13_18, D13_17, D13_16, D13_15, D13_14, D13_13, D13_12, 
    D13_11, D13_10, D13_9, D13_8, D13_7, D13_6, D13_5, D13_4, D13_3, D13_2, 
    D13_1, D13_0, D14_31, D14_30, D14_29, D14_28, D14_27, D14_26, D14_25, 
    D14_24, D14_23, D14_22, D14_21, D14_20, D14_19, D14_18, D14_17, D14_16, 
    D14_15, D14_14, D14_13, D14_12, D14_11, D14_10, D14_9, D14_8, D14_7, D14_6, 
    D14_5, D14_4, D14_3, D14_2, D14_1, D14_0, D15_31, D15_30, D15_29, D15_28, 
    D15_27, D15_26, D15_25, D15_24, D15_23, D15_22, D15_21, D15_20, D15_19, 
    D15_18, D15_17, D15_16, D15_15, D15_14, D15_13, D15_12, D15_11, D15_10, 
    D15_9, D15_8, D15_7, D15_6, D15_5, D15_4, D15_3, D15_2, D15_1, D15_0, 
    D16_31, D16_30, D16_29, D16_28, D16_27, D16_26, D16_25, D16_24, D16_23, 
    D16_22, D16_21, D16_20, D16_19, D16_18, D16_17, D16_16, D16_15, D16_14, 
    D16_13, D16_12, D16_11, D16_10, D16_9, D16_8, D16_7, D16_6, D16_5, D16_4, 
    D16_3, D16_2, D16_1, D16_0, D17_31, D17_30, D17_29, D17_28, D17_27, D17_26, 
    D17_25, D17_24, D17_23, D17_22, D17_21, D17_20, D17_19, D17_18, D17_17, 
    D17_16, D17_15, D17_14, D17_13, D17_12, D17_11, D17_10, D17_9, D17_8, 
    D17_7, D17_6, D17_5, D17_4, D17_3, D17_2, D17_1, D17_0, D18_31, D18_30, 
    D18_29, D18_28, D18_27, D18_26, D18_25, D18_24, D18_23, D18_22, D18_21, 
    D18_20, D18_19, D18_18, D18_17, D18_16, D18_15, D18_14, D18_13, D18_12, 
    D18_11, D18_10, D18_9, D18_8, D18_7, D18_6, D18_5, D18_4, D18_3, D18_2, 
    D18_1, D18_0, D19_31, D19_30, D19_29, D19_28, D19_27, D19_26, D19_25, 
    D19_24, D19_23, D19_22, D19_21, D19_20, D19_19, D19_18, D19_17, D19_16, 
    D19_15, D19_14, D19_13, D19_12, D19_11, D19_10, D19_9, D19_8, D19_7, D19_6, 
    D19_5, D19_4, D19_3, D19_2, D19_1, D19_0, D20_31, D20_30, D20_29, D20_28, 
    D20_27, D20_26, D20_25, D20_24, D20_23, D20_22, D20_21, D20_20, D20_19, 
    D20_18, D20_17, D20_16, D20_15, D20_14, D20_13, D20_12, D20_11, D20_10, 
    D20_9, D20_8, D20_7, D20_6, D20_5, D20_4, D20_3, D20_2, D20_1, D20_0, 
    D21_31, D21_30, D21_29, D21_28, D21_27, D21_26, D21_25, D21_24, D21_23, 
    D21_22, D21_21, D21_20, D21_19, D21_18, D21_17, D21_16, D21_15, D21_14, 
    D21_13, D21_12, D21_11, D21_10, D21_9, D21_8, D21_7, D21_6, D21_5, D21_4, 
    D21_3, D21_2, D21_1, D21_0, D22_31, D22_30, D22_29, D22_28, D22_27, D22_26, 
    D22_25, D22_24, D22_23, D22_22, D22_21, D22_20, D22_19, D22_18, D22_17, 
    D22_16, D22_15, D22_14, D22_13, D22_12, D22_11, D22_10, D22_9, D22_8, 
    D22_7, D22_6, D22_5, D22_4, D22_3, D22_2, D22_1, D22_0, D23_31, D23_30, 
    D23_29, D23_28, D23_27, D23_26, D23_25, D23_24, D23_23, D23_22, D23_21, 
    D23_20, D23_19, D23_18, D23_17, D23_16, D23_15, D23_14, D23_13, D23_12, 
    D23_11, D23_10, D23_9, D23_8, D23_7, D23_6, D23_5, D23_4, D23_3, D23_2, 
    D23_1, D23_0, D24_31, D24_30, D24_29, D24_28, D24_27, D24_26, D24_25, 
    D24_24, D24_23, D24_22, D24_21, D24_20, D24_19, D24_18, D24_17, D24_16, 
    D24_15, D24_14, D24_13, D24_12, D24_11, D24_10, D24_9, D24_8, D24_7, D24_6, 
    D24_5, D24_4, D24_3, D24_2, D24_1, D24_0, D25_31, D25_30, D25_29, D25_28, 
    D25_27, D25_26, D25_25, D25_24, D25_23, D25_22, D25_21, D25_20, D25_19, 
    D25_18, D25_17, D25_16, D25_15, D25_14, D25_13, D25_12, D25_11, D25_10, 
    D25_9, D25_8, D25_7, D25_6, D25_5, D25_4, D25_3, D25_2, D25_1, D25_0, 
    D26_31, D26_30, D26_29, D26_28, D26_27, D26_26, D26_25, D26_24, D26_23, 
    D26_22, D26_21, D26_20, D26_19, D26_18, D26_17, D26_16, D26_15, D26_14, 
    D26_13, D26_12, D26_11, D26_10, D26_9, D26_8, D26_7, D26_6, D26_5, D26_4, 
    D26_3, D26_2, D26_1, D26_0, D27_31, D27_30, D27_29, D27_28, D27_27, D27_26, 
    D27_25, D27_24, D27_23, D27_22, D27_21, D27_20, D27_19, D27_18, D27_17, 
    D27_16, D27_15, D27_14, D27_13, D27_12, D27_11, D27_10, D27_9, D27_8, 
    D27_7, D27_6, D27_5, D27_4, D27_3, D27_2, D27_1, D27_0, D28_31, D28_30, 
    D28_29, D28_28, D28_27, D28_26, D28_25, D28_24, D28_23, D28_22, D28_21, 
    D28_20, D28_19, D28_18, D28_17, D28_16, D28_15, D28_14, D28_13, D28_12, 
    D28_11, D28_10, D28_9, D28_8, D28_7, D28_6, D28_5, D28_4, D28_3, D28_2, 
    D28_1, D28_0, D29_31, D29_30, D29_29, D29_28, D29_27, D29_26, D29_25, 
    D29_24, D29_23, D29_22, D29_21, D29_20, D29_19, D29_18, D29_17, D29_16, 
    D29_15, D29_14, D29_13, D29_12, D29_11, D29_10, D29_9, D29_8, D29_7, D29_6, 
    D29_5, D29_4, D29_3, D29_2, D29_1, D29_0, D30_31, D30_30, D30_29, D30_28, 
    D30_27, D30_26, D30_25, D30_24, D30_23, D30_22, D30_21, D30_20, D30_19, 
    D30_18, D30_17, D30_16, D30_15, D30_14, D30_13, D30_12, D30_11, D30_10, 
    D30_9, D30_8, D30_7, D30_6, D30_5, D30_4, D30_3, D30_2, D30_1, D30_0, 
    D31_31, D31_30, D31_29, D31_28, D31_27, D31_26, D31_25, D31_24, D31_23, 
    D31_22, D31_21, D31_20, D31_19, D31_18, D31_17, D31_16, D31_15, D31_14, 
    D31_13, D31_12, D31_11, D31_10, D31_9, D31_8, D31_7, D31_6, D31_5, D31_4, 
    D31_3, D31_2, D31_1, D31_0, S0, S1, S2, S3, S4, Z_31, Z_30, Z_29, Z_28, 
    Z_27, Z_26, Z_25, Z_24, Z_23, Z_22, Z_21, Z_20, Z_19, Z_18, Z_17, Z_16, 
    Z_15, Z_14, Z_13, Z_12, Z_11, Z_10, Z_9, Z_8, Z_7, Z_6, Z_5, Z_4, Z_3, Z_2, 
    Z_1, Z_0 );
input  D0_31, D0_30, D0_29, D0_28, D0_27, D0_26, D0_25, D0_24, D0_23, D0_22, 
    D0_21, D0_20, D0_19, D0_18, D0_17, D0_16, D0_15, D0_14, D0_13, D0_12, 
    D0_11, D0_10, D0_9, D0_8, D0_7, D0_6, D0_5, D0_4, D0_3, D0_2, D0_1, D0_0, 
    D1_31, D1_30, D1_29, D1_28, D1_27, D1_26, D1_25, D1_24, D1_23, D1_22, 
    D1_21, D1_20, D1_19, D1_18, D1_17, D1_16, D1_15, D1_14, D1_13, D1_12, 
    D1_11, D1_10, D1_9, D1_8, D1_7, D1_6, D1_5, D1_4, D1_3, D1_2, D1_1, D1_0, 
    D2_31, D2_30, D2_29, D2_28, D2_27, D2_26, D2_25, D2_24, D2_23, D2_22, 
    D2_21, D2_20, D2_19, D2_18, D2_17, D2_16, D2_15, D2_14, D2_13, D2_12, 
    D2_11, D2_10, D2_9, D2_8, D2_7, D2_6, D2_5, D2_4, D2_3, D2_2, D2_1, D2_0, 
    D3_31, D3_30, D3_29, D3_28, D3_27, D3_26, D3_25, D3_24, D3_23, D3_22, 
    D3_21, D3_20, D3_19, D3_18, D3_17, D3_16, D3_15, D3_14, D3_13, D3_12, 
    D3_11, D3_10, D3_9, D3_8, D3_7, D3_6, D3_5, D3_4, D3_3, D3_2, D3_1, D3_0, 
    D4_31, D4_30, D4_29, D4_28, D4_27, D4_26, D4_25, D4_24, D4_23, D4_22, 
    D4_21, D4_20, D4_19, D4_18, D4_17, D4_16, D4_15, D4_14, D4_13, D4_12, 
    D4_11, D4_10, D4_9, D4_8, D4_7, D4_6, D4_5, D4_4, D4_3, D4_2, D4_1, D4_0, 
    D5_31, D5_30, D5_29, D5_28, D5_27, D5_26, D5_25, D5_24, D5_23, D5_22, 
    D5_21, D5_20, D5_19, D5_18, D5_17, D5_16, D5_15, D5_14, D5_13, D5_12, 
    D5_11, D5_10, D5_9, D5_8, D5_7, D5_6, D5_5, D5_4, D5_3, D5_2, D5_1, D5_0, 
    D6_31, D6_30, D6_29, D6_28, D6_27, D6_26, D6_25, D6_24, D6_23, D6_22, 
    D6_21, D6_20, D6_19, D6_18, D6_17, D6_16, D6_15, D6_14, D6_13, D6_12, 
    D6_11, D6_10, D6_9, D6_8, D6_7, D6_6, D6_5, D6_4, D6_3, D6_2, D6_1, D6_0, 
    D7_31, D7_30, D7_29, D7_28, D7_27, D7_26, D7_25, D7_24, D7_23, D7_22, 
    D7_21, D7_20, D7_19, D7_18, D7_17, D7_16, D7_15, D7_14, D7_13, D7_12, 
    D7_11, D7_10, D7_9, D7_8, D7_7, D7_6, D7_5, D7_4, D7_3, D7_2, D7_1, D7_0, 
    D8_31, D8_30, D8_29, D8_28, D8_27, D8_26, D8_25, D8_24, D8_23, D8_22, 
    D8_21, D8_20, D8_19, D8_18, D8_17, D8_16, D8_15, D8_14, D8_13, D8_12, 
    D8_11, D8_10, D8_9, D8_8, D8_7, D8_6, D8_5, D8_4, D8_3, D8_2, D8_1, D8_0, 
    D9_31, D9_30, D9_29, D9_28, D9_27, D9_26, D9_25, D9_24, D9_23, D9_22, 
    D9_21, D9_20, D9_19, D9_18, D9_17, D9_16, D9_15, D9_14, D9_13, D9_12, 
    D9_11, D9_10, D9_9, D9_8, D9_7, D9_6, D9_5, D9_4, D9_3, D9_2, D9_1, D9_0, 
    D10_31, D10_30, D10_29, D10_28, D10_27, D10_26, D10_25, D10_24, D10_23, 
    D10_22, D10_21, D10_20, D10_19, D10_18, D10_17, D10_16, D10_15, D10_14, 
    D10_13, D10_12, D10_11, D10_10, D10_9, D10_8, D10_7, D10_6, D10_5, D10_4, 
    D10_3, D10_2, D10_1, D10_0, D11_31, D11_30, D11_29, D11_28, D11_27, D11_26, 
    D11_25, D11_24, D11_23, D11_22, D11_21, D11_20, D11_19, D11_18, D11_17, 
    D11_16, D11_15, D11_14, D11_13, D11_12, D11_11, D11_10, D11_9, D11_8, 
    D11_7, D11_6, D11_5, D11_4, D11_3, D11_2, D11_1, D11_0, D12_31, D12_30, 
    D12_29, D12_28, D12_27, D12_26, D12_25, D12_24, D12_23, D12_22, D12_21, 
    D12_20, D12_19, D12_18, D12_17, D12_16, D12_15, D12_14, D12_13, D12_12, 
    D12_11, D12_10, D12_9, D12_8, D12_7, D12_6, D12_5, D12_4, D12_3, D12_2, 
    D12_1, D12_0, D13_31, D13_30, D13_29, D13_28, D13_27, D13_26, D13_25, 
    D13_24, D13_23, D13_22, D13_21, D13_20, D13_19, D13_18, D13_17, D13_16, 
    D13_15, D13_14, D13_13, D13_12, D13_11, D13_10, D13_9, D13_8, D13_7, D13_6, 
    D13_5, D13_4, D13_3, D13_2, D13_1, D13_0, D14_31, D14_30, D14_29, D14_28, 
    D14_27, D14_26, D14_25, D14_24, D14_23, D14_22, D14_21, D14_20, D14_19, 
    D14_18, D14_17, D14_16, D14_15, D14_14, D14_13, D14_12, D14_11, D14_10, 
    D14_9, D14_8, D14_7, D14_6, D14_5, D14_4, D14_3, D14_2, D14_1, D14_0, 
    D15_31, D15_30, D15_29, D15_28, D15_27, D15_26, D15_25, D15_24, D15_23, 
    D15_22, D15_21, D15_20, D15_19, D15_18, D15_17, D15_16, D15_15, D15_14, 
    D15_13, D15_12, D15_11, D15_10, D15_9, D15_8, D15_7, D15_6, D15_5, D15_4, 
    D15_3, D15_2, D15_1, D15_0, D16_31, D16_30, D16_29, D16_28, D16_27, D16_26, 
    D16_25, D16_24, D16_23, D16_22, D16_21, D16_20, D16_19, D16_18, D16_17, 
    D16_16, D16_15, D16_14, D16_13, D16_12, D16_11, D16_10, D16_9, D16_8, 
    D16_7, D16_6, D16_5, D16_4, D16_3, D16_2, D16_1, D16_0, D17_31, D17_30, 
    D17_29, D17_28, D17_27, D17_26, D17_25, D17_24, D17_23, D17_22, D17_21, 
    D17_20, D17_19, D17_18, D17_17, D17_16, D17_15, D17_14, D17_13, D17_12, 
    D17_11, D17_10, D17_9, D17_8, D17_7, D17_6, D17_5, D17_4, D17_3, D17_2, 
    D17_1, D17_0, D18_31, D18_30, D18_29, D18_28, D18_27, D18_26, D18_25, 
    D18_24, D18_23, D18_22, D18_21, D18_20, D18_19, D18_18, D18_17, D18_16, 
    D18_15, D18_14, D18_13, D18_12, D18_11, D18_10, D18_9, D18_8, D18_7, D18_6, 
    D18_5, D18_4, D18_3, D18_2, D18_1, D18_0, D19_31, D19_30, D19_29, D19_28, 
    D19_27, D19_26, D19_25, D19_24, D19_23, D19_22, D19_21, D19_20, D19_19, 
    D19_18, D19_17, D19_16, D19_15, D19_14, D19_13, D19_12, D19_11, D19_10, 
    D19_9, D19_8, D19_7, D19_6, D19_5, D19_4, D19_3, D19_2, D19_1, D19_0, 
    D20_31, D20_30, D20_29, D20_28, D20_27, D20_26, D20_25, D20_24, D20_23, 
    D20_22, D20_21, D20_20, D20_19, D20_18, D20_17, D20_16, D20_15, D20_14, 
    D20_13, D20_12, D20_11, D20_10, D20_9, D20_8, D20_7, D20_6, D20_5, D20_4, 
    D20_3, D20_2, D20_1, D20_0, D21_31, D21_30, D21_29, D21_28, D21_27, D21_26, 
    D21_25, D21_24, D21_23, D21_22, D21_21, D21_20, D21_19, D21_18, D21_17, 
    D21_16, D21_15, D21_14, D21_13, D21_12, D21_11, D21_10, D21_9, D21_8, 
    D21_7, D21_6, D21_5, D21_4, D21_3, D21_2, D21_1, D21_0, D22_31, D22_30, 
    D22_29, D22_28, D22_27, D22_26, D22_25, D22_24, D22_23, D22_22, D22_21, 
    D22_20, D22_19, D22_18, D22_17, D22_16, D22_15, D22_14, D22_13, D22_12, 
    D22_11, D22_10, D22_9, D22_8, D22_7, D22_6, D22_5, D22_4, D22_3, D22_2, 
    D22_1, D22_0, D23_31, D23_30, D23_29, D23_28, D23_27, D23_26, D23_25, 
    D23_24, D23_23, D23_22, D23_21, D23_20, D23_19, D23_18, D23_17, D23_16, 
    D23_15, D23_14, D23_13, D23_12, D23_11, D23_10, D23_9, D23_8, D23_7, D23_6, 
    D23_5, D23_4, D23_3, D23_2, D23_1, D23_0, D24_31, D24_30, D24_29, D24_28, 
    D24_27, D24_26, D24_25, D24_24, D24_23, D24_22, D24_21, D24_20, D24_19, 
    D24_18, D24_17, D24_16, D24_15, D24_14, D24_13, D24_12, D24_11, D24_10, 
    D24_9, D24_8, D24_7, D24_6, D24_5, D24_4, D24_3, D24_2, D24_1, D24_0, 
    D25_31, D25_30, D25_29, D25_28, D25_27, D25_26, D25_25, D25_24, D25_23, 
    D25_22, D25_21, D25_20, D25_19, D25_18, D25_17, D25_16, D25_15, D25_14, 
    D25_13, D25_12, D25_11, D25_10, D25_9, D25_8, D25_7, D25_6, D25_5, D25_4, 
    D25_3, D25_2, D25_1, D25_0, D26_31, D26_30, D26_29, D26_28, D26_27, D26_26, 
    D26_25, D26_24, D26_23, D26_22, D26_21, D26_20, D26_19, D26_18, D26_17, 
    D26_16, D26_15, D26_14, D26_13, D26_12, D26_11, D26_10, D26_9, D26_8, 
    D26_7, D26_6, D26_5, D26_4, D26_3, D26_2, D26_1, D26_0, D27_31, D27_30, 
    D27_29, D27_28, D27_27, D27_26, D27_25, D27_24, D27_23, D27_22, D27_21, 
    D27_20, D27_19, D27_18, D27_17, D27_16, D27_15, D27_14, D27_13, D27_12, 
    D27_11, D27_10, D27_9, D27_8, D27_7, D27_6, D27_5, D27_4, D27_3, D27_2, 
    D27_1, D27_0, D28_31, D28_30, D28_29, D28_28, D28_27, D28_26, D28_25, 
    D28_24, D28_23, D28_22, D28_21, D28_20, D28_19, D28_18, D28_17, D28_16, 
    D28_15, D28_14, D28_13, D28_12, D28_11, D28_10, D28_9, D28_8, D28_7, D28_6, 
    D28_5, D28_4, D28_3, D28_2, D28_1, D28_0, D29_31, D29_30, D29_29, D29_28, 
    D29_27, D29_26, D29_25, D29_24, D29_23, D29_22, D29_21, D29_20, D29_19, 
    D29_18, D29_17, D29_16, D29_15, D29_14, D29_13, D29_12, D29_11, D29_10, 
    D29_9, D29_8, D29_7, D29_6, D29_5, D29_4, D29_3, D29_2, D29_1, D29_0, 
    D30_31, D30_30, D30_29, D30_28, D30_27, D30_26, D30_25, D30_24, D30_23, 
    D30_22, D30_21, D30_20, D30_19, D30_18, D30_17, D30_16, D30_15, D30_14, 
    D30_13, D30_12, D30_11, D30_10, D30_9, D30_8, D30_7, D30_6, D30_5, D30_4, 
    D30_3, D30_2, D30_1, D30_0, D31_31, D31_30, D31_29, D31_28, D31_27, D31_26, 
    D31_25, D31_24, D31_23, D31_22, D31_21, D31_20, D31_19, D31_18, D31_17, 
    D31_16, D31_15, D31_14, D31_13, D31_12, D31_11, D31_10, D31_9, D31_8, 
    D31_7, D31_6, D31_5, D31_4, D31_3, D31_2, D31_1, D31_0, S0, S1, S2, S3, S4;
output Z_31, Z_30, Z_29, Z_28, Z_27, Z_26, Z_25, Z_24, Z_23, Z_22, Z_21, Z_20, 
    Z_19, Z_18, Z_17, Z_16, Z_15, Z_14, Z_13, Z_12, Z_11, Z_10, Z_9, Z_8, Z_7, 
    Z_6, Z_5, Z_4, Z_3, Z_2, Z_1, Z_0;
    wire n111, n11, n32, n250, n38, n67, n227, n68, n228, n69, n229, n70, n230, 
        n71, n231, n73, n233, n75, n235, n76, n236, n77, n237, n78, n238, n122, 
        n24, n47, n79, n143, n175, n4, n1, n48, n80, n144, n112, n176, n10, 
        n49, n81, n145, n113, n177, n2, n50, n82, n146, n114, n178, n52, n84, 
        n148, n116, n180, n53, n85, n149, n117, n181, n54, n86, n150, n118, 
        n182, n3, n55, n87, n151, n119, n183, n56, n88, n152, n120, n184, n57, 
        n89, n153, n121, n185, n154, n15, n34, n58, n90, n186, n60, n92, n156, 
        n124, n188, n61, n93, n157, n125, n189, n9, n62, n94, n158, n126, n190, 
        n63, n95, n159, n127, n191, n64, n96, n160, n128, n192, n66, n98, n162, 
        n130, n194, n99, n163, n131, n195, n100, n164, n132, n196, n101, n165, 
        n133, n197, n23, n30, n103, n167, n135, n199, n72, n104, n168, n136, 
        n200, n105, n169, n137, n201, n107, n171, n139, n203, n108, n172, n140, 
        n204, n110, n174, n142, n206, n26, n83, n17, n33, n19, n18, n28, n29, 
        n31, n20, n35, n97, n102, n16, n106, n123, n109, n115, n91, n129, n41, 
        n13, n134, n138, n141, n147, n25, n211, n243, n307, n275, n339, n155, 
        n161, n51, n179, n166, n170, n14, n173, n214, n246, n310, n278, n342, 
        n36, n5, n187, n37, n193, n198, n202, n22, n205, n232, n264, n328, 
        n296, n360, n207, n239, n303, n271, n335, n209, n241, n305, n273, n337, 
        n210, n242, n306, n274, n338, n212, n244, n308, n276, n340, n213, n245, 
        n309, n277, n341, n215, n247, n311, n279, n343, n216, n248, n312, n280, 
        n344, n217, n249, n313, n281, n345, n218, n314, n282, n346, n59, n220, 
        n252, n316, n284, n348, n221, n253, n317, n285, n349, n222, n254, n318, 
        n286, n350, n223, n255, n319, n287, n351, n224, n256, n320, n288, n352, 
        n225, n257, n321, n289, n353, n226, n258, n322, n290, n354, n259, n323, 
        n291, n355, n260, n324, n292, n356, n261, n325, n293, n357, n219, n251, 
        n315, n283, n347, n263, n327, n295, n359, n265, n329, n297, n361, n267, 
        n331, n299, n363, n268, n332, n300, n364, n270, n334, n302, n366, n240, 
        n74, n234, n39, n262, n266, n330, n298, n362, n269, n21, n40, n272, 
        n65, n12, n27, n326, n294, n358, n301, n42, n304, n333, n365, n43, n44, 
        n336, n45, n46, n7, n208, n6, n8;
    mux4_2 U1 ( .x(n111), .d0(D4_0), .d1(D12_0), .d2(D20_0), .d3(D28_0), .sl0(
        n11), .sl1(n32) );
    mux4_2 U10 ( .x(n250), .d0(D1_11), .d1(D9_11), .d2(D17_11), .d3(D25_11), 
        .sl0(n11), .sl1(n38) );
    mux2_4 U100 ( .x(Z_20), .d0(n67), .sl(S0), .d1(n227) );
    mux2_4 U101 ( .x(Z_21), .d0(n68), .sl(S0), .d1(n228) );
    mux2_4 U102 ( .x(Z_22), .d0(n69), .sl(S0), .d1(n229) );
    mux2_4 U103 ( .x(Z_23), .d0(n70), .sl(S0), .d1(n230) );
    mux2_4 U104 ( .x(Z_24), .d0(n71), .sl(S0), .d1(n231) );
    mux2_4 U105 ( .x(Z_26), .d0(n73), .sl(S0), .d1(n233) );
    mux2_4 U106 ( .x(Z_28), .d0(n75), .sl(S0), .d1(n235) );
    mux2_4 U107 ( .x(Z_29), .d0(n76), .sl(S0), .d1(n236) );
    mux2_4 U108 ( .x(Z_30), .d0(n77), .sl(S0), .d1(n237) );
    mux2_4 U109 ( .x(Z_31), .d0(n78), .sl(S0), .d1(n238) );
    mux4_2 U11 ( .x(n122), .d0(D4_11), .d1(D12_11), .d2(D20_11), .d3(D28_11), 
        .sl0(n24), .sl1(n32) );
    mux4_3 U110 ( .x(n47), .d0(n79), .d1(n143), .d2(n111), .d3(n175), .sl0(n4), 
        .sl1(n1) );
    mux4_3 U111 ( .x(n48), .d0(n80), .d1(n144), .d2(n112), .d3(n176), .sl0(n10
        ), .sl1(n1) );
    mux4_3 U112 ( .x(n49), .d0(n81), .d1(n145), .d2(n113), .d3(n177), .sl0(n4), 
        .sl1(n2) );
    mux4_3 U113 ( .x(n50), .d0(n82), .d1(n146), .d2(n114), .d3(n178), .sl0(n4), 
        .sl1(n2) );
    mux4_3 U114 ( .x(n52), .d0(n84), .d1(n148), .d2(n116), .d3(n180), .sl0(n4), 
        .sl1(n2) );
    mux4_3 U115 ( .x(n53), .d0(n85), .d1(n149), .d2(n117), .d3(n181), .sl0(n4), 
        .sl1(n2) );
    mux4_3 U116 ( .x(n54), .d0(n86), .d1(n150), .d2(n118), .d3(n182), .sl0(n3), 
        .sl1(n2) );
    mux4_3 U117 ( .x(n55), .d0(n87), .d1(n151), .d2(n119), .d3(n183), .sl0(n3), 
        .sl1(n1) );
    mux4_3 U118 ( .x(n56), .d0(n88), .d1(n152), .d2(n120), .d3(n184), .sl0(n4), 
        .sl1(n2) );
    mux4_3 U119 ( .x(n57), .d0(n89), .d1(n153), .d2(n121), .d3(n185), .sl0(n4), 
        .sl1(n1) );
    mux4_2 U12 ( .x(n154), .d0(D2_11), .d1(D10_11), .d2(D18_11), .d3(D26_11), 
        .sl0(n15), .sl1(n34) );
    mux4_3 U120 ( .x(n58), .d0(n90), .d1(n154), .d2(n122), .d3(n186), .sl0(n3), 
        .sl1(n1) );
    mux4_3 U121 ( .x(n60), .d0(n92), .d1(n156), .d2(n124), .d3(n188), .sl0(n3), 
        .sl1(n2) );
    mux4_3 U122 ( .x(n61), .d0(n93), .d1(n157), .d2(n125), .d3(n189), .sl0(n9), 
        .sl1(n2) );
    mux4_3 U123 ( .x(n62), .d0(n94), .d1(n158), .d2(n126), .d3(n190), .sl0(n4), 
        .sl1(n2) );
    mux4_3 U124 ( .x(n63), .d0(n95), .d1(n159), .d2(n127), .d3(n191), .sl0(n9), 
        .sl1(n2) );
    mux4_3 U125 ( .x(n64), .d0(n96), .d1(n160), .d2(n128), .d3(n192), .sl0(n4), 
        .sl1(n2) );
    mux4_3 U126 ( .x(n66), .d0(n98), .d1(n162), .d2(n130), .d3(n194), .sl0(n9), 
        .sl1(n1) );
    mux4_3 U127 ( .x(n67), .d0(n99), .d1(n163), .d2(n131), .d3(n195), .sl0(n3), 
        .sl1(n2) );
    mux4_3 U128 ( .x(n68), .d0(n100), .d1(n164), .d2(n132), .d3(n196), .sl0(n3
        ), .sl1(n1) );
    mux4_3 U129 ( .x(n69), .d0(n101), .d1(n165), .d2(n133), .d3(n197), .sl0(n9
        ), .sl1(n1) );
    mux4_2 U13 ( .x(n90), .d0(D0_11), .d1(D8_11), .d2(D16_11), .d3(D24_11), 
        .sl0(n23), .sl1(n30) );
    mux4_3 U130 ( .x(n71), .d0(n103), .d1(n167), .d2(n135), .d3(n199), .sl0(n4
        ), .sl1(n1) );
    mux4_3 U131 ( .x(n72), .d0(n104), .d1(n168), .d2(n136), .d3(n200), .sl0(n9
        ), .sl1(n2) );
    mux4_3 U132 ( .x(n73), .d0(n105), .d1(n169), .d2(n137), .d3(n201), .sl0(
        n10), .sl1(n1) );
    mux4_3 U133 ( .x(n75), .d0(n107), .d1(n171), .d2(n139), .d3(n203), .sl0(
        n10), .sl1(n1) );
    mux4_3 U134 ( .x(n76), .d0(n108), .d1(n172), .d2(n140), .d3(n204), .sl0(
        n10), .sl1(n1) );
    mux4_3 U135 ( .x(n78), .d0(n110), .d1(n174), .d2(n142), .d3(n206), .sl0(n9
        ), .sl1(n1) );
    mux4_3 U136 ( .x(n80), .d0(D0_1), .d1(D8_1), .d2(D16_1), .d3(D24_1), .sl0(
        n11), .sl1(n30) );
    mux4_3 U137 ( .x(n81), .d0(D0_2), .d1(D8_2), .d2(D16_2), .d3(D24_2), .sl0(
        n26), .sl1(n30) );
    mux4_3 U138 ( .x(n82), .d0(D0_3), .d1(D8_3), .d2(D16_3), .d3(D24_3), .sl0(
        n26), .sl1(n30) );
    mux4_3 U139 ( .x(n83), .d0(D0_4), .d1(D8_4), .d2(D16_4), .d3(D24_4), .sl0(
        n17), .sl1(n30) );
    mux4_2 U14 ( .x(n136), .d0(D4_25), .d1(D12_25), .d2(D20_25), .d3(D28_25), 
        .sl0(n15), .sl1(n33) );
    mux4_3 U140 ( .x(n84), .d0(D0_5), .d1(D8_5), .d2(D16_5), .d3(D24_5), .sl0(
        n19), .sl1(n30) );
    mux4_3 U141 ( .x(n85), .d0(D0_6), .d1(D8_6), .d2(D16_6), .d3(D24_6), .sl0(
        n23), .sl1(n30) );
    mux4_3 U142 ( .x(n86), .d0(D0_7), .d1(D8_7), .d2(D16_7), .d3(D24_7), .sl0(
        n17), .sl1(n30) );
    mux4_3 U143 ( .x(n88), .d0(D0_9), .d1(D8_9), .d2(D16_9), .d3(D24_9), .sl0(
        n18), .sl1(n30) );
    mux4_3 U144 ( .x(n89), .d0(D0_10), .d1(D8_10), .d2(D16_10), .d3(D24_10), 
        .sl0(n28), .sl1(n30) );
    mux4_3 U145 ( .x(n92), .d0(D0_13), .d1(D8_13), .d2(D16_13), .d3(D24_13), 
        .sl0(n17), .sl1(n30) );
    mux4_3 U146 ( .x(n93), .d0(D0_14), .d1(D8_14), .d2(D16_14), .d3(D24_14), 
        .sl0(n23), .sl1(n30) );
    mux4_3 U147 ( .x(n94), .d0(D0_15), .d1(D8_15), .d2(D16_15), .d3(D24_15), 
        .sl0(n29), .sl1(n30) );
    mux4_3 U148 ( .x(n95), .d0(D0_16), .d1(D8_16), .d2(D16_16), .d3(D24_16), 
        .sl0(n11), .sl1(n31) );
    mux4_3 U149 ( .x(n96), .d0(D0_17), .d1(D8_17), .d2(D16_17), .d3(D24_17), 
        .sl0(n20), .sl1(n31) );
    mux4_2 U15 ( .x(n168), .d0(D2_25), .d1(D10_25), .d2(D18_25), .d3(D26_25), 
        .sl0(n19), .sl1(n35) );
    mux4_3 U150 ( .x(n97), .d0(D0_18), .d1(D8_18), .d2(D16_18), .d3(D24_18), 
        .sl0(n17), .sl1(n31) );
    mux4_3 U151 ( .x(n98), .d0(D0_19), .d1(D8_19), .d2(D16_19), .d3(D24_19), 
        .sl0(n18), .sl1(n31) );
    mux4_3 U152 ( .x(n99), .d0(D0_20), .d1(D8_20), .d2(D16_20), .d3(D24_20), 
        .sl0(n23), .sl1(n31) );
    mux4_3 U153 ( .x(n100), .d0(D0_21), .d1(D8_21), .d2(D16_21), .d3(D24_21), 
        .sl0(n18), .sl1(n31) );
    mux4_3 U154 ( .x(n101), .d0(D0_22), .d1(D8_22), .d2(D16_22), .d3(D24_22), 
        .sl0(n23), .sl1(n31) );
    mux4_3 U155 ( .x(n102), .d0(D0_23), .d1(D8_23), .d2(D16_23), .d3(D24_23), 
        .sl0(n28), .sl1(n31) );
    mux4_3 U156 ( .x(n103), .d0(D0_24), .d1(D8_24), .d2(D16_24), .d3(D24_24), 
        .sl0(n16), .sl1(n31) );
    mux4_3 U157 ( .x(n104), .d0(D0_25), .d1(D8_25), .d2(D16_25), .d3(D24_25), 
        .sl0(n29), .sl1(n31) );
    mux4_3 U158 ( .x(n105), .d0(D0_26), .d1(D8_26), .d2(D16_26), .d3(D24_26), 
        .sl0(n23), .sl1(n31) );
    mux4_3 U159 ( .x(n106), .d0(D0_27), .d1(D8_27), .d2(D16_27), .d3(D24_27), 
        .sl0(n23), .sl1(n31) );
    mux4_2 U16 ( .x(n123), .d0(D4_12), .d1(D12_12), .d2(D20_12), .d3(D28_12), 
        .sl0(n15), .sl1(n32) );
    mux4_3 U160 ( .x(n107), .d0(D0_28), .d1(D8_28), .d2(D16_28), .d3(D24_28), 
        .sl0(n23), .sl1(n31) );
    mux4_3 U161 ( .x(n108), .d0(D0_29), .d1(D8_29), .d2(D16_29), .d3(D24_29), 
        .sl0(n18), .sl1(n31) );
    mux4_3 U162 ( .x(n109), .d0(D0_30), .d1(D8_30), .d2(D16_30), .d3(D24_30), 
        .sl0(n23), .sl1(n31) );
    mux4_3 U163 ( .x(n110), .d0(D0_31), .d1(D8_31), .d2(D16_31), .d3(D24_31), 
        .sl0(n23), .sl1(n31) );
    mux4_3 U164 ( .x(n112), .d0(D4_1), .d1(D12_1), .d2(D20_1), .d3(D28_1), 
        .sl0(n16), .sl1(n32) );
    mux4_3 U165 ( .x(n113), .d0(D4_2), .d1(D12_2), .d2(D20_2), .d3(D28_2), 
        .sl0(n19), .sl1(n32) );
    mux4_3 U166 ( .x(n114), .d0(D4_3), .d1(D12_3), .d2(D20_3), .d3(D28_3), 
        .sl0(n23), .sl1(n32) );
    mux4_3 U167 ( .x(n115), .d0(D4_4), .d1(D12_4), .d2(D20_4), .d3(D28_4), 
        .sl0(n19), .sl1(n32) );
    mux4_3 U168 ( .x(n116), .d0(D4_5), .d1(D12_5), .d2(D20_5), .d3(D28_5), 
        .sl0(n11), .sl1(n32) );
    mux4_3 U169 ( .x(n117), .d0(D4_6), .d1(D12_6), .d2(D20_6), .d3(D28_6), 
        .sl0(n19), .sl1(n32) );
    mux4_2 U17 ( .x(n91), .d0(D0_12), .d1(D8_12), .d2(D16_12), .d3(D24_12), 
        .sl0(n17), .sl1(n30) );
    mux4_3 U170 ( .x(n118), .d0(D4_7), .d1(D12_7), .d2(D20_7), .d3(D28_7), 
        .sl0(n29), .sl1(n32) );
    mux4_3 U171 ( .x(n120), .d0(D4_9), .d1(D12_9), .d2(D20_9), .d3(D28_9), 
        .sl0(n11), .sl1(n32) );
    mux4_3 U172 ( .x(n121), .d0(D4_10), .d1(D12_10), .d2(D20_10), .d3(D28_10), 
        .sl0(n24), .sl1(n32) );
    mux4_3 U173 ( .x(n124), .d0(D4_13), .d1(D12_13), .d2(D20_13), .d3(D28_13), 
        .sl0(n26), .sl1(n32) );
    mux4_3 U174 ( .x(n125), .d0(D4_14), .d1(D12_14), .d2(D20_14), .d3(D28_14), 
        .sl0(n15), .sl1(n32) );
    mux4_3 U175 ( .x(n126), .d0(D4_15), .d1(D12_15), .d2(D20_15), .d3(D28_15), 
        .sl0(n24), .sl1(n32) );
    mux4_3 U176 ( .x(n127), .d0(D4_16), .d1(D12_16), .d2(D20_16), .d3(D28_16), 
        .sl0(n24), .sl1(n33) );
    mux4_3 U177 ( .x(n128), .d0(D4_17), .d1(D12_17), .d2(D20_17), .d3(D28_17), 
        .sl0(n15), .sl1(n33) );
    mux4_3 U178 ( .x(n129), .d0(D4_18), .d1(D12_18), .d2(D20_18), .d3(D28_18), 
        .sl0(n24), .sl1(n33) );
    mux4_3 U179 ( .x(n130), .d0(D4_19), .d1(D12_19), .d2(D20_19), .d3(D28_19), 
        .sl0(n29), .sl1(n33) );
    buf_8 U18 ( .x(n41), .a(S4) );
    mux4_3 U180 ( .x(n131), .d0(D4_20), .d1(D12_20), .d2(D20_20), .d3(D28_20), 
        .sl0(n24), .sl1(n33) );
    mux4_3 U181 ( .x(n132), .d0(D4_21), .d1(D12_21), .d2(D20_21), .d3(D28_21), 
        .sl0(n15), .sl1(n33) );
    mux4_3 U182 ( .x(n133), .d0(D4_22), .d1(D12_22), .d2(D20_22), .d3(D28_22), 
        .sl0(n13), .sl1(n33) );
    mux4_3 U183 ( .x(n134), .d0(D4_23), .d1(D12_23), .d2(D20_23), .d3(D28_23), 
        .sl0(n19), .sl1(n33) );
    mux4_3 U184 ( .x(n135), .d0(D4_24), .d1(D12_24), .d2(D20_24), .d3(D28_24), 
        .sl0(n15), .sl1(n33) );
    mux4_3 U185 ( .x(n137), .d0(D4_26), .d1(D12_26), .d2(D20_26), .d3(D28_26), 
        .sl0(n17), .sl1(n33) );
    mux4_3 U186 ( .x(n138), .d0(D4_27), .d1(D12_27), .d2(D20_27), .d3(D28_27), 
        .sl0(n24), .sl1(n33) );
    mux4_3 U187 ( .x(n139), .d0(D4_28), .d1(D12_28), .d2(D20_28), .d3(D28_28), 
        .sl0(n20), .sl1(n33) );
    mux4_3 U188 ( .x(n140), .d0(D4_29), .d1(D12_29), .d2(D20_29), .d3(D28_29), 
        .sl0(n24), .sl1(n33) );
    mux4_3 U189 ( .x(n141), .d0(D4_30), .d1(D12_30), .d2(D20_30), .d3(D28_30), 
        .sl0(n24), .sl1(n33) );
    buf_8 U19 ( .x(n35), .a(S4) );
    mux4_3 U190 ( .x(n142), .d0(D4_31), .d1(D12_31), .d2(D20_31), .d3(D28_31), 
        .sl0(n15), .sl1(n33) );
    mux4_3 U191 ( .x(n144), .d0(D2_1), .d1(D10_1), .d2(D18_1), .d3(D26_1), 
        .sl0(n26), .sl1(n34) );
    mux4_3 U192 ( .x(n145), .d0(D2_2), .d1(D10_2), .d2(D18_2), .d3(D26_2), 
        .sl0(n24), .sl1(n34) );
    mux4_3 U193 ( .x(n146), .d0(D2_3), .d1(D10_3), .d2(D18_3), .d3(D26_3), 
        .sl0(n24), .sl1(n34) );
    mux4_3 U194 ( .x(n147), .d0(D2_4), .d1(D10_4), .d2(D18_4), .d3(D26_4), 
        .sl0(n15), .sl1(n34) );
    mux4_3 U195 ( .x(n148), .d0(D2_5), .d1(D10_5), .d2(D18_5), .d3(D26_5), 
        .sl0(n24), .sl1(n34) );
    mux4_3 U196 ( .x(n149), .d0(D2_6), .d1(D10_6), .d2(D18_6), .d3(D26_6), 
        .sl0(n24), .sl1(n34) );
    mux4_3 U197 ( .x(n150), .d0(D2_7), .d1(D10_7), .d2(D18_7), .d3(D26_7), 
        .sl0(n20), .sl1(n34) );
    mux4_3 U198 ( .x(n151), .d0(D2_8), .d1(D10_8), .d2(D18_8), .d3(D26_8), 
        .sl0(n25), .sl1(n34) );
    mux4_3 U199 ( .x(n152), .d0(D2_9), .d1(D10_9), .d2(D18_9), .d3(D26_9), 
        .sl0(n15), .sl1(n34) );
    mux4_2 U2 ( .x(n143), .d0(D2_0), .d1(D10_0), .d2(D18_0), .d3(D26_0), .sl0(
        n15), .sl1(n34) );
    mux4_2 U20 ( .x(n211), .d0(n243), .d1(n307), .d2(n275), .d3(n339), .sl0(n4
        ), .sl1(n2) );
    mux4_3 U200 ( .x(n153), .d0(D2_10), .d1(D10_10), .d2(D18_10), .d3(D26_10), 
        .sl0(n20), .sl1(n34) );
    mux4_3 U201 ( .x(n155), .d0(D2_12), .d1(D10_12), .d2(D18_12), .d3(D26_12), 
        .sl0(n25), .sl1(n34) );
    mux4_3 U202 ( .x(n156), .d0(D2_13), .d1(D10_13), .d2(D18_13), .d3(D26_13), 
        .sl0(n13), .sl1(n34) );
    mux4_3 U203 ( .x(n157), .d0(D2_14), .d1(D10_14), .d2(D18_14), .d3(D26_14), 
        .sl0(n20), .sl1(n34) );
    mux4_3 U204 ( .x(n158), .d0(D2_15), .d1(D10_15), .d2(D18_15), .d3(D26_15), 
        .sl0(n28), .sl1(n34) );
    mux4_3 U205 ( .x(n159), .d0(D2_16), .d1(D10_16), .d2(D18_16), .d3(D26_16), 
        .sl0(n15), .sl1(n35) );
    mux4_3 U206 ( .x(n160), .d0(D2_17), .d1(D10_17), .d2(D18_17), .d3(D26_17), 
        .sl0(n25), .sl1(n35) );
    mux4_3 U207 ( .x(n161), .d0(D2_18), .d1(D10_18), .d2(D18_18), .d3(D26_18), 
        .sl0(n13), .sl1(n35) );
    mux4_3 U208 ( .x(n162), .d0(D2_19), .d1(D10_19), .d2(D18_19), .d3(D26_19), 
        .sl0(n25), .sl1(n35) );
    mux4_3 U209 ( .x(n163), .d0(D2_20), .d1(D10_20), .d2(D18_20), .d3(D26_20), 
        .sl0(n25), .sl1(n35) );
    mux4_2 U21 ( .x(n51), .d0(n83), .d1(n147), .d2(n115), .d3(n179), .sl0(n3), 
        .sl1(n2) );
    mux4_3 U210 ( .x(n164), .d0(D2_21), .d1(D10_21), .d2(D18_21), .d3(D26_21), 
        .sl0(n15), .sl1(n35) );
    mux4_3 U211 ( .x(n165), .d0(D2_22), .d1(D10_22), .d2(D18_22), .d3(D26_22), 
        .sl0(n15), .sl1(n35) );
    mux4_3 U212 ( .x(n166), .d0(D2_23), .d1(D10_23), .d2(D18_23), .d3(D26_23), 
        .sl0(n18), .sl1(n35) );
    mux4_3 U213 ( .x(n167), .d0(D2_24), .d1(D10_24), .d2(D18_24), .d3(D26_24), 
        .sl0(n25), .sl1(n35) );
    mux4_3 U214 ( .x(n169), .d0(D2_26), .d1(D10_26), .d2(D18_26), .d3(D26_26), 
        .sl0(n25), .sl1(n35) );
    mux4_3 U215 ( .x(n170), .d0(D2_27), .d1(D10_27), .d2(D18_27), .d3(D26_27), 
        .sl0(n20), .sl1(n35) );
    mux4_3 U216 ( .x(n171), .d0(D2_28), .d1(D10_28), .d2(D18_28), .d3(D26_28), 
        .sl0(n14), .sl1(n35) );
    mux4_3 U217 ( .x(n172), .d0(D2_29), .d1(D10_29), .d2(D18_29), .d3(D26_29), 
        .sl0(n14), .sl1(n35) );
    mux4_3 U218 ( .x(n173), .d0(D2_30), .d1(D10_30), .d2(D18_30), .d3(D26_30), 
        .sl0(n14), .sl1(n35) );
    mux4_3 U219 ( .x(n174), .d0(D2_31), .d1(D10_31), .d2(D18_31), .d3(D26_31), 
        .sl0(n25), .sl1(n35) );
    mux4_2 U22 ( .x(n214), .d0(n246), .d1(n310), .d2(n278), .d3(n342), .sl0(n3
        ), .sl1(n2) );
    mux4_3 U220 ( .x(n175), .d0(D6_0), .d1(D14_0), .d2(D22_0), .d3(D30_0), 
        .sl0(n25), .sl1(n36) );
    mux4_3 U221 ( .x(n176), .d0(D6_1), .d1(D14_1), .d2(D22_1), .d3(D30_1), 
        .sl0(n29), .sl1(n36) );
    mux4_3 U222 ( .x(n177), .d0(D6_2), .d1(D14_2), .d2(D22_2), .d3(D30_2), 
        .sl0(n25), .sl1(n36) );
    mux4_3 U223 ( .x(n178), .d0(D6_3), .d1(D14_3), .d2(D22_3), .d3(D30_3), 
        .sl0(n25), .sl1(n36) );
    mux4_3 U224 ( .x(n179), .d0(D6_4), .d1(D14_4), .d2(D22_4), .d3(D30_4), 
        .sl0(n14), .sl1(n36) );
    mux4_3 U225 ( .x(n180), .d0(D6_5), .d1(D14_5), .d2(D22_5), .d3(D30_5), 
        .sl0(n29), .sl1(n36) );
    mux4_3 U226 ( .x(n181), .d0(D6_6), .d1(D14_6), .d2(D22_6), .d3(D30_6), 
        .sl0(n14), .sl1(n36) );
    mux4_3 U227 ( .x(n182), .d0(D6_7), .d1(D14_7), .d2(D22_7), .d3(D30_7), 
        .sl0(n14), .sl1(n36) );
    mux4_3 U228 ( .x(n184), .d0(D6_9), .d1(D14_9), .d2(D22_9), .d3(D30_9), 
        .sl0(n18), .sl1(n36) );
    mux4_3 U229 ( .x(n185), .d0(D6_10), .d1(D14_10), .d2(D22_10), .d3(D30_10), 
        .sl0(n19), .sl1(n36) );
    inv_3 U23 ( .x(Z_1), .a(n5) );
    mux4_3 U230 ( .x(n186), .d0(D6_11), .d1(D14_11), .d2(D22_11), .d3(D30_11), 
        .sl0(n14), .sl1(n36) );
    mux4_3 U231 ( .x(n187), .d0(D6_12), .d1(D14_12), .d2(D22_12), .d3(D30_12), 
        .sl0(n25), .sl1(n36) );
    mux4_3 U232 ( .x(n188), .d0(D6_13), .d1(D14_13), .d2(D22_13), .d3(D30_13), 
        .sl0(n18), .sl1(n36) );
    mux4_3 U233 ( .x(n189), .d0(D6_14), .d1(D14_14), .d2(D22_14), .d3(D30_14), 
        .sl0(n25), .sl1(n36) );
    mux4_3 U234 ( .x(n190), .d0(D6_15), .d1(D14_15), .d2(D22_15), .d3(D30_15), 
        .sl0(n25), .sl1(n36) );
    mux4_3 U235 ( .x(n191), .d0(D6_16), .d1(D14_16), .d2(D22_16), .d3(D30_16), 
        .sl0(n14), .sl1(n37) );
    mux4_3 U236 ( .x(n192), .d0(D6_17), .d1(D14_17), .d2(D22_17), .d3(D30_17), 
        .sl0(n11), .sl1(n37) );
    mux4_3 U237 ( .x(n193), .d0(D6_18), .d1(D14_18), .d2(D22_18), .d3(D30_18), 
        .sl0(n28), .sl1(n37) );
    mux4_3 U238 ( .x(n194), .d0(D6_19), .d1(D14_19), .d2(D22_19), .d3(D30_19), 
        .sl0(n14), .sl1(n37) );
    mux4_3 U239 ( .x(n195), .d0(D6_20), .d1(D14_20), .d2(D22_20), .d3(D30_20), 
        .sl0(n14), .sl1(n37) );
    mux4_3 U240 ( .x(n196), .d0(D6_21), .d1(D14_21), .d2(D22_21), .d3(D30_21), 
        .sl0(n14), .sl1(n37) );
    mux4_3 U241 ( .x(n197), .d0(D6_22), .d1(D14_22), .d2(D22_22), .d3(D30_22), 
        .sl0(n14), .sl1(n37) );
    mux4_3 U242 ( .x(n198), .d0(D6_23), .d1(D14_23), .d2(D22_23), .d3(D30_23), 
        .sl0(n28), .sl1(n37) );
    mux4_3 U243 ( .x(n199), .d0(D6_24), .d1(D14_24), .d2(D22_24), .d3(D30_24), 
        .sl0(n16), .sl1(n37) );
    mux4_3 U244 ( .x(n200), .d0(D6_25), .d1(D14_25), .d2(D22_25), .d3(D30_25), 
        .sl0(n13), .sl1(n37) );
    mux4_3 U245 ( .x(n201), .d0(D6_26), .d1(D14_26), .d2(D22_26), .d3(D30_26), 
        .sl0(n29), .sl1(n37) );
    mux4_3 U246 ( .x(n202), .d0(D6_27), .d1(D14_27), .d2(D22_27), .d3(D30_27), 
        .sl0(n22), .sl1(n37) );
    mux4_3 U247 ( .x(n203), .d0(D6_28), .d1(D14_28), .d2(D22_28), .d3(D30_28), 
        .sl0(n14), .sl1(n37) );
    mux4_3 U248 ( .x(n204), .d0(D6_29), .d1(D14_29), .d2(D22_29), .d3(D30_29), 
        .sl0(n18), .sl1(n37) );
    mux4_3 U249 ( .x(n205), .d0(D6_30), .d1(D14_30), .d2(D22_30), .d3(D30_30), 
        .sl0(n29), .sl1(n37) );
    mux4_2 U25 ( .x(n232), .d0(n264), .d1(n328), .d2(n296), .d3(n360), .sl0(n3
        ), .sl1(n2) );
    mux4_3 U250 ( .x(n206), .d0(D6_31), .d1(D14_31), .d2(D22_31), .d3(D30_31), 
        .sl0(n26), .sl1(n37) );
    mux4_3 U251 ( .x(n207), .d0(n239), .d1(n303), .d2(n271), .d3(n335), .sl0(
        n4), .sl1(n1) );
    mux4_3 U252 ( .x(n209), .d0(n241), .d1(n305), .d2(n273), .d3(n337), .sl0(
        n4), .sl1(n2) );
    mux4_3 U253 ( .x(n210), .d0(n242), .d1(n306), .d2(n274), .d3(n338), .sl0(
        n4), .sl1(n2) );
    mux4_3 U254 ( .x(n212), .d0(n244), .d1(n308), .d2(n276), .d3(n340), .sl0(
        n3), .sl1(n1) );
    mux4_3 U255 ( .x(n213), .d0(n245), .d1(n309), .d2(n277), .d3(n341), .sl0(
        n3), .sl1(n1) );
    mux4_3 U256 ( .x(n215), .d0(n247), .d1(n311), .d2(n279), .d3(n343), .sl0(
        n9), .sl1(n1) );
    mux4_3 U257 ( .x(n216), .d0(n248), .d1(n312), .d2(n280), .d3(n344), .sl0(
        n9), .sl1(n1) );
    mux4_3 U258 ( .x(n217), .d0(n249), .d1(n313), .d2(n281), .d3(n345), .sl0(
        n9), .sl1(n1) );
    mux4_3 U259 ( .x(n218), .d0(n250), .d1(n314), .d2(n282), .d3(n346), .sl0(
        n3), .sl1(n1) );
    mux4_2 U26 ( .x(n59), .d0(n91), .d1(n155), .d2(n123), .d3(n187), .sl0(n3), 
        .sl1(n2) );
    mux4_3 U260 ( .x(n220), .d0(n252), .d1(n316), .d2(n284), .d3(n348), .sl0(
        n3), .sl1(n2) );
    mux4_3 U261 ( .x(n221), .d0(n253), .d1(n317), .d2(n285), .d3(n349), .sl0(
        n9), .sl1(n2) );
    mux4_3 U262 ( .x(n222), .d0(n254), .d1(n318), .d2(n286), .d3(n350), .sl0(
        n3), .sl1(n2) );
    mux4_3 U263 ( .x(n223), .d0(n255), .d1(n319), .d2(n287), .d3(n351), .sl0(
        n4), .sl1(n1) );
    mux4_3 U264 ( .x(n224), .d0(n256), .d1(n320), .d2(n288), .d3(n352), .sl0(
        n4), .sl1(n2) );
    mux4_3 U265 ( .x(n225), .d0(n257), .d1(n321), .d2(n289), .d3(n353), .sl0(
        n9), .sl1(n2) );
    mux4_3 U266 ( .x(n226), .d0(n258), .d1(n322), .d2(n290), .d3(n354), .sl0(
        n9), .sl1(n1) );
    mux4_3 U267 ( .x(n227), .d0(n259), .d1(n323), .d2(n291), .d3(n355), .sl0(
        n3), .sl1(n2) );
    mux4_3 U268 ( .x(n228), .d0(n260), .d1(n324), .d2(n292), .d3(n356), .sl0(
        n9), .sl1(n1) );
    mux4_3 U269 ( .x(n229), .d0(n261), .d1(n325), .d2(n293), .d3(n357), .sl0(
        n3), .sl1(n1) );
    mux4_2 U27 ( .x(n219), .d0(n251), .d1(n315), .d2(n283), .d3(n347), .sl0(n9
        ), .sl1(n2) );
    mux4_3 U270 ( .x(n231), .d0(n263), .d1(n327), .d2(n295), .d3(n359), .sl0(
        n4), .sl1(n1) );
    mux4_3 U271 ( .x(n233), .d0(n265), .d1(n329), .d2(n297), .d3(n361), .sl0(
        n10), .sl1(n1) );
    mux4_3 U272 ( .x(n235), .d0(n267), .d1(n331), .d2(n299), .d3(n363), .sl0(
        n10), .sl1(n1) );
    mux4_3 U273 ( .x(n236), .d0(n268), .d1(n332), .d2(n300), .d3(n364), .sl0(
        n10), .sl1(n1) );
    mux4_3 U274 ( .x(n238), .d0(n270), .d1(n334), .d2(n302), .d3(n366), .sl0(
        n4), .sl1(n1) );
    mux4_3 U275 ( .x(n239), .d0(D1_0), .d1(D9_0), .d2(D17_0), .d3(D25_0), 
        .sl0(n13), .sl1(n38) );
    mux4_3 U276 ( .x(n240), .d0(D1_1), .d1(D9_1), .d2(D17_1), .d3(D25_1), 
        .sl0(n13), .sl1(n38) );
    mux4_3 U277 ( .x(n241), .d0(D1_2), .d1(D9_2), .d2(D17_2), .d3(D25_2), 
        .sl0(n26), .sl1(n38) );
    mux4_3 U278 ( .x(n242), .d0(D1_3), .d1(D9_3), .d2(D17_3), .d3(D25_3), 
        .sl0(n20), .sl1(n38) );
    mux4_3 U279 ( .x(n243), .d0(D1_4), .d1(D9_4), .d2(D17_4), .d3(D25_4), 
        .sl0(n28), .sl1(n38) );
    mux2_2 U28 ( .x(Z_27), .d0(n74), .sl(S0), .d1(n234) );
    mux4_3 U280 ( .x(n244), .d0(D1_5), .d1(D9_5), .d2(D17_5), .d3(D25_5), 
        .sl0(n29), .sl1(n38) );
    mux4_3 U281 ( .x(n245), .d0(D1_6), .d1(D9_6), .d2(D17_6), .d3(D25_6), 
        .sl0(n28), .sl1(n38) );
    mux4_3 U282 ( .x(n246), .d0(D1_7), .d1(D9_7), .d2(D17_7), .d3(D25_7), 
        .sl0(n26), .sl1(n38) );
    mux4_3 U283 ( .x(n247), .d0(D1_8), .d1(D9_8), .d2(D17_8), .d3(D25_8), 
        .sl0(n29), .sl1(n38) );
    mux4_3 U284 ( .x(n248), .d0(D1_9), .d1(D9_9), .d2(D17_9), .d3(D25_9), 
        .sl0(n17), .sl1(n38) );
    mux4_3 U285 ( .x(n249), .d0(D1_10), .d1(D9_10), .d2(D17_10), .d3(D25_10), 
        .sl0(n19), .sl1(n38) );
    mux4_3 U286 ( .x(n251), .d0(D1_12), .d1(D9_12), .d2(D17_12), .d3(D25_12), 
        .sl0(n20), .sl1(n38) );
    mux4_3 U287 ( .x(n252), .d0(D1_13), .d1(D9_13), .d2(D17_13), .d3(D25_13), 
        .sl0(n26), .sl1(n38) );
    mux4_3 U288 ( .x(n253), .d0(D1_14), .d1(D9_14), .d2(D17_14), .d3(D25_14), 
        .sl0(n29), .sl1(n38) );
    mux4_3 U289 ( .x(n254), .d0(D1_15), .d1(D9_15), .d2(D17_15), .d3(D25_15), 
        .sl0(n20), .sl1(n38) );
    mux4_2 U29 ( .x(n74), .d0(n106), .d1(n170), .d2(n138), .d3(n202), .sl0(n9), 
        .sl1(n2) );
    mux4_3 U290 ( .x(n255), .d0(D1_16), .d1(D9_16), .d2(D17_16), .d3(D25_16), 
        .sl0(n26), .sl1(n39) );
    mux4_3 U291 ( .x(n256), .d0(D1_17), .d1(D9_17), .d2(D17_17), .d3(D25_17), 
        .sl0(n29), .sl1(n39) );
    mux4_3 U292 ( .x(n257), .d0(D1_18), .d1(D9_18), .d2(D17_18), .d3(D25_18), 
        .sl0(n19), .sl1(n39) );
    mux4_3 U293 ( .x(n258), .d0(D1_19), .d1(D9_19), .d2(D17_19), .d3(D25_19), 
        .sl0(n16), .sl1(n39) );
    mux4_3 U294 ( .x(n259), .d0(D1_20), .d1(D9_20), .d2(D17_20), .d3(D25_20), 
        .sl0(n17), .sl1(n39) );
    mux4_3 U295 ( .x(n260), .d0(D1_21), .d1(D9_21), .d2(D17_21), .d3(D25_21), 
        .sl0(n28), .sl1(n39) );
    mux4_3 U296 ( .x(n261), .d0(D1_22), .d1(D9_22), .d2(D17_22), .d3(D25_22), 
        .sl0(n19), .sl1(n39) );
    mux4_3 U297 ( .x(n262), .d0(D1_23), .d1(D9_23), .d2(D17_23), .d3(D25_23), 
        .sl0(n13), .sl1(n39) );
    mux4_3 U298 ( .x(n263), .d0(D1_24), .d1(D9_24), .d2(D17_24), .d3(D25_24), 
        .sl0(n26), .sl1(n39) );
    mux4_3 U299 ( .x(n264), .d0(D1_25), .d1(D9_25), .d2(D17_25), .d3(D25_25), 
        .sl0(n25), .sl1(n39) );
    mux4_2 U3 ( .x(n79), .d0(D0_0), .d1(D8_0), .d2(D16_0), .d3(D24_0), .sl0(
        n17), .sl1(n30) );
    mux4_2 U30 ( .x(n234), .d0(n266), .d1(n330), .d2(n298), .d3(n362), .sl0(n4
        ), .sl1(n2) );
    mux4_3 U300 ( .x(n265), .d0(D1_26), .d1(D9_26), .d2(D17_26), .d3(D25_26), 
        .sl0(n13), .sl1(n39) );
    mux4_3 U301 ( .x(n266), .d0(D1_27), .d1(D9_27), .d2(D17_27), .d3(D25_27), 
        .sl0(n16), .sl1(n39) );
    mux4_3 U302 ( .x(n267), .d0(D1_28), .d1(D9_28), .d2(D17_28), .d3(D25_28), 
        .sl0(n20), .sl1(n39) );
    mux4_3 U303 ( .x(n268), .d0(D1_29), .d1(D9_29), .d2(D17_29), .d3(D25_29), 
        .sl0(n13), .sl1(n39) );
    mux4_3 U304 ( .x(n269), .d0(D1_30), .d1(D9_30), .d2(D17_30), .d3(D25_30), 
        .sl0(n21), .sl1(n39) );
    mux4_3 U305 ( .x(n270), .d0(D1_31), .d1(D9_31), .d2(D17_31), .d3(D25_31), 
        .sl0(n19), .sl1(n39) );
    mux4_3 U306 ( .x(n271), .d0(D5_0), .d1(D13_0), .d2(D21_0), .d3(D29_0), 
        .sl0(n20), .sl1(n40) );
    mux4_3 U307 ( .x(n272), .d0(D5_1), .d1(D13_1), .d2(D21_1), .d3(D29_1), 
        .sl0(n11), .sl1(n40) );
    mux4_3 U308 ( .x(n273), .d0(D5_2), .d1(D13_2), .d2(D21_2), .d3(D29_2), 
        .sl0(n13), .sl1(n40) );
    mux4_3 U309 ( .x(n274), .d0(D5_3), .d1(D13_3), .d2(D21_3), .d3(D29_3), 
        .sl0(n11), .sl1(n40) );
    mux4_2 U31 ( .x(n65), .d0(n97), .d1(n161), .d2(n129), .d3(n193), .sl0(n3), 
        .sl1(n2) );
    mux4_3 U310 ( .x(n275), .d0(D5_4), .d1(D13_4), .d2(D21_4), .d3(D29_4), 
        .sl0(n21), .sl1(n40) );
    mux4_3 U311 ( .x(n276), .d0(D5_5), .d1(D13_5), .d2(D21_5), .d3(D29_5), 
        .sl0(n18), .sl1(n40) );
    mux4_3 U312 ( .x(n277), .d0(D5_6), .d1(D13_6), .d2(D21_6), .d3(D29_6), 
        .sl0(n17), .sl1(n40) );
    mux4_3 U313 ( .x(n278), .d0(D5_7), .d1(D13_7), .d2(D21_7), .d3(D29_7), 
        .sl0(n21), .sl1(n40) );
    mux4_3 U314 ( .x(n280), .d0(D5_9), .d1(D13_9), .d2(D21_9), .d3(D29_9), 
        .sl0(n12), .sl1(n40) );
    mux4_3 U315 ( .x(n281), .d0(D5_10), .d1(D13_10), .d2(D21_10), .d3(D29_10), 
        .sl0(n12), .sl1(n40) );
    mux4_3 U316 ( .x(n283), .d0(D5_12), .d1(D13_12), .d2(D21_12), .d3(D29_12), 
        .sl0(n21), .sl1(n40) );
    mux4_3 U317 ( .x(n284), .d0(D5_13), .d1(D13_13), .d2(D21_13), .d3(D29_13), 
        .sl0(n21), .sl1(n40) );
    mux4_3 U318 ( .x(n285), .d0(D5_14), .d1(D13_14), .d2(D21_14), .d3(D29_14), 
        .sl0(n27), .sl1(n40) );
    mux4_3 U319 ( .x(n286), .d0(D5_15), .d1(D13_15), .d2(D21_15), .d3(D29_15), 
        .sl0(n12), .sl1(n40) );
    mux4_2 U32 ( .x(n230), .d0(n262), .d1(n326), .d2(n294), .d3(n358), .sl0(n3
        ), .sl1(n2) );
    mux4_3 U320 ( .x(n287), .d0(D5_16), .d1(D13_16), .d2(D21_16), .d3(D29_16), 
        .sl0(n12), .sl1(n41) );
    mux4_3 U321 ( .x(n288), .d0(D5_17), .d1(D13_17), .d2(D21_17), .d3(D29_17), 
        .sl0(n21), .sl1(n41) );
    mux4_3 U322 ( .x(n289), .d0(D5_18), .d1(D13_18), .d2(D21_18), .d3(D29_18), 
        .sl0(n12), .sl1(n41) );
    mux4_3 U323 ( .x(n290), .d0(D5_19), .d1(D13_19), .d2(D21_19), .d3(D29_19), 
        .sl0(n27), .sl1(n41) );
    mux4_3 U324 ( .x(n291), .d0(D5_20), .d1(D13_20), .d2(D21_20), .d3(D29_20), 
        .sl0(n21), .sl1(n41) );
    mux4_3 U325 ( .x(n292), .d0(D5_21), .d1(D13_21), .d2(D21_21), .d3(D29_21), 
        .sl0(n27), .sl1(n41) );
    mux4_3 U326 ( .x(n293), .d0(D5_22), .d1(D13_22), .d2(D21_22), .d3(D29_22), 
        .sl0(n27), .sl1(n41) );
    mux4_3 U327 ( .x(n294), .d0(D5_23), .d1(D13_23), .d2(D21_23), .d3(D29_23), 
        .sl0(n12), .sl1(n41) );
    mux4_3 U328 ( .x(n295), .d0(D5_24), .d1(D13_24), .d2(D21_24), .d3(D29_24), 
        .sl0(n27), .sl1(n41) );
    mux4_3 U329 ( .x(n296), .d0(D5_25), .d1(D13_25), .d2(D21_25), .d3(D29_25), 
        .sl0(n27), .sl1(n41) );
    mux4_2 U33 ( .x(n70), .d0(n102), .d1(n166), .d2(n134), .d3(n198), .sl0(n3), 
        .sl1(n2) );
    mux4_3 U330 ( .x(n297), .d0(D5_26), .d1(D13_26), .d2(D21_26), .d3(D29_26), 
        .sl0(n27), .sl1(n41) );
    mux4_3 U331 ( .x(n298), .d0(D5_27), .d1(D13_27), .d2(D21_27), .d3(D29_27), 
        .sl0(n27), .sl1(n41) );
    mux4_3 U332 ( .x(n299), .d0(D5_28), .d1(D13_28), .d2(D21_28), .d3(D29_28), 
        .sl0(n27), .sl1(n41) );
    mux4_3 U333 ( .x(n300), .d0(D5_29), .d1(D13_29), .d2(D21_29), .d3(D29_29), 
        .sl0(n21), .sl1(n41) );
    mux4_3 U334 ( .x(n301), .d0(D5_30), .d1(D13_30), .d2(D21_30), .d3(D29_30), 
        .sl0(n21), .sl1(n41) );
    mux4_3 U335 ( .x(n302), .d0(D5_31), .d1(D13_31), .d2(D21_31), .d3(D29_31), 
        .sl0(n27), .sl1(n41) );
    mux4_3 U336 ( .x(n303), .d0(D3_0), .d1(D11_0), .d2(D19_0), .d3(D27_0), 
        .sl0(n12), .sl1(n42) );
    mux4_3 U337 ( .x(n304), .d0(D3_1), .d1(D11_1), .d2(D19_1), .d3(D27_1), 
        .sl0(n27), .sl1(n42) );
    mux4_3 U338 ( .x(n305), .d0(D3_2), .d1(D11_2), .d2(D19_2), .d3(D27_2), 
        .sl0(n27), .sl1(n42) );
    mux4_3 U339 ( .x(n306), .d0(D3_3), .d1(D11_3), .d2(D19_3), .d3(D27_3), 
        .sl0(n27), .sl1(n42) );
    mux4_2 U34 ( .x(n237), .d0(n269), .d1(n333), .d2(n301), .d3(n365), .sl0(
        n10), .sl1(n1) );
    mux4_3 U340 ( .x(n307), .d0(D3_4), .d1(D11_4), .d2(D19_4), .d3(D27_4), 
        .sl0(n12), .sl1(n42) );
    mux4_3 U341 ( .x(n308), .d0(D3_5), .d1(D11_5), .d2(D19_5), .d3(D27_5), 
        .sl0(n21), .sl1(n42) );
    mux4_3 U342 ( .x(n309), .d0(D3_6), .d1(D11_6), .d2(D19_6), .d3(D27_6), 
        .sl0(n27), .sl1(n42) );
    mux4_3 U343 ( .x(n310), .d0(D3_7), .d1(D11_7), .d2(D19_7), .d3(D27_7), 
        .sl0(n12), .sl1(n42) );
    mux4_3 U344 ( .x(n312), .d0(D3_9), .d1(D11_9), .d2(D19_9), .d3(D27_9), 
        .sl0(n21), .sl1(n42) );
    mux4_3 U345 ( .x(n313), .d0(D3_10), .d1(D11_10), .d2(D19_10), .d3(D27_10), 
        .sl0(n12), .sl1(n42) );
    mux4_3 U346 ( .x(n314), .d0(D3_11), .d1(D11_11), .d2(D19_11), .d3(D27_11), 
        .sl0(n12), .sl1(n42) );
    mux4_3 U347 ( .x(n315), .d0(D3_12), .d1(D11_12), .d2(D19_12), .d3(D27_12), 
        .sl0(n12), .sl1(n42) );
    mux4_3 U348 ( .x(n316), .d0(D3_13), .d1(D11_13), .d2(D19_13), .d3(D27_13), 
        .sl0(n16), .sl1(n42) );
    mux4_3 U349 ( .x(n317), .d0(D3_14), .d1(D11_14), .d2(D19_14), .d3(D27_14), 
        .sl0(n12), .sl1(n42) );
    mux4_2 U35 ( .x(n77), .d0(n109), .d1(n173), .d2(n141), .d3(n205), .sl0(n10
        ), .sl1(n1) );
    mux4_3 U350 ( .x(n318), .d0(D3_15), .d1(D11_15), .d2(D19_15), .d3(D27_15), 
        .sl0(n13), .sl1(n42) );
    mux4_3 U351 ( .x(n319), .d0(D3_16), .d1(D11_16), .d2(D19_16), .d3(D27_16), 
        .sl0(n16), .sl1(n43) );
    mux4_3 U352 ( .x(n320), .d0(D3_17), .d1(D11_17), .d2(D19_17), .d3(D27_17), 
        .sl0(n21), .sl1(n43) );
    mux4_3 U353 ( .x(n321), .d0(D3_18), .d1(D11_18), .d2(D19_18), .d3(D27_18), 
        .sl0(n21), .sl1(n43) );
    mux4_3 U354 ( .x(n322), .d0(D3_19), .d1(D11_19), .d2(D19_19), .d3(D27_19), 
        .sl0(n22), .sl1(n43) );
    mux4_3 U355 ( .x(n323), .d0(D3_20), .d1(D11_20), .d2(D19_20), .d3(D27_20), 
        .sl0(n22), .sl1(n43) );
    mux4_3 U356 ( .x(n324), .d0(D3_21), .d1(D11_21), .d2(D19_21), .d3(D27_21), 
        .sl0(n22), .sl1(n43) );
    mux4_3 U357 ( .x(n325), .d0(D3_22), .d1(D11_22), .d2(D19_22), .d3(D27_22), 
        .sl0(n16), .sl1(n43) );
    mux4_3 U358 ( .x(n326), .d0(D3_23), .d1(D11_23), .d2(D19_23), .d3(D27_23), 
        .sl0(n28), .sl1(n43) );
    mux4_3 U359 ( .x(n327), .d0(D3_24), .d1(D11_24), .d2(D19_24), .d3(D27_24), 
        .sl0(n22), .sl1(n43) );
    buf_10 U36 ( .x(n1), .a(S2) );
    mux4_3 U360 ( .x(n328), .d0(D3_25), .d1(D11_25), .d2(D19_25), .d3(D27_25), 
        .sl0(n26), .sl1(n43) );
    mux4_3 U361 ( .x(n329), .d0(D3_26), .d1(D11_26), .d2(D19_26), .d3(D27_26), 
        .sl0(n11), .sl1(n43) );
    mux4_3 U362 ( .x(n330), .d0(D3_27), .d1(D11_27), .d2(D19_27), .d3(D27_27), 
        .sl0(n18), .sl1(n43) );
    mux4_3 U363 ( .x(n331), .d0(D3_28), .d1(D11_28), .d2(D19_28), .d3(D27_28), 
        .sl0(n11), .sl1(n43) );
    mux4_3 U364 ( .x(n332), .d0(D3_29), .d1(D11_29), .d2(D19_29), .d3(D27_29), 
        .sl0(n20), .sl1(n43) );
    mux4_3 U365 ( .x(n333), .d0(D3_30), .d1(D11_30), .d2(D19_30), .d3(D27_30), 
        .sl0(n18), .sl1(n43) );
    mux4_3 U366 ( .x(n334), .d0(D3_31), .d1(D11_31), .d2(D19_31), .d3(D27_31), 
        .sl0(n20), .sl1(n43) );
    mux4_3 U367 ( .x(n335), .d0(D7_0), .d1(D15_0), .d2(D23_0), .d3(D31_0), 
        .sl0(n22), .sl1(n44) );
    mux4_3 U368 ( .x(n336), .d0(D7_1), .d1(D15_1), .d2(D23_1), .d3(D31_1), 
        .sl0(n29), .sl1(n44) );
    mux4_3 U369 ( .x(n337), .d0(D7_2), .d1(D15_2), .d2(D23_2), .d3(D31_2), 
        .sl0(n22), .sl1(n44) );
    buf_7 U37 ( .x(n2), .a(S2) );
    mux4_3 U370 ( .x(n338), .d0(D7_3), .d1(D15_3), .d2(D23_3), .d3(D31_3), 
        .sl0(n28), .sl1(n44) );
    mux4_3 U371 ( .x(n339), .d0(D7_4), .d1(D15_4), .d2(D23_4), .d3(D31_4), 
        .sl0(n22), .sl1(n44) );
    mux4_3 U372 ( .x(n340), .d0(D7_5), .d1(D15_5), .d2(D23_5), .d3(D31_5), 
        .sl0(n16), .sl1(n44) );
    mux4_3 U373 ( .x(n341), .d0(D7_6), .d1(D15_6), .d2(D23_6), .d3(D31_6), 
        .sl0(n11), .sl1(n44) );
    mux4_3 U374 ( .x(n342), .d0(D7_7), .d1(D15_7), .d2(D23_7), .d3(D31_7), 
        .sl0(n22), .sl1(n44) );
    mux4_3 U375 ( .x(n343), .d0(D7_8), .d1(D15_8), .d2(D23_8), .d3(D31_8), 
        .sl0(n29), .sl1(n44) );
    mux4_3 U376 ( .x(n344), .d0(D7_9), .d1(D15_9), .d2(D23_9), .d3(D31_9), 
        .sl0(n22), .sl1(n44) );
    mux4_3 U377 ( .x(n345), .d0(D7_10), .d1(D15_10), .d2(D23_10), .d3(D31_10), 
        .sl0(n22), .sl1(n44) );
    mux4_3 U378 ( .x(n346), .d0(D7_11), .d1(D15_11), .d2(D23_11), .d3(D31_11), 
        .sl0(n16), .sl1(n44) );
    mux4_3 U379 ( .x(n347), .d0(D7_12), .d1(D15_12), .d2(D23_12), .d3(D31_12), 
        .sl0(n26), .sl1(n44) );
    mux4_3 U380 ( .x(n348), .d0(D7_13), .d1(D15_13), .d2(D23_13), .d3(D31_13), 
        .sl0(n18), .sl1(n44) );
    mux4_3 U381 ( .x(n349), .d0(D7_14), .d1(D15_14), .d2(D23_14), .d3(D31_14), 
        .sl0(n17), .sl1(n44) );
    mux4_3 U382 ( .x(n350), .d0(D7_15), .d1(D15_15), .d2(D23_15), .d3(D31_15), 
        .sl0(n22), .sl1(n44) );
    mux4_3 U383 ( .x(n351), .d0(D7_16), .d1(D15_16), .d2(D23_16), .d3(D31_16), 
        .sl0(n17), .sl1(n45) );
    mux4_3 U384 ( .x(n352), .d0(D7_17), .d1(D15_17), .d2(D23_17), .d3(D31_17), 
        .sl0(n22), .sl1(n45) );
    mux4_3 U385 ( .x(n353), .d0(D7_18), .d1(D15_18), .d2(D23_18), .d3(D31_18), 
        .sl0(n20), .sl1(n45) );
    mux4_3 U386 ( .x(n354), .d0(D7_19), .d1(D15_19), .d2(D23_19), .d3(D31_19), 
        .sl0(n22), .sl1(n45) );
    mux4_3 U387 ( .x(n355), .d0(D7_20), .d1(D15_20), .d2(D23_20), .d3(D31_20), 
        .sl0(n13), .sl1(n45) );
    mux4_3 U388 ( .x(n356), .d0(D7_21), .d1(D15_21), .d2(D23_21), .d3(D31_21), 
        .sl0(n13), .sl1(n45) );
    mux4_3 U389 ( .x(n357), .d0(D7_22), .d1(D15_22), .d2(D23_22), .d3(D31_22), 
        .sl0(n19), .sl1(n45) );
    buf_14 U39 ( .x(n16), .a(n46) );
    mux4_3 U390 ( .x(n358), .d0(D7_23), .d1(D15_23), .d2(D23_23), .d3(D31_23), 
        .sl0(n13), .sl1(n45) );
    mux4_3 U391 ( .x(n359), .d0(D7_24), .d1(D15_24), .d2(D23_24), .d3(D31_24), 
        .sl0(n23), .sl1(n45) );
    mux4_3 U392 ( .x(n360), .d0(D7_25), .d1(D15_25), .d2(D23_25), .d3(D31_25), 
        .sl0(n23), .sl1(n45) );
    mux4_3 U393 ( .x(n361), .d0(D7_26), .d1(D15_26), .d2(D23_26), .d3(D31_26), 
        .sl0(n17), .sl1(n45) );
    mux4_3 U394 ( .x(n362), .d0(D7_27), .d1(D15_27), .d2(D23_27), .d3(D31_27), 
        .sl0(n18), .sl1(n45) );
    mux4_3 U395 ( .x(n363), .d0(D7_28), .d1(D15_28), .d2(D23_28), .d3(D31_28), 
        .sl0(n16), .sl1(n45) );
    mux4_3 U396 ( .x(n364), .d0(D7_29), .d1(D15_29), .d2(D23_29), .d3(D31_29), 
        .sl0(n16), .sl1(n45) );
    mux4_3 U397 ( .x(n365), .d0(D7_30), .d1(D15_30), .d2(D23_30), .d3(D31_30), 
        .sl0(n26), .sl1(n45) );
    mux4_3 U398 ( .x(n366), .d0(D7_31), .d1(D15_31), .d2(D23_31), .d3(D31_31), 
        .sl0(n11), .sl1(n45) );
    mux2_3 U399 ( .x(Z_0), .d0(n47), .sl(S0), .d1(n207) );
    mux4_2 U4 ( .x(n279), .d0(D5_8), .d1(D13_8), .d2(D21_8), .d3(D29_8), .sl0(
        n19), .sl1(n40) );
    buf_12 U40 ( .x(n28), .a(n46) );
    buf_14 U400 ( .x(n19), .a(n46) );
    inv_16 U401 ( .x(n7), .a(S3) );
    mux2_4 U402 ( .x(Z_25), .d0(n72), .sl(S0), .d1(n232) );
    buf_14 U41 ( .x(n42), .a(S4) );
    buf_10 U42 ( .x(n36), .a(S4) );
    buf_14 U43 ( .x(n37), .a(S4) );
    buf_10 U44 ( .x(n34), .a(S4) );
    buf_10 U45 ( .x(n30), .a(S4) );
    buf_10 U46 ( .x(n40), .a(S4) );
    buf_14 U47 ( .x(n31), .a(S4) );
    buf_12 U48 ( .x(n32), .a(S4) );
    buf_10 U49 ( .x(n33), .a(S4) );
    mux4_2 U5 ( .x(n311), .d0(D3_8), .d1(D11_8), .d2(D19_8), .d3(D27_8), .sl0(
        n21), .sl1(n42) );
    mux4_3 U50 ( .x(n208), .d0(n240), .d1(n304), .d2(n272), .d3(n336), .sl0(S1
        ), .sl1(n1) );
    buf_16 U51 ( .x(n4), .a(S1) );
    buf_16 U52 ( .x(n3), .a(S1) );
    buf_10 U53 ( .x(n10), .a(S1) );
    mux2i_3 U54 ( .x(n5), .d0(n208), .sl(n6), .d1(n48) );
    inv_2 U55 ( .x(n6), .a(S0) );
    inv_16 U56 ( .x(n8), .a(n7) );
    buf_10 U57 ( .x(n9), .a(S1) );
    buf_16 U58 ( .x(n11), .a(n46) );
    buf_16 U59 ( .x(n12), .a(n8) );
    mux4_2 U6 ( .x(n183), .d0(D6_8), .d1(D14_8), .d2(D22_8), .d3(D30_8), .sl0(
        n14), .sl1(n36) );
    buf_16 U60 ( .x(n13), .a(n46) );
    buf_16 U61 ( .x(n14), .a(n8) );
    buf_16 U62 ( .x(n15), .a(n8) );
    buf_16 U63 ( .x(n17), .a(n46) );
    buf_16 U64 ( .x(n18), .a(n46) );
    buf_16 U66 ( .x(n20), .a(n46) );
    buf_16 U67 ( .x(n21), .a(n8) );
    buf_16 U68 ( .x(n22), .a(n8) );
    buf_16 U69 ( .x(n23), .a(n8) );
    mux4_2 U7 ( .x(n119), .d0(D4_8), .d1(D12_8), .d2(D20_8), .d3(D28_8), .sl0(
        n24), .sl1(n32) );
    buf_16 U70 ( .x(n24), .a(n8) );
    buf_16 U71 ( .x(n25), .a(n8) );
    buf_16 U72 ( .x(n26), .a(n46) );
    buf_16 U73 ( .x(n27), .a(n8) );
    buf_16 U74 ( .x(n29), .a(n46) );
    buf_16 U75 ( .x(n38), .a(S4) );
    buf_16 U76 ( .x(n39), .a(S4) );
    buf_16 U77 ( .x(n43), .a(S4) );
    buf_16 U78 ( .x(n44), .a(S4) );
    buf_16 U79 ( .x(n45), .a(S4) );
    mux4_2 U8 ( .x(n87), .d0(D0_8), .d1(D8_8), .d2(D16_8), .d3(D24_8), .sl0(
        n23), .sl1(n30) );
    inv_16 U80 ( .x(n46), .a(n7) );
    mux2_4 U82 ( .x(Z_2), .d0(n49), .sl(S0), .d1(n209) );
    mux2_4 U83 ( .x(Z_3), .d0(n50), .sl(S0), .d1(n210) );
    mux2_4 U84 ( .x(Z_4), .d0(n51), .sl(S0), .d1(n211) );
    mux2_4 U85 ( .x(Z_5), .d0(n52), .sl(S0), .d1(n212) );
    mux2_4 U86 ( .x(Z_6), .d0(n53), .sl(S0), .d1(n213) );
    mux2_4 U87 ( .x(Z_7), .d0(n54), .sl(S0), .d1(n214) );
    mux2_4 U88 ( .x(Z_8), .d0(n55), .sl(S0), .d1(n215) );
    mux2_4 U89 ( .x(Z_9), .d0(n56), .sl(S0), .d1(n216) );
    mux4_2 U9 ( .x(n282), .d0(D5_11), .d1(D13_11), .d2(D21_11), .d3(D29_11), 
        .sl0(n12), .sl1(n40) );
    mux2_4 U90 ( .x(Z_10), .d0(n57), .sl(S0), .d1(n217) );
    mux2_4 U91 ( .x(Z_11), .d0(n58), .sl(S0), .d1(n218) );
    mux2_4 U92 ( .x(Z_12), .d0(n59), .sl(S0), .d1(n219) );
    mux2_4 U93 ( .x(Z_13), .d0(n60), .sl(S0), .d1(n220) );
    mux2_4 U94 ( .x(Z_14), .d0(n61), .sl(S0), .d1(n221) );
    mux2_4 U95 ( .x(Z_15), .d0(n62), .sl(S0), .d1(n222) );
    mux2_4 U96 ( .x(Z_16), .d0(n63), .sl(S0), .d1(n223) );
    mux2_4 U97 ( .x(Z_17), .d0(n64), .sl(S0), .d1(n224) );
    mux2_4 U98 ( .x(Z_18), .d0(n65), .sl(S0), .d1(n225) );
    mux2_4 U99 ( .x(Z_19), .d0(n66), .sl(S0), .d1(n226) );
endmodule


module DLX_sync_MUX_OP_32_5_32_test_1 ( D0_31, D0_30, D0_29, D0_28, D0_27, 
    D0_26, D0_25, D0_24, D0_23, D0_22, D0_21, D0_20, D0_19, D0_18, D0_17, 
    D0_16, D0_15, D0_14, D0_13, D0_12, D0_11, D0_10, D0_9, D0_8, D0_7, D0_6, 
    D0_5, D0_4, D0_3, D0_2, D0_1, D0_0, D1_31, D1_30, D1_29, D1_28, D1_27, 
    D1_26, D1_25, D1_24, D1_23, D1_22, D1_21, D1_20, D1_19, D1_18, D1_17, 
    D1_16, D1_15, D1_14, D1_13, D1_12, D1_11, D1_10, D1_9, D1_8, D1_7, D1_6, 
    D1_5, D1_4, D1_3, D1_2, D1_1, D1_0, D2_31, D2_30, D2_29, D2_28, D2_27, 
    D2_26, D2_25, D2_24, D2_23, D2_22, D2_21, D2_20, D2_19, D2_18, D2_17, 
    D2_16, D2_15, D2_14, D2_13, D2_12, D2_11, D2_10, D2_9, D2_8, D2_7, D2_6, 
    D2_5, D2_4, D2_3, D2_2, D2_1, D2_0, D3_31, D3_30, D3_29, D3_28, D3_27, 
    D3_26, D3_25, D3_24, D3_23, D3_22, D3_21, D3_20, D3_19, D3_18, D3_17, 
    D3_16, D3_15, D3_14, D3_13, D3_12, D3_11, D3_10, D3_9, D3_8, D3_7, D3_6, 
    D3_5, D3_4, D3_3, D3_2, D3_1, D3_0, D4_31, D4_30, D4_29, D4_28, D4_27, 
    D4_26, D4_25, D4_24, D4_23, D4_22, D4_21, D4_20, D4_19, D4_18, D4_17, 
    D4_16, D4_15, D4_14, D4_13, D4_12, D4_11, D4_10, D4_9, D4_8, D4_7, D4_6, 
    D4_5, D4_4, D4_3, D4_2, D4_1, D4_0, D5_31, D5_30, D5_29, D5_28, D5_27, 
    D5_26, D5_25, D5_24, D5_23, D5_22, D5_21, D5_20, D5_19, D5_18, D5_17, 
    D5_16, D5_15, D5_14, D5_13, D5_12, D5_11, D5_10, D5_9, D5_8, D5_7, D5_6, 
    D5_5, D5_4, D5_3, D5_2, D5_1, D5_0, D6_31, D6_30, D6_29, D6_28, D6_27, 
    D6_26, D6_25, D6_24, D6_23, D6_22, D6_21, D6_20, D6_19, D6_18, D6_17, 
    D6_16, D6_15, D6_14, D6_13, D6_12, D6_11, D6_10, D6_9, D6_8, D6_7, D6_6, 
    D6_5, D6_4, D6_3, D6_2, D6_1, D6_0, D7_31, D7_30, D7_29, D7_28, D7_27, 
    D7_26, D7_25, D7_24, D7_23, D7_22, D7_21, D7_20, D7_19, D7_18, D7_17, 
    D7_16, D7_15, D7_14, D7_13, D7_12, D7_11, D7_10, D7_9, D7_8, D7_7, D7_6, 
    D7_5, D7_4, D7_3, D7_2, D7_1, D7_0, D8_31, D8_30, D8_29, D8_28, D8_27, 
    D8_26, D8_25, D8_24, D8_23, D8_22, D8_21, D8_20, D8_19, D8_18, D8_17, 
    D8_16, D8_15, D8_14, D8_13, D8_12, D8_11, D8_10, D8_9, D8_8, D8_7, D8_6, 
    D8_5, D8_4, D8_3, D8_2, D8_1, D8_0, D9_31, D9_30, D9_29, D9_28, D9_27, 
    D9_26, D9_25, D9_24, D9_23, D9_22, D9_21, D9_20, D9_19, D9_18, D9_17, 
    D9_16, D9_15, D9_14, D9_13, D9_12, D9_11, D9_10, D9_9, D9_8, D9_7, D9_6, 
    D9_5, D9_4, D9_3, D9_2, D9_1, D9_0, D10_31, D10_30, D10_29, D10_28, D10_27, 
    D10_26, D10_25, D10_24, D10_23, D10_22, D10_21, D10_20, D10_19, D10_18, 
    D10_17, D10_16, D10_15, D10_14, D10_13, D10_12, D10_11, D10_10, D10_9, 
    D10_8, D10_7, D10_6, D10_5, D10_4, D10_3, D10_2, D10_1, D10_0, D11_31, 
    D11_30, D11_29, D11_28, D11_27, D11_26, D11_25, D11_24, D11_23, D11_22, 
    D11_21, D11_20, D11_19, D11_18, D11_17, D11_16, D11_15, D11_14, D11_13, 
    D11_12, D11_11, D11_10, D11_9, D11_8, D11_7, D11_6, D11_5, D11_4, D11_3, 
    D11_2, D11_1, D11_0, D12_31, D12_30, D12_29, D12_28, D12_27, D12_26, 
    D12_25, D12_24, D12_23, D12_22, D12_21, D12_20, D12_19, D12_18, D12_17, 
    D12_16, D12_15, D12_14, D12_13, D12_12, D12_11, D12_10, D12_9, D12_8, 
    D12_7, D12_6, D12_5, D12_4, D12_3, D12_2, D12_1, D12_0, D13_31, D13_30, 
    D13_29, D13_28, D13_27, D13_26, D13_25, D13_24, D13_23, D13_22, D13_21, 
    D13_20, D13_19, D13_18, D13_17, D13_16, D13_15, D13_14, D13_13, D13_12, 
    D13_11, D13_10, D13_9, D13_8, D13_7, D13_6, D13_5, D13_4, D13_3, D13_2, 
    D13_1, D13_0, D14_31, D14_30, D14_29, D14_28, D14_27, D14_26, D14_25, 
    D14_24, D14_23, D14_22, D14_21, D14_20, D14_19, D14_18, D14_17, D14_16, 
    D14_15, D14_14, D14_13, D14_12, D14_11, D14_10, D14_9, D14_8, D14_7, D14_6, 
    D14_5, D14_4, D14_3, D14_2, D14_1, D14_0, D15_31, D15_30, D15_29, D15_28, 
    D15_27, D15_26, D15_25, D15_24, D15_23, D15_22, D15_21, D15_20, D15_19, 
    D15_18, D15_17, D15_16, D15_15, D15_14, D15_13, D15_12, D15_11, D15_10, 
    D15_9, D15_8, D15_7, D15_6, D15_5, D15_4, D15_3, D15_2, D15_1, D15_0, 
    D16_31, D16_30, D16_29, D16_28, D16_27, D16_26, D16_25, D16_24, D16_23, 
    D16_22, D16_21, D16_20, D16_19, D16_18, D16_17, D16_16, D16_15, D16_14, 
    D16_13, D16_12, D16_11, D16_10, D16_9, D16_8, D16_7, D16_6, D16_5, D16_4, 
    D16_3, D16_2, D16_1, D16_0, D17_31, D17_30, D17_29, D17_28, D17_27, D17_26, 
    D17_25, D17_24, D17_23, D17_22, D17_21, D17_20, D17_19, D17_18, D17_17, 
    D17_16, D17_15, D17_14, D17_13, D17_12, D17_11, D17_10, D17_9, D17_8, 
    D17_7, D17_6, D17_5, D17_4, D17_3, D17_2, D17_1, D17_0, D18_31, D18_30, 
    D18_29, D18_28, D18_27, D18_26, D18_25, D18_24, D18_23, D18_22, D18_21, 
    D18_20, D18_19, D18_18, D18_17, D18_16, D18_15, D18_14, D18_13, D18_12, 
    D18_11, D18_10, D18_9, D18_8, D18_7, D18_6, D18_5, D18_4, D18_3, D18_2, 
    D18_1, D18_0, D19_31, D19_30, D19_29, D19_28, D19_27, D19_26, D19_25, 
    D19_24, D19_23, D19_22, D19_21, D19_20, D19_19, D19_18, D19_17, D19_16, 
    D19_15, D19_14, D19_13, D19_12, D19_11, D19_10, D19_9, D19_8, D19_7, D19_6, 
    D19_5, D19_4, D19_3, D19_2, D19_1, D19_0, D20_31, D20_30, D20_29, D20_28, 
    D20_27, D20_26, D20_25, D20_24, D20_23, D20_22, D20_21, D20_20, D20_19, 
    D20_18, D20_17, D20_16, D20_15, D20_14, D20_13, D20_12, D20_11, D20_10, 
    D20_9, D20_8, D20_7, D20_6, D20_5, D20_4, D20_3, D20_2, D20_1, D20_0, 
    D21_31, D21_30, D21_29, D21_28, D21_27, D21_26, D21_25, D21_24, D21_23, 
    D21_22, D21_21, D21_20, D21_19, D21_18, D21_17, D21_16, D21_15, D21_14, 
    D21_13, D21_12, D21_11, D21_10, D21_9, D21_8, D21_7, D21_6, D21_5, D21_4, 
    D21_3, D21_2, D21_1, D21_0, D22_31, D22_30, D22_29, D22_28, D22_27, D22_26, 
    D22_25, D22_24, D22_23, D22_22, D22_21, D22_20, D22_19, D22_18, D22_17, 
    D22_16, D22_15, D22_14, D22_13, D22_12, D22_11, D22_10, D22_9, D22_8, 
    D22_7, D22_6, D22_5, D22_4, D22_3, D22_2, D22_1, D22_0, D23_31, D23_30, 
    D23_29, D23_28, D23_27, D23_26, D23_25, D23_24, D23_23, D23_22, D23_21, 
    D23_20, D23_19, D23_18, D23_17, D23_16, D23_15, D23_14, D23_13, D23_12, 
    D23_11, D23_10, D23_9, D23_8, D23_7, D23_6, D23_5, D23_4, D23_3, D23_2, 
    D23_1, D23_0, D24_31, D24_30, D24_29, D24_28, D24_27, D24_26, D24_25, 
    D24_24, D24_23, D24_22, D24_21, D24_20, D24_19, D24_18, D24_17, D24_16, 
    D24_15, D24_14, D24_13, D24_12, D24_11, D24_10, D24_9, D24_8, D24_7, D24_6, 
    D24_5, D24_4, D24_3, D24_2, D24_1, D24_0, D25_31, D25_30, D25_29, D25_28, 
    D25_27, D25_26, D25_25, D25_24, D25_23, D25_22, D25_21, D25_20, D25_19, 
    D25_18, D25_17, D25_16, D25_15, D25_14, D25_13, D25_12, D25_11, D25_10, 
    D25_9, D25_8, D25_7, D25_6, D25_5, D25_4, D25_3, D25_2, D25_1, D25_0, 
    D26_31, D26_30, D26_29, D26_28, D26_27, D26_26, D26_25, D26_24, D26_23, 
    D26_22, D26_21, D26_20, D26_19, D26_18, D26_17, D26_16, D26_15, D26_14, 
    D26_13, D26_12, D26_11, D26_10, D26_9, D26_8, D26_7, D26_6, D26_5, D26_4, 
    D26_3, D26_2, D26_1, D26_0, D27_31, D27_30, D27_29, D27_28, D27_27, D27_26, 
    D27_25, D27_24, D27_23, D27_22, D27_21, D27_20, D27_19, D27_18, D27_17, 
    D27_16, D27_15, D27_14, D27_13, D27_12, D27_11, D27_10, D27_9, D27_8, 
    D27_7, D27_6, D27_5, D27_4, D27_3, D27_2, D27_1, D27_0, D28_31, D28_30, 
    D28_29, D28_28, D28_27, D28_26, D28_25, D28_24, D28_23, D28_22, D28_21, 
    D28_20, D28_19, D28_18, D28_17, D28_16, D28_15, D28_14, D28_13, D28_12, 
    D28_11, D28_10, D28_9, D28_8, D28_7, D28_6, D28_5, D28_4, D28_3, D28_2, 
    D28_1, D28_0, D29_31, D29_30, D29_29, D29_28, D29_27, D29_26, D29_25, 
    D29_24, D29_23, D29_22, D29_21, D29_20, D29_19, D29_18, D29_17, D29_16, 
    D29_15, D29_14, D29_13, D29_12, D29_11, D29_10, D29_9, D29_8, D29_7, D29_6, 
    D29_5, D29_4, D29_3, D29_2, D29_1, D29_0, D30_31, D30_30, D30_29, D30_28, 
    D30_27, D30_26, D30_25, D30_24, D30_23, D30_22, D30_21, D30_20, D30_19, 
    D30_18, D30_17, D30_16, D30_15, D30_14, D30_13, D30_12, D30_11, D30_10, 
    D30_9, D30_8, D30_7, D30_6, D30_5, D30_4, D30_3, D30_2, D30_1, D30_0, 
    D31_31, D31_30, D31_29, D31_28, D31_27, D31_26, D31_25, D31_24, D31_23, 
    D31_22, D31_21, D31_20, D31_19, D31_18, D31_17, D31_16, D31_15, D31_14, 
    D31_13, D31_12, D31_11, D31_10, D31_9, D31_8, D31_7, D31_6, D31_5, D31_4, 
    D31_3, D31_2, D31_1, D31_0, S0, S1, S2, S3, S4, Z_31, Z_30, Z_29, Z_28, 
    Z_27, Z_26, Z_25, Z_24, Z_23, Z_22, Z_21, Z_20, Z_19, Z_18, Z_17, Z_16, 
    Z_15, Z_14, Z_13, Z_12, Z_11, Z_10, Z_9, Z_8, Z_7, Z_6, Z_5, Z_4, Z_3, Z_2, 
    Z_1, Z_0 );
input  D0_31, D0_30, D0_29, D0_28, D0_27, D0_26, D0_25, D0_24, D0_23, D0_22, 
    D0_21, D0_20, D0_19, D0_18, D0_17, D0_16, D0_15, D0_14, D0_13, D0_12, 
    D0_11, D0_10, D0_9, D0_8, D0_7, D0_6, D0_5, D0_4, D0_3, D0_2, D0_1, D0_0, 
    D1_31, D1_30, D1_29, D1_28, D1_27, D1_26, D1_25, D1_24, D1_23, D1_22, 
    D1_21, D1_20, D1_19, D1_18, D1_17, D1_16, D1_15, D1_14, D1_13, D1_12, 
    D1_11, D1_10, D1_9, D1_8, D1_7, D1_6, D1_5, D1_4, D1_3, D1_2, D1_1, D1_0, 
    D2_31, D2_30, D2_29, D2_28, D2_27, D2_26, D2_25, D2_24, D2_23, D2_22, 
    D2_21, D2_20, D2_19, D2_18, D2_17, D2_16, D2_15, D2_14, D2_13, D2_12, 
    D2_11, D2_10, D2_9, D2_8, D2_7, D2_6, D2_5, D2_4, D2_3, D2_2, D2_1, D2_0, 
    D3_31, D3_30, D3_29, D3_28, D3_27, D3_26, D3_25, D3_24, D3_23, D3_22, 
    D3_21, D3_20, D3_19, D3_18, D3_17, D3_16, D3_15, D3_14, D3_13, D3_12, 
    D3_11, D3_10, D3_9, D3_8, D3_7, D3_6, D3_5, D3_4, D3_3, D3_2, D3_1, D3_0, 
    D4_31, D4_30, D4_29, D4_28, D4_27, D4_26, D4_25, D4_24, D4_23, D4_22, 
    D4_21, D4_20, D4_19, D4_18, D4_17, D4_16, D4_15, D4_14, D4_13, D4_12, 
    D4_11, D4_10, D4_9, D4_8, D4_7, D4_6, D4_5, D4_4, D4_3, D4_2, D4_1, D4_0, 
    D5_31, D5_30, D5_29, D5_28, D5_27, D5_26, D5_25, D5_24, D5_23, D5_22, 
    D5_21, D5_20, D5_19, D5_18, D5_17, D5_16, D5_15, D5_14, D5_13, D5_12, 
    D5_11, D5_10, D5_9, D5_8, D5_7, D5_6, D5_5, D5_4, D5_3, D5_2, D5_1, D5_0, 
    D6_31, D6_30, D6_29, D6_28, D6_27, D6_26, D6_25, D6_24, D6_23, D6_22, 
    D6_21, D6_20, D6_19, D6_18, D6_17, D6_16, D6_15, D6_14, D6_13, D6_12, 
    D6_11, D6_10, D6_9, D6_8, D6_7, D6_6, D6_5, D6_4, D6_3, D6_2, D6_1, D6_0, 
    D7_31, D7_30, D7_29, D7_28, D7_27, D7_26, D7_25, D7_24, D7_23, D7_22, 
    D7_21, D7_20, D7_19, D7_18, D7_17, D7_16, D7_15, D7_14, D7_13, D7_12, 
    D7_11, D7_10, D7_9, D7_8, D7_7, D7_6, D7_5, D7_4, D7_3, D7_2, D7_1, D7_0, 
    D8_31, D8_30, D8_29, D8_28, D8_27, D8_26, D8_25, D8_24, D8_23, D8_22, 
    D8_21, D8_20, D8_19, D8_18, D8_17, D8_16, D8_15, D8_14, D8_13, D8_12, 
    D8_11, D8_10, D8_9, D8_8, D8_7, D8_6, D8_5, D8_4, D8_3, D8_2, D8_1, D8_0, 
    D9_31, D9_30, D9_29, D9_28, D9_27, D9_26, D9_25, D9_24, D9_23, D9_22, 
    D9_21, D9_20, D9_19, D9_18, D9_17, D9_16, D9_15, D9_14, D9_13, D9_12, 
    D9_11, D9_10, D9_9, D9_8, D9_7, D9_6, D9_5, D9_4, D9_3, D9_2, D9_1, D9_0, 
    D10_31, D10_30, D10_29, D10_28, D10_27, D10_26, D10_25, D10_24, D10_23, 
    D10_22, D10_21, D10_20, D10_19, D10_18, D10_17, D10_16, D10_15, D10_14, 
    D10_13, D10_12, D10_11, D10_10, D10_9, D10_8, D10_7, D10_6, D10_5, D10_4, 
    D10_3, D10_2, D10_1, D10_0, D11_31, D11_30, D11_29, D11_28, D11_27, D11_26, 
    D11_25, D11_24, D11_23, D11_22, D11_21, D11_20, D11_19, D11_18, D11_17, 
    D11_16, D11_15, D11_14, D11_13, D11_12, D11_11, D11_10, D11_9, D11_8, 
    D11_7, D11_6, D11_5, D11_4, D11_3, D11_2, D11_1, D11_0, D12_31, D12_30, 
    D12_29, D12_28, D12_27, D12_26, D12_25, D12_24, D12_23, D12_22, D12_21, 
    D12_20, D12_19, D12_18, D12_17, D12_16, D12_15, D12_14, D12_13, D12_12, 
    D12_11, D12_10, D12_9, D12_8, D12_7, D12_6, D12_5, D12_4, D12_3, D12_2, 
    D12_1, D12_0, D13_31, D13_30, D13_29, D13_28, D13_27, D13_26, D13_25, 
    D13_24, D13_23, D13_22, D13_21, D13_20, D13_19, D13_18, D13_17, D13_16, 
    D13_15, D13_14, D13_13, D13_12, D13_11, D13_10, D13_9, D13_8, D13_7, D13_6, 
    D13_5, D13_4, D13_3, D13_2, D13_1, D13_0, D14_31, D14_30, D14_29, D14_28, 
    D14_27, D14_26, D14_25, D14_24, D14_23, D14_22, D14_21, D14_20, D14_19, 
    D14_18, D14_17, D14_16, D14_15, D14_14, D14_13, D14_12, D14_11, D14_10, 
    D14_9, D14_8, D14_7, D14_6, D14_5, D14_4, D14_3, D14_2, D14_1, D14_0, 
    D15_31, D15_30, D15_29, D15_28, D15_27, D15_26, D15_25, D15_24, D15_23, 
    D15_22, D15_21, D15_20, D15_19, D15_18, D15_17, D15_16, D15_15, D15_14, 
    D15_13, D15_12, D15_11, D15_10, D15_9, D15_8, D15_7, D15_6, D15_5, D15_4, 
    D15_3, D15_2, D15_1, D15_0, D16_31, D16_30, D16_29, D16_28, D16_27, D16_26, 
    D16_25, D16_24, D16_23, D16_22, D16_21, D16_20, D16_19, D16_18, D16_17, 
    D16_16, D16_15, D16_14, D16_13, D16_12, D16_11, D16_10, D16_9, D16_8, 
    D16_7, D16_6, D16_5, D16_4, D16_3, D16_2, D16_1, D16_0, D17_31, D17_30, 
    D17_29, D17_28, D17_27, D17_26, D17_25, D17_24, D17_23, D17_22, D17_21, 
    D17_20, D17_19, D17_18, D17_17, D17_16, D17_15, D17_14, D17_13, D17_12, 
    D17_11, D17_10, D17_9, D17_8, D17_7, D17_6, D17_5, D17_4, D17_3, D17_2, 
    D17_1, D17_0, D18_31, D18_30, D18_29, D18_28, D18_27, D18_26, D18_25, 
    D18_24, D18_23, D18_22, D18_21, D18_20, D18_19, D18_18, D18_17, D18_16, 
    D18_15, D18_14, D18_13, D18_12, D18_11, D18_10, D18_9, D18_8, D18_7, D18_6, 
    D18_5, D18_4, D18_3, D18_2, D18_1, D18_0, D19_31, D19_30, D19_29, D19_28, 
    D19_27, D19_26, D19_25, D19_24, D19_23, D19_22, D19_21, D19_20, D19_19, 
    D19_18, D19_17, D19_16, D19_15, D19_14, D19_13, D19_12, D19_11, D19_10, 
    D19_9, D19_8, D19_7, D19_6, D19_5, D19_4, D19_3, D19_2, D19_1, D19_0, 
    D20_31, D20_30, D20_29, D20_28, D20_27, D20_26, D20_25, D20_24, D20_23, 
    D20_22, D20_21, D20_20, D20_19, D20_18, D20_17, D20_16, D20_15, D20_14, 
    D20_13, D20_12, D20_11, D20_10, D20_9, D20_8, D20_7, D20_6, D20_5, D20_4, 
    D20_3, D20_2, D20_1, D20_0, D21_31, D21_30, D21_29, D21_28, D21_27, D21_26, 
    D21_25, D21_24, D21_23, D21_22, D21_21, D21_20, D21_19, D21_18, D21_17, 
    D21_16, D21_15, D21_14, D21_13, D21_12, D21_11, D21_10, D21_9, D21_8, 
    D21_7, D21_6, D21_5, D21_4, D21_3, D21_2, D21_1, D21_0, D22_31, D22_30, 
    D22_29, D22_28, D22_27, D22_26, D22_25, D22_24, D22_23, D22_22, D22_21, 
    D22_20, D22_19, D22_18, D22_17, D22_16, D22_15, D22_14, D22_13, D22_12, 
    D22_11, D22_10, D22_9, D22_8, D22_7, D22_6, D22_5, D22_4, D22_3, D22_2, 
    D22_1, D22_0, D23_31, D23_30, D23_29, D23_28, D23_27, D23_26, D23_25, 
    D23_24, D23_23, D23_22, D23_21, D23_20, D23_19, D23_18, D23_17, D23_16, 
    D23_15, D23_14, D23_13, D23_12, D23_11, D23_10, D23_9, D23_8, D23_7, D23_6, 
    D23_5, D23_4, D23_3, D23_2, D23_1, D23_0, D24_31, D24_30, D24_29, D24_28, 
    D24_27, D24_26, D24_25, D24_24, D24_23, D24_22, D24_21, D24_20, D24_19, 
    D24_18, D24_17, D24_16, D24_15, D24_14, D24_13, D24_12, D24_11, D24_10, 
    D24_9, D24_8, D24_7, D24_6, D24_5, D24_4, D24_3, D24_2, D24_1, D24_0, 
    D25_31, D25_30, D25_29, D25_28, D25_27, D25_26, D25_25, D25_24, D25_23, 
    D25_22, D25_21, D25_20, D25_19, D25_18, D25_17, D25_16, D25_15, D25_14, 
    D25_13, D25_12, D25_11, D25_10, D25_9, D25_8, D25_7, D25_6, D25_5, D25_4, 
    D25_3, D25_2, D25_1, D25_0, D26_31, D26_30, D26_29, D26_28, D26_27, D26_26, 
    D26_25, D26_24, D26_23, D26_22, D26_21, D26_20, D26_19, D26_18, D26_17, 
    D26_16, D26_15, D26_14, D26_13, D26_12, D26_11, D26_10, D26_9, D26_8, 
    D26_7, D26_6, D26_5, D26_4, D26_3, D26_2, D26_1, D26_0, D27_31, D27_30, 
    D27_29, D27_28, D27_27, D27_26, D27_25, D27_24, D27_23, D27_22, D27_21, 
    D27_20, D27_19, D27_18, D27_17, D27_16, D27_15, D27_14, D27_13, D27_12, 
    D27_11, D27_10, D27_9, D27_8, D27_7, D27_6, D27_5, D27_4, D27_3, D27_2, 
    D27_1, D27_0, D28_31, D28_30, D28_29, D28_28, D28_27, D28_26, D28_25, 
    D28_24, D28_23, D28_22, D28_21, D28_20, D28_19, D28_18, D28_17, D28_16, 
    D28_15, D28_14, D28_13, D28_12, D28_11, D28_10, D28_9, D28_8, D28_7, D28_6, 
    D28_5, D28_4, D28_3, D28_2, D28_1, D28_0, D29_31, D29_30, D29_29, D29_28, 
    D29_27, D29_26, D29_25, D29_24, D29_23, D29_22, D29_21, D29_20, D29_19, 
    D29_18, D29_17, D29_16, D29_15, D29_14, D29_13, D29_12, D29_11, D29_10, 
    D29_9, D29_8, D29_7, D29_6, D29_5, D29_4, D29_3, D29_2, D29_1, D29_0, 
    D30_31, D30_30, D30_29, D30_28, D30_27, D30_26, D30_25, D30_24, D30_23, 
    D30_22, D30_21, D30_20, D30_19, D30_18, D30_17, D30_16, D30_15, D30_14, 
    D30_13, D30_12, D30_11, D30_10, D30_9, D30_8, D30_7, D30_6, D30_5, D30_4, 
    D30_3, D30_2, D30_1, D30_0, D31_31, D31_30, D31_29, D31_28, D31_27, D31_26, 
    D31_25, D31_24, D31_23, D31_22, D31_21, D31_20, D31_19, D31_18, D31_17, 
    D31_16, D31_15, D31_14, D31_13, D31_12, D31_11, D31_10, D31_9, D31_8, 
    D31_7, D31_6, D31_5, D31_4, D31_3, D31_2, D31_1, D31_0, S0, S1, S2, S3, S4;
output Z_31, Z_30, Z_29, Z_28, Z_27, Z_26, Z_25, Z_24, Z_23, Z_22, Z_21, Z_20, 
    Z_19, Z_18, Z_17, Z_16, Z_15, Z_14, Z_13, Z_12, Z_11, Z_10, Z_9, Z_8, Z_7, 
    Z_6, Z_5, Z_4, Z_3, Z_2, Z_1, Z_0;
    wire n342, n18, n40, n299, n8, n37, n249, n22, n34, n185, n15, n32, n121, 
        n11, n28, n153, n20, n30, n89, n19, n26, n350, n24, n41, n286, n23, 
        n318, n39, n254, n35, n190, n21, n33, n331, n126, n29, n158, n31, n94, 
        n27, n344, n7, n280, n36, n312, n38, n248, n16, n184, n120, n152, n267, 
        n9, n88, n13, n349, n285, n317, n253, n189, n125, n14, n157, n93, n358, 
        n203, n294, n326, n262, n198, n10, n134, n166, n102, n340, n276, n308, 
        n139, n244, n180, n116, n148, n84, n339, n275, n307, n17, n243, n179, 
        n171, n115, n147, n83, n12, n362, n298, n330, n266, n3, n202, n138, 
        n107, n170, n106, n74, n5, n353, n25, n289, n321, n257, n193, n129, 
        n161, n352, n97, n347, n283, n315, n251, n187, n123, n155, n91, n346, 
        n288, n282, n314, n250, n218, n4, n186, n122, n154, n90, n58, n355, 
        n320, n291, n323, n259, n195, n131, n163, n99, n337, n273, n305, n278, 
        n256, n241, n177, n113, n145, n81, n357, n293, n325, n261, n197, n192, 
        n133, n165, n101, n348, n284, n316, n252, n188, n124, n156, n128, n92, 
        n335, n271, n303, n239, n175, n111, n143, n79, n43, n160, n360, n296, 
        n328, n264, n232, n200, n136, n168, n104, n72, n96, n361, n297, n329, 
        n265, n233, n201, n137, n169, n105, n73, n343, n295, n135, n167, n279, 
        n103, n332, n268, n300, n236, n311, n172, n108, n140, n76, n54, n214, 
        n75, n235, n247, n64, n224, n55, n215, n45, n205, n66, n226, n50, n210, 
        n63, n223, n53, n213, n48, n208, n68, n228, n57, n217, n183, n62, n222, 
        n56, n216, n61, n221, n70, n230, n52, n212, n51, n211, n234, n65, n225, 
        n59, n219, n310, n119, n67, n227, n49, n209, n69, n229, n60, n220, n47, 
        n207, n44, n204, n2, n1, n151, n87, n333, n42, n46, n206, n71, n231, 
        n77, n141, n109, n173, n1425, n78, n142, n110, n174, n80, n144, n112, 
        n176, n269, n82, n146, n114, n178, n85, n149, n117, n181, n86, n150, 
        n118, n182, n301, n95, n159, n127, n191, n98, n162, n130, n194, n100, 
        n164, n132, n196, n237, n199, n238, n302, n270, n334, n240, n304, n272, 
        n336, n242, n306, n274, n338, n245, n309, n277, n341, n246, n313, n281, 
        n345, n255, n319, n287, n351, n258, n322, n290, n354, n260, n324, n292, 
        n356, n263, n327, n359, n363;
    mux4_1 U1 ( .x(n342), .d0(D7_10), .d1(D15_10), .d2(D23_10), .d3(D31_10), 
        .sl0(n18), .sl1(n40) );
    mux4_1 U10 ( .x(n299), .d0(D5_31), .d1(D13_31), .d2(D21_31), .d3(D29_31), 
        .sl0(n8), .sl1(n37) );
    mux4_1 U100 ( .x(n249), .d0(D1_13), .d1(D9_13), .d2(D17_13), .d3(D25_13), 
        .sl0(n22), .sl1(n34) );
    mux4_1 U101 ( .x(n185), .d0(D6_13), .d1(D14_13), .d2(D22_13), .d3(D30_13), 
        .sl0(n15), .sl1(n32) );
    mux4_1 U102 ( .x(n121), .d0(D4_13), .d1(D12_13), .d2(D20_13), .d3(D28_13), 
        .sl0(n11), .sl1(n28) );
    mux4_1 U103 ( .x(n153), .d0(D2_13), .d1(D10_13), .d2(D18_13), .d3(D26_13), 
        .sl0(n20), .sl1(n30) );
    mux4_1 U104 ( .x(n89), .d0(D0_13), .d1(D8_13), .d2(D16_13), .d3(D24_13), 
        .sl0(n19), .sl1(n26) );
    mux4_1 U105 ( .x(n350), .d0(D7_18), .d1(D15_18), .d2(D23_18), .d3(D31_18), 
        .sl0(n24), .sl1(n41) );
    mux4_1 U106 ( .x(n286), .d0(D5_18), .d1(D13_18), .d2(D21_18), .d3(D29_18), 
        .sl0(n23), .sl1(n37) );
    mux4_1 U107 ( .x(n318), .d0(D3_18), .d1(D11_18), .d2(D19_18), .d3(D27_18), 
        .sl0(n18), .sl1(n39) );
    mux4_1 U108 ( .x(n254), .d0(D1_18), .d1(D9_18), .d2(D17_18), .d3(D25_18), 
        .sl0(n22), .sl1(n35) );
    mux4_1 U109 ( .x(n190), .d0(D6_18), .d1(D14_18), .d2(D22_18), .d3(D30_18), 
        .sl0(n21), .sl1(n33) );
    mux4_1 U11 ( .x(n331), .d0(D3_31), .d1(D11_31), .d2(D19_31), .d3(D27_31), 
        .sl0(n18), .sl1(n39) );
    mux4_1 U110 ( .x(n126), .d0(D4_18), .d1(D12_18), .d2(D20_18), .d3(D28_18), 
        .sl0(n20), .sl1(n29) );
    mux4_1 U111 ( .x(n158), .d0(D2_18), .d1(D10_18), .d2(D18_18), .d3(D26_18), 
        .sl0(n11), .sl1(n31) );
    mux4_1 U112 ( .x(n94), .d0(D0_18), .d1(D8_18), .d2(D16_18), .d3(D24_18), 
        .sl0(n19), .sl1(n27) );
    mux4_1 U113 ( .x(n344), .d0(D7_12), .d1(D15_12), .d2(D23_12), .d3(D31_12), 
        .sl0(n7), .sl1(n40) );
    mux4_1 U114 ( .x(n280), .d0(D5_12), .d1(D13_12), .d2(D21_12), .d3(D29_12), 
        .sl0(n8), .sl1(n36) );
    mux4_1 U115 ( .x(n312), .d0(D3_12), .d1(D11_12), .d2(D19_12), .d3(D27_12), 
        .sl0(n8), .sl1(n38) );
    mux4_1 U116 ( .x(n248), .d0(D1_12), .d1(D9_12), .d2(D17_12), .d3(D25_12), 
        .sl0(n16), .sl1(n34) );
    mux4_1 U117 ( .x(n184), .d0(D6_12), .d1(D14_12), .d2(D22_12), .d3(D30_12), 
        .sl0(n15), .sl1(n32) );
    mux4_1 U118 ( .x(n120), .d0(D4_12), .d1(D12_12), .d2(D20_12), .d3(D28_12), 
        .sl0(n20), .sl1(n28) );
    mux4_1 U119 ( .x(n152), .d0(D2_12), .d1(D10_12), .d2(D18_12), .d3(D26_12), 
        .sl0(n20), .sl1(n30) );
    mux4_1 U12 ( .x(n267), .d0(D1_31), .d1(D9_31), .d2(D17_31), .d3(D25_31), 
        .sl0(n9), .sl1(n35) );
    mux4_1 U120 ( .x(n88), .d0(D0_12), .d1(D8_12), .d2(D16_12), .d3(D24_12), 
        .sl0(n13), .sl1(n26) );
    mux4_1 U121 ( .x(n349), .d0(D7_17), .d1(D15_17), .d2(D23_17), .d3(D31_17), 
        .sl0(n18), .sl1(n41) );
    mux4_1 U122 ( .x(n285), .d0(D5_17), .d1(D13_17), .d2(D21_17), .d3(D29_17), 
        .sl0(n8), .sl1(n37) );
    mux4_1 U123 ( .x(n317), .d0(D3_17), .d1(D11_17), .d2(D19_17), .d3(D27_17), 
        .sl0(n8), .sl1(n39) );
    mux4_1 U124 ( .x(n253), .d0(D1_17), .d1(D9_17), .d2(D17_17), .d3(D25_17), 
        .sl0(n16), .sl1(n35) );
    mux4_1 U125 ( .x(n189), .d0(D6_17), .d1(D14_17), .d2(D22_17), .d3(D30_17), 
        .sl0(n15), .sl1(n33) );
    mux4_1 U126 ( .x(n125), .d0(D4_17), .d1(D12_17), .d2(D20_17), .d3(D28_17), 
        .sl0(n14), .sl1(n29) );
    mux4_1 U127 ( .x(n157), .d0(D2_17), .d1(D10_17), .d2(D18_17), .d3(D26_17), 
        .sl0(n11), .sl1(n31) );
    mux4_1 U128 ( .x(n93), .d0(D0_17), .d1(D8_17), .d2(D16_17), .d3(D24_17), 
        .sl0(n13), .sl1(n27) );
    mux4_1 U129 ( .x(n358), .d0(D7_26), .d1(D15_26), .d2(D23_26), .d3(D31_26), 
        .sl0(n7), .sl1(n41) );
    mux4_1 U13 ( .x(n203), .d0(D6_31), .d1(D14_31), .d2(D22_31), .d3(D30_31), 
        .sl0(n16), .sl1(n33) );
    mux4_1 U130 ( .x(n294), .d0(D5_26), .d1(D13_26), .d2(D21_26), .d3(D29_26), 
        .sl0(n8), .sl1(n37) );
    mux4_1 U131 ( .x(n326), .d0(D3_26), .d1(D11_26), .d2(D19_26), .d3(D27_26), 
        .sl0(n18), .sl1(n39) );
    mux4_1 U132 ( .x(n262), .d0(D1_26), .d1(D9_26), .d2(D17_26), .d3(D25_26), 
        .sl0(n16), .sl1(n35) );
    mux4_1 U133 ( .x(n198), .d0(D6_26), .d1(D14_26), .d2(D22_26), .d3(D30_26), 
        .sl0(n10), .sl1(n33) );
    mux4_1 U134 ( .x(n134), .d0(D4_26), .d1(D12_26), .d2(D20_26), .d3(D28_26), 
        .sl0(n14), .sl1(n29) );
    mux4_1 U135 ( .x(n166), .d0(D2_26), .d1(D10_26), .d2(D18_26), .d3(D26_26), 
        .sl0(n21), .sl1(n31) );
    mux4_1 U136 ( .x(n102), .d0(D0_26), .d1(D8_26), .d2(D16_26), .d3(D24_26), 
        .sl0(n13), .sl1(n27) );
    mux4_1 U137 ( .x(n340), .d0(D7_8), .d1(D15_8), .d2(D23_8), .d3(D31_8), 
        .sl0(n24), .sl1(n40) );
    mux4_1 U138 ( .x(n276), .d0(D5_8), .d1(D13_8), .d2(D21_8), .d3(D29_8), 
        .sl0(n23), .sl1(n36) );
    mux4_1 U139 ( .x(n308), .d0(D3_8), .d1(D11_8), .d2(D19_8), .d3(D27_8), 
        .sl0(n8), .sl1(n38) );
    mux4_1 U14 ( .x(n139), .d0(D4_31), .d1(D12_31), .d2(D20_31), .d3(D28_31), 
        .sl0(n14), .sl1(n29) );
    mux4_1 U140 ( .x(n244), .d0(D1_8), .d1(D9_8), .d2(D17_8), .d3(D25_8), 
        .sl0(n16), .sl1(n34) );
    mux4_1 U141 ( .x(n180), .d0(D6_8), .d1(D14_8), .d2(D22_8), .d3(D30_8), 
        .sl0(n21), .sl1(n32) );
    mux4_1 U142 ( .x(n116), .d0(D4_8), .d1(D12_8), .d2(D20_8), .d3(D28_8), 
        .sl0(n20), .sl1(n28) );
    mux4_1 U143 ( .x(n148), .d0(D2_8), .d1(D10_8), .d2(D18_8), .d3(D26_8), 
        .sl0(n11), .sl1(n30) );
    mux4_1 U144 ( .x(n84), .d0(D0_8), .d1(D8_8), .d2(D16_8), .d3(D24_8), .sl0(
        n19), .sl1(n26) );
    mux4_1 U145 ( .x(n339), .d0(D7_7), .d1(D15_7), .d2(D23_7), .d3(D31_7), 
        .sl0(n18), .sl1(n40) );
    mux4_1 U146 ( .x(n275), .d0(D5_7), .d1(D13_7), .d2(D21_7), .d3(D29_7), 
        .sl0(n16), .sl1(n36) );
    mux4_1 U147 ( .x(n307), .d0(D3_7), .d1(D11_7), .d2(D19_7), .d3(D27_7), 
        .sl0(n17), .sl1(n38) );
    mux4_1 U148 ( .x(n243), .d0(D1_7), .d1(D9_7), .d2(D17_7), .d3(D25_7), 
        .sl0(n16), .sl1(n34) );
    mux4_1 U149 ( .x(n179), .d0(D6_7), .d1(D14_7), .d2(D22_7), .d3(D30_7), 
        .sl0(n15), .sl1(n32) );
    mux4_1 U15 ( .x(n171), .d0(D2_31), .d1(D10_31), .d2(D18_31), .d3(D26_31), 
        .sl0(n15), .sl1(n31) );
    mux4_1 U150 ( .x(n115), .d0(D4_7), .d1(D12_7), .d2(D20_7), .d3(D28_7), 
        .sl0(n14), .sl1(n28) );
    mux4_1 U151 ( .x(n147), .d0(D2_7), .d1(D10_7), .d2(D18_7), .d3(D26_7), 
        .sl0(n20), .sl1(n30) );
    mux4_1 U152 ( .x(n83), .d0(D0_7), .d1(D8_7), .d2(D16_7), .d3(D24_7), .sl0(
        n12), .sl1(n26) );
    mux4_1 U153 ( .x(n362), .d0(D7_30), .d1(D15_30), .d2(D23_30), .d3(D31_30), 
        .sl0(n19), .sl1(n41) );
    mux4_1 U154 ( .x(n298), .d0(D5_30), .d1(D13_30), .d2(D21_30), .d3(D29_30), 
        .sl0(n23), .sl1(n37) );
    mux4_1 U155 ( .x(n330), .d0(D3_30), .d1(D11_30), .d2(D19_30), .d3(D27_30), 
        .sl0(n7), .sl1(n39) );
    mux4_1 U156 ( .x(n266), .d0(D1_30), .d1(D9_30), .d2(D17_30), .d3(D25_30), 
        .sl0(n16), .sl1(n35) );
    buf_3 U157 ( .x(n3), .a(S1) );
    mux4_1 U158 ( .x(n202), .d0(D6_30), .d1(D14_30), .d2(D22_30), .d3(D30_30), 
        .sl0(n22), .sl1(n33) );
    mux4_1 U159 ( .x(n138), .d0(D4_30), .d1(D12_30), .d2(D20_30), .d3(D28_30), 
        .sl0(n11), .sl1(n29) );
    mux4_1 U16 ( .x(n107), .d0(D0_31), .d1(D8_31), .d2(D16_31), .d3(D24_31), 
        .sl0(n12), .sl1(n27) );
    mux4_1 U160 ( .x(n170), .d0(D2_30), .d1(D10_30), .d2(D18_30), .d3(D26_30), 
        .sl0(n10), .sl1(n31) );
    mux4_1 U161 ( .x(n106), .d0(D0_30), .d1(D8_30), .d2(D16_30), .d3(D24_30), 
        .sl0(n19), .sl1(n27) );
    mux4_2 U162 ( .x(n74), .d0(n106), .d1(n170), .d2(n138), .d3(n202), .sl0(n3
        ), .sl1(n5) );
    mux4_1 U163 ( .x(n353), .d0(D7_21), .d1(D15_21), .d2(D23_21), .d3(D31_21), 
        .sl0(n25), .sl1(n41) );
    mux4_1 U164 ( .x(n289), .d0(D5_21), .d1(D13_21), .d2(D21_21), .d3(D29_21), 
        .sl0(n8), .sl1(n37) );
    mux4_1 U165 ( .x(n321), .d0(D3_21), .d1(D11_21), .d2(D19_21), .d3(D27_21), 
        .sl0(n18), .sl1(n39) );
    mux4_1 U166 ( .x(n257), .d0(D1_21), .d1(D9_21), .d2(D17_21), .d3(D25_21), 
        .sl0(n22), .sl1(n35) );
    mux4_1 U167 ( .x(n193), .d0(D6_21), .d1(D14_21), .d2(D22_21), .d3(D30_21), 
        .sl0(n10), .sl1(n33) );
    mux4_1 U168 ( .x(n129), .d0(D4_21), .d1(D12_21), .d2(D20_21), .d3(D28_21), 
        .sl0(n20), .sl1(n29) );
    mux4_1 U169 ( .x(n161), .d0(D2_21), .d1(D10_21), .d2(D18_21), .d3(D26_21), 
        .sl0(n21), .sl1(n31) );
    mux4_1 U17 ( .x(n352), .d0(D7_20), .d1(D15_20), .d2(D23_20), .d3(D31_20), 
        .sl0(n18), .sl1(n41) );
    mux4_1 U170 ( .x(n97), .d0(D0_21), .d1(D8_21), .d2(D16_21), .d3(D24_21), 
        .sl0(n19), .sl1(n27) );
    mux4_1 U171 ( .x(n347), .d0(D7_15), .d1(D15_15), .d2(D23_15), .d3(D31_15), 
        .sl0(n24), .sl1(n40) );
    mux4_1 U172 ( .x(n283), .d0(D5_15), .d1(D13_15), .d2(D21_15), .d3(D29_15), 
        .sl0(n23), .sl1(n36) );
    mux4_1 U173 ( .x(n315), .d0(D3_15), .d1(D11_15), .d2(D19_15), .d3(D27_15), 
        .sl0(n24), .sl1(n38) );
    mux4_1 U174 ( .x(n251), .d0(D1_15), .d1(D9_15), .d2(D17_15), .d3(D25_15), 
        .sl0(n22), .sl1(n34) );
    mux4_1 U175 ( .x(n187), .d0(D6_15), .d1(D14_15), .d2(D22_15), .d3(D30_15), 
        .sl0(n15), .sl1(n32) );
    mux4_1 U176 ( .x(n123), .d0(D4_15), .d1(D12_15), .d2(D20_15), .d3(D28_15), 
        .sl0(n20), .sl1(n28) );
    mux4_1 U177 ( .x(n155), .d0(D2_15), .d1(D10_15), .d2(D18_15), .d3(D26_15), 
        .sl0(n15), .sl1(n30) );
    mux4_1 U178 ( .x(n91), .d0(D0_15), .d1(D8_15), .d2(D16_15), .d3(D24_15), 
        .sl0(n13), .sl1(n26) );
    mux4_1 U179 ( .x(n346), .d0(D7_14), .d1(D15_14), .d2(D23_14), .d3(D31_14), 
        .sl0(n7), .sl1(n40) );
    mux4_1 U18 ( .x(n288), .d0(D5_20), .d1(D13_20), .d2(D21_20), .d3(D29_20), 
        .sl0(n17), .sl1(n37) );
    mux4_1 U180 ( .x(n282), .d0(D5_14), .d1(D13_14), .d2(D21_14), .d3(D29_14), 
        .sl0(n17), .sl1(n36) );
    mux4_1 U181 ( .x(n314), .d0(D3_14), .d1(D11_14), .d2(D19_14), .d3(D27_14), 
        .sl0(n17), .sl1(n38) );
    mux4_1 U182 ( .x(n250), .d0(D1_14), .d1(D9_14), .d2(D17_14), .d3(D25_14), 
        .sl0(n9), .sl1(n34) );
    mux4_2 U183 ( .x(n218), .d0(n250), .d1(n314), .d2(n282), .d3(n346), .sl0(
        n4), .sl1(n5) );
    mux4_1 U184 ( .x(n186), .d0(D6_14), .d1(D14_14), .d2(D22_14), .d3(D30_14), 
        .sl0(n15), .sl1(n32) );
    mux4_1 U185 ( .x(n122), .d0(D4_14), .d1(D12_14), .d2(D20_14), .d3(D28_14), 
        .sl0(n14), .sl1(n28) );
    mux4_1 U186 ( .x(n154), .d0(D2_14), .d1(D10_14), .d2(D18_14), .d3(D26_14), 
        .sl0(n11), .sl1(n30) );
    mux4_1 U187 ( .x(n90), .d0(D0_14), .d1(D8_14), .d2(D16_14), .d3(D24_14), 
        .sl0(n12), .sl1(n26) );
    mux4_2 U188 ( .x(n58), .d0(n90), .d1(n154), .d2(n122), .d3(n186), .sl0(n4), 
        .sl1(n5) );
    mux4_1 U189 ( .x(n355), .d0(D7_23), .d1(D15_23), .d2(D23_23), .d3(D31_23), 
        .sl0(n18), .sl1(n41) );
    mux4_1 U19 ( .x(n320), .d0(D3_20), .d1(D11_20), .d2(D19_20), .d3(D27_20), 
        .sl0(n8), .sl1(n39) );
    mux4_1 U190 ( .x(n291), .d0(D5_23), .d1(D13_23), .d2(D21_23), .d3(D29_23), 
        .sl0(n17), .sl1(n37) );
    mux4_1 U191 ( .x(n323), .d0(D3_23), .d1(D11_23), .d2(D19_23), .d3(D27_23), 
        .sl0(n7), .sl1(n39) );
    mux4_1 U192 ( .x(n259), .d0(D1_23), .d1(D9_23), .d2(D17_23), .d3(D25_23), 
        .sl0(n22), .sl1(n35) );
    mux4_1 U193 ( .x(n195), .d0(D6_23), .d1(D14_23), .d2(D22_23), .d3(D30_23), 
        .sl0(n21), .sl1(n33) );
    mux4_1 U194 ( .x(n131), .d0(D4_23), .d1(D12_23), .d2(D20_23), .d3(D28_23), 
        .sl0(n14), .sl1(n29) );
    mux4_1 U195 ( .x(n163), .d0(D2_23), .d1(D10_23), .d2(D18_23), .d3(D26_23), 
        .sl0(n15), .sl1(n31) );
    mux4_1 U196 ( .x(n99), .d0(D0_23), .d1(D8_23), .d2(D16_23), .d3(D24_23), 
        .sl0(n19), .sl1(n27) );
    mux4_1 U197 ( .x(n337), .d0(D7_5), .d1(D15_5), .d2(D23_5), .d3(D31_5), 
        .sl0(n7), .sl1(n40) );
    mux4_1 U198 ( .x(n273), .d0(D5_5), .d1(D13_5), .d2(D21_5), .d3(D29_5), 
        .sl0(n23), .sl1(n36) );
    mux4_1 U199 ( .x(n305), .d0(D3_5), .d1(D11_5), .d2(D19_5), .d3(D27_5), 
        .sl0(n8), .sl1(n38) );
    mux4_1 U2 ( .x(n278), .d0(D5_10), .d1(D13_10), .d2(D21_10), .d3(D29_10), 
        .sl0(n17), .sl1(n36) );
    mux4_1 U20 ( .x(n256), .d0(D1_20), .d1(D9_20), .d2(D17_20), .d3(D25_20), 
        .sl0(n16), .sl1(n35) );
    mux4_1 U200 ( .x(n241), .d0(D1_5), .d1(D9_5), .d2(D17_5), .d3(D25_5), 
        .sl0(n22), .sl1(n34) );
    mux4_1 U201 ( .x(n177), .d0(D6_5), .d1(D14_5), .d2(D22_5), .d3(D30_5), 
        .sl0(n21), .sl1(n32) );
    mux4_1 U202 ( .x(n113), .d0(D4_5), .d1(D12_5), .d2(D20_5), .d3(D28_5), 
        .sl0(n12), .sl1(n28) );
    mux4_1 U203 ( .x(n145), .d0(D2_5), .d1(D10_5), .d2(D18_5), .d3(D26_5), 
        .sl0(n11), .sl1(n30) );
    mux4_1 U204 ( .x(n81), .d0(D0_5), .d1(D8_5), .d2(D16_5), .d3(D24_5), .sl0(
        n19), .sl1(n26) );
    mux4_1 U205 ( .x(n357), .d0(D7_25), .d1(D15_25), .d2(D23_25), .d3(D31_25), 
        .sl0(n7), .sl1(n41) );
    mux4_1 U206 ( .x(n293), .d0(D5_25), .d1(D13_25), .d2(D21_25), .d3(D29_25), 
        .sl0(n17), .sl1(n37) );
    mux4_1 U207 ( .x(n325), .d0(D3_25), .d1(D11_25), .d2(D19_25), .d3(D27_25), 
        .sl0(n7), .sl1(n39) );
    mux4_1 U208 ( .x(n261), .d0(D1_25), .d1(D9_25), .d2(D17_25), .d3(D25_25), 
        .sl0(n22), .sl1(n35) );
    mux4_1 U209 ( .x(n197), .d0(D6_25), .d1(D14_25), .d2(D22_25), .d3(D30_25), 
        .sl0(n10), .sl1(n33) );
    mux4_1 U21 ( .x(n192), .d0(D6_20), .d1(D14_20), .d2(D22_20), .d3(D30_20), 
        .sl0(n21), .sl1(n33) );
    mux4_1 U210 ( .x(n133), .d0(D4_25), .d1(D12_25), .d2(D20_25), .d3(D28_25), 
        .sl0(n20), .sl1(n29) );
    mux4_1 U211 ( .x(n165), .d0(D2_25), .d1(D10_25), .d2(D18_25), .d3(D26_25), 
        .sl0(n15), .sl1(n31) );
    mux4_1 U212 ( .x(n101), .d0(D0_25), .d1(D8_25), .d2(D16_25), .d3(D24_25), 
        .sl0(n12), .sl1(n27) );
    mux4_1 U213 ( .x(n348), .d0(D7_16), .d1(D15_16), .d2(D23_16), .d3(D31_16), 
        .sl0(n7), .sl1(n41) );
    mux4_1 U214 ( .x(n284), .d0(D5_16), .d1(D13_16), .d2(D21_16), .d3(D29_16), 
        .sl0(n17), .sl1(n37) );
    mux4_1 U215 ( .x(n316), .d0(D3_16), .d1(D11_16), .d2(D19_16), .d3(D27_16), 
        .sl0(n24), .sl1(n39) );
    mux4_1 U216 ( .x(n252), .d0(D1_16), .d1(D9_16), .d2(D17_16), .d3(D25_16), 
        .sl0(n9), .sl1(n35) );
    mux4_1 U217 ( .x(n188), .d0(D6_16), .d1(D14_16), .d2(D22_16), .d3(D30_16), 
        .sl0(n21), .sl1(n33) );
    mux4_1 U218 ( .x(n124), .d0(D4_16), .d1(D12_16), .d2(D20_16), .d3(D28_16), 
        .sl0(n11), .sl1(n29) );
    mux4_1 U219 ( .x(n156), .d0(D2_16), .d1(D10_16), .d2(D18_16), .d3(D26_16), 
        .sl0(n15), .sl1(n31) );
    mux4_1 U22 ( .x(n128), .d0(D4_20), .d1(D12_20), .d2(D20_20), .d3(D28_20), 
        .sl0(n14), .sl1(n29) );
    mux4_1 U220 ( .x(n92), .d0(D0_16), .d1(D8_16), .d2(D16_16), .d3(D24_16), 
        .sl0(n13), .sl1(n27) );
    mux4_1 U221 ( .x(n335), .d0(D7_3), .d1(D15_3), .d2(D23_3), .d3(D31_3), 
        .sl0(n24), .sl1(n40) );
    mux4_1 U222 ( .x(n271), .d0(D5_3), .d1(D13_3), .d2(D21_3), .d3(D29_3), 
        .sl0(n23), .sl1(n36) );
    mux4_1 U223 ( .x(n303), .d0(D3_3), .d1(D11_3), .d2(D19_3), .d3(D27_3), 
        .sl0(n23), .sl1(n38) );
    mux4_1 U224 ( .x(n239), .d0(D1_3), .d1(D9_3), .d2(D17_3), .d3(D25_3), 
        .sl0(n9), .sl1(n34) );
    mux4_1 U225 ( .x(n175), .d0(D6_3), .d1(D14_3), .d2(D22_3), .d3(D30_3), 
        .sl0(n10), .sl1(n32) );
    mux4_1 U226 ( .x(n111), .d0(D4_3), .d1(D12_3), .d2(D20_3), .d3(D28_3), 
        .sl0(n19), .sl1(n28) );
    mux4_1 U227 ( .x(n143), .d0(D2_3), .d1(D10_3), .d2(D18_3), .d3(D26_3), 
        .sl0(n14), .sl1(n30) );
    mux4_1 U228 ( .x(n79), .d0(D0_3), .d1(D8_3), .d2(D16_3), .d3(D24_3), .sl0(
        n13), .sl1(n26) );
    buf_3 U229 ( .x(n25), .a(n43) );
    mux4_1 U23 ( .x(n160), .d0(D2_20), .d1(D10_20), .d2(D18_20), .d3(D26_20), 
        .sl0(n11), .sl1(n31) );
    mux4_1 U230 ( .x(n360), .d0(D7_28), .d1(D15_28), .d2(D23_28), .d3(D31_28), 
        .sl0(n25), .sl1(n41) );
    mux4_1 U231 ( .x(n296), .d0(D5_28), .d1(D13_28), .d2(D21_28), .d3(D29_28), 
        .sl0(n17), .sl1(n37) );
    mux4_1 U232 ( .x(n328), .d0(D3_28), .d1(D11_28), .d2(D19_28), .d3(D27_28), 
        .sl0(n24), .sl1(n39) );
    mux4_1 U233 ( .x(n264), .d0(D1_28), .d1(D9_28), .d2(D17_28), .d3(D25_28), 
        .sl0(n9), .sl1(n35) );
    mux4_2 U234 ( .x(n232), .d0(n264), .d1(n328), .d2(n296), .d3(n360), .sl0(
        n3), .sl1(n5) );
    mux4_1 U235 ( .x(n200), .d0(D6_28), .d1(D14_28), .d2(D22_28), .d3(D30_28), 
        .sl0(n16), .sl1(n33) );
    mux4_1 U236 ( .x(n136), .d0(D4_28), .d1(D12_28), .d2(D20_28), .d3(D28_28), 
        .sl0(n20), .sl1(n29) );
    mux4_1 U237 ( .x(n168), .d0(D2_28), .d1(D10_28), .d2(D18_28), .d3(D26_28), 
        .sl0(n21), .sl1(n31) );
    mux4_1 U238 ( .x(n104), .d0(D0_28), .d1(D8_28), .d2(D16_28), .d3(D24_28), 
        .sl0(n13), .sl1(n27) );
    mux4_2 U239 ( .x(n72), .d0(n104), .d1(n168), .d2(n136), .d3(n200), .sl0(n3
        ), .sl1(n5) );
    mux4_1 U24 ( .x(n96), .d0(D0_20), .d1(D8_20), .d2(D16_20), .d3(D24_20), 
        .sl0(n12), .sl1(n27) );
    mux4_1 U240 ( .x(n361), .d0(D7_29), .d1(D15_29), .d2(D23_29), .d3(D31_29), 
        .sl0(n25), .sl1(n41) );
    mux4_1 U241 ( .x(n297), .d0(D5_29), .d1(D13_29), .d2(D21_29), .d3(D29_29), 
        .sl0(n23), .sl1(n37) );
    mux4_1 U242 ( .x(n329), .d0(D3_29), .d1(D11_29), .d2(D19_29), .d3(D27_29), 
        .sl0(n24), .sl1(n39) );
    mux4_1 U243 ( .x(n265), .d0(D1_29), .d1(D9_29), .d2(D17_29), .d3(D25_29), 
        .sl0(n22), .sl1(n35) );
    mux4_2 U244 ( .x(n233), .d0(n265), .d1(n329), .d2(n297), .d3(n361), .sl0(
        n3), .sl1(n5) );
    mux4_1 U245 ( .x(n201), .d0(D6_29), .d1(D14_29), .d2(D22_29), .d3(D30_29), 
        .sl0(n22), .sl1(n33) );
    mux4_1 U246 ( .x(n137), .d0(D4_29), .d1(D12_29), .d2(D20_29), .d3(D28_29), 
        .sl0(n11), .sl1(n29) );
    mux4_1 U247 ( .x(n169), .d0(D2_29), .d1(D10_29), .d2(D18_29), .d3(D26_29), 
        .sl0(n10), .sl1(n31) );
    mux4_1 U248 ( .x(n105), .d0(D0_29), .d1(D8_29), .d2(D16_29), .d3(D24_29), 
        .sl0(n19), .sl1(n27) );
    mux4_2 U249 ( .x(n73), .d0(n105), .d1(n169), .d2(n137), .d3(n201), .sl0(n3
        ), .sl1(n5) );
    mux4_1 U25 ( .x(n343), .d0(D7_11), .d1(D15_11), .d2(D23_11), .d3(D31_11), 
        .sl0(n7), .sl1(n40) );
    buf_3 U250 ( .x(n41), .a(S4) );
    buf_3 U251 ( .x(n37), .a(S4) );
    mux4_1 U252 ( .x(n295), .d0(D5_27), .d1(D13_27), .d2(D21_27), .d3(D29_27), 
        .sl0(n23), .sl1(n37) );
    buf_3 U253 ( .x(n39), .a(S4) );
    buf_3 U254 ( .x(n35), .a(S4) );
    buf_3 U255 ( .x(n33), .a(S4) );
    buf_3 U256 ( .x(n29), .a(S4) );
    mux4_1 U257 ( .x(n135), .d0(D4_27), .d1(D12_27), .d2(D20_27), .d3(D28_27), 
        .sl0(n11), .sl1(n29) );
    buf_3 U258 ( .x(n31), .a(S4) );
    mux4_1 U259 ( .x(n167), .d0(D2_27), .d1(D10_27), .d2(D18_27), .d3(D26_27), 
        .sl0(n10), .sl1(n31) );
    mux4_1 U26 ( .x(n279), .d0(D5_11), .d1(D13_11), .d2(D21_11), .d3(D29_11), 
        .sl0(n23), .sl1(n36) );
    buf_3 U260 ( .x(n27), .a(S4) );
    mux4_1 U261 ( .x(n103), .d0(D0_27), .d1(D8_27), .d2(D16_27), .d3(D24_27), 
        .sl0(n13), .sl1(n27) );
    buf_3 U262 ( .x(n40), .a(S4) );
    mux4_1 U263 ( .x(n332), .d0(D7_0), .d1(D15_0), .d2(D23_0), .d3(D31_0), 
        .sl0(n24), .sl1(n40) );
    buf_3 U264 ( .x(n36), .a(S4) );
    mux4_1 U265 ( .x(n268), .d0(D5_0), .d1(D13_0), .d2(D21_0), .d3(D29_0), 
        .sl0(n16), .sl1(n36) );
    buf_3 U266 ( .x(n38), .a(S4) );
    mux4_1 U267 ( .x(n300), .d0(D3_0), .d1(D11_0), .d2(D19_0), .d3(D27_0), 
        .sl0(n17), .sl1(n38) );
    buf_3 U268 ( .x(n34), .a(S4) );
    mux4_1 U269 ( .x(n236), .d0(D1_0), .d1(D9_0), .d2(D17_0), .d3(D25_0), 
        .sl0(n16), .sl1(n34) );
    mux4_1 U27 ( .x(n311), .d0(D3_11), .d1(D11_11), .d2(D19_11), .d3(D27_11), 
        .sl0(n8), .sl1(n38) );
    buf_3 U270 ( .x(n32), .a(S4) );
    mux4_1 U271 ( .x(n172), .d0(D6_0), .d1(D14_0), .d2(D22_0), .d3(D30_0), 
        .sl0(n10), .sl1(n32) );
    buf_3 U272 ( .x(n28), .a(S4) );
    mux4_1 U273 ( .x(n108), .d0(D4_0), .d1(D12_0), .d2(D20_0), .d3(D28_0), 
        .sl0(n12), .sl1(n28) );
    buf_3 U274 ( .x(n30), .a(S4) );
    mux4_1 U275 ( .x(n140), .d0(D2_0), .d1(D10_0), .d2(D18_0), .d3(D26_0), 
        .sl0(n14), .sl1(n30) );
    buf_3 U276 ( .x(n26), .a(S4) );
    mux4_1 U277 ( .x(n76), .d0(D0_0), .d1(D8_0), .d2(D16_0), .d3(D24_0), .sl0(
        n13), .sl1(n26) );
    mux2_2 U278 ( .x(Z_10), .d0(n54), .sl(S0), .d1(n214) );
    mux2_2 U279 ( .x(Z_31), .d0(n75), .sl(S0), .d1(n235) );
    mux4_1 U28 ( .x(n247), .d0(D1_11), .d1(D9_11), .d2(D17_11), .d3(D25_11), 
        .sl0(n16), .sl1(n34) );
    mux2_2 U280 ( .x(Z_20), .d0(n64), .sl(S0), .d1(n224) );
    mux2_2 U281 ( .x(Z_11), .d0(n55), .sl(S0), .d1(n215) );
    mux2_2 U282 ( .x(Z_1), .d0(n45), .sl(S0), .d1(n205) );
    mux2_2 U283 ( .x(Z_22), .d0(n66), .sl(S0), .d1(n226) );
    mux2_2 U284 ( .x(Z_6), .d0(n50), .sl(S0), .d1(n210) );
    mux2_2 U285 ( .x(Z_19), .d0(n63), .sl(S0), .d1(n223) );
    mux2_2 U286 ( .x(Z_9), .d0(n53), .sl(S0), .d1(n213) );
    mux2_2 U287 ( .x(Z_4), .d0(n48), .sl(S0), .d1(n208) );
    mux2_2 U288 ( .x(Z_24), .d0(n68), .sl(S0), .d1(n228) );
    mux2_2 U289 ( .x(Z_13), .d0(n57), .sl(S0), .d1(n217) );
    mux4_1 U29 ( .x(n183), .d0(D6_11), .d1(D14_11), .d2(D22_11), .d3(D30_11), 
        .sl0(n21), .sl1(n32) );
    mux2_2 U290 ( .x(Z_18), .d0(n62), .sl(S0), .d1(n222) );
    mux2_2 U291 ( .x(Z_12), .d0(n56), .sl(S0), .d1(n216) );
    mux2_2 U292 ( .x(Z_17), .d0(n61), .sl(S0), .d1(n221) );
    mux2_2 U293 ( .x(Z_26), .d0(n70), .sl(S0), .d1(n230) );
    mux2_2 U294 ( .x(Z_8), .d0(n52), .sl(S0), .d1(n212) );
    mux2_2 U295 ( .x(Z_7), .d0(n51), .sl(S0), .d1(n211) );
    mux2_2 U296 ( .x(Z_30), .d0(n74), .sl(S0), .d1(n234) );
    mux2_2 U297 ( .x(Z_21), .d0(n65), .sl(S0), .d1(n225) );
    mux2_2 U298 ( .x(Z_15), .d0(n59), .sl(S0), .d1(n219) );
    mux2_2 U299 ( .x(Z_14), .d0(n58), .sl(S0), .d1(n218) );
    mux4_1 U3 ( .x(n310), .d0(D3_10), .d1(D11_10), .d2(D19_10), .d3(D27_10), 
        .sl0(n24), .sl1(n38) );
    mux4_1 U30 ( .x(n119), .d0(D4_11), .d1(D12_11), .d2(D20_11), .d3(D28_11), 
        .sl0(n12), .sl1(n28) );
    mux2_2 U300 ( .x(Z_23), .d0(n67), .sl(S0), .d1(n227) );
    mux2_2 U301 ( .x(Z_5), .d0(n49), .sl(S0), .d1(n209) );
    mux2_2 U302 ( .x(Z_25), .d0(n69), .sl(S0), .d1(n229) );
    mux2_2 U303 ( .x(Z_16), .d0(n60), .sl(S0), .d1(n220) );
    mux2_2 U304 ( .x(Z_3), .d0(n47), .sl(S0), .d1(n207) );
    mux2_2 U305 ( .x(Z_28), .d0(n72), .sl(S0), .d1(n232) );
    mux2_2 U306 ( .x(Z_29), .d0(n73), .sl(S0), .d1(n233) );
    mux2_2 U307 ( .x(Z_0), .d0(n44), .sl(S0), .d1(n204) );
    buf_10 U308 ( .x(n2), .a(S1) );
    buf_10 U309 ( .x(n1), .a(S1) );
    mux4_1 U31 ( .x(n151), .d0(D2_11), .d1(D10_11), .d2(D18_11), .d3(D26_11), 
        .sl0(n20), .sl1(n30) );
    buf_4 U310 ( .x(n4), .a(S1) );
    buf_16 U313 ( .x(n7), .a(n43) );
    buf_16 U314 ( .x(n8), .a(n43) );
    buf_16 U315 ( .x(n9), .a(n43) );
    buf_16 U316 ( .x(n10), .a(n43) );
    buf_16 U317 ( .x(n11), .a(n43) );
    buf_16 U318 ( .x(n12), .a(n43) );
    buf_16 U319 ( .x(n13), .a(n43) );
    mux4_1 U32 ( .x(n87), .d0(D0_11), .d1(D8_11), .d2(D16_11), .d3(D24_11), 
        .sl0(n12), .sl1(n26) );
    buf_16 U320 ( .x(n14), .a(n43) );
    buf_16 U321 ( .x(n15), .a(n43) );
    buf_16 U322 ( .x(n16), .a(n43) );
    buf_16 U323 ( .x(n17), .a(n43) );
    buf_16 U324 ( .x(n18), .a(n43) );
    buf_16 U325 ( .x(n19), .a(n43) );
    buf_16 U326 ( .x(n20), .a(n43) );
    buf_16 U327 ( .x(n21), .a(n43) );
    buf_16 U328 ( .x(n22), .a(n43) );
    buf_16 U329 ( .x(n23), .a(n43) );
    mux4_1 U33 ( .x(n333), .d0(D7_1), .d1(D15_1), .d2(D23_1), .d3(D31_1), 
        .sl0(n18), .sl1(n40) );
    buf_16 U330 ( .x(n24), .a(n43) );
    inv_16 U331 ( .x(n43), .a(n42) );
    inv_16 U332 ( .x(n42), .a(S3) );
    mux2_4 U333 ( .x(Z_2), .d0(n46), .sl(S0), .d1(n206) );
    mux2_4 U334 ( .x(Z_27), .d0(n71), .sl(S0), .d1(n231) );
    mux4_3 U335 ( .x(n44), .d0(n76), .d1(n140), .d2(n108), .d3(n172), .sl0(n1), 
        .sl1(n5) );
    mux4_3 U336 ( .x(n45), .d0(n77), .d1(n141), .d2(n109), .d3(n173), .sl0(n2), 
        .sl1(n1425) );
    mux4_3 U337 ( .x(n46), .d0(n78), .d1(n142), .d2(n110), .d3(n174), .sl0(n4), 
        .sl1(n1425) );
    mux4_3 U338 ( .x(n47), .d0(n79), .d1(n143), .d2(n111), .d3(n175), .sl0(n2), 
        .sl1(n1425) );
    mux4_3 U339 ( .x(n48), .d0(n80), .d1(n144), .d2(n112), .d3(n176), .sl0(n1), 
        .sl1(n1425) );
    mux4_1 U34 ( .x(n269), .d0(D5_1), .d1(D13_1), .d2(D21_1), .d3(D29_1), 
        .sl0(n9), .sl1(n36) );
    mux4_3 U340 ( .x(n49), .d0(n81), .d1(n145), .d2(n113), .d3(n177), .sl0(n4), 
        .sl1(n1425) );
    mux4_3 U341 ( .x(n50), .d0(n82), .d1(n146), .d2(n114), .d3(n178), .sl0(n4), 
        .sl1(n1425) );
    mux4_3 U342 ( .x(n51), .d0(n83), .d1(n147), .d2(n115), .d3(n179), .sl0(n2), 
        .sl1(n1425) );
    mux4_3 U343 ( .x(n52), .d0(n84), .d1(n148), .d2(n116), .d3(n180), .sl0(n1), 
        .sl1(n1425) );
    mux4_3 U344 ( .x(n53), .d0(n85), .d1(n149), .d2(n117), .d3(n181), .sl0(n3), 
        .sl1(n1425) );
    mux4_3 U345 ( .x(n54), .d0(n86), .d1(n150), .d2(n118), .d3(n182), .sl0(n1), 
        .sl1(n1425) );
    mux4_3 U346 ( .x(n55), .d0(n87), .d1(n151), .d2(n119), .d3(n183), .sl0(n2), 
        .sl1(n1425) );
    mux4_3 U347 ( .x(n56), .d0(n88), .d1(n152), .d2(n120), .d3(n184), .sl0(n2), 
        .sl1(n1425) );
    mux4_3 U348 ( .x(n57), .d0(n89), .d1(n153), .d2(n121), .d3(n185), .sl0(n4), 
        .sl1(n5) );
    mux4_3 U349 ( .x(n59), .d0(n91), .d1(n155), .d2(n123), .d3(n187), .sl0(n1), 
        .sl1(n1425) );
    mux4_1 U35 ( .x(n301), .d0(D3_1), .d1(D11_1), .d2(D19_1), .d3(D27_1), 
        .sl0(n17), .sl1(n38) );
    mux4_3 U350 ( .x(n60), .d0(n92), .d1(n156), .d2(n124), .d3(n188), .sl0(n1), 
        .sl1(n1425) );
    mux4_3 U351 ( .x(n61), .d0(n93), .d1(n157), .d2(n125), .d3(n189), .sl0(n2), 
        .sl1(n1425) );
    mux4_3 U352 ( .x(n62), .d0(n94), .d1(n158), .d2(n126), .d3(n190), .sl0(n4), 
        .sl1(n5) );
    mux4_3 U353 ( .x(n63), .d0(n95), .d1(n159), .d2(n127), .d3(n191), .sl0(n3), 
        .sl1(n1425) );
    mux4_3 U354 ( .x(n64), .d0(n96), .d1(n160), .d2(n128), .d3(n192), .sl0(n4), 
        .sl1(n1425) );
    mux4_3 U355 ( .x(n65), .d0(n97), .d1(n161), .d2(n129), .d3(n193), .sl0(n2), 
        .sl1(n1425) );
    mux4_3 U356 ( .x(n66), .d0(n98), .d1(n162), .d2(n130), .d3(n194), .sl0(n2), 
        .sl1(n1425) );
    mux4_3 U357 ( .x(n67), .d0(n99), .d1(n163), .d2(n131), .d3(n195), .sl0(n1), 
        .sl1(n1425) );
    mux4_3 U358 ( .x(n68), .d0(n100), .d1(n164), .d2(n132), .d3(n196), .sl0(n4
        ), .sl1(n5) );
    mux4_3 U359 ( .x(n69), .d0(n101), .d1(n165), .d2(n133), .d3(n197), .sl0(n2
        ), .sl1(n5) );
    mux4_1 U36 ( .x(n237), .d0(D1_1), .d1(D9_1), .d2(D17_1), .d3(D25_1), .sl0(
        n9), .sl1(n34) );
    mux4_3 U360 ( .x(n70), .d0(n102), .d1(n166), .d2(n134), .d3(n198), .sl0(n2
        ), .sl1(n1425) );
    mux4_3 U361 ( .x(n71), .d0(n103), .d1(n167), .d2(n135), .d3(n199), .sl0(n3
        ), .sl1(n5) );
    mux4_3 U362 ( .x(n75), .d0(n107), .d1(n171), .d2(n139), .d3(n203), .sl0(n4
        ), .sl1(n1425) );
    mux4_3 U363 ( .x(n199), .d0(D6_27), .d1(D14_27), .d2(D22_27), .d3(D30_27), 
        .sl0(n21), .sl1(n33) );
    mux4_3 U364 ( .x(n204), .d0(n236), .d1(n300), .d2(n268), .d3(n332), .sl0(
        n4), .sl1(n5) );
    mux4_3 U365 ( .x(n205), .d0(n237), .d1(n301), .d2(n269), .d3(n333), .sl0(
        n3), .sl1(n5) );
    mux4_3 U366 ( .x(n206), .d0(n238), .d1(n302), .d2(n270), .d3(n334), .sl0(
        n3), .sl1(n5) );
    mux4_3 U367 ( .x(n207), .d0(n239), .d1(n303), .d2(n271), .d3(n335), .sl0(
        n1), .sl1(n5) );
    mux4_3 U368 ( .x(n208), .d0(n240), .d1(n304), .d2(n272), .d3(n336), .sl0(
        n4), .sl1(n1425) );
    mux4_3 U369 ( .x(n209), .d0(n241), .d1(n305), .d2(n273), .d3(n337), .sl0(
        n2), .sl1(n5) );
    mux4_1 U37 ( .x(n173), .d0(D6_1), .d1(D14_1), .d2(D22_1), .d3(D30_1), 
        .sl0(n21), .sl1(n32) );
    mux4_3 U370 ( .x(n210), .d0(n242), .d1(n306), .d2(n274), .d3(n338), .sl0(
        n2), .sl1(n1425) );
    mux4_3 U371 ( .x(n211), .d0(n243), .d1(n307), .d2(n275), .d3(n339), .sl0(
        n4), .sl1(n5) );
    mux4_3 U372 ( .x(n212), .d0(n244), .d1(n308), .d2(n276), .d3(n340), .sl0(
        n2), .sl1(n5) );
    mux4_3 U373 ( .x(n213), .d0(n245), .d1(n309), .d2(n277), .d3(n341), .sl0(
        n3), .sl1(n1425) );
    mux4_3 U374 ( .x(n214), .d0(n246), .d1(n310), .d2(n278), .d3(n342), .sl0(
        n3), .sl1(n1425) );
    mux4_3 U375 ( .x(n215), .d0(n247), .d1(n311), .d2(n279), .d3(n343), .sl0(
        n2), .sl1(n1425) );
    mux4_3 U376 ( .x(n216), .d0(n248), .d1(n312), .d2(n280), .d3(n344), .sl0(
        n1), .sl1(n1425) );
    mux4_3 U377 ( .x(n217), .d0(n249), .d1(n313), .d2(n281), .d3(n345), .sl0(
        n1), .sl1(n5) );
    mux4_3 U378 ( .x(n219), .d0(n251), .d1(n315), .d2(n283), .d3(n347), .sl0(
        n4), .sl1(n1425) );
    mux4_3 U379 ( .x(n220), .d0(n252), .d1(n316), .d2(n284), .d3(n348), .sl0(
        n2), .sl1(n5) );
    mux4_1 U38 ( .x(n109), .d0(D4_1), .d1(D12_1), .d2(D20_1), .d3(D28_1), 
        .sl0(n13), .sl1(n28) );
    mux4_3 U380 ( .x(n221), .d0(n253), .d1(n317), .d2(n285), .d3(n349), .sl0(
        n2), .sl1(n5) );
    mux4_3 U381 ( .x(n222), .d0(n254), .d1(n318), .d2(n286), .d3(n350), .sl0(
        n4), .sl1(n5) );
    mux4_3 U382 ( .x(n223), .d0(n255), .d1(n319), .d2(n287), .d3(n351), .sl0(
        n3), .sl1(n1425) );
    mux4_3 U383 ( .x(n224), .d0(n256), .d1(n320), .d2(n288), .d3(n352), .sl0(
        n1), .sl1(n1425) );
    mux4_3 U384 ( .x(n225), .d0(n257), .d1(n321), .d2(n289), .d3(n353), .sl0(
        n1), .sl1(n5) );
    mux4_3 U385 ( .x(n226), .d0(n258), .d1(n322), .d2(n290), .d3(n354), .sl0(
        n4), .sl1(n5) );
    mux4_3 U386 ( .x(n227), .d0(n259), .d1(n323), .d2(n291), .d3(n355), .sl0(
        n1), .sl1(n5) );
    mux4_3 U387 ( .x(n228), .d0(n260), .d1(n324), .d2(n292), .d3(n356), .sl0(
        n1), .sl1(n5) );
    mux4_3 U388 ( .x(n229), .d0(n261), .d1(n325), .d2(n293), .d3(n357), .sl0(
        n1), .sl1(n5) );
    mux4_3 U389 ( .x(n230), .d0(n262), .d1(n326), .d2(n294), .d3(n358), .sl0(
        n4), .sl1(n5) );
    mux4_1 U39 ( .x(n141), .d0(D2_1), .d1(D10_1), .d2(D18_1), .d3(D26_1), 
        .sl0(n20), .sl1(n30) );
    mux4_3 U390 ( .x(n231), .d0(n263), .d1(n327), .d2(n295), .d3(n359), .sl0(
        n3), .sl1(n5) );
    mux4_3 U391 ( .x(n234), .d0(n266), .d1(n330), .d2(n298), .d3(n362), .sl0(
        n3), .sl1(n5) );
    mux4_3 U392 ( .x(n235), .d0(n267), .d1(n331), .d2(n299), .d3(n363), .sl0(
        n1), .sl1(n1425) );
    mux4_3 U393 ( .x(n263), .d0(D1_27), .d1(D9_27), .d2(D17_27), .d3(D25_27), 
        .sl0(n22), .sl1(n35) );
    mux4_3 U394 ( .x(n327), .d0(D3_27), .d1(D11_27), .d2(D19_27), .d3(D27_27), 
        .sl0(n7), .sl1(n39) );
    mux4_3 U395 ( .x(n359), .d0(D7_27), .d1(D15_27), .d2(D23_27), .d3(D31_27), 
        .sl0(n19), .sl1(n41) );
    buf_3 U396 ( .x(n1425), .a(S2) );
    buf_3 U397 ( .x(n5), .a(S2) );
    mux4_1 U4 ( .x(n246), .d0(D1_10), .d1(D9_10), .d2(D17_10), .d3(D25_10), 
        .sl0(n9), .sl1(n34) );
    mux4_1 U40 ( .x(n77), .d0(D0_1), .d1(D8_1), .d2(D16_1), .d3(D24_1), .sl0(
        n13), .sl1(n26) );
    mux4_1 U41 ( .x(n354), .d0(D7_22), .d1(D15_22), .d2(D23_22), .d3(D31_22), 
        .sl0(n7), .sl1(n41) );
    mux4_1 U42 ( .x(n290), .d0(D5_22), .d1(D13_22), .d2(D21_22), .d3(D29_22), 
        .sl0(n23), .sl1(n37) );
    mux4_1 U43 ( .x(n322), .d0(D3_22), .d1(D11_22), .d2(D19_22), .d3(D27_22), 
        .sl0(n24), .sl1(n39) );
    mux4_1 U44 ( .x(n258), .d0(D1_22), .d1(D9_22), .d2(D17_22), .d3(D25_22), 
        .sl0(n9), .sl1(n35) );
    mux4_1 U45 ( .x(n194), .d0(D6_22), .d1(D14_22), .d2(D22_22), .d3(D30_22), 
        .sl0(n10), .sl1(n33) );
    mux4_1 U46 ( .x(n130), .d0(D4_22), .d1(D12_22), .d2(D20_22), .d3(D28_22), 
        .sl0(n11), .sl1(n29) );
    mux4_1 U47 ( .x(n162), .d0(D2_22), .d1(D10_22), .d2(D18_22), .d3(D26_22), 
        .sl0(n10), .sl1(n31) );
    mux4_1 U48 ( .x(n98), .d0(D0_22), .d1(D8_22), .d2(D16_22), .d3(D24_22), 
        .sl0(n13), .sl1(n27) );
    mux4_1 U49 ( .x(n334), .d0(D7_2), .d1(D15_2), .d2(D23_2), .d3(D31_2), 
        .sl0(n24), .sl1(n40) );
    mux4_1 U5 ( .x(n182), .d0(D6_10), .d1(D14_10), .d2(D22_10), .d3(D30_10), 
        .sl0(n15), .sl1(n32) );
    mux4_1 U50 ( .x(n270), .d0(D5_2), .d1(D13_2), .d2(D21_2), .d3(D29_2), 
        .sl0(n22), .sl1(n36) );
    mux4_1 U51 ( .x(n302), .d0(D3_2), .d1(D11_2), .d2(D19_2), .d3(D27_2), 
        .sl0(n17), .sl1(n38) );
    mux4_1 U52 ( .x(n238), .d0(D1_2), .d1(D9_2), .d2(D17_2), .d3(D25_2), .sl0(
        n22), .sl1(n34) );
    mux4_1 U53 ( .x(n174), .d0(D6_2), .d1(D14_2), .d2(D22_2), .d3(D30_2), 
        .sl0(n10), .sl1(n32) );
    mux4_1 U54 ( .x(n110), .d0(D4_2), .d1(D12_2), .d2(D20_2), .d3(D28_2), 
        .sl0(n12), .sl1(n28) );
    mux4_1 U55 ( .x(n142), .d0(D2_2), .d1(D10_2), .d2(D18_2), .d3(D26_2), 
        .sl0(n11), .sl1(n30) );
    mux4_1 U56 ( .x(n78), .d0(D0_2), .d1(D8_2), .d2(D16_2), .d3(D24_2), .sl0(
        n12), .sl1(n26) );
    mux4_1 U57 ( .x(n338), .d0(D7_6), .d1(D15_6), .d2(D23_6), .d3(D31_6), 
        .sl0(n18), .sl1(n40) );
    mux4_1 U58 ( .x(n274), .d0(D5_6), .d1(D13_6), .d2(D21_6), .d3(D29_6), 
        .sl0(n9), .sl1(n36) );
    mux4_1 U59 ( .x(n306), .d0(D3_6), .d1(D11_6), .d2(D19_6), .d3(D27_6), 
        .sl0(n23), .sl1(n38) );
    mux4_1 U6 ( .x(n118), .d0(D4_10), .d1(D12_10), .d2(D20_10), .d3(D28_10), 
        .sl0(n14), .sl1(n28) );
    mux4_1 U60 ( .x(n242), .d0(D1_6), .d1(D9_6), .d2(D17_6), .d3(D25_6), .sl0(
        n16), .sl1(n34) );
    mux4_1 U61 ( .x(n178), .d0(D6_6), .d1(D14_6), .d2(D22_6), .d3(D30_6), 
        .sl0(n10), .sl1(n32) );
    mux4_1 U62 ( .x(n114), .d0(D4_6), .d1(D12_6), .d2(D20_6), .d3(D28_6), 
        .sl0(n19), .sl1(n28) );
    mux4_1 U63 ( .x(n146), .d0(D2_6), .d1(D10_6), .d2(D18_6), .d3(D26_6), 
        .sl0(n14), .sl1(n30) );
    mux4_1 U64 ( .x(n82), .d0(D0_6), .d1(D8_6), .d2(D16_6), .d3(D24_6), .sl0(
        n12), .sl1(n26) );
    mux4_1 U65 ( .x(n351), .d0(D7_19), .d1(D15_19), .d2(D23_19), .d3(D31_19), 
        .sl0(n7), .sl1(n41) );
    mux4_1 U66 ( .x(n287), .d0(D5_19), .d1(D13_19), .d2(D21_19), .d3(D29_19), 
        .sl0(n17), .sl1(n37) );
    mux4_1 U67 ( .x(n319), .d0(D3_19), .d1(D11_19), .d2(D19_19), .d3(D27_19), 
        .sl0(n24), .sl1(n39) );
    mux4_1 U68 ( .x(n255), .d0(D1_19), .d1(D9_19), .d2(D17_19), .d3(D25_19), 
        .sl0(n9), .sl1(n35) );
    mux4_1 U69 ( .x(n191), .d0(D6_19), .d1(D14_19), .d2(D22_19), .d3(D30_19), 
        .sl0(n10), .sl1(n33) );
    mux4_1 U7 ( .x(n150), .d0(D2_10), .d1(D10_10), .d2(D18_10), .d3(D26_10), 
        .sl0(n14), .sl1(n30) );
    mux4_1 U70 ( .x(n127), .d0(D4_19), .d1(D12_19), .d2(D20_19), .d3(D28_19), 
        .sl0(n11), .sl1(n29) );
    mux4_1 U71 ( .x(n159), .d0(D2_19), .d1(D10_19), .d2(D18_19), .d3(D26_19), 
        .sl0(n21), .sl1(n31) );
    mux4_1 U72 ( .x(n95), .d0(D0_19), .d1(D8_19), .d2(D16_19), .d3(D24_19), 
        .sl0(n12), .sl1(n27) );
    mux4_1 U73 ( .x(n341), .d0(D7_9), .d1(D15_9), .d2(D23_9), .d3(D31_9), 
        .sl0(n24), .sl1(n40) );
    mux4_1 U74 ( .x(n277), .d0(D5_9), .d1(D13_9), .d2(D21_9), .d3(D29_9), 
        .sl0(n8), .sl1(n36) );
    mux4_1 U75 ( .x(n309), .d0(D3_9), .d1(D11_9), .d2(D19_9), .d3(D27_9), 
        .sl0(n23), .sl1(n38) );
    mux4_1 U76 ( .x(n245), .d0(D1_9), .d1(D9_9), .d2(D17_9), .d3(D25_9), .sl0(
        n22), .sl1(n34) );
    mux4_1 U77 ( .x(n181), .d0(D6_9), .d1(D14_9), .d2(D22_9), .d3(D30_9), 
        .sl0(n10), .sl1(n32) );
    mux4_1 U78 ( .x(n117), .d0(D4_9), .d1(D12_9), .d2(D20_9), .d3(D28_9), 
        .sl0(n20), .sl1(n28) );
    mux4_1 U79 ( .x(n149), .d0(D2_9), .d1(D10_9), .d2(D18_9), .d3(D26_9), 
        .sl0(n14), .sl1(n30) );
    mux4_1 U8 ( .x(n86), .d0(D0_10), .d1(D8_10), .d2(D16_10), .d3(D24_10), 
        .sl0(n19), .sl1(n26) );
    mux4_1 U80 ( .x(n85), .d0(D0_9), .d1(D8_9), .d2(D16_9), .d3(D24_9), .sl0(
        n13), .sl1(n26) );
    mux4_1 U81 ( .x(n336), .d0(D7_4), .d1(D15_4), .d2(D23_4), .d3(D31_4), 
        .sl0(n7), .sl1(n40) );
    mux4_1 U82 ( .x(n272), .d0(D5_4), .d1(D13_4), .d2(D21_4), .d3(D29_4), 
        .sl0(n9), .sl1(n36) );
    mux4_1 U83 ( .x(n304), .d0(D3_4), .d1(D11_4), .d2(D19_4), .d3(D27_4), 
        .sl0(n8), .sl1(n38) );
    mux4_1 U84 ( .x(n240), .d0(D1_4), .d1(D9_4), .d2(D17_4), .d3(D25_4), .sl0(
        n9), .sl1(n34) );
    mux4_1 U85 ( .x(n176), .d0(D6_4), .d1(D14_4), .d2(D22_4), .d3(D30_4), 
        .sl0(n15), .sl1(n32) );
    mux4_1 U86 ( .x(n112), .d0(D4_4), .d1(D12_4), .d2(D20_4), .d3(D28_4), 
        .sl0(n13), .sl1(n28) );
    mux4_1 U87 ( .x(n144), .d0(D2_4), .d1(D10_4), .d2(D18_4), .d3(D26_4), 
        .sl0(n20), .sl1(n30) );
    mux4_1 U88 ( .x(n80), .d0(D0_4), .d1(D8_4), .d2(D16_4), .d3(D24_4), .sl0(
        n19), .sl1(n26) );
    mux4_1 U89 ( .x(n356), .d0(D7_24), .d1(D15_24), .d2(D23_24), .d3(D31_24), 
        .sl0(n18), .sl1(n41) );
    mux4_1 U9 ( .x(n363), .d0(D7_31), .d1(D15_31), .d2(D23_31), .d3(D31_31), 
        .sl0(n25), .sl1(n41) );
    mux4_1 U90 ( .x(n292), .d0(D5_24), .d1(D13_24), .d2(D21_24), .d3(D29_24), 
        .sl0(n23), .sl1(n37) );
    mux4_1 U91 ( .x(n324), .d0(D3_24), .d1(D11_24), .d2(D19_24), .d3(D27_24), 
        .sl0(n18), .sl1(n39) );
    mux4_1 U92 ( .x(n260), .d0(D1_24), .d1(D9_24), .d2(D17_24), .d3(D25_24), 
        .sl0(n9), .sl1(n35) );
    mux4_1 U93 ( .x(n196), .d0(D6_24), .d1(D14_24), .d2(D22_24), .d3(D30_24), 
        .sl0(n21), .sl1(n33) );
    mux4_1 U94 ( .x(n132), .d0(D4_24), .d1(D12_24), .d2(D20_24), .d3(D28_24), 
        .sl0(n14), .sl1(n29) );
    mux4_1 U95 ( .x(n164), .d0(D2_24), .d1(D10_24), .d2(D18_24), .d3(D26_24), 
        .sl0(n15), .sl1(n31) );
    mux4_1 U96 ( .x(n100), .d0(D0_24), .d1(D8_24), .d2(D16_24), .d3(D24_24), 
        .sl0(n12), .sl1(n27) );
    mux4_1 U97 ( .x(n345), .d0(D7_13), .d1(D15_13), .d2(D23_13), .d3(D31_13), 
        .sl0(n18), .sl1(n40) );
    mux4_1 U98 ( .x(n281), .d0(D5_13), .d1(D13_13), .d2(D21_13), .d3(D29_13), 
        .sl0(n8), .sl1(n36) );
    mux4_1 U99 ( .x(n313), .d0(D3_13), .d1(D11_13), .d2(D19_13), .d3(D27_13), 
        .sl0(n17), .sl1(n38) );
endmodule


module ID_DW01_sub_32_2_test_1 ( A, B, CI, DIFF, CO );
input  [31:0] A;
input  [31:0] B;
output [31:0] DIFF;
input  CI;
output CO;
    wire A_1, A_0, n176, n67, n157, n81, n170, n155, n63, n130, n62, n129, n71, 
        n167, n64, n136, n95, n96, n97, n90, n177, n124, n142, n169, n137, n65, 
        n161, n70, n162, n135, n165, n104, n68, n69, n199, n87, n160, n173, 
        n174, n99, n188, n149, n198, n197, n189, n187, n182, n181, n180, n179, 
        n193, n72, n166, n164, n163, n84, n191, n184, n83, n195, n76, n77, n78, 
        n86, n88, n112, n113, n114, n139, n140, n141, n192, n190, n144, n172, 
        n171, n200, n74, n85, n201, n98, n101, n146, n202, n105, n194, n106, 
        n153, n110, n203, n151, n178, n122, n150, n120, n111, n109, n107, n102, 
        n123, n125, n89, n196, n126, n127, n128, n159, n132, n75, n91, n94, 
        n186, n100, n143, n152, n121, n148, n147, n145, n175, n119, n133, n117, 
        n118, n134, n103, n50, n156, n66, n73, n204, n206, n205, n116, n115, 
        n56, n154, n168, n108, n185, n183, n131, n80, n92, n93, n82, n57, n79, 
        n158, n52, n138, n55, n58, n59, n60, n61;
    assign A_1 = A[1];
    assign A_0 = A[0];
    assign DIFF[1] = A_1;
    assign DIFF[0] = A_0;
    nor2_1 U10 ( .x(n176), .a(A[29]), .b(A[28]) );
    nor2i_2 U100 ( .x(n67), .a(n157), .b(n81) );
    nor2_1 U101 ( .x(n170), .a(A[9]), .b(A[8]) );
    nor2_1 U102 ( .x(n155), .a(A[6]), .b(A[10]) );
    oa21_4 U103 ( .x(DIFF[6]), .a(n63), .b(n130), .c(n62) );
    nand2_0 U104 ( .x(n62), .a(n129), .b(n71) );
    nand2_1 U105 ( .x(n63), .a(n167), .b(n64) );
    inv_1 U106 ( .x(n64), .a(n136) );
    oai21_5 U108 ( .x(DIFF[17]), .a(n95), .b(n96), .c(n97) );
    inv_0 U109 ( .x(n90), .a(A[15]) );
    nand2i_2 U11 ( .x(n177), .a(A[27]), .b(n124) );
    nand3i_1 U110 ( .x(n142), .a(A[15]), .b(n169), .c(n137) );
    mux2_2 U111 ( .x(n65), .d0(n161), .sl(n167), .d1(n136) );
    nand2i_1 U112 ( .x(n136), .a(A[4]), .b(n137) );
    inv_1 U113 ( .x(n161), .a(n70) );
    nand2i_0 U114 ( .x(n162), .a(A[8]), .b(n135) );
    inv_2 U115 ( .x(DIFF[2]), .a(A[2]) );
    nor2_0 U116 ( .x(n165), .a(A[2]), .b(A[3]) );
    inv_0 U118 ( .x(n104), .a(A[20]) );
    oai21_1 U119 ( .x(DIFF[4]), .a(n68), .b(n69), .c(n70) );
    inv_0 U120 ( .x(n129), .a(A[6]) );
    nand2i_2 U121 ( .x(n199), .a(A[12]), .b(n157) );
    inv_0 U122 ( .x(n87), .a(A[13]) );
    nand2i_2 U123 ( .x(n70), .a(A[4]), .b(n160) );
    nor2_1 U124 ( .x(n173), .a(A[10]), .b(A[13]) );
    nand3i_1 U125 ( .x(n174), .a(A[14]), .b(n99), .c(n173) );
    nor2_1 U126 ( .x(n188), .a(A[13]), .b(A[14]) );
    inv_2 U127 ( .x(n149), .a(A[3]) );
    nand2i_0 U129 ( .x(n198), .a(A[11]), .b(n197) );
    nand3i_0 U130 ( .x(n189), .a(A[11]), .b(n188), .c(n187) );
    nand4i_1 U131 ( .x(n182), .a(A[11]), .b(n181), .c(n180), .d(n179) );
    nor2_0 U133 ( .x(n193), .a(A[9]), .b(A[8]) );
    nand4i_1 U134 ( .x(n72), .a(A[7]), .b(n165), .c(n166), .d(n69) );
    nand2i_0 U135 ( .x(n164), .a(A[7]), .b(n163) );
    inv_0 U136 ( .x(n84), .a(A[12]) );
    nor2_0 U137 ( .x(n197), .a(A[12]), .b(A[13]) );
    nor2_0 U138 ( .x(n191), .a(A[12]), .b(A[11]) );
    nor2_0 U139 ( .x(n184), .a(A[12]), .b(A[11]) );
    nand2i_0 U14 ( .x(n83), .a(n157), .b(n81) );
    nor2_0 U140 ( .x(n180), .a(A[15]), .b(A[12]) );
    inv_0 U141 ( .x(n167), .a(A[5]) );
    nor2_0 U142 ( .x(n166), .a(A[6]), .b(A[5]) );
    nor3_0 U143 ( .x(n195), .a(A[4]), .b(A[6]), .c(A[5]) );
    oai21_4 U146 ( .x(DIFF[9]), .a(n76), .b(n77), .c(n78) );
    oai21_4 U147 ( .x(DIFF[13]), .a(n86), .b(n87), .c(n88) );
    oai21_4 U148 ( .x(DIFF[24]), .a(n112), .b(n113), .c(n114) );
    nand2i_4 U149 ( .x(n139), .a(n140), .b(n141) );
    nor2i_1 U15 ( .x(n192), .a(n191), .b(n190) );
    and3i_3 U150 ( .x(n144), .a(n174), .b(n172), .c(n171) );
    inv_5 U151 ( .x(n68), .a(n200) );
    nand2i_4 U152 ( .x(n74), .a(n162), .b(n130) );
    nand2i_4 U153 ( .x(n78), .a(n164), .b(n130) );
    nand2i_4 U154 ( .x(n85), .a(n199), .b(n201) );
    inv_5 U155 ( .x(n86), .a(n85) );
    nand2i_4 U156 ( .x(n88), .a(n198), .b(n201) );
    inv_5 U157 ( .x(n98), .a(n97) );
    nand2i_4 U158 ( .x(n101), .a(A[19]), .b(n146) );
    inv_5 U159 ( .x(n202), .a(n105) );
    nand2i_0 U16 ( .x(n194), .a(A[7]), .b(n193) );
    nand2_5 U160 ( .x(n106), .a(n202), .b(n153) );
    nand2_5 U161 ( .x(n110), .a(n203), .b(n151) );
    nand2i_4 U162 ( .x(n114), .a(n178), .b(n203) );
    nand2i_4 U165 ( .x(n122), .a(n150), .b(n120) );
    nand2i_4 U166 ( .x(n111), .a(n151), .b(n109) );
    nand2i_4 U167 ( .x(n107), .a(n153), .b(n105) );
    nand2_5 U168 ( .x(DIFF[19]), .a(n101), .b(n102) );
    oai21_5 U169 ( .x(DIFF[28]), .a(n123), .b(n124), .c(n125) );
    nand4i_1 U17 ( .x(n89), .a(n194), .b(n192), .c(n196), .d(n195) );
    oai21_5 U170 ( .x(DIFF[29]), .a(n126), .b(n127), .c(n128) );
    exnor2_5 U171 ( .x(DIFF[30]), .a(n159), .b(n132) );
    nand2_5 U172 ( .x(DIFF[8]), .a(n74), .b(n75) );
    nand2i_5 U173 ( .x(n91), .a(n189), .b(n201) );
    nand2i_5 U174 ( .x(n94), .a(n186), .b(n201) );
    nand2i_5 U175 ( .x(n97), .a(n182), .b(n201) );
    nand3i_5 U176 ( .x(n100), .a(n142), .b(n143), .c(n144) );
    nand2i_6 U178 ( .x(n105), .a(n152), .b(n146) );
    inv_2 U18 ( .x(n69), .a(A[4]) );
    inv_6 U180 ( .x(n123), .a(n121) );
    nand2i_6 U181 ( .x(n125), .a(n177), .b(n148) );
    nand2i_6 U182 ( .x(n128), .a(n147), .b(n148) );
    nor2i_5 U183 ( .x(n143), .a(n170), .b(n199) );
    nand2_3 U185 ( .x(n145), .a(n175), .b(n119) );
    nor2_1 U187 ( .x(n133), .a(A[5]), .b(A[6]) );
    ao21_4 U188 ( .x(DIFF[26]), .a(n117), .b(A[26]), .c(n148) );
    inv_2 U189 ( .x(n118), .a(n117) );
    inv_4 U190 ( .x(n119), .a(A[26]) );
    nand2i_4 U191 ( .x(n120), .a(n145), .b(n146) );
    inv_7 U192 ( .x(n148), .a(n120) );
    nand2i_1 U193 ( .x(n117), .a(n139), .b(n146) );
    nand3_1 U194 ( .x(n71), .a(n69), .b(n133), .c(n134) );
    nor2_0 U195 ( .x(n172), .a(A[5]), .b(A[6]) );
    nand2_1 U196 ( .x(n102), .a(A[19]), .b(n100) );
    inv_8 U197 ( .x(n146), .a(n100) );
    oai21_2 U198 ( .x(DIFF[20]), .a(n104), .b(n103), .c(n105) );
    nand4_5 U199 ( .x(n81), .a(n68), .b(n50), .c(n155), .d(n156) );
    nand2i_2 U20 ( .x(n75), .a(n66), .b(n72) );
    inv_4 U200 ( .x(n130), .a(n71) );
    nand2i_1 U201 ( .x(n73), .a(n135), .b(n71) );
    aoi21_6 U202 ( .x(n204), .a(n206), .b(n205), .c(n118) );
    inv_7 U203 ( .x(DIFF[25]), .a(n204) );
    inv_2 U204 ( .x(n205), .a(n116) );
    inv_10 U205 ( .x(n206), .a(n115) );
    inv_7 U206 ( .x(n115), .a(n114) );
    nor2_3 U207 ( .x(n56), .a(A[20]), .b(A[19]) );
    nand2i_2 U208 ( .x(n152), .a(A[20]), .b(n154) );
    nor2_2 U209 ( .x(n168), .a(A[25]), .b(A[24]) );
    inv_2 U21 ( .x(n175), .a(n139) );
    nand2i_0 U210 ( .x(n178), .a(A[24]), .b(n151) );
    inv_6 U211 ( .x(n96), .a(A[17]) );
    nor2_1 U212 ( .x(n179), .a(A[17]), .b(A[16]) );
    inv_3 U213 ( .x(n66), .a(A[8]) );
    nor2_1 U214 ( .x(n163), .a(A[9]), .b(A[8]) );
    inv_4 U215 ( .x(n108), .a(A[22]) );
    nand3_1 U22 ( .x(n186), .a(n185), .b(n183), .c(n184) );
    nor2_0 U24 ( .x(n181), .a(A[14]), .b(A[13]) );
    nor2i_1 U26 ( .x(n131), .a(n132), .b(n128) );
    inv_1 U27 ( .x(n80), .a(A[10]) );
    nand2_3 U28 ( .x(n121), .a(n148), .b(n150) );
    nand2_2 U29 ( .x(DIFF[27]), .a(n121), .b(n122) );
    nand2_2 U30 ( .x(DIFF[7]), .a(n72), .b(n73) );
    inv_2 U31 ( .x(n126), .a(n125) );
    inv_2 U34 ( .x(n95), .a(n94) );
    inv_2 U35 ( .x(n92), .a(n91) );
    oai21_1 U36 ( .x(DIFF[16]), .a(n92), .b(n93), .c(n94) );
    nand2_2 U37 ( .x(DIFF[11]), .a(n82), .b(n83) );
    inv_2 U38 ( .x(n82), .a(n67) );
    inv_5 U39 ( .x(n203), .a(n109) );
    nor2_0 U4 ( .x(n187), .a(A[15]), .b(A[12]) );
    oai21_3 U40 ( .x(DIFF[15]), .a(n57), .b(n90), .c(n91) );
    inv_2 U41 ( .x(n79), .a(n78) );
    inv_2 U42 ( .x(n76), .a(n74) );
    inv_2 U44 ( .x(n112), .a(n110) );
    nand2_2 U45 ( .x(DIFF[21]), .a(n106), .b(n107) );
    oai21_2 U46 ( .x(DIFF[18]), .a(n98), .b(n99), .c(n100) );
    nand2_2 U47 ( .x(DIFF[23]), .a(n110), .b(n111) );
    inv_2 U48 ( .x(n159), .a(n128) );
    exnor2_1 U49 ( .x(DIFF[31]), .a(n131), .b(n158) );
    nand2i_2 U5 ( .x(n190), .a(A[2]), .b(n149) );
    inv_3 U50 ( .x(DIFF[5]), .a(n65) );
    inv_2 U51 ( .x(n99), .a(A[18]) );
    inv_0 U52 ( .x(n113), .a(A[24]) );
    inv_0 U53 ( .x(n116), .a(A[25]) );
    inv_2 U54 ( .x(n151), .a(A[23]) );
    inv_2 U55 ( .x(n135), .a(A[7]) );
    inv_2 U57 ( .x(n150), .a(A[27]) );
    inv_2 U58 ( .x(n124), .a(A[28]) );
    inv_2 U59 ( .x(n127), .a(A[29]) );
    nand2i_2 U6 ( .x(n140), .a(A[23]), .b(n168) );
    inv_2 U60 ( .x(n132), .a(A[30]) );
    inv_2 U61 ( .x(n158), .a(A[31]) );
    and3_5 U62 ( .x(n50), .a(n135), .b(n66), .c(n77) );
    ao21_6 U63 ( .x(DIFF[22]), .a(n106), .b(n52), .c(n203) );
    inv_2 U64 ( .x(n52), .a(n108) );
    nand2i_4 U66 ( .x(n109), .a(n138), .b(n146) );
    oai21_3 U69 ( .x(DIFF[12]), .a(n84), .b(n67), .c(n85) );
    nor2_0 U7 ( .x(n185), .a(A[13]), .b(A[14]) );
    nor2_1 U70 ( .x(n156), .a(A[4]), .b(A[5]) );
    inv_3 U71 ( .x(n77), .a(A[9]) );
    inv_5 U72 ( .x(n57), .a(n89) );
    nand3_2 U73 ( .x(n138), .a(n153), .b(n108), .c(n56) );
    or2_2 U75 ( .x(n55), .a(A[7]), .b(A[4]) );
    inv_2 U76 ( .x(n171), .a(n55) );
    inv_10 U77 ( .x(n201), .a(n81) );
    inv_2 U8 ( .x(n141), .a(n138) );
    nor2_0 U81 ( .x(n183), .a(A[16]), .b(A[15]) );
    inv_0 U82 ( .x(n93), .a(A[16]) );
    nor2_3 U83 ( .x(n137), .a(A[2]), .b(A[3]) );
    nor2_1 U84 ( .x(n134), .a(A[2]), .b(A[3]) );
    inv_0 U85 ( .x(n154), .a(A[19]) );
    ao21_3 U86 ( .x(DIFF[14]), .a(n88), .b(A[14]), .c(n57) );
    nand2i_2 U87 ( .x(n58), .a(A[16]), .b(n96) );
    inv_2 U88 ( .x(n169), .a(n58) );
    oai21_1 U89 ( .x(DIFF[3]), .a(n149), .b(n59), .c(n200) );
    nand2i_2 U9 ( .x(n147), .a(A[27]), .b(n176) );
    inv_0 U90 ( .x(n59), .a(A[2]) );
    and3_2 U91 ( .x(n196), .a(n60), .b(n80), .c(n61) );
    inv_0 U92 ( .x(n60), .a(A[13]) );
    inv_0 U93 ( .x(n61), .a(A[14]) );
    inv_6 U94 ( .x(n103), .a(n101) );
    nand2i_4 U95 ( .x(n200), .a(A[2]), .b(n149) );
    nor2_1 U96 ( .x(n160), .a(A[2]), .b(A[3]) );
    inv_2 U97 ( .x(n153), .a(A[21]) );
    inv_5 U98 ( .x(n157), .a(A[11]) );
    oai21_1 U99 ( .x(DIFF[10]), .a(n79), .b(n80), .c(n81) );
endmodule


module ID_DW01_sub_32_0_test_1 ( A, B, CI, DIFF, CO );
input  [31:0] A;
input  [31:0] B;
output [31:0] DIFF;
input  CI;
output CO;
    wire A_1, A_0, n123, n162, n121, n110, n177, n116, n130, n131, n132, n127, 
        n160, n124, n57, n125, n161, n55, n87, n88, n56, n91, n142, n166, n80, 
        n79, n168, n58, n140, n139, n136, n90, n103, n96, n64, n182, n115, n54, 
        n143, n178, n138, n148, n149, n170, n147, n179, n73, n61, n106, n119, 
        n120, n70, n146, n118, n107, n65, n66, n151, n153, n137, n67, n141, 
        n111, n84, n169, n71, n112, n113, n114, n172, n176, n82, n99, n100, 
        n101, n117, n133, n134, n128, n156, n157, n150, n181, n158, n97, n76, 
        n129, n77, n159, n126, n122, n163, n164, n98, n165, n85, n86, n94, n93, 
        n109, n95, n154, n155, n78, n81, n50, n72, n174, n60, n183, n83, n175, 
        n171, n108, n102, n104, n68, n135, n92, n75, n167, n152, n53, n51, 
        n105, n145, n69, n144, n173, n63, n62, n59, n52, n180, n89;
    assign A_1 = A[1];
    assign A_0 = A[0];
    assign DIFF[1] = A_1;
    assign DIFF[0] = A_0;
    nand2i_1 U10 ( .x(n123), .a(n162), .b(n121) );
    nand2_4 U100 ( .x(n110), .a(n177), .b(n116) );
    nor2i_2 U101 ( .x(n130), .a(n131), .b(n132) );
    nand2i_2 U102 ( .x(n127), .a(n160), .b(n124) );
    nor2i_5 U103 ( .x(n57), .a(n162), .b(n121) );
    nand2i_2 U104 ( .x(n125), .a(n161), .b(n55) );
    nand2_5 U105 ( .x(DIFF[25]), .a(n55), .b(n123) );
    ao21_6 U106 ( .x(DIFF[8]), .a(A[8]), .b(n87), .c(n88) );
    inv_2 U107 ( .x(n56), .a(n121) );
    nand2i_4 U108 ( .x(n124), .a(A[26]), .b(n57) );
    or3i_5 U109 ( .x(n91), .a(n142), .b(n166), .c(n80) );
    inv_10 U11 ( .x(n79), .a(A[4]) );
    nand2i_4 U110 ( .x(n168), .a(n80), .b(n142) );
    inv_0 U111 ( .x(n162), .a(A[25]) );
    nand3i_1 U112 ( .x(n58), .a(A[7]), .b(n140), .c(n139) );
    inv_10 U113 ( .x(n142), .a(n136) );
    nand2i_4 U115 ( .x(n166), .a(A[9]), .b(n90) );
    inv_5 U116 ( .x(n103), .a(A[15]) );
    nand2i_4 U117 ( .x(n96), .a(n64), .b(n182) );
    nor3_2 U118 ( .x(n115), .a(n54), .b(A[19]), .c(n143) );
    inv_7 U119 ( .x(n178), .a(n54) );
    nor2i_2 U12 ( .x(n138), .a(n148), .b(n149) );
    nor2_3 U120 ( .x(n170), .a(n54), .b(n147) );
    nand2i_1 U121 ( .x(n179), .a(A[15]), .b(n73) );
    nand2_5 U123 ( .x(n61), .a(n106), .b(n103) );
    nand2_6 U124 ( .x(DIFF[23]), .a(n119), .b(n120) );
    nand2_1 U125 ( .x(n70), .a(n146), .b(n142) );
    nand2_6 U126 ( .x(n118), .a(n170), .b(n116) );
    nand2i_4 U127 ( .x(n107), .a(n54), .b(n116) );
    nor2i_3 U128 ( .x(n65), .a(n66), .b(n151) );
    inv_5 U129 ( .x(n153), .a(n65) );
    nor2i_3 U13 ( .x(n137), .a(n138), .b(n70) );
    inv_0 U131 ( .x(n67), .a(A[6]) );
    mux2i_3 U132 ( .x(DIFF[9]), .d0(n141), .sl(A[9]), .d1(n88) );
    nand2_8 U133 ( .x(n111), .a(n146), .b(n142) );
    nor2_1 U134 ( .x(n84), .a(A[2]), .b(A[4]) );
    nor2_1 U135 ( .x(n169), .a(A[2]), .b(A[4]) );
    nand2_0 U136 ( .x(n71), .a(n146), .b(n142) );
    oai22_2 U137 ( .x(DIFF[18]), .a(n112), .b(n71), .c(n113), .d(n114) );
    nand2i_4 U138 ( .x(n143), .a(A[17]), .b(n114) );
    nand3i_3 U139 ( .x(n172), .a(n143), .b(n178), .c(n116) );
    nor2_0 U14 ( .x(n176), .a(A[2]), .b(A[4]) );
    nand2_8 U140 ( .x(n112), .a(n178), .b(n148) );
    inv_0 U141 ( .x(n82), .a(A[5]) );
    oai21_4 U142 ( .x(DIFF[14]), .a(n99), .b(n100), .c(n101) );
    aoai211_4 U143 ( .x(DIFF[20]), .a(n115), .b(n116), .c(n117), .d(n118) );
    nor2i_5 U144 ( .x(n133), .a(n134), .b(n128) );
    nand2_5 U145 ( .x(n128), .a(n156), .b(n157) );
    nor2_5 U146 ( .x(n150), .a(n149), .b(n147) );
    nand2i_4 U147 ( .x(n181), .a(A[2]), .b(n158) );
    nand2i_4 U148 ( .x(n97), .a(A[13]), .b(n116) );
    inv_5 U149 ( .x(n156), .a(n76) );
    nand3i_3 U15 ( .x(n147), .a(A[19]), .b(n117), .c(n148) );
    nand2i_4 U150 ( .x(n129), .a(n157), .b(n76) );
    nand2i_4 U151 ( .x(n77), .a(n159), .b(n126) );
    nand2i_4 U152 ( .x(n122), .a(n163), .b(n119) );
    nand2i_4 U153 ( .x(n120), .a(n164), .b(n153) );
    nand2i_4 U154 ( .x(n98), .a(n165), .b(n96) );
    nand2_6 U155 ( .x(DIFF[26]), .a(n124), .b(n125) );
    nand2_6 U156 ( .x(DIFF[28]), .a(n76), .b(n77) );
    nand2_6 U157 ( .x(DIFF[29]), .a(n128), .b(n129) );
    aoai211_5 U158 ( .x(DIFF[7]), .a(n84), .b(n85), .c(n86), .d(n87) );
    inv_6 U159 ( .x(n94), .a(n93) );
    nor2i_2 U16 ( .x(n177), .a(n109), .b(n54) );
    inv_10 U160 ( .x(n95), .a(A[12]) );
    nand2_8 U161 ( .x(n132), .a(n150), .b(n116) );
    nand2i_6 U162 ( .x(n126), .a(A[27]), .b(n154) );
    nand2i_6 U163 ( .x(n76), .a(A[28]), .b(n155) );
    inv_6 U164 ( .x(n78), .a(n181) );
    inv_6 U165 ( .x(n148), .a(n143) );
    nor2_6 U166 ( .x(n140), .a(A[6]), .b(A[5]) );
    inv_5 U167 ( .x(n81), .a(n80) );
    mux2i_5 U168 ( .x(DIFF[19]), .d0(n137), .sl(n50), .d1(n172) );
    nand2_4 U169 ( .x(n72), .a(n79), .b(n174) );
    mux2_6 U170 ( .x(DIFF[6]), .d0(n60), .sl(n183), .d1(n83) );
    inv_0 U171 ( .x(n183), .a(n67) );
    nand2_1 U172 ( .x(n83), .a(n169), .b(n175) );
    and2_1 U173 ( .x(n60), .a(n176), .b(n175) );
    inv_6 U174 ( .x(n117), .a(A[20]) );
    inv_7 U175 ( .x(n114), .a(A[18]) );
    inv_5 U176 ( .x(n109), .a(A[17]) );
    inv_3 U177 ( .x(n139), .a(A[8]) );
    inv_1 U178 ( .x(n66), .a(A[22]) );
    inv_0 U18 ( .x(n131), .a(A[21]) );
    inv_5 U19 ( .x(n171), .a(n118) );
    inv_5 U20 ( .x(n108), .a(n107) );
    nor2_4 U22 ( .x(n174), .a(A[3]), .b(A[2]) );
    inv_0 U23 ( .x(n161), .a(A[26]) );
    inv_5 U24 ( .x(n154), .a(n124) );
    inv_4 U25 ( .x(n102), .a(n101) );
    oai21_2 U26 ( .x(DIFF[15]), .a(n102), .b(n103), .c(n104) );
    inv_2 U28 ( .x(n99), .a(n97) );
    inv_5 U29 ( .x(n88), .a(n168) );
    ao21_1 U30 ( .x(DIFF[3]), .a(A[3]), .b(A[2]), .c(n78) );
    inv_0 U31 ( .x(DIFF[2]), .a(A[2]) );
    nand2i_2 U32 ( .x(n55), .a(A[25]), .b(n56) );
    inv_4 U33 ( .x(n119), .a(n68) );
    inv_4 U34 ( .x(n113), .a(n110) );
    nor2i_3 U35 ( .x(n68), .a(n164), .b(n153) );
    inv_0 U36 ( .x(n135), .a(A[9]) );
    inv_7 U37 ( .x(n155), .a(n126) );
    oai21_1 U39 ( .x(DIFF[4]), .a(n78), .b(n79), .c(n72) );
    oai21_5 U4 ( .x(DIFF[11]), .a(n92), .b(n75), .c(n93) );
    nand2_3 U40 ( .x(DIFF[13]), .a(n97), .b(n98) );
    inv_7 U41 ( .x(n86), .a(A[7]) );
    exnor2_1 U42 ( .x(DIFF[31]), .a(n133), .b(n167) );
    inv_5 U43 ( .x(n106), .a(A[16]) );
    inv_2 U44 ( .x(n90), .a(A[10]) );
    inv_0 U45 ( .x(n163), .a(A[24]) );
    inv_8 U46 ( .x(n100), .a(A[14]) );
    inv_7 U48 ( .x(n165), .a(A[13]) );
    inv_2 U49 ( .x(n160), .a(A[27]) );
    nand2i_5 U5 ( .x(n151), .a(A[21]), .b(n152) );
    inv_2 U50 ( .x(n159), .a(A[28]) );
    inv_2 U51 ( .x(n157), .a(A[29]) );
    inv_2 U52 ( .x(n167), .a(A[31]) );
    inv_3 U53 ( .x(n75), .a(A[11]) );
    exnor2_5 U54 ( .x(DIFF[30]), .a(n128), .b(n53) );
    buf_1 U55 ( .x(n51), .a(n90) );
    mux2i_3 U56 ( .x(DIFF[21]), .d0(n132), .sl(A[21]), .d1(n171) );
    oai21_5 U57 ( .x(DIFF[16]), .a(n105), .b(n106), .c(n107) );
    nor2_8 U58 ( .x(n145), .a(A[9]), .b(A[10]) );
    nor2_1 U59 ( .x(n175), .a(A[5]), .b(A[3]) );
    inv_10 U6 ( .x(n152), .a(n132) );
    oai21_2 U60 ( .x(DIFF[5]), .a(n81), .b(n82), .c(n83) );
    nand2i_4 U62 ( .x(n141), .a(n72), .b(n142) );
    mux2i_3 U63 ( .x(DIFF[22]), .d0(n130), .sl(n66), .d1(n151) );
    inv_6 U64 ( .x(n105), .a(n104) );
    inv_5 U65 ( .x(n158), .a(A[3]) );
    inv_1 U67 ( .x(n64), .a(n69) );
    inv_1 U68 ( .x(n69), .a(n144) );
    nor3_1 U69 ( .x(n85), .a(A[3]), .b(A[6]), .c(A[5]) );
    nand4i_1 U70 ( .x(n87), .a(A[5]), .b(n173), .c(n174), .d(n79) );
    nor3_5 U71 ( .x(n146), .a(n144), .b(n63), .c(n62) );
    nand2i_3 U72 ( .x(n62), .a(A[2]), .b(n158) );
    nand2_6 U73 ( .x(n101), .a(n73), .b(n116) );
    nand2_6 U74 ( .x(n59), .a(n165), .b(n100) );
    inv_7 U75 ( .x(n73), .a(n59) );
    and4i_1 U76 ( .x(n52), .a(n151), .b(n163), .c(n164), .d(n66) );
    inv_3 U77 ( .x(n121), .a(n52) );
    inv_2 U78 ( .x(n164), .a(A[23]) );
    nor2_3 U79 ( .x(n180), .a(n72), .b(n166) );
    inv_2 U8 ( .x(n50), .a(A[19]) );
    oai21_5 U80 ( .x(DIFF[12]), .a(n94), .b(n95), .c(n96) );
    inv_6 U81 ( .x(n63), .a(n79) );
    nand2_3 U82 ( .x(n80), .a(n79), .b(n174) );
    nand2_6 U83 ( .x(DIFF[27]), .a(n126), .b(n127) );
    nand3_3 U84 ( .x(n93), .a(n142), .b(n75), .c(n180) );
    nand3i_5 U85 ( .x(n144), .a(A[11]), .b(n95), .c(n145) );
    nand3_4 U86 ( .x(n136), .a(n86), .b(n139), .c(n140) );
    nand2i_3 U88 ( .x(n104), .a(n179), .b(n116) );
    inv_2 U89 ( .x(n53), .a(n134) );
    nand2_6 U9 ( .x(DIFF[24]), .a(n121), .b(n122) );
    inv_2 U90 ( .x(n134), .a(A[30]) );
    nor2_2 U91 ( .x(n173), .a(A[7]), .b(A[6]) );
    inv_6 U92 ( .x(n92), .a(n91) );
    nand2i_6 U93 ( .x(n149), .a(n61), .b(n73) );
    nand2i_6 U94 ( .x(n54), .a(n61), .b(n73) );
    inv_16 U95 ( .x(n116), .a(n111) );
    inv_4 U96 ( .x(n182), .a(n141) );
    oai21_2 U97 ( .x(DIFF[10]), .a(n89), .b(n51), .c(n91) );
    nor3i_2 U98 ( .x(n89), .a(n135), .b(n72), .c(n58) );
    oai21_4 U99 ( .x(DIFF[17]), .a(n108), .b(n109), .c(n110) );
endmodule


module ID_DW01_sub_32_1_test_1 ( A, B, CI, DIFF, CO );
input  [31:0] A;
input  [31:0] B;
output [31:0] DIFF;
input  CI;
output CO;
    wire A_1, A_0, n166, n167, n58, n59, n154, n155, n156, n78, n157, n83, n60, 
        n161, n129, n79, n134, n131, n62, n132, n128, n136, n54, n174, n173, 
        n135, n94, n168, n151, n175, n92, n90, n116, n117, n143, n170, n140, 
        n114, n68, n65, n66, n133, n125, n85, n130, n153, n70, n63, n162, n158, 
        n93, n64, n67, n127, n69, n176, n72, n164, n165, n82, n152, n76, n77, 
        n91, n98, n99, n100, n101, n102, n103, n104, n105, n106, n109, n110, 
        n111, n74, n163, n178, n75, n51, n86, n88, n172, n137, n171, n107, 
        n139, n113, n148, n108, n149, n84, n81, n80, n112, n118, n119, n120, 
        n160, n124, n138, n142, n55, n56, n87, n61, n122, n146, n177, n145, 
        n179, n147, n115, n73, n96, n97, n150, n141, n121, n123, n159, n144, 
        n95, n89, n57, n71, n126, n52, n53, n169;
    assign A_1 = A[1];
    assign A_0 = A[0];
    assign DIFF[1] = A_1;
    assign DIFF[0] = A_0;
    nor2_0 U10 ( .x(n166), .a(A[2]), .b(A[3]) );
    nor2_2 U100 ( .x(n167), .a(A[2]), .b(A[3]) );
    and4i_4 U101 ( .x(n58), .a(n59), .b(n154), .c(n155), .d(n156) );
    inv_4 U102 ( .x(n78), .a(n58) );
    inv_2 U103 ( .x(n59), .a(n157) );
    ao21_4 U104 ( .x(DIFF[14]), .a(n83), .b(A[14]), .c(n60) );
    nor2_1 U105 ( .x(n161), .a(A[2]), .b(A[3]) );
    nor2_5 U106 ( .x(n60), .a(n129), .b(n79) );
    inv_10 U107 ( .x(n134), .a(n79) );
    nor2_1 U108 ( .x(n131), .a(A[6]), .b(A[10]) );
    aoi21_1 U109 ( .x(n62), .a(n132), .b(n166), .c(n128) );
    inv_0 U11 ( .x(n136), .a(n54) );
    nand2i_0 U110 ( .x(n174), .a(A[15]), .b(n173) );
    nand3i_1 U111 ( .x(n135), .a(A[15]), .b(n94), .c(n168) );
    inv_0 U112 ( .x(n151), .a(A[15]) );
    nor2_0 U113 ( .x(n175), .a(A[15]), .b(A[16]) );
    nand2_1 U114 ( .x(n92), .a(A[17]), .b(n90) );
    inv_2 U116 ( .x(DIFF[2]), .a(A[2]) );
    nand2_6 U117 ( .x(DIFF[27]), .a(n116), .b(n117) );
    nand2i_6 U118 ( .x(n116), .a(A[27]), .b(n143) );
    nor2_0 U119 ( .x(n170), .a(A[21]), .b(A[20]) );
    nand2i_0 U12 ( .x(n140), .a(A[25]), .b(n114) );
    ao21_1 U120 ( .x(DIFF[3]), .a(A[3]), .b(A[2]), .c(n68) );
    and4i_3 U121 ( .x(n65), .a(n66), .b(n131), .c(n132), .d(n133) );
    nor2_0 U122 ( .x(n125), .a(A[5]), .b(A[6]) );
    nand3i_1 U123 ( .x(n129), .a(A[13]), .b(n85), .c(n130) );
    inv_0 U124 ( .x(n153), .a(A[13]) );
    nand2i_2 U125 ( .x(n70), .a(n63), .b(n161) );
    mux2i_2 U126 ( .x(DIFF[11]), .d0(n162), .sl(A[11]), .d1(n134) );
    nor2_0 U128 ( .x(n173), .a(A[17]), .b(A[16]) );
    inv_0 U129 ( .x(n158), .a(A[10]) );
    oai21_2 U13 ( .x(DIFF[18]), .a(n93), .b(n94), .c(n64) );
    nand2_1 U130 ( .x(n67), .a(n127), .b(n69) );
    inv_2 U131 ( .x(n155), .a(n67) );
    inv_0 U132 ( .x(n176), .a(A[11]) );
    nand2i_2 U133 ( .x(n162), .a(A[10]), .b(n58) );
    nand4i_1 U134 ( .x(n72), .a(A[7]), .b(n164), .c(n165), .d(n69) );
    oai21_1 U135 ( .x(n82), .a(A[11]), .b(n79), .c(A[12]) );
    nand2i_0 U136 ( .x(n152), .a(A[12]), .b(n176) );
    nor2_0 U137 ( .x(n165), .a(A[6]), .b(A[5]) );
    oai21_4 U138 ( .x(DIFF[4]), .a(n68), .b(n69), .c(n70) );
    oai21_4 U139 ( .x(DIFF[9]), .a(n76), .b(n77), .c(n78) );
    inv_2 U14 ( .x(n93), .a(n91) );
    oai21_4 U140 ( .x(DIFF[20]), .a(n98), .b(n99), .c(n100) );
    oai21_4 U141 ( .x(DIFF[21]), .a(n101), .b(n102), .c(n103) );
    oai21_4 U142 ( .x(DIFF[22]), .a(n104), .b(n105), .c(n106) );
    oai21_4 U143 ( .x(DIFF[24]), .a(n109), .b(n110), .c(n111) );
    nand2i_4 U144 ( .x(n74), .a(n163), .b(n178) );
    nand2i_4 U145 ( .x(n75), .a(n51), .b(n72) );
    nand2i_4 U146 ( .x(n86), .a(A[15]), .b(n60) );
    inv_5 U147 ( .x(n88), .a(n86) );
    nand2i_4 U148 ( .x(n91), .a(n174), .b(n60) );
    nand2i_4 U149 ( .x(n100), .a(n172), .b(n137) );
    nand2_2 U15 ( .x(DIFF[17]), .a(n91), .b(n92) );
    nand2i_4 U150 ( .x(n103), .a(n171), .b(n137) );
    nand2i_4 U151 ( .x(n107), .a(A[23]), .b(n139) );
    nand2i_4 U152 ( .x(n113), .a(n148), .b(n111) );
    nand2i_4 U153 ( .x(n108), .a(n149), .b(n106) );
    nand2i_4 U154 ( .x(n84), .a(n153), .b(n81) );
    nand2i_4 U155 ( .x(n80), .a(n158), .b(n78) );
    nand2_5 U156 ( .x(DIFF[23]), .a(n107), .b(n108) );
    nand2_5 U157 ( .x(DIFF[25]), .a(n112), .b(n113) );
    oai21_5 U158 ( .x(DIFF[28]), .a(n118), .b(n119), .c(n120) );
    exnor2_5 U159 ( .x(DIFF[30]), .a(n160), .b(n124) );
    nand2i_2 U16 ( .x(n138), .a(A[23]), .b(n110) );
    nand2i_6 U160 ( .x(n81), .a(n152), .b(n134) );
    nand2i_6 U161 ( .x(n111), .a(n138), .b(n139) );
    nand2i_6 U162 ( .x(n120), .a(n142), .b(n143) );
    mux2i_1 U163 ( .x(n55), .d0(n56), .sl(A[5]), .d1(n70) );
    inv_0 U164 ( .x(n99), .a(A[20]) );
    inv_0 U165 ( .x(n94), .a(A[18]) );
    inv_2 U166 ( .x(n110), .a(A[24]) );
    nor2_1 U167 ( .x(n168), .a(A[17]), .b(A[16]) );
    inv_4 U168 ( .x(n51), .a(A[8]) );
    nand2i_1 U169 ( .x(n163), .a(A[8]), .b(n127) );
    nand2i_2 U17 ( .x(n87), .a(n151), .b(n61) );
    inv_5 U170 ( .x(n105), .a(A[22]) );
    nand2_3 U18 ( .x(DIFF[8]), .a(n74), .b(n75) );
    inv_4 U19 ( .x(n76), .a(n74) );
    nand2i_0 U20 ( .x(n171), .a(A[19]), .b(n170) );
    nand2i_0 U21 ( .x(n172), .a(A[19]), .b(n99) );
    nand2i_2 U23 ( .x(n122), .a(n146), .b(n120) );
    nand2i_2 U24 ( .x(n177), .a(A[2]), .b(n145) );
    inv_5 U25 ( .x(n179), .a(n81) );
    nand2i_2 U26 ( .x(n117), .a(n147), .b(n115) );
    inv_2 U27 ( .x(n118), .a(n116) );
    nand2_2 U28 ( .x(DIFF[7]), .a(n72), .b(n73) );
    nand2i_2 U29 ( .x(n96), .a(A[19]), .b(n137) );
    nand2_2 U30 ( .x(DIFF[19]), .a(n96), .b(n97) );
    nand2i_2 U31 ( .x(n97), .a(n150), .b(n64) );
    inv_2 U32 ( .x(n98), .a(n96) );
    inv_5 U33 ( .x(n141), .a(n111) );
    inv_7 U34 ( .x(n139), .a(n106) );
    nand2_2 U35 ( .x(DIFF[15]), .a(n86), .b(n87) );
    inv_4 U36 ( .x(n68), .a(n177) );
    inv_2 U37 ( .x(n101), .a(n100) );
    inv_0 U38 ( .x(n85), .a(A[14]) );
    inv_2 U39 ( .x(n109), .a(n107) );
    nand2_2 U4 ( .x(DIFF[10]), .a(n80), .b(n79) );
    inv_2 U40 ( .x(n104), .a(n103) );
    nand2_2 U41 ( .x(DIFF[29]), .a(n121), .b(n122) );
    inv_3 U42 ( .x(n127), .a(A[7]) );
    exnor2_1 U43 ( .x(DIFF[31]), .a(n123), .b(n159) );
    nor2i_1 U44 ( .x(n123), .a(n124), .b(n121) );
    inv_2 U45 ( .x(n144), .a(n120) );
    nand2i_2 U46 ( .x(n121), .a(A[29]), .b(n144) );
    inv_2 U47 ( .x(n160), .a(n121) );
    inv_0 U48 ( .x(n114), .a(A[26]) );
    inv_0 U5 ( .x(n150), .a(A[19]) );
    inv_0 U51 ( .x(n148), .a(A[25]) );
    inv_0 U52 ( .x(n102), .a(A[21]) );
    inv_2 U54 ( .x(n149), .a(A[23]) );
    inv_2 U55 ( .x(n147), .a(A[27]) );
    inv_2 U56 ( .x(n119), .a(A[28]) );
    inv_2 U57 ( .x(n146), .a(A[29]) );
    inv_2 U58 ( .x(n124), .a(A[30]) );
    inv_2 U59 ( .x(n159), .a(A[31]) );
    nand2i_2 U6 ( .x(n142), .a(A[27]), .b(n119) );
    inv_4 U60 ( .x(n63), .a(n69) );
    ao21_4 U61 ( .x(DIFF[26]), .a(n112), .b(A[26]), .c(n143) );
    inv_2 U62 ( .x(n61), .a(n60) );
    nand2i_2 U63 ( .x(n64), .a(n135), .b(n60) );
    nand2i_3 U64 ( .x(n95), .a(n135), .b(n60) );
    nand3i_2 U65 ( .x(n90), .a(n129), .b(n175), .c(n134) );
    inv_8 U66 ( .x(n79), .a(n65) );
    oai21_5 U67 ( .x(DIFF[16]), .a(n88), .b(n89), .c(n90) );
    nor2_2 U68 ( .x(n132), .a(A[4]), .b(A[5]) );
    inv_5 U7 ( .x(n69), .a(A[4]) );
    nor2_0 U70 ( .x(n154), .a(A[5]), .b(A[6]) );
    inv_5 U71 ( .x(n143), .a(n115) );
    nand2i_5 U72 ( .x(n112), .a(A[25]), .b(n141) );
    nand2_8 U73 ( .x(DIFF[13]), .a(n83), .b(n84) );
    nand2i_5 U74 ( .x(n83), .a(A[13]), .b(n179) );
    and2_2 U75 ( .x(n156), .a(n77), .b(n51) );
    inv_4 U76 ( .x(n77), .a(A[9]) );
    nor2_5 U77 ( .x(n133), .a(A[2]), .b(A[3]) );
    inv_2 U78 ( .x(n57), .a(n63) );
    inv_3 U79 ( .x(n145), .a(A[3]) );
    nand3_1 U8 ( .x(n71), .a(n69), .b(n125), .c(n126) );
    nor2_1 U80 ( .x(n157), .a(A[2]), .b(A[3]) );
    nor2_1 U81 ( .x(n164), .a(A[2]), .b(A[3]) );
    nand2i_2 U82 ( .x(n73), .a(n127), .b(n71) );
    inv_4 U83 ( .x(n178), .a(n71) );
    inv_0 U84 ( .x(n89), .a(A[16]) );
    or2_6 U85 ( .x(DIFF[6]), .a(n178), .b(n62) );
    nand3_1 U86 ( .x(n66), .a(n127), .b(n51), .c(n77) );
    nand2_3 U87 ( .x(DIFF[12]), .a(n81), .b(n82) );
    nand4i_1 U88 ( .x(n115), .a(n140), .b(n52), .c(n137), .d(n54) );
    inv_2 U89 ( .x(n52), .a(n138) );
    inv_0 U9 ( .x(n128), .a(A[6]) );
    inv_7 U90 ( .x(n137), .a(n95) );
    nor2_3 U91 ( .x(n126), .a(A[2]), .b(A[3]) );
    nand2_8 U92 ( .x(n106), .a(n53), .b(n137) );
    inv_2 U93 ( .x(n53), .a(n136) );
    and3_1 U94 ( .x(n54), .a(n150), .b(n105), .c(n169) );
    nor2_0 U95 ( .x(n169), .a(A[21]), .b(A[20]) );
    nor2_1 U97 ( .x(n130), .a(A[12]), .b(A[11]) );
    inv_5 U98 ( .x(DIFF[5]), .a(n55) );
    and2_5 U99 ( .x(n56), .a(n57), .b(n167) );
endmodule


module ID_DW01_add_32_0_test_1 ( A, B, CI, SUM, CO );
input  [31:0] A;
input  [31:0] B;
output [31:0] SUM;
input  CI;
output CO;
    wire n353, n70, n320, n99, n325, n321, n330, n173, n413, n172, n291, n137, 
        n369, n370, n371, n249, n237, n158, n397, n238, n180, n181, n182, n279, 
        n408, n414, n327, n243, n329, n96, n398, n233, n232, n245, n231, n244, 
        n190, n384, n227, n121, n226, n396, n395, n393, n270, n272, n394, n273, 
        n286, n287, n367, n368, n134, n366, n139, n347, n83, n364, n365, n263, 
        n262, n274, n346, n339, n338, n344, n334, n248, n335, n246, n333, n235, 
        n200, n341, n323, n342, n343, n146, n332, n239, n254, n380, n152, n62, 
        n316, n412, n258, n315, n314, n265, n199, n271, n289, n136, n293, n135, 
        n372, n373, n234, n355, n125, n351, n264, n277, n356, n357, n358, n282, 
        n124, n406, n285, n119, n348, n196, n281, n354, n108, n225, n165, n164, 
        n283, n116, n378, n167, n115, n247, n170, n420, n111, n252, n213, n129, 
        n131, n205, n98, n322, n391, n390, n102, n100, n269, n382, n85, n86, 
        n69, n88, n308, n381, n123, n130, n132, n127, n51, n95, n97, n110, 
        n166, n192, n193, n113, n169, n109, n219, n154, n295, n401, n155, n156, 
        n78, n52, n203, n422, n421, n77, n305, n216, n145, n301, n259, n376, 
        n410, n147, n204, n93, n94, n92, n241, n66, n151, n73, n74, n299, n153, 
        n240, n168, n214, n133, n82, n84, n159, n220, n157, n400, n221, n399, 
        n256, n253, n257, n208, n212, n59, n107, n91, n222, n171, n120, n387, 
        n149, n122, n297, n298, n426, n148, n217, n176, n175, n150, n385, n303, 
        n81, n142, n141, n229, n224, n223, n106, n76, n215, n138, n140, n174, 
        n389, n104, n105, n383, n250, n317, n392, n319, n304, n290, n53, n195, 
        n71, n72, n54, n63, n191, n178, n126, n128, n407, n55, n112, n56, n186, 
        n187, n188, n57, n68, n403, n296, n179, n177, n64, n202, n160, n161, 
        n162, n75, n306, n58, n292, n87, n61, n117, n209, n206, n60, n345, n67, 
        n424, n207, n388, n218, n402, n379, n326, n114, n374, n65, n211, n411, 
        n419, n276, n251, n415, n331, n101, n103, n118, n201, n163, n189, n194, 
        n197, n198, n242, n266, n278, n307, n309, n310, n284, n324, n328, n336, 
        n337, n340, n352, n184, n261, n362, n185, n363, n236, n375, n405, n409, 
        n267, n417, n416, n349, n418, n288, n90, n302, n89, n311, n79, n313, 
        n80, n275, n228, n294, n386, n210, n423, n425, n183, n404, n350, n280, 
        n312, n318, n268, n361, n50, n49, n359, n360, n260, n230, n300, n144, 
        n143, n377, n255;
    nand2_2 U10 ( .x(n353), .a(B[30]), .b(n70) );
    inv_2 U100 ( .x(n320), .a(n99) );
    nand2i_2 U101 ( .x(n325), .a(n320), .b(n321) );
    nand2i_2 U102 ( .x(n330), .a(n173), .b(n413) );
    nand2_0 U103 ( .x(n172), .a(A[10]), .b(B[10]) );
    inv_2 U104 ( .x(n291), .a(n137) );
    nand2i_2 U105 ( .x(n369), .a(n370), .b(n371) );
    nand2i_3 U106 ( .x(n249), .a(A[15]), .b(n237) );
    nand2_0 U107 ( .x(n158), .a(B[15]), .b(A[15]) );
    nand2i_2 U108 ( .x(n397), .a(A[14]), .b(n238) );
    nor2i_1 U109 ( .x(n180), .a(n181), .b(n182) );
    nand2i_2 U11 ( .x(n279), .a(n70), .b(n408) );
    inv_5 U110 ( .x(n182), .a(n414) );
    nand2i_2 U111 ( .x(n327), .a(B[10]), .b(n243) );
    inv_2 U112 ( .x(n329), .a(n172) );
    nand2_2 U113 ( .x(n96), .a(A[8]), .b(B[8]) );
    ao21_1 U114 ( .x(n398), .a(n233), .b(n232), .c(n96) );
    nand2i_2 U115 ( .x(n245), .a(B[8]), .b(n231) );
    nand2i_2 U116 ( .x(n244), .a(n190), .b(n245) );
    nand2i_2 U117 ( .x(n384), .a(B[3]), .b(n227) );
    inv_1 U118 ( .x(n227), .a(A[3]) );
    nand2_0 U119 ( .x(n121), .a(A[3]), .b(B[3]) );
    nand2_2 U12 ( .x(n408), .a(B[27]), .b(B[26]) );
    inv_2 U120 ( .x(n226), .a(B[2]) );
    inv_5 U121 ( .x(n396), .a(n395) );
    nand2_2 U122 ( .x(n393), .a(B[25]), .b(n70) );
    inv_5 U123 ( .x(n270), .a(B[25]) );
    inv_2 U124 ( .x(n272), .a(B[24]) );
    nand2i_2 U125 ( .x(n394), .a(B[24]), .b(n273) );
    nand2_2 U126 ( .x(n371), .a(n286), .b(n287) );
    inv_2 U127 ( .x(n367), .a(n371) );
    inv_2 U128 ( .x(n368), .a(n134) );
    nor2i_1 U129 ( .x(n366), .a(n139), .b(n368) );
    nand2_0 U13 ( .x(n347), .a(B[27]), .b(B[26]) );
    nor2i_1 U130 ( .x(n83), .a(n366), .b(n367) );
    nand2_2 U131 ( .x(n364), .a(n365), .b(n263) );
    nand2i_2 U132 ( .x(n262), .a(A[21]), .b(n274) );
    inv_2 U133 ( .x(n274), .a(B[21]) );
    nand2_2 U134 ( .x(n137), .a(B[21]), .b(A[21]) );
    oai31_2 U135 ( .x(n346), .a(n339), .b(n182), .c(n338), .d(n344) );
    inv_7 U136 ( .x(n334), .a(n248) );
    inv_5 U137 ( .x(n335), .a(n246) );
    nand2_2 U138 ( .x(n333), .a(n334), .b(n335) );
    inv_2 U139 ( .x(n235), .a(A[20]) );
    nor2_1 U14 ( .x(n200), .a(A[22]), .b(B[22]) );
    aoi21_1 U140 ( .x(n341), .a(n323), .b(n342), .c(n343) );
    inv_2 U141 ( .x(n343), .a(n146) );
    inv_5 U142 ( .x(n332), .a(n239) );
    inv_2 U143 ( .x(n254), .a(B[17]) );
    inv_2 U144 ( .x(n380), .a(n152) );
    nand2_2 U145 ( .x(n152), .a(n62), .b(A[17]) );
    inv_1 U146 ( .x(n316), .a(n412) );
    inv_2 U147 ( .x(n258), .a(A[18]) );
    nor2i_1 U148 ( .x(n315), .a(n152), .b(n258) );
    nor2i_1 U149 ( .x(n314), .a(n315), .b(n316) );
    nor2_4 U15 ( .x(n265), .a(n199), .b(n200) );
    inv_2 U150 ( .x(n271), .a(B[23]) );
    inv_2 U151 ( .x(n370), .a(n139) );
    nand2_2 U152 ( .x(n139), .a(A[23]), .b(B[23]) );
    inv_2 U153 ( .x(n365), .a(n289) );
    nand2i_2 U154 ( .x(n289), .a(n136), .b(n262) );
    inv_2 U155 ( .x(n136), .a(n293) );
    nor2_1 U156 ( .x(n135), .a(n136), .b(n137) );
    nor2i_1 U157 ( .x(n372), .a(n373), .b(n135) );
    inv_2 U158 ( .x(n234), .a(B[30]) );
    nand2i_0 U159 ( .x(n355), .a(n125), .b(n351) );
    nand2i_4 U16 ( .x(n264), .a(B[24]), .b(n273) );
    inv_5 U160 ( .x(n351), .a(n277) );
    nor2i_1 U161 ( .x(n356), .a(n357), .b(n358) );
    inv_2 U162 ( .x(n357), .a(n282) );
    inv_2 U163 ( .x(n358), .a(n124) );
    inv_2 U164 ( .x(n406), .a(n285) );
    oai211_1 U165 ( .x(n119), .a(n348), .b(n196), .c(n281), .d(n354) );
    nand2_2 U166 ( .x(n108), .a(B[4]), .b(A[4]) );
    inv_2 U167 ( .x(n225), .a(B[4]) );
    inv_2 U168 ( .x(n165), .a(n181) );
    nand2_2 U169 ( .x(n164), .a(A[13]), .b(B[13]) );
    nand2_0 U17 ( .x(n283), .a(B[28]), .b(n70) );
    nand2i_0 U170 ( .x(n116), .a(n378), .b(n167) );
    nor2_0 U171 ( .x(n115), .a(n247), .b(n170) );
    inv_4 U172 ( .x(n247), .a(n420) );
    nand2i_2 U173 ( .x(n111), .a(B[11]), .b(n252) );
    exor2_1 U174 ( .x(n213), .a(B[27]), .b(n70) );
    inv_2 U175 ( .x(n129), .a(n131) );
    exor2_1 U176 ( .x(SUM[7]), .a(n205), .b(n98) );
    ao21_1 U177 ( .x(n205), .a(n322), .b(n391), .c(n390) );
    inv_2 U178 ( .x(n390), .a(n102) );
    nor2i_1 U179 ( .x(n98), .a(n99), .b(n100) );
    inv_5 U18 ( .x(n269), .a(B[28]) );
    inv_2 U180 ( .x(n100), .a(n382) );
    aoi21_1 U181 ( .x(n85), .a(n86), .b(n69), .c(n88) );
    exnor2_1 U182 ( .x(n308), .a(B[29]), .b(n70) );
    inv_2 U183 ( .x(n125), .a(n381) );
    nor2i_1 U184 ( .x(n123), .a(n124), .b(n125) );
    nor2i_1 U185 ( .x(n130), .a(n131), .b(n132) );
    inv_2 U186 ( .x(n132), .a(n127) );
    exnor2_1 U187 ( .x(SUM[8]), .a(n51), .b(n95) );
    nor2i_1 U188 ( .x(n95), .a(n96), .b(n97) );
    exnor2_1 U189 ( .x(SUM[12]), .a(n110), .b(n166) );
    nor2i_1 U19 ( .x(n192), .a(n137), .b(n193) );
    inv_2 U190 ( .x(n113), .a(n169) );
    nor2i_1 U191 ( .x(n166), .a(n167), .b(n109) );
    exor2_1 U192 ( .x(SUM[16]), .a(n219), .b(n154) );
    nand2i_2 U193 ( .x(n219), .a(n295), .b(n401) );
    nor2i_1 U194 ( .x(n154), .a(n155), .b(n156) );
    nand2i_2 U195 ( .x(n78), .a(n52), .b(n203) );
    inv_2 U196 ( .x(n422), .a(n421) );
    mux2i_1 U197 ( .x(n77), .d0(n422), .sl(A[19]), .d1(n305) );
    nand2_2 U198 ( .x(SUM[19]), .a(n77), .b(n78) );
    exor2_1 U199 ( .x(SUM[20]), .a(n216), .b(n145) );
    nand2i_2 U20 ( .x(n301), .a(A[18]), .b(n259) );
    nand2i_2 U200 ( .x(n216), .a(n376), .b(n410) );
    nor2i_1 U201 ( .x(n145), .a(n146), .b(n147) );
    inv_5 U202 ( .x(n147), .a(n342) );
    exor2_1 U203 ( .x(SUM[9]), .a(n204), .b(n93) );
    oai21_1 U204 ( .x(n204), .a(n51), .b(n97), .c(n96) );
    inv_2 U205 ( .x(n97), .a(n245) );
    nor2i_1 U206 ( .x(n93), .a(n94), .b(n92) );
    inv_2 U207 ( .x(n156), .a(n241) );
    exor2_1 U208 ( .x(SUM[17]), .a(n66), .b(n151) );
    nor2i_1 U209 ( .x(SUM[0]), .a(n73), .b(n74) );
    nor3_0 U21 ( .x(n299), .a(n153), .b(n156), .c(n240) );
    nand2_2 U210 ( .x(n73), .a(B[0]), .b(A[0]) );
    nor2i_1 U211 ( .x(n168), .a(n169), .b(n170) );
    inv_2 U212 ( .x(n170), .a(n111) );
    exor2_1 U213 ( .x(SUM[24]), .a(n214), .b(n133) );
    nand2i_2 U214 ( .x(n214), .a(n369), .b(n82) );
    nor2i_1 U215 ( .x(n133), .a(n134), .b(n84) );
    inv_2 U216 ( .x(n159), .a(n249) );
    exor2_1 U217 ( .x(SUM[15]), .a(n220), .b(n157) );
    inv_2 U218 ( .x(n400), .a(n221) );
    nand2i_2 U219 ( .x(n221), .a(n180), .b(n399) );
    ao221_2 U22 ( .x(n256), .a(n254), .b(n253), .c(n155), .d(n257), .e(n240)
         );
    ao21_3 U220 ( .x(n208), .a(n384), .b(n212), .c(n59) );
    nor2i_1 U221 ( .x(n107), .a(n108), .b(n91) );
    exor2_1 U222 ( .x(SUM[10]), .a(n222), .b(n171) );
    oai211_1 U223 ( .x(n222), .a(n51), .b(n244), .c(n398), .d(n94) );
    nor2i_1 U224 ( .x(n171), .a(n172), .b(n173) );
    inv_2 U225 ( .x(n173), .a(n327) );
    exor2_1 U226 ( .x(SUM[3]), .a(n212), .b(n120) );
    inv_2 U227 ( .x(n387), .a(n149) );
    nor2i_1 U228 ( .x(n120), .a(n121), .b(n122) );
    inv_2 U229 ( .x(n122), .a(n384) );
    nand2i_0 U23 ( .x(n297), .a(n298), .b(n256) );
    exor2_1 U230 ( .x(SUM[2]), .a(n426), .b(n148) );
    oai21_2 U231 ( .x(n217), .a(n176), .b(n73), .c(n175) );
    nor2i_1 U232 ( .x(n148), .a(n149), .b(n150) );
    inv_2 U233 ( .x(n150), .a(n385) );
    nand2i_2 U234 ( .x(n303), .a(n396), .b(n393) );
    inv_2 U235 ( .x(n84), .a(n394) );
    aoi21_1 U236 ( .x(n81), .a(n82), .b(n83), .c(n84) );
    exnor2_1 U237 ( .x(SUM[25]), .a(n81), .b(n303) );
    inv_2 U238 ( .x(n142), .a(n262) );
    nor2i_1 U239 ( .x(n141), .a(n137), .b(n142) );
    ao21_2 U24 ( .x(n229), .a(n224), .b(n223), .c(n106) );
    exor2_1 U240 ( .x(SUM[21]), .a(n69), .b(n141) );
    ao21_1 U241 ( .x(n76), .a(n152), .b(n412), .c(n301) );
    exor2_1 U242 ( .x(SUM[23]), .a(n215), .b(n138) );
    nor2i_1 U243 ( .x(n138), .a(n139), .b(n140) );
    exnor2_1 U244 ( .x(SUM[1]), .a(n174), .b(n73) );
    nor2i_0 U245 ( .x(n174), .a(n175), .b(n176) );
    inv_5 U247 ( .x(n106), .a(n389) );
    nor2i_0 U248 ( .x(n104), .a(n105), .b(n106) );
    inv_2 U249 ( .x(n383), .a(n108) );
    nand2_1 U25 ( .x(n94), .a(A[9]), .b(B[9]) );
    inv_0 U250 ( .x(n250), .a(A[12]) );
    aoi21_1 U251 ( .x(n51), .a(n317), .b(n392), .c(n319) );
    exnor2_3 U253 ( .x(n304), .a(n290), .b(n53) );
    inv_2 U254 ( .x(n53), .a(n195) );
    inv_2 U255 ( .x(n195), .a(B[22]) );
    inv_2 U256 ( .x(n71), .a(A[31]) );
    inv_2 U257 ( .x(n72), .a(A[31]) );
    buf_1 U258 ( .x(n54), .a(n63) );
    nand2_1 U259 ( .x(n146), .a(B[20]), .b(A[20]) );
    nor2_1 U26 ( .x(n191), .a(B[9]), .b(A[9]) );
    inv_0 U260 ( .x(n178), .a(B[5]) );
    exnor2_3 U261 ( .x(SUM[27]), .a(n126), .b(n213) );
    aoi21_3 U262 ( .x(n126), .a(n127), .b(n128), .c(n129) );
    inv_2 U263 ( .x(n407), .a(n128) );
    exor2_1 U264 ( .x(SUM[26]), .a(n128), .b(n130) );
    inv_0 U265 ( .x(n55), .a(n112) );
    inv_2 U266 ( .x(n56), .a(n55) );
    aoi31_6 U267 ( .x(n186), .a(n63), .b(n108), .c(n187), .d(n188) );
    nand2i_2 U268 ( .x(n293), .a(A[22]), .b(n195) );
    nand2_0 U269 ( .x(n373), .a(A[22]), .b(B[22]) );
    oai21_1 U27 ( .x(n413), .a(n191), .b(n96), .c(n94) );
    nor2i_2 U270 ( .x(n193), .a(A[22]), .b(n195) );
    and3i_1 U271 ( .x(n57), .a(n346), .b(n68), .c(n403) );
    oa31_4 U272 ( .x(n68), .a(n239), .b(n147), .c(n296), .d(n341) );
    nand3i_0 U273 ( .x(n392), .a(n179), .b(n108), .c(n63) );
    nand3i_0 U274 ( .x(n391), .a(n177), .b(n108), .c(n54) );
    oai21_5 U275 ( .x(n63), .a(A[4]), .b(n64), .c(n208) );
    nand2_1 U276 ( .x(n202), .a(B[18]), .b(A[18]) );
    nor2i_0 U277 ( .x(n160), .a(n161), .b(n162) );
    oai21_1 U278 ( .x(n220), .a(n162), .b(n400), .c(n161) );
    mux2i_2 U279 ( .x(n75), .d0(n306), .sl(n58), .d1(n314) );
    nand2i_2 U28 ( .x(n292), .a(n142), .b(n87) );
    inv_2 U280 ( .x(n58), .a(n61) );
    inv_2 U281 ( .x(n87), .a(n57) );
    nand2i_4 U282 ( .x(n420), .a(B[12]), .b(n250) );
    nor2_0 U283 ( .x(n109), .a(B[12]), .b(A[12]) );
    inv_2 U284 ( .x(n238), .a(B[14]) );
    nand2_2 U285 ( .x(n161), .a(B[14]), .b(A[14]) );
    exnor2_5 U286 ( .x(SUM[31]), .a(n117), .b(n209) );
    aoai211_1 U287 ( .x(n206), .a(n108), .b(n54), .c(n106), .d(n105) );
    inv_2 U288 ( .x(n59), .a(n121) );
    inv_0 U289 ( .x(n60), .a(A[11]) );
    inv_4 U29 ( .x(n345), .a(n256) );
    and3i_3 U290 ( .x(n67), .a(n346), .b(n68), .c(n403) );
    mux2i_1 U291 ( .x(SUM[29]), .d0(n123), .sl(n85), .d1(n308) );
    exor2_1 U292 ( .x(SUM[4]), .a(n424), .b(n107) );
    ao21_1 U293 ( .x(n207), .a(n388), .b(n424), .c(n383) );
    inv_0 U294 ( .x(n61), .a(n259) );
    buf_1 U295 ( .x(n62), .a(B[17]) );
    nand2i_4 U296 ( .x(n412), .a(n153), .b(n218) );
    inv_2 U297 ( .x(n153), .a(n402) );
    oai21_4 U298 ( .x(n379), .a(n186), .b(n325), .c(n326) );
    nand2i_3 U299 ( .x(n382), .a(A[7]), .b(n224) );
    inv_4 U30 ( .x(n259), .a(B[18]) );
    inv_0 U300 ( .x(n223), .a(A[7]) );
    inv_0 U301 ( .x(n231), .a(A[8]) );
    inv_2 U302 ( .x(n64), .a(n225) );
    exor2_1 U303 ( .x(SUM[11]), .a(n56), .b(n168) );
    aoi21_1 U304 ( .x(n110), .a(n111), .b(n56), .c(n113) );
    aoi21_1 U305 ( .x(n114), .a(n115), .b(n56), .c(n116) );
    nand2i_2 U306 ( .x(n399), .a(n246), .b(n112) );
    nand2i_4 U307 ( .x(n112), .a(n374), .b(n379) );
    inv_0 U308 ( .x(n243), .a(A[10]) );
    nand2_2 U31 ( .x(n257), .a(B[17]), .b(A[17]) );
    inv_2 U310 ( .x(n65), .a(n211) );
    exor2_1 U312 ( .x(n211), .a(B[30]), .b(n70) );
    aoai211_1 U313 ( .x(n66), .a(n411), .b(n401), .c(n156), .d(n155) );
    nand2i_2 U314 ( .x(n419), .a(A[24]), .b(n272) );
    nand2_1 U315 ( .x(n276), .a(A[24]), .b(B[24]) );
    nand2_0 U316 ( .x(n134), .a(A[24]), .b(B[24]) );
    inv_0 U317 ( .x(n273), .a(A[24]) );
    nand2_2 U318 ( .x(n187), .a(A[5]), .b(B[5]) );
    nor2i_0 U319 ( .x(n179), .a(A[5]), .b(n178) );
    inv_2 U32 ( .x(n253), .a(A[17]) );
    nor2i_0 U320 ( .x(n177), .a(A[5]), .b(n178) );
    nand2_0 U321 ( .x(n105), .a(A[5]), .b(B[5]) );
    nor2_0 U322 ( .x(n74), .a(A[0]), .b(B[0]) );
    inv_0 U323 ( .x(n251), .a(A[13]) );
    inv_0 U324 ( .x(n233), .a(A[9]) );
    nor2_1 U325 ( .x(n190), .a(B[9]), .b(A[9]) );
    nor2_0 U326 ( .x(n92), .a(B[9]), .b(A[9]) );
    inv_10 U327 ( .x(n69), .a(n67) );
    or3i_5 U328 ( .x(n403), .a(n415), .b(n333), .c(n331) );
    nand3i_2 U329 ( .x(n321), .a(n100), .b(A[6]), .c(B[6]) );
    inv_2 U33 ( .x(n298), .a(n202) );
    nand2_0 U330 ( .x(n102), .a(A[6]), .b(B[6]) );
    inv_0 U331 ( .x(n252), .a(A[11]) );
    nand2i_0 U332 ( .x(n388), .a(A[4]), .b(n225) );
    nor2_0 U333 ( .x(n91), .a(A[4]), .b(B[4]) );
    nand2i_2 U334 ( .x(n385), .a(A[2]), .b(n226) );
    nand2_2 U335 ( .x(n149), .a(B[2]), .b(A[2]) );
    nand2_2 U336 ( .x(n175), .a(A[1]), .b(B[1]) );
    inv_16 U337 ( .x(n70), .a(n71) );
    nor2i_5 U338 ( .x(n101), .a(n102), .b(n103) );
    aoi21_3 U339 ( .x(n117), .a(n118), .b(n69), .c(n119) );
    nor3_2 U34 ( .x(n201), .a(n147), .b(n202), .c(n203) );
    nor2i_5 U340 ( .x(n151), .a(n152), .b(n153) );
    nor2i_5 U341 ( .x(n163), .a(n164), .b(n165) );
    nor2_5 U342 ( .x(n189), .a(A[19]), .b(B[19]) );
    nor2_5 U343 ( .x(n194), .a(A[17]), .b(B[17]) );
    nor2_5 U344 ( .x(n196), .a(n197), .b(n198) );
    exor2_3 U345 ( .x(SUM[6]), .a(n206), .b(n101) );
    exor2_3 U346 ( .x(SUM[5]), .a(n207), .b(n104) );
    exor2_3 U347 ( .x(SUM[14]), .a(n221), .b(n160) );
    exnor2_5 U348 ( .x(SUM[13]), .a(n114), .b(n163) );
    inv_6 U349 ( .x(n237), .a(B[15]) );
    nand2_2 U35 ( .x(n167), .a(A[12]), .b(B[12]) );
    nand3i_5 U350 ( .x(n239), .a(n240), .b(n241), .c(n242) );
    ao21_4 U351 ( .x(n266), .a(n72), .b(n234), .c(n125) );
    oai211_4 U352 ( .x(n198), .a(n71), .b(n270), .c(n139), .d(n276) );
    nand2i_4 U353 ( .x(n277), .a(n278), .b(n279) );
    nand2i_4 U354 ( .x(n290), .a(n291), .b(n292) );
    exnor2_3 U355 ( .x(n306), .a(A[18]), .b(n307) );
    nor2i_5 U356 ( .x(n309), .a(n310), .b(n284) );
    nand2i_4 U358 ( .x(n188), .a(n103), .b(n324) );
    nor2i_5 U359 ( .x(n326), .a(n327), .b(n244) );
    nand2i_2 U36 ( .x(n328), .a(n329), .b(n330) );
    nand2i_4 U360 ( .x(n331), .a(n147), .b(n332) );
    nor2i_5 U361 ( .x(n336), .a(n167), .b(n337) );
    nand2_5 U362 ( .x(n339), .a(n334), .b(n332) );
    nor2_5 U363 ( .x(n340), .a(n147), .b(n203) );
    aoi21_3 U364 ( .x(n344), .a(n340), .b(n345), .c(n201) );
    nor2i_5 U365 ( .x(n118), .a(n86), .b(n266) );
    nand2_2 U366 ( .x(n352), .a(n353), .b(n283) );
    nor2_5 U367 ( .x(n184), .a(n261), .b(n362) );
    oai21_5 U368 ( .x(n185), .a(n362), .b(n285), .c(n363) );
    nand2i_4 U369 ( .x(n374), .a(n329), .b(n330) );
    inv_2 U37 ( .x(n236), .a(A[19]) );
    nand2_5 U370 ( .x(n375), .a(n335), .b(n334) );
    ao21_4 U371 ( .x(n212), .a(n217), .b(n385), .c(n387) );
    nand2i_4 U372 ( .x(n395), .a(n70), .b(n270) );
    inv_5 U373 ( .x(n337), .a(n164) );
    nand2i_4 U374 ( .x(n128), .a(n406), .b(n405) );
    nand2_2 U375 ( .x(n215), .a(n372), .b(n409) );
    nand2i_4 U376 ( .x(n414), .a(n378), .b(n336) );
    inv_5 U377 ( .x(n86), .a(n267) );
    nand2i_4 U378 ( .x(n417), .a(n169), .b(n416) );
    inv_5 U379 ( .x(n378), .a(n417) );
    nor2i_0 U38 ( .x(n323), .a(B[19]), .b(n236) );
    oai21_4 U380 ( .x(n349), .a(n396), .b(n418), .c(n393) );
    nand2i_4 U381 ( .x(n415), .a(n328), .b(n379) );
    nand2i_4 U382 ( .x(n307), .a(n380), .b(n412) );
    oai21_4 U383 ( .x(n288), .a(n396), .b(n418), .c(n393) );
    inv_5 U384 ( .x(n411), .a(n295) );
    nand2i_4 U385 ( .x(n90), .a(n269), .b(n302) );
    mux2i_3 U387 ( .x(n89), .d0(n309), .sl(n407), .d1(n311) );
    mux2i_3 U388 ( .x(n79), .d0(n313), .sl(A[22]), .d1(n304) );
    nand2_3 U389 ( .x(SUM[18]), .a(n75), .b(n76) );
    nor2_3 U39 ( .x(n242), .a(n189), .b(n194) );
    nand2_3 U390 ( .x(SUM[22]), .a(n79), .b(n80) );
    nand2_3 U391 ( .x(SUM[28]), .a(n89), .b(n90) );
    exor2_5 U392 ( .x(n209), .a(B[31]), .b(n70) );
    inv_6 U393 ( .x(n162), .a(n397) );
    nand2i_4 U394 ( .x(n409), .a(n289), .b(n69) );
    nand2i_5 U395 ( .x(n82), .a(n364), .b(n69) );
    aoai211_5 U397 ( .x(n285), .a(n286), .b(n287), .c(n198), .d(n288) );
    nand2i_6 U398 ( .x(n181), .a(B[13]), .b(n251) );
    nand3i_4 U399 ( .x(n246), .a(n247), .b(n111), .c(n181) );
    nand2i_5 U400 ( .x(n342), .a(B[20]), .b(n235) );
    nand2i_4 U401 ( .x(n338), .a(n147), .b(n181) );
    nand2i_5 U402 ( .x(n263), .a(A[23]), .b(n271) );
    nand4_5 U403 ( .x(n261), .a(n262), .b(n263), .c(n264), .d(n265) );
    nand2i_6 U404 ( .x(n284), .a(n70), .b(n269) );
    nand2i_5 U405 ( .x(n381), .a(B[29]), .b(n72) );
    inv_7 U406 ( .x(n286), .a(n275) );
    nand2i_5 U407 ( .x(n389), .a(B[5]), .b(n228) );
    inv_6 U408 ( .x(n240), .a(n301) );
    inv_6 U409 ( .x(n418), .a(n419) );
    inv_2 U41 ( .x(n296), .a(n294) );
    nor2_8 U410 ( .x(n199), .a(n70), .b(B[25]) );
    or2_6 U411 ( .x(n386), .a(B[1]), .b(A[1]) );
    nand2i_8 U412 ( .x(n405), .a(n261), .b(n69) );
    exnor2_5 U413 ( .x(SUM[30]), .a(n210), .b(n65) );
    aoai211_4 U414 ( .x(n218), .a(n411), .b(n401), .c(n156), .d(n155) );
    aoai211_3 U415 ( .x(n210), .a(n285), .b(n405), .c(n355), .d(n356) );
    nand2i_5 U416 ( .x(n401), .a(n375), .b(n112) );
    nor2i_2 U417 ( .x(n313), .a(B[22]), .b(n290) );
    nand2i_2 U418 ( .x(n80), .a(n293), .b(n290) );
    inv_3 U419 ( .x(n176), .a(n386) );
    oai31_2 U42 ( .x(n295), .a(n182), .b(n165), .c(n248), .d(n296) );
    inv_0 U420 ( .x(n423), .a(n208) );
    inv_2 U421 ( .x(n424), .a(n423) );
    inv_0 U422 ( .x(n425), .a(n217) );
    inv_2 U423 ( .x(n426), .a(n425) );
    inv_0 U44 ( .x(n140), .a(n263) );
    nor2_2 U45 ( .x(n183), .a(A[22]), .b(B[22]) );
    nand2i_2 U46 ( .x(n275), .a(n183), .b(n263) );
    nand2_0 U47 ( .x(n404), .a(A[22]), .b(B[22]) );
    nand2_2 U48 ( .x(n287), .a(n404), .b(n137) );
    and3i_1 U49 ( .x(n354), .a(n352), .b(n131), .c(n124) );
    nor2i_0 U5 ( .x(n157), .a(n158), .b(n159) );
    nand2_2 U50 ( .x(n131), .a(B[26]), .b(n70) );
    nand2_0 U51 ( .x(n124), .a(B[29]), .b(n70) );
    nand2_2 U52 ( .x(n281), .a(B[27]), .b(n70) );
    nand3_1 U53 ( .x(n348), .a(n349), .b(n350), .c(n351) );
    inv_4 U54 ( .x(n350), .a(n266) );
    nand2i_2 U55 ( .x(n416), .a(B[12]), .b(n250) );
    inv_2 U56 ( .x(n363), .a(n280) );
    nand2i_0 U57 ( .x(n312), .a(B[28]), .b(n70) );
    nand2_2 U58 ( .x(n280), .a(n281), .b(n131) );
    nor2_1 U59 ( .x(n311), .a(n280), .b(n312) );
    oai21_1 U6 ( .x(n294), .a(n159), .b(n161), .c(n158) );
    inv_2 U60 ( .x(n362), .a(n310) );
    nand2_2 U61 ( .x(n310), .a(n408), .b(n72) );
    nor2_0 U62 ( .x(n322), .a(n106), .b(n103) );
    inv_2 U63 ( .x(n228), .a(A[5]) );
    inv_3 U64 ( .x(n103), .a(n318) );
    inv_2 U65 ( .x(n278), .a(n284) );
    aoi21_1 U66 ( .x(n268), .a(n347), .b(n72), .c(n278) );
    nand2i_2 U67 ( .x(n267), .a(n261), .b(n268) );
    inv_2 U68 ( .x(n197), .a(n361) );
    nand2i_2 U69 ( .x(n282), .a(n280), .b(n283) );
    exnor2_2 U7 ( .x(n302), .a(n50), .b(n49) );
    nand2_2 U70 ( .x(n359), .a(n349), .b(n351) );
    nand2i_2 U71 ( .x(n361), .a(n192), .b(n286) );
    inv_2 U72 ( .x(n360), .a(n198) );
    aoai211_1 U73 ( .x(n88), .a(n360), .b(n361), .c(n359), .d(n357) );
    nand2i_2 U74 ( .x(n127), .a(n70), .b(n260) );
    inv_2 U75 ( .x(n260), .a(B[26]) );
    nand2i_0 U76 ( .x(n319), .a(n320), .b(n321) );
    nand2_0 U77 ( .x(n99), .a(B[7]), .b(A[7]) );
    nor2i_0 U78 ( .x(n317), .a(n318), .b(n229) );
    nand2i_2 U79 ( .x(n318), .a(B[6]), .b(n230) );
    inv_2 U8 ( .x(n49), .a(n71) );
    inv_0 U80 ( .x(n230), .a(A[6]) );
    inv_2 U81 ( .x(n224), .a(B[7]) );
    inv_2 U82 ( .x(n324), .a(n229) );
    inv_4 U83 ( .x(n203), .a(n300) );
    nand2i_2 U84 ( .x(n300), .a(A[19]), .b(n144) );
    nand2i_2 U85 ( .x(n421), .a(n144), .b(n52) );
    aoi21_1 U86 ( .x(n52), .a(n219), .b(n299), .c(n297) );
    exnor2_1 U87 ( .x(n305), .a(n52), .b(n144) );
    inv_5 U88 ( .x(n144), .a(B[19]) );
    nand2i_0 U89 ( .x(n410), .a(n239), .b(n219) );
    ao21_3 U9 ( .x(n50), .a(n184), .b(n69), .c(n185) );
    nand2i_2 U90 ( .x(n376), .a(n143), .b(n377) );
    nor2i_1 U91 ( .x(n143), .a(A[19]), .b(n144) );
    nand2i_2 U92 ( .x(n377), .a(n203), .b(n297) );
    inv_0 U93 ( .x(n232), .a(B[9]) );
    nand2i_2 U94 ( .x(n402), .a(A[17]), .b(n254) );
    inv_2 U95 ( .x(n255), .a(A[16]) );
    nand2i_2 U96 ( .x(n241), .a(B[16]), .b(n255) );
    nand2i_4 U97 ( .x(n248), .a(n162), .b(n249) );
    nand2_2 U98 ( .x(n155), .a(A[16]), .b(B[16]) );
    nand2i_2 U99 ( .x(n169), .a(n60), .b(B[11]) );
endmodule


module ID_DW01_add_32_2_test_1 ( A, B, CI, SUM, CO );
input  [31:0] A;
input  [31:0] B;
output [31:0] SUM;
input  CI;
output CO;
    wire n183, n158, n83, n160, n174, ___cell__37600_net131624, 
        ___cell__37600_net131625, n103, ___cell__37600_net131609, 
        ___cell__37600_net131611, ___cell__37600_net131612, 
        ___cell__37600_net131608, ___cell__37600_net131586, 
        ___cell__37600_net131802, ___cell__37600_net131575, n215, net152417, 
        ___cell__37600_net131806, n140, ___cell__37600_net131584, 
        ___cell__37600_net131756, n204, n137, n157, n210, net149842, 
        ___cell__37600_net131585, ___cell__37600_net131640, net148303, n141, 
        ___cell__37600_net131645, ___cell__37600_net131506, 
        ___cell__37600_net131507, ___cell__37600_net131508, 
        ___cell__37600_net131582, n151, n187, n188, n149, n171, n169, n54, 
        n197, n72, n52, n73, ___cell__37600_net131676, n209, 
        ___cell__11920_net39651, n208, ___cell__37600_net131623, 
        ___cell__37600_net131570, ___cell__37600_net131819, n116, n117, n122, 
        ___cell__37600_net131672, n163, n195, n114, n121, n207, n175, n184, 
        n161, n102, n185, n135, n50, ___cell__37600_net131622, 
        ___cell__37600_net131560, ___cell__37600_net131559, n56, n90, n51, 
        ___cell__37600_net131770, ___cell__37600_net131771, n112, n92, n74, 
        ___cell__37600_net131719, n65, n53, n126, n55, n68, n67, net149439, 
        ___cell__37600_net131851, n49, n62, n89, ___cell__37600_net131763, 
        net151798, n57, ___cell__37600_net131869, ___cell__37600_net131867, 
        ___cell__37600_net131866, net149697, ___cell__37600_net131766, 
        net149441, ___cell__37600_net131637, n96, n98, n95, 
        ___cell__37600_net131723, n88, n87, ___cell__37600_net131709, n63, 
        n106, n105, ___cell__37600_net131758, ___cell__37600_net131759, 
        ___cell__37600_net131760, n178, n108, n109, n58, net152263, n100, n110, 
        n59, n64, n104, ___cell__37600_net131873, ___cell__37600_net131767, 
        n91, ___cell__37600_net131861, ___cell__37600_net131620, net150527, 
        ___cell__37600_net131741, n132, n131, net151157, n193, n164, net150528, 
        n107, n101, n80, n79, n177, n60, n61, ___cell__37600_net131634, 
        ___cell__37600_net131562, n145, n125, n166, n162, n159, n99, n85, n66, 
        ___cell__37600_net131733, ___cell__37600_net131556, 
        ___cell__37600_net131596, n182, n128, n129, n75, 
        ___cell__37600_net131776, n70, n69, net149302, n71, n136, n124, 
        ___cell__37600_net131627, n76, n77, ___cell__37600_net131643, n144, 
        ___cell__37600_net131808, ___cell__37600_net131735, 
        ___cell__37600_net131734, ___cell__37600_net131809, 
        ___cell__37600_net131739, ___cell__37600_net131630, 
        ___cell__37600_net131736, ___cell__37600_net131737, 
        ___cell__37600_net131738, ___cell__37600_net131639, 
        ___cell__37600_net131846, n81, ___cell__37600_net131847, n139, n138, 
        n154, n201, n203, ___cell__37600_net131837, n181, 
        ___cell__37600_net131509, ___cell__37600_net131510, n213, n156, 
        ___cell__37600_net131583, n82, ___cell__37600_net131580, n86, n84, n94, 
        n97, n93, ___cell__37600_net131579, ___cell__37600_net131831, 
        ___cell__37600_net131749, ___cell__37600_net131730, n78, n111, 
        ___cell__37600_net131652, ___cell__37600_net131555, n119, n120, 
        ___cell__37600_net131553, ___cell__37600_net131571, n115, n196, 
        ___cell__37600_net131566, net152087, ___cell__37600_net131565, n217, 
        n113, n123, ___cell__37600_net131631, ___cell__37600_net131859, 
        ___cell__37600_net131635, ___cell__37600_net131680, 
        ___cell__37600_net131868, ___cell__37600_net131849, 
        ___cell__37600_net131638, ___cell__37600_net131636, n127, 
        ___cell__37600_net131821, ___cell__37600_net131844, 
        ___cell__37600_net131673, net150977, net151639, net151640, 
        ___cell__11920_net39652, net150978, n133, net152499, 
        ___cell__37600_net131568, n165, n199, n134, net151781, n152, n153, 
        n155, n186, n211, n143, ___cell__37600_net131841, n206, net151782, 
        n198, net151423, n170, n189, net149743, n118, n179, n180, n194, 
        ___cell__37600_net131561, n190, ___cell__37600_net131576, n200, 
        ___cell__37600_net131775, ___cell__37600_net131777, n148, n150, n212, 
        net152089, n214, n216, n192, n191, n205, n176, 
        ___cell__37600_net131811, ___cell__37600_net131858, 
        ___cell__37600_net131823, n130, n142, n147, n172, n167, 
        ___cell__37600_net131610, n146, n168, ___cell__37600_net131641, n173, 
        n202;
    inv_5 U10 ( .x(n183), .a(B[13]) );
    nor2i_1 U100 ( .x(n158), .a(n83), .b(n160) );
    exor2_1 U101 ( .x(SUM[14]), .a(n174), .b(n158) );
    exnor2_1 U102 ( .x(SUM[4]), .a(___cell__37600_net131624), .b(
        ___cell__37600_net131625) );
    inv_5 U103 ( .x(n103), .a(___cell__37600_net131609) );
    nor2i_0 U104 ( .x(___cell__37600_net131611), .a(___cell__37600_net131612), 
        .b(n103) );
    exor2_1 U105 ( .x(SUM[10]), .a(___cell__37600_net131608), .b(
        ___cell__37600_net131611) );
    inv_2 U106 ( .x(___cell__37600_net131586), .a(___cell__37600_net131802) );
    nor2i_1 U107 ( .x(___cell__37600_net131575), .a(n215), .b(net152417) );
    inv_5 U108 ( .x(net152417), .a(___cell__37600_net131806) );
    exnor2_1 U109 ( .x(SUM[2]), .a(n140), .b(___cell__37600_net131584) );
    or3i_3 U11 ( .x(___cell__37600_net131756), .a(n204), .b(n137), .c(n157) );
    nor2i_1 U110 ( .x(n140), .a(n210), .b(net149842) );
    nor2i_0 U111 ( .x(___cell__37600_net131584), .a(___cell__37600_net131585), 
        .b(___cell__37600_net131586) );
    exor2_1 U112 ( .x(___cell__37600_net131640), .a(net148303), .b(B[25]) );
    exnor2_1 U113 ( .x(SUM[21]), .a(n141), .b(___cell__37600_net131645) );
    aoi21_1 U114 ( .x(n141), .a(___cell__37600_net131506), .b(
        ___cell__37600_net131507), .c(___cell__37600_net131508) );
    inv_0 U115 ( .x(___cell__37600_net131508), .a(___cell__37600_net131582) );
    nand2i_2 U116 ( .x(n151), .a(n187), .b(n188) );
    inv_2 U117 ( .x(n149), .a(n151) );
    exnor2_1 U118 ( .x(SUM[18]), .a(n149), .b(n171) );
    exor2_1 U119 ( .x(n169), .a(B[23]), .b(n54) );
    inv_5 U12 ( .x(n157), .a(n197) );
    inv_2 U120 ( .x(n72), .a(n52) );
    inv_4 U121 ( .x(n73), .a(B[30]) );
    inv_2 U122 ( .x(___cell__37600_net131676), .a(B[29]) );
    exnor2_1 U123 ( .x(SUM[1]), .a(n209), .b(___cell__11920_net39651) );
    nor2i_1 U124 ( .x(n209), .a(n210), .b(n208) );
    exnor2_1 U125 ( .x(SUM[5]), .a(___cell__37600_net131623), .b(
        ___cell__37600_net131570) );
    inv_2 U126 ( .x(___cell__37600_net131623), .a(___cell__37600_net131819) );
    aoai211_1 U127 ( .x(___cell__37600_net131819), .a(___cell__37600_net131624
        ), .b(n116), .c(n117), .d(n122) );
    inv_2 U128 ( .x(___cell__37600_net131624), .a(___cell__37600_net131672) );
    inv_2 U129 ( .x(n116), .a(B[4]) );
    inv_10 U13 ( .x(n163), .a(n195) );
    inv_2 U130 ( .x(n114), .a(n121) );
    inv_2 U131 ( .x(n207), .a(n175) );
    inv_2 U132 ( .x(n184), .a(B[12]) );
    exor2_1 U133 ( .x(SUM[13]), .a(n175), .b(n161) );
    inv_2 U135 ( .x(n102), .a(A[11]) );
    inv_2 U136 ( .x(n117), .a(A[4]) );
    inv_0 U137 ( .x(n185), .a(A[12]) );
    inv_10 U138 ( .x(n135), .a(B[17]) );
    oa21_2 U139 ( .x(n50), .a(___cell__37600_net131622), .b(
        ___cell__37600_net131560), .c(___cell__37600_net131559) );
    inv_5 U14 ( .x(n56), .a(n90) );
    nand2_2 U140 ( .x(n51), .a(___cell__37600_net131770), .b(
        ___cell__37600_net131771) );
    inv_5 U141 ( .x(n112), .a(B[7]) );
    inv_2 U142 ( .x(n92), .a(A[21]) );
    exor2_1 U143 ( .x(n52), .a(n74), .b(n73) );
    oai22_3 U144 ( .x(___cell__37600_net131719), .a(A[17]), .b(B[17]), .c(A
        [16]), .d(B[16]) );
    inv_2 U145 ( .x(n65), .a(A[9]) );
    exnor2_1 U146 ( .x(n53), .a(B[29]), .b(net148303) );
    inv_2 U147 ( .x(n54), .a(n126) );
    inv_2 U148 ( .x(n126), .a(A[23]) );
    aoai211_3 U149 ( .x(n55), .a(n68), .b(n67), .c(net149439), .d(
        ___cell__37600_net131851) );
    inv_4 U15 ( .x(n49), .a(n62) );
    inv_2 U151 ( .x(n67), .a(B[28]) );
    or3i_2 U152 ( .x(n89), .a(___cell__37600_net131763), .b(net151798), .c(n57
        ) );
    aoai211_4 U153 ( .x(___cell__37600_net131869), .a(___cell__37600_net131867
        ), .b(___cell__37600_net131866), .c(net149697), .d(
        ___cell__37600_net131766) );
    oaoi211_4 U154 ( .x(net149439), .a(net149441), .b(A[28]), .c(
        ___cell__37600_net131637), .d(n51) );
    aoi21_3 U155 ( .x(net149697), .a(n56), .b(n96), .c(n98) );
    nand2i_1 U156 ( .x(n95), .a(B[21]), .b(___cell__37600_net131582) );
    or3i_5 U158 ( .x(n96), .a(___cell__37600_net131723), .b(n88), .c(n87) );
    nand2i_4 U159 ( .x(___cell__37600_net131609), .a(B[10]), .b(
        ___cell__37600_net131709) );
    nor2_6 U16 ( .x(n62), .a(B[24]), .b(n63) );
    nor2_3 U160 ( .x(n106), .a(n103), .b(n105) );
    nand3_3 U161 ( .x(n88), .a(___cell__37600_net131758), .b(
        ___cell__37600_net131759), .c(___cell__37600_net131760) );
    nand2i_4 U162 ( .x(___cell__37600_net131507), .a(A[20]), .b(n178) );
    nor2_2 U163 ( .x(n108), .a(n105), .b(___cell__37600_net131559) );
    inv_6 U164 ( .x(n105), .a(n109) );
    buf_1 U165 ( .x(n58), .a(net152263) );
    inv_5 U166 ( .x(n100), .a(n110) );
    ao31_3 U167 ( .x(n59), .a(n64), .b(n109), .c(___cell__37600_net131609), 
        .d(n104) );
    exnor2_2 U169 ( .x(SUM[30]), .a(___cell__37600_net131873), .b(n72) );
    inv_6 U17 ( .x(___cell__37600_net131767), .a(n62) );
    nand4_2 U170 ( .x(n91), .a(___cell__37600_net131861), .b(
        ___cell__37600_net131620), .c(___cell__37600_net131760), .d(
        ___cell__37600_net131719) );
    inv_2 U171 ( .x(net150527), .a(___cell__37600_net131741) );
    nand2_1 U172 ( .x(n132), .a(B[1]), .b(A[1]) );
    oai211_1 U173 ( .x(n131), .a(B[1]), .b(A[1]), .c(A[0]), .d(B[0]) );
    inv_0 U174 ( .x(net151157), .a(net149439) );
    exnor2_1 U175 ( .x(n193), .a(A[12]), .b(B[12]) );
    nor2_0 U176 ( .x(n164), .a(A[12]), .b(B[12]) );
    ao21_3 U177 ( .x(net150528), .a(n108), .b(n107), .c(n101) );
    nor2_2 U178 ( .x(n107), .a(n100), .b(n103) );
    ao221_4 U179 ( .x(___cell__37600_net131637), .a(___cell__37600_net131869), 
        .b(n80), .c(B[25]), .d(___cell__37600_net131869), .e(n79) );
    inv_2 U18 ( .x(n177), .a(B[27]) );
    nor2_0 U180 ( .x(n60), .a(n73), .b(n68) );
    inv_2 U181 ( .x(n61), .a(___cell__37600_net131634) );
    exor2_1 U182 ( .x(___cell__37600_net131634), .a(net148303), .b(B[28]) );
    exor2_1 U183 ( .x(SUM[6]), .a(___cell__37600_net131562), .b(n145) );
    inv_2 U184 ( .x(n63), .a(n125) );
    nor2_3 U185 ( .x(n137), .a(B[14]), .b(A[14]) );
    oai211_3 U186 ( .x(n204), .a(n163), .b(n166), .c(n162), .d(n159) );
    nand2_2 U187 ( .x(n162), .a(B[13]), .b(A[13]) );
    inv_0 U188 ( .x(n99), .a(n85) );
    nor2_3 U189 ( .x(n64), .a(n66), .b(n65) );
    nand2_1 U19 ( .x(___cell__37600_net131733), .a(A[4]), .b(B[4]) );
    inv_0 U190 ( .x(___cell__37600_net131556), .a(n64) );
    nor2i_0 U191 ( .x(n161), .a(n162), .b(n163) );
    oai21_1 U192 ( .x(n174), .a(n163), .b(n207), .c(n162) );
    nand2i_2 U193 ( .x(___cell__37600_net131596), .a(n182), .b(B[15]) );
    aoi21_3 U194 ( .x(___cell__37600_net131766), .a(n49), .b(n128), .c(n129)
         );
    inv_2 U195 ( .x(n68), .a(n75) );
    inv_0 U196 ( .x(___cell__37600_net131776), .a(___cell__37600_net131719) );
    exnor2_3 U197 ( .x(SUM[31]), .a(n70), .b(n69) );
    inv_2 U198 ( .x(n69), .a(net149302) );
    oaoi211_2 U199 ( .x(n70), .a(B[30]), .b(n71), .c(___cell__37600_net131873), 
        .d(n60) );
    inv_2 U20 ( .x(n136), .a(n135) );
    inv_1 U200 ( .x(n71), .a(n124) );
    inv_2 U201 ( .x(net149302), .a(___cell__37600_net131627) );
    inv_0 U202 ( .x(n74), .a(net148303) );
    inv_0 U203 ( .x(n75), .a(n124) );
    inv_2 U204 ( .x(___cell__37600_net131851), .a(n76) );
    inv_0 U205 ( .x(n77), .a(net148303) );
    exor2_1 U206 ( .x(SUM[23]), .a(___cell__37600_net131643), .b(n169) );
    nor2i_0 U207 ( .x(n144), .a(___cell__37600_net131559), .b(
        ___cell__37600_net131560) );
    oai211_2 U208 ( .x(___cell__37600_net131808), .a(___cell__37600_net131735), 
        .b(___cell__37600_net131734), .c(___cell__37600_net131809), .d(
        ___cell__37600_net131739) );
    oai211_2 U209 ( .x(___cell__37600_net131735), .a(___cell__37600_net131630), 
        .b(___cell__37600_net131736), .c(___cell__37600_net131737), .d(
        ___cell__37600_net131738) );
    nand2_2 U21 ( .x(___cell__37600_net131758), .a(A[17]), .b(n136) );
    inv_2 U210 ( .x(n80), .a(n124) );
    inv_0 U211 ( .x(___cell__37600_net131639), .a(___cell__37600_net131869) );
    nand2_1 U212 ( .x(___cell__37600_net131846), .a(B[25]), .b(net148303) );
    inv_0 U213 ( .x(n124), .a(A[31]) );
    inv_0 U214 ( .x(n81), .a(___cell__37600_net131847) );
    nand2_5 U215 ( .x(___cell__37600_net131760), .a(A[18]), .b(n139) );
    inv_3 U216 ( .x(n138), .a(B[18]) );
    nand2i_4 U217 ( .x(n188), .a(___cell__37600_net131719), .b(n154) );
    inv_0 U218 ( .x(n201), .a(n203) );
    nand2_0 U219 ( .x(___cell__37600_net131837), .a(A[18]), .b(n139) );
    nand2i_2 U22 ( .x(___cell__37600_net131861), .a(n181), .b(n203) );
    aoi21_1 U220 ( .x(___cell__37600_net131509), .a(___cell__37600_net131510), 
        .b(___cell__37600_net131506), .c(n213) );
    nor2i_1 U221 ( .x(n156), .a(___cell__37600_net131596), .b(n157) );
    nor2_0 U222 ( .x(___cell__37600_net131510), .a(___cell__37600_net131583), 
        .b(net151798) );
    inv_0 U223 ( .x(n82), .a(n159) );
    inv_2 U224 ( .x(n83), .a(n82) );
    inv_0 U225 ( .x(___cell__37600_net131643), .a(net149697) );
    inv_0 U226 ( .x(___cell__37600_net131580), .a(___cell__37600_net131763) );
    nand2_5 U227 ( .x(n87), .a(___cell__37600_net131756), .b(n86) );
    and2_3 U228 ( .x(n86), .a(___cell__37600_net131620), .b(
        ___cell__37600_net131596) );
    nor2i_3 U229 ( .x(n84), .a(___cell__37600_net131620), .b(net152263) );
    oa22_3 U23 ( .x(net152263), .a(B[18]), .b(A[18]), .c(B[19]), .d(A[19]) );
    nand2_1 U230 ( .x(n94), .a(___cell__37600_net131582), .b(n92) );
    inv_2 U231 ( .x(n97), .a(n93) );
    exor2_1 U232 ( .x(___cell__37600_net131645), .a(A[21]), .b(n97) );
    inv_0 U233 ( .x(n85), .a(A[22]) );
    nand2_1 U234 ( .x(___cell__37600_net131579), .a(A[22]), .b(B[22]) );
    ao211_5 U235 ( .x(___cell__37600_net131831), .a(net150527), .b(
        ___cell__37600_net131808), .c(net150528), .d(n59) );
    nand2i_4 U236 ( .x(___cell__37600_net131723), .a(___cell__37600_net131749), 
        .b(___cell__37600_net131831) );
    inv_0 U237 ( .x(___cell__37600_net131730), .a(___cell__37600_net131831) );
    and3i_2 U238 ( .x(n104), .a(n105), .b(n78), .c(A[10]) );
    inv_0 U239 ( .x(n111), .a(n102) );
    nand2_2 U24 ( .x(___cell__37600_net131582), .a(A[20]), .b(B[20]) );
    exor2_1 U240 ( .x(___cell__37600_net131652), .a(B[11]), .b(n111) );
    or3i_2 U241 ( .x(___cell__37600_net131741), .a(n106), .b(n100), .c(
        ___cell__37600_net131560) );
    oai21_1 U242 ( .x(___cell__37600_net131608), .a(n50), .b(n100), .c(
        ___cell__37600_net131556) );
    nor2i_0 U243 ( .x(___cell__37600_net131555), .a(___cell__37600_net131556), 
        .b(n100) );
    inv_0 U244 ( .x(___cell__37600_net131622), .a(___cell__37600_net131808) );
    aoi21_3 U245 ( .x(___cell__37600_net131739), .a(n119), .b(n120), .c(
        ___cell__37600_net131553) );
    nor2i_1 U246 ( .x(___cell__37600_net131553), .a(A[7]), .b(n112) );
    nand2i_6 U247 ( .x(___cell__37600_net131738), .a(A[7]), .b(n112) );
    aoi21_2 U248 ( .x(n120), .a(___cell__37600_net131571), .b(
        ___cell__37600_net131733), .c(n115) );
    nor2_1 U249 ( .x(n115), .a(B[5]), .b(A[5]) );
    nand2i_2 U25 ( .x(n196), .a(A[12]), .b(n184) );
    nor2_8 U250 ( .x(n119), .a(___cell__37600_net131566), .b(net152087) );
    aoi21_1 U251 ( .x(___cell__37600_net131565), .a(n217), .b(B[7]), .c(
        ___cell__37600_net131566) );
    nand2i_4 U252 ( .x(___cell__37600_net131734), .a(n114), .b(n113) );
    oai21_1 U253 ( .x(___cell__37600_net131562), .a(n114), .b(
        ___cell__37600_net131623), .c(___cell__37600_net131571) );
    nor2i_0 U254 ( .x(___cell__37600_net131570), .a(___cell__37600_net131571), 
        .b(n114) );
    aoi21_4 U255 ( .x(___cell__37600_net131737), .a(n116), .b(n117), .c(
        net152417) );
    aoai211_4 U256 ( .x(___cell__37600_net131873), .a(n123), .b(
        ___cell__37600_net131676), .c(___cell__37600_net131631), .d(
        ___cell__37600_net131859) );
    inv_2 U257 ( .x(n123), .a(A[31]) );
    aoai211_1 U259 ( .x(___cell__37600_net131635), .a(___cell__37600_net131680
        ), .b(n124), .c(___cell__37600_net131847), .d(___cell__37600_net131770
        ) );
    nand2_1 U26 ( .x(___cell__37600_net131770), .a(B[26]), .b(net148303) );
    inv_5 U260 ( .x(net149441), .a(___cell__37600_net131868) );
    nand2i_4 U261 ( .x(___cell__37600_net131868), .a(___cell__37600_net131680), 
        .b(___cell__37600_net131849) );
    inv_0 U262 ( .x(___cell__37600_net131847), .a(___cell__37600_net131637) );
    exor2_1 U263 ( .x(SUM[26]), .a(n81), .b(___cell__37600_net131638) );
    nand2_3 U264 ( .x(___cell__37600_net131636), .a(___cell__37600_net131771), 
        .b(___cell__37600_net131849) );
    exor2_2 U265 ( .x(___cell__37600_net131627), .a(net148303), .b(B[31]) );
    nor2i_6 U266 ( .x(n128), .a(A[23]), .b(n127) );
    inv_10 U267 ( .x(n127), .a(B[23]) );
    nand2i_4 U268 ( .x(___cell__37600_net131866), .a(n127), .b(
        ___cell__37600_net131767) );
    nand2i_4 U269 ( .x(___cell__37600_net131867), .a(n126), .b(
        ___cell__37600_net131767) );
    nand2_2 U27 ( .x(___cell__37600_net131771), .a(B[27]), .b(net148303) );
    inv_0 U270 ( .x(___cell__37600_net131821), .a(___cell__37600_net131767) );
    inv_0 U271 ( .x(n125), .a(A[24]) );
    nand2_2 U272 ( .x(___cell__37600_net131844), .a(A[24]), .b(B[24]) );
    inv_0 U273 ( .x(___cell__37600_net131673), .a(___cell__37600_net131630) );
    nand2_2 U274 ( .x(___cell__37600_net131585), .a(A[2]), .b(B[2]) );
    inv_0 U275 ( .x(net150977), .a(A[1]) );
    inv_0 U276 ( .x(net151639), .a(A[0]) );
    nand2_0 U277 ( .x(___cell__11920_net39651), .a(net151640), .b(B[0]) );
    nor2_0 U278 ( .x(___cell__11920_net39652), .a(B[0]), .b(net151640) );
    oa211_1 U279 ( .x(net149842), .a(B[1]), .b(net150978), .c(net151640), .d(B
        [0]) );
    nor2i_1 U28 ( .x(n76), .a(B[28]), .b(n77) );
    nand2i_4 U280 ( .x(___cell__37600_net131806), .a(B[3]), .b(n133) );
    exor2_1 U281 ( .x(___cell__37600_net131625), .a(A[4]), .b(B[4]) );
    oai21_1 U282 ( .x(___cell__37600_net131672), .a(___cell__37600_net131673), 
        .b(net152417), .c(n215) );
    exnor2_1 U283 ( .x(SUM[25]), .a(___cell__37600_net131639), .b(
        ___cell__37600_net131640) );
    exnor2_1 U284 ( .x(SUM[8]), .a(___cell__37600_net131622), .b(n144) );
    and2_2 U285 ( .x(net152499), .a(A[6]), .b(B[6]) );
    inv_0 U286 ( .x(___cell__37600_net131568), .a(net152499) );
    mux2i_1 U287 ( .x(SUM[12]), .d0(n165), .sl(___cell__37600_net131730), .d1(
        n193) );
    aoai211_1 U288 ( .x(n175), .a(n185), .b(n184), .c(___cell__37600_net131730
        ), .d(n166) );
    inv_6 U289 ( .x(___cell__37600_net131709), .a(A[10]) );
    inv_2 U29 ( .x(net148303), .a(n123) );
    nand3_0 U290 ( .x(n199), .a(___cell__37600_net131758), .b(
        ___cell__37600_net131759), .c(___cell__37600_net131760) );
    buf_3 U291 ( .x(n134), .a(B[8]) );
    exor2_1 U292 ( .x(SUM[3]), .a(___cell__37600_net131630), .b(
        ___cell__37600_net131575) );
    inv_2 U293 ( .x(n182), .a(A[15]) );
    inv_0 U294 ( .x(net151781), .a(___cell__37600_net131723) );
    aoi21_1 U296 ( .x(n152), .a(n153), .b(n154), .c(n155) );
    oai22_1 U297 ( .x(n187), .a(n135), .b(n186), .c(n201), .d(n211) );
    nand2i_0 U298 ( .x(n143), .a(n186), .b(n154) );
    inv_0 U299 ( .x(___cell__37600_net131841), .a(___cell__37600_net131620) );
    nand2i_2 U30 ( .x(___cell__37600_net131809), .a(___cell__37600_net131566), 
        .b(net152499) );
    nand2_1 U300 ( .x(___cell__37600_net131759), .a(A[16]), .b(B[16]) );
    nand2_0 U301 ( .x(n186), .a(A[16]), .b(B[16]) );
    inv_2 U303 ( .x(net151640), .a(net151639) );
    or3i_1 U305 ( .x(n206), .a(net151782), .b(n198), .c(n199) );
    inv_0 U306 ( .x(net151423), .a(___cell__37600_net131643) );
    exor2_1 U307 ( .x(n170), .a(B[19]), .b(A[19]) );
    inv_2 U308 ( .x(net150978), .a(net150977) );
    exnor2_1 U309 ( .x(n189), .a(A[9]), .b(net149743) );
    nand2i_2 U31 ( .x(n121), .a(B[5]), .b(n118) );
    inv_4 U310 ( .x(n139), .a(n138) );
    nand2_0 U311 ( .x(n198), .a(___cell__37600_net131756), .b(
        ___cell__37600_net131596) );
    nand2_2 U312 ( .x(___cell__37600_net131571), .a(A[5]), .b(B[5]) );
    inv_0 U313 ( .x(n179), .a(B[16]) );
    nand2i_0 U314 ( .x(n153), .a(B[16]), .b(n180) );
    ao21_3 U315 ( .x(n203), .a(A[16]), .b(B[16]), .c(B[17]) );
    inv_0 U316 ( .x(n160), .a(n194) );
    nand2_0 U317 ( .x(___cell__37600_net131612), .a(A[10]), .b(n78) );
    mux2i_1 U318 ( .x(SUM[7]), .d0(___cell__37600_net131565), .sl(
        ___cell__37600_net131561), .d1(n190) );
    exnor2_1 U319 ( .x(n190), .a(n217), .b(B[7]) );
    nand2_1 U32 ( .x(___cell__37600_net131576), .a(A[3]), .b(B[3]) );
    oai31_1 U320 ( .x(n200), .a(___cell__37600_net131775), .b(
        ___cell__37600_net131776), .c(___cell__37600_net131777), .d(n58) );
    nand2_0 U321 ( .x(n210), .a(net150978), .b(B[1]) );
    nor2_0 U322 ( .x(n208), .a(B[1]), .b(net150978) );
    nor2i_3 U323 ( .x(n148), .a(n139), .b(n149) );
    exor2_1 U324 ( .x(n171), .a(A[18]), .b(n139) );
    oaoi211_1 U325 ( .x(n150), .a(n139), .b(n151), .c(A[18]), .d(n148) );
    nand4_1 U326 ( .x(___cell__37600_net131749), .a(n197), .b(n195), .c(n196), 
        .d(n194) );
    nand2i_6 U327 ( .x(___cell__37600_net131849), .a(net148303), .b(n177) );
    nand2i_2 U328 ( .x(n154), .a(n198), .b(net151782) );
    inv_2 U329 ( .x(net151782), .a(net151781) );
    inv_7 U33 ( .x(___cell__37600_net131566), .a(___cell__37600_net131738) );
    inv_4 U330 ( .x(___cell__37600_net131631), .a(n55) );
    exnor2_1 U331 ( .x(SUM[29]), .a(n55), .b(n53) );
    inv_0 U332 ( .x(n211), .a(A[17]) );
    inv_2 U333 ( .x(n181), .a(A[17]) );
    exnor2_3 U334 ( .x(SUM[19]), .a(n150), .b(n170) );
    inv_0 U335 ( .x(n212), .a(net152089) );
    inv_2 U336 ( .x(n213), .a(n212) );
    oa211_4 U337 ( .x(net152089), .a(A[21]), .b(n97), .c(n94), .d(n95) );
    aoai211_2 U338 ( .x(___cell__37600_net131630), .a(n131), .b(n132), .c(
        ___cell__37600_net131586), .d(___cell__37600_net131585) );
    inv_0 U339 ( .x(n214), .a(___cell__37600_net131576) );
    buf_2 U34 ( .x(net149743), .a(B[9]) );
    inv_2 U340 ( .x(n215), .a(n214) );
    nand2_3 U341 ( .x(___cell__37600_net131620), .a(A[19]), .b(B[19]) );
    inv_0 U342 ( .x(n216), .a(A[7]) );
    inv_2 U343 ( .x(n217), .a(n216) );
    buf_2 U35 ( .x(n78), .a(B[10]) );
    nor2i_0 U36 ( .x(n101), .a(B[11]), .b(n102) );
    nor2i_0 U37 ( .x(n192), .a(n179), .b(n154) );
    exnor2_1 U38 ( .x(n191), .a(n154), .b(n179) );
    inv_2 U40 ( .x(___cell__37600_net131777), .a(___cell__37600_net131837) );
    inv_0 U41 ( .x(___cell__37600_net131775), .a(___cell__37600_net131861) );
    nand2i_2 U42 ( .x(n205), .a(n200), .b(n206) );
    inv_2 U43 ( .x(n176), .a(A[8]) );
    nand2i_2 U44 ( .x(___cell__37600_net131811), .a(B[8]), .b(n176) );
    nand2_2 U45 ( .x(___cell__37600_net131559), .a(A[8]), .b(n134) );
    inv_2 U46 ( .x(n180), .a(A[16]) );
    nand2_2 U47 ( .x(___cell__37600_net131858), .a(B[23]), .b(n54) );
    nand2i_4 U48 ( .x(n197), .a(B[15]), .b(n182) );
    inv_4 U49 ( .x(n113), .a(net152087) );
    oa21_3 U5 ( .x(n98), .a(net152089), .b(___cell__37600_net131823), .c(
        ___cell__37600_net131763) );
    nor2_6 U50 ( .x(net152087), .a(B[6]), .b(A[6]) );
    nand2_2 U51 ( .x(n159), .a(A[14]), .b(B[14]) );
    inv_2 U52 ( .x(n66), .a(net149743) );
    nand2i_2 U53 ( .x(n110), .a(B[9]), .b(n65) );
    inv_2 U54 ( .x(n133), .a(A[3]) );
    inv_2 U55 ( .x(___cell__37600_net131736), .a(___cell__37600_net131576) );
    inv_4 U56 ( .x(n130), .a(A[2]) );
    nand2i_2 U57 ( .x(___cell__37600_net131802), .a(B[2]), .b(n130) );
    inv_2 U58 ( .x(n129), .a(___cell__37600_net131844) );
    inv_5 U59 ( .x(n178), .a(B[20]) );
    or2_6 U6 ( .x(___cell__37600_net131763), .a(B[22]), .b(n99) );
    or3i_2 U60 ( .x(n90), .a(n91), .b(n84), .c(n89) );
    inv_2 U61 ( .x(n57), .a(___cell__37600_net131507) );
    inv_2 U62 ( .x(___cell__37600_net131823), .a(___cell__37600_net131579) );
    inv_3 U63 ( .x(n93), .a(B[21]) );
    nand2_2 U64 ( .x(___cell__37600_net131859), .a(B[29]), .b(net148303) );
    inv_2 U65 ( .x(n118), .a(A[5]) );
    nand2i_2 U66 ( .x(n122), .a(n116), .b(___cell__37600_net131672) );
    nand2_2 U67 ( .x(n166), .a(A[12]), .b(B[12]) );
    inv_5 U68 ( .x(___cell__37600_net131680), .a(B[26]) );
    exnor2_1 U69 ( .x(SUM[27]), .a(___cell__37600_net131635), .b(
        ___cell__37600_net131636) );
    nand2i_4 U7 ( .x(n109), .a(B[11]), .b(n102) );
    exnor2_1 U70 ( .x(SUM[28]), .a(net151157), .b(n61) );
    aoi21_1 U71 ( .x(___cell__37600_net131561), .a(___cell__37600_net131562), 
        .b(n113), .c(net152499) );
    inv_2 U72 ( .x(n79), .a(___cell__37600_net131846) );
    exor2_1 U73 ( .x(___cell__37600_net131638), .a(net148303), .b(B[26]) );
    nor2i_1 U74 ( .x(n165), .a(n166), .b(n164) );
    mux2i_1 U75 ( .x(n142), .d0(n191), .sl(A[16]), .d1(n192) );
    nand2_2 U76 ( .x(SUM[16]), .a(n142), .b(n143) );
    exor2_1 U77 ( .x(SUM[20]), .a(___cell__37600_net131506), .b(n147) );
    nand2i_2 U78 ( .x(___cell__37600_net131506), .a(___cell__37600_net131841), 
        .b(n205) );
    nor2i_1 U79 ( .x(n147), .a(___cell__37600_net131582), .b(
        ___cell__37600_net131583) );
    and2_3 U8 ( .x(net151798), .a(n92), .b(n93) );
    inv_2 U80 ( .x(___cell__37600_net131583), .a(___cell__37600_net131507) );
    inv_2 U81 ( .x(___cell__37600_net131560), .a(___cell__37600_net131811) );
    mux2i_1 U82 ( .x(SUM[9]), .d0(___cell__37600_net131555), .sl(n50), .d1(
        n189) );
    exor2_1 U83 ( .x(n172), .a(A[17]), .b(n136) );
    inv_2 U84 ( .x(n155), .a(n186) );
    exnor2_1 U85 ( .x(SUM[17]), .a(n152), .b(n172) );
    nor2i_1 U86 ( .x(SUM[0]), .a(___cell__11920_net39651), .b(
        ___cell__11920_net39652) );
    exnor2_1 U87 ( .x(SUM[11]), .a(n167), .b(___cell__37600_net131652) );
    aoi21_1 U88 ( .x(n167), .a(___cell__37600_net131608), .b(
        ___cell__37600_net131609), .c(___cell__37600_net131610) );
    inv_2 U89 ( .x(___cell__37600_net131610), .a(___cell__37600_net131612) );
    nand2i_3 U9 ( .x(n195), .a(A[13]), .b(n183) );
    exnor2_1 U90 ( .x(SUM[22]), .a(___cell__37600_net131509), .b(n146) );
    nor2i_1 U91 ( .x(n146), .a(___cell__37600_net131579), .b(
        ___cell__37600_net131580) );
    nand2i_0 U92 ( .x(n168), .a(___cell__37600_net131821), .b(
        ___cell__37600_net131844) );
    aoai211_1 U93 ( .x(___cell__37600_net131641), .a(n126), .b(n127), .c(
        net151423), .d(___cell__37600_net131858) );
    exnor2_1 U94 ( .x(SUM[24]), .a(___cell__37600_net131641), .b(n168) );
    exor2_1 U95 ( .x(SUM[15]), .a(n173), .b(n156) );
    oai21_1 U96 ( .x(n173), .a(n160), .b(n202), .c(n83) );
    inv_2 U97 ( .x(n194), .a(n137) );
    nor2i_0 U98 ( .x(n145), .a(___cell__37600_net131568), .b(net152087) );
    inv_2 U99 ( .x(n202), .a(n174) );
endmodule


module ID_DW01_add_32_1_test_1 ( A, B, CI, SUM, CO );
input  [31:0] A;
input  [31:0] B;
output [31:0] SUM;
input  CI;
output CO;
    wire n277, n217, n218, n106, n173, n170, n177, n178, n176, n191, n314, n79, 
        n316, n219, n105, n321, n62, n110, n302, n146, n308, n216, n149, n325, 
        n301, n282, n283, n152, n322, n127, n199, n53, n188, n189, n190, n66, 
        n55, n186, n187, n230, n232, n212, n145, n157, n158, n305, n150, n85, 
        n109, n226, n147, n265, n139, n135, n136, n137, n337, n210, n87, n209, 
        n328, n336, n239, n207, n88, n240, n267, n206, n117, n185, n98, n320, 
        n319, n99, n100, n245, n231, n211, n132, n89, n90, n148, n96, n97, 
        n263, n261, n114, n138, n115, n116, n140, n163, n327, n101, n111, n141, 
        n104, n213, n151, n229, n51, n153, n74, n123, n162, n313, n130, n124, 
        n125, n131, n311, n129, n80, n323, n250, n202, n254, n94, n275, n169, 
        n93, n345, n278, n91, n92, n347, n338, n269, n204, n307, n346, n262, 
        n70, n59, n154, n57, n156, n108, n225, n258, n289, n268, n107, n58, 
        n171, n75, n256, n259, n54, n172, n174, n304, n343, n317, n342, n279, 
        n95, n69, n183, n184, n306, n67, n68, n271, n56, n249, n248, n247, 
        n155, n175, n143, n237, n288, n287, n72, n60, n61, n159, n236, n280, 
        n63, n257, n266, n119, n341, n81, n233, n330, n82, n222, n293, n76, 
        n77, n64, n65, n179, n180, n181, n310, n198, n312, n142, n160, n329, 
        n201, n161, n331, n332, n71, n333, n295, n83, n120, n290, n73, n195, 
        n220, n228, n118, n324, n253, n192, n318, n334, n50, n164, n144, n78, 
        n128, n235, n86, n224, n281, n309, n167, n298, n299, n214, n84, n126, 
        n296, n165, n166, n168, n196, n197, n200, n203, n205, n303, n244, n238, 
        n133, n134, n270, n272, n274, n264, n291, n292, n251, n294, n297, n255, 
        n208, n315, n102, n326, n52, n335, n300, n339, n344, n284, n340, n103, 
        n276, n194, n193, n121, n122, n221, n285, n223, n252, n273, n182, n49, 
        n215, n234, n241, n242, n243, n260, n112, n227, n113, n246, n286;
    ao21_3 U10 ( .x(n277), .a(n217), .b(n218), .c(n106) );
    nand2i_2 U100 ( .x(n173), .a(B[30]), .b(n170) );
    nor2i_1 U101 ( .x(n177), .a(n178), .b(n176) );
    ao21_1 U102 ( .x(n191), .a(n314), .b(n79), .c(n316) );
    inv_2 U103 ( .x(n219), .a(A[4]) );
    inv_2 U104 ( .x(n316), .a(n105) );
    nand2_2 U105 ( .x(n105), .a(A[4]), .b(B[4]) );
    inv_2 U106 ( .x(n321), .a(n191) );
    inv_2 U107 ( .x(n106), .a(n314) );
    inv_5 U108 ( .x(n62), .a(B[13]) );
    nand2_0 U109 ( .x(n110), .a(n302), .b(n146) );
    nand2i_3 U11 ( .x(n308), .a(B[6]), .b(n216) );
    nand2i_2 U110 ( .x(n302), .a(n149), .b(n325) );
    nand2i_0 U111 ( .x(n301), .a(n282), .b(n283) );
    inv_2 U112 ( .x(n282), .a(n152) );
    inv_2 U113 ( .x(n322), .a(n127) );
    exnor2_3 U114 ( .x(SUM[27]), .a(n199), .b(n53) );
    exor2_1 U115 ( .x(SUM[7]), .a(n188), .b(n189) );
    ao21_1 U116 ( .x(n188), .a(n190), .b(n66), .c(n55) );
    exnor2_1 U117 ( .x(SUM[8]), .a(n186), .b(n187) );
    nand2i_2 U118 ( .x(n187), .a(n230), .b(n232) );
    exor2_1 U119 ( .x(SUM[12]), .a(n212), .b(n145) );
    nor2i_3 U12 ( .x(n157), .a(B[7]), .b(n158) );
    oai21_1 U120 ( .x(n212), .a(n305), .b(n150), .c(n85) );
    inv_2 U121 ( .x(n305), .a(n109) );
    inv_0 U122 ( .x(n150), .a(n226) );
    nor2i_0 U123 ( .x(n145), .a(n146), .b(n147) );
    inv_0 U124 ( .x(n147), .a(n325) );
    inv_2 U125 ( .x(n265), .a(n139) );
    nor2i_1 U126 ( .x(n135), .a(n136), .b(n137) );
    inv_2 U127 ( .x(n137), .a(n337) );
    exor2_1 U128 ( .x(n210), .a(B[19]), .b(n87) );
    nand2_2 U129 ( .x(n209), .a(n328), .b(n336) );
    inv_0 U13 ( .x(n239), .a(B[18]) );
    exor2_1 U130 ( .x(SUM[19]), .a(n209), .b(n210) );
    exor2_1 U131 ( .x(n207), .a(B[20]), .b(n88) );
    inv_2 U132 ( .x(n240), .a(B[19]) );
    inv_2 U133 ( .x(n328), .a(n267) );
    oai22_1 U134 ( .x(n206), .a(n328), .b(n240), .c(n117), .d(n170) );
    exor2_1 U136 ( .x(SUM[9]), .a(n185), .b(n98) );
    oai21_1 U137 ( .x(n185), .a(n320), .b(n230), .c(n232) );
    inv_2 U138 ( .x(n230), .a(n319) );
    nor2i_0 U139 ( .x(n98), .a(n99), .b(n100) );
    nand2_2 U14 ( .x(n245), .a(B[18]), .b(n88) );
    inv_5 U140 ( .x(n100), .a(n231) );
    exor2_1 U141 ( .x(SUM[17]), .a(n211), .b(n132) );
    nor2i_1 U142 ( .x(SUM[0]), .a(n89), .b(n90) );
    exor2_1 U143 ( .x(SUM[11]), .a(n109), .b(n148) );
    nand2_2 U144 ( .x(SUM[22]), .a(n96), .b(n97) );
    nand2i_2 U146 ( .x(n97), .a(n263), .b(n261) );
    exnor2_1 U147 ( .x(SUM[15]), .a(n114), .b(n138) );
    aoi21_1 U148 ( .x(n114), .a(n115), .b(n109), .c(n116) );
    nor2i_1 U149 ( .x(n138), .a(n139), .b(n140) );
    inv_2 U15 ( .x(n163), .a(B[13]) );
    inv_5 U150 ( .x(n140), .a(n327) );
    exor2_1 U151 ( .x(SUM[6]), .a(n190), .b(n101) );
    exnor2_1 U152 ( .x(SUM[14]), .a(n111), .b(n141) );
    exor2_1 U153 ( .x(SUM[4]), .a(n79), .b(n104) );
    nor2i_0 U154 ( .x(n104), .a(n105), .b(n106) );
    exor2_1 U155 ( .x(SUM[10]), .a(n213), .b(n151) );
    oai21_1 U156 ( .x(n213), .a(n320), .b(n229), .c(n51) );
    inv_2 U157 ( .x(n320), .a(n186) );
    nor2i_0 U158 ( .x(n151), .a(n152), .b(n153) );
    exor2_1 U159 ( .x(SUM[3]), .a(n74), .b(n123) );
    nor2i_1 U16 ( .x(n162), .a(A[13]), .b(n163) );
    inv_2 U160 ( .x(n313), .a(n130) );
    nor2i_1 U161 ( .x(n123), .a(n124), .b(n125) );
    inv_2 U162 ( .x(n131), .a(n311) );
    nor2i_1 U163 ( .x(n129), .a(n130), .b(n131) );
    exor2_1 U164 ( .x(SUM[2]), .a(n80), .b(n129) );
    inv_2 U165 ( .x(n323), .a(n250) );
    nand2i_2 U166 ( .x(n202), .a(n323), .b(n254) );
    mux2i_1 U167 ( .x(n94), .d0(n275), .sl(B[21]), .d1(n169) );
    inv_0 U169 ( .x(n93), .a(n345) );
    nor2_1 U17 ( .x(n278), .a(B[22]), .b(B[21]) );
    nand2_2 U170 ( .x(SUM[18]), .a(n91), .b(n92) );
    nand3i_1 U171 ( .x(n92), .a(n347), .b(n87), .c(n338) );
    inv_2 U172 ( .x(n338), .a(n269) );
    nand3i_1 U173 ( .x(n204), .a(n307), .b(n346), .c(n262) );
    inv_2 U174 ( .x(n307), .a(n263) );
    inv_3 U176 ( .x(n70), .a(n59) );
    nor2i_1 U177 ( .x(n154), .a(n57), .b(n156) );
    exnor2_1 U178 ( .x(SUM[1]), .a(n154), .b(n89) );
    inv_2 U179 ( .x(n108), .a(n225) );
    nand2i_3 U18 ( .x(n258), .a(n289), .b(n268) );
    aoi21_1 U180 ( .x(n107), .a(n108), .b(n109), .c(n110) );
    inv_0 U181 ( .x(n58), .a(A[14]) );
    oa21_1 U183 ( .x(n51), .a(n100), .b(n232), .c(n99) );
    exnor2_1 U184 ( .x(n53), .a(B[27]), .b(n87) );
    aoai211_4 U185 ( .x(n171), .a(n75), .b(n256), .c(n258), .d(n259) );
    exnor2_1 U187 ( .x(n54), .a(B[28]), .b(n87) );
    aoi22_2 U188 ( .x(n172), .a(B[30]), .b(n88), .c(n174), .d(n173) );
    nand2i_2 U189 ( .x(n109), .a(n301), .b(n304) );
    nand2_2 U19 ( .x(n289), .a(B[20]), .b(B[19]) );
    aoai211_3 U190 ( .x(n304), .a(n343), .b(n317), .c(n342), .d(n279) );
    oai21_1 U191 ( .x(SUM[21]), .a(n93), .b(n94), .c(n95) );
    inv_5 U192 ( .x(n69), .a(A[3]) );
    nor2i_2 U193 ( .x(n183), .a(B[21]), .b(n184) );
    nand3i_5 U194 ( .x(n306), .a(B[21]), .b(n184), .c(n345) );
    nand2_1 U195 ( .x(n152), .a(A[10]), .b(B[10]) );
    nor2i_3 U196 ( .x(n67), .a(n68), .b(A[1]) );
    oai21_3 U197 ( .x(n271), .a(n100), .b(n232), .c(n99) );
    inv_0 U198 ( .x(n56), .a(n218) );
    nand2i_0 U199 ( .x(n337), .a(B[16]), .b(n170) );
    or3i_2 U20 ( .x(n249), .a(n250), .b(n248), .c(n247) );
    nand2_0 U200 ( .x(n136), .a(B[16]), .b(n87) );
    buf_1 U201 ( .x(n57), .a(n155) );
    nor2_1 U202 ( .x(n175), .a(B[5]), .b(A[5]) );
    and2_5 U203 ( .x(n143), .a(n58), .b(n237) );
    and2_5 U204 ( .x(n256), .a(n288), .b(n287) );
    nand2i_2 U205 ( .x(n66), .a(B[6]), .b(n216) );
    inv_2 U206 ( .x(n72), .a(B[0]) );
    nor2i_5 U207 ( .x(n60), .a(n62), .b(n61) );
    inv_0 U208 ( .x(n159), .a(n60) );
    inv_2 U209 ( .x(n61), .a(n236) );
    nor2i_2 U21 ( .x(n279), .a(n280), .b(n229) );
    inv_0 U210 ( .x(n236), .a(A[13]) );
    or3i_2 U211 ( .x(n63), .a(n257), .b(n265), .c(n266) );
    or3i_3 U212 ( .x(n119), .a(n257), .b(n265), .c(n266) );
    inv_7 U213 ( .x(n342), .a(n341) );
    ao211_5 U214 ( .x(n75), .a(n304), .b(n81), .c(n233), .d(n140) );
    or3i_4 U215 ( .x(n330), .a(n82), .b(n222), .c(n293) );
    nor2_2 U216 ( .x(n76), .a(n69), .b(n77) );
    inv_0 U217 ( .x(n64), .a(B[13]) );
    inv_2 U218 ( .x(n65), .a(n64) );
    nand2i_0 U219 ( .x(n186), .a(n179), .b(n341) );
    nand2_2 U22 ( .x(n343), .a(n180), .b(n181) );
    nand2_2 U220 ( .x(n310), .a(n77), .b(n69) );
    exnor2_3 U221 ( .x(SUM[28]), .a(n198), .b(n54) );
    inv_3 U222 ( .x(n312), .a(n67) );
    inv_0 U223 ( .x(n89), .a(n70) );
    nor2i_0 U224 ( .x(n141), .a(n142), .b(n143) );
    oai31_1 U225 ( .x(n116), .a(n160), .b(n143), .c(n60), .d(n142) );
    nand2_5 U226 ( .x(n329), .a(n250), .b(n201) );
    nand4i_3 U227 ( .x(n174), .a(n161), .b(n330), .c(n331), .d(n332) );
    buf_4 U228 ( .x(n71), .a(B[12]) );
    nand2i_2 U229 ( .x(n333), .a(n295), .b(n82) );
    nand2_2 U23 ( .x(n283), .a(n271), .b(n280) );
    exnor2_1 U230 ( .x(SUM[25]), .a(n82), .b(n202) );
    inv_3 U231 ( .x(n83), .a(n184) );
    oai211_4 U232 ( .x(n201), .a(n184), .b(n120), .c(n290), .d(n345) );
    inv_2 U233 ( .x(n77), .a(B[3]) );
    exor2_1 U234 ( .x(n189), .a(B[7]), .b(A[7]) );
    inv_2 U235 ( .x(n158), .a(A[7]) );
    inv_0 U236 ( .x(n73), .a(n195) );
    inv_2 U237 ( .x(n74), .a(n73) );
    nand2_5 U238 ( .x(n232), .a(A[8]), .b(B[8]) );
    inv_4 U239 ( .x(n220), .a(A[8]) );
    nand2i_2 U24 ( .x(n280), .a(B[10]), .b(n228) );
    nor2i_1 U240 ( .x(n117), .a(n118), .b(n63) );
    exor2_1 U241 ( .x(SUM[16]), .a(n63), .b(n135) );
    nand2i_0 U242 ( .x(n336), .a(n170), .b(n63) );
    ao21_3 U243 ( .x(n211), .a(n337), .b(n63), .c(n324) );
    inv_0 U244 ( .x(n156), .a(n312) );
    ao211_3 U245 ( .x(n257), .a(n304), .b(n81), .c(n140), .d(n233) );
    nand2_2 U246 ( .x(n253), .a(B[27]), .b(n88) );
    inv_0 U247 ( .x(n124), .a(n76) );
    ao21_4 U248 ( .x(n192), .a(n310), .b(n195), .c(n76) );
    inv_0 U249 ( .x(n125), .a(n310) );
    inv_0 U25 ( .x(n228), .a(A[10]) );
    nand2_1 U250 ( .x(n318), .a(B[5]), .b(A[5]) );
    nand2_0 U251 ( .x(n178), .a(n56), .b(A[5]) );
    nor2_0 U252 ( .x(n176), .a(n56), .b(A[5]) );
    nand2i_2 U253 ( .x(n334), .a(n50), .b(n170) );
    inv_2 U254 ( .x(n248), .a(B[26]) );
    nor2_1 U255 ( .x(n164), .a(B[13]), .b(A[13]) );
    aoi21_1 U256 ( .x(n144), .a(A[13]), .b(n65), .c(n60) );
    inv_0 U257 ( .x(n78), .a(n192) );
    inv_2 U258 ( .x(n79), .a(n78) );
    nand2_3 U259 ( .x(n99), .a(A[9]), .b(B[9]) );
    inv_2 U26 ( .x(n128), .a(n334) );
    oai21_1 U260 ( .x(n80), .a(n156), .b(n89), .c(n57) );
    inv_4 U261 ( .x(n216), .a(A[6]) );
    inv_2 U262 ( .x(n235), .a(A[11]) );
    nand2_1 U263 ( .x(n149), .a(A[11]), .b(B[11]) );
    inv_0 U264 ( .x(n115), .a(n233) );
    nand2i_6 U265 ( .x(n327), .a(n86), .b(n224) );
    nand2i_2 U266 ( .x(n281), .a(n282), .b(n283) );
    oai211_1 U267 ( .x(n95), .a(n93), .b(n83), .c(n88), .d(B[21]) );
    nand2_1 U268 ( .x(n346), .a(n309), .b(n83) );
    aoi21_1 U269 ( .x(n167), .a(n298), .b(n83), .c(n299) );
    inv_2 U27 ( .x(n247), .a(B[27]) );
    oai211_4 U270 ( .x(n82), .a(n184), .b(n120), .c(n290), .d(n345) );
    nand2i_2 U271 ( .x(n311), .a(A[2]), .b(n214) );
    nand2_2 U272 ( .x(n130), .a(B[2]), .b(A[2]) );
    inv_0 U273 ( .x(n84), .a(n149) );
    inv_2 U274 ( .x(n85), .a(n84) );
    nor2_0 U275 ( .x(n90), .a(A[0]), .b(B[0]) );
    buf_2 U276 ( .x(n86), .a(A[31]) );
    buf_16 U277 ( .x(n88), .a(A[31]) );
    buf_16 U278 ( .x(n87), .a(A[31]) );
    nor2i_5 U279 ( .x(n126), .a(n127), .b(n128) );
    ao21_1 U28 ( .x(n296), .a(n170), .b(n247), .c(n128) );
    nor2_5 U280 ( .x(n165), .a(A[12]), .b(B[12]) );
    nor2i_3 U281 ( .x(n166), .a(n167), .b(n168) );
    exor2_3 U282 ( .x(SUM[5]), .a(n191), .b(n177) );
    exor2_3 U283 ( .x(SUM[29]), .a(n196), .b(n197) );
    exor2_3 U284 ( .x(SUM[26]), .a(n200), .b(n126) );
    exnor2_5 U285 ( .x(SUM[24]), .a(n166), .b(n203) );
    exnor2_3 U286 ( .x(SUM[23]), .a(n204), .b(n205) );
    exnor2_3 U287 ( .x(SUM[13]), .a(n107), .b(n144) );
    inv_6 U288 ( .x(n224), .a(B[15]) );
    nand2i_4 U289 ( .x(n225), .a(n165), .b(n226) );
    nand2i_3 U29 ( .x(n303), .a(n296), .b(n200) );
    oai211_4 U290 ( .x(n244), .a(n170), .b(n238), .c(n133), .d(n245) );
    oai21_5 U291 ( .x(n269), .a(n134), .b(n270), .c(n133) );
    exnor2_3 U292 ( .x(n272), .a(n269), .b(n88) );
    nor2i_5 U293 ( .x(n274), .a(n170), .b(n261) );
    aoi22_3 U294 ( .x(n259), .a(B[20]), .b(n88), .c(n87), .d(n264) );
    aoi21_3 U295 ( .x(n290), .a(n88), .b(n291), .c(n292) );
    nand2i_4 U296 ( .x(n293), .a(n251), .b(n294) );
    nand2_2 U297 ( .x(n297), .a(n253), .b(n255) );
    nand2i_4 U298 ( .x(n198), .a(n297), .b(n303) );
    inv_5 U299 ( .x(n168), .a(n262) );
    nand2_1 U30 ( .x(n255), .a(B[26]), .b(n87) );
    ao21_4 U300 ( .x(n195), .a(n208), .b(n311), .c(n313) );
    nand2i_4 U301 ( .x(n315), .a(B[7]), .b(n158) );
    oai211_4 U302 ( .x(n317), .a(n175), .b(n105), .c(n318), .d(n102) );
    nand2i_4 U303 ( .x(n319), .a(B[8]), .b(n220) );
    inv_5 U304 ( .x(n326), .a(n146) );
    nand2_5 U305 ( .x(n200), .a(n329), .b(n254) );
    aoai211_4 U306 ( .x(n196), .a(n52), .b(n329), .c(n170), .d(n333) );
    nand2i_4 U307 ( .x(n335), .a(n128), .b(n200) );
    nand2i_4 U308 ( .x(n199), .a(n322), .b(n335) );
    oai21_4 U309 ( .x(n205), .a(B[23]), .b(n88), .c(n300) );
    inv_2 U31 ( .x(n251), .a(B[28]) );
    inv_5 U310 ( .x(n270), .a(n211) );
    nand2_5 U311 ( .x(n341), .a(n339), .b(n315) );
    inv_5 U312 ( .x(n294), .a(n249) );
    or3i_5 U313 ( .x(n287), .a(n344), .b(n140), .c(n284) );
    nand2i_4 U314 ( .x(n288), .a(n142), .b(n327) );
    or3i_4 U315 ( .x(n340), .a(n192), .b(n103), .c(n277) );
    mux2i_3 U316 ( .x(n91), .d0(n276), .sl(n347), .d1(n272) );
    exor2_5 U317 ( .x(n203), .a(B[24]), .b(n87) );
    exor2_5 U318 ( .x(n197), .a(B[29]), .b(n88) );
    exor2_5 U319 ( .x(n194), .a(B[30]), .b(n88) );
    nand2i_0 U32 ( .x(n295), .a(n251), .b(n294) );
    exor2_5 U320 ( .x(n193), .a(B[31]), .b(n88) );
    nand2_8 U321 ( .x(n146), .a(n71), .b(A[12]) );
    inv_16 U322 ( .x(n170), .a(n87) );
    nand2i_6 U323 ( .x(n262), .a(n170), .b(n306) );
    aoi21_6 U324 ( .x(n120), .a(n121), .b(n122), .c(n87) );
    nand2_8 U325 ( .x(n254), .a(B[25]), .b(n88) );
    nor2i_6 U326 ( .x(n161), .a(n88), .b(n52) );
    nand2i_4 U327 ( .x(n331), .a(n170), .b(n82) );
    nand2i_5 U328 ( .x(n314), .a(B[4]), .b(n219) );
    nand2i_5 U329 ( .x(n231), .a(B[9]), .b(n221) );
    nand2_0 U33 ( .x(n127), .a(n50), .b(n87) );
    nand2i_5 U330 ( .x(n285), .a(A[14]), .b(n237) );
    nor2i_6 U331 ( .x(n122), .a(B[22]), .b(n223) );
    nand2i_5 U332 ( .x(n250), .a(n87), .b(n252) );
    nand2i_4 U333 ( .x(n339), .a(n157), .b(n340) );
    nand2i_4 U334 ( .x(n284), .a(n60), .b(n285) );
    exor2_2 U335 ( .x(SUM[20]), .a(n206), .b(n207) );
    inv_10 U336 ( .x(n184), .a(n171) );
    nand2i_4 U337 ( .x(n345), .a(n170), .b(n119) );
    mux2i_2 U338 ( .x(n96), .d0(n273), .sl(B[22]), .d1(n274) );
    exnor2_3 U339 ( .x(n273), .a(n261), .b(n170) );
    inv_1 U34 ( .x(n182), .a(n317) );
    nand2i_4 U340 ( .x(n59), .a(n72), .b(A[0]) );
    inv_0 U341 ( .x(n347), .a(n239) );
    inv_4 U342 ( .x(n68), .a(B[1]) );
    and2_4 U343 ( .x(n49), .a(A[1]), .b(B[1]) );
    inv_2 U35 ( .x(n215), .a(B[7]) );
    nand2i_2 U36 ( .x(n181), .a(n215), .b(n66) );
    nand2i_2 U37 ( .x(n180), .a(n158), .b(n66) );
    aoi21_1 U38 ( .x(n179), .a(n180), .b(n181), .c(n182) );
    inv_2 U39 ( .x(n234), .a(n71) );
    nand2i_2 U40 ( .x(n325), .a(A[12]), .b(n234) );
    inv_2 U41 ( .x(n238), .a(B[16]) );
    or3i_2 U42 ( .x(n241), .a(n242), .b(n238), .c(n239) );
    inv_2 U43 ( .x(n268), .a(n241) );
    ao21_1 U44 ( .x(n267), .a(n268), .b(n63), .c(n244) );
    inv_0 U45 ( .x(n118), .a(n264) );
    nand2i_3 U46 ( .x(n264), .a(n244), .b(n240) );
    nor2i_1 U47 ( .x(n132), .a(n133), .b(n134) );
    nand2_2 U48 ( .x(n133), .a(B[17]), .b(n86) );
    nand2i_2 U49 ( .x(n242), .a(n88), .b(n243) );
    exor2_2 U5 ( .x(SUM[30]), .a(n174), .b(n194) );
    inv_2 U50 ( .x(n243), .a(B[17]) );
    inv_2 U51 ( .x(n324), .a(n136) );
    nor2i_1 U52 ( .x(n148), .a(n85), .b(n150) );
    nand2i_2 U53 ( .x(n226), .a(B[11]), .b(n235) );
    nand2i_3 U54 ( .x(n261), .a(n183), .b(n262) );
    nor2_1 U56 ( .x(n298), .a(n260), .b(n223) );
    nand2_2 U57 ( .x(n299), .a(n263), .b(n300) );
    nand2i_4 U58 ( .x(n233), .a(n143), .b(n112) );
    inv_2 U59 ( .x(n112), .a(n227) );
    exnor2_3 U6 ( .x(SUM[31]), .a(n172), .b(n193) );
    or3i_4 U60 ( .x(n344), .a(n302), .b(n326), .c(n162) );
    nor2i_0 U61 ( .x(n101), .a(n102), .b(n103) );
    inv_2 U62 ( .x(n102), .a(n55) );
    and2_1 U63 ( .x(n55), .a(A[6]), .b(B[6]) );
    inv_5 U64 ( .x(n103), .a(n308) );
    aoai211_1 U65 ( .x(n190), .a(n217), .b(n218), .c(n321), .d(n178) );
    inv_2 U66 ( .x(n217), .a(A[5]) );
    inv_5 U67 ( .x(n218), .a(B[5]) );
    nand2_2 U68 ( .x(n142), .a(B[14]), .b(A[14]) );
    inv_5 U69 ( .x(n237), .a(B[14]) );
    aoi21_1 U70 ( .x(n111), .a(n112), .b(n109), .c(n113) );
    nand2i_2 U71 ( .x(n227), .a(n164), .b(n108) );
    nor2i_1 U72 ( .x(n113), .a(n159), .b(n160) );
    inv_0 U73 ( .x(n160), .a(n344) );
    inv_0 U74 ( .x(n153), .a(n280) );
    inv_2 U75 ( .x(n221), .a(A[9]) );
    nand2i_2 U76 ( .x(n229), .a(n230), .b(n231) );
    ao21_3 U77 ( .x(n208), .a(n312), .b(n70), .c(n49) );
    inv_2 U78 ( .x(n214), .a(B[2]) );
    inv_2 U79 ( .x(n252), .a(B[25]) );
    inv_0 U8 ( .x(n155), .a(n49) );
    nand2i_4 U80 ( .x(n291), .a(B[24]), .b(n278) );
    nor2i_5 U81 ( .x(n121), .a(B[24]), .b(n246) );
    inv_2 U82 ( .x(n246), .a(B[21]) );
    nor2i_0 U83 ( .x(n169), .a(n170), .b(n83) );
    exnor2_1 U84 ( .x(n275), .a(n83), .b(n170) );
    inv_2 U85 ( .x(n81), .a(n281) );
    inv_2 U86 ( .x(n286), .a(n288) );
    nand2i_2 U87 ( .x(n266), .a(n286), .b(n287) );
    nand2_2 U88 ( .x(n139), .a(B[15]), .b(n87) );
    inv_2 U89 ( .x(n134), .a(n242) );
    inv_2 U9 ( .x(n50), .a(n248) );
    nor2i_3 U90 ( .x(n276), .a(n269), .b(n87) );
    inv_2 U91 ( .x(n292), .a(n300) );
    nand2_2 U92 ( .x(n300), .a(B[23]), .b(n88) );
    inv_2 U93 ( .x(n223), .a(B[23]) );
    nand2_2 U94 ( .x(n263), .a(B[22]), .b(n88) );
    inv_2 U95 ( .x(n309), .a(n260) );
    nand2_2 U96 ( .x(n260), .a(B[21]), .b(B[22]) );
    nand2_2 U97 ( .x(n332), .a(B[29]), .b(n87) );
    inv_2 U98 ( .x(n222), .a(B[29]) );
    and4_4 U99 ( .x(n52), .a(n253), .b(n254), .c(n255), .d(n251) );
endmodule


module ID_test_1_desync ( INT, CLI, PIPEEMPTY, FREEZE, branch_address, 
    branch_sig, Imm, rt_addr, rd_addr, reg_dst, reg_write, mem_to_reg, 
    mem_write, mem_read, IR_opcode_field, IR_function_field, stall, counter, 
    reset, NPC, IR_latched_input, reg_out_A, reg_out_B, reg_write_WB, WB_data, 
    WB_data_old, test_si, test_so, test_se, sync_sel, global_g1, global_g2, 
    Ctrl__Regs_1__en1, Ctrl__Regs_1__en2 );
output [31:0] branch_address;
output [31:0] Imm;
output [4:0] rt_addr;
output [4:0] rd_addr;
output [5:0] IR_opcode_field;
output [5:0] IR_function_field;
output [1:0] counter;
input  [31:0] NPC;
input  [31:0] IR_latched_input;
output [31:0] reg_out_A;
output [31:0] reg_out_B;
input  [31:0] WB_data;
input  [31:0] WB_data_old;
input  INT, FREEZE, reset, reg_write_WB, test_si, test_se, sync_sel, global_g1, 
    global_g2, Ctrl__Regs_1__en1, Ctrl__Regs_1__en2;
output CLI, PIPEEMPTY, branch_sig, reg_dst, reg_write, mem_to_reg, mem_write, 
    mem_read, stall, test_so;
    wire _RegFile_0__0, _RegFile_0__1, _RegFile_0__2, _RegFile_0__3, 
        _RegFile_0__4, _RegFile_0__5, _RegFile_0__6, _RegFile_0__7, 
        _RegFile_0__8, _RegFile_0__9, _RegFile_0__10, _RegFile_0__11, 
        _RegFile_0__12, _RegFile_0__13, _RegFile_0__14, _RegFile_0__15, 
        _RegFile_0__16, _RegFile_0__17, _RegFile_0__18, _RegFile_0__19, 
        _RegFile_0__20, _RegFile_0__21, _RegFile_0__22, _RegFile_0__23, 
        _RegFile_0__24, _RegFile_0__25, _RegFile_0__26, _RegFile_0__27, 
        _RegFile_0__28, _RegFile_0__29, _RegFile_0__30, _RegFile_0__31, 
        _RegFile_1__0, _RegFile_1__1, _RegFile_1__2, _RegFile_1__3, 
        _RegFile_1__4, _RegFile_1__5, _RegFile_1__6, _RegFile_1__7, 
        _RegFile_1__8, _RegFile_1__9, _RegFile_1__10, _RegFile_1__11, 
        _RegFile_1__12, _RegFile_1__13, _RegFile_1__14, _RegFile_1__15, 
        _RegFile_1__16, _RegFile_1__17, _RegFile_1__18, _RegFile_1__19, 
        _RegFile_1__20, _RegFile_1__21, _RegFile_1__22, _RegFile_1__23, 
        _RegFile_1__24, _RegFile_1__25, _RegFile_1__26, _RegFile_1__27, 
        _RegFile_1__28, _RegFile_1__29, _RegFile_1__30, _RegFile_1__31, 
        _RegFile_2__0, _RegFile_2__1, _RegFile_2__2, _RegFile_2__3, 
        _RegFile_2__4, _RegFile_2__5, _RegFile_2__6, _RegFile_2__7, 
        _RegFile_2__8, _RegFile_2__9, _RegFile_2__10, _RegFile_2__11, 
        _RegFile_2__12, _RegFile_2__13, _RegFile_2__14, _RegFile_2__15, 
        _RegFile_2__16, _RegFile_2__17, _RegFile_2__18, _RegFile_2__19, 
        _RegFile_2__20, _RegFile_2__21, _RegFile_2__22, _RegFile_2__23, 
        _RegFile_2__24, _RegFile_2__25, _RegFile_2__26, _RegFile_2__27, 
        _RegFile_2__28, _RegFile_2__29, _RegFile_2__30, _RegFile_2__31, 
        _RegFile_3__0, _RegFile_3__1, _RegFile_3__2, _RegFile_3__3, 
        _RegFile_3__4, _RegFile_3__5, _RegFile_3__6, _RegFile_3__7, 
        _RegFile_3__8, _RegFile_3__9, _RegFile_3__10, _RegFile_3__11, 
        _RegFile_3__12, _RegFile_3__13, _RegFile_3__14, _RegFile_3__15, 
        _RegFile_3__16, _RegFile_3__17, _RegFile_3__18, _RegFile_3__19, 
        _RegFile_3__20, _RegFile_3__21, _RegFile_3__22, _RegFile_3__23, 
        _RegFile_3__24, _RegFile_3__25, _RegFile_3__26, _RegFile_3__27, 
        _RegFile_3__28, _RegFile_3__29, _RegFile_3__30, _RegFile_3__31, 
        _RegFile_4__0, _RegFile_4__1, _RegFile_4__2, _RegFile_4__3, 
        _RegFile_4__4, _RegFile_4__5, _RegFile_4__6, _RegFile_4__7, 
        _RegFile_4__8, _RegFile_4__9, _RegFile_4__10, _RegFile_4__11, 
        _RegFile_4__12, _RegFile_4__13, _RegFile_4__14, _RegFile_4__15, 
        _RegFile_4__16, _RegFile_4__17, _RegFile_4__18, _RegFile_4__19, 
        _RegFile_4__20, _RegFile_4__21, _RegFile_4__22, _RegFile_4__23, 
        _RegFile_4__24, _RegFile_4__25, _RegFile_4__26, _RegFile_4__27, 
        _RegFile_4__28, _RegFile_4__29, _RegFile_4__30, _RegFile_4__31, 
        _RegFile_5__0, _RegFile_5__1, _RegFile_5__2, _RegFile_5__3, 
        _RegFile_5__4, _RegFile_5__5, _RegFile_5__6, _RegFile_5__7, 
        _RegFile_5__8, _RegFile_5__9, _RegFile_5__10, _RegFile_5__11, 
        _RegFile_5__12, _RegFile_5__13, _RegFile_5__14, _RegFile_5__15, 
        _RegFile_5__16, _RegFile_5__17, _RegFile_5__18, _RegFile_5__19, 
        _RegFile_5__20, _RegFile_5__21, _RegFile_5__22, _RegFile_5__23, 
        _RegFile_5__24, _RegFile_5__25, _RegFile_5__26, _RegFile_5__27, 
        _RegFile_5__28, _RegFile_5__29, _RegFile_5__30, _RegFile_5__31, 
        _RegFile_6__0, _RegFile_6__1, _RegFile_6__2, _RegFile_6__3, 
        _RegFile_6__4, _RegFile_6__5, _RegFile_6__6, _RegFile_6__7, 
        _RegFile_6__8, _RegFile_6__9, _RegFile_6__10, _RegFile_6__11, 
        _RegFile_6__12, _RegFile_6__13, _RegFile_6__14, _RegFile_6__15, 
        _RegFile_6__16, _RegFile_6__17, _RegFile_6__18, _RegFile_6__19, 
        _RegFile_6__20, _RegFile_6__21, _RegFile_6__22, _RegFile_6__23, 
        _RegFile_6__24, _RegFile_6__25, _RegFile_6__26, _RegFile_6__27, 
        _RegFile_6__28, _RegFile_6__29, _RegFile_6__30, _RegFile_6__31, 
        _RegFile_7__0, _RegFile_7__1, _RegFile_7__2, _RegFile_7__3, 
        _RegFile_7__4, _RegFile_7__5, _RegFile_7__6, _RegFile_7__7, 
        _RegFile_7__8, _RegFile_7__9, _RegFile_7__10, _RegFile_7__11, 
        _RegFile_7__12, _RegFile_7__13, _RegFile_7__14, _RegFile_7__15, 
        _RegFile_7__16, _RegFile_7__17, _RegFile_7__18, _RegFile_7__19, 
        _RegFile_7__20, _RegFile_7__21, _RegFile_7__22, _RegFile_7__23, 
        _RegFile_7__24, _RegFile_7__25, _RegFile_7__26, _RegFile_7__27, 
        _RegFile_7__28, _RegFile_7__29, _RegFile_7__30, _RegFile_7__31, 
        _RegFile_8__0, _RegFile_8__1, _RegFile_8__2, _RegFile_8__3, 
        _RegFile_8__4, _RegFile_8__5, _RegFile_8__6, _RegFile_8__7, 
        _RegFile_8__8, _RegFile_8__9, _RegFile_8__10, _RegFile_8__11, 
        _RegFile_8__12, _RegFile_8__13, _RegFile_8__14, _RegFile_8__15, 
        _RegFile_8__16, _RegFile_8__17, _RegFile_8__18, _RegFile_8__19, 
        _RegFile_8__20, _RegFile_8__21, _RegFile_8__22, _RegFile_8__23, 
        _RegFile_8__24, _RegFile_8__25, _RegFile_8__26, _RegFile_8__27, 
        _RegFile_8__28, _RegFile_8__29, _RegFile_8__30, _RegFile_8__31, 
        _RegFile_9__0, _RegFile_9__1, _RegFile_9__2, _RegFile_9__3, 
        _RegFile_9__4, _RegFile_9__5, _RegFile_9__6, _RegFile_9__7, 
        _RegFile_9__8, _RegFile_9__9, _RegFile_9__10, _RegFile_9__11, 
        _RegFile_9__12, _RegFile_9__13, _RegFile_9__14, _RegFile_9__15, 
        _RegFile_9__16, _RegFile_9__17, _RegFile_9__18, _RegFile_9__19, 
        _RegFile_9__20, _RegFile_9__21, _RegFile_9__22, _RegFile_9__23, 
        _RegFile_9__24, _RegFile_9__25, _RegFile_9__26, _RegFile_9__27, 
        _RegFile_9__28, _RegFile_9__29, _RegFile_9__30, _RegFile_9__31, 
        _RegFile_10__0, _RegFile_10__1, _RegFile_10__2, _RegFile_10__3, 
        _RegFile_10__4, _RegFile_10__5, _RegFile_10__6, _RegFile_10__7, 
        _RegFile_10__8, _RegFile_10__9, _RegFile_10__10, _RegFile_10__11, 
        _RegFile_10__12, _RegFile_10__13, _RegFile_10__14, _RegFile_10__15, 
        _RegFile_10__16, _RegFile_10__17, _RegFile_10__18, _RegFile_10__19, 
        _RegFile_10__20, _RegFile_10__21, _RegFile_10__22, _RegFile_10__23, 
        _RegFile_10__24, _RegFile_10__25, _RegFile_10__26, _RegFile_10__27, 
        _RegFile_10__28, _RegFile_10__29, _RegFile_10__30, _RegFile_10__31, 
        _RegFile_11__0, _RegFile_11__1, _RegFile_11__2, _RegFile_11__3, 
        _RegFile_11__4, _RegFile_11__5, _RegFile_11__6, _RegFile_11__7, 
        _RegFile_11__8, _RegFile_11__9, _RegFile_11__10, _RegFile_11__11, 
        _RegFile_11__12, _RegFile_11__13, _RegFile_11__14, _RegFile_11__15, 
        _RegFile_11__16, _RegFile_11__17, _RegFile_11__18, _RegFile_11__19, 
        _RegFile_11__20, _RegFile_11__21, _RegFile_11__22, _RegFile_11__23, 
        _RegFile_11__24, _RegFile_11__25, _RegFile_11__26, _RegFile_11__27, 
        _RegFile_11__28, _RegFile_11__29, _RegFile_11__30, _RegFile_11__31, 
        _RegFile_12__0, _RegFile_12__1, _RegFile_12__2, _RegFile_12__3, 
        _RegFile_12__4, _RegFile_12__5, _RegFile_12__6, _RegFile_12__7, 
        _RegFile_12__8, _RegFile_12__9, _RegFile_12__10, _RegFile_12__11, 
        _RegFile_12__12, _RegFile_12__13, _RegFile_12__14, _RegFile_12__15, 
        _RegFile_12__16, _RegFile_12__17, _RegFile_12__18, _RegFile_12__19, 
        _RegFile_12__20, _RegFile_12__21, _RegFile_12__22, _RegFile_12__23, 
        _RegFile_12__24, _RegFile_12__25, _RegFile_12__26, _RegFile_12__27, 
        _RegFile_12__28, _RegFile_12__29, _RegFile_12__30, _RegFile_12__31, 
        _RegFile_13__0, _RegFile_13__1, _RegFile_13__2, _RegFile_13__3, 
        _RegFile_13__4, _RegFile_13__5, _RegFile_13__6, _RegFile_13__7, 
        _RegFile_13__8, _RegFile_13__9, _RegFile_13__10, _RegFile_13__11, 
        _RegFile_13__12, _RegFile_13__13, _RegFile_13__14, _RegFile_13__15, 
        _RegFile_13__16, _RegFile_13__17, _RegFile_13__18, _RegFile_13__19, 
        _RegFile_13__20, _RegFile_13__21, _RegFile_13__22, _RegFile_13__23, 
        _RegFile_13__24, _RegFile_13__25, _RegFile_13__26, _RegFile_13__27, 
        _RegFile_13__28, _RegFile_13__29, _RegFile_13__30, _RegFile_13__31, 
        _RegFile_14__0, _RegFile_14__1, _RegFile_14__2, _RegFile_14__3, 
        _RegFile_14__4, _RegFile_14__5, _RegFile_14__6, _RegFile_14__7, 
        _RegFile_14__8, _RegFile_14__9, _RegFile_14__10, _RegFile_14__11, 
        _RegFile_14__12, _RegFile_14__13, _RegFile_14__14, _RegFile_14__15, 
        _RegFile_14__16, _RegFile_14__17, _RegFile_14__18, _RegFile_14__19, 
        _RegFile_14__20, _RegFile_14__21, _RegFile_14__22, _RegFile_14__23, 
        _RegFile_14__24, _RegFile_14__25, _RegFile_14__26, _RegFile_14__27, 
        _RegFile_14__28, _RegFile_14__29, _RegFile_14__30, _RegFile_14__31, 
        _RegFile_15__0, _RegFile_15__1, _RegFile_15__2, _RegFile_15__3, 
        _RegFile_15__4, _RegFile_15__5, _RegFile_15__6, _RegFile_15__7, 
        _RegFile_15__8, _RegFile_15__9, _RegFile_15__10, _RegFile_15__11, 
        _RegFile_15__12, _RegFile_15__13, _RegFile_15__14, _RegFile_15__15, 
        _RegFile_15__16, _RegFile_15__17, _RegFile_15__18, _RegFile_15__19, 
        _RegFile_15__20, _RegFile_15__21, _RegFile_15__22, _RegFile_15__23, 
        _RegFile_15__24, _RegFile_15__25, _RegFile_15__26, _RegFile_15__27, 
        _RegFile_15__28, _RegFile_15__29, _RegFile_15__30, _RegFile_15__31, 
        _RegFile_16__0, _RegFile_16__1, _RegFile_16__2, _RegFile_16__3, 
        _RegFile_16__4, _RegFile_16__5, _RegFile_16__6, _RegFile_16__7, 
        _RegFile_16__8, _RegFile_16__9, _RegFile_16__10, _RegFile_16__11, 
        _RegFile_16__12, _RegFile_16__13, _RegFile_16__14, _RegFile_16__15, 
        _RegFile_16__16, _RegFile_16__17, _RegFile_16__18, _RegFile_16__19, 
        _RegFile_16__20, _RegFile_16__21, _RegFile_16__22, _RegFile_16__23, 
        _RegFile_16__24, _RegFile_16__25, _RegFile_16__26, _RegFile_16__27, 
        _RegFile_16__28, _RegFile_16__29, _RegFile_16__30, _RegFile_16__31, 
        _RegFile_17__0, _RegFile_17__1, _RegFile_17__2, _RegFile_17__3, 
        _RegFile_17__4, _RegFile_17__5, _RegFile_17__6, _RegFile_17__7, 
        _RegFile_17__8, _RegFile_17__9, _RegFile_17__10, _RegFile_17__11, 
        _RegFile_17__12, _RegFile_17__13, _RegFile_17__14, _RegFile_17__15, 
        _RegFile_17__16, _RegFile_17__17, _RegFile_17__18, _RegFile_17__19, 
        _RegFile_17__20, _RegFile_17__21, _RegFile_17__22, _RegFile_17__23, 
        _RegFile_17__24, _RegFile_17__25, _RegFile_17__26, _RegFile_17__27, 
        _RegFile_17__28, _RegFile_17__29, _RegFile_17__30, _RegFile_17__31, 
        _RegFile_18__0, _RegFile_18__1, _RegFile_18__2, _RegFile_18__3, 
        _RegFile_18__4, _RegFile_18__5, _RegFile_18__6, _RegFile_18__7, 
        _RegFile_18__8, _RegFile_18__9, _RegFile_18__10, _RegFile_18__11, 
        _RegFile_18__12, _RegFile_18__13, _RegFile_18__14, _RegFile_18__15, 
        _RegFile_18__16, _RegFile_18__17, _RegFile_18__18, _RegFile_18__19, 
        _RegFile_18__20, _RegFile_18__21, _RegFile_18__22, _RegFile_18__23, 
        _RegFile_18__24, _RegFile_18__25, _RegFile_18__26, _RegFile_18__27, 
        _RegFile_18__28, _RegFile_18__29, _RegFile_18__30, _RegFile_18__31, 
        _RegFile_19__0, _RegFile_19__1, _RegFile_19__2, _RegFile_19__3, 
        _RegFile_19__4, _RegFile_19__5, _RegFile_19__6, _RegFile_19__7, 
        _RegFile_19__8, _RegFile_19__9, _RegFile_19__10, _RegFile_19__11, 
        _RegFile_19__12, _RegFile_19__13, _RegFile_19__14, _RegFile_19__15, 
        _RegFile_19__16, _RegFile_19__17, _RegFile_19__18, _RegFile_19__19, 
        _RegFile_19__20, _RegFile_19__21, _RegFile_19__22, _RegFile_19__23, 
        _RegFile_19__24, _RegFile_19__25, _RegFile_19__26, _RegFile_19__27, 
        _RegFile_19__28, _RegFile_19__29, _RegFile_19__30, _RegFile_19__31, 
        _RegFile_20__0, _RegFile_20__1, _RegFile_20__2, _RegFile_20__3, 
        _RegFile_20__4, _RegFile_20__5, _RegFile_20__6, _RegFile_20__7, 
        _RegFile_20__8, _RegFile_20__9, _RegFile_20__10, _RegFile_20__11, 
        _RegFile_20__12, _RegFile_20__13, _RegFile_20__14, _RegFile_20__15, 
        _RegFile_20__16, _RegFile_20__17, _RegFile_20__18, _RegFile_20__19, 
        _RegFile_20__20, _RegFile_20__21, _RegFile_20__22, _RegFile_20__23, 
        _RegFile_20__24, _RegFile_20__25, _RegFile_20__26, _RegFile_20__27, 
        _RegFile_20__28, _RegFile_20__29, _RegFile_20__30, _RegFile_20__31, 
        _RegFile_21__0, _RegFile_21__1, _RegFile_21__2, _RegFile_21__3, 
        _RegFile_21__4, _RegFile_21__5, _RegFile_21__6, _RegFile_21__7, 
        _RegFile_21__8, _RegFile_21__9, _RegFile_21__10, _RegFile_21__11, 
        _RegFile_21__12, _RegFile_21__13, _RegFile_21__14, _RegFile_21__15, 
        _RegFile_21__16, _RegFile_21__17, _RegFile_21__18, _RegFile_21__19, 
        _RegFile_21__20, _RegFile_21__21, _RegFile_21__22, _RegFile_21__23, 
        _RegFile_21__24, _RegFile_21__25, _RegFile_21__26, _RegFile_21__27, 
        _RegFile_21__28, _RegFile_21__29, _RegFile_21__30, _RegFile_21__31, 
        _RegFile_22__0, _RegFile_22__1, _RegFile_22__2, _RegFile_22__3, 
        _RegFile_22__4, _RegFile_22__5, _RegFile_22__6, _RegFile_22__7, 
        _RegFile_22__8, _RegFile_22__9, _RegFile_22__10, _RegFile_22__11, 
        _RegFile_22__12, _RegFile_22__13, _RegFile_22__14, _RegFile_22__15, 
        _RegFile_22__16, _RegFile_22__17, _RegFile_22__18, _RegFile_22__19, 
        _RegFile_22__20, _RegFile_22__21, _RegFile_22__22, _RegFile_22__23, 
        _RegFile_22__24, _RegFile_22__25, _RegFile_22__26, _RegFile_22__27, 
        _RegFile_22__28, _RegFile_22__29, _RegFile_22__30, _RegFile_22__31, 
        _RegFile_23__0, _RegFile_23__1, _RegFile_23__2, _RegFile_23__3, 
        _RegFile_23__4, _RegFile_23__5, _RegFile_23__6, _RegFile_23__7, 
        _RegFile_23__8, _RegFile_23__9, _RegFile_23__10, _RegFile_23__11, 
        _RegFile_23__12, _RegFile_23__13, _RegFile_23__14, _RegFile_23__15, 
        _RegFile_23__16, _RegFile_23__17, _RegFile_23__18, _RegFile_23__19, 
        _RegFile_23__20, _RegFile_23__21, _RegFile_23__22, _RegFile_23__23, 
        _RegFile_23__24, _RegFile_23__25, _RegFile_23__26, _RegFile_23__27, 
        _RegFile_23__28, _RegFile_23__29, _RegFile_23__30, _RegFile_23__31, 
        _RegFile_24__0, _RegFile_24__1, _RegFile_24__2, _RegFile_24__3, 
        _RegFile_24__4, _RegFile_24__5, _RegFile_24__6, _RegFile_24__7, 
        _RegFile_24__8, _RegFile_24__9, _RegFile_24__10, _RegFile_24__11, 
        _RegFile_24__12, _RegFile_24__13, _RegFile_24__14, _RegFile_24__15, 
        _RegFile_24__16, _RegFile_24__17, _RegFile_24__18, _RegFile_24__19, 
        _RegFile_24__20, _RegFile_24__21, _RegFile_24__22, _RegFile_24__23, 
        _RegFile_24__24, _RegFile_24__25, _RegFile_24__26, _RegFile_24__27, 
        _RegFile_24__28, _RegFile_24__29, _RegFile_24__30, _RegFile_24__31, 
        _RegFile_25__0, _RegFile_25__1, _RegFile_25__2, _RegFile_25__3, 
        _RegFile_25__4, _RegFile_25__5, _RegFile_25__6, _RegFile_25__7, 
        _RegFile_25__8, _RegFile_25__9, _RegFile_25__10, _RegFile_25__11, 
        _RegFile_25__12, _RegFile_25__13, _RegFile_25__14, _RegFile_25__15, 
        _RegFile_25__16, _RegFile_25__17, _RegFile_25__18, _RegFile_25__19, 
        _RegFile_25__20, _RegFile_25__21, _RegFile_25__22, _RegFile_25__23, 
        _RegFile_25__24, _RegFile_25__25, _RegFile_25__26, _RegFile_25__27, 
        _RegFile_25__28, _RegFile_25__29, _RegFile_25__30, _RegFile_25__31, 
        _RegFile_26__0, _RegFile_26__1, _RegFile_26__2, _RegFile_26__3, 
        _RegFile_26__4, _RegFile_26__5, _RegFile_26__6, _RegFile_26__7, 
        _RegFile_26__8, _RegFile_26__9, _RegFile_26__10, _RegFile_26__11, 
        _RegFile_26__12, _RegFile_26__13, _RegFile_26__14, _RegFile_26__15, 
        _RegFile_26__16, _RegFile_26__17, _RegFile_26__18, _RegFile_26__19, 
        _RegFile_26__20, _RegFile_26__21, _RegFile_26__22, _RegFile_26__23, 
        _RegFile_26__24, _RegFile_26__25, _RegFile_26__26, _RegFile_26__27, 
        _RegFile_26__28, _RegFile_26__29, _RegFile_26__30, _RegFile_26__31, 
        _RegFile_27__0, _RegFile_27__1, _RegFile_27__2, _RegFile_27__3, 
        _RegFile_27__4, _RegFile_27__5, _RegFile_27__6, _RegFile_27__7, 
        _RegFile_27__8, _RegFile_27__9, _RegFile_27__10, _RegFile_27__11, 
        _RegFile_27__12, _RegFile_27__13, _RegFile_27__14, _RegFile_27__15, 
        _RegFile_27__16, _RegFile_27__17, _RegFile_27__18, _RegFile_27__19, 
        _RegFile_27__20, _RegFile_27__21, _RegFile_27__22, _RegFile_27__23, 
        _RegFile_27__24, _RegFile_27__25, _RegFile_27__26, _RegFile_27__27, 
        _RegFile_27__28, _RegFile_27__29, _RegFile_27__30, _RegFile_27__31, 
        _RegFile_28__0, _RegFile_28__1, _RegFile_28__2, _RegFile_28__3, 
        _RegFile_28__4, _RegFile_28__5, _RegFile_28__6, _RegFile_28__7, 
        _RegFile_28__8, _RegFile_28__9, _RegFile_28__10, _RegFile_28__11, 
        _RegFile_28__12, _RegFile_28__13, _RegFile_28__14, _RegFile_28__15, 
        _RegFile_28__16, _RegFile_28__17, _RegFile_28__18, _RegFile_28__19, 
        _RegFile_28__20, _RegFile_28__21, _RegFile_28__22, _RegFile_28__23, 
        _RegFile_28__24, _RegFile_28__25, _RegFile_28__26, _RegFile_28__27, 
        _RegFile_28__28, _RegFile_28__29, _RegFile_28__30, _RegFile_28__31, 
        _RegFile_29__0, _RegFile_29__1, _RegFile_29__2, _RegFile_29__3, 
        _RegFile_29__4, _RegFile_29__5, _RegFile_29__6, _RegFile_29__7, 
        _RegFile_29__8, _RegFile_29__9, _RegFile_29__10, _RegFile_29__11, 
        _RegFile_29__12, _RegFile_29__13, _RegFile_29__14, _RegFile_29__15, 
        _RegFile_29__16, _RegFile_29__17, _RegFile_29__18, _RegFile_29__19, 
        _RegFile_29__20, _RegFile_29__21, _RegFile_29__22, _RegFile_29__23, 
        _RegFile_29__24, _RegFile_29__25, _RegFile_29__26, _RegFile_29__27, 
        _RegFile_29__28, _RegFile_29__29, _RegFile_29__30, _RegFile_29__31, 
        _RegFile_30__0, _RegFile_30__1, _RegFile_30__2, _RegFile_30__3, 
        _RegFile_30__4, _RegFile_30__5, _RegFile_30__6, _RegFile_30__7, 
        _RegFile_30__8, _RegFile_30__9, _RegFile_30__10, _RegFile_30__11, 
        _RegFile_30__12, _RegFile_30__13, _RegFile_30__14, _RegFile_30__15, 
        _RegFile_30__16, _RegFile_30__17, _RegFile_30__18, _RegFile_30__19, 
        _RegFile_30__20, _RegFile_30__21, _RegFile_30__22, _RegFile_30__23, 
        _RegFile_30__24, _RegFile_30__25, _RegFile_30__26, _RegFile_30__27, 
        _RegFile_30__28, _RegFile_30__29, _RegFile_30__30, _RegFile_30__31, 
        _RegFile_31__0, _RegFile_31__1, _RegFile_31__2, _RegFile_31__3, 
        _RegFile_31__4, _RegFile_31__5, _RegFile_31__6, _RegFile_31__7, 
        _RegFile_31__8, _RegFile_31__9, _RegFile_31__10, _RegFile_31__11, 
        _RegFile_31__12, _RegFile_31__13, _RegFile_31__14, _RegFile_31__15, 
        _RegFile_31__16, _RegFile_31__17, _RegFile_31__18, _RegFile_31__19, 
        _RegFile_31__20, _RegFile_31__21, _RegFile_31__22, _RegFile_31__23, 
        _RegFile_31__24, _RegFile_31__25, _RegFile_31__26, _RegFile_31__27, 
        _RegFile_31__28, _RegFile_31__29, _RegFile_31__30, _RegFile_31__31, 
        n804, n896, n694, n332, n331, N468, N467, N466, N465, N464, N463, N462, 
        N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, 
        N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, 
        N437, n857, n339, n848, n337, n802, N535, N534, N533, N532, N531, N530, 
        N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, 
        N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, 
        N505, N504, CLI_reg__m2s, n2641, n953, n4386, Cause_Reg_reg_0__m2s, 
        n2642, Cause_Reg_0, n627, Cause_Reg_reg_10__m2s, n2652, n618, 
        Cause_Reg_10, n617, Cause_Reg_reg_11__m2s, n2653, Cause_Reg_11, n616, 
        Cause_Reg_reg_12__m2s, n2654, Cause_Reg_12, n615, 
        Cause_Reg_reg_13__m2s, n2655, Cause_Reg_13, n614, 
        Cause_Reg_reg_14__m2s, n2656, Cause_Reg_14, n613, 
        Cause_Reg_reg_15__m2s, n2657, n952, Cause_Reg_15, n612, 
        Cause_Reg_reg_16__m2s, n2658, Cause_Reg_16, n611, 
        Cause_Reg_reg_17__m2s, n2659, Cause_Reg_17, n610, 
        Cause_Reg_reg_18__m2s, n2660, Cause_Reg_18, n609, 
        Cause_Reg_reg_19__m2s, n2661, Cause_Reg_19, n608, Cause_Reg_reg_1__m2s, 
        n2643, Cause_Reg_1, n626, Cause_Reg_reg_20__m2s, n2662, Cause_Reg_20, 
        n607, Cause_Reg_reg_21__m2s, n2663, Cause_Reg_21, n606, 
        Cause_Reg_reg_22__m2s, n2664, Cause_Reg_22, n605, 
        Cause_Reg_reg_23__m2s, n2665, Cause_Reg_23, n604, 
        Cause_Reg_reg_24__m2s, n2666, Cause_Reg_24, n603, 
        Cause_Reg_reg_25__m2s, n2667, Cause_Reg_25, n602, 
        Cause_Reg_reg_26__m2s, n2668, Cause_Reg_26, n601, 
        Cause_Reg_reg_27__m2s, n2669, Cause_Reg_27, n600, 
        Cause_Reg_reg_28__m2s, n2670, Cause_Reg_28, n599, 
        Cause_Reg_reg_29__m2s, n2671, n954, Cause_Reg_29, n598, 
        Cause_Reg_reg_2__m2s, n2644, Cause_Reg_2, n625, Cause_Reg_reg_30__m2s, 
        n2672, Cause_Reg_30, n597, Cause_Reg_reg_31__m2s, n2673, Cause_Reg_31, 
        n596, Cause_Reg_reg_3__m2s, n2645, Cause_Reg_3, n624, 
        Cause_Reg_reg_4__m2s, n2646, Cause_Reg_4, n623, Cause_Reg_reg_5__m2s, 
        n2647, Cause_Reg_5, n622, Cause_Reg_reg_6__m2s, n2648, Cause_Reg_6, 
        n621, Cause_Reg_reg_7__m2s, n2649, Cause_Reg_7, n620, 
        Cause_Reg_reg_8__m2s, n2650, Cause_Reg_8, n619, Cause_Reg_reg_9__m2s, 
        n2651, Cause_Reg_9, EPC_reg_0__m2s, n2674, EPC_0, n595, 
        EPC_reg_10__m2s, n2684, EPC_9, EPC_10, n593, EPC_reg_11__m2s, n2685, 
        EPC_11, n592, EPC_reg_12__m2s, n2686, EPC_12, n591, EPC_reg_13__m2s, 
        n2687, n951, EPC_13, n590, EPC_reg_14__m2s, n2688, EPC_14, n589, 
        EPC_reg_15__m2s, n2689, EPC_15, n588, EPC_reg_16__m2s, n2690, EPC_16, 
        n587, EPC_reg_17__m2s, n2691, EPC_17, n586, EPC_reg_18__m2s, n2692, 
        EPC_18, n585, EPC_reg_19__m2s, n2693, EPC_19, n584, EPC_reg_1__m2s, 
        n2675, EPC_1, n594, EPC_reg_20__m2s, n2694, EPC_20, n583, 
        EPC_reg_21__m2s, n2695, EPC_21, n4383, EPC_reg_22__m2s, n2696, EPC_22, 
        n4382, EPC_reg_23__m2s, n2697, EPC_23, n4381, EPC_reg_24__m2s, n2698, 
        EPC_24, n4380, EPC_reg_25__m2s, n2699, EPC_25, n4379, EPC_reg_26__m2s, 
        n2700, EPC_26, n582, EPC_reg_27__m2s, n2701, n955, EPC_27, n581, 
        EPC_reg_28__m2s, n2702, EPC_28, n580, EPC_reg_29__m2s, n2703, EPC_29, 
        n579, EPC_reg_2__m2s, n2676, EPC_2, n4385, EPC_reg_30__m2s, n2704, 
        EPC_30, n662, EPC_reg_31__m2s, _EPC_reg_31_net69891, EPC_31, n578, 
        EPC_reg_3__m2s, n2677, EPC_3, n4384, EPC_reg_4__m2s, n2678, EPC_4, 
        n577, EPC_reg_5__m2s, n2679, EPC_5, n576, EPC_reg_6__m2s, n2680, EPC_6, 
        n575, EPC_reg_7__m2s, n2681, EPC_7, n574, EPC_reg_8__m2s, n2682, EPC_8, 
        n573, EPC_reg_9__m2s, n2683, n572, IR_function_field_reg_0__m2s, n3764, 
        n1859, IR_function_field_reg_1__m2s, n3765, n1860, 
        IR_function_field_reg_2__m2s, n3766, n1861, 
        IR_function_field_reg_3__m2s, n3767, n950, n1862, 
        IR_function_field_reg_4__m2s, n3768, n1863, 
        IR_function_field_reg_5__m2s, n3769, n4378, IR_opcode_field_reg_0__m2s, 
        n3770, n911, n4454, n4377, IR_opcode_field_reg_1__m2s, n3771, n4453, 
        n4376, IR_opcode_field_reg_2__m2s, n3772, n4452, n4375, 
        IR_opcode_field_reg_3__m2s, n3773, n4374, IR_opcode_field_reg_4__m2s, 
        n3774, n4373, IR_opcode_field_reg_5__m2s, n3775, n4372, Imm_reg_0__m2s, 
        n3791, n914, N6328, n813, Imm_reg_10__m2s, n3801, n873, N6348, n4371, 
        Imm_reg_11__m2s, n3802, n949, N6350, n786, Imm_reg_12__m2s, n3803, 
        N6352, n779, Imm_reg_13__m2s, n3804, n916, N6354, n4370, 
        Imm_reg_14__m2s, n3805, N6356, n647, Imm_reg_15__m2s, n3806, N6358, 
        n829, Imm_reg_16__m2s, n3807, N6360, n648, Imm_reg_17__m2s, n3808, 
        N6362, n803, Imm_reg_18__m2s, n3809, N6364, n778, Imm_reg_19__m2s, 
        n3810, N6366, n775, Imm_reg_1__m2s, n3792, n915, n720, Imm_reg_20__m2s, 
        n3811, N6368, n732, Imm_reg_21__m2s, n3812, N6370, n649, 
        Imm_reg_22__m2s, n3813, n789, Imm_reg_23__m2s, n3814, n912, n827, 
        Imm_reg_24__m2s, n3815, N6376, n654, Imm_reg_25__m2s, n3816, n816, 
        Imm_reg_26__m2s, n3817, N6380, n735, Imm_reg_27__m2s, n3818, N6382, 
        n765, Imm_reg_28__m2s, n3819, N6384, n696, Imm_reg_29__m2s, n3820, 
        N6386, n762, Imm_reg_2__m2s, n3793, N6332, n870, Imm_reg_30__m2s, 
        n3821, N6388, n701, Imm_reg_31__m2s, n3822, N6390, n4369, 
        Imm_reg_3__m2s, n3794, N6334, n886, Imm_reg_4__m2s, n3795, N6336, n871, 
        Imm_reg_5__m2s, n3796, N6338, n845, Imm_reg_6__m2s, n3797, N6340, n643, 
        Imm_reg_7__m2s, n3798, N6342, n734, Imm_reg_8__m2s, n3799, N6344, n872, 
        Imm_reg_9__m2s, n3800, N6346, n554, n1547, n1382, n1767, n3936, n3940, 
        n3285, n1830, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3294, 
        n1983, n1801, n1399, n3295, n1960, n1778, n3296, n1961, n1779, n3297, 
        n1962, n1780, n3298, n1963, n1781, n3299, n1964, n1782, n3300, n1965, 
        n1783, n3301, n1966, n1784, n3302, n1967, n1785, n3303, n1968, n1786, 
        n3304, n1969, n1787, n1520, n1515, n1521, n3305, n1970, n1788, n3306, 
        n1971, n1789, n3307, n1972, n1790, n3308, n1973, n1791, n3309, n1974, 
        n1792, n3310, n1975, n1793, n3311, n1976, n1794, n3312, n1977, n1795, 
        n3313, n1978, n1796, n3314, n1979, n1797, n1518, n1519, n3315, n1980, 
        n1798, n1768, n3935, n3317, n1829, n3318, n3319, n3320, n3321, n3322, 
        n3323, n3324, n796, n795, ___cell__36997_net129977, 
        ___cell__36997_net129979, ___cell__36997_net130187, n3326, n1959, 
        n3327, n1936, n3328, n1937, n3329, n1938, n3330, n1939, n3331, n1940, 
        n3332, n1941, n3333, n1942, n3334, n1943, n3335, n1944, n693, n3336, 
        n1945, n3337, n1946, n3338, n1947, n3339, n1948, n3340, n1949, n3341, 
        n1950, n3342, n1951, n3343, n1952, n3344, n1953, n3345, n1954, n704, 
        ___cell__36997_net126612, n3346, n1955, n959, n957, n3347, n1956, n946, 
        n939, n1769, n3927, n3349, n1828, n3350, n3351, n3352, n3353, n1262, 
        n1263, n3354, n3355, n3356, n3358, n1935, n3359, n1912, n3360, n1913, 
        n3361, n1914, n3362, n1915, n3363, n1916, n3364, n1917, n1261, n1314, 
        n883, n564, n3365, n1918, n3366, n1919, n3367, n1920, n3368, n1921, 
        n3369, n1922, n3370, n1923, n3371, n1924, n3372, n1925, n3373, n1926, 
        n3374, n1927, n3944, WB_index_0, WB_index_4, WB_index_1, n3375, n1928, 
        n3376, n1929, n3377, n1930, n3378, n1931, n958, n945, n3379, n1932, 
        n1770, n3937, n3939, n3381, n1827, n3382, n3383, n3958, n3943, n3928, 
        n3384, n3385, n3386, n3387, n3388, n3390, n1911, n3391, n1888, n3392, 
        n1889, n3393, n1890, n3394, n1891, n3942, n3929, n3395, n1892, n3396, 
        n1893, n3397, n1894, n3398, n1895, n3399, n1896, n3400, n1897, n3401, 
        n1898, n3402, n1899, n3403, n1900, n3404, n1901, n3941, n3405, n1902, 
        n3406, n1903, n3407, n1904, n3408, n1905, n3409, n1906, n3410, n1907, 
        n3411, n1908, n1771, n3413, n1857, n3414, WB_index_2, WB_index_3, 
        n3415, n3416, n3417, n3418, n3419, n691, n3420, n692, n3422, n2631, 
        n3423, n2608, n3424, n2609, n3425, n2610, n3925, n3426, n2611, n3427, 
        n2612, n3428, n2613, n3429, n2614, n3430, n2615, n3431, n2616, n3432, 
        n2617, n3433, n2618, n3434, n2619, n3435, n2620, n3938, n3926, n3436, 
        n2621, n3437, n2622, n3438, n2623, n3439, n2624, n3440, n2625, n3441, 
        n2626, n3442, n2627, n3443, n2628, n1741, n3445, n1856, 
        ___cell__6171_net27367, n3446, n3447, n3448, n3449, n3450, n3451, 
        n3452, n3454, n2607, n3455, n2584, n3456, n2585, n3457, n2586, n3458, 
        n2587, n3459, n2588, n3460, n2589, n3461, n2590, n3462, n2591, n3463, 
        n2592, n3464, n2593, n3465, n2594, n3466, n2595, n3467, n2596, n3468, 
        n2597, n3469, n2598, n3470, n2599, n3471, n2600, n3472, n2601, n3473, 
        n2602, n3474, n2603, n3475, n2604, n920, n989, n3934, n555, n1742, 
        n3477, n1855, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3486, 
        n2583, n750, n1602, n1395, n1511, n3487, n2560, n3488, n2561, n3489, 
        n2562, n3490, n2563, n3491, n2564, n3492, n2565, n3493, n2566, n3494, 
        n2567, n3495, n2568, n3496, n2569, n1600, n1411, n3497, n2570, n3498, 
        n2571, n3499, n2572, n3500, n2573, n3501, n2574, n3502, n2575, n3503, 
        n2576, n3504, n2577, n3505, n2578, n3506, n2579, n1648, n1392, n3507, 
        n2580, n1743, n3509, n1854, n3510, n3511, n3512, n3513, n3514, n3515, 
        n3516, n1646, n1354, n3518, n2559, n3519, n2536, n3520, n2537, n3521, 
        n2538, n3522, n2539, n3523, n2540, n3524, n2541, n3525, n2542, n3526, 
        n2543, n3527, n2544, n1740, n3528, n2545, n3529, n2546, n3530, n2547, 
        n3531, n2548, n3532, n2549, n3533, n2550, n3534, n2551, n3535, n2552, 
        n3536, n2553, n3537, n2554, n1512, n1303, n3538, n2555, n3539, n2556, 
        n1744, n3541, n1853, n3542, n3543, n3544, n3545, n3546, n3547, n1644, 
        n1400, n3548, n3550, n2535, n3551, n2512, n3552, n2513, n3553, n2514, 
        n3554, n2515, n3555, n2516, n3556, n2517, n3557, n2518, n3558, n2519, 
        n1642, n1406, n3559, n2520, n3560, n2521, n3561, n2522, n3562, n2523, 
        n3563, n2524, n3564, n2525, n3565, n2526, n3566, n2527, n3567, n2528, 
        n3568, n2529, n1640, n1359, n3569, n2530, n3570, n2531, n978, n983, 
        n3571, n2532, n1745, n3573, n1852, n3574, n3575, n3576, n3577, n1638, 
        n1304, n3578, n3579, n3580, n924, n937, n3582, n2511, n3583, n2488, 
        n3584, n2489, n3585, n2490, n3586, n2491, n3587, n2492, n1636, n1376, 
        n3588, n2493, n3589, n2494, n3590, n2495, n3591, n2496, n3592, n2497, 
        n3593, n2498, n3594, n2499, n3595, n2500, n3596, n2501, n3597, n2502, 
        n1634, n1349, n3598, n2503, n3599, n2504, n3600, n2505, n3601, n2506, 
        n3602, n2507, n977, n923, n3603, n2508, n925, n1746, n3605, n1851, 
        n1632, n1340, n927, n936, n3606, n3607, n3608, n3609, n3610, n3611, 
        n3612, n3614, n2487, n3615, n2464, n1630, n1383, n3616, n2465, n3617, 
        n2466, n3618, n2467, n3619, n2468, n3620, n2469, n3621, n2470, n3622, 
        n2471, n3623, n2472, n3624, n2473, n3625, n2474, n1628, n1381, n3626, 
        n2475, n3627, n2476, n3628, n2477, n3629, n2478, n3630, n2479, n3631, 
        n2480, n3632, n2481, n3633, n2482, n3634, n2483, n3635, n2484, n1626, 
        n1379, n1747, n3637, n1848, n3638, n3639, n3640, n3641, n3642, n3643, 
        n3644, n3646, n2415, n1624, n1374, n3647, n2392, n3648, n2393, n3649, 
        n2394, n3650, n2395, n3651, n2396, n930, n987, n3652, n2397, n3653, 
        n2398, n3654, n2399, n3655, n2400, n1622, n1403, n3656, n2401, n3657, 
        n2402, n3658, n2403, n3659, n2404, n3660, n2405, n3661, n2406, n3662, 
        n2407, n3663, n2408, n3664, n2409, n3665, n2410, n1620, n1409, n3666, 
        n2411, n3667, n2412, n929, n1750, n3669, n1837, n3670, n3671, n3672, 
        n3673, n3674, n1618, n1338, n3675, n3676, n1603, n1601, n3678, n2151, 
        n3679, n2128, n3680, n2129, n3681, n2130, n3682, n2131, n3683, n2132, 
        n3684, n2133, n3945, n3933, opcode_of_MEM_4, n1616, n1361, n3685, 
        n2134, n3686, n2135, n3687, n2136, n3688, n2137, n3689, n2138, n962, 
        n984, n3690, n2139, n3691, n2140, n3692, n2141, n3693, n2142, n1614, 
        n1346, n3694, n2143, n3695, n2144, n3696, n2145, n3697, n2146, n3698, 
        n2147, n963, n3699, n2148, n1761, n3701, n1826, n690, n3702, n688, 
        n1612, n1357, n3703, n3704, n3705, n687, n3706, n689, n3707, n3708, 
        n1800, n1772, n3930, n3733, n1423, n1424, _current_IR_reg_1_net49291, 
        n800, ___cell__36997_net130681, n801, n1610, n1343, current_IR_1, 
        n3734, n1421, n1422, n3736, n1418, n1419, n3738, n631, n1596, n3740, 
        n630, n1593, n3741, n629, n1592, n3742, n632, n1597, n3746, n569, 
        n1413, n3748, n645, n1330, n3749, n1332, n1333, n1608, n1363, n3756, 
        n1323, n1324, n3759, n1318, n1319, n1066, n1718, n1065, 
        ___cell__36997_net126621, n1074, n642, n1107, n2637, n1098, n2635, 
        n1086, n2636, n3778, n1085, n1302, n1305, n1097, n1716, n1485, n1069, 
        n1719, n3784, n1061, n1076, n1070, n1802, n3785, n1775, n1063, n917, 
        n990, n1077, n561, n1122, n671, n705, n1606, ___cell__36997_net129389, 
        n1133, n558, n3790, n1132, n918, n988, n919, n1213, net150785, n1650, 
        n1773, n856, n340, n1682, n3891, n1000, n1484, 
        ___cell__36997_net127190, n1307, n679, n913, n1728, reg_dst_of_EX_0, 
        n1530, n1529, n993, n991, n992, n1726, n1725, n2638, n3931, n1727, 
        n1729, n843, n847, n1532, n1552, n1553, n1595, n1594, current_IR_7, 
        n1534, n1531, n1536, n3967, n1316, n851, n1535, n1439, n1311, n1461, 
        n1287, n1283, current_IR_0, current_IR_2, current_IR_4, current_IR_17, 
        current_IR_24, current_IR_27, n1686, n1417, n1416, n1415, n1414, n1412, 
        n1331, n1527, n1526, n1525, n1524, ___cell__36997_net129786, n556, 
        opcode_of_MEM_2, n628, n3946, opcode_of_MEM_1, n3947, n1691, n772, 
        n637, n1410, ___cell__36997_net129354, n640, n1380, n1647, n1645, 
        n1643, n1641, n1639, n1637, n1635, n1633, n1071, n1631, n1629, n1627, 
        n1625, n1623, n1621, n1619, n1617, n1615, n1613, n1735, n1687, n1575, 
        n1611, n1609, n1607, n1604, n1605, n1799, n1599, n1514, n1803, n932, 
        n1734, n1574, n1573, n967, n922, n966, n975, n974, n976, n968, n947, 
        n938, n969, n948, n964, n1858, n926, n972, n986, n961, n892, n934, 
        n921, n970, n971, n981, n980, n935, n985, n979, n982, n973, n956, n650, 
        n882, n1517, n881, n653, n1367, n1368, n335, n879, net152024, n728, 
        ___cell__36997_net130705, net148858, net148913, n1328, n1326, n3978, 
        n668, ___cell__36997_net129247, n1277, n1325, n1688, n1083, n672, 
        n1384, n1385, n673, n1386, n1387, n674, n1339, reg_dst_of_EX_3, n702, 
        n1336, n1337, n698, n675, ___cell__36997_net130713, N6039, n333, n676, 
        N6040, n1522, n1523, n1445, n744, n3948, ___cell__36997_net125928, 
        n1516, n680, n1559, ___cell__36997_net129626, n3954, n682, n782, n1466, 
        n1706, n639, n1014, n663, n1703, n1701, n1702, n1710, n1128, n1020, 
        n1003, n1024, n1344, n1144, n797, net150625, n683, n850, n684, n1377, 
        n1378, n685, n686, n1390, n1397, reg_dst_of_MEM_2, n1724, n1371, n1366, 
        n1657, reg_dst_of_MEM_0, reg_dst_of_MEM_1, n3953, n3952, n695, n1161, 
        net150626, n1181, n1165, n1149, n1169, n1225, n1533, reg_dst_of_MEM_3, 
        reg_dst_of_MEM_4, n1209, n1229, n1201, n1157, n1189, n1177, n1245, 
        n1205, n1153, n1173, n1089, n559, n697, n1431, n1432, n1430, n1096, 
        net149679, n780, n787, n1704, n1372, n1130, n994, n1028, n699, n1347, 
        n1072, n560, n1009, n1348, n1459, n855, n714, n747, n1026, n998, n1006, 
        n1722, n2634, n1143, n1498, n863, n700, n1456, n1457, n1458, n1444, 
        n1455, N6723, n995, n1126, n3737, n565, n1427, n1562, n634, n1695, 
        n756, n822, n1446, ___cell__36997_net125989, ___cell__36997_net129381, 
        ___cell__36997_net125941, ___cell__36997_net129378, n859, n757, n752, 
        n3760, n566, n1442, reg_dst_of_EX_4, n1570, n1571, n708, n703, n1731, 
        n3998, n1565, n1685, n739, n815, n3752, n567, n1260, n1428, n1315, 
        n1111, n707, N6718, n3985, ___cell__36997_net130580, n996, n709, n710, 
        n1694, n715, n761, n1434, n724, n3747, n568, n1449, N6721, n1777, 
        n1238, n769, n736, n1087, n1141, n1355, n1356, n711, n1429, n753, 
        n3745, n570, n825, n1737, n826, n1451, n1500, N5378, n1075, n807, n759, 
        n760, current_IR_23, n1264, n1265, n712, n823, n1437, n713, n1487, 
        n846, n3743, n571, ___cell__36997_net129632, n812, net148863, N6731, 
        n1004, n1404, N6719, n1131, n841, n1081, n767, 
        ___cell__36997_net130567, n1082, n1491, n1467, n1435, n717, n1548, 
        n718, n719, n1581, n1321, ___cell__36997_net130125, n721, n861, n755, 
        n1560, n1561, n1080, n722, n3763, n633, n725, n1137, 
        ___cell__36997_net130709, N5449, n1101, n1100, n3853, n1139, n1138, 
        n1140, n810, n865, n726, n1543, N6722, n636, n1127, N6729, n999, n3990, 
        n1730, n3783, n1774, n1059, n1040, n1079, n1043, n3782, n1057, n3786, 
        n3789, n3992, n1112, N6725, n1243, n1038, n1078, current_IR_30, n2707, 
        n729, n1134, n742, n1312, n837, n731, n771, ___cell__36997_net130572, 
        n2706, n1473, n1090, n1689, n1477, n733, n1280, n799, n1110, n1479, 
        n1585, n1582, n1438, n738, n791, n3753, n646, net149236, current_IR_31, 
        n1463, n1578, n666, n1327, n740, n1590, n741, n1454, n1591, n745, n743, 
        n3735, n651, n1420, n1266, n1267, n835, ___cell__36997_net130214, 
        N6023, n811, n1228, N5361, N6028, n1200, N5355, N6022, n1696, n1557, 
        n334, n3744, n652, n1008, n1732, n1538, n1736, n1483, n1476, n1489, 
        n1440, n1441, n1443, n746, n1545, n1313, reg_dst_of_EX_2, n1697, n748, 
        n884, net149681, n1084, n3755, n659, n1495, N5382, n1174, n766, N5424, 
        n1182, N5436, n1216, N5434, n1214, N5432, n1190, N5430, n1154, N5420, 
        n1580, n1568, n3754, n661, n1178, N5425, n1268, n2705, n1091, n1447, 
        ___cell__36997_net130306, n1468, n1469, n1436, n3852, n1142, n665, 
        n1693, n338, n1352, n1044, n1219, n1350, n768, n660, n1183, N6735, 
        n1010, N6732, n1005, n1167, n3757, N6733, n1007, N6734, n1163, n1341, 
        n1342, n1106, n1488, n832, n777, n1222, N6036, n1295, n1334, net149680, 
        n1335, n3901, n1672, n1212, N5364, n862, N6031, n1272, n1566, n1448, 
        n1108, net152025, n716, n1236, n1508, n758, net151343, n867, n868, 
        current_IR_19, n1016, n1733, n1037, n764, n3922, n1649, n763, n1309, 
        n887, n1480, n1554, n1497, N6047, n1804, ___cell__36997_net129624, 
        ___cell__36997_net129625, n3777, n1094, n1113, n1114, n1152, N5352, 
        n895, N6019, IR_latched_1, n3959, ___cell__36997_net129524, n3911, 
        n1662, n3949, n3950, n3750, current_IR_18, n1329, n3969, n773, n1317, 
        n842, n854, n1237, ___cell__36997_net126604, n1278, n1598, n2633, 
        n1471, n1499, N5446, n776, n1147, N6045, ___cell__36997_net129239, 
        n1300, N6029, n783, n3842, n784, n1223, n1221, n1220, n1067, n3902, 
        n1671, n1490, n785, n1699, n1684, n655, n818, n3989, n1539, 
        _counter_reg_0_net48671, ___cell__36997_net127189, 
        _counter_reg_1_net48651, n790, n4011, n798, ___cell__36997_net129477, 
        n1109, n1717, n1258, n3762, n658, n1310, n3955, n878, n889, n808, 
        n1496, N6048, n3780, n809, n1051, IR_latched_8, n1049, n1537, 
        ___cell__36997_net127155, n1492, n1240, N6021, n1198, n1505, n1217, 
        n1510, n1041, n1073, n1255, net148865, N6020, n1250, n1501, n1194, 
        n1507, n1136, n1293, net148916, n1294, n1275, n1276, n1282, 
        ___cell__36997_net130217, n849, current_IR_3, n1546, n1032, n1551, 
        n866, n1253, n737, n1588, slot_num_0, n1589, slot_num_1, n1576, 
        IR_latched_13, n1714, n557, n3972, n1047, n817, n820, n3758, n852, 
        n1068, n1426, n3781, n1055, n1425, n1712, n1713, n1474, n1475, n1690, 
        n1039, n2708, n1035, n1036, n834, net151366, n836, n840, n1462, n670, 
        n1104, n1776, n888, n1308, n3776, n1095, n1464, n1567, n1088, n3788, 
        n3986, IR_latched_5, n1541, n3779, n3892, n1681, n1011, IR_latched_11, 
        n1172, N5356, n1270, n3847, n1193, n1192, n1195, n1711, n1708, n1705, 
        n1218, N5366, n3968, n3823, n3827, n1239, n1241, n1242, n3826, n1254, 
        n1256, n1257, IR_latched_12, n1284, n1285, n1549, n1540, n1279, n1550, 
        n1482, n1544, n997, n1018, n1196, n1235, N5447, n1150, n1233, n1191, 
        n1159, n1247, n1175, n1179, n1252, n3913, n1660, n1203, n1171, n1031, 
        n1215, n1231, n638, n1211, n1155, n1227, n1001, n1207, n1248, N5445, 
        n3956, n860, n3845, n1232, n1234, n3995, n1042, n1045, n1046, n1048, 
        n1680, n1050, n1052, n1058, n1060, n1064, n1062, IR_latched_0, n3893, 
        n1493, ___cell__36997_net129654, n2632, n669, n3897, n1676, n562, 
        n1433, IR_latched_15, n1579, n3923, opcode_of_MEM_3, N6744, n1023, 
        ___cell__36997_net129657, n1146, n1187, n1503, n1199, n1504, n1251, 
        n1502, n1180, N5368, n1297, n1188, N5362, n1506, n1156, N5351, n1301, 
        n1509, N5353, N5354, n1168, N5359, N6026, n1160, N5367, N6034, n1224, 
        N5363, N6030, n1587, n1151, N5371, N6038, n1053, n1054, n1033, N6745, 
        n678, n1025, n3910, n1663, n1542, n1002, n3957, n1118, N6743, n1022, 
        n1120, n1056, net148915, n1322, n1700, n1572, n3787, N5440, 
        ___cell__36997_net130212, n1290, N5442, n1286, n1162, N5435, n1158, 
        N5419, n1166, N5433, n1170, N5427, n1230, N5429, n1206, N5428, n3900, 
        n1673, n1226, N5431, n1202, N5423, N5437, n1185, n3971, n3974, n3965, 
        n3970, n3964, n1034, n1099, n1103, n1105, n1115, n1116, n1117, n1119, 
        n1249, n1121, n1123, n1124, n1125, n3851, n1145, n3844, n1148, n3825, 
        n3824, n3840, n3838, n1164, N6044, n3832, n3829, n3841, n3835, n3828, 
        n3833, n1204, n3843, n1208, n1210, n3837, n3924, N5377, n3839, n3836, 
        n3834, n3831, n1246, n1244, n3850, n1184, n1281, n1292, n1296, n3895, 
        n1678, n1345, n1351, n1353, n1358, n1360, n1364, n1365, n1369, n1370, 
        n1373, n1388, n1389, n1393, n1394, n1398, n1401, n1402, n1405, n1407, 
        n1408, n3915, n1658, IR_latched_14, current_IR_9, current_IR_8, n1450, 
        n1452, n1478, n1486, n1273, N5381, N6042, N5369, n1563, n1569, n3751, 
        n657, n3761, n656, n3421, n2630, n3444, n2629, n3453, n2606, n3476, 
        n2605, n3485, n2582, n3508, n2581, n3517, n2558, N5439, n3540, n2557, 
        n3549, n2534, n3572, n2533, n3581, n2510, n3604, n2509, n3613, n2486, 
        n3636, n2485, n2717, n2462, n1850, n2740, n2461, n2749, n2438, n1849, 
        n3904, n1669, n2772, n2437, n3645, n2414, n3668, n2413, n2781, n2390, 
        n1847, n2804, n2389, n2813, n2366, n1846, n2836, n2365, n2845, n2342, 
        n1845, n2868, n2341, n2877, n2318, n1844, n2900, n2317, n2909, n2294, 
        n1843, n2932, n2293, n2941, n2270, n1842, n2964, n2269, n2973, n2246, 
        n1841, n2996, n2245, n3005, n2222, n1840, n3028, n2221, n3037, n2198, 
        n1839, n3909, n1664, n3060, n2197, n3069, n2174, n1838, n3092, n2173, 
        n3677, n2150, n3700, n2149, n3101, n2126, n1836, n3124, n2125, n3133, 
        n2102, n1835, n3156, n2101, n3165, n2078, n1834, n3188, n2077, n3197, 
        n2054, n1833, n3220, n2053, n3229, n2030, n1832, n3252, n2029, n3261, 
        n2006, n1831, n3284, n2005, n3293, n1982, n3316, n1981, n3325, n1958, 
        n3348, n1957, n3357, n1934, n3380, n1933, n3389, n1910, n3412, n1909, 
        n3710, n1887, n3709, n1886, n3732, n1885, n3731, n1884, n3730, n1883, 
        n3729, n1882, n3728, n1881, n3727, n1880, n3726, n1879, n3725, n1878, 
        n3724, n1877, n3723, n1876, n3722, n1875, n3721, n1874, n3720, n1873, 
        n3719, n1872, n3718, n1871, n3717, n1870, n3716, n1869, n3715, n1868, 
        n3714, n1867, n3713, n1866, n3712, n1865, n3711, n1864, n1558, 
        ___cell__36997_net130191, n1707, n3903, n1670, n1709, n1654, n1748, 
        n1749, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n3932, 
        n3908, n1665, n1759, n1760, n1762, n1763, n1764, n1765, n1766, n336, 
        n3917, n1655, n3980, n3983, n3973, n3962, n3963, n3981, n3960, n3951, 
        n1494, n1259, n1470, n1481, n1093, n1465, n1460, n1723, n3739, n1513, 
        n1721, N13832, opcode_of_WB_5, n3889, n3887, n3890, n1683, n635, n3899, 
        n1674, n667, n3898, n1675, n749, n3997, n1197, n4005, n831, n3921, 
        n1651, IR_latched_2, n1715, n3984, n1375, n641, 
        ___cell__36997_net126005, n794, n3977, n3830, n1176, N5357, n1269, 
        n833, n4007, n644, n3987, n3988, current_IR_21, N5426, N6025, n853, 
        n3912, n1661, n3854, n1135, n3996, n3991, current_IR_29, n4432, n681, 
        N5358, ___cell__36997_net129384, n1362, n1453, n1698, n1564, n3846, 
        n3848, n3993, N5438, N5370, N6037, _branch_address_reg_31_net46811, 
        N5450, n664, n792, N5365, n1299, N6032, n4457, N5380, n1271, N5375, 
        N5441, n1288, n1289, N5448, n3849, n1186, n1291, n793, n805, n3966, 
        N6033, N6043, n4004, n4003, n3999, n4001, n4000, n4002, current_IR_6, 
        N6027, N5360, n3982, n4442, n3905, N5443, N6046, n4008, N6024, n770, 
        reg_dst_of_EX_1, n3906, n1667, n563, n4009, n4012, n4455, n4456, n4390, 
        n4458, n4394, n4410, n1668, n4434, n4422, n4430, n4388, n4392, n4396, 
        n4398, n3918, n4400, n3894, n4402, n3907, n4404, n3916, n4406, n3896, 
        n4408, n3914, n4412, n4414, n4416, n4418, n4420, n4424, n4426, n4428, 
        n1659, n4436, n4438, n3920, n4440, n3919, n4444, n4446, n4448, n4450, 
        n1274, n3961, N5422, N5421, N5444, N5376, N5372, N6041, N5374, N6749, 
        ___cell__36997_net127210, ___cell__36997_net129388, n1528, n677, 
        IR_latched_10, n1102, n910, N6049, n3979, n1677, N6742, n1021, N6746, 
        n1027, n1656, n1666, N6748, n1030, n909, n1679, N6739, n1015, n1029, 
        N6747, n1017, N6740, N6741, n1019, N6738, n1013, IR_latched_9, n1653, 
        N6736, n1652, n1129, n1306, N6724, N6737, n1012, current_IR_10, N6727, 
        n1396, N6730, N6728, n1391, IR_latched_3, N6726, N6720, IR_latched_4, 
        n2640, intr_slot, n1092, delay_slot, n1739, n824, n2709, n2710, n2711, 
        n2712, n2713, n2714, n2715, n1692, n2716, n2718, n2463, n2719, n2440, 
        n2720, n2441, n2721, n2442, n2722, n2443, n2723, n2444, n2724, n2445, 
        n2725, n2446, n2726, n2447, n2727, n2448, n2728, n2449, n2729, n2450, 
        n2730, n2451, n2731, n2452, n2732, n2453, n2733, n2454, n2734, n2455, 
        n2735, n2456, n2736, n2457, n2737, n2458, n2738, n2459, n2739, n2460, 
        n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2750, n2439, 
        n2751, n2416, n2752, n2417, n2753, n2418, n2754, n2419, n2755, n2420, 
        n2756, n2421, n2757, n2422, n1584, n2758, n2423, n2759, n2424, n2760, 
        n2425, n2761, n2426, n2762, n2427, n2763, n2428, n2764, n2429, n2765, 
        n2430, n2766, n2431, n2767, n2432, n1583, n2768, n2433, n2769, n2434, 
        n2770, n2435, n2771, n2436, n928, n2773, n2774, n2775, n2776, n2777, 
        n2778, n2779, n2780, n2782, n2391, n2783, n2368, n2784, n2369, n2785, 
        n2370, n2786, n2371, n2787, n2372, n1320, n1586, n2788, n2373, n2789, 
        n2374, n2790, n2375, n2791, n2376, n2792, n2377, n2793, n2378, n2794, 
        n2379, n2795, n2380, n2796, n2381, n2797, n2382, n2798, n2383, n2799, 
        n2384, n2800, n2385, n2801, n2386, n2802, n2387, n2803, n2388, n2805, 
        n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2814, n2367, n2815, 
        n2344, n2816, n2345, n2817, n2346, n2818, n2347, n2819, n2348, n2820, 
        n2349, n2821, n2350, n2822, n2351, n2823, n2352, n2824, n2353, n2825, 
        n2354, n2826, n2355, n2827, n2356, n2828, n2357, n2829, n2358, n2830, 
        n2359, n2831, n2360, n2832, n2361, n2833, n2362, n2834, n2363, n2835, 
        n2364, n931, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, 
        n2846, n2343, n2847, n2320, n2848, n2321, n2849, n2322, n2850, n2323, 
        n2851, n2324, n2852, n2325, n2853, n2326, n2854, n2327, n2855, n2328, 
        n2856, n2329, n2857, n2330, n2858, n2331, opcode_of_MEM_5, n2859, 
        n2332, n2860, n2333, n2861, n2334, n2862, n2335, n2863, n2336, n2864, 
        n2337, n2865, n2338, n2866, n2339, n2867, n2340, n2869, n2870, n2871, 
        n2872, n2873, n2874, n2875, n2876, n2878, n2319, n2879, n2296, n2880, 
        n2297, n2881, n2298, n2882, n2299, n2883, n2300, n2884, n2301, n2885, 
        n2302, n2886, n2303, n2887, n2304, n2888, n2305, n2889, n2306, n2890, 
        n2307, n2891, n2308, n2892, n2309, n2893, n2310, n2894, n2311, n2895, 
        n2312, n2896, n2313, n2897, n2314, n2898, n2315, n2899, n2316, n933, 
        n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2910, n2295, 
        n2911, n2272, n2912, n2273, n2913, n2274, n2914, n2275, n2915, n2276, 
        n2916, n2277, n2917, n2278, n2918, n2279, n2919, n2280, n3888, n2920, 
        n2281, n2921, n2282, n2922, n2283, n2923, n2284, n2924, n2285, n2925, 
        n2286, n2926, n2287, n2927, n2288, n2928, n2289, n2929, n2290, n2930, 
        n2291, n2931, n2292, n2933, n2934, n2935, n2936, n2937, n2938, n2939, 
        n2940, n2942, n2271, n2943, n2248, n2944, n2249, n2945, n2250, n2946, 
        n2251, n2947, n2252, n2948, n2253, n2949, n2254, n2950, n2255, n2951, 
        n2256, n2952, n2257, n2953, n2258, n2954, n2259, n2955, n2260, n2956, 
        n2261, n2957, n2262, n2958, n2263, n2959, n2264, n2960, n2265, n2961, 
        n2266, n2962, n2267, n2963, n2268, n2965, n2966, n2967, n2968, n2969, 
        n2970, n2971, n2972, n2974, n2247, n2975, n2224, n2976, n2225, n2977, 
        n2226, n2978, n2227, n2979, n2228, n2980, n2229, n2981, n2230, n2982, 
        n2231, n2983, n2232, n2984, n2233, n2985, n2234, n2986, n2235, n2987, 
        n2236, n2988, n2237, n2989, n2238, n2990, n2239, n2991, n2240, n2992, 
        n2241, n2993, n2242, n2994, n2243, n2995, n2244, n2997, n2998, n2999, 
        n3000, n3001, n1720, n3002, n3003, n3004, n3006, n2223, n3007, n2200, 
        n3008, n2201, n3009, n2202, n3010, n2203, n3011, n2204, n3012, n2205, 
        n3013, n2206, n3014, n2207, n3015, n2208, n3016, n2209, n3017, n2210, 
        n3018, n2211, n3019, n2212, n3020, n2213, n3021, n2214, n3022, n2215, 
        n3023, n2216, n3024, n2217, n3025, n2218, n3026, n2219, n3027, n2220, 
        n3029, n3030, n3031, n3032, N5379, n3033, n3034, n3035, n3036, n3038, 
        n2199, n3039, n2176, n3040, n2177, n3041, n2178, n3042, n2179, n3043, 
        n2180, n1738, n3044, n2181, n3045, n2182, n3046, n2183, n3047, n2184, 
        n3048, n2185, n3049, n2186, n3050, n2187, n3051, n2188, n3052, n2189, 
        n3053, n2190, n3054, n2191, n3055, n2192, n3056, n2193, n3057, n2194, 
        n3058, n2195, n965, n3059, n2196, n3061, n3062, n1472, n3063, n3064, 
        n3065, n3066, n3067, n3068, n3070, n2175, n3071, n2152, n3072, n2153, 
        n3073, n2154, n3074, n2155, n3075, n2156, n3076, n2157, n3077, n2158, 
        n3078, n2159, n3079, n2160, n3080, n2161, n3081, n2162, n3082, n2163, 
        n3083, n2164, n3084, n2165, n3085, n2166, n3086, n2167, n3087, n2168, 
        n3088, n2169, n3089, n2170, n3090, n2171, n3091, n2172, n3093, n1298, 
        N6035, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3102, n2127, 
        n3103, n2104, n3104, n2105, n3105, n2106, n3106, n2107, n3107, n2108, 
        n3108, n2109, n3109, n2110, n3110, n2111, n3111, n2112, n3112, n2113, 
        n3113, n2114, n3114, n2115, N6018, n3115, n2116, n3116, n2117, n3117, 
        n2118, n3118, n2119, n3119, n2120, n3120, n2121, n3121, n2122, n3122, 
        n2123, n3123, n2124, n940, N5373, n3125, n3126, n3127, n3128, n3129, 
        n3130, n3131, n3132, n3134, n2103, n3135, n2080, n3136, n2081, n3137, 
        n2082, n3138, n2083, n3139, n2084, n3140, n2085, n3141, n2086, n3142, 
        n2087, n3143, n2088, n3144, n2089, n3145, n2090, n3146, n2091, n3147, 
        n2092, n3148, n2093, n3149, n2094, n3150, n2095, n3151, n2096, n3152, 
        n2097, n3153, n2098, n3154, n2099, n3155, n2100, n941, n3157, n3158, 
        n3159, n3160, n3161, n3162, n3163, n3164, n3166, n2079, n3167, n2056, 
        n3168, n2057, n3169, n2058, n3170, n2059, n3171, n2060, n3172, n2061, 
        n3173, n2062, n3174, n2063, n3175, n2064, n3176, n2065, n3177, n2066, 
        n3178, n2067, n3179, n2068, n3180, n2069, n3181, n2070, n3182, n2071, 
        n3183, n2072, n3184, n2073, n3185, n2074, n3186, n2075, n3187, n2076, 
        n942, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3198, 
        n2055, n3199, n2032, n3200, n2033, n3201, n2034, n3202, n2035, n3203, 
        n2036, n3204, n2037, n2639, n3205, n2038, n3206, n2039, n3207, n2040, 
        n3208, n2041, n3209, n2042, n3210, n2043, n3211, n2044, n3212, n2045, 
        n3213, n2046, n3214, n2047, n3215, n2048, n3216, n2049, n3217, n2050, 
        n3218, n2051, n3219, n2052, n943, n3221, n3222, n3223, n3224, n3225, 
        n3226, n3227, n3228, n960, n3230, n2031, n3231, n2008, n3232, n2009, 
        n3233, n2010, n3234, n2011, n3235, n2012, n3236, n2013, n3237, n2014, 
        n3238, n2015, n3239, n2016, n3240, n2017, n3241, n2018, n3242, n2019, 
        n3243, n2020, n3244, n2021, n3245, n2022, n3246, n2023, n3247, n2024, 
        n3248, n2025, n3249, n2026, n3250, n2027, n3251, n2028, n944, n3253, 
        n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3262, n2007, n3263, 
        n1984, n3264, n1985, n3265, n1986, n3266, n1987, n3267, n1988, n3268, 
        n1989, n3269, n1990, n3270, n1991, n3271, n1992, n3272, n1993, n3273, 
        n1994, n3274, n1995, n3275, n1996, n3276, n1997, n3277, n1998, n3278, 
        n1999, n3279, n2000, n3280, n2001, n3281, n2002, n3282, n2003, n3283, 
        n2004, WB_index_reg_0__m2s, WB_index_reg_1__m2s, WB_index_reg_2__m2s, 
        WB_index_reg_3__m2s, WB_index_reg_4__m2s, _RegFile_reg_0__0__m2s, 
        n4368, _RegFile_reg_0__10__m2s, _RegFile_reg_0__11__m2s, 
        _RegFile_reg_0__12__m2s, _RegFile_reg_0__13__m2s, 
        _RegFile_reg_0__14__m2s, _RegFile_reg_0__15__m2s, 
        _RegFile_reg_0__16__m2s, _RegFile_reg_0__17__m2s, 
        _RegFile_reg_0__18__m2s, _RegFile_reg_0__19__m2s, 
        _RegFile_reg_0__1__m2s, n4367, _RegFile_reg_0__20__m2s, 
        _RegFile_reg_0__21__m2s, _RegFile_reg_0__22__m2s, 
        _RegFile_reg_0__23__m2s, _RegFile_reg_0__24__m2s, 
        _RegFile_reg_0__25__m2s, _RegFile_reg_0__26__m2s, 
        _RegFile_reg_0__27__m2s, _RegFile_reg_0__28__m2s, 
        _RegFile_reg_0__29__m2s, _RegFile_reg_0__2__m2s, n4366, 
        _RegFile_reg_0__30__m2s, _RegFile_reg_0__31__m2s, 
        _RegFile_reg_0__3__m2s, n4365, _RegFile_reg_0__4__m2s, n4364, 
        _RegFile_reg_0__5__m2s, n4363, _RegFile_reg_0__6__m2s, n4362, 
        _RegFile_reg_0__7__m2s, n4361, _RegFile_reg_0__8__m2s, 
        _RegFile_reg_0__9__m2s, _RegFile_reg_10__0__m2s, n4288, 
        _RegFile_reg_10__10__m2s, _RegFile_reg_10__11__m2s, 
        _RegFile_reg_10__12__m2s, _RegFile_reg_10__13__m2s, 
        _RegFile_reg_10__14__m2s, _RegFile_reg_10__15__m2s, 
        _RegFile_reg_10__16__m2s, _RegFile_reg_10__17__m2s, 
        _RegFile_reg_10__18__m2s, _RegFile_reg_10__19__m2s, 
        _RegFile_reg_10__1__m2s, n4287, _RegFile_reg_10__20__m2s, 
        _RegFile_reg_10__21__m2s, _RegFile_reg_10__22__m2s, 
        _RegFile_reg_10__23__m2s, _RegFile_reg_10__24__m2s, 
        _RegFile_reg_10__25__m2s, _RegFile_reg_10__26__m2s, 
        _RegFile_reg_10__27__m2s, _RegFile_reg_10__28__m2s, 
        _RegFile_reg_10__29__m2s, _RegFile_reg_10__2__m2s, n4286, 
        _RegFile_reg_10__30__m2s, _RegFile_reg_10__31__m2s, 
        _RegFile_reg_10__3__m2s, n4285, _RegFile_reg_10__4__m2s, n4284, 
        _RegFile_reg_10__5__m2s, n4283, _RegFile_reg_10__6__m2s, n4282, 
        _RegFile_reg_10__7__m2s, n4281, _RegFile_reg_10__8__m2s, 
        _RegFile_reg_10__9__m2s, _RegFile_reg_11__0__m2s, n4280, 
        _RegFile_reg_11__10__m2s, _RegFile_reg_11__11__m2s, 
        _RegFile_reg_11__12__m2s, _RegFile_reg_11__13__m2s, 
        _RegFile_reg_11__14__m2s, _RegFile_reg_11__15__m2s, 
        _RegFile_reg_11__16__m2s, _RegFile_reg_11__17__m2s, 
        _RegFile_reg_11__18__m2s, _RegFile_reg_11__19__m2s, 
        _RegFile_reg_11__1__m2s, n4279, _RegFile_reg_11__20__m2s, 
        _RegFile_reg_11__21__m2s, _RegFile_reg_11__22__m2s, 
        _RegFile_reg_11__23__m2s, _RegFile_reg_11__24__m2s, 
        _RegFile_reg_11__25__m2s, _RegFile_reg_11__26__m2s, 
        _RegFile_reg_11__27__m2s, _RegFile_reg_11__28__m2s, 
        _RegFile_reg_11__29__m2s, _RegFile_reg_11__2__m2s, n4278, 
        _RegFile_reg_11__30__m2s, _RegFile_reg_11__31__m2s, 
        _RegFile_reg_11__3__m2s, n4277, _RegFile_reg_11__4__m2s, n4276, 
        _RegFile_reg_11__5__m2s, n4275, _RegFile_reg_11__6__m2s, n4274, 
        _RegFile_reg_11__7__m2s, n4273, _RegFile_reg_11__8__m2s, 
        _RegFile_reg_11__9__m2s, _RegFile_reg_12__0__m2s, n4272, 
        _RegFile_reg_12__10__m2s, _RegFile_reg_12__11__m2s, 
        _RegFile_reg_12__12__m2s, _RegFile_reg_12__13__m2s, 
        _RegFile_reg_12__14__m2s, _RegFile_reg_12__15__m2s, 
        _RegFile_reg_12__16__m2s, _RegFile_reg_12__17__m2s, 
        _RegFile_reg_12__18__m2s, _RegFile_reg_12__19__m2s, 
        _RegFile_reg_12__1__m2s, n4271, _RegFile_reg_12__20__m2s, 
        _RegFile_reg_12__21__m2s, _RegFile_reg_12__22__m2s, 
        _RegFile_reg_12__23__m2s, _RegFile_reg_12__24__m2s, 
        _RegFile_reg_12__25__m2s, _RegFile_reg_12__26__m2s, 
        _RegFile_reg_12__27__m2s, _RegFile_reg_12__28__m2s, 
        _RegFile_reg_12__29__m2s, _RegFile_reg_12__2__m2s, n4270, 
        _RegFile_reg_12__30__m2s, _RegFile_reg_12__31__m2s, 
        _RegFile_reg_12__3__m2s, n4269, _RegFile_reg_12__4__m2s, n4268, 
        _RegFile_reg_12__5__m2s, n4267, _RegFile_reg_12__6__m2s, n4266, 
        _RegFile_reg_12__7__m2s, n4265, _RegFile_reg_12__8__m2s, 
        _RegFile_reg_12__9__m2s, _RegFile_reg_13__0__m2s, n4264, 
        _RegFile_reg_13__10__m2s, _RegFile_reg_13__11__m2s, 
        _RegFile_reg_13__12__m2s, _RegFile_reg_13__13__m2s, 
        _RegFile_reg_13__14__m2s, _RegFile_reg_13__15__m2s, 
        _RegFile_reg_13__16__m2s, _RegFile_reg_13__17__m2s, 
        _RegFile_reg_13__18__m2s, _RegFile_reg_13__19__m2s, 
        _RegFile_reg_13__1__m2s, n4263, _RegFile_reg_13__20__m2s, 
        _RegFile_reg_13__21__m2s, _RegFile_reg_13__22__m2s, 
        _RegFile_reg_13__23__m2s, _RegFile_reg_13__24__m2s, 
        _RegFile_reg_13__25__m2s, _RegFile_reg_13__26__m2s, 
        _RegFile_reg_13__27__m2s, _RegFile_reg_13__28__m2s, 
        _RegFile_reg_13__29__m2s, _RegFile_reg_13__2__m2s, n4262, 
        _RegFile_reg_13__30__m2s, _RegFile_reg_13__31__m2s, 
        _RegFile_reg_13__3__m2s, n4261, _RegFile_reg_13__4__m2s, n4260, 
        _RegFile_reg_13__5__m2s, n4259, _RegFile_reg_13__6__m2s, n4258, 
        _RegFile_reg_13__7__m2s, n4257, _RegFile_reg_13__8__m2s, 
        _RegFile_reg_13__9__m2s, _RegFile_reg_14__0__m2s, n4256, 
        _RegFile_reg_14__10__m2s, _RegFile_reg_14__11__m2s, 
        _RegFile_reg_14__12__m2s, _RegFile_reg_14__13__m2s, 
        _RegFile_reg_14__14__m2s, _RegFile_reg_14__15__m2s, 
        _RegFile_reg_14__16__m2s, _RegFile_reg_14__17__m2s, 
        _RegFile_reg_14__18__m2s, _RegFile_reg_14__19__m2s, 
        _RegFile_reg_14__1__m2s, n4255, _RegFile_reg_14__20__m2s, 
        _RegFile_reg_14__21__m2s, _RegFile_reg_14__22__m2s, 
        _RegFile_reg_14__23__m2s, _RegFile_reg_14__24__m2s, 
        _RegFile_reg_14__25__m2s, _RegFile_reg_14__26__m2s, 
        _RegFile_reg_14__27__m2s, _RegFile_reg_14__28__m2s, 
        _RegFile_reg_14__29__m2s, _RegFile_reg_14__2__m2s, n4254, 
        _RegFile_reg_14__30__m2s, _RegFile_reg_14__31__m2s, 
        _RegFile_reg_14__3__m2s, n4253, _RegFile_reg_14__4__m2s, n4252, 
        _RegFile_reg_14__5__m2s, n4251, _RegFile_reg_14__6__m2s, n4250, 
        _RegFile_reg_14__7__m2s, n4249, _RegFile_reg_14__8__m2s, 
        _RegFile_reg_14__9__m2s, _RegFile_reg_15__0__m2s, n4248, 
        _RegFile_reg_15__10__m2s, _RegFile_reg_15__11__m2s, 
        _RegFile_reg_15__12__m2s, _RegFile_reg_15__13__m2s, 
        _RegFile_reg_15__14__m2s, _RegFile_reg_15__15__m2s, 
        _RegFile_reg_15__16__m2s, _RegFile_reg_15__17__m2s, 
        _RegFile_reg_15__18__m2s, _RegFile_reg_15__19__m2s, 
        _RegFile_reg_15__1__m2s, n4247, _RegFile_reg_15__20__m2s, 
        _RegFile_reg_15__21__m2s, _RegFile_reg_15__22__m2s, 
        _RegFile_reg_15__23__m2s, _RegFile_reg_15__24__m2s, 
        _RegFile_reg_15__25__m2s, _RegFile_reg_15__26__m2s, 
        _RegFile_reg_15__27__m2s, _RegFile_reg_15__28__m2s, 
        _RegFile_reg_15__29__m2s, _RegFile_reg_15__2__m2s, n4246, 
        _RegFile_reg_15__30__m2s, _RegFile_reg_15__31__m2s, 
        _RegFile_reg_15__3__m2s, n4245, _RegFile_reg_15__4__m2s, n4244, 
        _RegFile_reg_15__5__m2s, n4243, _RegFile_reg_15__6__m2s, n4242, 
        _RegFile_reg_15__7__m2s, n4241, _RegFile_reg_15__8__m2s, 
        _RegFile_reg_15__9__m2s, _RegFile_reg_16__0__m2s, n4240, 
        _RegFile_reg_16__10__m2s, _RegFile_reg_16__11__m2s, 
        _RegFile_reg_16__12__m2s, _RegFile_reg_16__13__m2s, 
        _RegFile_reg_16__14__m2s, _RegFile_reg_16__15__m2s, 
        _RegFile_reg_16__16__m2s, _RegFile_reg_16__17__m2s, 
        _RegFile_reg_16__18__m2s, _RegFile_reg_16__19__m2s, 
        _RegFile_reg_16__1__m2s, n4239, _RegFile_reg_16__20__m2s, 
        _RegFile_reg_16__21__m2s, _RegFile_reg_16__22__m2s, 
        _RegFile_reg_16__23__m2s, _RegFile_reg_16__24__m2s, 
        _RegFile_reg_16__25__m2s, _RegFile_reg_16__26__m2s, 
        _RegFile_reg_16__27__m2s, _RegFile_reg_16__28__m2s, 
        _RegFile_reg_16__29__m2s, _RegFile_reg_16__2__m2s, n4238, 
        _RegFile_reg_16__30__m2s, _RegFile_reg_16__31__m2s, 
        _RegFile_reg_16__3__m2s, n4237, _RegFile_reg_16__4__m2s, n4236, 
        _RegFile_reg_16__5__m2s, n4235, _RegFile_reg_16__6__m2s, n4234, 
        _RegFile_reg_16__7__m2s, n4233, _RegFile_reg_16__8__m2s, 
        _RegFile_reg_16__9__m2s, _RegFile_reg_17__0__m2s, n4232, 
        _RegFile_reg_17__10__m2s, _RegFile_reg_17__11__m2s, 
        _RegFile_reg_17__12__m2s, _RegFile_reg_17__13__m2s, 
        _RegFile_reg_17__14__m2s, _RegFile_reg_17__15__m2s, 
        _RegFile_reg_17__16__m2s, _RegFile_reg_17__17__m2s, 
        _RegFile_reg_17__18__m2s, _RegFile_reg_17__19__m2s, 
        _RegFile_reg_17__1__m2s, n4231, _RegFile_reg_17__20__m2s, 
        _RegFile_reg_17__21__m2s, _RegFile_reg_17__22__m2s, 
        _RegFile_reg_17__23__m2s, _RegFile_reg_17__24__m2s, 
        _RegFile_reg_17__25__m2s, _RegFile_reg_17__26__m2s, 
        _RegFile_reg_17__27__m2s, _RegFile_reg_17__28__m2s, 
        _RegFile_reg_17__29__m2s, _RegFile_reg_17__2__m2s, n4230, 
        _RegFile_reg_17__30__m2s, _RegFile_reg_17__31__m2s, 
        _RegFile_reg_17__3__m2s, n4229, _RegFile_reg_17__4__m2s, n4228, 
        _RegFile_reg_17__5__m2s, n4227, _RegFile_reg_17__6__m2s, n4226, 
        _RegFile_reg_17__7__m2s, n4225, _RegFile_reg_17__8__m2s, 
        _RegFile_reg_17__9__m2s, _RegFile_reg_18__0__m2s, n4224, 
        _RegFile_reg_18__10__m2s, _RegFile_reg_18__11__m2s, 
        _RegFile_reg_18__12__m2s, _RegFile_reg_18__13__m2s, 
        _RegFile_reg_18__14__m2s, _RegFile_reg_18__15__m2s, 
        _RegFile_reg_18__16__m2s, _RegFile_reg_18__17__m2s, 
        _RegFile_reg_18__18__m2s, _RegFile_reg_18__19__m2s, 
        _RegFile_reg_18__1__m2s, n4223, _RegFile_reg_18__20__m2s, 
        _RegFile_reg_18__21__m2s, _RegFile_reg_18__22__m2s, 
        _RegFile_reg_18__23__m2s, _RegFile_reg_18__24__m2s, 
        _RegFile_reg_18__25__m2s, _RegFile_reg_18__26__m2s, 
        _RegFile_reg_18__27__m2s, _RegFile_reg_18__28__m2s, 
        _RegFile_reg_18__29__m2s, _RegFile_reg_18__2__m2s, n4222, 
        _RegFile_reg_18__30__m2s, _RegFile_reg_18__31__m2s, 
        _RegFile_reg_18__3__m2s, n4221, _RegFile_reg_18__4__m2s, n4220, 
        _RegFile_reg_18__5__m2s, n4219, _RegFile_reg_18__6__m2s, n4218, 
        _RegFile_reg_18__7__m2s, n4217, _RegFile_reg_18__8__m2s, 
        _RegFile_reg_18__9__m2s, _RegFile_reg_19__0__m2s, n4216, 
        _RegFile_reg_19__10__m2s, _RegFile_reg_19__11__m2s, 
        _RegFile_reg_19__12__m2s, _RegFile_reg_19__13__m2s, 
        _RegFile_reg_19__14__m2s, _RegFile_reg_19__15__m2s, 
        _RegFile_reg_19__16__m2s, _RegFile_reg_19__17__m2s, 
        _RegFile_reg_19__18__m2s, _RegFile_reg_19__19__m2s, 
        _RegFile_reg_19__1__m2s, n4215, _RegFile_reg_19__20__m2s, 
        _RegFile_reg_19__21__m2s, _RegFile_reg_19__22__m2s, 
        _RegFile_reg_19__23__m2s, _RegFile_reg_19__24__m2s, 
        _RegFile_reg_19__25__m2s, _RegFile_reg_19__26__m2s, 
        _RegFile_reg_19__27__m2s, _RegFile_reg_19__28__m2s, 
        _RegFile_reg_19__29__m2s, _RegFile_reg_19__2__m2s, n4214, 
        _RegFile_reg_19__30__m2s, _RegFile_reg_19__31__m2s, 
        _RegFile_reg_19__3__m2s, n4213, _RegFile_reg_19__4__m2s, n4212, 
        _RegFile_reg_19__5__m2s, n4211, _RegFile_reg_19__6__m2s, n4210, 
        _RegFile_reg_19__7__m2s, n4209, _RegFile_reg_19__8__m2s, 
        _RegFile_reg_19__9__m2s, _RegFile_reg_1__0__m2s, n4360, 
        _RegFile_reg_1__10__m2s, _RegFile_reg_1__11__m2s, 
        _RegFile_reg_1__12__m2s, _RegFile_reg_1__13__m2s, 
        _RegFile_reg_1__14__m2s, _RegFile_reg_1__15__m2s, 
        _RegFile_reg_1__16__m2s, _RegFile_reg_1__17__m2s, 
        _RegFile_reg_1__18__m2s, _RegFile_reg_1__19__m2s, 
        _RegFile_reg_1__1__m2s, n4359, _RegFile_reg_1__20__m2s, 
        _RegFile_reg_1__21__m2s, _RegFile_reg_1__22__m2s, 
        _RegFile_reg_1__23__m2s, _RegFile_reg_1__24__m2s, 
        _RegFile_reg_1__25__m2s, _RegFile_reg_1__26__m2s, 
        _RegFile_reg_1__27__m2s, _RegFile_reg_1__28__m2s, 
        _RegFile_reg_1__29__m2s, _RegFile_reg_1__2__m2s, n4358, 
        _RegFile_reg_1__30__m2s, _RegFile_reg_1__31__m2s, 
        _RegFile_reg_1__3__m2s, n4357, _RegFile_reg_1__4__m2s, n4356, 
        _RegFile_reg_1__5__m2s, n4355, _RegFile_reg_1__6__m2s, n4354, 
        _RegFile_reg_1__7__m2s, n4353, _RegFile_reg_1__8__m2s, 
        _RegFile_reg_1__9__m2s, _RegFile_reg_20__0__m2s, n4208, 
        _RegFile_reg_20__10__m2s, _RegFile_reg_20__11__m2s, 
        _RegFile_reg_20__12__m2s, _RegFile_reg_20__13__m2s, 
        _RegFile_reg_20__14__m2s, _RegFile_reg_20__15__m2s, 
        _RegFile_reg_20__16__m2s, _RegFile_reg_20__17__m2s, 
        _RegFile_reg_20__18__m2s, _RegFile_reg_20__19__m2s, 
        _RegFile_reg_20__1__m2s, n4207, _RegFile_reg_20__20__m2s, 
        _RegFile_reg_20__21__m2s, _RegFile_reg_20__22__m2s, 
        _RegFile_reg_20__23__m2s, _RegFile_reg_20__24__m2s, 
        _RegFile_reg_20__25__m2s, _RegFile_reg_20__26__m2s, 
        _RegFile_reg_20__27__m2s, _RegFile_reg_20__28__m2s, 
        _RegFile_reg_20__29__m2s, _RegFile_reg_20__2__m2s, n4206, 
        _RegFile_reg_20__30__m2s, _RegFile_reg_20__31__m2s, 
        _RegFile_reg_20__3__m2s, n4205, _RegFile_reg_20__4__m2s, n4204, 
        _RegFile_reg_20__5__m2s, n4203, _RegFile_reg_20__6__m2s, n4202, 
        _RegFile_reg_20__7__m2s, n4201, _RegFile_reg_20__8__m2s, 
        _RegFile_reg_20__9__m2s, _RegFile_reg_21__0__m2s, n4200, 
        _RegFile_reg_21__10__m2s, _RegFile_reg_21__11__m2s, 
        _RegFile_reg_21__12__m2s, _RegFile_reg_21__13__m2s, 
        _RegFile_reg_21__14__m2s, _RegFile_reg_21__15__m2s, 
        _RegFile_reg_21__16__m2s, _RegFile_reg_21__17__m2s, 
        _RegFile_reg_21__18__m2s, _RegFile_reg_21__19__m2s, 
        _RegFile_reg_21__1__m2s, n4199, _RegFile_reg_21__20__m2s, 
        _RegFile_reg_21__21__m2s, _RegFile_reg_21__22__m2s, 
        _RegFile_reg_21__23__m2s, _RegFile_reg_21__24__m2s, 
        _RegFile_reg_21__25__m2s, _RegFile_reg_21__26__m2s, 
        _RegFile_reg_21__27__m2s, _RegFile_reg_21__28__m2s, 
        _RegFile_reg_21__29__m2s, _RegFile_reg_21__2__m2s, n4198, 
        _RegFile_reg_21__30__m2s, _RegFile_reg_21__31__m2s, 
        _RegFile_reg_21__3__m2s, n4197, _RegFile_reg_21__4__m2s, n4196, 
        _RegFile_reg_21__5__m2s, n4195, _RegFile_reg_21__6__m2s, n4194, 
        _RegFile_reg_21__7__m2s, n4193, _RegFile_reg_21__8__m2s, 
        _RegFile_reg_21__9__m2s, _RegFile_reg_22__0__m2s, n4192, 
        _RegFile_reg_22__10__m2s, _RegFile_reg_22__11__m2s, 
        _RegFile_reg_22__12__m2s, _RegFile_reg_22__13__m2s, 
        _RegFile_reg_22__14__m2s, _RegFile_reg_22__15__m2s, 
        _RegFile_reg_22__16__m2s, _RegFile_reg_22__17__m2s, 
        _RegFile_reg_22__18__m2s, _RegFile_reg_22__19__m2s, 
        _RegFile_reg_22__1__m2s, n4191, _RegFile_reg_22__20__m2s, 
        _RegFile_reg_22__21__m2s, _RegFile_reg_22__22__m2s, 
        _RegFile_reg_22__23__m2s, _RegFile_reg_22__24__m2s, 
        _RegFile_reg_22__25__m2s, _RegFile_reg_22__26__m2s, 
        _RegFile_reg_22__27__m2s, _RegFile_reg_22__28__m2s, 
        _RegFile_reg_22__29__m2s, _RegFile_reg_22__2__m2s, n4190, 
        _RegFile_reg_22__30__m2s, _RegFile_reg_22__31__m2s, 
        _RegFile_reg_22__3__m2s, n4189, _RegFile_reg_22__4__m2s, n4188, 
        _RegFile_reg_22__5__m2s, n4187, _RegFile_reg_22__6__m2s, n4186, 
        _RegFile_reg_22__7__m2s, n4185, _RegFile_reg_22__8__m2s, 
        _RegFile_reg_22__9__m2s, _RegFile_reg_23__0__m2s, n4184, 
        _RegFile_reg_23__10__m2s, _RegFile_reg_23__11__m2s, 
        _RegFile_reg_23__12__m2s, _RegFile_reg_23__13__m2s, 
        _RegFile_reg_23__14__m2s, _RegFile_reg_23__15__m2s, 
        _RegFile_reg_23__16__m2s, _RegFile_reg_23__17__m2s, 
        _RegFile_reg_23__18__m2s, _RegFile_reg_23__19__m2s, 
        _RegFile_reg_23__1__m2s, n4183, _RegFile_reg_23__20__m2s, 
        _RegFile_reg_23__21__m2s, _RegFile_reg_23__22__m2s, 
        _RegFile_reg_23__23__m2s, _RegFile_reg_23__24__m2s, 
        _RegFile_reg_23__25__m2s, _RegFile_reg_23__26__m2s, 
        _RegFile_reg_23__27__m2s, _RegFile_reg_23__28__m2s, 
        _RegFile_reg_23__29__m2s, _RegFile_reg_23__2__m2s, n4182, 
        _RegFile_reg_23__30__m2s, _RegFile_reg_23__31__m2s, 
        _RegFile_reg_23__3__m2s, n4181, _RegFile_reg_23__4__m2s, n4180, 
        _RegFile_reg_23__5__m2s, n4179, _RegFile_reg_23__6__m2s, n4178, 
        _RegFile_reg_23__7__m2s, n4177, _RegFile_reg_23__8__m2s, 
        _RegFile_reg_23__9__m2s, _RegFile_reg_24__0__m2s, n4176, 
        _RegFile_reg_24__10__m2s, _RegFile_reg_24__11__m2s, 
        _RegFile_reg_24__12__m2s, _RegFile_reg_24__13__m2s, 
        _RegFile_reg_24__14__m2s, _RegFile_reg_24__15__m2s, 
        _RegFile_reg_24__16__m2s, _RegFile_reg_24__17__m2s, 
        _RegFile_reg_24__18__m2s, _RegFile_reg_24__19__m2s, 
        _RegFile_reg_24__1__m2s, n4175, _RegFile_reg_24__20__m2s, 
        _RegFile_reg_24__21__m2s, _RegFile_reg_24__22__m2s, 
        _RegFile_reg_24__23__m2s, _RegFile_reg_24__24__m2s, 
        _RegFile_reg_24__25__m2s, _RegFile_reg_24__26__m2s, 
        _RegFile_reg_24__27__m2s, _RegFile_reg_24__28__m2s, 
        _RegFile_reg_24__29__m2s, _RegFile_reg_24__2__m2s, n4174, 
        _RegFile_reg_24__30__m2s, _RegFile_reg_24__31__m2s, 
        _RegFile_reg_24__3__m2s, n4173, _RegFile_reg_24__4__m2s, n4172, 
        _RegFile_reg_24__5__m2s, n4171, _RegFile_reg_24__6__m2s, n4170, 
        _RegFile_reg_24__7__m2s, n4169, _RegFile_reg_24__8__m2s, 
        _RegFile_reg_24__9__m2s, _RegFile_reg_25__0__m2s, n4168, 
        _RegFile_reg_25__10__m2s, _RegFile_reg_25__11__m2s, 
        _RegFile_reg_25__12__m2s, _RegFile_reg_25__13__m2s, 
        _RegFile_reg_25__14__m2s, _RegFile_reg_25__15__m2s, 
        _RegFile_reg_25__16__m2s, _RegFile_reg_25__17__m2s, 
        _RegFile_reg_25__18__m2s, _RegFile_reg_25__19__m2s, 
        _RegFile_reg_25__1__m2s, n4167, _RegFile_reg_25__20__m2s, 
        _RegFile_reg_25__21__m2s, _RegFile_reg_25__22__m2s, 
        _RegFile_reg_25__23__m2s, _RegFile_reg_25__24__m2s, 
        _RegFile_reg_25__25__m2s, _RegFile_reg_25__26__m2s, 
        _RegFile_reg_25__27__m2s, _RegFile_reg_25__28__m2s, 
        _RegFile_reg_25__29__m2s, _RegFile_reg_25__2__m2s, n4166, 
        _RegFile_reg_25__30__m2s, _RegFile_reg_25__31__m2s, 
        _RegFile_reg_25__3__m2s, n4165, _RegFile_reg_25__4__m2s, n4164, 
        _RegFile_reg_25__5__m2s, n4163, _RegFile_reg_25__6__m2s, n4162, 
        _RegFile_reg_25__7__m2s, n4161, _RegFile_reg_25__8__m2s, 
        _RegFile_reg_25__9__m2s, _RegFile_reg_26__0__m2s, n4160, 
        _RegFile_reg_26__10__m2s, _RegFile_reg_26__11__m2s, 
        _RegFile_reg_26__12__m2s, _RegFile_reg_26__13__m2s, 
        _RegFile_reg_26__14__m2s, _RegFile_reg_26__15__m2s, 
        _RegFile_reg_26__16__m2s, _RegFile_reg_26__17__m2s, 
        _RegFile_reg_26__18__m2s, _RegFile_reg_26__19__m2s, 
        _RegFile_reg_26__1__m2s, n4159, _RegFile_reg_26__20__m2s, 
        _RegFile_reg_26__21__m2s, _RegFile_reg_26__22__m2s, 
        _RegFile_reg_26__23__m2s, _RegFile_reg_26__24__m2s, 
        _RegFile_reg_26__25__m2s, _RegFile_reg_26__26__m2s, 
        _RegFile_reg_26__27__m2s, _RegFile_reg_26__28__m2s, 
        _RegFile_reg_26__29__m2s, _RegFile_reg_26__2__m2s, n4158, 
        _RegFile_reg_26__30__m2s, _RegFile_reg_26__31__m2s, 
        _RegFile_reg_26__3__m2s, n4157, _RegFile_reg_26__4__m2s, n4156, 
        _RegFile_reg_26__5__m2s, n4155, _RegFile_reg_26__6__m2s, n4154, 
        _RegFile_reg_26__7__m2s, n4153, _RegFile_reg_26__8__m2s, 
        _RegFile_reg_26__9__m2s, _RegFile_reg_27__0__m2s, n4152, 
        _RegFile_reg_27__10__m2s, _RegFile_reg_27__11__m2s, 
        _RegFile_reg_27__12__m2s, _RegFile_reg_27__13__m2s, 
        _RegFile_reg_27__14__m2s, _RegFile_reg_27__15__m2s, 
        _RegFile_reg_27__16__m2s, _RegFile_reg_27__17__m2s, 
        _RegFile_reg_27__18__m2s, _RegFile_reg_27__19__m2s, 
        _RegFile_reg_27__1__m2s, n4151, _RegFile_reg_27__20__m2s, 
        _RegFile_reg_27__21__m2s, _RegFile_reg_27__22__m2s, 
        _RegFile_reg_27__23__m2s, _RegFile_reg_27__24__m2s, 
        _RegFile_reg_27__25__m2s, _RegFile_reg_27__26__m2s, 
        _RegFile_reg_27__27__m2s, _RegFile_reg_27__28__m2s, 
        _RegFile_reg_27__29__m2s, _RegFile_reg_27__2__m2s, n4150, 
        _RegFile_reg_27__30__m2s, _RegFile_reg_27__31__m2s, 
        _RegFile_reg_27__3__m2s, n4149, _RegFile_reg_27__4__m2s, n4148, 
        _RegFile_reg_27__5__m2s, n4147, _RegFile_reg_27__6__m2s, n4146, 
        _RegFile_reg_27__7__m2s, n4145, _RegFile_reg_27__8__m2s, 
        _RegFile_reg_27__9__m2s, _RegFile_reg_28__0__m2s, n4144, 
        _RegFile_reg_28__10__m2s, _RegFile_reg_28__11__m2s, 
        _RegFile_reg_28__12__m2s, _RegFile_reg_28__13__m2s, 
        _RegFile_reg_28__14__m2s, _RegFile_reg_28__15__m2s, 
        _RegFile_reg_28__16__m2s, _RegFile_reg_28__17__m2s, 
        _RegFile_reg_28__18__m2s, _RegFile_reg_28__19__m2s, 
        _RegFile_reg_28__1__m2s, n4143, _RegFile_reg_28__20__m2s, 
        _RegFile_reg_28__21__m2s, _RegFile_reg_28__22__m2s, 
        _RegFile_reg_28__23__m2s, _RegFile_reg_28__24__m2s, 
        _RegFile_reg_28__25__m2s, _RegFile_reg_28__26__m2s, 
        _RegFile_reg_28__27__m2s, _RegFile_reg_28__28__m2s, 
        _RegFile_reg_28__29__m2s, _RegFile_reg_28__2__m2s, n4142, 
        _RegFile_reg_28__30__m2s, _RegFile_reg_28__31__m2s, 
        _RegFile_reg_28__3__m2s, n4141, _RegFile_reg_28__4__m2s, n4140, 
        _RegFile_reg_28__5__m2s, n4139, _RegFile_reg_28__6__m2s, n4138, 
        _RegFile_reg_28__7__m2s, n4137, _RegFile_reg_28__8__m2s, 
        _RegFile_reg_28__9__m2s, _RegFile_reg_29__0__m2s, n4136, 
        _RegFile_reg_29__10__m2s, _RegFile_reg_29__11__m2s, 
        _RegFile_reg_29__12__m2s, _RegFile_reg_29__13__m2s, 
        _RegFile_reg_29__14__m2s, _RegFile_reg_29__15__m2s, 
        _RegFile_reg_29__16__m2s, _RegFile_reg_29__17__m2s, 
        _RegFile_reg_29__18__m2s, _RegFile_reg_29__19__m2s, 
        _RegFile_reg_29__1__m2s, n4135, _RegFile_reg_29__20__m2s, 
        _RegFile_reg_29__21__m2s, _RegFile_reg_29__22__m2s, 
        _RegFile_reg_29__23__m2s, _RegFile_reg_29__24__m2s, 
        _RegFile_reg_29__25__m2s, _RegFile_reg_29__26__m2s, 
        _RegFile_reg_29__27__m2s, _RegFile_reg_29__28__m2s, 
        _RegFile_reg_29__29__m2s, _RegFile_reg_29__2__m2s, n4134, 
        _RegFile_reg_29__30__m2s, _RegFile_reg_29__31__m2s, 
        _RegFile_reg_29__3__m2s, n4133, _RegFile_reg_29__4__m2s, n4132, 
        _RegFile_reg_29__5__m2s, n4131, _RegFile_reg_29__6__m2s, n4130, 
        _RegFile_reg_29__7__m2s, n4129, _RegFile_reg_29__8__m2s, 
        _RegFile_reg_29__9__m2s, _RegFile_reg_2__0__m2s, n4352, 
        _RegFile_reg_2__10__m2s, _RegFile_reg_2__11__m2s, 
        _RegFile_reg_2__12__m2s, _RegFile_reg_2__13__m2s, 
        _RegFile_reg_2__14__m2s, _RegFile_reg_2__15__m2s, 
        _RegFile_reg_2__16__m2s, _RegFile_reg_2__17__m2s, 
        _RegFile_reg_2__18__m2s, _RegFile_reg_2__19__m2s, 
        _RegFile_reg_2__1__m2s, n4351, _RegFile_reg_2__20__m2s, 
        _RegFile_reg_2__21__m2s, _RegFile_reg_2__22__m2s, 
        _RegFile_reg_2__23__m2s, _RegFile_reg_2__24__m2s, 
        _RegFile_reg_2__25__m2s, _RegFile_reg_2__26__m2s, 
        _RegFile_reg_2__27__m2s, _RegFile_reg_2__28__m2s, 
        _RegFile_reg_2__29__m2s, _RegFile_reg_2__2__m2s, n4350, 
        _RegFile_reg_2__30__m2s, _RegFile_reg_2__31__m2s, 
        _RegFile_reg_2__3__m2s, n4349, _RegFile_reg_2__4__m2s, n4348, 
        _RegFile_reg_2__5__m2s, n4347, _RegFile_reg_2__6__m2s, n4346, 
        _RegFile_reg_2__7__m2s, n4345, _RegFile_reg_2__8__m2s, 
        _RegFile_reg_2__9__m2s, _RegFile_reg_30__0__m2s, n4128, 
        _RegFile_reg_30__10__m2s, _RegFile_reg_30__11__m2s, 
        _RegFile_reg_30__12__m2s, _RegFile_reg_30__13__m2s, 
        _RegFile_reg_30__14__m2s, _RegFile_reg_30__15__m2s, 
        _RegFile_reg_30__16__m2s, _RegFile_reg_30__17__m2s, 
        _RegFile_reg_30__18__m2s, _RegFile_reg_30__19__m2s, 
        _RegFile_reg_30__1__m2s, n4127, _RegFile_reg_30__20__m2s, 
        _RegFile_reg_30__21__m2s, _RegFile_reg_30__22__m2s, 
        _RegFile_reg_30__23__m2s, _RegFile_reg_30__24__m2s, 
        _RegFile_reg_30__25__m2s, _RegFile_reg_30__26__m2s, 
        _RegFile_reg_30__27__m2s, _RegFile_reg_30__28__m2s, 
        _RegFile_reg_30__29__m2s, _RegFile_reg_30__2__m2s, n4126, 
        _RegFile_reg_30__30__m2s, _RegFile_reg_30__31__m2s, 
        _RegFile_reg_30__3__m2s, n4125, _RegFile_reg_30__4__m2s, n4124, 
        _RegFile_reg_30__5__m2s, n4123, _RegFile_reg_30__6__m2s, n4122, 
        _RegFile_reg_30__7__m2s, n4121, _RegFile_reg_30__8__m2s, 
        _RegFile_reg_30__9__m2s, _RegFile_reg_31__0__m2s, n4120, 
        _RegFile_reg_31__10__m2s, _RegFile_reg_31__11__m2s, 
        _RegFile_reg_31__12__m2s, _RegFile_reg_31__13__m2s, 
        _RegFile_reg_31__14__m2s, _RegFile_reg_31__15__m2s, 
        _RegFile_reg_31__16__m2s, _RegFile_reg_31__17__m2s, 
        _RegFile_reg_31__18__m2s, _RegFile_reg_31__19__m2s, 
        _RegFile_reg_31__1__m2s, n4119, _RegFile_reg_31__20__m2s, 
        _RegFile_reg_31__21__m2s, _RegFile_reg_31__22__m2s, 
        _RegFile_reg_31__23__m2s, _RegFile_reg_31__24__m2s, 
        _RegFile_reg_31__25__m2s, _RegFile_reg_31__26__m2s, 
        _RegFile_reg_31__27__m2s, _RegFile_reg_31__28__m2s, 
        _RegFile_reg_31__29__m2s, _RegFile_reg_31__2__m2s, n4118, 
        _RegFile_reg_31__30__m2s, _RegFile_reg_31__31__m2s, 
        _RegFile_reg_31__3__m2s, n4117, _RegFile_reg_31__4__m2s, n4116, 
        _RegFile_reg_31__5__m2s, n4115, _RegFile_reg_31__6__m2s, n4114, 
        _RegFile_reg_31__7__m2s, n4113, _RegFile_reg_31__8__m2s, 
        _RegFile_reg_31__9__m2s, _RegFile_reg_3__0__m2s, n4344, 
        _RegFile_reg_3__10__m2s, _RegFile_reg_3__11__m2s, 
        _RegFile_reg_3__12__m2s, _RegFile_reg_3__13__m2s, 
        _RegFile_reg_3__14__m2s, _RegFile_reg_3__15__m2s, 
        _RegFile_reg_3__16__m2s, _RegFile_reg_3__17__m2s, 
        _RegFile_reg_3__18__m2s, _RegFile_reg_3__19__m2s, 
        _RegFile_reg_3__1__m2s, n4343, _RegFile_reg_3__20__m2s, 
        _RegFile_reg_3__21__m2s, _RegFile_reg_3__22__m2s, 
        _RegFile_reg_3__23__m2s, _RegFile_reg_3__24__m2s, 
        _RegFile_reg_3__25__m2s, _RegFile_reg_3__26__m2s, 
        _RegFile_reg_3__27__m2s, _RegFile_reg_3__28__m2s, 
        _RegFile_reg_3__29__m2s, _RegFile_reg_3__2__m2s, n4342, 
        _RegFile_reg_3__30__m2s, _RegFile_reg_3__31__m2s, 
        _RegFile_reg_3__3__m2s, n4341, _RegFile_reg_3__4__m2s, n4340, 
        _RegFile_reg_3__5__m2s, n4339, _RegFile_reg_3__6__m2s, n4338, 
        _RegFile_reg_3__7__m2s, n4337, _RegFile_reg_3__8__m2s, 
        _RegFile_reg_3__9__m2s, _RegFile_reg_4__0__m2s, n4336, 
        _RegFile_reg_4__10__m2s, _RegFile_reg_4__11__m2s, 
        _RegFile_reg_4__12__m2s, _RegFile_reg_4__13__m2s, 
        _RegFile_reg_4__14__m2s, _RegFile_reg_4__15__m2s, 
        _RegFile_reg_4__16__m2s, _RegFile_reg_4__17__m2s, 
        _RegFile_reg_4__18__m2s, _RegFile_reg_4__19__m2s, 
        _RegFile_reg_4__1__m2s, n4335, _RegFile_reg_4__20__m2s, 
        _RegFile_reg_4__21__m2s, _RegFile_reg_4__22__m2s, 
        _RegFile_reg_4__23__m2s, _RegFile_reg_4__24__m2s, 
        _RegFile_reg_4__25__m2s, _RegFile_reg_4__26__m2s, 
        _RegFile_reg_4__27__m2s, _RegFile_reg_4__28__m2s, 
        _RegFile_reg_4__29__m2s, _RegFile_reg_4__2__m2s, n4334, 
        _RegFile_reg_4__30__m2s, _RegFile_reg_4__31__m2s, 
        _RegFile_reg_4__3__m2s, n4333, _RegFile_reg_4__4__m2s, n4332, 
        _RegFile_reg_4__5__m2s, n4331, _RegFile_reg_4__6__m2s, n4330, 
        _RegFile_reg_4__7__m2s, n4329, _RegFile_reg_4__8__m2s, 
        _RegFile_reg_4__9__m2s, _RegFile_reg_5__0__m2s, n4328, 
        _RegFile_reg_5__10__m2s, _RegFile_reg_5__11__m2s, 
        _RegFile_reg_5__12__m2s, _RegFile_reg_5__13__m2s, 
        _RegFile_reg_5__14__m2s, _RegFile_reg_5__15__m2s, 
        _RegFile_reg_5__16__m2s, _RegFile_reg_5__17__m2s, 
        _RegFile_reg_5__18__m2s, _RegFile_reg_5__19__m2s, 
        _RegFile_reg_5__1__m2s, n4327, _RegFile_reg_5__20__m2s, 
        _RegFile_reg_5__21__m2s, _RegFile_reg_5__22__m2s, 
        _RegFile_reg_5__23__m2s, _RegFile_reg_5__24__m2s, 
        _RegFile_reg_5__25__m2s, _RegFile_reg_5__26__m2s, 
        _RegFile_reg_5__27__m2s, _RegFile_reg_5__28__m2s, 
        _RegFile_reg_5__29__m2s, _RegFile_reg_5__2__m2s, n4326, 
        _RegFile_reg_5__30__m2s, _RegFile_reg_5__31__m2s, 
        _RegFile_reg_5__3__m2s, n4325, _RegFile_reg_5__4__m2s, n4324, 
        _RegFile_reg_5__5__m2s, n4323, _RegFile_reg_5__6__m2s, n4322, 
        _RegFile_reg_5__7__m2s, n4321, _RegFile_reg_5__8__m2s, 
        _RegFile_reg_5__9__m2s, _RegFile_reg_6__0__m2s, n4320, 
        _RegFile_reg_6__10__m2s, _RegFile_reg_6__11__m2s, 
        _RegFile_reg_6__12__m2s, _RegFile_reg_6__13__m2s, 
        _RegFile_reg_6__14__m2s, _RegFile_reg_6__15__m2s, 
        _RegFile_reg_6__16__m2s, _RegFile_reg_6__17__m2s, 
        _RegFile_reg_6__18__m2s, _RegFile_reg_6__19__m2s, 
        _RegFile_reg_6__1__m2s, n4319, _RegFile_reg_6__20__m2s, 
        _RegFile_reg_6__21__m2s, _RegFile_reg_6__22__m2s, 
        _RegFile_reg_6__23__m2s, _RegFile_reg_6__24__m2s, 
        _RegFile_reg_6__25__m2s, _RegFile_reg_6__26__m2s, 
        _RegFile_reg_6__27__m2s, _RegFile_reg_6__28__m2s, 
        _RegFile_reg_6__29__m2s, _RegFile_reg_6__2__m2s, n4318, 
        _RegFile_reg_6__30__m2s, _RegFile_reg_6__31__m2s, 
        _RegFile_reg_6__3__m2s, n4317, _RegFile_reg_6__4__m2s, n4316, 
        _RegFile_reg_6__5__m2s, n4315, _RegFile_reg_6__6__m2s, n4314, 
        _RegFile_reg_6__7__m2s, n4313, _RegFile_reg_6__8__m2s, 
        _RegFile_reg_6__9__m2s, _RegFile_reg_7__0__m2s, n4312, 
        _RegFile_reg_7__10__m2s, _RegFile_reg_7__11__m2s, 
        _RegFile_reg_7__12__m2s, _RegFile_reg_7__13__m2s, 
        _RegFile_reg_7__14__m2s, _RegFile_reg_7__15__m2s, 
        _RegFile_reg_7__16__m2s, _RegFile_reg_7__17__m2s, 
        _RegFile_reg_7__18__m2s, _RegFile_reg_7__19__m2s, 
        _RegFile_reg_7__1__m2s, n4311, _RegFile_reg_7__20__m2s, 
        _RegFile_reg_7__21__m2s, _RegFile_reg_7__22__m2s, 
        _RegFile_reg_7__23__m2s, _RegFile_reg_7__24__m2s, 
        _RegFile_reg_7__25__m2s, _RegFile_reg_7__26__m2s, 
        _RegFile_reg_7__27__m2s, _RegFile_reg_7__28__m2s, 
        _RegFile_reg_7__29__m2s, _RegFile_reg_7__2__m2s, n4310, 
        _RegFile_reg_7__30__m2s, _RegFile_reg_7__31__m2s, 
        _RegFile_reg_7__3__m2s, n4309, _RegFile_reg_7__4__m2s, n4308, 
        _RegFile_reg_7__5__m2s, n4307, _RegFile_reg_7__6__m2s, n4306, 
        _RegFile_reg_7__7__m2s, n4305, _RegFile_reg_7__8__m2s, 
        _RegFile_reg_7__9__m2s, _RegFile_reg_8__0__m2s, n4304, 
        _RegFile_reg_8__10__m2s, _RegFile_reg_8__11__m2s, 
        _RegFile_reg_8__12__m2s, _RegFile_reg_8__13__m2s, 
        _RegFile_reg_8__14__m2s, _RegFile_reg_8__15__m2s, 
        _RegFile_reg_8__16__m2s, _RegFile_reg_8__17__m2s, 
        _RegFile_reg_8__18__m2s, _RegFile_reg_8__19__m2s, 
        _RegFile_reg_8__1__m2s, n4303, _RegFile_reg_8__20__m2s, 
        _RegFile_reg_8__21__m2s, _RegFile_reg_8__22__m2s, 
        _RegFile_reg_8__23__m2s, _RegFile_reg_8__24__m2s, 
        _RegFile_reg_8__25__m2s, _RegFile_reg_8__26__m2s, 
        _RegFile_reg_8__27__m2s, _RegFile_reg_8__28__m2s, 
        _RegFile_reg_8__29__m2s, _RegFile_reg_8__2__m2s, n4302, 
        _RegFile_reg_8__30__m2s, _RegFile_reg_8__31__m2s, 
        _RegFile_reg_8__3__m2s, n4301, _RegFile_reg_8__4__m2s, n4300, 
        _RegFile_reg_8__5__m2s, n4299, _RegFile_reg_8__6__m2s, n4298, 
        _RegFile_reg_8__7__m2s, n4297, _RegFile_reg_8__8__m2s, 
        _RegFile_reg_8__9__m2s, _RegFile_reg_9__0__m2s, n4296, 
        _RegFile_reg_9__10__m2s, _RegFile_reg_9__11__m2s, 
        _RegFile_reg_9__12__m2s, _RegFile_reg_9__13__m2s, 
        _RegFile_reg_9__14__m2s, _RegFile_reg_9__15__m2s, 
        _RegFile_reg_9__16__m2s, _RegFile_reg_9__17__m2s, 
        _RegFile_reg_9__18__m2s, _RegFile_reg_9__19__m2s, 
        _RegFile_reg_9__1__m2s, n4295, _RegFile_reg_9__20__m2s, 
        _RegFile_reg_9__21__m2s, _RegFile_reg_9__22__m2s, 
        _RegFile_reg_9__23__m2s, _RegFile_reg_9__24__m2s, 
        _RegFile_reg_9__25__m2s, _RegFile_reg_9__26__m2s, 
        _RegFile_reg_9__27__m2s, _RegFile_reg_9__28__m2s, 
        _RegFile_reg_9__29__m2s, _RegFile_reg_9__2__m2s, n4294, 
        _RegFile_reg_9__30__m2s, _RegFile_reg_9__31__m2s, 
        _RegFile_reg_9__3__m2s, n4293, _RegFile_reg_9__4__m2s, n4292, 
        _RegFile_reg_9__5__m2s, n4291, _RegFile_reg_9__6__m2s, n4290, 
        _RegFile_reg_9__7__m2s, n4289, _RegFile_reg_9__8__m2s, 
        _RegFile_reg_9__9__m2s, N5350, N5349, N5348, N5347, N5346, N5345, 
        N5344, N5343, N5342, N5341, N5340, N5339, N5338, N5337, N5336, N5335, 
        N5334, N5333, N5332, N5331, N5330, N5329, N5328, N5327, N5326, N5325, 
        N5324, N5323, N5322, N5321, N5320, N5319, N5418, N5417, N5416, N5415, 
        N5414, N5413, N5412, N5411, N5410, N5409, N5408, N5407, N5406, N5405, 
        N5404, N5403, N5402, N5401, N5400, N5399, N5398, N5397, N5396, N5395, 
        N5394, N5393, N5392, N5391, N5390, N5389, N5388, N5387, N6017, N6016, 
        N6015, N6014, N6013, N6012, N6011, N6010, N6009, N6008, N6007, N6006, 
        N6005, N6004, N6003, N6002, N6001, N6000, N5999, N5998, N5997, N5996, 
        N5995, N5994, N5993, N5992, N5991, N5990, N5989, N5988, N5987, N5986, 
        branch_address_reg_0__m2s, n4112, branch_address_reg_10__m2s, n4104, 
        n4103, branch_address_reg_11__m2s, n4102, branch_address_reg_12__m2s, 
        n4101, branch_address_reg_13__m2s, n4100, branch_address_reg_14__m2s, 
        n4099, branch_address_reg_15__m2s, n4098, branch_address_reg_16__m2s, 
        n4097, branch_address_reg_17__m2s, n4096, branch_address_reg_18__m2s, 
        n4095, branch_address_reg_19__m2s, n4094, branch_address_reg_1__m2s, 
        n4111, branch_address_reg_20__m2s, n4093, branch_address_reg_21__m2s, 
        n4092, branch_address_reg_22__m2s, n4091, branch_address_reg_23__m2s, 
        n4090, branch_address_reg_24__m2s, n4089, branch_address_reg_25__m2s, 
        n4088, branch_address_reg_26__m2s, n4087, branch_address_reg_27__m2s, 
        n4086, branch_address_reg_28__m2s, n4085, branch_address_reg_29__m2s, 
        n4084, branch_address_reg_2__m2s, n4110, branch_address_reg_30__m2s, 
        n4083, branch_address_reg_31__m2s, branch_address_reg_3__m2s, n4109, 
        branch_address_reg_4__m2s, n4108, branch_address_reg_5__m2s, n4107, 
        branch_address_reg_6__m2s, n4106, branch_address_reg_7__m2s, 
        branch_address_reg_8__m2s, n4105, branch_address_reg_9__m2s, 
        branch_sig_reg__m2s, counter_reg_0__m2s, counter_reg_1__m2s, 
        current_IR_reg_0__m2s, n4082, current_IR_reg_10__m2s, 
        current_IR_reg_11__m2s, n4076, current_IR_reg_12__m2s, n4075, 
        current_IR_reg_13__m2s, n4074, current_IR_reg_14__m2s, n4073, 
        current_IR_reg_15__m2s, n4072, current_IR_reg_16__m2s, 
        current_IR_reg_17__m2s, n4071, current_IR_reg_18__m2s, n4070, 
        current_IR_reg_19__m2s, current_IR_reg_1__m2s, n4081, 
        current_IR_reg_20__m2s, n4069, current_IR_reg_21__m2s, 
        current_IR_reg_22__m2s, current_IR_reg_23__m2s, current_IR_reg_24__m2s, 
        n4068, current_IR_reg_25__m2s, n4067, current_IR_reg_26__m2s, n4066, 
        current_IR_reg_27__m2s, n4065, current_IR_reg_28__m2s, n4064, 
        current_IR_reg_29__m2s, current_IR_reg_2__m2s, n4080, 
        current_IR_reg_30__m2s, current_IR_reg_31__m2s, current_IR_reg_3__m2s, 
        current_IR_reg_4__m2s, n4079, current_IR_reg_5__m2s, n4078, 
        current_IR_reg_6__m2s, current_IR_reg_7__m2s, n4077, 
        current_IR_reg_8__m2s, current_IR_reg_9__m2s, delay_slot_reg__m2s, 
        intr_slot_reg__m2s, mem_read_reg__m2s, mem_to_reg_reg__m2s, 
        mem_write_reg__m2s, opcode_of_MEM_reg_0__m2s, opcode_of_MEM_0, 
        opcode_of_MEM_reg_1__m2s, n4063, opcode_of_MEM_reg_2__m2s, 
        opcode_of_MEM_reg_3__m2s, opcode_of_MEM_reg_4__m2s, n4062, 
        opcode_of_MEM_reg_5__m2s, n4061, opcode_of_WB_reg_0__m2s, n4060, 
        opcode_of_WB_reg_1__m2s, n4059, opcode_of_WB_reg_2__m2s, n4058, 
        opcode_of_WB_reg_3__m2s, n4057, opcode_of_WB_reg_4__m2s, n4056, 
        opcode_of_WB_reg_5__m2s, n4055, rd_addr_reg_0__m2s, rd_addr_reg_1__m2s, 
        rd_addr_reg_2__m2s, rd_addr_reg_3__m2s, n4054, rd_addr_reg_4__m2s, 
        reg_dst_of_MEM_reg_0__m2s, n4053, reg_dst_of_MEM_reg_1__m2s, n4052, 
        reg_dst_of_MEM_reg_2__m2s, reg_dst_of_MEM_reg_3__m2s, 
        reg_dst_of_MEM_reg_4__m2s, reg_dst_reg__m2s, reg_out_A_reg_0__m2s, 
        n4051, reg_out_A_reg_10__m2s, n4042, n4041, reg_out_A_reg_11__m2s, 
        n4040, reg_out_A_reg_12__m2s, n4039, reg_out_A_reg_13__m2s, n4038, 
        reg_out_A_reg_14__m2s, n4037, reg_out_A_reg_15__m2s, n4036, 
        reg_out_A_reg_16__m2s, n4035, reg_out_A_reg_17__m2s, n4034, 
        reg_out_A_reg_18__m2s, n4033, reg_out_A_reg_19__m2s, n4032, 
        reg_out_A_reg_1__m2s, n4050, reg_out_A_reg_20__m2s, n4031, 
        reg_out_A_reg_21__m2s, n4030, reg_out_A_reg_22__m2s, n4029, 
        reg_out_A_reg_23__m2s, n4028, reg_out_A_reg_24__m2s, n4027, 
        reg_out_A_reg_25__m2s, n4026, reg_out_A_reg_26__m2s, n4025, 
        reg_out_A_reg_27__m2s, n4024, reg_out_A_reg_28__m2s, n4023, 
        reg_out_A_reg_29__m2s, n4022, reg_out_A_reg_2__m2s, n4049, 
        reg_out_A_reg_30__m2s, n4021, reg_out_A_reg_31__m2s, n4020, 
        reg_out_A_reg_3__m2s, n4048, reg_out_A_reg_4__m2s, n4047, 
        reg_out_A_reg_5__m2s, n4046, reg_out_A_reg_6__m2s, n4045, 
        reg_out_A_reg_7__m2s, n4044, reg_out_A_reg_8__m2s, n4043, 
        reg_out_A_reg_9__m2s, reg_out_B_reg_0__m2s, n4393, 
        reg_out_B_reg_10__m2s, n4389, n4413, reg_out_B_reg_11__m2s, n4395, 
        reg_out_B_reg_12__m2s, n4433, reg_out_B_reg_13__m2s, n4425, 
        reg_out_B_reg_14__m2s, n4421, reg_out_B_reg_15__m2s, n4403, 
        reg_out_B_reg_16__m2s, n4411, reg_out_B_reg_17__m2s, n4443, 
        reg_out_B_reg_18__m2s, n4427, reg_out_B_reg_19__m2s, n4423, 
        reg_out_B_reg_1__m2s, n4445, reg_out_B_reg_20__m2s, n4391, 
        reg_out_B_reg_21__m2s, n4437, reg_out_B_reg_22__m2s, n4447, 
        reg_out_B_reg_23__m2s, n4415, reg_out_B_reg_24__m2s, n4417, 
        reg_out_B_reg_25__m2s, n4435, reg_out_B_reg_26__m2s, n4407, 
        reg_out_B_reg_27__m2s, n4431, reg_out_B_reg_28__m2s, n4401, 
        reg_out_B_reg_29__m2s, n4397, reg_out_B_reg_2__m2s, n4439, 
        reg_out_B_reg_30__m2s, n4449, reg_out_B_reg_31__m2s, n4451, 
        reg_out_B_reg_3__m2s, n4441, reg_out_B_reg_4__m2s, n4399, 
        reg_out_B_reg_5__m2s, n4419, reg_out_B_reg_6__m2s, n4405, 
        reg_out_B_reg_7__m2s, n4429, reg_out_B_reg_8__m2s, n4409, 
        reg_out_B_reg_9__m2s, reg_write_reg__m2s, rt_addr_reg_0__m2s, 
        rt_addr_reg_1__m2s, rt_addr_reg_2__m2s, rt_addr_reg_3__m2s, 
        rt_addr_reg_4__m2s, slot_num_reg_0__m2s, n4019, slot_num_reg_1__m2s, 
        stall_reg__m2s;
    assign test_so = stall;
    DLX_sync_MUX_OP_32_5_32_2_test_1 C440 ( .D0_31(_RegFile_0__0), .D0_30(
        _RegFile_0__1), .D0_29(_RegFile_0__2), .D0_28(_RegFile_0__3), .D0_27(
        _RegFile_0__4), .D0_26(_RegFile_0__5), .D0_25(_RegFile_0__6), .D0_24(
        _RegFile_0__7), .D0_23(_RegFile_0__8), .D0_22(_RegFile_0__9), .D0_21(
        _RegFile_0__10), .D0_20(_RegFile_0__11), .D0_19(_RegFile_0__12), 
        .D0_18(_RegFile_0__13), .D0_17(_RegFile_0__14), .D0_16(_RegFile_0__15), 
        .D0_15(_RegFile_0__16), .D0_14(_RegFile_0__17), .D0_13(_RegFile_0__18), 
        .D0_12(_RegFile_0__19), .D0_11(_RegFile_0__20), .D0_10(_RegFile_0__21), 
        .D0_9(_RegFile_0__22), .D0_8(_RegFile_0__23), .D0_7(_RegFile_0__24), 
        .D0_6(_RegFile_0__25), .D0_5(_RegFile_0__26), .D0_4(_RegFile_0__27), 
        .D0_3(_RegFile_0__28), .D0_2(_RegFile_0__29), .D0_1(_RegFile_0__30), 
        .D0_0(_RegFile_0__31), .D1_31(_RegFile_1__0), .D1_30(_RegFile_1__1), 
        .D1_29(_RegFile_1__2), .D1_28(_RegFile_1__3), .D1_27(_RegFile_1__4), 
        .D1_26(_RegFile_1__5), .D1_25(_RegFile_1__6), .D1_24(_RegFile_1__7), 
        .D1_23(_RegFile_1__8), .D1_22(_RegFile_1__9), .D1_21(_RegFile_1__10), 
        .D1_20(_RegFile_1__11), .D1_19(_RegFile_1__12), .D1_18(_RegFile_1__13), 
        .D1_17(_RegFile_1__14), .D1_16(_RegFile_1__15), .D1_15(_RegFile_1__16), 
        .D1_14(_RegFile_1__17), .D1_13(_RegFile_1__18), .D1_12(_RegFile_1__19), 
        .D1_11(_RegFile_1__20), .D1_10(_RegFile_1__21), .D1_9(_RegFile_1__22), 
        .D1_8(_RegFile_1__23), .D1_7(_RegFile_1__24), .D1_6(_RegFile_1__25), 
        .D1_5(_RegFile_1__26), .D1_4(_RegFile_1__27), .D1_3(_RegFile_1__28), 
        .D1_2(_RegFile_1__29), .D1_1(_RegFile_1__30), .D1_0(_RegFile_1__31), 
        .D2_31(_RegFile_2__0), .D2_30(_RegFile_2__1), .D2_29(_RegFile_2__2), 
        .D2_28(_RegFile_2__3), .D2_27(_RegFile_2__4), .D2_26(_RegFile_2__5), 
        .D2_25(_RegFile_2__6), .D2_24(_RegFile_2__7), .D2_23(_RegFile_2__8), 
        .D2_22(_RegFile_2__9), .D2_21(_RegFile_2__10), .D2_20(_RegFile_2__11), 
        .D2_19(_RegFile_2__12), .D2_18(_RegFile_2__13), .D2_17(_RegFile_2__14), 
        .D2_16(_RegFile_2__15), .D2_15(_RegFile_2__16), .D2_14(_RegFile_2__17), 
        .D2_13(_RegFile_2__18), .D2_12(_RegFile_2__19), .D2_11(_RegFile_2__20), 
        .D2_10(_RegFile_2__21), .D2_9(_RegFile_2__22), .D2_8(_RegFile_2__23), 
        .D2_7(_RegFile_2__24), .D2_6(_RegFile_2__25), .D2_5(_RegFile_2__26), 
        .D2_4(_RegFile_2__27), .D2_3(_RegFile_2__28), .D2_2(_RegFile_2__29), 
        .D2_1(_RegFile_2__30), .D2_0(_RegFile_2__31), .D3_31(_RegFile_3__0), 
        .D3_30(_RegFile_3__1), .D3_29(_RegFile_3__2), .D3_28(_RegFile_3__3), 
        .D3_27(_RegFile_3__4), .D3_26(_RegFile_3__5), .D3_25(_RegFile_3__6), 
        .D3_24(_RegFile_3__7), .D3_23(_RegFile_3__8), .D3_22(_RegFile_3__9), 
        .D3_21(_RegFile_3__10), .D3_20(_RegFile_3__11), .D3_19(_RegFile_3__12), 
        .D3_18(_RegFile_3__13), .D3_17(_RegFile_3__14), .D3_16(_RegFile_3__15), 
        .D3_15(_RegFile_3__16), .D3_14(_RegFile_3__17), .D3_13(_RegFile_3__18), 
        .D3_12(_RegFile_3__19), .D3_11(_RegFile_3__20), .D3_10(_RegFile_3__21), 
        .D3_9(_RegFile_3__22), .D3_8(_RegFile_3__23), .D3_7(_RegFile_3__24), 
        .D3_6(_RegFile_3__25), .D3_5(_RegFile_3__26), .D3_4(_RegFile_3__27), 
        .D3_3(_RegFile_3__28), .D3_2(_RegFile_3__29), .D3_1(_RegFile_3__30), 
        .D3_0(_RegFile_3__31), .D4_31(_RegFile_4__0), .D4_30(_RegFile_4__1), 
        .D4_29(_RegFile_4__2), .D4_28(_RegFile_4__3), .D4_27(_RegFile_4__4), 
        .D4_26(_RegFile_4__5), .D4_25(_RegFile_4__6), .D4_24(_RegFile_4__7), 
        .D4_23(_RegFile_4__8), .D4_22(_RegFile_4__9), .D4_21(_RegFile_4__10), 
        .D4_20(_RegFile_4__11), .D4_19(_RegFile_4__12), .D4_18(_RegFile_4__13), 
        .D4_17(_RegFile_4__14), .D4_16(_RegFile_4__15), .D4_15(_RegFile_4__16), 
        .D4_14(_RegFile_4__17), .D4_13(_RegFile_4__18), .D4_12(_RegFile_4__19), 
        .D4_11(_RegFile_4__20), .D4_10(_RegFile_4__21), .D4_9(_RegFile_4__22), 
        .D4_8(_RegFile_4__23), .D4_7(_RegFile_4__24), .D4_6(_RegFile_4__25), 
        .D4_5(_RegFile_4__26), .D4_4(_RegFile_4__27), .D4_3(_RegFile_4__28), 
        .D4_2(_RegFile_4__29), .D4_1(_RegFile_4__30), .D4_0(_RegFile_4__31), 
        .D5_31(_RegFile_5__0), .D5_30(_RegFile_5__1), .D5_29(_RegFile_5__2), 
        .D5_28(_RegFile_5__3), .D5_27(_RegFile_5__4), .D5_26(_RegFile_5__5), 
        .D5_25(_RegFile_5__6), .D5_24(_RegFile_5__7), .D5_23(_RegFile_5__8), 
        .D5_22(_RegFile_5__9), .D5_21(_RegFile_5__10), .D5_20(_RegFile_5__11), 
        .D5_19(_RegFile_5__12), .D5_18(_RegFile_5__13), .D5_17(_RegFile_5__14), 
        .D5_16(_RegFile_5__15), .D5_15(_RegFile_5__16), .D5_14(_RegFile_5__17), 
        .D5_13(_RegFile_5__18), .D5_12(_RegFile_5__19), .D5_11(_RegFile_5__20), 
        .D5_10(_RegFile_5__21), .D5_9(_RegFile_5__22), .D5_8(_RegFile_5__23), 
        .D5_7(_RegFile_5__24), .D5_6(_RegFile_5__25), .D5_5(_RegFile_5__26), 
        .D5_4(_RegFile_5__27), .D5_3(_RegFile_5__28), .D5_2(_RegFile_5__29), 
        .D5_1(_RegFile_5__30), .D5_0(_RegFile_5__31), .D6_31(_RegFile_6__0), 
        .D6_30(_RegFile_6__1), .D6_29(_RegFile_6__2), .D6_28(_RegFile_6__3), 
        .D6_27(_RegFile_6__4), .D6_26(_RegFile_6__5), .D6_25(_RegFile_6__6), 
        .D6_24(_RegFile_6__7), .D6_23(_RegFile_6__8), .D6_22(_RegFile_6__9), 
        .D6_21(_RegFile_6__10), .D6_20(_RegFile_6__11), .D6_19(_RegFile_6__12), 
        .D6_18(_RegFile_6__13), .D6_17(_RegFile_6__14), .D6_16(_RegFile_6__15), 
        .D6_15(_RegFile_6__16), .D6_14(_RegFile_6__17), .D6_13(_RegFile_6__18), 
        .D6_12(_RegFile_6__19), .D6_11(_RegFile_6__20), .D6_10(_RegFile_6__21), 
        .D6_9(_RegFile_6__22), .D6_8(_RegFile_6__23), .D6_7(_RegFile_6__24), 
        .D6_6(_RegFile_6__25), .D6_5(_RegFile_6__26), .D6_4(_RegFile_6__27), 
        .D6_3(_RegFile_6__28), .D6_2(_RegFile_6__29), .D6_1(_RegFile_6__30), 
        .D6_0(_RegFile_6__31), .D7_31(_RegFile_7__0), .D7_30(_RegFile_7__1), 
        .D7_29(_RegFile_7__2), .D7_28(_RegFile_7__3), .D7_27(_RegFile_7__4), 
        .D7_26(_RegFile_7__5), .D7_25(_RegFile_7__6), .D7_24(_RegFile_7__7), 
        .D7_23(_RegFile_7__8), .D7_22(_RegFile_7__9), .D7_21(_RegFile_7__10), 
        .D7_20(_RegFile_7__11), .D7_19(_RegFile_7__12), .D7_18(_RegFile_7__13), 
        .D7_17(_RegFile_7__14), .D7_16(_RegFile_7__15), .D7_15(_RegFile_7__16), 
        .D7_14(_RegFile_7__17), .D7_13(_RegFile_7__18), .D7_12(_RegFile_7__19), 
        .D7_11(_RegFile_7__20), .D7_10(_RegFile_7__21), .D7_9(_RegFile_7__22), 
        .D7_8(_RegFile_7__23), .D7_7(_RegFile_7__24), .D7_6(_RegFile_7__25), 
        .D7_5(_RegFile_7__26), .D7_4(_RegFile_7__27), .D7_3(_RegFile_7__28), 
        .D7_2(_RegFile_7__29), .D7_1(_RegFile_7__30), .D7_0(_RegFile_7__31), 
        .D8_31(_RegFile_8__0), .D8_30(_RegFile_8__1), .D8_29(_RegFile_8__2), 
        .D8_28(_RegFile_8__3), .D8_27(_RegFile_8__4), .D8_26(_RegFile_8__5), 
        .D8_25(_RegFile_8__6), .D8_24(_RegFile_8__7), .D8_23(_RegFile_8__8), 
        .D8_22(_RegFile_8__9), .D8_21(_RegFile_8__10), .D8_20(_RegFile_8__11), 
        .D8_19(_RegFile_8__12), .D8_18(_RegFile_8__13), .D8_17(_RegFile_8__14), 
        .D8_16(_RegFile_8__15), .D8_15(_RegFile_8__16), .D8_14(_RegFile_8__17), 
        .D8_13(_RegFile_8__18), .D8_12(_RegFile_8__19), .D8_11(_RegFile_8__20), 
        .D8_10(_RegFile_8__21), .D8_9(_RegFile_8__22), .D8_8(_RegFile_8__23), 
        .D8_7(_RegFile_8__24), .D8_6(_RegFile_8__25), .D8_5(_RegFile_8__26), 
        .D8_4(_RegFile_8__27), .D8_3(_RegFile_8__28), .D8_2(_RegFile_8__29), 
        .D8_1(_RegFile_8__30), .D8_0(_RegFile_8__31), .D9_31(_RegFile_9__0), 
        .D9_30(_RegFile_9__1), .D9_29(_RegFile_9__2), .D9_28(_RegFile_9__3), 
        .D9_27(_RegFile_9__4), .D9_26(_RegFile_9__5), .D9_25(_RegFile_9__6), 
        .D9_24(_RegFile_9__7), .D9_23(_RegFile_9__8), .D9_22(_RegFile_9__9), 
        .D9_21(_RegFile_9__10), .D9_20(_RegFile_9__11), .D9_19(_RegFile_9__12), 
        .D9_18(_RegFile_9__13), .D9_17(_RegFile_9__14), .D9_16(_RegFile_9__15), 
        .D9_15(_RegFile_9__16), .D9_14(_RegFile_9__17), .D9_13(_RegFile_9__18), 
        .D9_12(_RegFile_9__19), .D9_11(_RegFile_9__20), .D9_10(_RegFile_9__21), 
        .D9_9(_RegFile_9__22), .D9_8(_RegFile_9__23), .D9_7(_RegFile_9__24), 
        .D9_6(_RegFile_9__25), .D9_5(_RegFile_9__26), .D9_4(_RegFile_9__27), 
        .D9_3(_RegFile_9__28), .D9_2(_RegFile_9__29), .D9_1(_RegFile_9__30), 
        .D9_0(_RegFile_9__31), .D10_31(_RegFile_10__0), .D10_30(_RegFile_10__1
        ), .D10_29(_RegFile_10__2), .D10_28(_RegFile_10__3), .D10_27(
        _RegFile_10__4), .D10_26(_RegFile_10__5), .D10_25(_RegFile_10__6), 
        .D10_24(_RegFile_10__7), .D10_23(_RegFile_10__8), .D10_22(
        _RegFile_10__9), .D10_21(_RegFile_10__10), .D10_20(_RegFile_10__11), 
        .D10_19(_RegFile_10__12), .D10_18(_RegFile_10__13), .D10_17(
        _RegFile_10__14), .D10_16(_RegFile_10__15), .D10_15(_RegFile_10__16), 
        .D10_14(_RegFile_10__17), .D10_13(_RegFile_10__18), .D10_12(
        _RegFile_10__19), .D10_11(_RegFile_10__20), .D10_10(_RegFile_10__21), 
        .D10_9(_RegFile_10__22), .D10_8(_RegFile_10__23), .D10_7(
        _RegFile_10__24), .D10_6(_RegFile_10__25), .D10_5(_RegFile_10__26), 
        .D10_4(_RegFile_10__27), .D10_3(_RegFile_10__28), .D10_2(
        _RegFile_10__29), .D10_1(_RegFile_10__30), .D10_0(_RegFile_10__31), 
        .D11_31(_RegFile_11__0), .D11_30(_RegFile_11__1), .D11_29(
        _RegFile_11__2), .D11_28(_RegFile_11__3), .D11_27(_RegFile_11__4), 
        .D11_26(_RegFile_11__5), .D11_25(_RegFile_11__6), .D11_24(
        _RegFile_11__7), .D11_23(_RegFile_11__8), .D11_22(_RegFile_11__9), 
        .D11_21(_RegFile_11__10), .D11_20(_RegFile_11__11), .D11_19(
        _RegFile_11__12), .D11_18(_RegFile_11__13), .D11_17(_RegFile_11__14), 
        .D11_16(_RegFile_11__15), .D11_15(_RegFile_11__16), .D11_14(
        _RegFile_11__17), .D11_13(_RegFile_11__18), .D11_12(_RegFile_11__19), 
        .D11_11(_RegFile_11__20), .D11_10(_RegFile_11__21), .D11_9(
        _RegFile_11__22), .D11_8(_RegFile_11__23), .D11_7(_RegFile_11__24), 
        .D11_6(_RegFile_11__25), .D11_5(_RegFile_11__26), .D11_4(
        _RegFile_11__27), .D11_3(_RegFile_11__28), .D11_2(_RegFile_11__29), 
        .D11_1(_RegFile_11__30), .D11_0(_RegFile_11__31), .D12_31(
        _RegFile_12__0), .D12_30(_RegFile_12__1), .D12_29(_RegFile_12__2), 
        .D12_28(_RegFile_12__3), .D12_27(_RegFile_12__4), .D12_26(
        _RegFile_12__5), .D12_25(_RegFile_12__6), .D12_24(_RegFile_12__7), 
        .D12_23(_RegFile_12__8), .D12_22(_RegFile_12__9), .D12_21(
        _RegFile_12__10), .D12_20(_RegFile_12__11), .D12_19(_RegFile_12__12), 
        .D12_18(_RegFile_12__13), .D12_17(_RegFile_12__14), .D12_16(
        _RegFile_12__15), .D12_15(_RegFile_12__16), .D12_14(_RegFile_12__17), 
        .D12_13(_RegFile_12__18), .D12_12(_RegFile_12__19), .D12_11(
        _RegFile_12__20), .D12_10(_RegFile_12__21), .D12_9(_RegFile_12__22), 
        .D12_8(_RegFile_12__23), .D12_7(_RegFile_12__24), .D12_6(
        _RegFile_12__25), .D12_5(_RegFile_12__26), .D12_4(_RegFile_12__27), 
        .D12_3(_RegFile_12__28), .D12_2(_RegFile_12__29), .D12_1(
        _RegFile_12__30), .D12_0(_RegFile_12__31), .D13_31(_RegFile_13__0), 
        .D13_30(_RegFile_13__1), .D13_29(_RegFile_13__2), .D13_28(
        _RegFile_13__3), .D13_27(_RegFile_13__4), .D13_26(_RegFile_13__5), 
        .D13_25(_RegFile_13__6), .D13_24(_RegFile_13__7), .D13_23(
        _RegFile_13__8), .D13_22(_RegFile_13__9), .D13_21(_RegFile_13__10), 
        .D13_20(_RegFile_13__11), .D13_19(_RegFile_13__12), .D13_18(
        _RegFile_13__13), .D13_17(_RegFile_13__14), .D13_16(_RegFile_13__15), 
        .D13_15(_RegFile_13__16), .D13_14(_RegFile_13__17), .D13_13(
        _RegFile_13__18), .D13_12(_RegFile_13__19), .D13_11(_RegFile_13__20), 
        .D13_10(_RegFile_13__21), .D13_9(_RegFile_13__22), .D13_8(
        _RegFile_13__23), .D13_7(_RegFile_13__24), .D13_6(_RegFile_13__25), 
        .D13_5(_RegFile_13__26), .D13_4(_RegFile_13__27), .D13_3(
        _RegFile_13__28), .D13_2(_RegFile_13__29), .D13_1(_RegFile_13__30), 
        .D13_0(_RegFile_13__31), .D14_31(_RegFile_14__0), .D14_30(
        _RegFile_14__1), .D14_29(_RegFile_14__2), .D14_28(_RegFile_14__3), 
        .D14_27(_RegFile_14__4), .D14_26(_RegFile_14__5), .D14_25(
        _RegFile_14__6), .D14_24(_RegFile_14__7), .D14_23(_RegFile_14__8), 
        .D14_22(_RegFile_14__9), .D14_21(_RegFile_14__10), .D14_20(
        _RegFile_14__11), .D14_19(_RegFile_14__12), .D14_18(_RegFile_14__13), 
        .D14_17(_RegFile_14__14), .D14_16(_RegFile_14__15), .D14_15(
        _RegFile_14__16), .D14_14(_RegFile_14__17), .D14_13(_RegFile_14__18), 
        .D14_12(_RegFile_14__19), .D14_11(_RegFile_14__20), .D14_10(
        _RegFile_14__21), .D14_9(_RegFile_14__22), .D14_8(_RegFile_14__23), 
        .D14_7(_RegFile_14__24), .D14_6(_RegFile_14__25), .D14_5(
        _RegFile_14__26), .D14_4(_RegFile_14__27), .D14_3(_RegFile_14__28), 
        .D14_2(_RegFile_14__29), .D14_1(_RegFile_14__30), .D14_0(
        _RegFile_14__31), .D15_31(_RegFile_15__0), .D15_30(_RegFile_15__1), 
        .D15_29(_RegFile_15__2), .D15_28(_RegFile_15__3), .D15_27(
        _RegFile_15__4), .D15_26(_RegFile_15__5), .D15_25(_RegFile_15__6), 
        .D15_24(_RegFile_15__7), .D15_23(_RegFile_15__8), .D15_22(
        _RegFile_15__9), .D15_21(_RegFile_15__10), .D15_20(_RegFile_15__11), 
        .D15_19(_RegFile_15__12), .D15_18(_RegFile_15__13), .D15_17(
        _RegFile_15__14), .D15_16(_RegFile_15__15), .D15_15(_RegFile_15__16), 
        .D15_14(_RegFile_15__17), .D15_13(_RegFile_15__18), .D15_12(
        _RegFile_15__19), .D15_11(_RegFile_15__20), .D15_10(_RegFile_15__21), 
        .D15_9(_RegFile_15__22), .D15_8(_RegFile_15__23), .D15_7(
        _RegFile_15__24), .D15_6(_RegFile_15__25), .D15_5(_RegFile_15__26), 
        .D15_4(_RegFile_15__27), .D15_3(_RegFile_15__28), .D15_2(
        _RegFile_15__29), .D15_1(_RegFile_15__30), .D15_0(_RegFile_15__31), 
        .D16_31(_RegFile_16__0), .D16_30(_RegFile_16__1), .D16_29(
        _RegFile_16__2), .D16_28(_RegFile_16__3), .D16_27(_RegFile_16__4), 
        .D16_26(_RegFile_16__5), .D16_25(_RegFile_16__6), .D16_24(
        _RegFile_16__7), .D16_23(_RegFile_16__8), .D16_22(_RegFile_16__9), 
        .D16_21(_RegFile_16__10), .D16_20(_RegFile_16__11), .D16_19(
        _RegFile_16__12), .D16_18(_RegFile_16__13), .D16_17(_RegFile_16__14), 
        .D16_16(_RegFile_16__15), .D16_15(_RegFile_16__16), .D16_14(
        _RegFile_16__17), .D16_13(_RegFile_16__18), .D16_12(_RegFile_16__19), 
        .D16_11(_RegFile_16__20), .D16_10(_RegFile_16__21), .D16_9(
        _RegFile_16__22), .D16_8(_RegFile_16__23), .D16_7(_RegFile_16__24), 
        .D16_6(_RegFile_16__25), .D16_5(_RegFile_16__26), .D16_4(
        _RegFile_16__27), .D16_3(_RegFile_16__28), .D16_2(_RegFile_16__29), 
        .D16_1(_RegFile_16__30), .D16_0(_RegFile_16__31), .D17_31(
        _RegFile_17__0), .D17_30(_RegFile_17__1), .D17_29(_RegFile_17__2), 
        .D17_28(_RegFile_17__3), .D17_27(_RegFile_17__4), .D17_26(
        _RegFile_17__5), .D17_25(_RegFile_17__6), .D17_24(_RegFile_17__7), 
        .D17_23(_RegFile_17__8), .D17_22(_RegFile_17__9), .D17_21(
        _RegFile_17__10), .D17_20(_RegFile_17__11), .D17_19(_RegFile_17__12), 
        .D17_18(_RegFile_17__13), .D17_17(_RegFile_17__14), .D17_16(
        _RegFile_17__15), .D17_15(_RegFile_17__16), .D17_14(_RegFile_17__17), 
        .D17_13(_RegFile_17__18), .D17_12(_RegFile_17__19), .D17_11(
        _RegFile_17__20), .D17_10(_RegFile_17__21), .D17_9(_RegFile_17__22), 
        .D17_8(_RegFile_17__23), .D17_7(_RegFile_17__24), .D17_6(
        _RegFile_17__25), .D17_5(_RegFile_17__26), .D17_4(_RegFile_17__27), 
        .D17_3(_RegFile_17__28), .D17_2(_RegFile_17__29), .D17_1(
        _RegFile_17__30), .D17_0(_RegFile_17__31), .D18_31(_RegFile_18__0), 
        .D18_30(_RegFile_18__1), .D18_29(_RegFile_18__2), .D18_28(
        _RegFile_18__3), .D18_27(_RegFile_18__4), .D18_26(_RegFile_18__5), 
        .D18_25(_RegFile_18__6), .D18_24(_RegFile_18__7), .D18_23(
        _RegFile_18__8), .D18_22(_RegFile_18__9), .D18_21(_RegFile_18__10), 
        .D18_20(_RegFile_18__11), .D18_19(_RegFile_18__12), .D18_18(
        _RegFile_18__13), .D18_17(_RegFile_18__14), .D18_16(_RegFile_18__15), 
        .D18_15(_RegFile_18__16), .D18_14(_RegFile_18__17), .D18_13(
        _RegFile_18__18), .D18_12(_RegFile_18__19), .D18_11(_RegFile_18__20), 
        .D18_10(_RegFile_18__21), .D18_9(_RegFile_18__22), .D18_8(
        _RegFile_18__23), .D18_7(_RegFile_18__24), .D18_6(_RegFile_18__25), 
        .D18_5(_RegFile_18__26), .D18_4(_RegFile_18__27), .D18_3(
        _RegFile_18__28), .D18_2(_RegFile_18__29), .D18_1(_RegFile_18__30), 
        .D18_0(_RegFile_18__31), .D19_31(_RegFile_19__0), .D19_30(
        _RegFile_19__1), .D19_29(_RegFile_19__2), .D19_28(_RegFile_19__3), 
        .D19_27(_RegFile_19__4), .D19_26(_RegFile_19__5), .D19_25(
        _RegFile_19__6), .D19_24(_RegFile_19__7), .D19_23(_RegFile_19__8), 
        .D19_22(_RegFile_19__9), .D19_21(_RegFile_19__10), .D19_20(
        _RegFile_19__11), .D19_19(_RegFile_19__12), .D19_18(_RegFile_19__13), 
        .D19_17(_RegFile_19__14), .D19_16(_RegFile_19__15), .D19_15(
        _RegFile_19__16), .D19_14(_RegFile_19__17), .D19_13(_RegFile_19__18), 
        .D19_12(_RegFile_19__19), .D19_11(_RegFile_19__20), .D19_10(
        _RegFile_19__21), .D19_9(_RegFile_19__22), .D19_8(_RegFile_19__23), 
        .D19_7(_RegFile_19__24), .D19_6(_RegFile_19__25), .D19_5(
        _RegFile_19__26), .D19_4(_RegFile_19__27), .D19_3(_RegFile_19__28), 
        .D19_2(_RegFile_19__29), .D19_1(_RegFile_19__30), .D19_0(
        _RegFile_19__31), .D20_31(_RegFile_20__0), .D20_30(_RegFile_20__1), 
        .D20_29(_RegFile_20__2), .D20_28(_RegFile_20__3), .D20_27(
        _RegFile_20__4), .D20_26(_RegFile_20__5), .D20_25(_RegFile_20__6), 
        .D20_24(_RegFile_20__7), .D20_23(_RegFile_20__8), .D20_22(
        _RegFile_20__9), .D20_21(_RegFile_20__10), .D20_20(_RegFile_20__11), 
        .D20_19(_RegFile_20__12), .D20_18(_RegFile_20__13), .D20_17(
        _RegFile_20__14), .D20_16(_RegFile_20__15), .D20_15(_RegFile_20__16), 
        .D20_14(_RegFile_20__17), .D20_13(_RegFile_20__18), .D20_12(
        _RegFile_20__19), .D20_11(_RegFile_20__20), .D20_10(_RegFile_20__21), 
        .D20_9(_RegFile_20__22), .D20_8(_RegFile_20__23), .D20_7(
        _RegFile_20__24), .D20_6(_RegFile_20__25), .D20_5(_RegFile_20__26), 
        .D20_4(_RegFile_20__27), .D20_3(_RegFile_20__28), .D20_2(
        _RegFile_20__29), .D20_1(_RegFile_20__30), .D20_0(_RegFile_20__31), 
        .D21_31(_RegFile_21__0), .D21_30(_RegFile_21__1), .D21_29(
        _RegFile_21__2), .D21_28(_RegFile_21__3), .D21_27(_RegFile_21__4), 
        .D21_26(_RegFile_21__5), .D21_25(_RegFile_21__6), .D21_24(
        _RegFile_21__7), .D21_23(_RegFile_21__8), .D21_22(_RegFile_21__9), 
        .D21_21(_RegFile_21__10), .D21_20(_RegFile_21__11), .D21_19(
        _RegFile_21__12), .D21_18(_RegFile_21__13), .D21_17(_RegFile_21__14), 
        .D21_16(_RegFile_21__15), .D21_15(_RegFile_21__16), .D21_14(
        _RegFile_21__17), .D21_13(_RegFile_21__18), .D21_12(_RegFile_21__19), 
        .D21_11(_RegFile_21__20), .D21_10(_RegFile_21__21), .D21_9(
        _RegFile_21__22), .D21_8(_RegFile_21__23), .D21_7(_RegFile_21__24), 
        .D21_6(_RegFile_21__25), .D21_5(_RegFile_21__26), .D21_4(
        _RegFile_21__27), .D21_3(_RegFile_21__28), .D21_2(_RegFile_21__29), 
        .D21_1(_RegFile_21__30), .D21_0(_RegFile_21__31), .D22_31(
        _RegFile_22__0), .D22_30(_RegFile_22__1), .D22_29(_RegFile_22__2), 
        .D22_28(_RegFile_22__3), .D22_27(_RegFile_22__4), .D22_26(
        _RegFile_22__5), .D22_25(_RegFile_22__6), .D22_24(_RegFile_22__7), 
        .D22_23(_RegFile_22__8), .D22_22(_RegFile_22__9), .D22_21(
        _RegFile_22__10), .D22_20(_RegFile_22__11), .D22_19(_RegFile_22__12), 
        .D22_18(_RegFile_22__13), .D22_17(_RegFile_22__14), .D22_16(
        _RegFile_22__15), .D22_15(_RegFile_22__16), .D22_14(_RegFile_22__17), 
        .D22_13(_RegFile_22__18), .D22_12(_RegFile_22__19), .D22_11(
        _RegFile_22__20), .D22_10(_RegFile_22__21), .D22_9(_RegFile_22__22), 
        .D22_8(_RegFile_22__23), .D22_7(_RegFile_22__24), .D22_6(
        _RegFile_22__25), .D22_5(_RegFile_22__26), .D22_4(_RegFile_22__27), 
        .D22_3(_RegFile_22__28), .D22_2(_RegFile_22__29), .D22_1(
        _RegFile_22__30), .D22_0(_RegFile_22__31), .D23_31(_RegFile_23__0), 
        .D23_30(_RegFile_23__1), .D23_29(_RegFile_23__2), .D23_28(
        _RegFile_23__3), .D23_27(_RegFile_23__4), .D23_26(_RegFile_23__5), 
        .D23_25(_RegFile_23__6), .D23_24(_RegFile_23__7), .D23_23(
        _RegFile_23__8), .D23_22(_RegFile_23__9), .D23_21(_RegFile_23__10), 
        .D23_20(_RegFile_23__11), .D23_19(_RegFile_23__12), .D23_18(
        _RegFile_23__13), .D23_17(_RegFile_23__14), .D23_16(_RegFile_23__15), 
        .D23_15(_RegFile_23__16), .D23_14(_RegFile_23__17), .D23_13(
        _RegFile_23__18), .D23_12(_RegFile_23__19), .D23_11(_RegFile_23__20), 
        .D23_10(_RegFile_23__21), .D23_9(_RegFile_23__22), .D23_8(
        _RegFile_23__23), .D23_7(_RegFile_23__24), .D23_6(_RegFile_23__25), 
        .D23_5(_RegFile_23__26), .D23_4(_RegFile_23__27), .D23_3(
        _RegFile_23__28), .D23_2(_RegFile_23__29), .D23_1(_RegFile_23__30), 
        .D23_0(_RegFile_23__31), .D24_31(_RegFile_24__0), .D24_30(
        _RegFile_24__1), .D24_29(_RegFile_24__2), .D24_28(_RegFile_24__3), 
        .D24_27(_RegFile_24__4), .D24_26(_RegFile_24__5), .D24_25(
        _RegFile_24__6), .D24_24(_RegFile_24__7), .D24_23(_RegFile_24__8), 
        .D24_22(_RegFile_24__9), .D24_21(_RegFile_24__10), .D24_20(
        _RegFile_24__11), .D24_19(_RegFile_24__12), .D24_18(_RegFile_24__13), 
        .D24_17(_RegFile_24__14), .D24_16(_RegFile_24__15), .D24_15(
        _RegFile_24__16), .D24_14(_RegFile_24__17), .D24_13(_RegFile_24__18), 
        .D24_12(_RegFile_24__19), .D24_11(_RegFile_24__20), .D24_10(
        _RegFile_24__21), .D24_9(_RegFile_24__22), .D24_8(_RegFile_24__23), 
        .D24_7(_RegFile_24__24), .D24_6(_RegFile_24__25), .D24_5(
        _RegFile_24__26), .D24_4(_RegFile_24__27), .D24_3(_RegFile_24__28), 
        .D24_2(_RegFile_24__29), .D24_1(_RegFile_24__30), .D24_0(
        _RegFile_24__31), .D25_31(_RegFile_25__0), .D25_30(_RegFile_25__1), 
        .D25_29(_RegFile_25__2), .D25_28(_RegFile_25__3), .D25_27(
        _RegFile_25__4), .D25_26(_RegFile_25__5), .D25_25(_RegFile_25__6), 
        .D25_24(_RegFile_25__7), .D25_23(_RegFile_25__8), .D25_22(
        _RegFile_25__9), .D25_21(_RegFile_25__10), .D25_20(_RegFile_25__11), 
        .D25_19(_RegFile_25__12), .D25_18(_RegFile_25__13), .D25_17(
        _RegFile_25__14), .D25_16(_RegFile_25__15), .D25_15(_RegFile_25__16), 
        .D25_14(_RegFile_25__17), .D25_13(_RegFile_25__18), .D25_12(
        _RegFile_25__19), .D25_11(_RegFile_25__20), .D25_10(_RegFile_25__21), 
        .D25_9(_RegFile_25__22), .D25_8(_RegFile_25__23), .D25_7(
        _RegFile_25__24), .D25_6(_RegFile_25__25), .D25_5(_RegFile_25__26), 
        .D25_4(_RegFile_25__27), .D25_3(_RegFile_25__28), .D25_2(
        _RegFile_25__29), .D25_1(_RegFile_25__30), .D25_0(_RegFile_25__31), 
        .D26_31(_RegFile_26__0), .D26_30(_RegFile_26__1), .D26_29(
        _RegFile_26__2), .D26_28(_RegFile_26__3), .D26_27(_RegFile_26__4), 
        .D26_26(_RegFile_26__5), .D26_25(_RegFile_26__6), .D26_24(
        _RegFile_26__7), .D26_23(_RegFile_26__8), .D26_22(_RegFile_26__9), 
        .D26_21(_RegFile_26__10), .D26_20(_RegFile_26__11), .D26_19(
        _RegFile_26__12), .D26_18(_RegFile_26__13), .D26_17(_RegFile_26__14), 
        .D26_16(_RegFile_26__15), .D26_15(_RegFile_26__16), .D26_14(
        _RegFile_26__17), .D26_13(_RegFile_26__18), .D26_12(_RegFile_26__19), 
        .D26_11(_RegFile_26__20), .D26_10(_RegFile_26__21), .D26_9(
        _RegFile_26__22), .D26_8(_RegFile_26__23), .D26_7(_RegFile_26__24), 
        .D26_6(_RegFile_26__25), .D26_5(_RegFile_26__26), .D26_4(
        _RegFile_26__27), .D26_3(_RegFile_26__28), .D26_2(_RegFile_26__29), 
        .D26_1(_RegFile_26__30), .D26_0(_RegFile_26__31), .D27_31(
        _RegFile_27__0), .D27_30(_RegFile_27__1), .D27_29(_RegFile_27__2), 
        .D27_28(_RegFile_27__3), .D27_27(_RegFile_27__4), .D27_26(
        _RegFile_27__5), .D27_25(_RegFile_27__6), .D27_24(_RegFile_27__7), 
        .D27_23(_RegFile_27__8), .D27_22(_RegFile_27__9), .D27_21(
        _RegFile_27__10), .D27_20(_RegFile_27__11), .D27_19(_RegFile_27__12), 
        .D27_18(_RegFile_27__13), .D27_17(_RegFile_27__14), .D27_16(
        _RegFile_27__15), .D27_15(_RegFile_27__16), .D27_14(_RegFile_27__17), 
        .D27_13(_RegFile_27__18), .D27_12(_RegFile_27__19), .D27_11(
        _RegFile_27__20), .D27_10(_RegFile_27__21), .D27_9(_RegFile_27__22), 
        .D27_8(_RegFile_27__23), .D27_7(_RegFile_27__24), .D27_6(
        _RegFile_27__25), .D27_5(_RegFile_27__26), .D27_4(_RegFile_27__27), 
        .D27_3(_RegFile_27__28), .D27_2(_RegFile_27__29), .D27_1(
        _RegFile_27__30), .D27_0(_RegFile_27__31), .D28_31(_RegFile_28__0), 
        .D28_30(_RegFile_28__1), .D28_29(_RegFile_28__2), .D28_28(
        _RegFile_28__3), .D28_27(_RegFile_28__4), .D28_26(_RegFile_28__5), 
        .D28_25(_RegFile_28__6), .D28_24(_RegFile_28__7), .D28_23(
        _RegFile_28__8), .D28_22(_RegFile_28__9), .D28_21(_RegFile_28__10), 
        .D28_20(_RegFile_28__11), .D28_19(_RegFile_28__12), .D28_18(
        _RegFile_28__13), .D28_17(_RegFile_28__14), .D28_16(_RegFile_28__15), 
        .D28_15(_RegFile_28__16), .D28_14(_RegFile_28__17), .D28_13(
        _RegFile_28__18), .D28_12(_RegFile_28__19), .D28_11(_RegFile_28__20), 
        .D28_10(_RegFile_28__21), .D28_9(_RegFile_28__22), .D28_8(
        _RegFile_28__23), .D28_7(_RegFile_28__24), .D28_6(_RegFile_28__25), 
        .D28_5(_RegFile_28__26), .D28_4(_RegFile_28__27), .D28_3(
        _RegFile_28__28), .D28_2(_RegFile_28__29), .D28_1(_RegFile_28__30), 
        .D28_0(_RegFile_28__31), .D29_31(_RegFile_29__0), .D29_30(
        _RegFile_29__1), .D29_29(_RegFile_29__2), .D29_28(_RegFile_29__3), 
        .D29_27(_RegFile_29__4), .D29_26(_RegFile_29__5), .D29_25(
        _RegFile_29__6), .D29_24(_RegFile_29__7), .D29_23(_RegFile_29__8), 
        .D29_22(_RegFile_29__9), .D29_21(_RegFile_29__10), .D29_20(
        _RegFile_29__11), .D29_19(_RegFile_29__12), .D29_18(_RegFile_29__13), 
        .D29_17(_RegFile_29__14), .D29_16(_RegFile_29__15), .D29_15(
        _RegFile_29__16), .D29_14(_RegFile_29__17), .D29_13(_RegFile_29__18), 
        .D29_12(_RegFile_29__19), .D29_11(_RegFile_29__20), .D29_10(
        _RegFile_29__21), .D29_9(_RegFile_29__22), .D29_8(_RegFile_29__23), 
        .D29_7(_RegFile_29__24), .D29_6(_RegFile_29__25), .D29_5(
        _RegFile_29__26), .D29_4(_RegFile_29__27), .D29_3(_RegFile_29__28), 
        .D29_2(_RegFile_29__29), .D29_1(_RegFile_29__30), .D29_0(
        _RegFile_29__31), .D30_31(_RegFile_30__0), .D30_30(_RegFile_30__1), 
        .D30_29(_RegFile_30__2), .D30_28(_RegFile_30__3), .D30_27(
        _RegFile_30__4), .D30_26(_RegFile_30__5), .D30_25(_RegFile_30__6), 
        .D30_24(_RegFile_30__7), .D30_23(_RegFile_30__8), .D30_22(
        _RegFile_30__9), .D30_21(_RegFile_30__10), .D30_20(_RegFile_30__11), 
        .D30_19(_RegFile_30__12), .D30_18(_RegFile_30__13), .D30_17(
        _RegFile_30__14), .D30_16(_RegFile_30__15), .D30_15(_RegFile_30__16), 
        .D30_14(_RegFile_30__17), .D30_13(_RegFile_30__18), .D30_12(
        _RegFile_30__19), .D30_11(_RegFile_30__20), .D30_10(_RegFile_30__21), 
        .D30_9(_RegFile_30__22), .D30_8(_RegFile_30__23), .D30_7(
        _RegFile_30__24), .D30_6(_RegFile_30__25), .D30_5(_RegFile_30__26), 
        .D30_4(_RegFile_30__27), .D30_3(_RegFile_30__28), .D30_2(
        _RegFile_30__29), .D30_1(_RegFile_30__30), .D30_0(_RegFile_30__31), 
        .D31_31(_RegFile_31__0), .D31_30(_RegFile_31__1), .D31_29(
        _RegFile_31__2), .D31_28(_RegFile_31__3), .D31_27(_RegFile_31__4), 
        .D31_26(_RegFile_31__5), .D31_25(_RegFile_31__6), .D31_24(
        _RegFile_31__7), .D31_23(_RegFile_31__8), .D31_22(_RegFile_31__9), 
        .D31_21(_RegFile_31__10), .D31_20(_RegFile_31__11), .D31_19(
        _RegFile_31__12), .D31_18(_RegFile_31__13), .D31_17(_RegFile_31__14), 
        .D31_16(_RegFile_31__15), .D31_15(_RegFile_31__16), .D31_14(
        _RegFile_31__17), .D31_13(_RegFile_31__18), .D31_12(_RegFile_31__19), 
        .D31_11(_RegFile_31__20), .D31_10(_RegFile_31__21), .D31_9(
        _RegFile_31__22), .D31_8(_RegFile_31__23), .D31_7(_RegFile_31__24), 
        .D31_6(_RegFile_31__25), .D31_5(_RegFile_31__26), .D31_4(
        _RegFile_31__27), .D31_3(_RegFile_31__28), .D31_2(_RegFile_31__29), 
        .D31_1(_RegFile_31__30), .D31_0(_RegFile_31__31), .S0(n804), .S1(n896), 
        .S2(n694), .S3(n332), .S4(n331), .Z_31(N468), .Z_30(N467), .Z_29(N466), 
        .Z_28(N465), .Z_27(N464), .Z_26(N463), .Z_25(N462), .Z_24(N461), 
        .Z_23(N460), .Z_22(N459), .Z_21(N458), .Z_20(N457), .Z_19(N456), 
        .Z_18(N455), .Z_17(N454), .Z_16(N453), .Z_15(N452), .Z_14(N451), 
        .Z_13(N450), .Z_12(N449), .Z_11(N448), .Z_10(N447), .Z_9(N446), .Z_8(
        N445), .Z_7(N444), .Z_6(N443), .Z_5(N442), .Z_4(N441), .Z_3(N440), 
        .Z_2(N439), .Z_1(N438), .Z_0(N437) );
    DLX_sync_MUX_OP_32_5_32_test_1 C476 ( .D0_31(_RegFile_0__0), .D0_30(
        _RegFile_0__1), .D0_29(_RegFile_0__2), .D0_28(_RegFile_0__3), .D0_27(
        _RegFile_0__4), .D0_26(_RegFile_0__5), .D0_25(_RegFile_0__6), .D0_24(
        _RegFile_0__7), .D0_23(_RegFile_0__8), .D0_22(_RegFile_0__9), .D0_21(
        _RegFile_0__10), .D0_20(_RegFile_0__11), .D0_19(_RegFile_0__12), 
        .D0_18(_RegFile_0__13), .D0_17(_RegFile_0__14), .D0_16(_RegFile_0__15), 
        .D0_15(_RegFile_0__16), .D0_14(_RegFile_0__17), .D0_13(_RegFile_0__18), 
        .D0_12(_RegFile_0__19), .D0_11(_RegFile_0__20), .D0_10(_RegFile_0__21), 
        .D0_9(_RegFile_0__22), .D0_8(_RegFile_0__23), .D0_7(_RegFile_0__24), 
        .D0_6(_RegFile_0__25), .D0_5(_RegFile_0__26), .D0_4(_RegFile_0__27), 
        .D0_3(_RegFile_0__28), .D0_2(_RegFile_0__29), .D0_1(_RegFile_0__30), 
        .D0_0(_RegFile_0__31), .D1_31(_RegFile_1__0), .D1_30(_RegFile_1__1), 
        .D1_29(_RegFile_1__2), .D1_28(_RegFile_1__3), .D1_27(_RegFile_1__4), 
        .D1_26(_RegFile_1__5), .D1_25(_RegFile_1__6), .D1_24(_RegFile_1__7), 
        .D1_23(_RegFile_1__8), .D1_22(_RegFile_1__9), .D1_21(_RegFile_1__10), 
        .D1_20(_RegFile_1__11), .D1_19(_RegFile_1__12), .D1_18(_RegFile_1__13), 
        .D1_17(_RegFile_1__14), .D1_16(_RegFile_1__15), .D1_15(_RegFile_1__16), 
        .D1_14(_RegFile_1__17), .D1_13(_RegFile_1__18), .D1_12(_RegFile_1__19), 
        .D1_11(_RegFile_1__20), .D1_10(_RegFile_1__21), .D1_9(_RegFile_1__22), 
        .D1_8(_RegFile_1__23), .D1_7(_RegFile_1__24), .D1_6(_RegFile_1__25), 
        .D1_5(_RegFile_1__26), .D1_4(_RegFile_1__27), .D1_3(_RegFile_1__28), 
        .D1_2(_RegFile_1__29), .D1_1(_RegFile_1__30), .D1_0(_RegFile_1__31), 
        .D2_31(_RegFile_2__0), .D2_30(_RegFile_2__1), .D2_29(_RegFile_2__2), 
        .D2_28(_RegFile_2__3), .D2_27(_RegFile_2__4), .D2_26(_RegFile_2__5), 
        .D2_25(_RegFile_2__6), .D2_24(_RegFile_2__7), .D2_23(_RegFile_2__8), 
        .D2_22(_RegFile_2__9), .D2_21(_RegFile_2__10), .D2_20(_RegFile_2__11), 
        .D2_19(_RegFile_2__12), .D2_18(_RegFile_2__13), .D2_17(_RegFile_2__14), 
        .D2_16(_RegFile_2__15), .D2_15(_RegFile_2__16), .D2_14(_RegFile_2__17), 
        .D2_13(_RegFile_2__18), .D2_12(_RegFile_2__19), .D2_11(_RegFile_2__20), 
        .D2_10(_RegFile_2__21), .D2_9(_RegFile_2__22), .D2_8(_RegFile_2__23), 
        .D2_7(_RegFile_2__24), .D2_6(_RegFile_2__25), .D2_5(_RegFile_2__26), 
        .D2_4(_RegFile_2__27), .D2_3(_RegFile_2__28), .D2_2(_RegFile_2__29), 
        .D2_1(_RegFile_2__30), .D2_0(_RegFile_2__31), .D3_31(_RegFile_3__0), 
        .D3_30(_RegFile_3__1), .D3_29(_RegFile_3__2), .D3_28(_RegFile_3__3), 
        .D3_27(_RegFile_3__4), .D3_26(_RegFile_3__5), .D3_25(_RegFile_3__6), 
        .D3_24(_RegFile_3__7), .D3_23(_RegFile_3__8), .D3_22(_RegFile_3__9), 
        .D3_21(_RegFile_3__10), .D3_20(_RegFile_3__11), .D3_19(_RegFile_3__12), 
        .D3_18(_RegFile_3__13), .D3_17(_RegFile_3__14), .D3_16(_RegFile_3__15), 
        .D3_15(_RegFile_3__16), .D3_14(_RegFile_3__17), .D3_13(_RegFile_3__18), 
        .D3_12(_RegFile_3__19), .D3_11(_RegFile_3__20), .D3_10(_RegFile_3__21), 
        .D3_9(_RegFile_3__22), .D3_8(_RegFile_3__23), .D3_7(_RegFile_3__24), 
        .D3_6(_RegFile_3__25), .D3_5(_RegFile_3__26), .D3_4(_RegFile_3__27), 
        .D3_3(_RegFile_3__28), .D3_2(_RegFile_3__29), .D3_1(_RegFile_3__30), 
        .D3_0(_RegFile_3__31), .D4_31(_RegFile_4__0), .D4_30(_RegFile_4__1), 
        .D4_29(_RegFile_4__2), .D4_28(_RegFile_4__3), .D4_27(_RegFile_4__4), 
        .D4_26(_RegFile_4__5), .D4_25(_RegFile_4__6), .D4_24(_RegFile_4__7), 
        .D4_23(_RegFile_4__8), .D4_22(_RegFile_4__9), .D4_21(_RegFile_4__10), 
        .D4_20(_RegFile_4__11), .D4_19(_RegFile_4__12), .D4_18(_RegFile_4__13), 
        .D4_17(_RegFile_4__14), .D4_16(_RegFile_4__15), .D4_15(_RegFile_4__16), 
        .D4_14(_RegFile_4__17), .D4_13(_RegFile_4__18), .D4_12(_RegFile_4__19), 
        .D4_11(_RegFile_4__20), .D4_10(_RegFile_4__21), .D4_9(_RegFile_4__22), 
        .D4_8(_RegFile_4__23), .D4_7(_RegFile_4__24), .D4_6(_RegFile_4__25), 
        .D4_5(_RegFile_4__26), .D4_4(_RegFile_4__27), .D4_3(_RegFile_4__28), 
        .D4_2(_RegFile_4__29), .D4_1(_RegFile_4__30), .D4_0(_RegFile_4__31), 
        .D5_31(_RegFile_5__0), .D5_30(_RegFile_5__1), .D5_29(_RegFile_5__2), 
        .D5_28(_RegFile_5__3), .D5_27(_RegFile_5__4), .D5_26(_RegFile_5__5), 
        .D5_25(_RegFile_5__6), .D5_24(_RegFile_5__7), .D5_23(_RegFile_5__8), 
        .D5_22(_RegFile_5__9), .D5_21(_RegFile_5__10), .D5_20(_RegFile_5__11), 
        .D5_19(_RegFile_5__12), .D5_18(_RegFile_5__13), .D5_17(_RegFile_5__14), 
        .D5_16(_RegFile_5__15), .D5_15(_RegFile_5__16), .D5_14(_RegFile_5__17), 
        .D5_13(_RegFile_5__18), .D5_12(_RegFile_5__19), .D5_11(_RegFile_5__20), 
        .D5_10(_RegFile_5__21), .D5_9(_RegFile_5__22), .D5_8(_RegFile_5__23), 
        .D5_7(_RegFile_5__24), .D5_6(_RegFile_5__25), .D5_5(_RegFile_5__26), 
        .D5_4(_RegFile_5__27), .D5_3(_RegFile_5__28), .D5_2(_RegFile_5__29), 
        .D5_1(_RegFile_5__30), .D5_0(_RegFile_5__31), .D6_31(_RegFile_6__0), 
        .D6_30(_RegFile_6__1), .D6_29(_RegFile_6__2), .D6_28(_RegFile_6__3), 
        .D6_27(_RegFile_6__4), .D6_26(_RegFile_6__5), .D6_25(_RegFile_6__6), 
        .D6_24(_RegFile_6__7), .D6_23(_RegFile_6__8), .D6_22(_RegFile_6__9), 
        .D6_21(_RegFile_6__10), .D6_20(_RegFile_6__11), .D6_19(_RegFile_6__12), 
        .D6_18(_RegFile_6__13), .D6_17(_RegFile_6__14), .D6_16(_RegFile_6__15), 
        .D6_15(_RegFile_6__16), .D6_14(_RegFile_6__17), .D6_13(_RegFile_6__18), 
        .D6_12(_RegFile_6__19), .D6_11(_RegFile_6__20), .D6_10(_RegFile_6__21), 
        .D6_9(_RegFile_6__22), .D6_8(_RegFile_6__23), .D6_7(_RegFile_6__24), 
        .D6_6(_RegFile_6__25), .D6_5(_RegFile_6__26), .D6_4(_RegFile_6__27), 
        .D6_3(_RegFile_6__28), .D6_2(_RegFile_6__29), .D6_1(_RegFile_6__30), 
        .D6_0(_RegFile_6__31), .D7_31(_RegFile_7__0), .D7_30(_RegFile_7__1), 
        .D7_29(_RegFile_7__2), .D7_28(_RegFile_7__3), .D7_27(_RegFile_7__4), 
        .D7_26(_RegFile_7__5), .D7_25(_RegFile_7__6), .D7_24(_RegFile_7__7), 
        .D7_23(_RegFile_7__8), .D7_22(_RegFile_7__9), .D7_21(_RegFile_7__10), 
        .D7_20(_RegFile_7__11), .D7_19(_RegFile_7__12), .D7_18(_RegFile_7__13), 
        .D7_17(_RegFile_7__14), .D7_16(_RegFile_7__15), .D7_15(_RegFile_7__16), 
        .D7_14(_RegFile_7__17), .D7_13(_RegFile_7__18), .D7_12(_RegFile_7__19), 
        .D7_11(_RegFile_7__20), .D7_10(_RegFile_7__21), .D7_9(_RegFile_7__22), 
        .D7_8(_RegFile_7__23), .D7_7(_RegFile_7__24), .D7_6(_RegFile_7__25), 
        .D7_5(_RegFile_7__26), .D7_4(_RegFile_7__27), .D7_3(_RegFile_7__28), 
        .D7_2(_RegFile_7__29), .D7_1(_RegFile_7__30), .D7_0(_RegFile_7__31), 
        .D8_31(_RegFile_8__0), .D8_30(_RegFile_8__1), .D8_29(_RegFile_8__2), 
        .D8_28(_RegFile_8__3), .D8_27(_RegFile_8__4), .D8_26(_RegFile_8__5), 
        .D8_25(_RegFile_8__6), .D8_24(_RegFile_8__7), .D8_23(_RegFile_8__8), 
        .D8_22(_RegFile_8__9), .D8_21(_RegFile_8__10), .D8_20(_RegFile_8__11), 
        .D8_19(_RegFile_8__12), .D8_18(_RegFile_8__13), .D8_17(_RegFile_8__14), 
        .D8_16(_RegFile_8__15), .D8_15(_RegFile_8__16), .D8_14(_RegFile_8__17), 
        .D8_13(_RegFile_8__18), .D8_12(_RegFile_8__19), .D8_11(_RegFile_8__20), 
        .D8_10(_RegFile_8__21), .D8_9(_RegFile_8__22), .D8_8(_RegFile_8__23), 
        .D8_7(_RegFile_8__24), .D8_6(_RegFile_8__25), .D8_5(_RegFile_8__26), 
        .D8_4(_RegFile_8__27), .D8_3(_RegFile_8__28), .D8_2(_RegFile_8__29), 
        .D8_1(_RegFile_8__30), .D8_0(_RegFile_8__31), .D9_31(_RegFile_9__0), 
        .D9_30(_RegFile_9__1), .D9_29(_RegFile_9__2), .D9_28(_RegFile_9__3), 
        .D9_27(_RegFile_9__4), .D9_26(_RegFile_9__5), .D9_25(_RegFile_9__6), 
        .D9_24(_RegFile_9__7), .D9_23(_RegFile_9__8), .D9_22(_RegFile_9__9), 
        .D9_21(_RegFile_9__10), .D9_20(_RegFile_9__11), .D9_19(_RegFile_9__12), 
        .D9_18(_RegFile_9__13), .D9_17(_RegFile_9__14), .D9_16(_RegFile_9__15), 
        .D9_15(_RegFile_9__16), .D9_14(_RegFile_9__17), .D9_13(_RegFile_9__18), 
        .D9_12(_RegFile_9__19), .D9_11(_RegFile_9__20), .D9_10(_RegFile_9__21), 
        .D9_9(_RegFile_9__22), .D9_8(_RegFile_9__23), .D9_7(_RegFile_9__24), 
        .D9_6(_RegFile_9__25), .D9_5(_RegFile_9__26), .D9_4(_RegFile_9__27), 
        .D9_3(_RegFile_9__28), .D9_2(_RegFile_9__29), .D9_1(_RegFile_9__30), 
        .D9_0(_RegFile_9__31), .D10_31(_RegFile_10__0), .D10_30(_RegFile_10__1
        ), .D10_29(_RegFile_10__2), .D10_28(_RegFile_10__3), .D10_27(
        _RegFile_10__4), .D10_26(_RegFile_10__5), .D10_25(_RegFile_10__6), 
        .D10_24(_RegFile_10__7), .D10_23(_RegFile_10__8), .D10_22(
        _RegFile_10__9), .D10_21(_RegFile_10__10), .D10_20(_RegFile_10__11), 
        .D10_19(_RegFile_10__12), .D10_18(_RegFile_10__13), .D10_17(
        _RegFile_10__14), .D10_16(_RegFile_10__15), .D10_15(_RegFile_10__16), 
        .D10_14(_RegFile_10__17), .D10_13(_RegFile_10__18), .D10_12(
        _RegFile_10__19), .D10_11(_RegFile_10__20), .D10_10(_RegFile_10__21), 
        .D10_9(_RegFile_10__22), .D10_8(_RegFile_10__23), .D10_7(
        _RegFile_10__24), .D10_6(_RegFile_10__25), .D10_5(_RegFile_10__26), 
        .D10_4(_RegFile_10__27), .D10_3(_RegFile_10__28), .D10_2(
        _RegFile_10__29), .D10_1(_RegFile_10__30), .D10_0(_RegFile_10__31), 
        .D11_31(_RegFile_11__0), .D11_30(_RegFile_11__1), .D11_29(
        _RegFile_11__2), .D11_28(_RegFile_11__3), .D11_27(_RegFile_11__4), 
        .D11_26(_RegFile_11__5), .D11_25(_RegFile_11__6), .D11_24(
        _RegFile_11__7), .D11_23(_RegFile_11__8), .D11_22(_RegFile_11__9), 
        .D11_21(_RegFile_11__10), .D11_20(_RegFile_11__11), .D11_19(
        _RegFile_11__12), .D11_18(_RegFile_11__13), .D11_17(_RegFile_11__14), 
        .D11_16(_RegFile_11__15), .D11_15(_RegFile_11__16), .D11_14(
        _RegFile_11__17), .D11_13(_RegFile_11__18), .D11_12(_RegFile_11__19), 
        .D11_11(_RegFile_11__20), .D11_10(_RegFile_11__21), .D11_9(
        _RegFile_11__22), .D11_8(_RegFile_11__23), .D11_7(_RegFile_11__24), 
        .D11_6(_RegFile_11__25), .D11_5(_RegFile_11__26), .D11_4(
        _RegFile_11__27), .D11_3(_RegFile_11__28), .D11_2(_RegFile_11__29), 
        .D11_1(_RegFile_11__30), .D11_0(_RegFile_11__31), .D12_31(
        _RegFile_12__0), .D12_30(_RegFile_12__1), .D12_29(_RegFile_12__2), 
        .D12_28(_RegFile_12__3), .D12_27(_RegFile_12__4), .D12_26(
        _RegFile_12__5), .D12_25(_RegFile_12__6), .D12_24(_RegFile_12__7), 
        .D12_23(_RegFile_12__8), .D12_22(_RegFile_12__9), .D12_21(
        _RegFile_12__10), .D12_20(_RegFile_12__11), .D12_19(_RegFile_12__12), 
        .D12_18(_RegFile_12__13), .D12_17(_RegFile_12__14), .D12_16(
        _RegFile_12__15), .D12_15(_RegFile_12__16), .D12_14(_RegFile_12__17), 
        .D12_13(_RegFile_12__18), .D12_12(_RegFile_12__19), .D12_11(
        _RegFile_12__20), .D12_10(_RegFile_12__21), .D12_9(_RegFile_12__22), 
        .D12_8(_RegFile_12__23), .D12_7(_RegFile_12__24), .D12_6(
        _RegFile_12__25), .D12_5(_RegFile_12__26), .D12_4(_RegFile_12__27), 
        .D12_3(_RegFile_12__28), .D12_2(_RegFile_12__29), .D12_1(
        _RegFile_12__30), .D12_0(_RegFile_12__31), .D13_31(_RegFile_13__0), 
        .D13_30(_RegFile_13__1), .D13_29(_RegFile_13__2), .D13_28(
        _RegFile_13__3), .D13_27(_RegFile_13__4), .D13_26(_RegFile_13__5), 
        .D13_25(_RegFile_13__6), .D13_24(_RegFile_13__7), .D13_23(
        _RegFile_13__8), .D13_22(_RegFile_13__9), .D13_21(_RegFile_13__10), 
        .D13_20(_RegFile_13__11), .D13_19(_RegFile_13__12), .D13_18(
        _RegFile_13__13), .D13_17(_RegFile_13__14), .D13_16(_RegFile_13__15), 
        .D13_15(_RegFile_13__16), .D13_14(_RegFile_13__17), .D13_13(
        _RegFile_13__18), .D13_12(_RegFile_13__19), .D13_11(_RegFile_13__20), 
        .D13_10(_RegFile_13__21), .D13_9(_RegFile_13__22), .D13_8(
        _RegFile_13__23), .D13_7(_RegFile_13__24), .D13_6(_RegFile_13__25), 
        .D13_5(_RegFile_13__26), .D13_4(_RegFile_13__27), .D13_3(
        _RegFile_13__28), .D13_2(_RegFile_13__29), .D13_1(_RegFile_13__30), 
        .D13_0(_RegFile_13__31), .D14_31(_RegFile_14__0), .D14_30(
        _RegFile_14__1), .D14_29(_RegFile_14__2), .D14_28(_RegFile_14__3), 
        .D14_27(_RegFile_14__4), .D14_26(_RegFile_14__5), .D14_25(
        _RegFile_14__6), .D14_24(_RegFile_14__7), .D14_23(_RegFile_14__8), 
        .D14_22(_RegFile_14__9), .D14_21(_RegFile_14__10), .D14_20(
        _RegFile_14__11), .D14_19(_RegFile_14__12), .D14_18(_RegFile_14__13), 
        .D14_17(_RegFile_14__14), .D14_16(_RegFile_14__15), .D14_15(
        _RegFile_14__16), .D14_14(_RegFile_14__17), .D14_13(_RegFile_14__18), 
        .D14_12(_RegFile_14__19), .D14_11(_RegFile_14__20), .D14_10(
        _RegFile_14__21), .D14_9(_RegFile_14__22), .D14_8(_RegFile_14__23), 
        .D14_7(_RegFile_14__24), .D14_6(_RegFile_14__25), .D14_5(
        _RegFile_14__26), .D14_4(_RegFile_14__27), .D14_3(_RegFile_14__28), 
        .D14_2(_RegFile_14__29), .D14_1(_RegFile_14__30), .D14_0(
        _RegFile_14__31), .D15_31(_RegFile_15__0), .D15_30(_RegFile_15__1), 
        .D15_29(_RegFile_15__2), .D15_28(_RegFile_15__3), .D15_27(
        _RegFile_15__4), .D15_26(_RegFile_15__5), .D15_25(_RegFile_15__6), 
        .D15_24(_RegFile_15__7), .D15_23(_RegFile_15__8), .D15_22(
        _RegFile_15__9), .D15_21(_RegFile_15__10), .D15_20(_RegFile_15__11), 
        .D15_19(_RegFile_15__12), .D15_18(_RegFile_15__13), .D15_17(
        _RegFile_15__14), .D15_16(_RegFile_15__15), .D15_15(_RegFile_15__16), 
        .D15_14(_RegFile_15__17), .D15_13(_RegFile_15__18), .D15_12(
        _RegFile_15__19), .D15_11(_RegFile_15__20), .D15_10(_RegFile_15__21), 
        .D15_9(_RegFile_15__22), .D15_8(_RegFile_15__23), .D15_7(
        _RegFile_15__24), .D15_6(_RegFile_15__25), .D15_5(_RegFile_15__26), 
        .D15_4(_RegFile_15__27), .D15_3(_RegFile_15__28), .D15_2(
        _RegFile_15__29), .D15_1(_RegFile_15__30), .D15_0(_RegFile_15__31), 
        .D16_31(_RegFile_16__0), .D16_30(_RegFile_16__1), .D16_29(
        _RegFile_16__2), .D16_28(_RegFile_16__3), .D16_27(_RegFile_16__4), 
        .D16_26(_RegFile_16__5), .D16_25(_RegFile_16__6), .D16_24(
        _RegFile_16__7), .D16_23(_RegFile_16__8), .D16_22(_RegFile_16__9), 
        .D16_21(_RegFile_16__10), .D16_20(_RegFile_16__11), .D16_19(
        _RegFile_16__12), .D16_18(_RegFile_16__13), .D16_17(_RegFile_16__14), 
        .D16_16(_RegFile_16__15), .D16_15(_RegFile_16__16), .D16_14(
        _RegFile_16__17), .D16_13(_RegFile_16__18), .D16_12(_RegFile_16__19), 
        .D16_11(_RegFile_16__20), .D16_10(_RegFile_16__21), .D16_9(
        _RegFile_16__22), .D16_8(_RegFile_16__23), .D16_7(_RegFile_16__24), 
        .D16_6(_RegFile_16__25), .D16_5(_RegFile_16__26), .D16_4(
        _RegFile_16__27), .D16_3(_RegFile_16__28), .D16_2(_RegFile_16__29), 
        .D16_1(_RegFile_16__30), .D16_0(_RegFile_16__31), .D17_31(
        _RegFile_17__0), .D17_30(_RegFile_17__1), .D17_29(_RegFile_17__2), 
        .D17_28(_RegFile_17__3), .D17_27(_RegFile_17__4), .D17_26(
        _RegFile_17__5), .D17_25(_RegFile_17__6), .D17_24(_RegFile_17__7), 
        .D17_23(_RegFile_17__8), .D17_22(_RegFile_17__9), .D17_21(
        _RegFile_17__10), .D17_20(_RegFile_17__11), .D17_19(_RegFile_17__12), 
        .D17_18(_RegFile_17__13), .D17_17(_RegFile_17__14), .D17_16(
        _RegFile_17__15), .D17_15(_RegFile_17__16), .D17_14(_RegFile_17__17), 
        .D17_13(_RegFile_17__18), .D17_12(_RegFile_17__19), .D17_11(
        _RegFile_17__20), .D17_10(_RegFile_17__21), .D17_9(_RegFile_17__22), 
        .D17_8(_RegFile_17__23), .D17_7(_RegFile_17__24), .D17_6(
        _RegFile_17__25), .D17_5(_RegFile_17__26), .D17_4(_RegFile_17__27), 
        .D17_3(_RegFile_17__28), .D17_2(_RegFile_17__29), .D17_1(
        _RegFile_17__30), .D17_0(_RegFile_17__31), .D18_31(_RegFile_18__0), 
        .D18_30(_RegFile_18__1), .D18_29(_RegFile_18__2), .D18_28(
        _RegFile_18__3), .D18_27(_RegFile_18__4), .D18_26(_RegFile_18__5), 
        .D18_25(_RegFile_18__6), .D18_24(_RegFile_18__7), .D18_23(
        _RegFile_18__8), .D18_22(_RegFile_18__9), .D18_21(_RegFile_18__10), 
        .D18_20(_RegFile_18__11), .D18_19(_RegFile_18__12), .D18_18(
        _RegFile_18__13), .D18_17(_RegFile_18__14), .D18_16(_RegFile_18__15), 
        .D18_15(_RegFile_18__16), .D18_14(_RegFile_18__17), .D18_13(
        _RegFile_18__18), .D18_12(_RegFile_18__19), .D18_11(_RegFile_18__20), 
        .D18_10(_RegFile_18__21), .D18_9(_RegFile_18__22), .D18_8(
        _RegFile_18__23), .D18_7(_RegFile_18__24), .D18_6(_RegFile_18__25), 
        .D18_5(_RegFile_18__26), .D18_4(_RegFile_18__27), .D18_3(
        _RegFile_18__28), .D18_2(_RegFile_18__29), .D18_1(_RegFile_18__30), 
        .D18_0(_RegFile_18__31), .D19_31(_RegFile_19__0), .D19_30(
        _RegFile_19__1), .D19_29(_RegFile_19__2), .D19_28(_RegFile_19__3), 
        .D19_27(_RegFile_19__4), .D19_26(_RegFile_19__5), .D19_25(
        _RegFile_19__6), .D19_24(_RegFile_19__7), .D19_23(_RegFile_19__8), 
        .D19_22(_RegFile_19__9), .D19_21(_RegFile_19__10), .D19_20(
        _RegFile_19__11), .D19_19(_RegFile_19__12), .D19_18(_RegFile_19__13), 
        .D19_17(_RegFile_19__14), .D19_16(_RegFile_19__15), .D19_15(
        _RegFile_19__16), .D19_14(_RegFile_19__17), .D19_13(_RegFile_19__18), 
        .D19_12(_RegFile_19__19), .D19_11(_RegFile_19__20), .D19_10(
        _RegFile_19__21), .D19_9(_RegFile_19__22), .D19_8(_RegFile_19__23), 
        .D19_7(_RegFile_19__24), .D19_6(_RegFile_19__25), .D19_5(
        _RegFile_19__26), .D19_4(_RegFile_19__27), .D19_3(_RegFile_19__28), 
        .D19_2(_RegFile_19__29), .D19_1(_RegFile_19__30), .D19_0(
        _RegFile_19__31), .D20_31(_RegFile_20__0), .D20_30(_RegFile_20__1), 
        .D20_29(_RegFile_20__2), .D20_28(_RegFile_20__3), .D20_27(
        _RegFile_20__4), .D20_26(_RegFile_20__5), .D20_25(_RegFile_20__6), 
        .D20_24(_RegFile_20__7), .D20_23(_RegFile_20__8), .D20_22(
        _RegFile_20__9), .D20_21(_RegFile_20__10), .D20_20(_RegFile_20__11), 
        .D20_19(_RegFile_20__12), .D20_18(_RegFile_20__13), .D20_17(
        _RegFile_20__14), .D20_16(_RegFile_20__15), .D20_15(_RegFile_20__16), 
        .D20_14(_RegFile_20__17), .D20_13(_RegFile_20__18), .D20_12(
        _RegFile_20__19), .D20_11(_RegFile_20__20), .D20_10(_RegFile_20__21), 
        .D20_9(_RegFile_20__22), .D20_8(_RegFile_20__23), .D20_7(
        _RegFile_20__24), .D20_6(_RegFile_20__25), .D20_5(_RegFile_20__26), 
        .D20_4(_RegFile_20__27), .D20_3(_RegFile_20__28), .D20_2(
        _RegFile_20__29), .D20_1(_RegFile_20__30), .D20_0(_RegFile_20__31), 
        .D21_31(_RegFile_21__0), .D21_30(_RegFile_21__1), .D21_29(
        _RegFile_21__2), .D21_28(_RegFile_21__3), .D21_27(_RegFile_21__4), 
        .D21_26(_RegFile_21__5), .D21_25(_RegFile_21__6), .D21_24(
        _RegFile_21__7), .D21_23(_RegFile_21__8), .D21_22(_RegFile_21__9), 
        .D21_21(_RegFile_21__10), .D21_20(_RegFile_21__11), .D21_19(
        _RegFile_21__12), .D21_18(_RegFile_21__13), .D21_17(_RegFile_21__14), 
        .D21_16(_RegFile_21__15), .D21_15(_RegFile_21__16), .D21_14(
        _RegFile_21__17), .D21_13(_RegFile_21__18), .D21_12(_RegFile_21__19), 
        .D21_11(_RegFile_21__20), .D21_10(_RegFile_21__21), .D21_9(
        _RegFile_21__22), .D21_8(_RegFile_21__23), .D21_7(_RegFile_21__24), 
        .D21_6(_RegFile_21__25), .D21_5(_RegFile_21__26), .D21_4(
        _RegFile_21__27), .D21_3(_RegFile_21__28), .D21_2(_RegFile_21__29), 
        .D21_1(_RegFile_21__30), .D21_0(_RegFile_21__31), .D22_31(
        _RegFile_22__0), .D22_30(_RegFile_22__1), .D22_29(_RegFile_22__2), 
        .D22_28(_RegFile_22__3), .D22_27(_RegFile_22__4), .D22_26(
        _RegFile_22__5), .D22_25(_RegFile_22__6), .D22_24(_RegFile_22__7), 
        .D22_23(_RegFile_22__8), .D22_22(_RegFile_22__9), .D22_21(
        _RegFile_22__10), .D22_20(_RegFile_22__11), .D22_19(_RegFile_22__12), 
        .D22_18(_RegFile_22__13), .D22_17(_RegFile_22__14), .D22_16(
        _RegFile_22__15), .D22_15(_RegFile_22__16), .D22_14(_RegFile_22__17), 
        .D22_13(_RegFile_22__18), .D22_12(_RegFile_22__19), .D22_11(
        _RegFile_22__20), .D22_10(_RegFile_22__21), .D22_9(_RegFile_22__22), 
        .D22_8(_RegFile_22__23), .D22_7(_RegFile_22__24), .D22_6(
        _RegFile_22__25), .D22_5(_RegFile_22__26), .D22_4(_RegFile_22__27), 
        .D22_3(_RegFile_22__28), .D22_2(_RegFile_22__29), .D22_1(
        _RegFile_22__30), .D22_0(_RegFile_22__31), .D23_31(_RegFile_23__0), 
        .D23_30(_RegFile_23__1), .D23_29(_RegFile_23__2), .D23_28(
        _RegFile_23__3), .D23_27(_RegFile_23__4), .D23_26(_RegFile_23__5), 
        .D23_25(_RegFile_23__6), .D23_24(_RegFile_23__7), .D23_23(
        _RegFile_23__8), .D23_22(_RegFile_23__9), .D23_21(_RegFile_23__10), 
        .D23_20(_RegFile_23__11), .D23_19(_RegFile_23__12), .D23_18(
        _RegFile_23__13), .D23_17(_RegFile_23__14), .D23_16(_RegFile_23__15), 
        .D23_15(_RegFile_23__16), .D23_14(_RegFile_23__17), .D23_13(
        _RegFile_23__18), .D23_12(_RegFile_23__19), .D23_11(_RegFile_23__20), 
        .D23_10(_RegFile_23__21), .D23_9(_RegFile_23__22), .D23_8(
        _RegFile_23__23), .D23_7(_RegFile_23__24), .D23_6(_RegFile_23__25), 
        .D23_5(_RegFile_23__26), .D23_4(_RegFile_23__27), .D23_3(
        _RegFile_23__28), .D23_2(_RegFile_23__29), .D23_1(_RegFile_23__30), 
        .D23_0(_RegFile_23__31), .D24_31(_RegFile_24__0), .D24_30(
        _RegFile_24__1), .D24_29(_RegFile_24__2), .D24_28(_RegFile_24__3), 
        .D24_27(_RegFile_24__4), .D24_26(_RegFile_24__5), .D24_25(
        _RegFile_24__6), .D24_24(_RegFile_24__7), .D24_23(_RegFile_24__8), 
        .D24_22(_RegFile_24__9), .D24_21(_RegFile_24__10), .D24_20(
        _RegFile_24__11), .D24_19(_RegFile_24__12), .D24_18(_RegFile_24__13), 
        .D24_17(_RegFile_24__14), .D24_16(_RegFile_24__15), .D24_15(
        _RegFile_24__16), .D24_14(_RegFile_24__17), .D24_13(_RegFile_24__18), 
        .D24_12(_RegFile_24__19), .D24_11(_RegFile_24__20), .D24_10(
        _RegFile_24__21), .D24_9(_RegFile_24__22), .D24_8(_RegFile_24__23), 
        .D24_7(_RegFile_24__24), .D24_6(_RegFile_24__25), .D24_5(
        _RegFile_24__26), .D24_4(_RegFile_24__27), .D24_3(_RegFile_24__28), 
        .D24_2(_RegFile_24__29), .D24_1(_RegFile_24__30), .D24_0(
        _RegFile_24__31), .D25_31(_RegFile_25__0), .D25_30(_RegFile_25__1), 
        .D25_29(_RegFile_25__2), .D25_28(_RegFile_25__3), .D25_27(
        _RegFile_25__4), .D25_26(_RegFile_25__5), .D25_25(_RegFile_25__6), 
        .D25_24(_RegFile_25__7), .D25_23(_RegFile_25__8), .D25_22(
        _RegFile_25__9), .D25_21(_RegFile_25__10), .D25_20(_RegFile_25__11), 
        .D25_19(_RegFile_25__12), .D25_18(_RegFile_25__13), .D25_17(
        _RegFile_25__14), .D25_16(_RegFile_25__15), .D25_15(_RegFile_25__16), 
        .D25_14(_RegFile_25__17), .D25_13(_RegFile_25__18), .D25_12(
        _RegFile_25__19), .D25_11(_RegFile_25__20), .D25_10(_RegFile_25__21), 
        .D25_9(_RegFile_25__22), .D25_8(_RegFile_25__23), .D25_7(
        _RegFile_25__24), .D25_6(_RegFile_25__25), .D25_5(_RegFile_25__26), 
        .D25_4(_RegFile_25__27), .D25_3(_RegFile_25__28), .D25_2(
        _RegFile_25__29), .D25_1(_RegFile_25__30), .D25_0(_RegFile_25__31), 
        .D26_31(_RegFile_26__0), .D26_30(_RegFile_26__1), .D26_29(
        _RegFile_26__2), .D26_28(_RegFile_26__3), .D26_27(_RegFile_26__4), 
        .D26_26(_RegFile_26__5), .D26_25(_RegFile_26__6), .D26_24(
        _RegFile_26__7), .D26_23(_RegFile_26__8), .D26_22(_RegFile_26__9), 
        .D26_21(_RegFile_26__10), .D26_20(_RegFile_26__11), .D26_19(
        _RegFile_26__12), .D26_18(_RegFile_26__13), .D26_17(_RegFile_26__14), 
        .D26_16(_RegFile_26__15), .D26_15(_RegFile_26__16), .D26_14(
        _RegFile_26__17), .D26_13(_RegFile_26__18), .D26_12(_RegFile_26__19), 
        .D26_11(_RegFile_26__20), .D26_10(_RegFile_26__21), .D26_9(
        _RegFile_26__22), .D26_8(_RegFile_26__23), .D26_7(_RegFile_26__24), 
        .D26_6(_RegFile_26__25), .D26_5(_RegFile_26__26), .D26_4(
        _RegFile_26__27), .D26_3(_RegFile_26__28), .D26_2(_RegFile_26__29), 
        .D26_1(_RegFile_26__30), .D26_0(_RegFile_26__31), .D27_31(
        _RegFile_27__0), .D27_30(_RegFile_27__1), .D27_29(_RegFile_27__2), 
        .D27_28(_RegFile_27__3), .D27_27(_RegFile_27__4), .D27_26(
        _RegFile_27__5), .D27_25(_RegFile_27__6), .D27_24(_RegFile_27__7), 
        .D27_23(_RegFile_27__8), .D27_22(_RegFile_27__9), .D27_21(
        _RegFile_27__10), .D27_20(_RegFile_27__11), .D27_19(_RegFile_27__12), 
        .D27_18(_RegFile_27__13), .D27_17(_RegFile_27__14), .D27_16(
        _RegFile_27__15), .D27_15(_RegFile_27__16), .D27_14(_RegFile_27__17), 
        .D27_13(_RegFile_27__18), .D27_12(_RegFile_27__19), .D27_11(
        _RegFile_27__20), .D27_10(_RegFile_27__21), .D27_9(_RegFile_27__22), 
        .D27_8(_RegFile_27__23), .D27_7(_RegFile_27__24), .D27_6(
        _RegFile_27__25), .D27_5(_RegFile_27__26), .D27_4(_RegFile_27__27), 
        .D27_3(_RegFile_27__28), .D27_2(_RegFile_27__29), .D27_1(
        _RegFile_27__30), .D27_0(_RegFile_27__31), .D28_31(_RegFile_28__0), 
        .D28_30(_RegFile_28__1), .D28_29(_RegFile_28__2), .D28_28(
        _RegFile_28__3), .D28_27(_RegFile_28__4), .D28_26(_RegFile_28__5), 
        .D28_25(_RegFile_28__6), .D28_24(_RegFile_28__7), .D28_23(
        _RegFile_28__8), .D28_22(_RegFile_28__9), .D28_21(_RegFile_28__10), 
        .D28_20(_RegFile_28__11), .D28_19(_RegFile_28__12), .D28_18(
        _RegFile_28__13), .D28_17(_RegFile_28__14), .D28_16(_RegFile_28__15), 
        .D28_15(_RegFile_28__16), .D28_14(_RegFile_28__17), .D28_13(
        _RegFile_28__18), .D28_12(_RegFile_28__19), .D28_11(_RegFile_28__20), 
        .D28_10(_RegFile_28__21), .D28_9(_RegFile_28__22), .D28_8(
        _RegFile_28__23), .D28_7(_RegFile_28__24), .D28_6(_RegFile_28__25), 
        .D28_5(_RegFile_28__26), .D28_4(_RegFile_28__27), .D28_3(
        _RegFile_28__28), .D28_2(_RegFile_28__29), .D28_1(_RegFile_28__30), 
        .D28_0(_RegFile_28__31), .D29_31(_RegFile_29__0), .D29_30(
        _RegFile_29__1), .D29_29(_RegFile_29__2), .D29_28(_RegFile_29__3), 
        .D29_27(_RegFile_29__4), .D29_26(_RegFile_29__5), .D29_25(
        _RegFile_29__6), .D29_24(_RegFile_29__7), .D29_23(_RegFile_29__8), 
        .D29_22(_RegFile_29__9), .D29_21(_RegFile_29__10), .D29_20(
        _RegFile_29__11), .D29_19(_RegFile_29__12), .D29_18(_RegFile_29__13), 
        .D29_17(_RegFile_29__14), .D29_16(_RegFile_29__15), .D29_15(
        _RegFile_29__16), .D29_14(_RegFile_29__17), .D29_13(_RegFile_29__18), 
        .D29_12(_RegFile_29__19), .D29_11(_RegFile_29__20), .D29_10(
        _RegFile_29__21), .D29_9(_RegFile_29__22), .D29_8(_RegFile_29__23), 
        .D29_7(_RegFile_29__24), .D29_6(_RegFile_29__25), .D29_5(
        _RegFile_29__26), .D29_4(_RegFile_29__27), .D29_3(_RegFile_29__28), 
        .D29_2(_RegFile_29__29), .D29_1(_RegFile_29__30), .D29_0(
        _RegFile_29__31), .D30_31(_RegFile_30__0), .D30_30(_RegFile_30__1), 
        .D30_29(_RegFile_30__2), .D30_28(_RegFile_30__3), .D30_27(
        _RegFile_30__4), .D30_26(_RegFile_30__5), .D30_25(_RegFile_30__6), 
        .D30_24(_RegFile_30__7), .D30_23(_RegFile_30__8), .D30_22(
        _RegFile_30__9), .D30_21(_RegFile_30__10), .D30_20(_RegFile_30__11), 
        .D30_19(_RegFile_30__12), .D30_18(_RegFile_30__13), .D30_17(
        _RegFile_30__14), .D30_16(_RegFile_30__15), .D30_15(_RegFile_30__16), 
        .D30_14(_RegFile_30__17), .D30_13(_RegFile_30__18), .D30_12(
        _RegFile_30__19), .D30_11(_RegFile_30__20), .D30_10(_RegFile_30__21), 
        .D30_9(_RegFile_30__22), .D30_8(_RegFile_30__23), .D30_7(
        _RegFile_30__24), .D30_6(_RegFile_30__25), .D30_5(_RegFile_30__26), 
        .D30_4(_RegFile_30__27), .D30_3(_RegFile_30__28), .D30_2(
        _RegFile_30__29), .D30_1(_RegFile_30__30), .D30_0(_RegFile_30__31), 
        .D31_31(_RegFile_31__0), .D31_30(_RegFile_31__1), .D31_29(
        _RegFile_31__2), .D31_28(_RegFile_31__3), .D31_27(_RegFile_31__4), 
        .D31_26(_RegFile_31__5), .D31_25(_RegFile_31__6), .D31_24(
        _RegFile_31__7), .D31_23(_RegFile_31__8), .D31_22(_RegFile_31__9), 
        .D31_21(_RegFile_31__10), .D31_20(_RegFile_31__11), .D31_19(
        _RegFile_31__12), .D31_18(_RegFile_31__13), .D31_17(_RegFile_31__14), 
        .D31_16(_RegFile_31__15), .D31_15(_RegFile_31__16), .D31_14(
        _RegFile_31__17), .D31_13(_RegFile_31__18), .D31_12(_RegFile_31__19), 
        .D31_11(_RegFile_31__20), .D31_10(_RegFile_31__21), .D31_9(
        _RegFile_31__22), .D31_8(_RegFile_31__23), .D31_7(_RegFile_31__24), 
        .D31_6(_RegFile_31__25), .D31_5(_RegFile_31__26), .D31_4(
        _RegFile_31__27), .D31_3(_RegFile_31__28), .D31_2(_RegFile_31__29), 
        .D31_1(_RegFile_31__30), .D31_0(_RegFile_31__31), .S0(n857), .S1(n339), 
        .S2(n848), .S3(n337), .S4(n802), .Z_31(N535), .Z_30(N534), .Z_29(N533), 
        .Z_28(N532), .Z_27(N531), .Z_26(N530), .Z_25(N529), .Z_24(N528), 
        .Z_23(N527), .Z_22(N526), .Z_21(N525), .Z_20(N524), .Z_19(N523), 
        .Z_18(N522), .Z_17(N521), .Z_16(N520), .Z_15(N519), .Z_14(N518), 
        .Z_13(N517), .Z_12(N516), .Z_11(N515), .Z_10(N514), .Z_9(N513), .Z_8(
        N512), .Z_7(N511), .Z_6(N510), .Z_5(N509), .Z_4(N508), .Z_3(N507), 
        .Z_2(N506), .Z_1(N505), .Z_0(N504) );
    smlatnr_1 CLI_reg__master ( .q(CLI_reg__m2s), .d(n2641), .sdi(test_si), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n953), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 CLI_reg__slave ( .q(CLI), .qb(n4386), .d(CLI_reg__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n953), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 Cause_Reg_reg_0__master ( .q(Cause_Reg_reg_0__m2s), .d(n2642), 
        .sdi(n4386), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n953), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 Cause_Reg_reg_0__slave ( .q(Cause_Reg_0), .qb(n627), .d(
        Cause_Reg_reg_0__m2s), .g(Ctrl__Regs_1__en2), .rb(n953), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 Cause_Reg_reg_10__master ( .q(Cause_Reg_reg_10__m2s), .d(n2652), 
        .sdi(n618), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n953), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 Cause_Reg_reg_10__slave ( .q(Cause_Reg_10), .qb(n617), .d(
        Cause_Reg_reg_10__m2s), .g(Ctrl__Regs_1__en2), .rb(n953), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 Cause_Reg_reg_11__master ( .q(Cause_Reg_reg_11__m2s), .d(n2653), 
        .sdi(n617), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n953), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 Cause_Reg_reg_11__slave ( .q(Cause_Reg_11), .qb(n616), .d(
        Cause_Reg_reg_11__m2s), .g(Ctrl__Regs_1__en2), .rb(n953), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 Cause_Reg_reg_12__master ( .q(Cause_Reg_reg_12__m2s), .d(n2654), 
        .sdi(n616), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n953), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 Cause_Reg_reg_12__slave ( .q(Cause_Reg_12), .qb(n615), .d(
        Cause_Reg_reg_12__m2s), .g(Ctrl__Regs_1__en2), .rb(n953), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 Cause_Reg_reg_13__master ( .q(Cause_Reg_reg_13__m2s), .d(n2655), 
        .sdi(n615), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n953), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 Cause_Reg_reg_13__slave ( .q(Cause_Reg_13), .qb(n614), .d(
        Cause_Reg_reg_13__m2s), .g(Ctrl__Regs_1__en2), .rb(n953), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 Cause_Reg_reg_14__master ( .q(Cause_Reg_reg_14__m2s), .d(n2656), 
        .sdi(n614), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n953), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 Cause_Reg_reg_14__slave ( .q(Cause_Reg_14), .qb(n613), .d(
        Cause_Reg_reg_14__m2s), .g(Ctrl__Regs_1__en2), .rb(n953), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 Cause_Reg_reg_15__master ( .q(Cause_Reg_reg_15__m2s), .d(n2657), 
        .sdi(n613), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n952), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 Cause_Reg_reg_15__slave ( .q(Cause_Reg_15), .qb(n612), .d(
        Cause_Reg_reg_15__m2s), .g(Ctrl__Regs_1__en2), .rb(n952), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 Cause_Reg_reg_16__master ( .q(Cause_Reg_reg_16__m2s), .d(n2658), 
        .sdi(n612), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n953), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 Cause_Reg_reg_16__slave ( .q(Cause_Reg_16), .qb(n611), .d(
        Cause_Reg_reg_16__m2s), .g(Ctrl__Regs_1__en2), .rb(n953), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 Cause_Reg_reg_17__master ( .q(Cause_Reg_reg_17__m2s), .d(n2659), 
        .sdi(n611), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n952), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 Cause_Reg_reg_17__slave ( .q(Cause_Reg_17), .qb(n610), .d(
        Cause_Reg_reg_17__m2s), .g(Ctrl__Regs_1__en2), .rb(n952), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 Cause_Reg_reg_18__master ( .q(Cause_Reg_reg_18__m2s), .d(n2660), 
        .sdi(n610), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n953), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 Cause_Reg_reg_18__slave ( .q(Cause_Reg_18), .qb(n609), .d(
        Cause_Reg_reg_18__m2s), .g(Ctrl__Regs_1__en2), .rb(n953), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 Cause_Reg_reg_19__master ( .q(Cause_Reg_reg_19__m2s), .d(n2661), 
        .sdi(n609), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n952), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 Cause_Reg_reg_19__slave ( .q(Cause_Reg_19), .qb(n608), .d(
        Cause_Reg_reg_19__m2s), .g(Ctrl__Regs_1__en2), .rb(n952), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 Cause_Reg_reg_1__master ( .q(Cause_Reg_reg_1__m2s), .d(n2643), 
        .sdi(n627), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n953), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 Cause_Reg_reg_1__slave ( .q(Cause_Reg_1), .qb(n626), .d(
        Cause_Reg_reg_1__m2s), .g(Ctrl__Regs_1__en2), .rb(n953), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 Cause_Reg_reg_20__master ( .q(Cause_Reg_reg_20__m2s), .d(n2662), 
        .sdi(n608), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n952), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 Cause_Reg_reg_20__slave ( .q(Cause_Reg_20), .qb(n607), .d(
        Cause_Reg_reg_20__m2s), .g(Ctrl__Regs_1__en2), .rb(n952), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 Cause_Reg_reg_21__master ( .q(Cause_Reg_reg_21__m2s), .d(n2663), 
        .sdi(n607), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n953), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 Cause_Reg_reg_21__slave ( .q(Cause_Reg_21), .qb(n606), .d(
        Cause_Reg_reg_21__m2s), .g(Ctrl__Regs_1__en2), .rb(n953), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 Cause_Reg_reg_22__master ( .q(Cause_Reg_reg_22__m2s), .d(n2664), 
        .sdi(n606), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n952), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 Cause_Reg_reg_22__slave ( .q(Cause_Reg_22), .qb(n605), .d(
        Cause_Reg_reg_22__m2s), .g(Ctrl__Regs_1__en2), .rb(n952), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 Cause_Reg_reg_23__master ( .q(Cause_Reg_reg_23__m2s), .d(n2665), 
        .sdi(n605), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n953), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 Cause_Reg_reg_23__slave ( .q(Cause_Reg_23), .qb(n604), .d(
        Cause_Reg_reg_23__m2s), .g(Ctrl__Regs_1__en2), .rb(n953), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 Cause_Reg_reg_24__master ( .q(Cause_Reg_reg_24__m2s), .d(n2666), 
        .sdi(n604), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n952), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 Cause_Reg_reg_24__slave ( .q(Cause_Reg_24), .qb(n603), .d(
        Cause_Reg_reg_24__m2s), .g(Ctrl__Regs_1__en2), .rb(n952), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 Cause_Reg_reg_25__master ( .q(Cause_Reg_reg_25__m2s), .d(n2667), 
        .sdi(n603), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n953), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 Cause_Reg_reg_25__slave ( .q(Cause_Reg_25), .qb(n602), .d(
        Cause_Reg_reg_25__m2s), .g(Ctrl__Regs_1__en2), .rb(n953), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 Cause_Reg_reg_26__master ( .q(Cause_Reg_reg_26__m2s), .d(n2668), 
        .sdi(n602), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n952), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 Cause_Reg_reg_26__slave ( .q(Cause_Reg_26), .qb(n601), .d(
        Cause_Reg_reg_26__m2s), .g(Ctrl__Regs_1__en2), .rb(n952), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 Cause_Reg_reg_27__master ( .q(Cause_Reg_reg_27__m2s), .d(n2669), 
        .sdi(n601), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n953), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 Cause_Reg_reg_27__slave ( .q(Cause_Reg_27), .qb(n600), .d(
        Cause_Reg_reg_27__m2s), .g(Ctrl__Regs_1__en2), .rb(n953), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 Cause_Reg_reg_28__master ( .q(Cause_Reg_reg_28__m2s), .d(n2670), 
        .sdi(n600), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n952), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 Cause_Reg_reg_28__slave ( .q(Cause_Reg_28), .qb(n599), .d(
        Cause_Reg_reg_28__m2s), .g(Ctrl__Regs_1__en2), .rb(n952), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 Cause_Reg_reg_29__master ( .q(Cause_Reg_reg_29__m2s), .d(n2671), 
        .sdi(n599), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n954), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 Cause_Reg_reg_29__slave ( .q(Cause_Reg_29), .qb(n598), .d(
        Cause_Reg_reg_29__m2s), .g(Ctrl__Regs_1__en2), .rb(n954), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 Cause_Reg_reg_2__master ( .q(Cause_Reg_reg_2__m2s), .d(n2644), 
        .sdi(n626), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n953), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 Cause_Reg_reg_2__slave ( .q(Cause_Reg_2), .qb(n625), .d(
        Cause_Reg_reg_2__m2s), .g(Ctrl__Regs_1__en2), .rb(n953), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 Cause_Reg_reg_30__master ( .q(Cause_Reg_reg_30__m2s), .d(n2672), 
        .sdi(n598), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n954), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 Cause_Reg_reg_30__slave ( .q(Cause_Reg_30), .qb(n597), .d(
        Cause_Reg_reg_30__m2s), .g(Ctrl__Regs_1__en2), .rb(n954), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 Cause_Reg_reg_31__master ( .q(Cause_Reg_reg_31__m2s), .d(n2673), 
        .sdi(n597), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n952), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 Cause_Reg_reg_31__slave ( .q(Cause_Reg_31), .qb(n596), .d(
        Cause_Reg_reg_31__m2s), .g(Ctrl__Regs_1__en2), .rb(n952), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 Cause_Reg_reg_3__master ( .q(Cause_Reg_reg_3__m2s), .d(n2645), 
        .sdi(n625), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n952), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 Cause_Reg_reg_3__slave ( .q(Cause_Reg_3), .qb(n624), .d(
        Cause_Reg_reg_3__m2s), .g(Ctrl__Regs_1__en2), .rb(n952), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 Cause_Reg_reg_4__master ( .q(Cause_Reg_reg_4__m2s), .d(n2646), 
        .sdi(n624), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n954), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 Cause_Reg_reg_4__slave ( .q(Cause_Reg_4), .qb(n623), .d(
        Cause_Reg_reg_4__m2s), .g(Ctrl__Regs_1__en2), .rb(n954), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 Cause_Reg_reg_5__master ( .q(Cause_Reg_reg_5__m2s), .d(n2647), 
        .sdi(n623), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n952), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 Cause_Reg_reg_5__slave ( .q(Cause_Reg_5), .qb(n622), .d(
        Cause_Reg_reg_5__m2s), .g(Ctrl__Regs_1__en2), .rb(n952), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 Cause_Reg_reg_6__master ( .q(Cause_Reg_reg_6__m2s), .d(n2648), 
        .sdi(n622), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n954), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 Cause_Reg_reg_6__slave ( .q(Cause_Reg_6), .qb(n621), .d(
        Cause_Reg_reg_6__m2s), .g(Ctrl__Regs_1__en2), .rb(n954), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 Cause_Reg_reg_7__master ( .q(Cause_Reg_reg_7__m2s), .d(n2649), 
        .sdi(n621), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n952), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 Cause_Reg_reg_7__slave ( .q(Cause_Reg_7), .qb(n620), .d(
        Cause_Reg_reg_7__m2s), .g(Ctrl__Regs_1__en2), .rb(n952), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 Cause_Reg_reg_8__master ( .q(Cause_Reg_reg_8__m2s), .d(n2650), 
        .sdi(n620), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n954), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 Cause_Reg_reg_8__slave ( .q(Cause_Reg_8), .qb(n619), .d(
        Cause_Reg_reg_8__m2s), .g(Ctrl__Regs_1__en2), .rb(n954), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 Cause_Reg_reg_9__master ( .q(Cause_Reg_reg_9__m2s), .d(n2651), 
        .sdi(n619), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n952), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 Cause_Reg_reg_9__slave ( .q(Cause_Reg_9), .qb(n618), .d(
        Cause_Reg_reg_9__m2s), .g(Ctrl__Regs_1__en2), .rb(n952), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 EPC_reg_0__master ( .q(EPC_reg_0__m2s), .d(n2674), .sdi(n596), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n954), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 EPC_reg_0__slave ( .q(EPC_0), .qb(n595), .d(EPC_reg_0__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n954), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 EPC_reg_10__master ( .q(EPC_reg_10__m2s), .d(n2684), .sdi(EPC_9), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n954), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 EPC_reg_10__slave ( .q(EPC_10), .qb(n593), .d(EPC_reg_10__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n954), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 EPC_reg_11__master ( .q(EPC_reg_11__m2s), .d(n2685), .sdi(EPC_10
        ), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n952), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 EPC_reg_11__slave ( .q(EPC_11), .qb(n592), .d(EPC_reg_11__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n952), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 EPC_reg_12__master ( .q(EPC_reg_12__m2s), .d(n2686), .sdi(EPC_11
        ), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n954), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 EPC_reg_12__slave ( .q(EPC_12), .qb(n591), .d(EPC_reg_12__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n954), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 EPC_reg_13__master ( .q(EPC_reg_13__m2s), .d(n2687), .sdi(EPC_12
        ), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n951), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 EPC_reg_13__slave ( .q(EPC_13), .qb(n590), .d(EPC_reg_13__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n951), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 EPC_reg_14__master ( .q(EPC_reg_14__m2s), .d(n2688), .sdi(EPC_13
        ), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n954), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 EPC_reg_14__slave ( .q(EPC_14), .qb(n589), .d(EPC_reg_14__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n954), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 EPC_reg_15__master ( .q(EPC_reg_15__m2s), .d(n2689), .sdi(EPC_14
        ), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n951), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 EPC_reg_15__slave ( .q(EPC_15), .qb(n588), .d(EPC_reg_15__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n951), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 EPC_reg_16__master ( .q(EPC_reg_16__m2s), .d(n2690), .sdi(n588), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n954), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 EPC_reg_16__slave ( .q(EPC_16), .qb(n587), .d(EPC_reg_16__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n954), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 EPC_reg_17__master ( .q(EPC_reg_17__m2s), .d(n2691), .sdi(EPC_16
        ), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n951), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 EPC_reg_17__slave ( .q(EPC_17), .qb(n586), .d(EPC_reg_17__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n951), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 EPC_reg_18__master ( .q(EPC_reg_18__m2s), .d(n2692), .sdi(EPC_17
        ), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n954), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 EPC_reg_18__slave ( .q(EPC_18), .qb(n585), .d(EPC_reg_18__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n954), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 EPC_reg_19__master ( .q(EPC_reg_19__m2s), .d(n2693), .sdi(EPC_18
        ), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n951), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 EPC_reg_19__slave ( .q(EPC_19), .qb(n584), .d(EPC_reg_19__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n951), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 EPC_reg_1__master ( .q(EPC_reg_1__m2s), .d(n2675), .sdi(EPC_0), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n952), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 EPC_reg_1__slave ( .q(EPC_1), .qb(n594), .d(EPC_reg_1__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n952), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 EPC_reg_20__master ( .q(EPC_reg_20__m2s), .d(n2694), .sdi(EPC_19
        ), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n951), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 EPC_reg_20__slave ( .q(EPC_20), .qb(n583), .d(EPC_reg_20__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n951), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 EPC_reg_21__master ( .q(EPC_reg_21__m2s), .d(n2695), .sdi(EPC_20
        ), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n954), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 EPC_reg_21__slave ( .q(EPC_21), .qb(n4383), .d(EPC_reg_21__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n954), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 EPC_reg_22__master ( .q(EPC_reg_22__m2s), .d(n2696), .sdi(n4383), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n951), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 EPC_reg_22__slave ( .q(EPC_22), .qb(n4382), .d(EPC_reg_22__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n951), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 EPC_reg_23__master ( .q(EPC_reg_23__m2s), .d(n2697), .sdi(n4382), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n954), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 EPC_reg_23__slave ( .q(EPC_23), .qb(n4381), .d(EPC_reg_23__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n954), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 EPC_reg_24__master ( .q(EPC_reg_24__m2s), .d(n2698), .sdi(n4381), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n951), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 EPC_reg_24__slave ( .q(EPC_24), .qb(n4380), .d(EPC_reg_24__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n951), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 EPC_reg_25__master ( .q(EPC_reg_25__m2s), .d(n2699), .sdi(n4380), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n954), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 EPC_reg_25__slave ( .q(EPC_25), .qb(n4379), .d(EPC_reg_25__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n954), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 EPC_reg_26__master ( .q(EPC_reg_26__m2s), .d(n2700), .sdi(n4379), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n951), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 EPC_reg_26__slave ( .q(EPC_26), .qb(n582), .d(EPC_reg_26__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n951), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 EPC_reg_27__master ( .q(EPC_reg_27__m2s), .d(n2701), .sdi(n582), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n955), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 EPC_reg_27__slave ( .q(EPC_27), .qb(n581), .d(EPC_reg_27__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n955), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 EPC_reg_28__master ( .q(EPC_reg_28__m2s), .d(n2702), .sdi(n581), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n951), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 EPC_reg_28__slave ( .q(EPC_28), .qb(n580), .d(EPC_reg_28__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n951), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 EPC_reg_29__master ( .q(EPC_reg_29__m2s), .d(n2703), .sdi(n580), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n955), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 EPC_reg_29__slave ( .q(EPC_29), .qb(n579), .d(EPC_reg_29__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n955), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 EPC_reg_2__master ( .q(EPC_reg_2__m2s), .d(n2676), .sdi(EPC_1), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n954), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 EPC_reg_2__slave ( .q(EPC_2), .qb(n4385), .d(EPC_reg_2__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n954), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 EPC_reg_30__master ( .q(EPC_reg_30__m2s), .d(n2704), .sdi(n579), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n955), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 EPC_reg_30__slave ( .q(EPC_30), .qb(n662), .d(EPC_reg_30__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n955), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 EPC_reg_31__master ( .q(EPC_reg_31__m2s), .d(
        _EPC_reg_31_net69891), .sdi(EPC_30), .se(test_se), .g(
        Ctrl__Regs_1__en1), .rb(n951), .glob_g(global_g1), .sync_sel(sync_sel)
         );
    mlatnr_2 EPC_reg_31__slave ( .q(EPC_31), .qb(n578), .d(EPC_reg_31__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n951), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 EPC_reg_3__master ( .q(EPC_reg_3__m2s), .d(n2677), .sdi(n4385), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n951), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 EPC_reg_3__slave ( .q(EPC_3), .qb(n4384), .d(EPC_reg_3__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n951), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 EPC_reg_4__master ( .q(EPC_reg_4__m2s), .d(n2678), .sdi(n4384), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n955), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 EPC_reg_4__slave ( .q(EPC_4), .qb(n577), .d(EPC_reg_4__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n955), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 EPC_reg_5__master ( .q(EPC_reg_5__m2s), .d(n2679), .sdi(EPC_4), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n951), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 EPC_reg_5__slave ( .q(EPC_5), .qb(n576), .d(EPC_reg_5__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n951), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 EPC_reg_6__master ( .q(EPC_reg_6__m2s), .d(n2680), .sdi(EPC_5), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n955), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 EPC_reg_6__slave ( .q(EPC_6), .qb(n575), .d(EPC_reg_6__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n955), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 EPC_reg_7__master ( .q(EPC_reg_7__m2s), .d(n2681), .sdi(EPC_6), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n951), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 EPC_reg_7__slave ( .q(EPC_7), .qb(n574), .d(EPC_reg_7__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n951), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 EPC_reg_8__master ( .q(EPC_reg_8__m2s), .d(n2682), .sdi(EPC_7), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n955), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 EPC_reg_8__slave ( .q(EPC_8), .qb(n573), .d(EPC_reg_8__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n955), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 EPC_reg_9__master ( .q(EPC_reg_9__m2s), .d(n2683), .sdi(EPC_8), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n951), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 EPC_reg_9__slave ( .q(EPC_9), .qb(n572), .d(EPC_reg_9__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n951), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 IR_function_field_reg_0__master ( .q(
        IR_function_field_reg_0__m2s), .d(n3764), .sdi(EPC_31), .se(test_se), 
        .g(Ctrl__Regs_1__en1), .rb(n955), .glob_g(global_g1), .sync_sel(
        sync_sel) );
    mlatnr_2 IR_function_field_reg_0__slave ( .q(IR_function_field[0]), .qb(
        n1859), .d(IR_function_field_reg_0__m2s), .g(Ctrl__Regs_1__en2), .rb(
        n955), .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_function_field_reg_1__master ( .q(
        IR_function_field_reg_1__m2s), .d(n3765), .sdi(n1859), .se(test_se), 
        .g(Ctrl__Regs_1__en1), .rb(n951), .glob_g(global_g1), .sync_sel(
        sync_sel) );
    mlatnr_2 IR_function_field_reg_1__slave ( .q(IR_function_field[1]), .qb(
        n1860), .d(IR_function_field_reg_1__m2s), .g(Ctrl__Regs_1__en2), .rb(
        n951), .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_function_field_reg_2__master ( .q(
        IR_function_field_reg_2__m2s), .d(n3766), .sdi(n1860), .se(test_se), 
        .g(Ctrl__Regs_1__en1), .rb(n955), .glob_g(global_g1), .sync_sel(
        sync_sel) );
    mlatnr_2 IR_function_field_reg_2__slave ( .q(IR_function_field[2]), .qb(
        n1861), .d(IR_function_field_reg_2__m2s), .g(Ctrl__Regs_1__en2), .rb(
        n955), .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_function_field_reg_3__master ( .q(
        IR_function_field_reg_3__m2s), .d(n3767), .sdi(n1861), .se(test_se), 
        .g(Ctrl__Regs_1__en1), .rb(n950), .glob_g(global_g1), .sync_sel(
        sync_sel) );
    mlatnr_2 IR_function_field_reg_3__slave ( .q(IR_function_field[3]), .qb(
        n1862), .d(IR_function_field_reg_3__m2s), .g(Ctrl__Regs_1__en2), .rb(
        n950), .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_function_field_reg_4__master ( .q(
        IR_function_field_reg_4__m2s), .d(n3768), .sdi(n1862), .se(test_se), 
        .g(Ctrl__Regs_1__en1), .rb(n955), .glob_g(global_g1), .sync_sel(
        sync_sel) );
    mlatnr_2 IR_function_field_reg_4__slave ( .q(IR_function_field[4]), .qb(
        n1863), .d(IR_function_field_reg_4__m2s), .g(Ctrl__Regs_1__en2), .rb(
        n955), .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_function_field_reg_5__master ( .q(
        IR_function_field_reg_5__m2s), .d(n3769), .sdi(n1863), .se(test_se), 
        .g(Ctrl__Regs_1__en1), .rb(n950), .glob_g(global_g1), .sync_sel(
        sync_sel) );
    mlatnr_2 IR_function_field_reg_5__slave ( .q(IR_function_field[5]), .qb(
        n4378), .d(IR_function_field_reg_5__m2s), .g(Ctrl__Regs_1__en2), .rb(
        n950), .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_opcode_field_reg_0__master ( .q(IR_opcode_field_reg_0__m2s), 
        .d(n3770), .sdi(n4378), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n911), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_4 IR_opcode_field_reg_0__slave ( .q(n4454), .qb(n4377), .d(
        IR_opcode_field_reg_0__m2s), .g(Ctrl__Regs_1__en2), .rb(n911), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_opcode_field_reg_1__master ( .q(IR_opcode_field_reg_1__m2s), 
        .d(n3771), .sdi(n4377), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n911), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_4 IR_opcode_field_reg_1__slave ( .q(n4453), .qb(n4376), .d(
        IR_opcode_field_reg_1__m2s), .g(Ctrl__Regs_1__en2), .rb(n911), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_opcode_field_reg_2__master ( .q(IR_opcode_field_reg_2__m2s), 
        .d(n3772), .sdi(n4376), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n955), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_4 IR_opcode_field_reg_2__slave ( .q(n4452), .qb(n4375), .d(
        IR_opcode_field_reg_2__m2s), .g(Ctrl__Regs_1__en2), .rb(n955), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_opcode_field_reg_3__master ( .q(IR_opcode_field_reg_3__m2s), 
        .d(n3773), .sdi(n4375), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_4 IR_opcode_field_reg_3__slave ( .q(IR_opcode_field[3]), .qb(n4374), 
        .d(IR_opcode_field_reg_3__m2s), .g(Ctrl__Regs_1__en2), .rb(n950), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_opcode_field_reg_4__master ( .q(IR_opcode_field_reg_4__m2s), 
        .d(n3774), .sdi(n4374), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n955), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_4 IR_opcode_field_reg_4__slave ( .q(IR_opcode_field[4]), .qb(n4373), 
        .d(IR_opcode_field_reg_4__m2s), .g(Ctrl__Regs_1__en2), .rb(n955), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_opcode_field_reg_5__master ( .q(IR_opcode_field_reg_5__m2s), 
        .d(n3775), .sdi(n4373), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_4 IR_opcode_field_reg_5__slave ( .q(IR_opcode_field[5]), .qb(n4372), 
        .d(IR_opcode_field_reg_5__m2s), .g(Ctrl__Regs_1__en2), .rb(n950), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_1 Imm_reg_0__master ( .q(Imm_reg_0__m2s), .d(n3791), .sdi(n4372), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n914), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 Imm_reg_0__slave ( .q(N6328), .qb(n813), .d(Imm_reg_0__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n914), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 Imm_reg_10__master ( .q(Imm_reg_10__m2s), .d(n3801), .sdi(n873), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n914), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_4 Imm_reg_10__slave ( .q(N6348), .qb(n4371), .d(Imm_reg_10__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n914), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 Imm_reg_11__master ( .q(Imm_reg_11__m2s), .d(n3802), .sdi(n4371), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 Imm_reg_11__slave ( .q(N6350), .qb(n786), .d(Imm_reg_11__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 Imm_reg_12__master ( .q(Imm_reg_12__m2s), .d(n3803), .sdi(n786), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_4 Imm_reg_12__slave ( .q(N6352), .qb(n779), .d(Imm_reg_12__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 Imm_reg_13__master ( .q(Imm_reg_13__m2s), .d(n3804), .sdi(n779), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n916), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_4 Imm_reg_13__slave ( .q(N6354), .qb(n4370), .d(Imm_reg_13__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n916), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 Imm_reg_14__master ( .q(Imm_reg_14__m2s), .d(n3805), .sdi(n4370), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_4 Imm_reg_14__slave ( .q(N6356), .qb(n647), .d(Imm_reg_14__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 Imm_reg_15__master ( .q(Imm_reg_15__m2s), .d(n3806), .sdi(n647), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_4 Imm_reg_15__slave ( .q(N6358), .qb(n829), .d(Imm_reg_15__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 Imm_reg_16__master ( .q(Imm_reg_16__m2s), .d(n3807), .sdi(n829), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n911), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_4 Imm_reg_16__slave ( .q(N6360), .qb(n648), .d(Imm_reg_16__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n911), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 Imm_reg_17__master ( .q(Imm_reg_17__m2s), .d(n3808), .sdi(n648), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_4 Imm_reg_17__slave ( .q(N6362), .qb(n803), .d(Imm_reg_17__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 Imm_reg_18__master ( .q(Imm_reg_18__m2s), .d(n3809), .sdi(n803), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_4 Imm_reg_18__slave ( .q(N6364), .qb(n778), .d(Imm_reg_18__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 Imm_reg_19__master ( .q(Imm_reg_19__m2s), .d(n3810), .sdi(n778), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n911), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 Imm_reg_19__slave ( .q(N6366), .qb(n775), .d(Imm_reg_19__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n911), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 Imm_reg_1__master ( .q(Imm_reg_1__m2s), .d(n3792), .sdi(n813), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n915), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_4 Imm_reg_1__slave ( .q(Imm[1]), .qb(n720), .d(Imm_reg_1__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n915), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 Imm_reg_20__master ( .q(Imm_reg_20__m2s), .d(n3811), .sdi(n775), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n911), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 Imm_reg_20__slave ( .q(N6368), .qb(n732), .d(Imm_reg_20__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n911), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 Imm_reg_21__master ( .q(Imm_reg_21__m2s), .d(n3812), .sdi(n732), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 Imm_reg_21__slave ( .q(N6370), .qb(n649), .d(Imm_reg_21__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 Imm_reg_22__master ( .q(Imm_reg_22__m2s), .d(n3813), .sdi(n649), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n911), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_4 Imm_reg_22__slave ( .q(Imm[22]), .qb(n789), .d(Imm_reg_22__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n911), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 Imm_reg_23__master ( .q(Imm_reg_23__m2s), .d(n3814), .sdi(n789), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n912), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 Imm_reg_23__slave ( .q(Imm[23]), .qb(n827), .d(Imm_reg_23__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n912), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 Imm_reg_24__master ( .q(Imm_reg_24__m2s), .d(n3815), .sdi(n827), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n911), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 Imm_reg_24__slave ( .q(N6376), .qb(n654), .d(Imm_reg_24__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n911), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 Imm_reg_25__master ( .q(Imm_reg_25__m2s), .d(n3816), .sdi(n654), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n951), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 Imm_reg_25__slave ( .q(Imm[25]), .qb(n816), .d(Imm_reg_25__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n951), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 Imm_reg_26__master ( .q(Imm_reg_26__m2s), .d(n3817), .sdi(n816), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n912), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 Imm_reg_26__slave ( .q(N6380), .qb(n735), .d(Imm_reg_26__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n912), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 Imm_reg_27__master ( .q(Imm_reg_27__m2s), .d(n3818), .sdi(n735), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 Imm_reg_27__slave ( .q(N6382), .qb(n765), .d(Imm_reg_27__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 Imm_reg_28__master ( .q(Imm_reg_28__m2s), .d(n3819), .sdi(n765), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 Imm_reg_28__slave ( .q(N6384), .qb(n696), .d(Imm_reg_28__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 Imm_reg_29__master ( .q(Imm_reg_29__m2s), .d(n3820), .sdi(n696), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n914), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 Imm_reg_29__slave ( .q(N6386), .qb(n762), .d(Imm_reg_29__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n914), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 Imm_reg_2__master ( .q(Imm_reg_2__m2s), .d(n3793), .sdi(n720), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n914), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 Imm_reg_2__slave ( .q(N6332), .qb(n870), .d(Imm_reg_2__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n914), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 Imm_reg_30__master ( .q(Imm_reg_30__m2s), .d(n3821), .sdi(n762), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n914), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 Imm_reg_30__slave ( .q(N6388), .qb(n701), .d(Imm_reg_30__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n914), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 Imm_reg_31__master ( .q(Imm_reg_31__m2s), .d(n3822), .sdi(n701), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n911), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_4 Imm_reg_31__slave ( .q(N6390), .qb(n4369), .d(Imm_reg_31__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n911), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 Imm_reg_3__master ( .q(Imm_reg_3__m2s), .d(n3794), .sdi(n870), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n914), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_4 Imm_reg_3__slave ( .q(N6334), .qb(n886), .d(Imm_reg_3__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n914), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 Imm_reg_4__master ( .q(Imm_reg_4__m2s), .d(n3795), .sdi(n886), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_4 Imm_reg_4__slave ( .q(N6336), .qb(n871), .d(Imm_reg_4__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n949), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 Imm_reg_5__master ( .q(Imm_reg_5__m2s), .d(n3796), .sdi(n871), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n914), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_4 Imm_reg_5__slave ( .q(N6338), .qb(n845), .d(Imm_reg_5__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n914), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 Imm_reg_6__master ( .q(Imm_reg_6__m2s), .d(n3797), .sdi(n845), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n914), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_4 Imm_reg_6__slave ( .q(N6340), .qb(n643), .d(Imm_reg_6__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n914), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 Imm_reg_7__master ( .q(Imm_reg_7__m2s), .d(n3798), .sdi(n643), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n914), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_4 Imm_reg_7__slave ( .q(N6342), .qb(n734), .d(Imm_reg_7__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n914), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 Imm_reg_8__master ( .q(Imm_reg_8__m2s), .d(n3799), .sdi(n734), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n911), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_4 Imm_reg_8__slave ( .q(N6344), .qb(n872), .d(Imm_reg_8__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n911), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 Imm_reg_9__master ( .q(Imm_reg_9__m2s), .d(n3800), .sdi(n872), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 Imm_reg_9__slave ( .q(N6346), .qb(n873), .d(Imm_reg_9__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n949), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    inv_2 U10 ( .x(n554), .a(n1547) );
    inv_2 U100 ( .x(n1382), .a(N449) );
    or2_2 U1000 ( .x(n1767), .a(n3936), .b(n3940) );
    mux2_2 U1001 ( .x(n3285), .d0(_RegFile_13__0), .sl(n1830), .d1(WB_data[0])
         );
    mux2_2 U1002 ( .x(n3286), .d0(_RegFile_13__1), .sl(n1830), .d1(WB_data[1])
         );
    mux2_2 U1003 ( .x(n3287), .d0(_RegFile_13__2), .sl(n1830), .d1(WB_data[2])
         );
    mux2_2 U1004 ( .x(n3288), .d0(_RegFile_13__3), .sl(n1830), .d1(WB_data[3])
         );
    mux2_2 U1005 ( .x(n3289), .d0(_RegFile_13__4), .sl(n1830), .d1(WB_data[4])
         );
    mux2_2 U1006 ( .x(n3290), .d0(_RegFile_13__5), .sl(n1830), .d1(WB_data[5])
         );
    mux2_2 U1007 ( .x(n3291), .d0(_RegFile_13__6), .sl(n1830), .d1(WB_data[6])
         );
    mux2_2 U1008 ( .x(n3292), .d0(_RegFile_13__7), .sl(n1830), .d1(WB_data[7])
         );
    mux2i_1 U1009 ( .x(n3294), .d0(n1983), .sl(n1830), .d1(n1801) );
    inv_2 U101 ( .x(n1399), .a(N456) );
    mux2i_1 U1010 ( .x(n3295), .d0(n1960), .sl(n1830), .d1(n1778) );
    mux2i_1 U1011 ( .x(n3296), .d0(n1961), .sl(n1830), .d1(n1779) );
    mux2i_1 U1012 ( .x(n3297), .d0(n1962), .sl(n1830), .d1(n1780) );
    mux2i_1 U1013 ( .x(n3298), .d0(n1963), .sl(n1830), .d1(n1781) );
    mux2i_1 U1014 ( .x(n3299), .d0(n1964), .sl(n1830), .d1(n1782) );
    mux2i_1 U1015 ( .x(n3300), .d0(n1965), .sl(n1830), .d1(n1783) );
    mux2i_1 U1016 ( .x(n3301), .d0(n1966), .sl(n1830), .d1(n1784) );
    mux2i_1 U1017 ( .x(n3302), .d0(n1967), .sl(n1830), .d1(n1785) );
    mux2i_1 U1018 ( .x(n3303), .d0(n1968), .sl(n1830), .d1(n1786) );
    mux2i_1 U1019 ( .x(n3304), .d0(n1969), .sl(n1830), .d1(n1787) );
    nand2i_2 U102 ( .x(n1520), .a(n1515), .b(n1521) );
    mux2i_1 U1020 ( .x(n3305), .d0(n1970), .sl(n1830), .d1(n1788) );
    mux2i_1 U1021 ( .x(n3306), .d0(n1971), .sl(n1830), .d1(n1789) );
    mux2i_1 U1022 ( .x(n3307), .d0(n1972), .sl(n1830), .d1(n1790) );
    mux2i_1 U1023 ( .x(n3308), .d0(n1973), .sl(n1830), .d1(n1791) );
    mux2i_1 U1024 ( .x(n3309), .d0(n1974), .sl(n1830), .d1(n1792) );
    mux2i_1 U1025 ( .x(n3310), .d0(n1975), .sl(n1830), .d1(n1793) );
    mux2i_1 U1026 ( .x(n3311), .d0(n1976), .sl(n1830), .d1(n1794) );
    mux2i_1 U1027 ( .x(n3312), .d0(n1977), .sl(n1830), .d1(n1795) );
    mux2i_1 U1028 ( .x(n3313), .d0(n1978), .sl(n1830), .d1(n1796) );
    mux2i_1 U1029 ( .x(n3314), .d0(n1979), .sl(n1830), .d1(n1797) );
    nand2i_2 U103 ( .x(n1518), .a(n1515), .b(n1519) );
    mux2i_1 U1030 ( .x(n3315), .d0(n1980), .sl(n1830), .d1(n1798) );
    or2_2 U1031 ( .x(n1768), .a(n3935), .b(n3940) );
    mux2_2 U1032 ( .x(n3317), .d0(_RegFile_12__0), .sl(n1829), .d1(WB_data[0])
         );
    mux2_2 U1033 ( .x(n3318), .d0(_RegFile_12__1), .sl(n1829), .d1(WB_data[1])
         );
    mux2_2 U1034 ( .x(n3319), .d0(_RegFile_12__2), .sl(n1829), .d1(WB_data[2])
         );
    mux2_2 U1035 ( .x(n3320), .d0(_RegFile_12__3), .sl(n1829), .d1(WB_data[3])
         );
    mux2_2 U1036 ( .x(n3321), .d0(_RegFile_12__4), .sl(n1829), .d1(WB_data[4])
         );
    mux2_2 U1037 ( .x(n3322), .d0(_RegFile_12__5), .sl(n1829), .d1(WB_data[5])
         );
    mux2_2 U1038 ( .x(n3323), .d0(_RegFile_12__6), .sl(n1829), .d1(WB_data[6])
         );
    mux2_2 U1039 ( .x(n3324), .d0(_RegFile_12__7), .sl(n1829), .d1(WB_data[7])
         );
    and4i_3 U104 ( .x(n796), .a(n795), .b(___cell__36997_net129977), .c(
        ___cell__36997_net129979), .d(___cell__36997_net130187) );
    mux2i_1 U1040 ( .x(n3326), .d0(n1959), .sl(n1829), .d1(n1801) );
    mux2i_1 U1041 ( .x(n3327), .d0(n1936), .sl(n1829), .d1(n1778) );
    mux2i_1 U1042 ( .x(n3328), .d0(n1937), .sl(n1829), .d1(n1779) );
    mux2i_1 U1043 ( .x(n3329), .d0(n1938), .sl(n1829), .d1(n1780) );
    mux2i_1 U1044 ( .x(n3330), .d0(n1939), .sl(n1829), .d1(n1781) );
    mux2i_1 U1045 ( .x(n3331), .d0(n1940), .sl(n1829), .d1(n1782) );
    mux2i_1 U1046 ( .x(n3332), .d0(n1941), .sl(n1829), .d1(n1783) );
    mux2i_1 U1047 ( .x(n3333), .d0(n1942), .sl(n1829), .d1(n1784) );
    mux2i_1 U1048 ( .x(n3334), .d0(n1943), .sl(n1829), .d1(n1785) );
    mux2i_1 U1049 ( .x(n3335), .d0(n1944), .sl(n1829), .d1(n1786) );
    inv_2 U105 ( .x(n694), .a(n693) );
    mux2i_1 U1050 ( .x(n3336), .d0(n1945), .sl(n1829), .d1(n1787) );
    mux2i_1 U1051 ( .x(n3337), .d0(n1946), .sl(n1829), .d1(n1788) );
    mux2i_1 U1052 ( .x(n3338), .d0(n1947), .sl(n1829), .d1(n1789) );
    mux2i_1 U1053 ( .x(n3339), .d0(n1948), .sl(n1829), .d1(n1790) );
    mux2i_1 U1054 ( .x(n3340), .d0(n1949), .sl(n1829), .d1(n1791) );
    mux2i_1 U1055 ( .x(n3341), .d0(n1950), .sl(n1829), .d1(n1792) );
    mux2i_1 U1056 ( .x(n3342), .d0(n1951), .sl(n1829), .d1(n1793) );
    mux2i_1 U1057 ( .x(n3343), .d0(n1952), .sl(n1829), .d1(n1794) );
    mux2i_1 U1058 ( .x(n3344), .d0(n1953), .sl(n1829), .d1(n1795) );
    mux2i_1 U1059 ( .x(n3345), .d0(n1954), .sl(n1829), .d1(n1796) );
    inv_5 U106 ( .x(n704), .a(___cell__36997_net126612) );
    mux2i_1 U1060 ( .x(n3346), .d0(n1955), .sl(n1829), .d1(n1797) );
    buf_3 U1061 ( .x(n959), .a(n957) );
    mux2i_1 U1062 ( .x(n3347), .d0(n1956), .sl(n1829), .d1(n1798) );
    buf_3 U1063 ( .x(n946), .a(n939) );
    or2_2 U1064 ( .x(n1769), .a(n3927), .b(n3940) );
    mux2_2 U1065 ( .x(n3349), .d0(_RegFile_11__0), .sl(n1828), .d1(WB_data[0])
         );
    mux2_2 U1066 ( .x(n3350), .d0(_RegFile_11__1), .sl(n1828), .d1(WB_data[1])
         );
    mux2_2 U1067 ( .x(n3351), .d0(_RegFile_11__2), .sl(n1828), .d1(WB_data[2])
         );
    mux2_2 U1068 ( .x(n3352), .d0(_RegFile_11__3), .sl(n1828), .d1(WB_data[3])
         );
    mux2_2 U1069 ( .x(n3353), .d0(_RegFile_11__4), .sl(n1828), .d1(WB_data[4])
         );
    nor2i_1 U107 ( .x(n1262), .a(___cell__36997_net126612), .b(n1263) );
    mux2_2 U1070 ( .x(n3354), .d0(_RegFile_11__5), .sl(n1828), .d1(WB_data[5])
         );
    mux2_2 U1071 ( .x(n3355), .d0(_RegFile_11__6), .sl(n1828), .d1(WB_data[6])
         );
    mux2_2 U1072 ( .x(n3356), .d0(_RegFile_11__7), .sl(n1828), .d1(WB_data[7])
         );
    mux2i_1 U1073 ( .x(n3358), .d0(n1935), .sl(n1828), .d1(n1801) );
    mux2i_1 U1074 ( .x(n3359), .d0(n1912), .sl(n1828), .d1(n1778) );
    mux2i_1 U1075 ( .x(n3360), .d0(n1913), .sl(n1828), .d1(n1779) );
    mux2i_1 U1076 ( .x(n3361), .d0(n1914), .sl(n1828), .d1(n1780) );
    mux2i_1 U1077 ( .x(n3362), .d0(n1915), .sl(n1828), .d1(n1781) );
    mux2i_1 U1078 ( .x(n3363), .d0(n1916), .sl(n1828), .d1(n1782) );
    mux2i_1 U1079 ( .x(n3364), .d0(n1917), .sl(n1828), .d1(n1783) );
    oai211_1 U108 ( .x(n1261), .a(n1314), .b(n883), .c(FREEZE), .d(n564) );
    mux2i_1 U1080 ( .x(n3365), .d0(n1918), .sl(n1828), .d1(n1784) );
    mux2i_1 U1081 ( .x(n3366), .d0(n1919), .sl(n1828), .d1(n1785) );
    mux2i_1 U1082 ( .x(n3367), .d0(n1920), .sl(n1828), .d1(n1786) );
    mux2i_1 U1083 ( .x(n3368), .d0(n1921), .sl(n1828), .d1(n1787) );
    mux2i_1 U1084 ( .x(n3369), .d0(n1922), .sl(n1828), .d1(n1788) );
    mux2i_1 U1085 ( .x(n3370), .d0(n1923), .sl(n1828), .d1(n1789) );
    mux2i_1 U1086 ( .x(n3371), .d0(n1924), .sl(n1828), .d1(n1790) );
    mux2i_1 U1087 ( .x(n3372), .d0(n1925), .sl(n1828), .d1(n1791) );
    mux2i_1 U1088 ( .x(n3373), .d0(n1926), .sl(n1828), .d1(n1792) );
    mux2i_1 U1089 ( .x(n3374), .d0(n1927), .sl(n1828), .d1(n1793) );
    nand3_1 U109 ( .x(n3944), .a(WB_index_0), .b(WB_index_4), .c(WB_index_1)
         );
    mux2i_1 U1090 ( .x(n3375), .d0(n1928), .sl(n1828), .d1(n1794) );
    mux2i_1 U1091 ( .x(n3376), .d0(n1929), .sl(n1828), .d1(n1795) );
    mux2i_1 U1092 ( .x(n3377), .d0(n1930), .sl(n1828), .d1(n1796) );
    mux2i_1 U1093 ( .x(n3378), .d0(n1931), .sl(n1828), .d1(n1797) );
    buf_3 U1094 ( .x(n958), .a(n945) );
    mux2i_1 U1095 ( .x(n3379), .d0(n1932), .sl(n1828), .d1(n1798) );
    or2_2 U1096 ( .x(n1770), .a(n3937), .b(n3939) );
    mux2_2 U1097 ( .x(n3381), .d0(_RegFile_10__0), .sl(n1827), .d1(WB_data[0])
         );
    mux2_2 U1098 ( .x(n3382), .d0(_RegFile_10__1), .sl(n1827), .d1(WB_data[1])
         );
    mux2_2 U1099 ( .x(n3383), .d0(_RegFile_10__2), .sl(n1827), .d1(WB_data[2])
         );
    buf_3 U11 ( .x(reg_out_A[23]), .a(n3958) );
    nand3_1 U110 ( .x(n3943), .a(WB_index_4), .b(n3928), .c(WB_index_1) );
    mux2_2 U1100 ( .x(n3384), .d0(_RegFile_10__3), .sl(n1827), .d1(WB_data[3])
         );
    mux2_2 U1101 ( .x(n3385), .d0(_RegFile_10__4), .sl(n1827), .d1(WB_data[4])
         );
    mux2_2 U1102 ( .x(n3386), .d0(_RegFile_10__5), .sl(n1827), .d1(WB_data[5])
         );
    mux2_2 U1103 ( .x(n3387), .d0(_RegFile_10__6), .sl(n1827), .d1(WB_data[6])
         );
    mux2_2 U1104 ( .x(n3388), .d0(_RegFile_10__7), .sl(n1827), .d1(WB_data[7])
         );
    mux2i_1 U1105 ( .x(n3390), .d0(n1911), .sl(n1827), .d1(n1801) );
    mux2i_1 U1106 ( .x(n3391), .d0(n1888), .sl(n1827), .d1(n1778) );
    mux2i_1 U1107 ( .x(n3392), .d0(n1889), .sl(n1827), .d1(n1779) );
    mux2i_1 U1108 ( .x(n3393), .d0(n1890), .sl(n1827), .d1(n1780) );
    mux2i_1 U1109 ( .x(n3394), .d0(n1891), .sl(n1827), .d1(n1781) );
    nand3_1 U111 ( .x(n3942), .a(WB_index_4), .b(n3929), .c(WB_index_0) );
    mux2i_1 U1110 ( .x(n3395), .d0(n1892), .sl(n1827), .d1(n1782) );
    mux2i_1 U1111 ( .x(n3396), .d0(n1893), .sl(n1827), .d1(n1783) );
    mux2i_1 U1112 ( .x(n3397), .d0(n1894), .sl(n1827), .d1(n1784) );
    mux2i_1 U1113 ( .x(n3398), .d0(n1895), .sl(n1827), .d1(n1785) );
    mux2i_1 U1114 ( .x(n3399), .d0(n1896), .sl(n1827), .d1(n1786) );
    mux2i_1 U1115 ( .x(n3400), .d0(n1897), .sl(n1827), .d1(n1787) );
    mux2i_1 U1116 ( .x(n3401), .d0(n1898), .sl(n1827), .d1(n1788) );
    mux2i_1 U1117 ( .x(n3402), .d0(n1899), .sl(n1827), .d1(n1789) );
    mux2i_1 U1118 ( .x(n3403), .d0(n1900), .sl(n1827), .d1(n1790) );
    mux2i_1 U1119 ( .x(n3404), .d0(n1901), .sl(n1827), .d1(n1791) );
    nand3_1 U112 ( .x(n3941), .a(n3929), .b(n3928), .c(WB_index_4) );
    mux2i_1 U1120 ( .x(n3405), .d0(n1902), .sl(n1827), .d1(n1792) );
    mux2i_1 U1121 ( .x(n3406), .d0(n1903), .sl(n1827), .d1(n1793) );
    mux2i_1 U1122 ( .x(n3407), .d0(n1904), .sl(n1827), .d1(n1794) );
    mux2i_1 U1123 ( .x(n3408), .d0(n1905), .sl(n1827), .d1(n1795) );
    mux2i_1 U1124 ( .x(n3409), .d0(n1906), .sl(n1827), .d1(n1796) );
    mux2i_1 U1125 ( .x(n3410), .d0(n1907), .sl(n1827), .d1(n1797) );
    mux2i_1 U1126 ( .x(n3411), .d0(n1908), .sl(n1827), .d1(n1798) );
    or2_2 U1127 ( .x(n1771), .a(n3936), .b(n3939) );
    mux2_2 U1128 ( .x(n3413), .d0(_RegFile_9__0), .sl(n1857), .d1(WB_data[0])
         );
    mux2_2 U1129 ( .x(n3414), .d0(_RegFile_9__1), .sl(n1857), .d1(WB_data[1])
         );
    nand3_1 U113 ( .x(n3940), .a(WB_index_2), .b(WB_index_3), .c(reg_write_WB)
         );
    mux2_2 U1130 ( .x(n3415), .d0(_RegFile_9__2), .sl(n1857), .d1(WB_data[2])
         );
    mux2_2 U1131 ( .x(n3416), .d0(_RegFile_9__3), .sl(n1857), .d1(WB_data[3])
         );
    mux2_2 U1132 ( .x(n3417), .d0(_RegFile_9__4), .sl(n1857), .d1(WB_data[4])
         );
    mux2_2 U1133 ( .x(n3418), .d0(_RegFile_9__5), .sl(n1857), .d1(WB_data[5])
         );
    mux2_2 U1134 ( .x(n3419), .d0(_RegFile_9__6), .sl(n1857), .d1(n691) );
    mux2_2 U1135 ( .x(n3420), .d0(_RegFile_9__7), .sl(n1857), .d1(n692) );
    mux2i_1 U1136 ( .x(n3422), .d0(n2631), .sl(n1857), .d1(n1801) );
    mux2i_1 U1137 ( .x(n3423), .d0(n2608), .sl(n1857), .d1(n1778) );
    mux2i_1 U1138 ( .x(n3424), .d0(n2609), .sl(n1857), .d1(n1779) );
    mux2i_1 U1139 ( .x(n3425), .d0(n2610), .sl(n1857), .d1(n1780) );
    nand3_1 U114 ( .x(n3939), .a(reg_write_WB), .b(n3925), .c(WB_index_3) );
    mux2i_1 U1140 ( .x(n3426), .d0(n2611), .sl(n1857), .d1(n1781) );
    mux2i_1 U1141 ( .x(n3427), .d0(n2612), .sl(n1857), .d1(n1782) );
    mux2i_1 U1142 ( .x(n3428), .d0(n2613), .sl(n1857), .d1(n1783) );
    mux2i_1 U1143 ( .x(n3429), .d0(n2614), .sl(n1857), .d1(n1784) );
    mux2i_1 U1144 ( .x(n3430), .d0(n2615), .sl(n1857), .d1(n1785) );
    mux2i_1 U1145 ( .x(n3431), .d0(n2616), .sl(n1857), .d1(n1786) );
    mux2i_1 U1146 ( .x(n3432), .d0(n2617), .sl(n1857), .d1(n1787) );
    mux2i_1 U1147 ( .x(n3433), .d0(n2618), .sl(n1857), .d1(n1788) );
    mux2i_1 U1148 ( .x(n3434), .d0(n2619), .sl(n1857), .d1(n1789) );
    mux2i_1 U1149 ( .x(n3435), .d0(n2620), .sl(n1857), .d1(n1790) );
    nand3_1 U115 ( .x(n3938), .a(reg_write_WB), .b(n3926), .c(WB_index_2) );
    mux2i_1 U1150 ( .x(n3436), .d0(n2621), .sl(n1857), .d1(n1791) );
    mux2i_1 U1151 ( .x(n3437), .d0(n2622), .sl(n1857), .d1(n1792) );
    mux2i_1 U1152 ( .x(n3438), .d0(n2623), .sl(n1857), .d1(n1793) );
    mux2i_1 U1153 ( .x(n3439), .d0(n2624), .sl(n1857), .d1(n1794) );
    mux2i_1 U1154 ( .x(n3440), .d0(n2625), .sl(n1857), .d1(n1795) );
    mux2i_1 U1155 ( .x(n3441), .d0(n2626), .sl(n1857), .d1(n1796) );
    mux2i_1 U1156 ( .x(n3442), .d0(n2627), .sl(n1857), .d1(n1797) );
    mux2i_1 U1157 ( .x(n3443), .d0(n2628), .sl(n1857), .d1(n1798) );
    or2_2 U1158 ( .x(n1741), .a(n3935), .b(n3939) );
    mux2_2 U1159 ( .x(n3445), .d0(_RegFile_8__0), .sl(n1856), .d1(WB_data[0])
         );
    nand3_1 U116 ( .x(n3937), .a(WB_index_0), .b(___cell__6171_net27367), .c(
        WB_index_1) );
    mux2_2 U1160 ( .x(n3446), .d0(_RegFile_8__1), .sl(n1856), .d1(WB_data[1])
         );
    mux2_2 U1161 ( .x(n3447), .d0(_RegFile_8__2), .sl(n1856), .d1(WB_data[2])
         );
    mux2_2 U1162 ( .x(n3448), .d0(_RegFile_8__3), .sl(n1856), .d1(WB_data[3])
         );
    mux2_2 U1163 ( .x(n3449), .d0(_RegFile_8__4), .sl(n1856), .d1(WB_data[4])
         );
    mux2_2 U1164 ( .x(n3450), .d0(_RegFile_8__5), .sl(n1856), .d1(WB_data[5])
         );
    mux2_2 U1165 ( .x(n3451), .d0(_RegFile_8__6), .sl(n1856), .d1(n691) );
    mux2_2 U1166 ( .x(n3452), .d0(_RegFile_8__7), .sl(n1856), .d1(WB_data[7])
         );
    mux2i_1 U1167 ( .x(n3454), .d0(n2607), .sl(n1856), .d1(n1801) );
    mux2i_1 U1168 ( .x(n3455), .d0(n2584), .sl(n1856), .d1(n1778) );
    mux2i_1 U1169 ( .x(n3456), .d0(n2585), .sl(n1856), .d1(n1779) );
    nand3_1 U117 ( .x(n3936), .a(___cell__6171_net27367), .b(n3928), .c(
        WB_index_1) );
    mux2i_1 U1170 ( .x(n3457), .d0(n2586), .sl(n1856), .d1(n1780) );
    mux2i_1 U1171 ( .x(n3458), .d0(n2587), .sl(n1856), .d1(n1781) );
    mux2i_1 U1172 ( .x(n3459), .d0(n2588), .sl(n1856), .d1(n1782) );
    mux2i_1 U1173 ( .x(n3460), .d0(n2589), .sl(n1856), .d1(n1783) );
    mux2i_1 U1174 ( .x(n3461), .d0(n2590), .sl(n1856), .d1(n1784) );
    mux2i_1 U1175 ( .x(n3462), .d0(n2591), .sl(n1856), .d1(n1785) );
    mux2i_1 U1176 ( .x(n3463), .d0(n2592), .sl(n1856), .d1(n1786) );
    mux2i_1 U1177 ( .x(n3464), .d0(n2593), .sl(n1856), .d1(n1787) );
    mux2i_1 U1178 ( .x(n3465), .d0(n2594), .sl(n1856), .d1(n1788) );
    mux2i_1 U1179 ( .x(n3466), .d0(n2595), .sl(n1856), .d1(n1789) );
    nand3_1 U118 ( .x(n3935), .a(n3929), .b(___cell__6171_net27367), .c(
        WB_index_0) );
    mux2i_1 U1180 ( .x(n3467), .d0(n2596), .sl(n1856), .d1(n1790) );
    mux2i_1 U1181 ( .x(n3468), .d0(n2597), .sl(n1856), .d1(n1791) );
    mux2i_1 U1182 ( .x(n3469), .d0(n2598), .sl(n1856), .d1(n1792) );
    mux2i_1 U1183 ( .x(n3470), .d0(n2599), .sl(n1856), .d1(n1793) );
    mux2i_1 U1184 ( .x(n3471), .d0(n2600), .sl(n1856), .d1(n1794) );
    mux2i_1 U1185 ( .x(n3472), .d0(n2601), .sl(n1856), .d1(n1795) );
    mux2i_1 U1186 ( .x(n3473), .d0(n2602), .sl(n1856), .d1(n1796) );
    mux2i_1 U1187 ( .x(n3474), .d0(n2603), .sl(n1856), .d1(n1797) );
    mux2i_1 U1188 ( .x(n3475), .d0(n2604), .sl(n1856), .d1(n1798) );
    buf_3 U1189 ( .x(n920), .a(n989) );
    nand2_2 U119 ( .x(n3934), .a(reg_write_WB), .b(n555) );
    or2_2 U1190 ( .x(n1742), .a(n3927), .b(n3939) );
    mux2_2 U1191 ( .x(n3477), .d0(_RegFile_7__0), .sl(n1855), .d1(WB_data[0])
         );
    mux2_2 U1192 ( .x(n3478), .d0(_RegFile_7__1), .sl(n1855), .d1(WB_data[1])
         );
    mux2_2 U1193 ( .x(n3479), .d0(_RegFile_7__2), .sl(n1855), .d1(WB_data[2])
         );
    mux2_2 U1194 ( .x(n3480), .d0(_RegFile_7__3), .sl(n1855), .d1(WB_data[3])
         );
    mux2_2 U1195 ( .x(n3481), .d0(_RegFile_7__4), .sl(n1855), .d1(WB_data[4])
         );
    mux2_2 U1196 ( .x(n3482), .d0(_RegFile_7__5), .sl(n1855), .d1(WB_data[5])
         );
    mux2_2 U1197 ( .x(n3483), .d0(_RegFile_7__6), .sl(n1855), .d1(WB_data[6])
         );
    mux2_2 U1198 ( .x(n3484), .d0(_RegFile_7__7), .sl(n1855), .d1(n692) );
    mux2i_1 U1199 ( .x(n3486), .d0(n2583), .sl(n1855), .d1(n1801) );
    inv_6 U12 ( .x(reg_out_B[12]), .a(n750) );
    nand2i_2 U120 ( .x(n1602), .a(n1395), .b(n1511) );
    mux2i_1 U1200 ( .x(n3487), .d0(n2560), .sl(n1855), .d1(n1778) );
    mux2i_1 U1201 ( .x(n3488), .d0(n2561), .sl(n1855), .d1(n1779) );
    mux2i_1 U1202 ( .x(n3489), .d0(n2562), .sl(n1855), .d1(n1780) );
    mux2i_1 U1203 ( .x(n3490), .d0(n2563), .sl(n1855), .d1(n1781) );
    mux2i_1 U1204 ( .x(n3491), .d0(n2564), .sl(n1855), .d1(n1782) );
    mux2i_1 U1205 ( .x(n3492), .d0(n2565), .sl(n1855), .d1(n1783) );
    mux2i_1 U1206 ( .x(n3493), .d0(n2566), .sl(n1855), .d1(n1784) );
    mux2i_1 U1207 ( .x(n3494), .d0(n2567), .sl(n1855), .d1(n1785) );
    mux2i_1 U1208 ( .x(n3495), .d0(n2568), .sl(n1855), .d1(n1786) );
    mux2i_1 U1209 ( .x(n3496), .d0(n2569), .sl(n1855), .d1(n1787) );
    nand2i_2 U121 ( .x(n1600), .a(n1411), .b(n1511) );
    mux2i_1 U1210 ( .x(n3497), .d0(n2570), .sl(n1855), .d1(n1788) );
    mux2i_1 U1211 ( .x(n3498), .d0(n2571), .sl(n1855), .d1(n1789) );
    mux2i_1 U1212 ( .x(n3499), .d0(n2572), .sl(n1855), .d1(n1790) );
    mux2i_1 U1213 ( .x(n3500), .d0(n2573), .sl(n1855), .d1(n1791) );
    mux2i_1 U1214 ( .x(n3501), .d0(n2574), .sl(n1855), .d1(n1792) );
    mux2i_1 U1215 ( .x(n3502), .d0(n2575), .sl(n1855), .d1(n1793) );
    mux2i_1 U1216 ( .x(n3503), .d0(n2576), .sl(n1855), .d1(n1794) );
    mux2i_1 U1217 ( .x(n3504), .d0(n2577), .sl(n1855), .d1(n1795) );
    mux2i_1 U1218 ( .x(n3505), .d0(n2578), .sl(n1855), .d1(n1796) );
    mux2i_1 U1219 ( .x(n3506), .d0(n2579), .sl(n1855), .d1(n1797) );
    nand2i_2 U122 ( .x(n1648), .a(n1392), .b(n1511) );
    mux2i_1 U1220 ( .x(n3507), .d0(n2580), .sl(n1855), .d1(n1798) );
    or2_2 U1221 ( .x(n1743), .a(n3937), .b(n3938) );
    mux2_2 U1222 ( .x(n3509), .d0(_RegFile_6__0), .sl(n1854), .d1(WB_data[0])
         );
    mux2_2 U1223 ( .x(n3510), .d0(_RegFile_6__1), .sl(n1854), .d1(WB_data[1])
         );
    mux2_2 U1224 ( .x(n3511), .d0(_RegFile_6__2), .sl(n1854), .d1(WB_data[2])
         );
    mux2_2 U1225 ( .x(n3512), .d0(_RegFile_6__3), .sl(n1854), .d1(WB_data[3])
         );
    mux2_2 U1226 ( .x(n3513), .d0(_RegFile_6__4), .sl(n1854), .d1(WB_data[4])
         );
    mux2_2 U1227 ( .x(n3514), .d0(_RegFile_6__5), .sl(n1854), .d1(WB_data[5])
         );
    mux2_2 U1228 ( .x(n3515), .d0(_RegFile_6__6), .sl(n1854), .d1(WB_data[6])
         );
    mux2_2 U1229 ( .x(n3516), .d0(_RegFile_6__7), .sl(n1854), .d1(WB_data[7])
         );
    nand2i_2 U123 ( .x(n1646), .a(n1354), .b(n1511) );
    mux2i_1 U1230 ( .x(n3518), .d0(n2559), .sl(n1854), .d1(n1801) );
    mux2i_1 U1231 ( .x(n3519), .d0(n2536), .sl(n1854), .d1(n1778) );
    mux2i_1 U1232 ( .x(n3520), .d0(n2537), .sl(n1854), .d1(n1779) );
    mux2i_1 U1233 ( .x(n3521), .d0(n2538), .sl(n1854), .d1(n1780) );
    mux2i_1 U1234 ( .x(n3522), .d0(n2539), .sl(n1854), .d1(n1781) );
    mux2i_1 U1235 ( .x(n3523), .d0(n2540), .sl(n1854), .d1(n1782) );
    mux2i_1 U1236 ( .x(n3524), .d0(n2541), .sl(n1854), .d1(n1783) );
    mux2i_1 U1237 ( .x(n3525), .d0(n2542), .sl(n1854), .d1(n1784) );
    mux2i_1 U1238 ( .x(n3526), .d0(n2543), .sl(n1854), .d1(n1785) );
    mux2i_1 U1239 ( .x(n3527), .d0(n2544), .sl(n1854), .d1(n1786) );
    inv_8 U124 ( .x(n1740), .a(n1511) );
    mux2i_1 U1240 ( .x(n3528), .d0(n2545), .sl(n1854), .d1(n1787) );
    mux2i_1 U1241 ( .x(n3529), .d0(n2546), .sl(n1854), .d1(n1788) );
    mux2i_1 U1242 ( .x(n3530), .d0(n2547), .sl(n1854), .d1(n1789) );
    mux2i_1 U1243 ( .x(n3531), .d0(n2548), .sl(n1854), .d1(n1790) );
    mux2i_1 U1244 ( .x(n3532), .d0(n2549), .sl(n1854), .d1(n1791) );
    mux2i_1 U1245 ( .x(n3533), .d0(n2550), .sl(n1854), .d1(n1792) );
    mux2i_1 U1246 ( .x(n3534), .d0(n2551), .sl(n1854), .d1(n1793) );
    mux2i_1 U1247 ( .x(n3535), .d0(n2552), .sl(n1854), .d1(n1794) );
    mux2i_1 U1248 ( .x(n3536), .d0(n2553), .sl(n1854), .d1(n1795) );
    mux2i_1 U1249 ( .x(n3537), .d0(n2554), .sl(n1854), .d1(n1796) );
    inv_2 U125 ( .x(n1512), .a(n1303) );
    mux2i_1 U1250 ( .x(n3538), .d0(n2555), .sl(n1854), .d1(n1797) );
    mux2i_1 U1251 ( .x(n3539), .d0(n2556), .sl(n1854), .d1(n1798) );
    or2_2 U1252 ( .x(n1744), .a(n3936), .b(n3938) );
    mux2_2 U1253 ( .x(n3541), .d0(_RegFile_5__0), .sl(n1853), .d1(WB_data[0])
         );
    mux2_2 U1254 ( .x(n3542), .d0(_RegFile_5__1), .sl(n1853), .d1(WB_data[1])
         );
    mux2_2 U1255 ( .x(n3543), .d0(_RegFile_5__2), .sl(n1853), .d1(WB_data[2])
         );
    mux2_2 U1256 ( .x(n3544), .d0(_RegFile_5__3), .sl(n1853), .d1(WB_data[3])
         );
    mux2_2 U1257 ( .x(n3545), .d0(_RegFile_5__4), .sl(n1853), .d1(WB_data[4])
         );
    mux2_2 U1258 ( .x(n3546), .d0(_RegFile_5__5), .sl(n1853), .d1(WB_data[5])
         );
    mux2_2 U1259 ( .x(n3547), .d0(_RegFile_5__6), .sl(n1853), .d1(WB_data[6])
         );
    nand2i_2 U126 ( .x(n1644), .a(n1400), .b(n1511) );
    mux2_2 U1260 ( .x(n3548), .d0(_RegFile_5__7), .sl(n1853), .d1(WB_data[7])
         );
    mux2i_1 U1261 ( .x(n3550), .d0(n2535), .sl(n1853), .d1(n1801) );
    mux2i_1 U1262 ( .x(n3551), .d0(n2512), .sl(n1853), .d1(n1778) );
    mux2i_1 U1263 ( .x(n3552), .d0(n2513), .sl(n1853), .d1(n1779) );
    mux2i_1 U1264 ( .x(n3553), .d0(n2514), .sl(n1853), .d1(n1780) );
    mux2i_1 U1265 ( .x(n3554), .d0(n2515), .sl(n1853), .d1(n1781) );
    mux2i_1 U1266 ( .x(n3555), .d0(n2516), .sl(n1853), .d1(n1782) );
    mux2i_1 U1267 ( .x(n3556), .d0(n2517), .sl(n1853), .d1(n1783) );
    mux2i_1 U1268 ( .x(n3557), .d0(n2518), .sl(n1853), .d1(n1784) );
    mux2i_1 U1269 ( .x(n3558), .d0(n2519), .sl(n1853), .d1(n1785) );
    nand2i_2 U127 ( .x(n1642), .a(n1406), .b(n1511) );
    mux2i_1 U1270 ( .x(n3559), .d0(n2520), .sl(n1853), .d1(n1786) );
    mux2i_1 U1271 ( .x(n3560), .d0(n2521), .sl(n1853), .d1(n1787) );
    mux2i_1 U1272 ( .x(n3561), .d0(n2522), .sl(n1853), .d1(n1788) );
    mux2i_1 U1273 ( .x(n3562), .d0(n2523), .sl(n1853), .d1(n1789) );
    mux2i_1 U1274 ( .x(n3563), .d0(n2524), .sl(n1853), .d1(n1790) );
    mux2i_1 U1275 ( .x(n3564), .d0(n2525), .sl(n1853), .d1(n1791) );
    mux2i_1 U1276 ( .x(n3565), .d0(n2526), .sl(n1853), .d1(n1792) );
    mux2i_1 U1277 ( .x(n3566), .d0(n2527), .sl(n1853), .d1(n1793) );
    mux2i_1 U1278 ( .x(n3567), .d0(n2528), .sl(n1853), .d1(n1794) );
    mux2i_1 U1279 ( .x(n3568), .d0(n2529), .sl(n1853), .d1(n1795) );
    nand2i_2 U128 ( .x(n1640), .a(n1359), .b(n1511) );
    mux2i_1 U1280 ( .x(n3569), .d0(n2530), .sl(n1853), .d1(n1796) );
    mux2i_1 U1281 ( .x(n3570), .d0(n2531), .sl(n1853), .d1(n1797) );
    buf_3 U1282 ( .x(n978), .a(n983) );
    mux2i_1 U1283 ( .x(n3571), .d0(n2532), .sl(n1853), .d1(n1798) );
    or2_2 U1284 ( .x(n1745), .a(n3935), .b(n3938) );
    mux2_2 U1285 ( .x(n3573), .d0(_RegFile_4__0), .sl(n1852), .d1(WB_data[0])
         );
    mux2_2 U1286 ( .x(n3574), .d0(_RegFile_4__1), .sl(n1852), .d1(WB_data[1])
         );
    mux2_2 U1287 ( .x(n3575), .d0(_RegFile_4__2), .sl(n1852), .d1(WB_data[2])
         );
    mux2_2 U1288 ( .x(n3576), .d0(_RegFile_4__3), .sl(n1852), .d1(WB_data[3])
         );
    mux2_2 U1289 ( .x(n3577), .d0(_RegFile_4__4), .sl(n1852), .d1(WB_data[4])
         );
    nand2i_2 U129 ( .x(n1638), .a(n1304), .b(n1511) );
    mux2_2 U1290 ( .x(n3578), .d0(_RegFile_4__5), .sl(n1852), .d1(WB_data[5])
         );
    mux2_2 U1291 ( .x(n3579), .d0(_RegFile_4__6), .sl(n1852), .d1(WB_data[6])
         );
    mux2_2 U1292 ( .x(n3580), .d0(_RegFile_4__7), .sl(n1852), .d1(WB_data[7])
         );
    buf_3 U1293 ( .x(n924), .a(n937) );
    mux2i_1 U1294 ( .x(n3582), .d0(n2511), .sl(n1852), .d1(n1801) );
    mux2i_1 U1295 ( .x(n3583), .d0(n2488), .sl(n1852), .d1(n1778) );
    mux2i_1 U1296 ( .x(n3584), .d0(n2489), .sl(n1852), .d1(n1779) );
    mux2i_1 U1297 ( .x(n3585), .d0(n2490), .sl(n1852), .d1(n1780) );
    mux2i_1 U1298 ( .x(n3586), .d0(n2491), .sl(n1852), .d1(n1781) );
    mux2i_1 U1299 ( .x(n3587), .d0(n2492), .sl(n1852), .d1(n1782) );
    buf_3 U13 ( .x(Imm[27]), .a(N6382) );
    nand2i_2 U130 ( .x(n1636), .a(n1376), .b(n1303) );
    mux2i_1 U1300 ( .x(n3588), .d0(n2493), .sl(n1852), .d1(n1783) );
    mux2i_1 U1301 ( .x(n3589), .d0(n2494), .sl(n1852), .d1(n1784) );
    mux2i_1 U1302 ( .x(n3590), .d0(n2495), .sl(n1852), .d1(n1785) );
    mux2i_1 U1303 ( .x(n3591), .d0(n2496), .sl(n1852), .d1(n1786) );
    mux2i_1 U1304 ( .x(n3592), .d0(n2497), .sl(n1852), .d1(n1787) );
    mux2i_1 U1305 ( .x(n3593), .d0(n2498), .sl(n1852), .d1(n1788) );
    mux2i_1 U1306 ( .x(n3594), .d0(n2499), .sl(n1852), .d1(n1789) );
    mux2i_1 U1307 ( .x(n3595), .d0(n2500), .sl(n1852), .d1(n1790) );
    mux2i_1 U1308 ( .x(n3596), .d0(n2501), .sl(n1852), .d1(n1791) );
    mux2i_1 U1309 ( .x(n3597), .d0(n2502), .sl(n1852), .d1(n1792) );
    nand2i_2 U131 ( .x(n1634), .a(n1349), .b(n1303) );
    mux2i_1 U1310 ( .x(n3598), .d0(n2503), .sl(n1852), .d1(n1793) );
    mux2i_1 U1311 ( .x(n3599), .d0(n2504), .sl(n1852), .d1(n1794) );
    mux2i_1 U1312 ( .x(n3600), .d0(n2505), .sl(n1852), .d1(n1795) );
    mux2i_1 U1313 ( .x(n3601), .d0(n2506), .sl(n1852), .d1(n1796) );
    mux2i_1 U1314 ( .x(n3602), .d0(n2507), .sl(n1852), .d1(n1797) );
    buf_3 U1315 ( .x(n977), .a(n923) );
    mux2i_1 U1316 ( .x(n3603), .d0(n2508), .sl(n1852), .d1(n1798) );
    buf_3 U1317 ( .x(n925), .a(n937) );
    or2_2 U1318 ( .x(n1746), .a(n3927), .b(n3938) );
    mux2_2 U1319 ( .x(n3605), .d0(_RegFile_3__0), .sl(n1851), .d1(WB_data[0])
         );
    nand2i_2 U132 ( .x(n1632), .a(n1340), .b(n1303) );
    buf_3 U1320 ( .x(n927), .a(n936) );
    mux2_2 U1321 ( .x(n3606), .d0(_RegFile_3__1), .sl(n1851), .d1(WB_data[1])
         );
    mux2_2 U1322 ( .x(n3607), .d0(_RegFile_3__2), .sl(n1851), .d1(WB_data[2])
         );
    mux2_2 U1323 ( .x(n3608), .d0(_RegFile_3__3), .sl(n1851), .d1(WB_data[3])
         );
    mux2_2 U1324 ( .x(n3609), .d0(_RegFile_3__4), .sl(n1851), .d1(WB_data[4])
         );
    mux2_2 U1325 ( .x(n3610), .d0(_RegFile_3__5), .sl(n1851), .d1(WB_data[5])
         );
    mux2_2 U1326 ( .x(n3611), .d0(_RegFile_3__6), .sl(n1851), .d1(WB_data[6])
         );
    mux2_2 U1327 ( .x(n3612), .d0(_RegFile_3__7), .sl(n1851), .d1(WB_data[7])
         );
    mux2i_1 U1328 ( .x(n3614), .d0(n2487), .sl(n1851), .d1(n1801) );
    mux2i_1 U1329 ( .x(n3615), .d0(n2464), .sl(n1851), .d1(n1778) );
    nand2i_2 U133 ( .x(n1630), .a(n1383), .b(n1303) );
    mux2i_1 U1330 ( .x(n3616), .d0(n2465), .sl(n1851), .d1(n1779) );
    mux2i_1 U1331 ( .x(n3617), .d0(n2466), .sl(n1851), .d1(n1780) );
    mux2i_1 U1332 ( .x(n3618), .d0(n2467), .sl(n1851), .d1(n1781) );
    mux2i_1 U1333 ( .x(n3619), .d0(n2468), .sl(n1851), .d1(n1782) );
    mux2i_1 U1334 ( .x(n3620), .d0(n2469), .sl(n1851), .d1(n1783) );
    mux2i_1 U1335 ( .x(n3621), .d0(n2470), .sl(n1851), .d1(n1784) );
    mux2i_1 U1336 ( .x(n3622), .d0(n2471), .sl(n1851), .d1(n1785) );
    mux2i_1 U1337 ( .x(n3623), .d0(n2472), .sl(n1851), .d1(n1786) );
    mux2i_1 U1338 ( .x(n3624), .d0(n2473), .sl(n1851), .d1(n1787) );
    mux2i_1 U1339 ( .x(n3625), .d0(n2474), .sl(n1851), .d1(n1788) );
    nand2i_2 U134 ( .x(n1628), .a(n1381), .b(n1303) );
    mux2i_1 U1340 ( .x(n3626), .d0(n2475), .sl(n1851), .d1(n1789) );
    mux2i_1 U1341 ( .x(n3627), .d0(n2476), .sl(n1851), .d1(n1790) );
    mux2i_1 U1342 ( .x(n3628), .d0(n2477), .sl(n1851), .d1(n1791) );
    mux2i_1 U1343 ( .x(n3629), .d0(n2478), .sl(n1851), .d1(n1792) );
    mux2i_1 U1344 ( .x(n3630), .d0(n2479), .sl(n1851), .d1(n1793) );
    mux2i_1 U1345 ( .x(n3631), .d0(n2480), .sl(n1851), .d1(n1794) );
    mux2i_1 U1346 ( .x(n3632), .d0(n2481), .sl(n1851), .d1(n1795) );
    mux2i_1 U1347 ( .x(n3633), .d0(n2482), .sl(n1851), .d1(n1796) );
    mux2i_1 U1348 ( .x(n3634), .d0(n2483), .sl(n1851), .d1(n1797) );
    mux2i_1 U1349 ( .x(n3635), .d0(n2484), .sl(n1851), .d1(n1798) );
    nand2i_2 U135 ( .x(n1626), .a(n1379), .b(n1303) );
    or2_2 U1350 ( .x(n1747), .a(n3934), .b(n3937) );
    mux2_2 U1351 ( .x(n3637), .d0(_RegFile_2__0), .sl(n1848), .d1(WB_data[0])
         );
    mux2_2 U1352 ( .x(n3638), .d0(_RegFile_2__1), .sl(n1848), .d1(WB_data[1])
         );
    mux2_2 U1353 ( .x(n3639), .d0(_RegFile_2__2), .sl(n1848), .d1(WB_data[2])
         );
    mux2_2 U1354 ( .x(n3640), .d0(_RegFile_2__3), .sl(n1848), .d1(WB_data[3])
         );
    mux2_2 U1355 ( .x(n3641), .d0(_RegFile_2__4), .sl(n1848), .d1(WB_data[4])
         );
    mux2_2 U1356 ( .x(n3642), .d0(_RegFile_2__5), .sl(n1848), .d1(WB_data[5])
         );
    mux2_2 U1357 ( .x(n3643), .d0(_RegFile_2__6), .sl(n1848), .d1(WB_data[6])
         );
    mux2_2 U1358 ( .x(n3644), .d0(_RegFile_2__7), .sl(n1848), .d1(WB_data[7])
         );
    mux2i_1 U1359 ( .x(n3646), .d0(n2415), .sl(n1848), .d1(n1801) );
    nand2i_2 U136 ( .x(n1624), .a(n1374), .b(n1303) );
    mux2i_1 U1360 ( .x(n3647), .d0(n2392), .sl(n1848), .d1(n1778) );
    mux2i_1 U1361 ( .x(n3648), .d0(n2393), .sl(n1848), .d1(n1779) );
    mux2i_1 U1362 ( .x(n3649), .d0(n2394), .sl(n1848), .d1(n1780) );
    mux2i_1 U1363 ( .x(n3650), .d0(n2395), .sl(n1848), .d1(n1781) );
    mux2i_1 U1364 ( .x(n3651), .d0(n2396), .sl(n1848), .d1(n1782) );
    buf_3 U1365 ( .x(n930), .a(n987) );
    mux2i_1 U1366 ( .x(n3652), .d0(n2397), .sl(n1848), .d1(n1783) );
    mux2i_1 U1367 ( .x(n3653), .d0(n2398), .sl(n1848), .d1(n1784) );
    mux2i_1 U1368 ( .x(n3654), .d0(n2399), .sl(n1848), .d1(n1785) );
    mux2i_1 U1369 ( .x(n3655), .d0(n2400), .sl(n1848), .d1(n1786) );
    nand2i_2 U137 ( .x(n1622), .a(n1403), .b(n1303) );
    mux2i_1 U1370 ( .x(n3656), .d0(n2401), .sl(n1848), .d1(n1787) );
    mux2i_1 U1371 ( .x(n3657), .d0(n2402), .sl(n1848), .d1(n1788) );
    mux2i_1 U1372 ( .x(n3658), .d0(n2403), .sl(n1848), .d1(n1789) );
    mux2i_1 U1373 ( .x(n3659), .d0(n2404), .sl(n1848), .d1(n1790) );
    mux2i_1 U1374 ( .x(n3660), .d0(n2405), .sl(n1848), .d1(n1791) );
    mux2i_1 U1375 ( .x(n3661), .d0(n2406), .sl(n1848), .d1(n1792) );
    mux2i_1 U1376 ( .x(n3662), .d0(n2407), .sl(n1848), .d1(n1793) );
    mux2i_1 U1377 ( .x(n3663), .d0(n2408), .sl(n1848), .d1(n1794) );
    mux2i_1 U1378 ( .x(n3664), .d0(n2409), .sl(n1848), .d1(n1795) );
    mux2i_1 U1379 ( .x(n3665), .d0(n2410), .sl(n1848), .d1(n1796) );
    nand2i_2 U138 ( .x(n1620), .a(n1409), .b(n1303) );
    mux2i_1 U1380 ( .x(n3666), .d0(n2411), .sl(n1848), .d1(n1797) );
    mux2i_1 U1381 ( .x(n3667), .d0(n2412), .sl(n1848), .d1(n1798) );
    buf_3 U1382 ( .x(n929), .a(n987) );
    or2_2 U1383 ( .x(n1750), .a(n3934), .b(n3936) );
    mux2_2 U1384 ( .x(n3669), .d0(_RegFile_1__0), .sl(n1837), .d1(WB_data[0])
         );
    mux2_2 U1385 ( .x(n3670), .d0(_RegFile_1__1), .sl(n1837), .d1(WB_data[1])
         );
    mux2_2 U1386 ( .x(n3671), .d0(_RegFile_1__2), .sl(n1837), .d1(WB_data[2])
         );
    mux2_2 U1387 ( .x(n3672), .d0(_RegFile_1__3), .sl(n1837), .d1(WB_data[3])
         );
    mux2_2 U1388 ( .x(n3673), .d0(_RegFile_1__4), .sl(n1837), .d1(WB_data[4])
         );
    mux2_2 U1389 ( .x(n3674), .d0(_RegFile_1__5), .sl(n1837), .d1(WB_data[5])
         );
    nand2i_2 U139 ( .x(n1618), .a(n1338), .b(n1303) );
    mux2_2 U1390 ( .x(n3675), .d0(_RegFile_1__6), .sl(n1837), .d1(WB_data[6])
         );
    mux2_2 U1391 ( .x(n3676), .d0(_RegFile_1__7), .sl(n1837), .d1(WB_data[7])
         );
    inv_2 U1392 ( .x(n1603), .a(n1601) );
    mux2i_1 U1393 ( .x(n3678), .d0(n2151), .sl(n1837), .d1(n1801) );
    mux2i_1 U1394 ( .x(n3679), .d0(n2128), .sl(n1837), .d1(n1778) );
    mux2i_1 U1395 ( .x(n3680), .d0(n2129), .sl(n1837), .d1(n1779) );
    mux2i_1 U1396 ( .x(n3681), .d0(n2130), .sl(n1837), .d1(n1780) );
    mux2i_1 U1397 ( .x(n3682), .d0(n2131), .sl(n1837), .d1(n1781) );
    mux2i_1 U1398 ( .x(n3683), .d0(n2132), .sl(n1837), .d1(n1782) );
    mux2i_1 U1399 ( .x(n3684), .d0(n2133), .sl(n1837), .d1(n1783) );
    exor2_1 U14 ( .x(n3945), .a(n3933), .b(opcode_of_MEM_4) );
    nand2i_2 U140 ( .x(n1616), .a(n1361), .b(n1303) );
    mux2i_1 U1400 ( .x(n3685), .d0(n2134), .sl(n1837), .d1(n1784) );
    mux2i_1 U1401 ( .x(n3686), .d0(n2135), .sl(n1837), .d1(n1785) );
    mux2i_1 U1402 ( .x(n3687), .d0(n2136), .sl(n1837), .d1(n1786) );
    mux2i_1 U1403 ( .x(n3688), .d0(n2137), .sl(n1837), .d1(n1787) );
    mux2i_1 U1404 ( .x(n3689), .d0(n2138), .sl(n1837), .d1(n1788) );
    buf_3 U1405 ( .x(n962), .a(n984) );
    mux2i_1 U1406 ( .x(n3690), .d0(n2139), .sl(n1837), .d1(n1789) );
    mux2i_1 U1407 ( .x(n3691), .d0(n2140), .sl(n1837), .d1(n1790) );
    mux2i_1 U1408 ( .x(n3692), .d0(n2141), .sl(n1837), .d1(n1791) );
    mux2i_1 U1409 ( .x(n3693), .d0(n2142), .sl(n1837), .d1(n1792) );
    nand2i_2 U141 ( .x(n1614), .a(n1346), .b(n1303) );
    mux2i_1 U1410 ( .x(n3694), .d0(n2143), .sl(n1837), .d1(n1793) );
    mux2i_1 U1411 ( .x(n3695), .d0(n2144), .sl(n1837), .d1(n1794) );
    mux2i_1 U1412 ( .x(n3696), .d0(n2145), .sl(n1837), .d1(n1795) );
    mux2i_1 U1413 ( .x(n3697), .d0(n2146), .sl(n1837), .d1(n1796) );
    mux2i_1 U1414 ( .x(n3698), .d0(n2147), .sl(n1837), .d1(n1797) );
    buf_3 U1415 ( .x(n963), .a(n984) );
    mux2i_1 U1416 ( .x(n3699), .d0(n2148), .sl(n1837), .d1(n1798) );
    or2_2 U1417 ( .x(n1761), .a(n3934), .b(n3935) );
    mux2_2 U1418 ( .x(n3701), .d0(_RegFile_0__0), .sl(n1826), .d1(n690) );
    mux2_2 U1419 ( .x(n3702), .d0(_RegFile_0__1), .sl(n1826), .d1(n688) );
    nand2i_2 U142 ( .x(n1612), .a(n1357), .b(n1303) );
    mux2_2 U1420 ( .x(n3703), .d0(_RegFile_0__2), .sl(n1826), .d1(WB_data[2])
         );
    mux2_2 U1421 ( .x(n3704), .d0(_RegFile_0__3), .sl(n1826), .d1(WB_data[3])
         );
    mux2_2 U1422 ( .x(n3705), .d0(_RegFile_0__4), .sl(n1826), .d1(n687) );
    mux2_2 U1423 ( .x(n3706), .d0(_RegFile_0__5), .sl(n1826), .d1(n689) );
    mux2_2 U1424 ( .x(n3707), .d0(_RegFile_0__6), .sl(n1826), .d1(WB_data[6])
         );
    mux2_2 U1425 ( .x(n3708), .d0(_RegFile_0__7), .sl(n1826), .d1(WB_data[7])
         );
    inv_2 U1426 ( .x(n1800), .a(n1601) );
    nand2i_2 U1427 ( .x(n1772), .a(n3930), .b(reg_write_WB) );
    mux2i_1 U1428 ( .x(n3733), .d0(n1423), .sl(___cell__36997_net126612), .d1(
        n1424) );
    mux2i_2 U1429 ( .x(_current_IR_reg_1_net49291), .d0(n800), .sl(
        ___cell__36997_net130681), .d1(n801) );
    nand2i_2 U143 ( .x(n1610), .a(n1343), .b(n1303) );
    inv_2 U1430 ( .x(n800), .a(current_IR_1) );
    mux2i_1 U1431 ( .x(n3734), .d0(n1421), .sl(___cell__36997_net126612), .d1(
        n1422) );
    mux2i_1 U1432 ( .x(n3736), .d0(n1418), .sl(___cell__36997_net126612), .d1(
        n1419) );
    mux2i_1 U1433 ( .x(n3738), .d0(n631), .sl(___cell__36997_net126612), .d1(
        n1596) );
    mux2i_1 U1434 ( .x(n3740), .d0(n630), .sl(___cell__36997_net126612), .d1(
        n1593) );
    mux2i_1 U1435 ( .x(n3741), .d0(n629), .sl(___cell__36997_net130681), .d1(
        n1592) );
    mux2i_1 U1436 ( .x(n3742), .d0(n632), .sl(___cell__36997_net126612), .d1(
        n1597) );
    mux2i_1 U1437 ( .x(n3746), .d0(n569), .sl(___cell__36997_net126612), .d1(
        n1413) );
    mux2i_1 U1438 ( .x(n3748), .d0(n645), .sl(___cell__36997_net126612), .d1(
        n1330) );
    mux2i_1 U1439 ( .x(n3749), .d0(n1332), .sl(___cell__36997_net130681), .d1(
        n1333) );
    nand2i_2 U144 ( .x(n1608), .a(n1363), .b(n1303) );
    mux2i_1 U1440 ( .x(n3756), .d0(n1323), .sl(___cell__36997_net130681), .d1(
        n1324) );
    mux2i_1 U1441 ( .x(n3759), .d0(n1318), .sl(___cell__36997_net126612), .d1(
        n1319) );
    inv_5 U1442 ( .x(n1319), .a(IR_latched_input[27]) );
    nand2i_2 U1443 ( .x(n1066), .a(n1860), .b(n1718) );
    oai21_1 U1444 ( .x(n3765), .a(n1065), .b(___cell__36997_net126621), .c(
        n1066) );
    nand2i_2 U1445 ( .x(n1074), .a(n1863), .b(n642) );
    nand2i_2 U1446 ( .x(n1107), .a(n2637), .b(n1718) );
    nand2i_3 U1447 ( .x(n1098), .a(n2635), .b(n1718) );
    nand2i_2 U1448 ( .x(n1086), .a(n2636), .b(n642) );
    oai21_1 U1449 ( .x(n3778), .a(n1065), .b(n1085), .c(n1086) );
    nor3_1 U145 ( .x(n1302), .a(n1303), .b(n1304), .c(n1305) );
    nor2i_1 U1450 ( .x(n1097), .a(n1716), .b(n1485) );
    aoi21_1 U1451 ( .x(n1069), .a(rd_addr[1]), .b(n642), .c(n1719) );
    oai21_1 U1452 ( .x(n3784), .a(n1065), .b(n1061), .c(n1076) );
    aoi21_1 U1453 ( .x(n1076), .a(rd_addr[3]), .b(n642), .c(n1719) );
    aoi21_1 U1454 ( .x(n1070), .a(rd_addr[4]), .b(n1718), .c(n1802) );
    oai21_1 U1455 ( .x(n3785), .a(n1775), .b(n1063), .c(n1070) );
    buf_3 U1456 ( .x(n917), .a(n990) );
    nand2i_2 U1457 ( .x(n1077), .a(n561), .b(n642) );
    nand2i_2 U1458 ( .x(n1122), .a(n671), .b(n1718) );
    inv_5 U1459 ( .x(n1718), .a(n705) );
    nand2i_2 U146 ( .x(n1606), .a(___cell__36997_net129389), .b(n1303) );
    nand2i_2 U1460 ( .x(n1133), .a(n558), .b(n642) );
    oai21_1 U1461 ( .x(n3790), .a(n1132), .b(n1775), .c(n1133) );
    buf_3 U1462 ( .x(n918), .a(n988) );
    buf_3 U1463 ( .x(n919), .a(n988) );
    nand2i_2 U1464 ( .x(n1213), .a(n590), .b(net150785) );
    inv_5 U1465 ( .x(n1650), .a(n1773) );
    inv_2 U1466 ( .x(n856), .a(n340) );
    inv_2 U1467 ( .x(n1682), .a(N504) );
    mux2i_1 U1468 ( .x(n3891), .d0(n1682), .sl(n1650), .d1(
        ___cell__36997_net129389) );
    nor2i_1 U1469 ( .x(n1000), .a(___cell__36997_net130681), .b(n1484) );
    oai21_1 U147 ( .x(n1485), .a(___cell__36997_net127190), .b(n1263), .c(
        n1307) );
    inv_2 U1470 ( .x(n679), .a(n1000) );
    buf_3 U1471 ( .x(n912), .a(n951) );
    buf_3 U1472 ( .x(n913), .a(n952) );
    inv_2 U1473 ( .x(n1728), .a(reg_dst_of_EX_0) );
    buf_3 U1474 ( .x(n914), .a(n952) );
    inv_2 U1475 ( .x(n801), .a(IR_latched_input[1]) );
    inv_1 U1476 ( .x(n1530), .a(NPC[24]) );
    inv_0 U1477 ( .x(n1529), .a(NPC[25]) );
    and3i_1 U1478 ( .x(PIPEEMPTY), .a(n993), .b(n991), .c(n992) );
    nor2i_1 U1479 ( .x(n991), .a(n1726), .b(n1725) );
    nand2i_2 U148 ( .x(n1716), .a(n2638), .b(n1718) );
    inv_2 U1480 ( .x(n992), .a(n3930) );
    nand2_2 U1481 ( .x(n3930), .a(n3931), .b(n555) );
    inv_2 U1482 ( .x(n3931), .a(n3927) );
    nand2i_2 U1483 ( .x(n993), .a(n1727), .b(n1729) );
    inv_2 U1484 ( .x(n1354), .a(WB_data[11]) );
    inv_2 U1485 ( .x(n1359), .a(WB_data[14]) );
    inv_2 U1486 ( .x(n1383), .a(WB_data[19]) );
    inv_2 U1487 ( .x(n1374), .a(WB_data[22]) );
    inv_2 U1488 ( .x(n1346), .a(WB_data[27]) );
    inv_2 U1489 ( .x(n1343), .a(WB_data[29]) );
    inv_5 U149 ( .x(n843), .a(n847) );
    inv_2 U1490 ( .x(n1532), .a(NPC[22]) );
    inv_2 U1491 ( .x(n1395), .a(WB_data[8]) );
    inv_2 U1492 ( .x(n1552), .a(NPC[1]) );
    inv_2 U1493 ( .x(n1553), .a(NPC[0]) );
    inv_2 U1494 ( .x(n1363), .a(WB_data[30]) );
    inv_2 U1495 ( .x(n1595), .a(IR_latched_input[7]) );
    inv_2 U1496 ( .x(n1594), .a(current_IR_7) );
    inv_2 U1497 ( .x(n1534), .a(NPC[20]) );
    inv_2 U1498 ( .x(n1531), .a(NPC[23]) );
    inv_0 U1499 ( .x(n1536), .a(NPC[18]) );
    buf_14 U15 ( .x(reg_out_A[11]), .a(n3967) );
    inv_2 U150 ( .x(n1316), .a(IR_latched_input[28]) );
    inv_2 U1500 ( .x(n851), .a(IR_latched_input[26]) );
    inv_2 U1501 ( .x(___cell__36997_net129389), .a(WB_data[31]) );
    inv_0 U1502 ( .x(n1535), .a(NPC[19]) );
    inv_2 U1503 ( .x(n1361), .a(WB_data[26]) );
    inv_2 U1504 ( .x(n1439), .a(n4454) );
    inv_1 U1505 ( .x(n1311), .a(Imm[31]) );
    inv_2 U1506 ( .x(n1411), .a(WB_data[9]) );
    inv_2 U1507 ( .x(n1392), .a(WB_data[10]) );
    inv_2 U1508 ( .x(n1400), .a(WB_data[12]) );
    inv_2 U1509 ( .x(n1406), .a(WB_data[13]) );
    and2_3 U151 ( .x(n642), .a(n704), .b(n1461) );
    inv_2 U1510 ( .x(n1304), .a(WB_data[15]) );
    inv_2 U1511 ( .x(n1376), .a(WB_data[16]) );
    inv_2 U1512 ( .x(n1349), .a(WB_data[17]) );
    inv_2 U1513 ( .x(n1340), .a(WB_data[18]) );
    inv_2 U1514 ( .x(n1381), .a(WB_data[20]) );
    inv_2 U1515 ( .x(n1379), .a(WB_data[21]) );
    inv_2 U1516 ( .x(n1403), .a(WB_data[23]) );
    inv_2 U1517 ( .x(n1409), .a(WB_data[24]) );
    inv_2 U1518 ( .x(n1338), .a(WB_data[25]) );
    inv_2 U1519 ( .x(n1357), .a(WB_data[28]) );
    inv_2 U1520 ( .x(n1287), .a(EPC_23) );
    inv_2 U1521 ( .x(n1283), .a(EPC_25) );
    inv_2 U1522 ( .x(n1423), .a(current_IR_0) );
    inv_2 U1523 ( .x(n1421), .a(current_IR_2) );
    inv_5 U1524 ( .x(n1418), .a(current_IR_4) );
    inv_2 U1525 ( .x(n1332), .a(current_IR_17) );
    inv_2 U1526 ( .x(n1323), .a(current_IR_24) );
    inv_5 U1527 ( .x(n1318), .a(current_IR_27) );
    inv_2 U1528 ( .x(n1686), .a(WB_index_1) );
    inv_2 U1529 ( .x(n1424), .a(IR_latched_input[0]) );
    inv_2 U1530 ( .x(n1422), .a(IR_latched_input[2]) );
    inv_2 U1531 ( .x(n1417), .a(IR_latched_input[5]) );
    inv_2 U1532 ( .x(n1596), .a(IR_latched_input[6]) );
    inv_2 U1533 ( .x(n1593), .a(IR_latched_input[8]) );
    inv_2 U1534 ( .x(n1592), .a(IR_latched_input[9]) );
    inv_2 U1535 ( .x(n1416), .a(IR_latched_input[11]) );
    inv_2 U1536 ( .x(n1415), .a(IR_latched_input[12]) );
    inv_2 U1537 ( .x(n1414), .a(IR_latched_input[13]) );
    inv_2 U1538 ( .x(n1413), .a(IR_latched_input[14]) );
    inv_2 U1539 ( .x(n1412), .a(IR_latched_input[15]) );
    inv_2 U1540 ( .x(n1331), .a(IR_latched_input[20]) );
    inv_2 U1541 ( .x(n1324), .a(IR_latched_input[24]) );
    inv_2 U1542 ( .x(n1527), .a(NPC[27]) );
    inv_2 U1543 ( .x(n1526), .a(NPC[28]) );
    inv_2 U1544 ( .x(n1525), .a(NPC[29]) );
    inv_2 U1545 ( .x(n1524), .a(NPC[30]) );
    inv_2 U1546 ( .x(___cell__36997_net129786), .a(NPC[31]) );
    and2_1 U1547 ( .x(n555), .a(n3925), .b(n3926) );
    and2_1 U1548 ( .x(n556), .a(opcode_of_MEM_2), .b(opcode_of_MEM_4) );
    mux2i_1 U1549 ( .x(n628), .d0(n3946), .sl(opcode_of_MEM_1), .d1(n3947) );
    nor2i_6 U155 ( .x(n1691), .a(n772), .b(n340) );
    mux2_6 U1550 ( .x(n637), .d0(n1410), .sl(___cell__36997_net129354), .d1(
        n1411) );
    mux2_6 U1551 ( .x(n640), .d0(n1380), .sl(___cell__36997_net129354), .d1(
        n1381) );
    inv_16 U1552 ( .x(n1778), .a(n1647) );
    inv_16 U1553 ( .x(n1779), .a(n1645) );
    inv_16 U1554 ( .x(n1780), .a(n1643) );
    inv_16 U1555 ( .x(n1781), .a(n1641) );
    inv_16 U1556 ( .x(n1782), .a(n1639) );
    inv_16 U1557 ( .x(n1783), .a(n1637) );
    inv_16 U1558 ( .x(n1784), .a(n1635) );
    inv_16 U1559 ( .x(n1785), .a(n1633) );
    inv_5 U156 ( .x(n1071), .a(n339) );
    inv_16 U1560 ( .x(n1786), .a(n1631) );
    inv_16 U1561 ( .x(n1787), .a(n1629) );
    inv_16 U1562 ( .x(n1788), .a(n1627) );
    inv_16 U1563 ( .x(n1789), .a(n1625) );
    inv_16 U1564 ( .x(n1790), .a(n1623) );
    inv_16 U1565 ( .x(n1791), .a(n1621) );
    inv_16 U1566 ( .x(n1792), .a(n1619) );
    inv_16 U1567 ( .x(n1793), .a(n1617) );
    inv_16 U1568 ( .x(n1794), .a(n1615) );
    inv_16 U1569 ( .x(n1795), .a(n1613) );
    and3i_1 U157 ( .x(n1735), .a(n1687), .b(n1575), .c(reg_write_WB) );
    inv_16 U1570 ( .x(n1796), .a(n1611) );
    inv_16 U1571 ( .x(n1797), .a(n1609) );
    inv_16 U1572 ( .x(n1798), .a(n1607) );
    nand2_2 U1573 ( .x(n1604), .a(n1605), .b(n1606) );
    inv_5 U1574 ( .x(n1799), .a(n1604) );
    nand2_2 U1575 ( .x(n1599), .a(n1514), .b(n1600) );
    inv_5 U1576 ( .x(n1801), .a(n1599) );
    inv_16 U1577 ( .x(n1803), .a(n1520) );
    buf_3 U1578 ( .x(n949), .a(n932) );
    buf_3 U1579 ( .x(n950), .a(n932) );
    nand2_2 U158 ( .x(n1734), .a(n1574), .b(n1573) );
    buf_3 U1580 ( .x(n967), .a(n922) );
    buf_3 U1581 ( .x(n966), .a(n922) );
    buf_3 U1582 ( .x(n975), .a(n922) );
    buf_3 U1583 ( .x(n974), .a(n922) );
    buf_3 U1584 ( .x(n976), .a(n923) );
    buf_3 U1585 ( .x(n968), .a(n952) );
    buf_3 U1586 ( .x(n947), .a(n938) );
    buf_3 U1587 ( .x(n969), .a(n952) );
    buf_3 U1588 ( .x(n948), .a(n938) );
    buf_3 U1589 ( .x(n964), .a(n952) );
    exnor2_1 U159 ( .x(n1573), .a(n772), .b(n3926) );
    buf_3 U1590 ( .x(n983), .a(n1858) );
    buf_3 U1591 ( .x(n923), .a(n915) );
    buf_3 U1592 ( .x(n954), .a(n926) );
    buf_3 U1593 ( .x(n972), .a(n986) );
    buf_3 U1594 ( .x(n922), .a(n915) );
    buf_3 U1595 ( .x(n957), .a(n945) );
    buf_3 U1596 ( .x(n945), .a(n939) );
    buf_3 U1597 ( .x(n926), .a(n936) );
    buf_3 U1598 ( .x(n932), .a(n961) );
    buf_3 U1599 ( .x(n938), .a(n961) );
    buf_14 U16 ( .x(Imm[19]), .a(N6366) );
    buf_3 U160 ( .x(n892), .a(n339) );
    buf_3 U1600 ( .x(n939), .a(n961) );
    buf_3 U1601 ( .x(n934), .a(n984) );
    buf_3 U1602 ( .x(n984), .a(n936) );
    buf_3 U1603 ( .x(n961), .a(n988) );
    buf_3 U1604 ( .x(n937), .a(n987) );
    buf_3 U1605 ( .x(n915), .a(n951) );
    buf_3 U1606 ( .x(n988), .a(n921) );
    buf_3 U1607 ( .x(n952), .a(n936) );
    buf_3 U1608 ( .x(n951), .a(n936) );
    buf_3 U1609 ( .x(n987), .a(n921) );
    inv_2 U161 ( .x(n1333), .a(IR_latched_input[17]) );
    buf_3 U1610 ( .x(n970), .a(n972) );
    buf_3 U1611 ( .x(n971), .a(n972) );
    buf_3 U1612 ( .x(n921), .a(n989) );
    buf_3 U1613 ( .x(n990), .a(n970) );
    buf_3 U1614 ( .x(n916), .a(n990) );
    buf_3 U1615 ( .x(n981), .a(n980) );
    buf_3 U1616 ( .x(n989), .a(n971) );
    buf_3 U1617 ( .x(n935), .a(n988) );
    buf_3 U1618 ( .x(n936), .a(n987) );
    buf_3 U1619 ( .x(n980), .a(n983) );
    buf_3 U1620 ( .x(n985), .a(n935) );
    buf_3 U1621 ( .x(n979), .a(n983) );
    buf_3 U1622 ( .x(n982), .a(n964) );
    buf_3 U1623 ( .x(n911), .a(n951) );
    buf_3 U1624 ( .x(n973), .a(n954) );
    buf_3 U1625 ( .x(n953), .a(n926) );
    buf_3 U1626 ( .x(n986), .a(n981) );
    buf_3 U1627 ( .x(n956), .a(n986) );
    buf_3 U1628 ( .x(n955), .a(n986) );
    inv_2 U1631 ( .x(n1330), .a(IR_latched_input[16]) );
    ao22_2 U1633 ( .x(n650), .a(n883), .b(n882), .c(n1517), .d(n881) );
    mux2_5 U1634 ( .x(n653), .d0(n1367), .sl(___cell__36997_net129354), .d1(
        n1368) );
    inv_2 U1635 ( .x(n335), .a(n879) );
    inv_10 U1637 ( .x(net152024), .a(n728) );
    inv_6 U1638 ( .x(___cell__36997_net130705), .a(net148858) );
    inv_6 U1639 ( .x(net148913), .a(___cell__36997_net130705) );
    inv_2 U1640 ( .x(n1328), .a(IR_latched_input[22]) );
    inv_2 U1641 ( .x(n1326), .a(IR_latched_input[23]) );
    buf_16 U1642 ( .x(reg_out_B[17]), .a(n3978) );
    or2_2 U1644 ( .x(n668), .a(___cell__36997_net129247), .b(n1277) );
    inv_2 U1645 ( .x(n1325), .a(IR_latched_input[21]) );
    inv_12 U1646 ( .x(n1688), .a(n1083) );
    mux2_6 U1647 ( .x(n672), .d0(n1384), .sl(___cell__36997_net129354), .d1(
        n1385) );
    mux2_6 U1648 ( .x(n673), .d0(n1386), .sl(___cell__36997_net129354), .d1(
        n1387) );
    mux2_6 U1649 ( .x(n674), .d0(n1339), .sl(___cell__36997_net129354), .d1(
        n1340) );
    inv_2 U165 ( .x(reg_dst_of_EX_3), .a(n702) );
    mux2i_5 U1650 ( .x(n1336), .d0(n1337), .sl(___cell__36997_net129354), .d1(
        n1338) );
    inv_7 U1651 ( .x(n698), .a(n1336) );
    nand2_2 U1652 ( .x(n675), .a(___cell__36997_net130713), .b(N6039) );
    inv_2 U1653 ( .x(n693), .a(n333) );
    nand2_2 U1654 ( .x(n676), .a(___cell__36997_net130713), .b(N6040) );
    nand2i_4 U1655 ( .x(n1522), .a(n1523), .b(n1445) );
    inv_7 U1656 ( .x(n744), .a(n1522) );
    nand3i_2 U1657 ( .x(n3948), .a(___cell__36997_net125928), .b(n1000), .c(
        n744) );
    nand2i_2 U1658 ( .x(n1515), .a(n1516), .b(n1517) );
    or3i_5 U1659 ( .x(n680), .a(n744), .b(___cell__36997_net125928), .c(n679)
         );
    nand3_1 U166 ( .x(n1727), .a(n1559), .b(n702), .c(n1728) );
    inv_7 U1660 ( .x(___cell__36997_net125928), .a(___cell__36997_net129626)
         );
    buf_10 U1661 ( .x(reg_out_A[27]), .a(n3954) );
    inv_4 U1662 ( .x(n682), .a(n782) );
    inv_5 U1663 ( .x(n1466), .a(n782) );
    nand4_4 U1664 ( .x(n1706), .a(n639), .b(n640), .c(n1014), .d(n663) );
    nor2_6 U1665 ( .x(n1703), .a(n1701), .b(n1702) );
    nand4_5 U1666 ( .x(n1710), .a(n1128), .b(n637), .c(n1020), .d(n1003) );
    inv_6 U1667 ( .x(n1024), .a(n1344) );
    aoi22_1 U1668 ( .x(n1144), .a(n1344), .b(n797), .c(EPC_27), .d(net150625)
         );
    inv_0 U1669 ( .x(n683), .a(n847) );
    nand3_1 U167 ( .x(n3927), .a(___cell__6171_net27367), .b(n3928), .c(n3929)
         );
    inv_6 U1670 ( .x(n847), .a(n850) );
    inv_0 U1671 ( .x(n684), .a(n1377) );
    mux2i_2 U1672 ( .x(n1377), .d0(n1378), .sl(___cell__36997_net129354), .d1(
        n1379) );
    inv_4 U1673 ( .x(n1014), .a(n1377) );
    inv_2 U1674 ( .x(n685), .a(n1387) );
    inv_2 U1675 ( .x(n1387), .a(WB_data[3]) );
    inv_2 U1676 ( .x(n686), .a(n1390) );
    inv_2 U1677 ( .x(n1390), .a(WB_data[2]) );
    inv_2 U1678 ( .x(n687), .a(n1397) );
    inv_2 U1679 ( .x(n1397), .a(WB_data[4]) );
    nand2i_2 U168 ( .x(n1725), .a(reg_dst_of_MEM_2), .b(n1724) );
    inv_2 U1680 ( .x(n688), .a(n1371) );
    inv_2 U1681 ( .x(n1371), .a(WB_data[1]) );
    inv_2 U1682 ( .x(n689), .a(n1368) );
    inv_2 U1683 ( .x(n1368), .a(WB_data[5]) );
    inv_2 U1684 ( .x(n690), .a(n1366) );
    inv_2 U1685 ( .x(n1366), .a(WB_data[0]) );
    inv_2 U1686 ( .x(n691), .a(n1657) );
    inv_2 U1687 ( .x(n1657), .a(WB_data[6]) );
    inv_2 U1688 ( .x(n692), .a(n1385) );
    inv_2 U1689 ( .x(n1385), .a(WB_data[7]) );
    nor2_1 U169 ( .x(n1724), .a(reg_dst_of_MEM_0), .b(reg_dst_of_MEM_1) );
    buf_14 U1690 ( .x(reg_out_A[28]), .a(n3953) );
    buf_14 U1691 ( .x(reg_out_A[29]), .a(n3952) );
    inv_2 U1693 ( .x(n695), .a(n693) );
    nand2i_2 U1694 ( .x(n1161), .a(n587), .b(net150626) );
    nand2i_2 U1695 ( .x(n1181), .a(n586), .b(net150626) );
    nand2i_2 U1696 ( .x(n1165), .a(n589), .b(net150626) );
    nand2i_2 U1697 ( .x(n1149), .a(n583), .b(net150626) );
    nand2i_2 U1698 ( .x(n1169), .a(n573), .b(net150626) );
    nand2i_2 U1699 ( .x(n1225), .a(n591), .b(net150626) );
    inv_0 U17 ( .x(n1533), .a(NPC[21]) );
    nor2_1 U170 ( .x(n1726), .a(reg_dst_of_MEM_3), .b(reg_dst_of_MEM_4) );
    nand2i_2 U1700 ( .x(n1209), .a(n584), .b(net150626) );
    nand2i_2 U1701 ( .x(n1229), .a(n593), .b(net150626) );
    nand2i_2 U1702 ( .x(n1201), .a(n577), .b(net150626) );
    nand2i_2 U1703 ( .x(n1157), .a(n595), .b(net150626) );
    nand2i_2 U1704 ( .x(n1189), .a(n592), .b(net150626) );
    nand2i_2 U1705 ( .x(n1177), .a(n575), .b(net150626) );
    nand2i_2 U1706 ( .x(n1245), .a(n574), .b(net150626) );
    nand2i_2 U1707 ( .x(n1205), .a(n572), .b(net150626) );
    nand2i_2 U1708 ( .x(n1153), .a(n594), .b(net150626) );
    nand2i_2 U1709 ( .x(n1173), .a(n576), .b(net150626) );
    nand2i_2 U171 ( .x(n1089), .a(n559), .b(n642) );
    inv_5 U1711 ( .x(n1339), .a(N450) );
    inv_10 U1712 ( .x(n697), .a(n1431) );
    nand2i_8 U1713 ( .x(n1431), .a(n1432), .b(n1430) );
    inv_0 U1714 ( .x(n1096), .a(n1431) );
    and2_8 U1715 ( .x(net149679), .a(n780), .b(n787) );
    nand4i_4 U1716 ( .x(n1704), .a(n1372), .b(n1130), .c(n653), .d(n994) );
    nand4_5 U1718 ( .x(n1701), .a(n1024), .b(n1028), .c(n674), .d(n698) );
    inv_0 U1719 ( .x(n699), .a(n1347) );
    nand2i_2 U172 ( .x(n1072), .a(n560), .b(n1718) );
    inv_6 U1720 ( .x(n1009), .a(n1347) );
    mux2i_5 U1721 ( .x(n1347), .d0(n1348), .sl(___cell__36997_net129354), .d1(
        n1349) );
    nand3_4 U1722 ( .x(n1459), .a(n855), .b(n714), .c(n747) );
    nand4_5 U1723 ( .x(n1702), .a(n1026), .b(n998), .c(n1006), .d(n1009) );
    nand2i_0 U1724 ( .x(n1722), .a(n2634), .b(n1461) );
    nand2i_3 U1725 ( .x(n1143), .a(n1498), .b(n863) );
    nand4i_1 U1727 ( .x(n700), .a(n1456), .b(n1457), .c(n1458), .d(n1444) );
    inv_5 U1728 ( .x(n714), .a(n1455) );
    oai21_1 U1729 ( .x(N6723), .a(n653), .b(n995), .c(n1126) );
    mux2i_1 U173 ( .x(n3737), .d0(n565), .sl(___cell__36997_net130681), .d1(
        n1417) );
    exnor2_1 U1731 ( .x(___cell__36997_net129977), .a(n1427), .b(n3926) );
    exnor2_1 U1732 ( .x(n1562), .a(n1427), .b(n634) );
    exnor2_2 U1733 ( .x(n1695), .a(n1427), .b(n702) );
    nand2_6 U1734 ( .x(n756), .a(n822), .b(n1446) );
    inv_10 U1736 ( .x(___cell__36997_net125989), .a(___cell__36997_net129381)
         );
    inv_10 U1737 ( .x(___cell__36997_net125941), .a(___cell__36997_net129378)
         );
    aoi22_4 U1738 ( .x(n859), .a(n883), .b(n882), .c(n757), .d(n881) );
    inv_6 U1739 ( .x(n757), .a(n752) );
    mux2i_1 U174 ( .x(n3760), .d0(n566), .sl(___cell__36997_net130681), .d1(
        n1316) );
    exor2_5 U1740 ( .x(n1442), .a(reg_dst_of_EX_4), .b(n1132) );
    exnor2_6 U1741 ( .x(n1570), .a(n1571), .b(n708) );
    mux2i_2 U1743 ( .x(n702), .d0(rd_addr[3]), .sl(n703), .d1(rt_addr[3]) );
    nand2_0 U1744 ( .x(n1731), .a(n3998), .b(n1565) );
    exor2_1 U1745 ( .x(n1685), .a(n1686), .b(n1565) );
    nand2_3 U1747 ( .x(n1432), .a(n739), .b(n815) );
    nand2_8 U1749 ( .x(n705), .a(n704), .b(n1461) );
    mux2i_1 U175 ( .x(n3752), .d0(n567), .sl(___cell__36997_net130681), .d1(
        n1331) );
    inv_16 U1750 ( .x(n1461), .a(n1260) );
    nand2i_8 U1751 ( .x(n1428), .a(n1315), .b(n1111) );
    inv_0 U1752 ( .x(n707), .a(n683) );
    inv_2 U1753 ( .x(n708), .a(n707) );
    oai21_1 U1754 ( .x(N6718), .a(n3985), .b(___cell__36997_net130580), .c(
        n996) );
    inv_5 U1755 ( .x(n1337), .a(N443) );
    and2_8 U1756 ( .x(n709), .a(n710), .b(n1694) );
    nor3_2 U1757 ( .x(n710), .a(n333), .b(n715), .c(n761) );
    nand2_1 U1758 ( .x(n1434), .a(n739), .b(n850) );
    nand2_0 U1759 ( .x(n1516), .a(n724), .b(n683) );
    mux2i_1 U176 ( .x(n3747), .d0(n568), .sl(___cell__36997_net130681), .d1(
        n1412) );
    nand2i_3 U1761 ( .x(n1449), .a(n1446), .b(n822) );
    oai21_1 U1762 ( .x(N6721), .a(n673), .b(n1777), .c(n1238) );
    inv_6 U1763 ( .x(n769), .a(n736) );
    aoi21_1 U1764 ( .x(n1087), .a(rd_addr[2]), .b(n1718), .c(n1802) );
    aoi22_1 U1766 ( .x(n1141), .a(n1355), .b(n797), .c(EPC_28), .d(net150625)
         );
    mux2i_6 U1767 ( .x(n1355), .d0(n1356), .sl(___cell__36997_net129354), .d1(
        n1357) );
    nand2i_4 U1768 ( .x(n711), .a(n1429), .b(n753) );
    nand2i_4 U1769 ( .x(n752), .a(n1429), .b(n753) );
    mux2i_1 U177 ( .x(n3745), .d0(n570), .sl(___cell__36997_net130681), .d1(
        n1414) );
    aoi21_3 U1770 ( .x(n825), .a(n1737), .b(n826), .c(n1451) );
    inv_3 U1771 ( .x(n1500), .a(N5378) );
    aoi21_1 U1772 ( .x(n1075), .a(rd_addr[0]), .b(n1718), .c(n1802) );
    inv_0 U1773 ( .x(n807), .a(n1096) );
    inv_10 U1774 ( .x(n333), .a(n759) );
    mux2i_8 U1775 ( .x(n759), .d0(IR_latched_input[23]), .sl(n760), .d1(
        current_IR_23) );
    nor2i_2 U1776 ( .x(n1264), .a(n855), .b(n1265) );
    mux2i_8 U1777 ( .x(n712), .d0(n1318), .sl(n728), .d1(n1319) );
    and2_8 U1778 ( .x(n822), .a(n823), .b(n1437) );
    nand2i_0 U1779 ( .x(n713), .a(n1487), .b(n846) );
    mux2i_1 U178 ( .x(n3743), .d0(n571), .sl(___cell__36997_net130681), .d1(
        n1416) );
    inv_14 U1781 ( .x(n855), .a(n756) );
    nand4i_3 U1782 ( .x(n1455), .a(n1456), .b(n1457), .c(n1458), .d(n1444) );
    nand2_6 U1783 ( .x(___cell__36997_net129632), .a(n812), .b(net148863) );
    oai21_1 U1784 ( .x(N6731), .a(n1003), .b(n995), .c(n1004) );
    inv_8 U1785 ( .x(n1003), .a(n1404) );
    oai21_1 U1786 ( .x(N6719), .a(n1130), .b(n995), .c(n1131) );
    oai211_2 U1789 ( .x(n841), .a(n1081), .b(n843), .c(n767), .d(n724) );
    mux2i_1 U179 ( .x(n2647), .d0(n622), .sl(___cell__36997_net130567), .d1(
        n845) );
    oai21_1 U1790 ( .x(n3771), .a(n1081), .b(n1775), .c(n1082) );
    nand2i_1 U1791 ( .x(n1491), .a(n1688), .b(n1096) );
    inv_6 U1792 ( .x(n767), .a(n1688) );
    and2_1 U1794 ( .x(n812), .a(n1467), .b(n1688) );
    inv_10 U1795 ( .x(n1437), .a(n1435) );
    inv_2 U1796 ( .x(n717), .a(n1548) );
    inv_0 U1797 ( .x(n718), .a(n715) );
    inv_2 U1798 ( .x(n719), .a(n718) );
    inv_2 U1799 ( .x(n1445), .a(n855) );
    nor2_1 U18 ( .x(n1581), .a(IR_opcode_field[3]), .b(n1321) );
    mux2i_1 U180 ( .x(n2646), .d0(n623), .sl(___cell__36997_net130125), .d1(
        n871) );
    ao21_4 U1800 ( .x(n721), .a(n1737), .b(n861), .c(n755) );
    exor2_2 U1802 ( .x(n1560), .a(n1561), .b(n759) );
    aoi21_1 U1805 ( .x(n1080), .a(IR_function_field[5]), .b(n1718), .c(n1719)
         );
    inv_8 U1806 ( .x(n722), .a(N6376) );
    inv_16 U1807 ( .x(Imm[24]), .a(n722) );
    inv_3 U1808 ( .x(n1427), .a(n332) );
    mux2i_2 U181 ( .x(n3763), .d0(n633), .sl(___cell__36997_net130681), .d1(
        n725) );
    nand2_2 U1810 ( .x(n1137), .a(___cell__36997_net130709), .b(N5449) );
    nand2i_2 U1811 ( .x(n3810), .a(n1101), .b(n1100) );
    nand4_1 U1812 ( .x(n3853), .a(n1139), .b(n668), .c(n1138), .d(n1140) );
    inv_10 U1813 ( .x(n810), .a(NPC[3]) );
    inv_16 U1814 ( .x(n865), .a(NPC[2]) );
    inv_2 U1815 ( .x(n725), .a(n724) );
    inv_2 U1816 ( .x(n726), .a(n1543) );
    oai21_1 U1817 ( .x(N6722), .a(n636), .b(n1777), .c(n1127) );
    oai21_1 U1819 ( .x(N6729), .a(n998), .b(n1777), .c(n999) );
    inv_2 U182 ( .x(n1559), .a(reg_dst_of_EX_4) );
    nor2i_2 U1820 ( .x(n1694), .a(n879), .b(n3990) );
    nand2i_0 U1821 ( .x(n1730), .a(n3998), .b(n3990) );
    oai21_1 U1822 ( .x(n3783), .a(n1774), .b(n1059), .c(n1087) );
    oai21_1 U1823 ( .x(n3766), .a(n1774), .b(n1040), .c(n1079) );
    oai21_1 U1824 ( .x(n3768), .a(n1774), .b(n1043), .c(n1074) );
    oai21_1 U1825 ( .x(n3782), .a(n1774), .b(n1057), .c(n1069) );
    oai21_1 U1826 ( .x(n3786), .a(n856), .b(n1774), .c(n1077) );
    oai21_1 U1827 ( .x(n3789), .a(n772), .b(n1774), .c(n1122) );
    oai21_1 U1828 ( .x(n3773), .a(n3992), .b(n1774), .c(n1112) );
    oai21_1 U1829 ( .x(N6725), .a(n672), .b(n995), .c(n1243) );
    oai21_1 U183 ( .x(n3764), .a(n1065), .b(n1038), .c(n1078) );
    mux2i_8 U1830 ( .x(n1083), .d0(current_IR_30), .sl(net149679), .d1(
        IR_latched_input[30]) );
    nand2_1 U1831 ( .x(n2707), .a(n729), .b(n1134) );
    inv_2 U1832 ( .x(n729), .a(n742) );
    nor2i_2 U1833 ( .x(n1312), .a(n825), .b(n837) );
    inv_10 U1835 ( .x(n731), .a(n771) );
    inv_10 U1836 ( .x(___cell__36997_net130572), .a(n771) );
    or3i_1 U1837 ( .x(n2706), .a(n1134), .b(n1473), .c(n1090) );
    nand2i_6 U1838 ( .x(n1737), .a(n1689), .b(n1477) );
    nand2i_2 U184 ( .x(n1078), .a(n1859), .b(n642) );
    ao21_3 U1842 ( .x(n733), .a(net150625), .b(EPC_26), .c(n1280) );
    buf_10 U1843 ( .x(net150625), .a(n799) );
    nand2_0 U1844 ( .x(n1110), .a(n1718), .b(IR_opcode_field[5]) );
    mux2i_1 U1845 ( .x(n1479), .d0(n1585), .sl(IR_opcode_field[5]), .d1(n1582)
         );
    or3i_1 U1846 ( .x(n1438), .a(IR_opcode_field[3]), .b(IR_opcode_field[5]), 
        .c(IR_opcode_field[1]) );
    inv_10 U1848 ( .x(n738), .a(n791) );
    inv_10 U1849 ( .x(net148863), .a(n791) );
    mux2i_1 U185 ( .x(n3753), .d0(n646), .sl(___cell__36997_net126612), .d1(
        n1325) );
    mux2i_8 U1850 ( .x(n739), .d0(IR_latched_input[31]), .sl(net149236), .d1(
        current_IR_31) );
    nor2_4 U1851 ( .x(n1463), .a(n724), .b(n1578) );
    mux2i_8 U1852 ( .x(n761), .d0(n666), .sl(net149679), .d1(n1327) );
    inv_2 U1853 ( .x(n1327), .a(IR_latched_input[25]) );
    inv_16 U1855 ( .x(net149236), .a(___cell__36997_net130572) );
    nor2i_3 U1856 ( .x(n740), .a(n1590), .b(n741) );
    inv_5 U1857 ( .x(n741), .a(n1454) );
    inv_0 U1858 ( .x(n1591), .a(n1590) );
    oaoi211_1 U1859 ( .x(n742), .a(n745), .b(n744), .c(n743), .d(n883) );
    mux2i_1 U186 ( .x(n3735), .d0(n651), .sl(___cell__36997_net130681), .d1(
        n1420) );
    inv_2 U1860 ( .x(n743), .a(n1266) );
    inv_0 U1861 ( .x(n745), .a(n1461) );
    nor2i_0 U1862 ( .x(n1266), .a(n1267), .b(___cell__36997_net126612) );
    nand2_5 U1863 ( .x(n835), .a(___cell__36997_net130214), .b(N6023) );
    inv_16 U1864 ( .x(n811), .a(n810) );
    aoi22_2 U1865 ( .x(n1228), .a(N5361), .b(n863), .c(N6028), .d(
        ___cell__36997_net130713) );
    aoi22_2 U1866 ( .x(n1200), .a(N5355), .b(n863), .c(N6022), .d(
        ___cell__36997_net130713) );
    exor2_2 U1867 ( .x(n1696), .a(n1557), .b(n334) );
    inv_10 U1868 ( .x(n1565), .a(n334) );
    mux2i_1 U187 ( .x(n3744), .d0(n652), .sl(___cell__36997_net126612), .d1(
        n1415) );
    aoi222_1 U1871 ( .x(n1008), .a(NPC[16]), .b(n1802), .c(n1732), .d(EPC_16), 
        .e(Cause_Reg_16), .f(n1803) );
    inv_0 U1872 ( .x(n1538), .a(NPC[16]) );
    inv_7 U1873 ( .x(n1736), .a(n1459) );
    nand2i_1 U1875 ( .x(n1483), .a(n1476), .b(n1736) );
    nand2_5 U1876 ( .x(n1489), .a(n1736), .b(n1476) );
    nand4i_5 U1877 ( .x(n1440), .a(n1441), .b(n1444), .c(n1443), .d(n1442) );
    inv_2 U1878 ( .x(n746), .a(n1545) );
    and2_8 U1879 ( .x(n747), .a(n1440), .b(n1313) );
    inv_2 U188 ( .x(n1561), .a(reg_dst_of_EX_2) );
    inv_5 U1881 ( .x(n1517), .a(n711) );
    nor2_3 U1883 ( .x(n1697), .a(n748), .b(n1560) );
    inv_16 U1884 ( .x(n340), .a(n884) );
    inv_10 U1885 ( .x(n1523), .a(n1449) );
    inv_5 U1888 ( .x(n760), .a(net149681) );
    nand2_0 U1889 ( .x(n1084), .a(n642), .b(IR_opcode_field[4]) );
    mux2i_1 U189 ( .x(n3755), .d0(n659), .sl(___cell__36997_net126612), .d1(
        n1326) );
    nand2_1 U1890 ( .x(n1321), .a(IR_opcode_field[4]), .b(IR_opcode_field[2])
         );
    inv_3 U1891 ( .x(n1495), .a(N5382) );
    inv_6 U1892 ( .x(n753), .a(n1428) );
    aoi22_1 U1893 ( .x(n1174), .a(branch_address[5]), .b(n766), .c(N5424), .d(
        ___cell__36997_net130709) );
    aoi22_1 U1895 ( .x(n1182), .a(branch_address[17]), .b(n766), .c(N5436), 
        .d(___cell__36997_net130709) );
    aoi22_1 U1896 ( .x(n1216), .a(branch_address[15]), .b(n766), .c(N5434), 
        .d(___cell__36997_net130709) );
    aoi22_1 U1897 ( .x(n1214), .a(branch_address[13]), .b(n766), .c(N5432), 
        .d(___cell__36997_net130709) );
    aoi22_1 U1898 ( .x(n1190), .a(branch_address[11]), .b(n766), .c(N5430), 
        .d(___cell__36997_net130709) );
    aoi22_1 U1899 ( .x(n1154), .a(branch_address[1]), .b(n766), .c(N5420), .d(
        ___cell__36997_net130709) );
    nor2i_1 U19 ( .x(n1580), .a(n1439), .b(n1568) );
    mux2i_1 U190 ( .x(n3754), .d0(n661), .sl(___cell__36997_net130681), .d1(
        n1328) );
    aoi21_1 U1900 ( .x(n1178), .a(N5425), .b(___cell__36997_net130709), .c(
        n1268) );
    or3i_1 U1902 ( .x(n2705), .a(n1134), .b(n1473), .c(n1091) );
    nand2_5 U1903 ( .x(n1446), .a(n1447), .b(___cell__36997_net130306) );
    nand2i_5 U1904 ( .x(n1467), .a(n1468), .b(n1469) );
    inv_1 U1905 ( .x(n1468), .a(n1436) );
    nand4_1 U1906 ( .x(n3852), .a(n1142), .b(n665), .c(n1141), .d(n1143) );
    inv_2 U1907 ( .x(n755), .a(n1479) );
    exnor2_1 U1908 ( .x(n1693), .a(reg_dst_of_EX_2), .b(n338) );
    inv_8 U1909 ( .x(n998), .a(n1352) );
    oai21_1 U191 ( .x(n3769), .a(n1775), .b(n1044), .c(n1080) );
    inv_8 U1910 ( .x(n804), .a(n879) );
    buf_16 U1911 ( .x(Imm[3]), .a(N6334) );
    nand2i_2 U1912 ( .x(n1219), .a(n1006), .b(n797) );
    inv_8 U1913 ( .x(n1006), .a(n1350) );
    mux2i_8 U1915 ( .x(n768), .d0(IR_latched_input[22]), .sl(n769), .d1(n660)
         );
    nand2i_2 U1916 ( .x(n1183), .a(n699), .b(n797) );
    oai21_1 U1917 ( .x(N6735), .a(n699), .b(n1777), .c(n1010) );
    oai21_1 U1918 ( .x(N6732), .a(___cell__36997_net125941), .b(n1777), .c(
        n1005) );
    nand2i_2 U1919 ( .x(n1167), .a(___cell__36997_net125941), .b(n797) );
    mux2i_1 U192 ( .x(n3757), .d0(n666), .sl(___cell__36997_net126612), .d1(
        n1327) );
    oai21_1 U1920 ( .x(N6733), .a(n1006), .b(___cell__36997_net130580), .c(
        n1007) );
    oai21_1 U1921 ( .x(N6734), .a(n663), .b(n995), .c(n1008) );
    nand2i_2 U1922 ( .x(n1163), .a(n663), .b(n797) );
    mux2i_6 U1923 ( .x(n1341), .d0(n1342), .sl(___cell__36997_net129354), .d1(
        n1343) );
    nand2i_5 U1924 ( .x(n1106), .a(n1487), .b(n846) );
    nand2i_0 U1925 ( .x(n1085), .a(n1488), .b(n846) );
    inv_10 U1926 ( .x(n846), .a(n841) );
    mux2i_8 U1927 ( .x(n832), .d0(n1418), .sl(n777), .d1(n1419) );
    aoi21_2 U1928 ( .x(n1222), .a(N6036), .b(___cell__36997_net130713), .c(
        n1295) );
    mux2i_3 U1929 ( .x(n338), .d0(n1334), .sl(net149680), .d1(n1335) );
    mux2i_1 U193 ( .x(n3901), .d0(n1672), .sl(n1650), .d1(n1379) );
    inv_2 U1930 ( .x(n1335), .a(IR_latched_input[18]) );
    aoi22_3 U1931 ( .x(n1212), .a(N5364), .b(n862), .c(N6031), .d(
        ___cell__36997_net130713) );
    inv_16 U1932 ( .x(n862), .a(n1272) );
    exor2_1 U1933 ( .x(n1566), .a(reg_dst_of_MEM_0), .b(n884) );
    exor2_1 U1934 ( .x(n1575), .a(WB_index_0), .b(n856) );
    inv_10 U1935 ( .x(n1477), .a(n1448) );
    nand2_8 U1936 ( .x(n1448), .a(n1106), .b(n1108) );
    mux2i_8 U1937 ( .x(n896), .d0(n1328), .sl(net152024), .d1(n661) );
    inv_2 U1938 ( .x(net152025), .a(net152024) );
    nand2_8 U1939 ( .x(n1429), .a(n716), .b(n1688) );
    inv_2 U194 ( .x(n1672), .a(N514) );
    nand2i_4 U1940 ( .x(n1236), .a(n1508), .b(n862) );
    inv_16 U1941 ( .x(n797), .a(___cell__36997_net129632) );
    or2_3 U1943 ( .x(n758), .a(net151343), .b(n662) );
    inv_0 U1944 ( .x(net151343), .a(n799) );
    and2_6 U1945 ( .x(n867), .a(n868), .b(net148863) );
    mux2i_5 U1946 ( .x(n772), .d0(IR_latched_input[19]), .sl(n760), .d1(
        current_IR_19) );
    inv_2 U1947 ( .x(n1016), .a(n1372) );
    or2_4 U1948 ( .x(n1100), .a(n1733), .b(n1037) );
    or2_8 U1949 ( .x(n764), .a(n1733), .b(n1037) );
    mux2i_1 U195 ( .x(n3922), .d0(n1649), .sl(n1650), .d1(n1366) );
    or2_8 U1950 ( .x(n763), .a(n1733), .b(n1037) );
    nand2i_2 U1951 ( .x(n1733), .a(n1309), .b(n887) );
    oai21_5 U1952 ( .x(n1037), .a(n1484), .b(n1480), .c(n1554) );
    inv_3 U1953 ( .x(n1497), .a(N6047) );
    oai21_1 U1955 ( .x(n1804), .a(___cell__36997_net129624), .b(
        ___cell__36997_net129625), .c(___cell__36997_net130681) );
    mux2i_8 U1956 ( .x(n332), .d0(n1324), .sl(net149236), .d1(n1323) );
    oai21_1 U1957 ( .x(n3777), .a(n1094), .b(n1085), .c(n1098) );
    nand2i_2 U1958 ( .x(n1094), .a(___cell__36997_net127190), .b(n1480) );
    oai21_1 U1959 ( .x(n3772), .a(n1113), .b(n1065), .c(n1114) );
    inv_2 U196 ( .x(n1649), .a(N535) );
    oai21_1 U1960 ( .x(n1488), .a(n1081), .b(n1113), .c(n3992) );
    aoi22_2 U1961 ( .x(n1152), .a(N5352), .b(n895), .c(N6019), .d(
        ___cell__36997_net130214) );
    mux2i_8 U1964 ( .x(IR_latched_1), .d0(n801), .sl(net149236), .d1(n800) );
    buf_10 U1965 ( .x(reg_out_A[22]), .a(n3959) );
    ao22_6 U1968 ( .x(___cell__36997_net129524), .a(n721), .b(n1523), .c(n855), 
        .d(n740) );
    mux2i_1 U197 ( .x(n3911), .d0(n1662), .sl(n1650), .d1(n1354) );
    or2_8 U1970 ( .x(n771), .a(n3949), .b(n3950) );
    mux2i_1 U1971 ( .x(n3750), .d0(n1334), .sl(___cell__36997_net126612), .d1(
        n1335) );
    inv_2 U1972 ( .x(n1334), .a(current_IR_18) );
    inv_10 U1973 ( .x(n337), .a(n772) );
    inv_0 U1974 ( .x(n1329), .a(IR_latched_input[19]) );
    buf_16 U1975 ( .x(reg_out_A[9]), .a(n3969) );
    oai21_1 U1976 ( .x(n773), .a(n1317), .b(n847), .c(n1688) );
    inv_0 U1978 ( .x(n842), .a(n1688) );
    inv_2 U198 ( .x(n1662), .a(N524) );
    inv_4 U1980 ( .x(counter[1]), .a(n780) );
    oai21_4 U1981 ( .x(n1065), .a(n1484), .b(n1480), .c(
        ___cell__36997_net130681) );
    oai21_4 U1982 ( .x(n1775), .a(n1484), .b(n1480), .c(
        ___cell__36997_net126612) );
    oai21_4 U1983 ( .x(n1774), .a(n1484), .b(n1480), .c(
        ___cell__36997_net130681) );
    oai21_2 U1984 ( .x(n854), .a(n1484), .b(n1480), .c(n1554) );
    nor2i_0 U1985 ( .x(n1268), .a(branch_address[6]), .b(n738) );
    oai21_1 U1986 ( .x(n1237), .a(n738), .b(n1722), .c(
        ___cell__36997_net126604) );
    nor2i_0 U1987 ( .x(n1278), .a(branch_address[29]), .b(n738) );
    mux2i_1 U1988 ( .x(n1598), .d0(n2633), .sl(n738), .d1(n1471) );
    nor2i_0 U1989 ( .x(n1280), .a(branch_address[26]), .b(n738) );
    inv_2 U199 ( .x(n1499), .a(N5446) );
    inv_0 U1991 ( .x(n776), .a(net149680) );
    inv_2 U1992 ( .x(n777), .a(n776) );
    aoi22_2 U1993 ( .x(n1147), .a(branch_address[27]), .b(n766), .c(N6045), 
        .d(___cell__36997_net130713) );
    inv_14 U1994 ( .x(___cell__36997_net130713), .a(___cell__36997_net129239)
         );
    nor2i_1 U1995 ( .x(n1300), .a(N6029), .b(___cell__36997_net129239) );
    inv_2 U1997 ( .x(n783), .a(___cell__36997_net129247) );
    nand4_1 U1998 ( .x(n3842), .a(n1222), .b(n784), .c(n1223), .d(n1221) );
    inv_5 U1999 ( .x(n784), .a(n1220) );
    inv_4 U20 ( .x(n1067), .a(n850) );
    mux2i_1 U200 ( .x(n3902), .d0(n1671), .sl(n1650), .d1(n1381) );
    nand2i_4 U2000 ( .x(n1490), .a(n785), .b(n1699) );
    inv_3 U2001 ( .x(n785), .a(n855) );
    exnor2_3 U2002 ( .x(n1684), .a(n655), .b(n333) );
    mux2i_3 U2003 ( .x(n818), .d0(n773), .sl(n1578), .d1(n3989) );
    aoi222_1 U2004 ( .x(n1007), .a(NPC[15]), .b(n1719), .c(n1732), .d(EPC_15), 
        .e(Cause_Reg_15), .f(n1803) );
    inv_0 U2005 ( .x(n1539), .a(NPC[15]) );
    oaoi211_1 U2006 ( .x(_counter_reg_0_net48671), .a(___cell__36997_net127189
        ), .b(___cell__36997_net127190), .c(n777), .d(counter[0]) );
    nor2i_0 U2007 ( .x(_counter_reg_1_net48651), .a(n790), .b(n4011) );
    buf_1 U2008 ( .x(n790), .a(counter[1]) );
    nand2i_8 U2009 ( .x(___cell__36997_net129247), .a(___cell__36997_net129626
        ), .b(n738) );
    inv_2 U201 ( .x(n1671), .a(N515) );
    oai21_6 U2010 ( .x(n791), .a(___cell__36997_net129624), .b(
        ___cell__36997_net129625), .c(___cell__36997_net130681) );
    inv_16 U2011 ( .x(___cell__36997_net130681), .a(___cell__36997_net127190)
         );
    inv_10 U2012 ( .x(___cell__36997_net130214), .a(___cell__36997_net129239)
         );
    buf_16 U2014 ( .x(net150626), .a(n799) );
    inv_16 U2015 ( .x(___cell__36997_net129354), .a(n798) );
    exor2_3 U2017 ( .x(n795), .a(___cell__6171_net27367), .b(
        ___cell__36997_net129477) );
    inv_0 U2018 ( .x(___cell__36997_net126621), .a(IR_latched_1) );
    inv_10 U2019 ( .x(n1578), .a(n1111) );
    nor2i_1 U202 ( .x(n1109), .a(n1717), .b(n1485) );
    buf_16 U2020 ( .x(n802), .a(n1258) );
    oai21_1 U2021 ( .x(n3774), .a(n842), .b(n1775), .c(n1084) );
    mux2i_1 U2022 ( .x(n3762), .d0(n658), .sl(___cell__36997_net126612), .d1(
        n842) );
    and4i_1 U2023 ( .x(n1309), .a(n1310), .b(n842), .c(n725), .d(n683) );
    nand2_6 U2024 ( .x(n1435), .a(n859), .b(n1436) );
    buf_16 U2026 ( .x(reg_out_A[26]), .a(n3955) );
    buf_14 U2027 ( .x(n878), .a(n889) );
    inv_2 U2028 ( .x(n808), .a(n807) );
    inv_2 U2029 ( .x(n1496), .a(N6048) );
    oai21_1 U203 ( .x(n3780), .a(n1775), .b(n1108), .c(n1109) );
    inv_7 U2030 ( .x(n809), .a(n1051) );
    inv_10 U2031 ( .x(IR_latched_8), .a(n1049) );
    aoi222_1 U2032 ( .x(n1010), .a(NPC[17]), .b(n1719), .c(n1732), .d(EPC_17), 
        .e(Cause_Reg_17), .f(n1803) );
    inv_0 U2033 ( .x(n1537), .a(NPC[17]) );
    nand2_8 U2035 ( .x(___cell__36997_net127155), .a(net148863), .b(n1492) );
    aoi22_1 U2036 ( .x(n1240), .a(branch_address[3]), .b(n766), .c(N6021), .d(
        ___cell__36997_net130713) );
    nand2i_2 U2037 ( .x(n1140), .a(n1497), .b(___cell__36997_net130713) );
    nand2i_2 U2038 ( .x(n1198), .a(n1505), .b(___cell__36997_net130713) );
    nand2i_2 U2039 ( .x(n1217), .a(n1510), .b(___cell__36997_net130713) );
    oai21_1 U204 ( .x(n3767), .a(n1065), .b(n1041), .c(n1073) );
    aoi22_1 U2040 ( .x(n1255), .a(branch_address[2]), .b(net148865), .c(N6020), 
        .d(___cell__36997_net130713) );
    nand2i_2 U2041 ( .x(n1250), .a(n1501), .b(___cell__36997_net130713) );
    nand2i_2 U2043 ( .x(n1194), .a(n1507), .b(___cell__36997_net130713) );
    nand2i_2 U2044 ( .x(n1136), .a(n1496), .b(___cell__36997_net130713) );
    nor2_3 U2046 ( .x(n1293), .a(net148916), .b(n1294) );
    nor2_3 U2047 ( .x(n1275), .a(net148916), .b(n1276) );
    nor2_4 U2048 ( .x(n1282), .a(net148916), .b(n1283) );
    inv_3 U2049 ( .x(net150785), .a(net148916) );
    nand2i_2 U205 ( .x(n1073), .a(n1862), .b(n1718) );
    inv_14 U2050 ( .x(net148916), .a(___cell__36997_net130217) );
    mux2i_1 U2051 ( .x(n849), .d0(current_IR_3), .sl(n731), .d1(
        IR_latched_input[3]) );
    inv_0 U2052 ( .x(n1546), .a(NPC[8]) );
    aoi222_1 U2053 ( .x(n1032), .a(NPC[8]), .b(n1802), .c(n1732), .d(EPC_8), 
        .e(Cause_Reg_8), .f(n1803) );
    inv_0 U2054 ( .x(n1551), .a(n866) );
    aoi222_1 U2055 ( .x(n1253), .a(n737), .b(n1719), .c(n1732), .d(EPC_2), .e(
        Cause_Reg_2), .f(n1803) );
    mux2i_1 U2056 ( .x(n1091), .d0(n1588), .sl(slot_num_0), .d1(n1589) );
    exnor2_1 U2057 ( .x(n1314), .a(slot_num_1), .b(slot_num_0) );
    nand2i_0 U2058 ( .x(n1267), .a(slot_num_1), .b(slot_num_0) );
    nand2_2 U2059 ( .x(n1576), .a(slot_num_1), .b(slot_num_0) );
    inv_2 U206 ( .x(n1059), .a(IR_latched_13) );
    nor2i_1 U2060 ( .x(n1714), .a(slot_num_0), .b(n557) );
    buf_16 U2061 ( .x(reg_out_A[5]), .a(n3972) );
    inv_0 U2062 ( .x(n1047), .a(n817) );
    inv_0 U2064 ( .x(n820), .a(n809) );
    buf_16 U2065 ( .x(Imm[7]), .a(N6342) );
    inv_2 U2066 ( .x(n861), .a(n1438) );
    mux2i_1 U2067 ( .x(n3758), .d0(n852), .sl(___cell__36997_net130681), .d1(
        n1067) );
    oai21_1 U2068 ( .x(n3770), .a(n1067), .b(n1774), .c(n1068) );
    inv_5 U2069 ( .x(n1426), .a(n333) );
    oai21_1 U207 ( .x(n3781), .a(n1775), .b(n1055), .c(n1075) );
    nor2_0 U2070 ( .x(n1519), .a(n1730), .b(n1425) );
    nor2_0 U2071 ( .x(n1521), .a(n1731), .b(n1425) );
    nand2i_0 U2072 ( .x(n1712), .a(___cell__36997_net125928), .b(n1713) );
    inv_10 U2073 ( .x(n1713), .a(n1467) );
    inv_2 U2074 ( .x(n826), .a(n1474) );
    inv_5 U2075 ( .x(n1475), .a(n1451) );
    nand2i_2 U2076 ( .x(n1474), .a(opcode_of_MEM_1), .b(n1690) );
    nand2_1 U2077 ( .x(n1487), .a(n1578), .b(n1113) );
    nand2_0 U2078 ( .x(n1310), .a(n1578), .b(n1113) );
    nand3_0 U2079 ( .x(n1425), .a(n1426), .b(n1427), .c(
        ___cell__36997_net129477) );
    nand2i_2 U208 ( .x(n1039), .a(n720), .b(n1718) );
    ao21_1 U2081 ( .x(n2708), .a(___cell__36997_net130681), .b(n1035), .c(
        n1036) );
    and3i_5 U2082 ( .x(n834), .a(net151366), .b(n1489), .c(n1490) );
    inv_0 U2083 ( .x(n1035), .a(n834) );
    inv_10 U2084 ( .x(net151366), .a(___cell__36997_net127189) );
    inv_10 U2085 ( .x(___cell__36997_net127189), .a(___cell__36997_net129524)
         );
    inv_0 U2087 ( .x(n836), .a(n840) );
    inv_3 U2088 ( .x(n840), .a(n1462) );
    mux2i_6 U2089 ( .x(reg_dst_of_EX_2), .d0(n559), .sl(reg_dst), .d1(n670) );
    nor2_1 U209 ( .x(n1104), .a(n1776), .b(n654) );
    inv_0 U2090 ( .x(n1044), .a(n888) );
    inv_0 U2091 ( .x(n1308), .a(NPC[6]) );
    oai21_1 U2092 ( .x(n3776), .a(n1094), .b(n713), .c(n1107) );
    inv_0 U2093 ( .x(n1095), .a(n713) );
    buf_16 U2094 ( .x(Imm[21]), .a(N6370) );
    ao221_4 U2095 ( .x(n1689), .a(n1430), .b(n846), .c(n818), .d(n739), .e(
        n840) );
    nand3i_3 U2096 ( .x(n1462), .a(n712), .b(n1463), .c(n1464) );
    inv_10 U2097 ( .x(n1430), .a(n1428) );
    mux2i_8 U2098 ( .x(n1317), .d0(n1318), .sl(n728), .d1(n1319) );
    exor2_2 U2099 ( .x(n1567), .a(n1088), .b(reg_dst_of_MEM_2) );
    buf_14 U21 ( .x(Imm[9]), .a(N6346) );
    nand2i_2 U210 ( .x(n3815), .a(n1104), .b(n763) );
    exor2_1 U2100 ( .x(n1574), .a(WB_index_2), .b(n1088) );
    oai21_1 U2101 ( .x(n3788), .a(n3986), .b(n1065), .c(n1089) );
    nand4_5 U2102 ( .x(n1444), .a(n1088), .b(n1071), .c(n1691), .d(n1132) );
    buf_14 U2104 ( .x(n888), .a(IR_latched_5) );
    aoi22_1 U2105 ( .x(n1138), .a(n1341), .b(n797), .c(EPC_29), .d(net150625)
         );
    aoi222_1 U2106 ( .x(n1004), .a(NPC[13]), .b(n1719), .c(n1732), .d(EPC_13), 
        .e(Cause_Reg_13), .f(n1803) );
    inv_0 U2107 ( .x(n1541), .a(NPC[13]) );
    oai31_1 U2108 ( .x(n3779), .a(n1094), .b(n1095), .c(n808), .d(n1097) );
    nand2_6 U2109 ( .x(n1469), .a(n1466), .b(n808) );
    mux2i_1 U211 ( .x(n3892), .d0(n1681), .sl(n1650), .d1(n1363) );
    nand2i_8 U2110 ( .x(n1436), .a(n1067), .b(n697) );
    aoi222_1 U2111 ( .x(n1011), .a(NPC[18]), .b(n1802), .c(n1732), .d(EPC_18), 
        .e(Cause_Reg_18), .f(n1803) );
    inv_0 U2112 ( .x(n1055), .a(IR_latched_11) );
    aoi21_2 U2113 ( .x(n1172), .a(N5356), .b(n862), .c(n1270) );
    nand4_1 U2114 ( .x(n3847), .a(n1193), .b(n1192), .c(n1194), .d(n1195) );
    nand4_3 U2115 ( .x(n1571), .a(n1711), .b(n1708), .c(n1705), .d(n1703) );
    buf_16 U2116 ( .x(Imm[26]), .a(N6380) );
    aoi22_2 U2117 ( .x(n1218), .a(N5366), .b(n895), .c(EPC_15), .d(net150625)
         );
    buf_16 U2118 ( .x(reg_out_A[10]), .a(n3968) );
    nand3i_1 U2119 ( .x(n3823), .a(n1237), .b(net148916), .c(n1134) );
    inv_2 U212 ( .x(n1681), .a(N505) );
    mux2i_8 U2120 ( .x(n850), .d0(n851), .sl(net149236), .d1(n852) );
    nand4i_2 U2121 ( .x(n3827), .a(n1239), .b(n1240), .c(n1241), .d(n1242) );
    nand4i_2 U2122 ( .x(n3826), .a(n1254), .b(n1255), .c(n1256), .d(n1257) );
    mux2i_8 U2123 ( .x(IR_latched_12), .d0(n1415), .sl(net149236), .d1(n652)
         );
    nor2_4 U2125 ( .x(n1284), .a(net148913), .b(n1285) );
    inv_0 U2126 ( .x(n1549), .a(NPC[4]) );
    aoi222_1 U2127 ( .x(n1127), .a(NPC[4]), .b(n1719), .c(n1732), .d(EPC_4), 
        .e(Cause_Reg_4), .f(n1803) );
    aoi222_1 U2128 ( .x(n1005), .a(NPC[14]), .b(n1802), .c(n1732), .d(EPC_14), 
        .e(Cause_Reg_14), .f(n1803) );
    inv_0 U2129 ( .x(n1540), .a(NPC[14]) );
    or2_4 U213 ( .x(n665), .a(___cell__36997_net129247), .b(n1279) );
    aoi222_1 U2130 ( .x(n1238), .a(n811), .b(n1802), .c(n1732), .d(EPC_3), .e(
        Cause_Reg_3), .f(n1803) );
    inv_0 U2131 ( .x(n1550), .a(n811) );
    nand2i_2 U2132 ( .x(n1482), .a(n721), .b(n1523) );
    mux2i_2 U2133 ( .x(n1315), .d0(n566), .sl(n731), .d1(n1316) );
    inv_5 U2134 ( .x(n857), .a(n856) );
    inv_0 U2135 ( .x(n1544), .a(NPC[10]) );
    aoi222_1 U2136 ( .x(n997), .a(NPC[10]), .b(n1802), .c(n1732), .d(EPC_10), 
        .e(Cause_Reg_10), .f(n1803) );
    nand2i_1 U2137 ( .x(n1192), .a(n1018), .b(n797) );
    nand2i_1 U2138 ( .x(n1196), .a(n1020), .b(n797) );
    nand2i_1 U2139 ( .x(n1235), .a(n1016), .b(n797) );
    inv_2 U214 ( .x(n1279), .a(N5447) );
    nand2i_1 U2140 ( .x(n1150), .a(n640), .b(n797) );
    nand2i_1 U2141 ( .x(n1233), .a(n1014), .b(n797) );
    nand2i_1 U2142 ( .x(n1191), .a(n998), .b(n797) );
    nand2i_1 U2143 ( .x(n1159), .a(n3985), .b(n797) );
    nand2i_1 U2144 ( .x(n1247), .a(n672), .b(n797) );
    nand2i_1 U2145 ( .x(n1175), .a(n653), .b(n797) );
    nand2i_1 U2146 ( .x(n1179), .a(n1128), .b(n797) );
    nand2i_2 U2147 ( .x(n1257), .a(n1252), .b(n797) );
    nand2i_2 U2148 ( .x(n1242), .a(n673), .b(n797) );
    nand2i_2 U2149 ( .x(n1223), .a(n674), .b(n797) );
    mux2i_1 U215 ( .x(n3913), .d0(n1660), .sl(n1650), .d1(n1411) );
    nand2i_1 U2150 ( .x(n1203), .a(n636), .b(n797) );
    nand2i_1 U2151 ( .x(n1171), .a(n1031), .b(n797) );
    nand2i_1 U2152 ( .x(n1215), .a(n1003), .b(n797) );
    nand2i_1 U2153 ( .x(n1231), .a(n638), .b(n797) );
    nand2i_1 U2154 ( .x(n1211), .a(n639), .b(n797) );
    nand2i_1 U2155 ( .x(n1155), .a(n1130), .b(n797) );
    nand2i_1 U2156 ( .x(n1227), .a(n1001), .b(n797) );
    nand2i_1 U2157 ( .x(n1207), .a(n637), .b(n797) );
    aoi22_1 U2158 ( .x(n1248), .a(___cell__36997_net129381), .b(n797), .c(
        N5445), .d(___cell__36997_net130709) );
    buf_16 U2159 ( .x(reg_out_A[25]), .a(n3956) );
    inv_2 U216 ( .x(n1660), .a(N526) );
    aoi22_1 U2160 ( .x(n860), .a(n883), .b(n882), .c(n1517), .d(n881) );
    nand4_1 U2161 ( .x(n3845), .a(n1232), .b(n675), .c(n1233), .d(n1234) );
    oai22_1 U2162 ( .x(n3791), .a(n705), .b(n813), .c(n854), .d(n1038) );
    oai21_1 U2163 ( .x(n3792), .a(n3995), .b(___cell__36997_net126621), .c(
        n1039) );
    oai22_1 U2164 ( .x(n3793), .a(n1776), .b(n870), .c(n3995), .d(n1040) );
    oai21_1 U2165 ( .x(n3794), .a(n3995), .b(n1041), .c(n1042) );
    oai22_1 U2167 ( .x(n3796), .a(n1776), .b(n845), .c(n3995), .d(n1044) );
    oai21_1 U2168 ( .x(n3797), .a(n1045), .b(n3995), .c(n1046) );
    oai21_1 U2169 ( .x(n3798), .a(n1047), .b(n3995), .c(n1048) );
    inv_2 U217 ( .x(n1680), .a(N506) );
    oai21_1 U2170 ( .x(n3799), .a(n1049), .b(n3995), .c(n1050) );
    oai21_1 U2171 ( .x(n3800), .a(n820), .b(n3995), .c(n1052) );
    oai21_1 U2172 ( .x(n3803), .a(n1057), .b(n854), .c(n1058) );
    oai21_1 U2173 ( .x(n3804), .a(n1059), .b(n854), .c(n1060) );
    oai21_1 U2174 ( .x(n3806), .a(n1063), .b(n3995), .c(n1064) );
    oai21_1 U2175 ( .x(n3805), .a(n1061), .b(n854), .c(n1062) );
    inv_16 U2176 ( .x(n863), .a(n1272) );
    inv_16 U2177 ( .x(n1272), .a(n867) );
    mux2i_8 U2178 ( .x(IR_latched_0), .d0(n1423), .sl(net149681), .d1(n1424)
         );
    inv_16 U2179 ( .x(n866), .a(n865) );
    mux2i_1 U218 ( .x(n3893), .d0(n1680), .sl(n1650), .d1(n1343) );
    inv_2 U2180 ( .x(n868), .a(n1493) );
    nand2i_0 U2181 ( .x(n1493), .a(n1688), .b(n1468) );
    mux2i_1 U2182 ( .x(___cell__36997_net129654), .d0(n2632), .sl(n738), .d1(
        n1471) );
    buf_16 U2184 ( .x(Imm[20]), .a(N6368) );
    buf_16 U2185 ( .x(Imm[11]), .a(N6350) );
    buf_8 U2186 ( .x(n889), .a(n338) );
    mux2i_8 U2187 ( .x(n339), .d0(n1332), .sl(net149681), .d1(n1333) );
    mux2i_3 U2189 ( .x(reg_dst_of_EX_0), .d0(n561), .sl(reg_dst), .d1(n669) );
    mux2i_1 U219 ( .x(n3897), .d0(n1676), .sl(n1650), .d1(n1338) );
    mux2i_3 U2190 ( .x(reg_dst_of_EX_4), .d0(n558), .sl(reg_dst), .d1(n562) );
    inv_5 U2192 ( .x(n882), .a(n1433) );
    nand2i_2 U2193 ( .x(n1433), .a(CLI), .b(INT) );
    nand2_0 U2194 ( .x(n1717), .a(n642), .b(reg_dst) );
    inv_0 U2196 ( .x(n1543), .a(NPC[11]) );
    aoi222_1 U2197 ( .x(n999), .a(n726), .b(n1719), .c(n1732), .d(EPC_11), .e(
        Cause_Reg_11), .f(n1803) );
    mux2i_1 U2199 ( .x(IR_latched_15), .d0(n568), .sl(net149680), .d1(n1412)
         );
    nor3_1 U22 ( .x(n1579), .a(n3923), .b(opcode_of_MEM_3), .c(opcode_of_MEM_4
        ) );
    inv_2 U220 ( .x(n1676), .a(N510) );
    inv_0 U2200 ( .x(n1063), .a(n887) );
    oai21_1 U2201 ( .x(N6744), .a(___cell__36997_net125989), .b(n1777), .c(
        n1023) );
    nand2i_2 U2202 ( .x(___cell__36997_net129657), .a(n1495), .b(n867) );
    nand2i_2 U2203 ( .x(n1146), .a(n1500), .b(n863) );
    nand2i_2 U2204 ( .x(n1187), .a(n1503), .b(n862) );
    nand2i_2 U2205 ( .x(n1199), .a(n1504), .b(n863) );
    nand2i_2 U2206 ( .x(n1251), .a(n1502), .b(n862) );
    aoi21_1 U2208 ( .x(n1180), .a(N5368), .b(n863), .c(n1297) );
    aoi21_1 U2209 ( .x(n1188), .a(N5362), .b(n863), .c(n1300) );
    nand2i_2 U2210 ( .x(n1195), .a(n1506), .b(n862) );
    aoi21_1 U2211 ( .x(n1156), .a(N5351), .b(n863), .c(n1301) );
    nand2i_2 U2213 ( .x(n1234), .a(n1509), .b(n863) );
    aoi21_3 U2214 ( .x(n1256), .a(N5353), .b(n862), .c(n1293) );
    aoi21_3 U2215 ( .x(n1241), .a(N5354), .b(n863), .c(n1275) );
    aoi22_1 U2217 ( .x(n1168), .a(N5359), .b(n895), .c(N6026), .d(
        ___cell__36997_net130214) );
    aoi22_1 U2218 ( .x(n1160), .a(N5367), .b(n895), .c(N6034), .d(
        ___cell__36997_net130214) );
    aoi22_1 U2219 ( .x(n1224), .a(N5363), .b(n895), .c(N6030), .d(
        ___cell__36997_net130214) );
    mux2i_1 U222 ( .x(n1090), .d0(n1587), .sl(___cell__36997_net126612), .d1(
        n883) );
    aoi22_1 U2221 ( .x(n1151), .a(N5371), .b(n895), .c(N6038), .d(
        ___cell__36997_net130214) );
    oai21_1 U2222 ( .x(n3801), .a(n1053), .b(n3995), .c(n1054) );
    oai21_1 U2223 ( .x(n3775), .a(n725), .b(n1065), .c(n1110) );
    inv_0 U2224 ( .x(n1545), .a(NPC[9]) );
    aoi222_1 U2225 ( .x(n1033), .a(n746), .b(n1719), .c(n1732), .d(EPC_9), .e(
        Cause_Reg_9), .f(n1803) );
    mux2i_1 U2226 ( .x(IR_latched_5), .d0(n565), .sl(n731), .d1(n1417) );
    oai21_1 U2227 ( .x(N6745), .a(n1024), .b(n678), .c(n1025) );
    inv_0 U2228 ( .x(n1547), .a(NPC[7]) );
    aoi222_1 U2229 ( .x(n1243), .a(n554), .b(n1719), .c(n1732), .d(EPC_7), .e(
        Cause_Reg_7), .f(n1803) );
    mux2i_1 U223 ( .x(n3910), .d0(n1663), .sl(n1650), .d1(n1400) );
    inv_0 U2230 ( .x(n1542), .a(NPC[12]) );
    aoi222_1 U2231 ( .x(n1002), .a(NPC[12]), .b(n1802), .c(n1732), .d(EPC_12), 
        .e(Cause_Reg_12), .f(n1803) );
    buf_16 U2232 ( .x(reg_out_A[24]), .a(n3957) );
    exor2_1 U2233 ( .x(n1568), .a(IR_opcode_field[2]), .b(IR_opcode_field[4])
         );
    nand2i_2 U2234 ( .x(n3812), .a(n1118), .b(n763) );
    buf_16 U2235 ( .x(Imm[28]), .a(N6384) );
    oai21_1 U2236 ( .x(N6743), .a(n698), .b(n995), .c(n1022) );
    nand2i_2 U2237 ( .x(n3809), .a(n1120), .b(n1100) );
    oai21_1 U2238 ( .x(n3802), .a(n1055), .b(n854), .c(n1056) );
    inv_0 U2239 ( .x(n1548), .a(NPC[5]) );
    inv_2 U224 ( .x(n1663), .a(N523) );
    aoi222_1 U2240 ( .x(n1126), .a(n717), .b(n1802), .c(n1732), .d(EPC_5), .e(
        Cause_Reg_5), .f(n1803) );
    inv_7 U2242 ( .x(net148915), .a(___cell__36997_net130217) );
    nand2_0 U2243 ( .x(n1112), .a(n1718), .b(IR_opcode_field[3]) );
    inv_0 U2244 ( .x(n1322), .a(IR_opcode_field[3]) );
    nor2_0 U2245 ( .x(n1700), .a(IR_opcode_field[3]), .b(IR_opcode_field[4])
         );
    nand4i_1 U2247 ( .x(n1773), .a(n1734), .b(n1572), .c(n1735), .d(n1444) );
    oai21_1 U2248 ( .x(n3787), .a(n1071), .b(n1775), .c(n1072) );
    exor2_1 U2249 ( .x(n1687), .a(n1686), .b(n1071) );
    buf_16 U2250 ( .x(Imm[17]), .a(N6362) );
    buf_16 U2251 ( .x(Imm[15]), .a(N6358) );
    aoi221_1 U2252 ( .x(n1232), .a(N5440), .b(___cell__36997_net130212), .c(
        branch_address[21]), .d(net148865), .e(n1290) );
    aoi221_1 U2253 ( .x(n1193), .a(N5442), .b(___cell__36997_net130212), .c(
        branch_address[23]), .d(net148865), .e(n1286) );
    aoi22_1 U2254 ( .x(n1162), .a(branch_address[16]), .b(net148865), .c(N5435
        ), .d(___cell__36997_net130212) );
    aoi22_1 U2255 ( .x(n1158), .a(branch_address[0]), .b(net148865), .c(N5419), 
        .d(___cell__36997_net130212) );
    aoi22_1 U2256 ( .x(n1166), .a(branch_address[14]), .b(net148865), .c(N5433
        ), .d(___cell__36997_net130212) );
    aoi22_1 U2257 ( .x(n1170), .a(branch_address[8]), .b(net148865), .c(N5427), 
        .d(___cell__36997_net130212) );
    aoi22_1 U2258 ( .x(n1230), .a(branch_address[10]), .b(net148865), .c(N5429
        ), .d(___cell__36997_net130212) );
    aoi22_1 U2259 ( .x(n1206), .a(branch_address[9]), .b(net148865), .c(N5428), 
        .d(___cell__36997_net130709) );
    mux2i_1 U226 ( .x(n3900), .d0(n1673), .sl(n1650), .d1(n1374) );
    aoi22_1 U2260 ( .x(n1226), .a(branch_address[12]), .b(net148865), .c(N5431
        ), .d(___cell__36997_net130212) );
    aoi22_1 U2261 ( .x(n1202), .a(branch_address[4]), .b(net148865), .c(N5423), 
        .d(___cell__36997_net130212) );
    aoi22_1 U2262 ( .x(n1221), .a(branch_address[18]), .b(net148865), .c(N5437
        ), .d(___cell__36997_net130212) );
    aoi22_1 U2263 ( .x(n1185), .a(branch_address[25]), .b(net148865), .c(n1336
        ), .d(n797) );
    buf_16 U2265 ( .x(reg_out_A[7]), .a(n3971) );
    buf_16 U2266 ( .x(reg_out_A[3]), .a(n3974) );
    buf_16 U2267 ( .x(reg_out_A[16]), .a(n3965) );
    buf_16 U2268 ( .x(reg_out_A[8]), .a(n3970) );
    buf_16 U2269 ( .x(Imm[2]), .a(N6332) );
    inv_2 U227 ( .x(n1673), .a(N513) );
    buf_16 U2270 ( .x(Imm[4]), .a(N6336) );
    buf_16 U2271 ( .x(reg_out_A[17]), .a(n3964) );
    nand2_2 U2272 ( .x(n2641), .a(___cell__36997_net126604), .b(n1034) );
    nand2i_4 U2273 ( .x(n3807), .a(n1099), .b(n763) );
    nand2i_4 U2274 ( .x(n3813), .a(n1103), .b(n764) );
    nand2i_4 U2275 ( .x(n3822), .a(n1105), .b(n764) );
    nand2i_4 U2276 ( .x(n3820), .a(n1115), .b(n764) );
    nand2i_4 U2277 ( .x(n3821), .a(n1116), .b(n764) );
    nand2i_4 U2278 ( .x(n3818), .a(n1117), .b(n764) );
    nand2i_4 U2279 ( .x(n3816), .a(n1119), .b(n763) );
    inv_2 U228 ( .x(n1249), .a(n733) );
    nand2i_4 U2280 ( .x(n3819), .a(n1121), .b(n763) );
    nand2i_4 U2281 ( .x(n3808), .a(n1123), .b(n763) );
    nand2i_4 U2282 ( .x(n3817), .a(n1124), .b(n763) );
    nand2i_4 U2283 ( .x(n3814), .a(n1125), .b(n1100) );
    nand4_1 U2284 ( .x(n3851), .a(n1144), .b(n1147), .c(n1146), .d(n1145) );
    nand4_1 U2285 ( .x(n3844), .a(n1151), .b(n1149), .c(n1150), .d(n1148) );
    nand4_1 U2286 ( .x(n3825), .a(n1152), .b(n1153), .c(n1154), .d(n1155) );
    nand4_1 U2287 ( .x(n3824), .a(n1156), .b(n1157), .c(n1158), .d(n1159) );
    nand4_1 U2288 ( .x(n3840), .a(n1160), .b(n1161), .c(n1162), .d(n1163) );
    nand4_1 U2289 ( .x(n3838), .a(n1164), .b(n1165), .c(n1166), .d(n1167) );
    inv_2 U229 ( .x(n1501), .a(N6044) );
    nand4_1 U2290 ( .x(n3832), .a(n1168), .b(n1169), .c(n1170), .d(n1171) );
    nand4_1 U2291 ( .x(n3829), .a(n1172), .b(n1173), .c(n1174), .d(n1175) );
    nand4_1 U2293 ( .x(n3841), .a(n1180), .b(n1181), .c(n1182), .d(n1183) );
    nand4_1 U2294 ( .x(n3835), .a(n1188), .b(n1189), .c(n1190), .d(n1191) );
    nand4_1 U2296 ( .x(n3828), .a(n1200), .b(n1201), .c(n1202), .d(n1203) );
    nand4_1 U2297 ( .x(n3833), .a(n1204), .b(n1206), .c(n1207), .d(n1205) );
    nand4_1 U2298 ( .x(n3843), .a(n1208), .b(n1210), .c(n1209), .d(n1211) );
    nand4_1 U2299 ( .x(n3837), .a(n1212), .b(n1213), .c(n1214), .d(n1215) );
    oa21_2 U23 ( .x(n3923), .a(opcode_of_MEM_2), .b(n3924), .c(opcode_of_MEM_1
        ) );
    inv_2 U230 ( .x(n1502), .a(N5377) );
    nand4_1 U2300 ( .x(n3839), .a(n1218), .b(n1217), .c(n1216), .d(n1219) );
    nand4_1 U2301 ( .x(n3836), .a(n1224), .b(n1225), .c(n1226), .d(n1227) );
    nand4_1 U2302 ( .x(n3834), .a(n1228), .b(n1229), .c(n1230), .d(n1231) );
    nand4_1 U2304 ( .x(n3831), .a(n1246), .b(n1244), .c(n1245), .d(n1247) );
    nand4_1 U2305 ( .x(n3850), .a(n1248), .b(n1249), .c(n1250), .d(n1251) );
    nor2_5 U2306 ( .x(n1184), .a(___cell__36997_net129247), .b(n1281) );
    nor2_5 U2307 ( .x(n1254), .a(___cell__36997_net129247), .b(n1292) );
    nor2_5 U2308 ( .x(n1220), .a(n1272), .b(n1296) );
    nor2_5 U2309 ( .x(n1119), .a(n705), .b(n816) );
    mux2i_1 U231 ( .x(n3895), .d0(n1678), .sl(n1650), .d1(n1346) );
    nor2_5 U2310 ( .x(n1125), .a(n705), .b(n827) );
    nor2_5 U2311 ( .x(n1103), .a(n1776), .b(n789) );
    nor2_5 U2312 ( .x(n1118), .a(n705), .b(n649) );
    nor2_5 U2313 ( .x(n1123), .a(n705), .b(n803) );
    nor2_5 U2314 ( .x(n1099), .a(n1776), .b(n648) );
    mux2i_3 U2315 ( .x(n1258), .d0(n567), .sl(net149680), .d1(n1331) );
    mux2i_3 U2316 ( .x(n1344), .d0(n1345), .sl(___cell__36997_net129354), .d1(
        n1346) );
    mux2i_3 U2317 ( .x(n1350), .d0(n1351), .sl(___cell__36997_net129354), .d1(
        n1304) );
    mux2i_3 U2318 ( .x(n1352), .d0(n1353), .sl(___cell__36997_net129354), .d1(
        n1354) );
    mux2i_3 U2319 ( .x(___cell__36997_net129378), .d0(n1358), .sl(
        ___cell__36997_net129354), .d1(n1359) );
    inv_2 U232 ( .x(n1678), .a(N508) );
    mux2i_3 U2320 ( .x(___cell__36997_net129381), .d0(n1360), .sl(
        ___cell__36997_net129354), .d1(n1361) );
    mux2i_3 U2321 ( .x(n1364), .d0(n1365), .sl(___cell__36997_net129354), .d1(
        n1366) );
    mux2i_3 U2322 ( .x(n1369), .d0(n1370), .sl(___cell__36997_net129354), .d1(
        n1371) );
    mux2i_3 U2323 ( .x(n1372), .d0(n1373), .sl(___cell__36997_net129354), .d1(
        n1374) );
    mux2i_3 U2324 ( .x(n1388), .d0(n1389), .sl(___cell__36997_net129354), .d1(
        n1390) );
    mux2i_3 U2325 ( .x(n1393), .d0(n1394), .sl(___cell__36997_net129354), .d1(
        n1395) );
    mux2i_3 U2326 ( .x(n1398), .d0(n1399), .sl(___cell__36997_net129354), .d1(
        n1400) );
    mux2i_3 U2327 ( .x(n1401), .d0(n1402), .sl(___cell__36997_net129354), .d1(
        n1403) );
    mux2i_3 U2328 ( .x(n1404), .d0(n1405), .sl(___cell__36997_net129354), .d1(
        n1406) );
    mux2i_3 U2329 ( .x(n1407), .d0(n1408), .sl(___cell__36997_net129354), .d1(
        n1409) );
    mux2i_1 U233 ( .x(n3915), .d0(n1658), .sl(n1650), .d1(n1385) );
    mux2i_3 U2330 ( .x(IR_latched_14), .d0(n569), .sl(net149681), .d1(n1413)
         );
    mux2i_3 U2331 ( .x(IR_latched_13), .d0(n570), .sl(net149680), .d1(n1414)
         );
    mux2i_3 U2332 ( .x(IR_latched_11), .d0(n571), .sl(net149680), .d1(n1416)
         );
    mux2i_3 U2333 ( .x(n1051), .d0(current_IR_9), .sl(net149680), .d1(
        IR_latched_input[9]) );
    mux2i_3 U2334 ( .x(n1049), .d0(current_IR_8), .sl(n728), .d1(
        IR_latched_input[8]) );
    oai21_4 U2335 ( .x(n1451), .a(n1450), .b(n556), .c(n1452) );
    oai21_4 U2336 ( .x(n1476), .a(n1477), .b(n1478), .c(n1475) );
    nand2i_4 U2337 ( .x(n1108), .a(n1486), .b(n1430) );
    inv_6 U2338 ( .x(n1419), .a(IR_latched_input[4]) );
    inv_6 U2339 ( .x(n1273), .a(N5381) );
    inv_2 U234 ( .x(n1658), .a(N528) );
    inv_6 U2340 ( .x(n1505), .a(N6042) );
    inv_6 U2341 ( .x(n1296), .a(N5369) );
    exor2_3 U2342 ( .x(n1563), .a(reg_dst_of_MEM_0), .b(n879) );
    exor2_3 U2343 ( .x(n1457), .a(reg_dst_of_MEM_4), .b(n1132) );
    exor2_3 U2344 ( .x(n1569), .a(WB_index_2), .b(n1426) );
    exor2_3 U2345 ( .x(n1572), .a(WB_index_4), .b(n1132) );
    inv_6 U2346 ( .x(n1345), .a(N441) );
    inv_6 U2347 ( .x(n1348), .a(N451) );
    inv_6 U2348 ( .x(n1351), .a(N453) );
    inv_6 U2349 ( .x(n1353), .a(N457) );
    mux2i_1 U235 ( .x(n3751), .d0(n657), .sl(___cell__36997_net130681), .d1(
        n1329) );
    inv_6 U2350 ( .x(n1358), .a(N454) );
    inv_6 U2351 ( .x(n1360), .a(N442) );
    inv_6 U2354 ( .x(n1370), .a(N467) );
    inv_6 U2355 ( .x(n1373), .a(N446) );
    inv_6 U2356 ( .x(n1378), .a(N447) );
    inv_6 U2357 ( .x(n1384), .a(N461) );
    inv_6 U2358 ( .x(n1389), .a(N466) );
    inv_6 U2359 ( .x(n1394), .a(N460) );
    aoi222_1 U236 ( .x(n1023), .a(NPC[26]), .b(n1802), .c(n1732), .d(EPC_26), 
        .e(Cause_Reg_26), .f(n1803) );
    inv_6 U2360 ( .x(n1405), .a(N455) );
    inv_6 U2361 ( .x(n1408), .a(N444) );
    mux2i_3 U2362 ( .x(n3761), .d0(n656), .sl(___cell__36997_net126612), .d1(
        n3992) );
    mux2i_3 U2363 ( .x(n3421), .d0(n2630), .sl(n1857), .d1(n1800) );
    mux2i_3 U2364 ( .x(n3444), .d0(n2629), .sl(n1857), .d1(n1799) );
    mux2i_3 U2365 ( .x(n3453), .d0(n2606), .sl(n1856), .d1(n1603) );
    mux2i_3 U2366 ( .x(n3476), .d0(n2605), .sl(n1856), .d1(n1799) );
    mux2i_3 U2367 ( .x(n3485), .d0(n2582), .sl(n1855), .d1(n1800) );
    mux2i_3 U2368 ( .x(n3508), .d0(n2581), .sl(n1855), .d1(n1799) );
    mux2i_3 U2369 ( .x(n3517), .d0(n2558), .sl(n1854), .d1(n1603) );
    aoi22_2 U237 ( .x(n1148), .a(branch_address[20]), .b(n766), .c(N5439), .d(
        ___cell__36997_net130212) );
    mux2i_3 U2370 ( .x(n3540), .d0(n2557), .sl(n1854), .d1(n1799) );
    mux2i_3 U2371 ( .x(n3549), .d0(n2534), .sl(n1853), .d1(n1800) );
    mux2i_3 U2372 ( .x(n3572), .d0(n2533), .sl(n1853), .d1(n1799) );
    mux2i_3 U2373 ( .x(n3581), .d0(n2510), .sl(n1852), .d1(n1603) );
    mux2i_3 U2374 ( .x(n3604), .d0(n2509), .sl(n1852), .d1(n1799) );
    mux2i_3 U2375 ( .x(n3613), .d0(n2486), .sl(n1851), .d1(n1800) );
    mux2i_3 U2376 ( .x(n3636), .d0(n2485), .sl(n1851), .d1(n1799) );
    mux2i_3 U2377 ( .x(n2717), .d0(n2462), .sl(n1850), .d1(n1603) );
    mux2i_3 U2378 ( .x(n2740), .d0(n2461), .sl(n1850), .d1(n1799) );
    mux2i_3 U2379 ( .x(n2749), .d0(n2438), .sl(n1849), .d1(n1800) );
    mux2i_1 U238 ( .x(n3904), .d0(n1669), .sl(n1650), .d1(n1340) );
    mux2i_3 U2380 ( .x(n2772), .d0(n2437), .sl(n1849), .d1(n1799) );
    mux2i_3 U2381 ( .x(n3645), .d0(n2414), .sl(n1848), .d1(n1603) );
    mux2i_3 U2382 ( .x(n3668), .d0(n2413), .sl(n1848), .d1(n1799) );
    mux2i_3 U2383 ( .x(n2781), .d0(n2390), .sl(n1847), .d1(n1800) );
    mux2i_3 U2384 ( .x(n2804), .d0(n2389), .sl(n1847), .d1(n1799) );
    mux2i_3 U2385 ( .x(n2813), .d0(n2366), .sl(n1846), .d1(n1603) );
    mux2i_3 U2386 ( .x(n2836), .d0(n2365), .sl(n1846), .d1(n1799) );
    mux2i_3 U2387 ( .x(n2845), .d0(n2342), .sl(n1845), .d1(n1800) );
    mux2i_3 U2388 ( .x(n2868), .d0(n2341), .sl(n1845), .d1(n1799) );
    mux2i_3 U2389 ( .x(n2877), .d0(n2318), .sl(n1844), .d1(n1603) );
    inv_2 U239 ( .x(n1669), .a(N517) );
    mux2i_3 U2390 ( .x(n2900), .d0(n2317), .sl(n1844), .d1(n1799) );
    mux2i_3 U2391 ( .x(n2909), .d0(n2294), .sl(n1843), .d1(n1800) );
    mux2i_3 U2392 ( .x(n2932), .d0(n2293), .sl(n1843), .d1(n1799) );
    mux2i_3 U2393 ( .x(n2941), .d0(n2270), .sl(n1842), .d1(n1603) );
    mux2i_3 U2394 ( .x(n2964), .d0(n2269), .sl(n1842), .d1(n1799) );
    mux2i_3 U2395 ( .x(n2973), .d0(n2246), .sl(n1841), .d1(n1603) );
    mux2i_3 U2396 ( .x(n2996), .d0(n2245), .sl(n1841), .d1(n1799) );
    mux2i_3 U2397 ( .x(n3005), .d0(n2222), .sl(n1840), .d1(n1800) );
    mux2i_3 U2398 ( .x(n3028), .d0(n2221), .sl(n1840), .d1(n1799) );
    mux2i_3 U2399 ( .x(n3037), .d0(n2198), .sl(n1839), .d1(n1603) );
    nand2_2 U24 ( .x(n3946), .a(n3945), .b(n3924) );
    mux2i_1 U240 ( .x(n3909), .d0(n1664), .sl(n1650), .d1(n1406) );
    mux2i_3 U2400 ( .x(n3060), .d0(n2197), .sl(n1839), .d1(n1799) );
    mux2i_3 U2401 ( .x(n3069), .d0(n2174), .sl(n1838), .d1(n1800) );
    mux2i_3 U2402 ( .x(n3092), .d0(n2173), .sl(n1838), .d1(n1799) );
    mux2i_3 U2403 ( .x(n3677), .d0(n2150), .sl(n1837), .d1(n1800) );
    mux2i_3 U2404 ( .x(n3700), .d0(n2149), .sl(n1837), .d1(n1799) );
    mux2i_3 U2405 ( .x(n3101), .d0(n2126), .sl(n1836), .d1(n1603) );
    mux2i_3 U2406 ( .x(n3124), .d0(n2125), .sl(n1836), .d1(n1799) );
    mux2i_3 U2407 ( .x(n3133), .d0(n2102), .sl(n1835), .d1(n1800) );
    mux2i_3 U2408 ( .x(n3156), .d0(n2101), .sl(n1835), .d1(n1799) );
    mux2i_3 U2409 ( .x(n3165), .d0(n2078), .sl(n1834), .d1(n1603) );
    inv_2 U241 ( .x(n1664), .a(N522) );
    mux2i_3 U2410 ( .x(n3188), .d0(n2077), .sl(n1834), .d1(n1799) );
    mux2i_3 U2411 ( .x(n3197), .d0(n2054), .sl(n1833), .d1(n1800) );
    mux2i_3 U2412 ( .x(n3220), .d0(n2053), .sl(n1833), .d1(n1799) );
    mux2i_3 U2413 ( .x(n3229), .d0(n2030), .sl(n1832), .d1(n1603) );
    mux2i_3 U2414 ( .x(n3252), .d0(n2029), .sl(n1832), .d1(n1799) );
    mux2i_3 U2415 ( .x(n3261), .d0(n2006), .sl(n1831), .d1(n1800) );
    mux2i_3 U2416 ( .x(n3284), .d0(n2005), .sl(n1831), .d1(n1799) );
    mux2i_3 U2417 ( .x(n3293), .d0(n1982), .sl(n1830), .d1(n1603) );
    mux2i_3 U2418 ( .x(n3316), .d0(n1981), .sl(n1830), .d1(n1799) );
    mux2i_3 U2419 ( .x(n3325), .d0(n1958), .sl(n1829), .d1(n1603) );
    mux2i_3 U2420 ( .x(n3348), .d0(n1957), .sl(n1829), .d1(n1799) );
    mux2i_3 U2421 ( .x(n3357), .d0(n1934), .sl(n1828), .d1(n1800) );
    mux2i_3 U2422 ( .x(n3380), .d0(n1933), .sl(n1828), .d1(n1799) );
    mux2i_3 U2423 ( .x(n3389), .d0(n1910), .sl(n1827), .d1(n1800) );
    mux2i_3 U2424 ( .x(n3412), .d0(n1909), .sl(n1827), .d1(n1799) );
    mux2i_3 U2425 ( .x(n3710), .d0(n1887), .sl(n1826), .d1(n1801) );
    mux2i_3 U2426 ( .x(n3709), .d0(n1886), .sl(n1826), .d1(n1603) );
    mux2i_3 U2427 ( .x(n3732), .d0(n1885), .sl(n1826), .d1(n1799) );
    mux2i_3 U2428 ( .x(n3731), .d0(n1884), .sl(n1826), .d1(n1798) );
    mux2i_3 U2429 ( .x(n3730), .d0(n1883), .sl(n1826), .d1(n1797) );
    nand2i_2 U243 ( .x(n1046), .a(n643), .b(n1718) );
    mux2i_3 U2430 ( .x(n3729), .d0(n1882), .sl(n1826), .d1(n1796) );
    mux2i_3 U2431 ( .x(n3728), .d0(n1881), .sl(n1826), .d1(n1795) );
    mux2i_3 U2432 ( .x(n3727), .d0(n1880), .sl(n1826), .d1(n1794) );
    mux2i_3 U2433 ( .x(n3726), .d0(n1879), .sl(n1826), .d1(n1793) );
    mux2i_3 U2434 ( .x(n3725), .d0(n1878), .sl(n1826), .d1(n1792) );
    mux2i_3 U2435 ( .x(n3724), .d0(n1877), .sl(n1826), .d1(n1791) );
    mux2i_3 U2436 ( .x(n3723), .d0(n1876), .sl(n1826), .d1(n1790) );
    mux2i_3 U2437 ( .x(n3722), .d0(n1875), .sl(n1826), .d1(n1789) );
    mux2i_3 U2438 ( .x(n3721), .d0(n1874), .sl(n1826), .d1(n1788) );
    mux2i_3 U2439 ( .x(n3720), .d0(n1873), .sl(n1826), .d1(n1787) );
    mux2i_3 U2440 ( .x(n3719), .d0(n1872), .sl(n1826), .d1(n1786) );
    mux2i_3 U2441 ( .x(n3718), .d0(n1871), .sl(n1826), .d1(n1785) );
    mux2i_3 U2442 ( .x(n3717), .d0(n1870), .sl(n1826), .d1(n1784) );
    mux2i_3 U2443 ( .x(n3716), .d0(n1869), .sl(n1826), .d1(n1783) );
    mux2i_3 U2444 ( .x(n3715), .d0(n1868), .sl(n1826), .d1(n1782) );
    mux2i_3 U2445 ( .x(n3714), .d0(n1867), .sl(n1826), .d1(n1781) );
    mux2i_3 U2446 ( .x(n3713), .d0(n1866), .sl(n1826), .d1(n1780) );
    mux2i_3 U2447 ( .x(n3712), .d0(n1865), .sl(n1826), .d1(n1779) );
    mux2i_3 U2448 ( .x(n3711), .d0(n1864), .sl(n1826), .d1(n1778) );
    mux2i_3 U2449 ( .x(n2651), .d0(n618), .sl(___cell__36997_net130567), .d1(
        n873) );
    nand2i_2 U245 ( .x(n1048), .a(n734), .b(n642) );
    mux2i_3 U2450 ( .x(n2650), .d0(n619), .sl(___cell__36997_net130125), .d1(
        n872) );
    mux2i_3 U2451 ( .x(n2649), .d0(n620), .sl(___cell__36997_net130567), .d1(
        n734) );
    mux2i_3 U2452 ( .x(n2648), .d0(n621), .sl(___cell__36997_net130125), .d1(
        n643) );
    mux2i_3 U2453 ( .x(n2672), .d0(n597), .sl(___cell__36997_net130125), .d1(
        n701) );
    mux2i_3 U2454 ( .x(n2645), .d0(n624), .sl(___cell__36997_net130567), .d1(
        n886) );
    mux2i_3 U2455 ( .x(n2671), .d0(n598), .sl(___cell__36997_net130125), .d1(
        n762) );
    mux2i_3 U2456 ( .x(n2670), .d0(n599), .sl(___cell__36997_net130567), .d1(
        n696) );
    mux2i_3 U2457 ( .x(n2669), .d0(n600), .sl(___cell__36997_net130125), .d1(
        n765) );
    mux2i_3 U2458 ( .x(n2668), .d0(n601), .sl(___cell__36997_net130567), .d1(
        n735) );
    mux2i_3 U2459 ( .x(n2667), .d0(n602), .sl(___cell__36997_net130125), .d1(
        n816) );
    mux2i_3 U2460 ( .x(n2665), .d0(n604), .sl(___cell__36997_net130125), .d1(
        n827) );
    mux2i_3 U2461 ( .x(n2664), .d0(n605), .sl(___cell__36997_net130567), .d1(
        n789) );
    mux2i_3 U2462 ( .x(n2663), .d0(n606), .sl(___cell__36997_net130125), .d1(
        n649) );
    mux2i_3 U2463 ( .x(n2662), .d0(n607), .sl(___cell__36997_net130567), .d1(
        n732) );
    mux2i_3 U2464 ( .x(n2644), .d0(n625), .sl(___cell__36997_net130125), .d1(
        n870) );
    mux2i_3 U2465 ( .x(n2661), .d0(n608), .sl(___cell__36997_net130567), .d1(
        n775) );
    mux2i_3 U2466 ( .x(n2660), .d0(n609), .sl(___cell__36997_net130125), .d1(
        n778) );
    mux2i_3 U2467 ( .x(n2659), .d0(n610), .sl(___cell__36997_net130567), .d1(
        n803) );
    mux2i_3 U2468 ( .x(n2658), .d0(n611), .sl(___cell__36997_net130125), .d1(
        n648) );
    mux2i_3 U2469 ( .x(n2657), .d0(n612), .sl(___cell__36997_net130567), .d1(
        n829) );
    nand2i_4 U247 ( .x(n1058), .a(n779), .b(n642) );
    mux2i_3 U2470 ( .x(n2656), .d0(n613), .sl(___cell__36997_net130125), .d1(
        n647) );
    mux2i_3 U2471 ( .x(n2654), .d0(n615), .sl(___cell__36997_net130125), .d1(
        n779) );
    mux2i_3 U2472 ( .x(n2653), .d0(n616), .sl(___cell__36997_net130567), .d1(
        n786) );
    mux2i_3 U2473 ( .x(n2643), .d0(n626), .sl(___cell__36997_net130567), .d1(
        n720) );
    nand4_1 U2474 ( .x(n1486), .a(n739), .b(n1081), .c(n1067), .d(n767) );
    and4i_5 U2475 ( .x(n1447), .a(n1558), .b(n1697), .c(n1696), .d(n1695) );
    and3i_4 U2477 ( .x(___cell__36997_net130187), .a(n1685), .b(reg_write_WB), 
        .c(n1569) );
    nor2_5 U2478 ( .x(n1705), .a(___cell__36997_net130191), .b(n1704) );
    nor2_5 U2479 ( .x(n1708), .a(n1706), .b(n1707) );
    mux2i_1 U248 ( .x(n3903), .d0(n1670), .sl(n1650), .d1(n1383) );
    nor2_5 U2480 ( .x(n1711), .a(n1709), .b(n1710) );
    inv_6 U2481 ( .x(n1654), .a(N531) );
    inv_5 U2482 ( .x(n1857), .a(n1741) );
    inv_5 U2483 ( .x(n1856), .a(n1742) );
    inv_5 U2484 ( .x(n1855), .a(n1743) );
    inv_5 U2485 ( .x(n1854), .a(n1744) );
    inv_5 U2486 ( .x(n1853), .a(n1745) );
    inv_5 U2487 ( .x(n1852), .a(n1746) );
    inv_5 U2488 ( .x(n1851), .a(n1747) );
    inv_5 U2489 ( .x(n1850), .a(n1748) );
    inv_2 U249 ( .x(n1670), .a(N516) );
    inv_5 U2490 ( .x(n1849), .a(n1749) );
    inv_5 U2491 ( .x(n1848), .a(n1750) );
    inv_5 U2492 ( .x(n1847), .a(n1751) );
    inv_5 U2493 ( .x(n1846), .a(n1752) );
    inv_5 U2494 ( .x(n1845), .a(n1753) );
    inv_5 U2495 ( .x(n1844), .a(n1754) );
    inv_5 U2496 ( .x(n1843), .a(n1755) );
    inv_5 U2497 ( .x(n1842), .a(n1756) );
    inv_5 U2498 ( .x(n1841), .a(n1757) );
    inv_5 U2499 ( .x(n1840), .a(n1758) );
    nand2_2 U25 ( .x(n3947), .a(n556), .b(n3932) );
    mux2i_1 U250 ( .x(n3908), .d0(n1665), .sl(n1650), .d1(n1359) );
    inv_5 U2500 ( .x(n1839), .a(n1759) );
    inv_5 U2501 ( .x(n1838), .a(n1760) );
    inv_5 U2502 ( .x(n1837), .a(n1761) );
    inv_5 U2503 ( .x(n1836), .a(n1762) );
    inv_5 U2504 ( .x(n1835), .a(n1763) );
    inv_5 U2505 ( .x(n1834), .a(n1764) );
    inv_5 U2506 ( .x(n1833), .a(n1765) );
    inv_5 U2507 ( .x(n1832), .a(n1766) );
    inv_5 U2508 ( .x(n1831), .a(n1767) );
    inv_5 U2509 ( .x(n1830), .a(n1768) );
    inv_2 U251 ( .x(n1665), .a(N521) );
    inv_5 U2510 ( .x(n1829), .a(n1769) );
    inv_5 U2511 ( .x(n1828), .a(n1770) );
    inv_5 U2512 ( .x(n1827), .a(n1771) );
    inv_5 U2513 ( .x(n1826), .a(n1772) );
    buf_16 U2514 ( .x(n331), .a(n761) );
    buf_16 U2515 ( .x(n336), .a(n1258) );
    buf_16 U2516 ( .x(Imm[0]), .a(N6328) );
    buf_16 U2517 ( .x(Imm[5]), .a(N6338) );
    buf_16 U2518 ( .x(Imm[29]), .a(N6386) );
    buf_16 U2519 ( .x(Imm[30]), .a(N6388) );
    mux2i_1 U252 ( .x(n3917), .d0(n1655), .sl(n1650), .d1(n1368) );
    buf_16 U2520 ( .x(reg_out_B[4]), .a(n3980) );
    buf_16 U2521 ( .x(reg_out_B[1]), .a(n3983) );
    buf_16 U2522 ( .x(reg_out_A[4]), .a(n3973) );
    buf_16 U2523 ( .x(reg_out_A[19]), .a(n3962) );
    buf_16 U2524 ( .x(reg_out_A[18]), .a(n3963) );
    buf_16 U2525 ( .x(reg_out_B[3]), .a(n3981) );
    buf_16 U2526 ( .x(reg_out_A[21]), .a(n3960) );
    buf_16 U2527 ( .x(reg_out_A[30]), .a(n3951) );
    nand2i_5 U2528 ( .x(___cell__36997_net126604), .a(___cell__36997_net127190
        ), .b(n1484) );
    nand2i_6 U2529 ( .x(n1776), .a(___cell__36997_net130681), .b(n1461) );
    inv_2 U253 ( .x(n1655), .a(N530) );
    nand2i_5 U2531 ( .x(n1145), .a(n1499), .b(___cell__36997_net130212) );
    aoai211_5 U2532 ( .x(n1134), .a(n1570), .b(n1494), .c(n1712), .d(
        ___cell__36997_net126612) );
    nand2i_8 U2533 ( .x(___cell__36997_net127190), .a(n1259), .b(n1461) );
    inv_16 U2534 ( .x(___cell__36997_net126612), .a(___cell__36997_net127190)
         );
    inv_16 U2535 ( .x(n1132), .a(n336) );
    nand2i_6 U2536 ( .x(___cell__36997_net129626), .a(n1491), .b(n1437) );
    inv_14 U2537 ( .x(n1484), .a(n1471) );
    nand2i_6 U2538 ( .x(n1263), .a(n1470), .b(n860) );
    nand4i_5 U2539 ( .x(n1480), .a(n1264), .b(n1481), .c(n1482), .d(n1483) );
    nand2i_2 U254 ( .x(n1062), .a(n647), .b(n642) );
    inv_14 U2540 ( .x(n1802), .a(n1307) );
    nor2i_8 U2541 ( .x(n1554), .a(n1461), .b(n642) );
    inv_16 U2542 ( .x(n1732), .a(n1518) );
    nand2_8 U2543 ( .x(n1647), .a(n1514), .b(n1648) );
    nand2_8 U2544 ( .x(n1645), .a(n1514), .b(n1646) );
    nand2_8 U2545 ( .x(n1643), .a(n1514), .b(n1644) );
    nand2_8 U2546 ( .x(n1641), .a(n1514), .b(n1642) );
    nand2_8 U2547 ( .x(n1639), .a(n1514), .b(n1640) );
    nand2_8 U2548 ( .x(n1637), .a(n1514), .b(n1638) );
    nand2_8 U2549 ( .x(n1635), .a(n1605), .b(n1636) );
    ao21_1 U255 ( .x(n1473), .a(n1714), .b(___cell__36997_net127190), .c(n1093
        ) );
    nand2_8 U2550 ( .x(n1633), .a(n1605), .b(n1634) );
    nand2_8 U2551 ( .x(n1631), .a(n1605), .b(n1632) );
    nand2_8 U2552 ( .x(n1629), .a(n1605), .b(n1630) );
    nand2_8 U2553 ( .x(n1627), .a(n1605), .b(n1628) );
    nand2_8 U2554 ( .x(n1625), .a(n1605), .b(n1626) );
    nand2_8 U2555 ( .x(n1623), .a(n1605), .b(n1624) );
    nand2_8 U2556 ( .x(n1621), .a(n1605), .b(n1622) );
    nand2_8 U2557 ( .x(n1619), .a(n1605), .b(n1620) );
    nand2_8 U2558 ( .x(n1617), .a(n1605), .b(n1618) );
    nand2_8 U2559 ( .x(n1615), .a(n1605), .b(n1616) );
    inv_5 U256 ( .x(n1494), .a(n1465) );
    nand2_8 U2560 ( .x(n1613), .a(n1605), .b(n1614) );
    nand2_8 U2561 ( .x(n1611), .a(n1605), .b(n1612) );
    nand2_8 U2562 ( .x(n1609), .a(n1605), .b(n1610) );
    nand2_8 U2563 ( .x(n1607), .a(n1605), .b(n1608) );
    nand2_8 U2564 ( .x(n1601), .a(n1514), .b(n1602) );
    inv_16 U2565 ( .x(___cell__36997_net130217), .a(net148858) );
    inv_10 U2566 ( .x(n1492), .a(n1263) );
    nand3_4 U2567 ( .x(n1260), .a(n1460), .b(n564), .c(net152025) );
    nand2_8 U2568 ( .x(n1471), .a(n650), .b(n1436) );
    nand2i_8 U2569 ( .x(n1514), .a(n1723), .b(n1740) );
    mux2i_1 U257 ( .x(n3739), .d0(n1594), .sl(___cell__36997_net130681), .d1(
        n1595) );
    inv_16 U2570 ( .x(n1605), .a(n1513) );
    nand3i_5 U2571 ( .x(___cell__36997_net129625), .a(n1721), .b(n1465), .c(
        n834) );
    nand2i_6 U2572 ( .x(n1465), .a(n836), .b(n682) );
    nand2i_8 U2573 ( .x(n1511), .a(N13832), .b(n1512) );
    nand2i_8 U2574 ( .x(n1513), .a(n1302), .b(n1514) );
    nand4_5 U2575 ( .x(n1303), .a(opcode_of_WB_5), .b(n3889), .c(n3887), .d(
        n3890) );
    exnor2_5 U2577 ( .x(n1558), .a(n1559), .b(n331) );
    exor2_5 U2578 ( .x(n1683), .a(n635), .b(___cell__36997_net129477) );
    mux2i_1 U258 ( .x(n3899), .d0(n1674), .sl(n1650), .d1(n1403) );
    inv_2 U259 ( .x(n1674), .a(N512) );
    exnor2_1 U26 ( .x(n667), .a(reg_dst_of_MEM_1), .b(n1071) );
    mux2i_1 U260 ( .x(n3898), .d0(n1675), .sl(n1650), .d1(n1409) );
    inv_2 U261 ( .x(n1675), .a(N511) );
    inv_2 U2611 ( .x(n1858), .a(reset) );
    inv_2 U2612 ( .x(n848), .a(n1088) );
    inv_7 U2613 ( .x(n749), .a(n3997) );
    inv_7 U2614 ( .x(n1197), .a(n4005) );
    mux2i_1 U2615 ( .x(n815), .d0(n1318), .sl(net149681), .d1(n1319) );
    inv_10 U2616 ( .x(n1081), .a(n712) );
    inv_6 U2617 ( .x(n716), .a(n1317) );
    mux2i_3 U2618 ( .x(n887), .d0(n568), .sl(net149680), .d1(n1412) );
    mux2i_3 U2619 ( .x(n831), .d0(n1418), .sl(net149680), .d1(n1419) );
    mux2i_1 U262 ( .x(n3921), .d0(n1651), .sl(n1650), .d1(n1371) );
    mux2i_6 U2620 ( .x(IR_latched_2), .d0(n1422), .sl(net149236), .d1(n1421)
         );
    nand4_3 U2621 ( .x(n1709), .a(n1018), .b(n1001), .c(n636), .d(n1031) );
    inv_4 U2622 ( .x(n1367), .a(N463) );
    oa22_3 U2623 ( .x(n823), .a(n724), .b(n711), .c(n1688), .d(n1431) );
    nand4_4 U2624 ( .x(n1707), .a(n638), .b(n1252), .c(n673), .d(n672) );
    nand2_8 U2625 ( .x(___cell__36997_net129624), .a(n1713), .b(n1481) );
    nand2i_5 U2626 ( .x(n1481), .a(n1715), .b(n682) );
    mux2i_3 U2627 ( .x(n3984), .d0(n1376), .sl(n798), .d1(n1375) );
    inv_6 U2628 ( .x(n663), .a(n3984) );
    inv_5 U2629 ( .x(n1375), .a(N452) );
    inv_2 U263 ( .x(n1651), .a(N534) );
    buf_14 U2630 ( .x(net148858), .a(___cell__36997_net127155) );
    inv_6 U2631 ( .x(n799), .a(___cell__36997_net127155) );
    nand4_4 U2632 ( .x(___cell__36997_net130191), .a(n641), .b(
        ___cell__36997_net126005), .c(___cell__36997_net125989), .d(
        ___cell__36997_net125941) );
    nand2i_2 U2633 ( .x(n794), .a(n641), .b(n797) );
    inv_0 U2634 ( .x(n3985), .a(n1364) );
    inv_5 U2635 ( .x(n994), .a(n1364) );
    inv_5 U2636 ( .x(n1365), .a(N468) );
    inv_1 U2637 ( .x(n3986), .a(n848) );
    inv_10 U2638 ( .x(n1088), .a(n889) );
    buf_16 U2639 ( .x(reg_out_B[22]), .a(n3977) );
    nand2_2 U264 ( .x(n1114), .a(n642), .b(IR_opcode_field[2]) );
    nand4_1 U2640 ( .x(n3830), .a(n1176), .b(n1177), .c(n1178), .d(n1179) );
    aoi21_4 U2641 ( .x(n1176), .a(N5357), .b(n862), .c(n1269) );
    buf_2 U2642 ( .x(n833), .a(n339) );
    nand3_4 U2643 ( .x(n782), .a(n855), .b(n700), .c(n747) );
    nor3i_2 U2644 ( .x(n1699), .a(n1440), .b(n837), .c(n825) );
    inv_5 U2645 ( .x(n1269), .a(n4007) );
    mux2i_8 U2646 ( .x(n884), .d0(n644), .sl(n736), .d1(IR_latched_input[16])
         );
    inv_10 U2647 ( .x(n736), .a(net149236) );
    exnor2_3 U2648 ( .x(n3987), .a(n3988), .b(n879) );
    inv_4 U2649 ( .x(n748), .a(n3987) );
    aoi222_1 U265 ( .x(n1025), .a(NPC[27]), .b(n1719), .c(n1732), .d(EPC_27), 
        .e(Cause_Reg_27), .f(n1803) );
    inv_4 U2650 ( .x(n3988), .a(reg_dst_of_EX_0) );
    mux2i_8 U2651 ( .x(n879), .d0(IR_latched_input[21]), .sl(net149236), .d1(
        current_IR_21) );
    nor2_2 U2652 ( .x(n1464), .a(n1688), .b(n1113) );
    inv_7 U2653 ( .x(n1113), .a(n1315) );
    aoi22_2 U2654 ( .x(n1246), .a(N5426), .b(___cell__36997_net130212), .c(
        N6025), .d(___cell__36997_net130713) );
    aoi211_1 U2655 ( .x(n3989), .a(n1083), .b(n853), .c(n1081), .d(n1113) );
    inv_7 U2656 ( .x(n853), .a(n850) );
    inv_10 U2657 ( .x(n3990), .a(n768) );
    inv_6 U2658 ( .x(n334), .a(n768) );
    buf_10 U2659 ( .x(net149680), .a(___cell__36997_net130572) );
    mux2i_1 U266 ( .x(n3912), .d0(n1661), .sl(n1650), .d1(n1392) );
    buf_14 U2660 ( .x(net149681), .a(n731) );
    buf_4 U2661 ( .x(n837), .a(n1313) );
    nand4_3 U2662 ( .x(n3854), .a(n1135), .b(n758), .c(n1136), .d(n1137) );
    inv_7 U2663 ( .x(n1135), .a(n3996) );
    inv_0 U2664 ( .x(n3991), .a(n1111) );
    inv_2 U2665 ( .x(n3992), .a(n3991) );
    mux2i_6 U2666 ( .x(n1111), .d0(IR_latched_input[29]), .sl(net149236), .d1(
        current_IR_29) );
    and2_4 U2667 ( .x(n4432), .a(n3910), .b(n681) );
    aoi21_3 U2668 ( .x(n1244), .a(N5358), .b(n863), .c(n1598) );
    inv_6 U2669 ( .x(___cell__36997_net126005), .a(___cell__36997_net129384)
         );
    inv_2 U267 ( .x(n1661), .a(N525) );
    mux2i_5 U2670 ( .x(___cell__36997_net129384), .d0(n1362), .sl(
        ___cell__36997_net129354), .d1(n1363) );
    and4i_3 U2671 ( .x(n1453), .a(n1683), .b(n1698), .c(n1562), .d(n1564) );
    exor2_3 U2672 ( .x(n1564), .a(reg_dst_of_MEM_1), .b(n1565) );
    nand2i_4 U2673 ( .x(n1313), .a(n709), .b(n1453) );
    nand4_3 U2674 ( .x(n3846), .a(n749), .b(n1235), .c(n676), .d(n1236) );
    nand4_3 U2675 ( .x(n3848), .a(n1197), .b(n1196), .c(n1198), .d(n1199) );
    ao22_3 U2676 ( .x(n3993), .a(branch_address[19]), .b(n766), .c(N5438), .d(
        ___cell__36997_net130709) );
    inv_4 U2677 ( .x(n1210), .a(n3993) );
    inv_16 U2678 ( .x(___cell__36997_net130709), .a(___cell__36997_net129247)
         );
    aoi22_3 U2679 ( .x(n1208), .a(N5370), .b(n895), .c(N6037), .d(
        ___cell__36997_net130214) );
    inv_12 U268 ( .x(n724), .a(n739) );
    ao211_5 U2680 ( .x(_branch_address_reg_31_net46811), .a(N5450), .b(n783), 
        .c(n664), .d(n792) );
    aoi21_2 U2681 ( .x(n1164), .a(N5365), .b(n862), .c(n1299) );
    nor2i_1 U2682 ( .x(n1299), .a(N6032), .b(___cell__36997_net129239) );
    buf_8 U2683 ( .x(reg_out_B[6]), .a(n4457) );
    aoi21_3 U2684 ( .x(n1139), .a(N5380), .b(n862), .c(n1278) );
    oai21_5 U2685 ( .x(n3995), .a(n1484), .b(n1480), .c(n1554) );
    ao221_5 U2686 ( .x(n3996), .a(___cell__36997_net129384), .b(n797), .c(
        branch_address[30]), .d(n766), .e(n1271) );
    nor2_6 U2687 ( .x(n1271), .a(n1272), .b(n1273) );
    nor2_4 U2688 ( .x(n1286), .a(net148915), .b(n1287) );
    nor2_3 U2689 ( .x(n1295), .a(net148915), .b(n585) );
    inv_2 U269 ( .x(n1504), .a(N5375) );
    inv_5 U2690 ( .x(n1270), .a(n835) );
    ao221_5 U2691 ( .x(n3997), .a(N5441), .b(___cell__36997_net130709), .c(
        branch_address[22]), .d(n766), .e(n1288) );
    nor2_4 U2692 ( .x(n1288), .a(net148913), .b(n1289) );
    inv_16 U2693 ( .x(___cell__36997_net130212), .a(___cell__36997_net129247)
         );
    inv_3 U2694 ( .x(n1277), .a(N5448) );
    nand4i_2 U2695 ( .x(n3849), .a(n1184), .b(n1186), .c(n1185), .d(n1187) );
    nor2_6 U2696 ( .x(n1290), .a(net148916), .b(n1291) );
    nand4i_1 U2697 ( .x(n792), .a(___cell__36997_net129654), .b(
        ___cell__36997_net129657), .c(n794), .d(n793) );
    buf_2 U2698 ( .x(n3998), .a(n805) );
    buf_14 U2699 ( .x(Imm[14]), .a(N6356) );
    buf_14 U27 ( .x(reg_out_A[12]), .a(n3966) );
    inv_2 U270 ( .x(n1510), .a(N6033) );
    buf_14 U2700 ( .x(Imm[6]), .a(N6340) );
    oai22_2 U2701 ( .x(n3795), .a(n705), .b(n871), .c(n3995), .d(n1043) );
    aoi21_2 U2702 ( .x(n1186), .a(N6043), .b(___cell__36997_net130713), .c(
        n1282) );
    oa22_4 U2703 ( .x(n1204), .a(n4004), .b(n1272), .c(n4003), .d(
        ___cell__36997_net129239) );
    mux2i_8 U2704 ( .x(n3999), .d0(n4001), .sl(n4000), .d1(n4002) );
    inv_0 U2705 ( .x(n1045), .a(n3999) );
    inv_10 U2706 ( .x(n4000), .a(n728) );
    inv_2 U2707 ( .x(n4001), .a(IR_latched_input[6]) );
    inv_2 U2708 ( .x(n4002), .a(current_IR_6) );
    buf_14 U2709 ( .x(n728), .a(n731) );
    nand2i_2 U271 ( .x(n1079), .a(n1861), .b(n642) );
    inv_16 U2710 ( .x(n895), .a(n1272) );
    inv_0 U2711 ( .x(n4003), .a(N6027) );
    inv_0 U2712 ( .x(n4004), .a(N5360) );
    nand2_5 U2713 ( .x(___cell__36997_net129239), .a(net148863), .b(n1494) );
    buf_16 U2714 ( .x(Imm[13]), .a(N6354) );
    buf_8 U2715 ( .x(reg_out_B[2]), .a(n3982) );
    mux2i_8 U2716 ( .x(n817), .d0(n1595), .sl(net152024), .d1(n1594) );
    and2_4 U2717 ( .x(n4442), .a(n3905), .b(n680) );
    inv_8 U2718 ( .x(net148865), .a(n738) );
    ao221_5 U2719 ( .x(n4005), .a(N5443), .b(___cell__36997_net130709), .c(
        branch_address[24]), .d(n766), .e(n1284) );
    nor2_3 U272 ( .x(n1124), .a(n1776), .b(n735) );
    buf_8 U2720 ( .x(n766), .a(n1804) );
    aoi22_2 U2721 ( .x(n1142), .a(branch_address[28]), .b(net148865), .c(N6046
        ), .d(___cell__36997_net130214) );
    nor2i_5 U2722 ( .x(n1698), .a(n1563), .b(n1684) );
    buf_10 U2723 ( .x(Imm[16]), .a(N6360) );
    buf_14 U2724 ( .x(Imm[18]), .a(N6364) );
    buf_10 U2725 ( .x(IR_opcode_field[1]), .a(n4453) );
    inv_8 U2726 ( .x(n1130), .a(n1369) );
    nand2i_4 U2727 ( .x(n4007), .a(n4008), .b(___cell__36997_net130214) );
    inv_0 U2728 ( .x(n4008), .a(N6024) );
    exnor2_2 U2729 ( .x(n770), .a(reg_dst_of_EX_1), .b(n339) );
    mux2i_1 U273 ( .x(n3906), .d0(n1667), .sl(n1650), .d1(n1376) );
    nor3i_0 U2730 ( .x(n1729), .a(FREEZE), .b(reg_dst_of_EX_2), .c(
        reg_dst_of_EX_1) );
    inv_5 U2731 ( .x(n1557), .a(reg_dst_of_EX_1) );
    mux2i_5 U2732 ( .x(reg_dst_of_EX_1), .d0(n560), .sl(reg_dst), .d1(n563) );
    inv_6 U2733 ( .x(n4009), .a(n4452) );
    inv_10 U2734 ( .x(IR_opcode_field[2]), .a(n4009) );
    inv_3 U2735 ( .x(n4011), .a(n3950) );
    mux2_4 U2736 ( .x(n1128), .d0(n1657), .sl(n798), .d1(n4012) );
    inv_4 U2737 ( .x(n4012), .a(N462) );
    nand2i_6 U2738 ( .x(n798), .a(n709), .b(n796) );
    inv_10 U2739 ( .x(IR_opcode_field[0]), .a(n4377) );
    inv_2 U274 ( .x(n1667), .a(N519) );
    buf_16 U2740 ( .x(Imm[10]), .a(N6348) );
    buf_14 U2741 ( .x(reg_out_B[25]), .a(n4455) );
    buf_10 U2742 ( .x(Imm[12]), .a(N6352) );
    buf_10 U2743 ( .x(Imm[31]), .a(N6390) );
    buf_14 U2744 ( .x(Imm[8]), .a(N6344) );
    buf_10 U2745 ( .x(reg_out_B[19]), .a(n4456) );
    and2_4 U2746 ( .x(n4390), .a(n3902), .b(n680) );
    buf_10 U2747 ( .x(reg_out_B[0]), .a(n4458) );
    and2_4 U2748 ( .x(n4394), .a(n3911), .b(n680) );
    and2_4 U2749 ( .x(n4410), .a(n3906), .b(n680) );
    mux2i_1 U275 ( .x(n3905), .d0(n1668), .sl(n1650), .d1(n1349) );
    and2_4 U2750 ( .x(n4434), .a(n3897), .b(n680) );
    and2_4 U2751 ( .x(n4422), .a(n3903), .b(n680) );
    and2_4 U2752 ( .x(n4430), .a(n3895), .b(n680) );
    and2_1 U2753 ( .x(n4388), .a(n3913), .b(n680) );
    and2_1 U2754 ( .x(n4392), .a(n3922), .b(n680) );
    and2_1 U2755 ( .x(n4396), .a(n3893), .b(n681) );
    and2_1 U2756 ( .x(n4398), .a(n3918), .b(n681) );
    and2_1 U2757 ( .x(n4400), .a(n3894), .b(n680) );
    and2_1 U2758 ( .x(n4402), .a(n3907), .b(n680) );
    and2_1 U2759 ( .x(n4404), .a(n3916), .b(n680) );
    inv_2 U276 ( .x(n1668), .a(N518) );
    and2_1 U2760 ( .x(n4406), .a(n3896), .b(n680) );
    and2_1 U2761 ( .x(n4408), .a(n3914), .b(n680) );
    and2_1 U2762 ( .x(n4412), .a(n3912), .b(n680) );
    and2_1 U2763 ( .x(n4414), .a(n3899), .b(n680) );
    and2_1 U2764 ( .x(n4416), .a(n3898), .b(n680) );
    and2_1 U2765 ( .x(n4418), .a(n3917), .b(n680) );
    and2_1 U2766 ( .x(n4420), .a(n3908), .b(n680) );
    and2_1 U2767 ( .x(n4424), .a(n3909), .b(n680) );
    and2_1 U2768 ( .x(n4426), .a(n3904), .b(n680) );
    and2_1 U2769 ( .x(n4428), .a(n3915), .b(n680) );
    mux2i_1 U277 ( .x(n3914), .d0(n1659), .sl(n1650), .d1(n1395) );
    and2_1 U2770 ( .x(n4436), .a(n3901), .b(n681) );
    and2_1 U2771 ( .x(n4438), .a(n3920), .b(n681) );
    and2_1 U2772 ( .x(n4440), .a(n3919), .b(n681) );
    and2_1 U2773 ( .x(n4444), .a(n3921), .b(n681) );
    and2_1 U2774 ( .x(n4446), .a(n3900), .b(n681) );
    and2_1 U2775 ( .x(n4448), .a(n3892), .b(n681) );
    and2_1 U2776 ( .x(n4450), .a(n3891), .b(n680) );
    inv_2 U278 ( .x(n1659), .a(N527) );
    nor2_2 U279 ( .x(n1239), .a(___cell__36997_net129247), .b(n1274) );
    buf_14 U28 ( .x(reg_out_A[20]), .a(n3961) );
    inv_2 U280 ( .x(n1274), .a(N5422) );
    inv_2 U281 ( .x(n1292), .a(N5421) );
    inv_2 U282 ( .x(n1281), .a(N5444) );
    inv_2 U283 ( .x(n1503), .a(N5376) );
    inv_2 U284 ( .x(n1509), .a(N5372) );
    aoi222_1 U285 ( .x(n1022), .a(NPC[25]), .b(n1719), .c(n1732), .d(EPC_25), 
        .e(Cause_Reg_25), .f(n1803) );
    inv_2 U286 ( .x(n1507), .a(N6041) );
    inv_2 U287 ( .x(n1506), .a(N5374) );
    oai21_1 U288 ( .x(N6749), .a(n641), .b(___cell__36997_net130580), .c(
        ___cell__36997_net127210) );
    mux2_4 U289 ( .x(n641), .d0(___cell__36997_net129388), .sl(
        ___cell__36997_net129354), .d1(___cell__36997_net129389) );
    inv_0 U29 ( .x(n1528), .a(NPC[26]) );
    and2_1 U290 ( .x(n677), .a(n3948), .b(n1515) );
    aoi222_1 U291 ( .x(___cell__36997_net127210), .a(NPC[31]), .b(n1719), .c(
        n1732), .d(EPC_31), .e(Cause_Reg_31), .f(n1803) );
    nor2_1 U292 ( .x(n1120), .a(n1776), .b(n778) );
    inv_5 U293 ( .x(IR_latched_10), .a(n1053) );
    nand2i_2 U294 ( .x(n1054), .a(n4371), .b(n642) );
    nand2i_2 U295 ( .x(n1060), .a(n4370), .b(n1718) );
    nor2_1 U296 ( .x(n1102), .a(n1776), .b(n732) );
    nand2i_2 U297 ( .x(n3811), .a(n1102), .b(n764) );
    nand2i_2 U298 ( .x(n1056), .a(n786), .b(n1718) );
    buf_3 U299 ( .x(n910), .a(n951) );
    and2_5 U3 ( .x(n664), .a(___cell__36997_net130214), .b(N6049) );
    inv_2 U30 ( .x(n750), .a(n3979) );
    mux2i_1 U300 ( .x(n3896), .d0(n1677), .sl(n1650), .d1(n1361) );
    inv_2 U301 ( .x(n1677), .a(N509) );
    nor2_1 U302 ( .x(n1101), .a(n705), .b(n775) );
    nand2i_2 U303 ( .x(n1050), .a(n872), .b(n1718) );
    oai21_1 U306 ( .x(N6742), .a(n1020), .b(n678), .c(n1021) );
    inv_5 U307 ( .x(n1020), .a(n1407) );
    aoi222_1 U308 ( .x(n1021), .a(NPC[24]), .b(n1802), .c(n1732), .d(EPC_24), 
        .e(Cause_Reg_24), .f(n1803) );
    oai21_1 U309 ( .x(N6746), .a(n1026), .b(n995), .c(n1027) );
    inv_7 U310 ( .x(n1026), .a(n1355) );
    aoi222_1 U311 ( .x(n1027), .a(NPC[28]), .b(n1802), .c(n1732), .d(EPC_28), 
        .e(Cause_Reg_28), .f(n1803) );
    mux2i_1 U312 ( .x(n3916), .d0(n1656), .sl(n1650), .d1(n1657) );
    inv_2 U313 ( .x(n1656), .a(N529) );
    mux2i_1 U314 ( .x(n3907), .d0(n1666), .sl(n1650), .d1(n1304) );
    inv_2 U315 ( .x(n1666), .a(N520) );
    oai21_1 U316 ( .x(N6748), .a(___cell__36997_net126005), .b(n995), .c(n1030
        ) );
    inv_4 U318 ( .x(n1362), .a(N438) );
    aoi222_1 U319 ( .x(n1030), .a(NPC[30]), .b(n1802), .c(n1732), .d(EPC_30), 
        .e(Cause_Reg_30), .f(n1803) );
    inv_2 U32 ( .x(n1061), .a(IR_latched_14) );
    buf_3 U320 ( .x(n909), .a(n951) );
    mux2i_1 U321 ( .x(n3894), .d0(n1679), .sl(n1650), .d1(n1357) );
    inv_2 U322 ( .x(n1679), .a(N507) );
    oai21_1 U323 ( .x(N6739), .a(n684), .b(___cell__36997_net130580), .c(n1015
        ) );
    aoi222_1 U324 ( .x(n1015), .a(NPC[21]), .b(n1719), .c(n1732), .d(EPC_21), 
        .e(Cause_Reg_21), .f(n1803) );
    inv_2 U325 ( .x(___cell__36997_net130580), .a(n677) );
    aoi222_1 U326 ( .x(n1029), .a(NPC[29]), .b(n1719), .c(n1732), .d(EPC_29), 
        .e(Cause_Reg_29), .f(n1803) );
    inv_2 U327 ( .x(n678), .a(n677) );
    inv_4 U328 ( .x(n1342), .a(N439) );
    inv_7 U329 ( .x(n1028), .a(n1341) );
    inv_0 U33 ( .x(n1597), .a(IR_latched_input[10]) );
    oai21_1 U330 ( .x(N6747), .a(n1028), .b(n678), .c(n1029) );
    aoi222_1 U331 ( .x(n1017), .a(NPC[22]), .b(n1802), .c(n1732), .d(EPC_22), 
        .e(Cause_Reg_22), .f(n1803) );
    nand2_2 U332 ( .x(n995), .a(n3948), .b(n1515) );
    oai21_1 U333 ( .x(N6740), .a(n1016), .b(n995), .c(n1017) );
    oai21_1 U334 ( .x(N6741), .a(n1018), .b(n1777), .c(n1019) );
    inv_5 U335 ( .x(n1018), .a(n1401) );
    aoi222_1 U336 ( .x(n1019), .a(NPC[23]), .b(n1719), .c(n1732), .d(EPC_23), 
        .e(Cause_Reg_23), .f(n1803) );
    oai21_1 U337 ( .x(N6738), .a(n640), .b(n1777), .c(n1013) );
    nand2_2 U338 ( .x(n1777), .a(n3948), .b(n1515) );
    aoi222_1 U339 ( .x(n1013), .a(NPC[20]), .b(n1802), .c(n1732), .d(EPC_20), 
        .e(Cause_Reg_20), .f(n1803) );
    inv_2 U34 ( .x(IR_latched_9), .a(n1051) );
    mux2i_1 U340 ( .x(n3919), .d0(n1653), .sl(n1650), .d1(n1387) );
    inv_2 U341 ( .x(n1653), .a(N532) );
    oai21_1 U342 ( .x(N6736), .a(n674), .b(n678), .c(n1011) );
    nand2_2 U343 ( .x(n1082), .a(n1718), .b(IR_opcode_field[1]) );
    mux2i_1 U344 ( .x(n3920), .d0(n1652), .sl(n1650), .d1(n1390) );
    inv_2 U345 ( .x(n1652), .a(N533) );
    aoi221_1 U346 ( .x(n1129), .a(Cause_Reg_6), .b(n1803), .c(n1732), .d(EPC_6
        ), .e(n1306) );
    oai21_1 U347 ( .x(N6724), .a(n1128), .b(n678), .c(n1129) );
    oai21_1 U348 ( .x(N6737), .a(n639), .b(n995), .c(n1012) );
    mux2_4 U349 ( .x(n639), .d0(n1382), .sl(___cell__36997_net129354), .d1(
        n1383) );
    mux2i_2 U35 ( .x(n1053), .d0(current_IR_10), .sl(net149680), .d1(
        IR_latched_input[10]) );
    aoi222_1 U350 ( .x(n1012), .a(NPC[19]), .b(n1719), .c(n1732), .d(EPC_19), 
        .e(Cause_Reg_19), .f(n1803) );
    inv_2 U351 ( .x(n1410), .a(N459) );
    oai21_1 U352 ( .x(N6727), .a(n637), .b(___cell__36997_net130580), .c(n1033
        ) );
    inv_2 U353 ( .x(n1396), .a(N464) );
    mux2_4 U354 ( .x(n636), .d0(n1396), .sl(___cell__36997_net129354), .d1(
        n1397) );
    inv_5 U355 ( .x(n1001), .a(n1398) );
    oai21_1 U356 ( .x(N6730), .a(n1001), .b(___cell__36997_net130580), .c(
        n1002) );
    oai21_1 U357 ( .x(N6728), .a(n638), .b(n995), .c(n997) );
    mux2_4 U358 ( .x(n638), .d0(n1391), .sl(___cell__36997_net129354), .d1(
        n1392) );
    inv_2 U359 ( .x(n1391), .a(N458) );
    inv_4 U36 ( .x(IR_latched_3), .a(n849) );
    nand2_2 U361 ( .x(n1068), .a(n642), .b(IR_opcode_field[0]) );
    inv_2 U362 ( .x(n1386), .a(N465) );
    mux2i_1 U363 ( .x(n3918), .d0(n1654), .sl(n1650), .d1(n1397) );
    or3i_2 U364 ( .x(n681), .a(n744), .b(___cell__36997_net125928), .c(n679)
         );
    aoi222_1 U365 ( .x(n996), .a(NPC[0]), .b(n1719), .c(n1732), .d(EPC_0), .e(
        Cause_Reg_0), .f(n1803) );
    inv_5 U366 ( .x(n1031), .a(n1393) );
    oai21_1 U367 ( .x(N6726), .a(n1031), .b(n1777), .c(n1032) );
    inv_5 U368 ( .x(n1252), .a(n1388) );
    oai21_1 U369 ( .x(N6720), .a(n1252), .b(n1777), .c(n1253) );
    inv_0 U37 ( .x(n1420), .a(IR_latched_input[3]) );
    nor2_4 U370 ( .x(n1105), .a(n705), .b(n1311) );
    nor2_3 U371 ( .x(n1121), .a(n1776), .b(n696) );
    aoi222_1 U372 ( .x(n1131), .a(NPC[1]), .b(n1802), .c(n1732), .d(EPC_1), 
        .e(Cause_Reg_1), .f(n1803) );
    nand2i_2 U373 ( .x(n1064), .a(n829), .b(n1718) );
    nand2i_2 U374 ( .x(n1052), .a(n873), .b(n642) );
    nor2_1 U375 ( .x(n1117), .a(n705), .b(n765) );
    nor2_3 U376 ( .x(n1116), .a(n1776), .b(n701) );
    nor2_3 U377 ( .x(n1115), .a(n705), .b(n762) );
    nand2i_2 U378 ( .x(n1042), .a(n886), .b(n642) );
    inv_2 U379 ( .x(n1041), .a(IR_latched_3) );
    inv_14 U38 ( .x(n737), .a(n865) );
    inv_2 U380 ( .x(n1043), .a(IR_latched_4) );
    mux2i_3 U381 ( .x(IR_latched_4), .d0(n1418), .sl(net149680), .d1(n1419) );
    inv_4 U382 ( .x(counter[0]), .a(n4011) );
    ao21_1 U383 ( .x(n2640), .a(intr_slot), .b(n1092), .c(n1093) );
    nand2i_2 U384 ( .x(n1092), .a(delay_slot), .b(n1739) );
    inv_2 U385 ( .x(n1739), .a(n1267) );
    nand2i_2 U386 ( .x(n1093), .a(n1262), .b(___cell__36997_net126604) );
    oai21_1 U387 ( .x(n1034), .a(___cell__36997_net127190), .b(n1263), .c(CLI)
         );
    inv_5 U388 ( .x(___cell__36997_net130567), .a(___cell__36997_net126604) );
    mux2i_1 U389 ( .x(n2642), .d0(n627), .sl(___cell__36997_net130125), .d1(
        n813) );
    inv_0 U39 ( .x(n1040), .a(IR_latched_2) );
    mux2i_1 U390 ( .x(n2652), .d0(n617), .sl(___cell__36997_net130125), .d1(
        n4371) );
    mux2i_1 U391 ( .x(n2655), .d0(n614), .sl(___cell__36997_net130567), .d1(
        n4370) );
    mux2i_2 U392 ( .x(n2666), .d0(n603), .sl(___cell__36997_net130567), .d1(
        n654) );
    mux2i_1 U393 ( .x(n2673), .d0(n596), .sl(___cell__36997_net130567), .d1(
        n1311) );
    mux2i_1 U394 ( .x(n2674), .d0(n595), .sl(___cell__36997_net130125), .d1(
        n1553) );
    mux2i_1 U395 ( .x(n2675), .d0(n594), .sl(___cell__36997_net130567), .d1(
        n1552) );
    mux2i_1 U396 ( .x(n2676), .d0(n1294), .sl(___cell__36997_net130125), .d1(
        n1551) );
    inv_2 U397 ( .x(n1294), .a(EPC_2) );
    inv_2 U398 ( .x(n1276), .a(EPC_3) );
    mux2i_1 U399 ( .x(n2677), .d0(n1276), .sl(___cell__36997_net130567), .d1(
        n1550) );
    inv_0 U40 ( .x(n1038), .a(IR_latched_0) );
    mux2i_1 U400 ( .x(n2678), .d0(n577), .sl(___cell__36997_net130125), .d1(
        n1549) );
    mux2i_1 U401 ( .x(n2679), .d0(n576), .sl(___cell__36997_net130567), .d1(
        n1548) );
    mux2i_1 U402 ( .x(n2680), .d0(n575), .sl(___cell__36997_net130125), .d1(
        n1308) );
    mux2i_1 U403 ( .x(n2681), .d0(n574), .sl(___cell__36997_net130567), .d1(
        n1547) );
    mux2i_1 U404 ( .x(n2682), .d0(n573), .sl(___cell__36997_net130125), .d1(
        n1546) );
    mux2i_1 U405 ( .x(n2683), .d0(n572), .sl(___cell__36997_net130567), .d1(
        n1545) );
    mux2i_1 U406 ( .x(n2684), .d0(n593), .sl(___cell__36997_net130125), .d1(
        n1544) );
    mux2i_1 U407 ( .x(n2685), .d0(n592), .sl(___cell__36997_net130567), .d1(
        n1543) );
    mux2i_1 U408 ( .x(n2686), .d0(n591), .sl(___cell__36997_net130125), .d1(
        n1542) );
    mux2i_1 U409 ( .x(n2687), .d0(n590), .sl(___cell__36997_net130567), .d1(
        n1541) );
    inv_2 U41 ( .x(n824), .a(n1427) );
    mux2i_1 U410 ( .x(n2688), .d0(n589), .sl(___cell__36997_net130125), .d1(
        n1540) );
    mux2i_1 U411 ( .x(n2689), .d0(n588), .sl(___cell__36997_net130567), .d1(
        n1539) );
    mux2i_1 U412 ( .x(n2690), .d0(n587), .sl(___cell__36997_net130125), .d1(
        n1538) );
    mux2i_1 U413 ( .x(n2691), .d0(n586), .sl(___cell__36997_net130567), .d1(
        n1537) );
    mux2i_1 U414 ( .x(n2692), .d0(n585), .sl(___cell__36997_net130125), .d1(
        n1536) );
    mux2i_1 U415 ( .x(n2693), .d0(n584), .sl(___cell__36997_net130567), .d1(
        n1535) );
    mux2i_1 U416 ( .x(n2694), .d0(n583), .sl(___cell__36997_net130567), .d1(
        n1534) );
    mux2i_1 U417 ( .x(n2695), .d0(n1291), .sl(___cell__36997_net130125), .d1(
        n1533) );
    inv_2 U418 ( .x(n1291), .a(EPC_21) );
    mux2i_1 U419 ( .x(n2696), .d0(n1289), .sl(___cell__36997_net130567), .d1(
        n1532) );
    inv_2 U420 ( .x(n1289), .a(EPC_22) );
    mux2i_1 U421 ( .x(n2697), .d0(n1287), .sl(___cell__36997_net130125), .d1(
        n1531) );
    mux2i_1 U422 ( .x(n2698), .d0(n1285), .sl(___cell__36997_net130567), .d1(
        n1530) );
    inv_2 U423 ( .x(n1285), .a(EPC_24) );
    mux2i_1 U424 ( .x(n2699), .d0(n1283), .sl(___cell__36997_net130125), .d1(
        n1529) );
    mux2i_1 U425 ( .x(n2700), .d0(n582), .sl(___cell__36997_net130567), .d1(
        n1528) );
    mux2i_1 U426 ( .x(n2701), .d0(n581), .sl(___cell__36997_net130125), .d1(
        n1527) );
    mux2i_1 U427 ( .x(n2702), .d0(n580), .sl(___cell__36997_net130567), .d1(
        n1526) );
    mux2i_1 U428 ( .x(n2703), .d0(n579), .sl(___cell__36997_net130125), .d1(
        n1525) );
    mux2i_1 U429 ( .x(n2704), .d0(n662), .sl(___cell__36997_net130125), .d1(
        n1524) );
    inv_0 U43 ( .x(n805), .a(n879) );
    mux2i_1 U430 ( .x(_EPC_reg_31_net69891), .d0(n578), .sl(
        ___cell__36997_net130567), .d1(___cell__36997_net129786) );
    inv_5 U431 ( .x(___cell__36997_net130125), .a(___cell__36997_net126604) );
    nor2i_1 U432 ( .x(n1036), .a(n1260), .b(n1261) );
    mux2_2 U433 ( .x(n2709), .d0(_RegFile_31__0), .sl(n1850), .d1(WB_data[0])
         );
    mux2_2 U434 ( .x(n2710), .d0(_RegFile_31__1), .sl(n1850), .d1(WB_data[1])
         );
    mux2_2 U435 ( .x(n2711), .d0(_RegFile_31__2), .sl(n1850), .d1(WB_data[2])
         );
    mux2_2 U436 ( .x(n2712), .d0(_RegFile_31__3), .sl(n1850), .d1(WB_data[3])
         );
    mux2_2 U437 ( .x(n2713), .d0(_RegFile_31__4), .sl(n1850), .d1(WB_data[4])
         );
    mux2_2 U438 ( .x(n2714), .d0(_RegFile_31__5), .sl(n1850), .d1(WB_data[5])
         );
    mux2_2 U439 ( .x(n2715), .d0(_RegFile_31__6), .sl(n1850), .d1(WB_data[6])
         );
    and3_3 U44 ( .x(n1443), .a(n770), .b(n1693), .c(n1692) );
    mux2_2 U440 ( .x(n2716), .d0(_RegFile_31__7), .sl(n1850), .d1(WB_data[7])
         );
    mux2i_1 U441 ( .x(n2718), .d0(n2463), .sl(n1850), .d1(n1801) );
    mux2i_1 U442 ( .x(n2719), .d0(n2440), .sl(n1850), .d1(n1778) );
    mux2i_1 U443 ( .x(n2720), .d0(n2441), .sl(n1850), .d1(n1779) );
    mux2i_1 U444 ( .x(n2721), .d0(n2442), .sl(n1850), .d1(n1780) );
    mux2i_1 U445 ( .x(n2722), .d0(n2443), .sl(n1850), .d1(n1781) );
    mux2i_1 U446 ( .x(n2723), .d0(n2444), .sl(n1850), .d1(n1782) );
    mux2i_1 U447 ( .x(n2724), .d0(n2445), .sl(n1850), .d1(n1783) );
    mux2i_1 U448 ( .x(n2725), .d0(n2446), .sl(n1850), .d1(n1784) );
    mux2i_1 U449 ( .x(n2726), .d0(n2447), .sl(n1850), .d1(n1785) );
    mux2i_1 U450 ( .x(n2727), .d0(n2448), .sl(n1850), .d1(n1786) );
    mux2i_1 U451 ( .x(n2728), .d0(n2449), .sl(n1850), .d1(n1787) );
    mux2i_1 U452 ( .x(n2729), .d0(n2450), .sl(n1850), .d1(n1788) );
    mux2i_1 U453 ( .x(n2730), .d0(n2451), .sl(n1850), .d1(n1789) );
    mux2i_1 U454 ( .x(n2731), .d0(n2452), .sl(n1850), .d1(n1790) );
    mux2i_1 U455 ( .x(n2732), .d0(n2453), .sl(n1850), .d1(n1791) );
    mux2i_1 U456 ( .x(n2733), .d0(n2454), .sl(n1850), .d1(n1792) );
    mux2i_1 U457 ( .x(n2734), .d0(n2455), .sl(n1850), .d1(n1793) );
    mux2i_1 U458 ( .x(n2735), .d0(n2456), .sl(n1850), .d1(n1794) );
    mux2i_1 U459 ( .x(n2736), .d0(n2457), .sl(n1850), .d1(n1795) );
    exor2_1 U46 ( .x(n1692), .a(reg_dst_of_EX_0), .b(n884) );
    mux2i_1 U460 ( .x(n2737), .d0(n2458), .sl(n1850), .d1(n1796) );
    mux2i_1 U461 ( .x(n2738), .d0(n2459), .sl(n1850), .d1(n1797) );
    mux2i_1 U462 ( .x(n2739), .d0(n2460), .sl(n1850), .d1(n1798) );
    or2_2 U463 ( .x(n1748), .a(n3940), .b(n3944) );
    mux2_2 U464 ( .x(n2741), .d0(_RegFile_30__0), .sl(n1849), .d1(WB_data[0])
         );
    mux2_2 U465 ( .x(n2742), .d0(_RegFile_30__1), .sl(n1849), .d1(WB_data[1])
         );
    mux2_2 U466 ( .x(n2743), .d0(_RegFile_30__2), .sl(n1849), .d1(WB_data[2])
         );
    mux2_2 U467 ( .x(n2744), .d0(_RegFile_30__3), .sl(n1849), .d1(WB_data[3])
         );
    mux2_2 U468 ( .x(n2745), .d0(_RegFile_30__4), .sl(n1849), .d1(WB_data[4])
         );
    mux2_2 U469 ( .x(n2746), .d0(_RegFile_30__5), .sl(n1849), .d1(WB_data[5])
         );
    exnor2_1 U47 ( .x(n1441), .a(n772), .b(reg_dst_of_EX_3) );
    mux2_2 U470 ( .x(n2747), .d0(_RegFile_30__6), .sl(n1849), .d1(WB_data[6])
         );
    mux2_2 U471 ( .x(n2748), .d0(_RegFile_30__7), .sl(n1849), .d1(WB_data[7])
         );
    mux2i_1 U472 ( .x(n2750), .d0(n2439), .sl(n1849), .d1(n1801) );
    mux2i_1 U473 ( .x(n2751), .d0(n2416), .sl(n1849), .d1(n1778) );
    mux2i_1 U474 ( .x(n2752), .d0(n2417), .sl(n1849), .d1(n1779) );
    mux2i_1 U475 ( .x(n2753), .d0(n2418), .sl(n1849), .d1(n1780) );
    mux2i_1 U476 ( .x(n2754), .d0(n2419), .sl(n1849), .d1(n1781) );
    mux2i_1 U477 ( .x(n2755), .d0(n2420), .sl(n1849), .d1(n1782) );
    mux2i_1 U478 ( .x(n2756), .d0(n2421), .sl(n1849), .d1(n1783) );
    mux2i_1 U479 ( .x(n2757), .d0(n2422), .sl(n1849), .d1(n1784) );
    inv_2 U48 ( .x(n1584), .a(n1700) );
    mux2i_1 U480 ( .x(n2758), .d0(n2423), .sl(n1849), .d1(n1785) );
    mux2i_1 U481 ( .x(n2759), .d0(n2424), .sl(n1849), .d1(n1786) );
    mux2i_1 U482 ( .x(n2760), .d0(n2425), .sl(n1849), .d1(n1787) );
    mux2i_1 U483 ( .x(n2761), .d0(n2426), .sl(n1849), .d1(n1788) );
    mux2i_1 U484 ( .x(n2762), .d0(n2427), .sl(n1849), .d1(n1789) );
    mux2i_1 U485 ( .x(n2763), .d0(n2428), .sl(n1849), .d1(n1790) );
    mux2i_1 U486 ( .x(n2764), .d0(n2429), .sl(n1849), .d1(n1791) );
    mux2i_1 U487 ( .x(n2765), .d0(n2430), .sl(n1849), .d1(n1792) );
    mux2i_1 U488 ( .x(n2766), .d0(n2431), .sl(n1849), .d1(n1793) );
    mux2i_1 U489 ( .x(n2767), .d0(n2432), .sl(n1849), .d1(n1794) );
    nand2i_0 U49 ( .x(n1583), .a(IR_opcode_field[2]), .b(n4454) );
    mux2i_1 U490 ( .x(n2768), .d0(n2433), .sl(n1849), .d1(n1795) );
    mux2i_1 U491 ( .x(n2769), .d0(n2434), .sl(n1849), .d1(n1796) );
    mux2i_1 U492 ( .x(n2770), .d0(n2435), .sl(n1849), .d1(n1797) );
    mux2i_1 U493 ( .x(n2771), .d0(n2436), .sl(n1849), .d1(n1798) );
    buf_3 U494 ( .x(n928), .a(n987) );
    or2_2 U495 ( .x(n1749), .a(n3940), .b(n3943) );
    mux2_2 U496 ( .x(n2773), .d0(_RegFile_29__0), .sl(n1847), .d1(WB_data[0])
         );
    mux2_2 U497 ( .x(n2774), .d0(_RegFile_29__1), .sl(n1847), .d1(WB_data[1])
         );
    mux2_2 U498 ( .x(n2775), .d0(_RegFile_29__2), .sl(n1847), .d1(WB_data[2])
         );
    mux2_2 U499 ( .x(n2776), .d0(_RegFile_29__3), .sl(n1847), .d1(WB_data[3])
         );
    aoi21_1 U50 ( .x(n1582), .a(IR_opcode_field[1]), .b(n1583), .c(n1584) );
    mux2_2 U500 ( .x(n2777), .d0(_RegFile_29__4), .sl(n1847), .d1(WB_data[4])
         );
    mux2_2 U501 ( .x(n2778), .d0(_RegFile_29__5), .sl(n1847), .d1(WB_data[5])
         );
    mux2_2 U502 ( .x(n2779), .d0(_RegFile_29__6), .sl(n1847), .d1(WB_data[6])
         );
    mux2_2 U503 ( .x(n2780), .d0(_RegFile_29__7), .sl(n1847), .d1(WB_data[7])
         );
    mux2i_1 U504 ( .x(n2782), .d0(n2391), .sl(n1847), .d1(n1801) );
    mux2i_1 U505 ( .x(n2783), .d0(n2368), .sl(n1847), .d1(n1778) );
    mux2i_1 U506 ( .x(n2784), .d0(n2369), .sl(n1847), .d1(n1779) );
    mux2i_1 U507 ( .x(n2785), .d0(n2370), .sl(n1847), .d1(n1780) );
    mux2i_1 U508 ( .x(n2786), .d0(n2371), .sl(n1847), .d1(n1781) );
    mux2i_1 U509 ( .x(n2787), .d0(n2372), .sl(n1847), .d1(n1782) );
    nand2i_2 U51 ( .x(n1585), .a(n1320), .b(n1586) );
    mux2i_1 U510 ( .x(n2788), .d0(n2373), .sl(n1847), .d1(n1783) );
    mux2i_1 U511 ( .x(n2789), .d0(n2374), .sl(n1847), .d1(n1784) );
    mux2i_1 U512 ( .x(n2790), .d0(n2375), .sl(n1847), .d1(n1785) );
    mux2i_1 U513 ( .x(n2791), .d0(n2376), .sl(n1847), .d1(n1786) );
    mux2i_1 U514 ( .x(n2792), .d0(n2377), .sl(n1847), .d1(n1787) );
    mux2i_1 U515 ( .x(n2793), .d0(n2378), .sl(n1847), .d1(n1788) );
    mux2i_1 U516 ( .x(n2794), .d0(n2379), .sl(n1847), .d1(n1789) );
    mux2i_1 U517 ( .x(n2795), .d0(n2380), .sl(n1847), .d1(n1790) );
    mux2i_1 U518 ( .x(n2796), .d0(n2381), .sl(n1847), .d1(n1791) );
    mux2i_1 U519 ( .x(n2797), .d0(n2382), .sl(n1847), .d1(n1792) );
    nor2i_1 U52 ( .x(n1320), .a(n1321), .b(n1322) );
    mux2i_1 U520 ( .x(n2798), .d0(n2383), .sl(n1847), .d1(n1793) );
    mux2i_1 U521 ( .x(n2799), .d0(n2384), .sl(n1847), .d1(n1794) );
    mux2i_1 U522 ( .x(n2800), .d0(n2385), .sl(n1847), .d1(n1795) );
    mux2i_1 U523 ( .x(n2801), .d0(n2386), .sl(n1847), .d1(n1796) );
    mux2i_1 U524 ( .x(n2802), .d0(n2387), .sl(n1847), .d1(n1797) );
    mux2i_1 U525 ( .x(n2803), .d0(n2388), .sl(n1847), .d1(n1798) );
    or2_2 U526 ( .x(n1751), .a(n3940), .b(n3942) );
    mux2_2 U527 ( .x(n2805), .d0(_RegFile_28__0), .sl(n1846), .d1(WB_data[0])
         );
    mux2_2 U528 ( .x(n2806), .d0(_RegFile_28__1), .sl(n1846), .d1(WB_data[1])
         );
    mux2_2 U529 ( .x(n2807), .d0(_RegFile_28__2), .sl(n1846), .d1(WB_data[2])
         );
    mux2i_1 U53 ( .x(n1586), .d0(n1580), .sl(IR_opcode_field[1]), .d1(n1581)
         );
    mux2_2 U530 ( .x(n2808), .d0(_RegFile_28__3), .sl(n1846), .d1(WB_data[3])
         );
    mux2_2 U531 ( .x(n2809), .d0(_RegFile_28__4), .sl(n1846), .d1(WB_data[4])
         );
    mux2_2 U532 ( .x(n2810), .d0(_RegFile_28__5), .sl(n1846), .d1(WB_data[5])
         );
    mux2_2 U533 ( .x(n2811), .d0(_RegFile_28__6), .sl(n1846), .d1(WB_data[6])
         );
    mux2_2 U534 ( .x(n2812), .d0(_RegFile_28__7), .sl(n1846), .d1(WB_data[7])
         );
    mux2i_1 U535 ( .x(n2814), .d0(n2367), .sl(n1846), .d1(n1801) );
    mux2i_1 U536 ( .x(n2815), .d0(n2344), .sl(n1846), .d1(n1778) );
    mux2i_1 U537 ( .x(n2816), .d0(n2345), .sl(n1846), .d1(n1779) );
    mux2i_1 U538 ( .x(n2817), .d0(n2346), .sl(n1846), .d1(n1780) );
    mux2i_1 U539 ( .x(n2818), .d0(n2347), .sl(n1846), .d1(n1781) );
    inv_10 U54 ( .x(___cell__36997_net129477), .a(n331) );
    mux2i_1 U540 ( .x(n2819), .d0(n2348), .sl(n1846), .d1(n1782) );
    mux2i_1 U541 ( .x(n2820), .d0(n2349), .sl(n1846), .d1(n1783) );
    mux2i_1 U542 ( .x(n2821), .d0(n2350), .sl(n1846), .d1(n1784) );
    mux2i_1 U543 ( .x(n2822), .d0(n2351), .sl(n1846), .d1(n1785) );
    mux2i_1 U544 ( .x(n2823), .d0(n2352), .sl(n1846), .d1(n1786) );
    mux2i_1 U545 ( .x(n2824), .d0(n2353), .sl(n1846), .d1(n1787) );
    mux2i_1 U546 ( .x(n2825), .d0(n2354), .sl(n1846), .d1(n1788) );
    mux2i_1 U547 ( .x(n2826), .d0(n2355), .sl(n1846), .d1(n1789) );
    mux2i_1 U548 ( .x(n2827), .d0(n2356), .sl(n1846), .d1(n1790) );
    mux2i_1 U549 ( .x(n2828), .d0(n2357), .sl(n1846), .d1(n1791) );
    exor2_1 U55 ( .x(___cell__36997_net129979), .a(WB_index_0), .b(n879) );
    mux2i_1 U550 ( .x(n2829), .d0(n2358), .sl(n1846), .d1(n1792) );
    mux2i_1 U551 ( .x(n2830), .d0(n2359), .sl(n1846), .d1(n1793) );
    mux2i_1 U552 ( .x(n2831), .d0(n2360), .sl(n1846), .d1(n1794) );
    mux2i_1 U553 ( .x(n2832), .d0(n2361), .sl(n1846), .d1(n1795) );
    mux2i_1 U554 ( .x(n2833), .d0(n2362), .sl(n1846), .d1(n1796) );
    mux2i_1 U555 ( .x(n2834), .d0(n2363), .sl(n1846), .d1(n1797) );
    mux2i_1 U556 ( .x(n2835), .d0(n2364), .sl(n1846), .d1(n1798) );
    buf_3 U557 ( .x(n931), .a(n987) );
    or2_2 U558 ( .x(n1752), .a(n3940), .b(n3941) );
    mux2_2 U559 ( .x(n2837), .d0(_RegFile_27__0), .sl(n1845), .d1(WB_data[0])
         );
    buf_3 U56 ( .x(n715), .a(n332) );
    mux2_2 U560 ( .x(n2838), .d0(_RegFile_27__1), .sl(n1845), .d1(WB_data[1])
         );
    mux2_2 U561 ( .x(n2839), .d0(_RegFile_27__2), .sl(n1845), .d1(WB_data[2])
         );
    mux2_2 U562 ( .x(n2840), .d0(_RegFile_27__3), .sl(n1845), .d1(WB_data[3])
         );
    mux2_2 U563 ( .x(n2841), .d0(_RegFile_27__4), .sl(n1845), .d1(WB_data[4])
         );
    mux2_2 U564 ( .x(n2842), .d0(_RegFile_27__5), .sl(n1845), .d1(WB_data[5])
         );
    mux2_2 U565 ( .x(n2843), .d0(_RegFile_27__6), .sl(n1845), .d1(WB_data[6])
         );
    mux2_2 U566 ( .x(n2844), .d0(_RegFile_27__7), .sl(n1845), .d1(WB_data[7])
         );
    mux2i_1 U567 ( .x(n2846), .d0(n2343), .sl(n1845), .d1(n1801) );
    mux2i_1 U568 ( .x(n2847), .d0(n2320), .sl(n1845), .d1(n1778) );
    mux2i_1 U569 ( .x(n2848), .d0(n2321), .sl(n1845), .d1(n1779) );
    inv_5 U57 ( .x(___cell__36997_net130306), .a(n709) );
    mux2i_1 U570 ( .x(n2849), .d0(n2322), .sl(n1845), .d1(n1780) );
    mux2i_1 U571 ( .x(n2850), .d0(n2323), .sl(n1845), .d1(n1781) );
    mux2i_1 U572 ( .x(n2851), .d0(n2324), .sl(n1845), .d1(n1782) );
    mux2i_1 U573 ( .x(n2852), .d0(n2325), .sl(n1845), .d1(n1783) );
    mux2i_1 U574 ( .x(n2853), .d0(n2326), .sl(n1845), .d1(n1784) );
    mux2i_1 U575 ( .x(n2854), .d0(n2327), .sl(n1845), .d1(n1785) );
    mux2i_1 U576 ( .x(n2855), .d0(n2328), .sl(n1845), .d1(n1786) );
    mux2i_1 U577 ( .x(n2856), .d0(n2329), .sl(n1845), .d1(n1787) );
    mux2i_1 U578 ( .x(n2857), .d0(n2330), .sl(n1845), .d1(n1788) );
    mux2i_1 U579 ( .x(n2858), .d0(n2331), .sl(n1845), .d1(n1789) );
    mux2i_1 U58 ( .x(n1452), .d0(n628), .sl(opcode_of_MEM_5), .d1(n1579) );
    mux2i_1 U580 ( .x(n2859), .d0(n2332), .sl(n1845), .d1(n1790) );
    mux2i_1 U581 ( .x(n2860), .d0(n2333), .sl(n1845), .d1(n1791) );
    mux2i_1 U582 ( .x(n2861), .d0(n2334), .sl(n1845), .d1(n1792) );
    mux2i_1 U583 ( .x(n2862), .d0(n2335), .sl(n1845), .d1(n1793) );
    mux2i_1 U584 ( .x(n2863), .d0(n2336), .sl(n1845), .d1(n1794) );
    mux2i_1 U585 ( .x(n2864), .d0(n2337), .sl(n1845), .d1(n1795) );
    mux2i_1 U586 ( .x(n2865), .d0(n2338), .sl(n1845), .d1(n1796) );
    mux2i_1 U587 ( .x(n2866), .d0(n2339), .sl(n1845), .d1(n1797) );
    mux2i_1 U588 ( .x(n2867), .d0(n2340), .sl(n1845), .d1(n1798) );
    or2_2 U589 ( .x(n1753), .a(n3939), .b(n3944) );
    nand2i_2 U59 ( .x(n1478), .a(opcode_of_MEM_1), .b(n1690) );
    mux2_2 U590 ( .x(n2869), .d0(_RegFile_26__0), .sl(n1844), .d1(WB_data[0])
         );
    mux2_2 U591 ( .x(n2870), .d0(_RegFile_26__1), .sl(n1844), .d1(WB_data[1])
         );
    mux2_2 U592 ( .x(n2871), .d0(_RegFile_26__2), .sl(n1844), .d1(WB_data[2])
         );
    mux2_2 U593 ( .x(n2872), .d0(_RegFile_26__3), .sl(n1844), .d1(WB_data[3])
         );
    mux2_2 U594 ( .x(n2873), .d0(_RegFile_26__4), .sl(n1844), .d1(WB_data[4])
         );
    mux2_2 U595 ( .x(n2874), .d0(_RegFile_26__5), .sl(n1844), .d1(WB_data[5])
         );
    mux2_2 U596 ( .x(n2875), .d0(_RegFile_26__6), .sl(n1844), .d1(WB_data[6])
         );
    mux2_2 U597 ( .x(n2876), .d0(_RegFile_26__7), .sl(n1844), .d1(WB_data[7])
         );
    mux2i_1 U598 ( .x(n2878), .d0(n2319), .sl(n1844), .d1(n1801) );
    mux2i_1 U599 ( .x(n2879), .d0(n2296), .sl(n1844), .d1(n1778) );
    inv_2 U60 ( .x(n1690), .a(n1450) );
    mux2i_1 U600 ( .x(n2880), .d0(n2297), .sl(n1844), .d1(n1779) );
    mux2i_1 U601 ( .x(n2881), .d0(n2298), .sl(n1844), .d1(n1780) );
    mux2i_1 U602 ( .x(n2882), .d0(n2299), .sl(n1844), .d1(n1781) );
    mux2i_1 U603 ( .x(n2883), .d0(n2300), .sl(n1844), .d1(n1782) );
    mux2i_1 U604 ( .x(n2884), .d0(n2301), .sl(n1844), .d1(n1783) );
    mux2i_1 U605 ( .x(n2885), .d0(n2302), .sl(n1844), .d1(n1784) );
    mux2i_1 U606 ( .x(n2886), .d0(n2303), .sl(n1844), .d1(n1785) );
    mux2i_1 U607 ( .x(n2887), .d0(n2304), .sl(n1844), .d1(n1786) );
    mux2i_1 U608 ( .x(n2888), .d0(n2305), .sl(n1844), .d1(n1787) );
    mux2i_1 U609 ( .x(n2889), .d0(n2306), .sl(n1844), .d1(n1788) );
    nand2i_2 U61 ( .x(n1450), .a(opcode_of_MEM_5), .b(opcode_of_MEM_3) );
    mux2i_1 U610 ( .x(n2890), .d0(n2307), .sl(n1844), .d1(n1789) );
    mux2i_1 U611 ( .x(n2891), .d0(n2308), .sl(n1844), .d1(n1790) );
    mux2i_1 U612 ( .x(n2892), .d0(n2309), .sl(n1844), .d1(n1791) );
    mux2i_1 U613 ( .x(n2893), .d0(n2310), .sl(n1844), .d1(n1792) );
    mux2i_1 U614 ( .x(n2894), .d0(n2311), .sl(n1844), .d1(n1793) );
    mux2i_1 U615 ( .x(n2895), .d0(n2312), .sl(n1844), .d1(n1794) );
    mux2i_1 U616 ( .x(n2896), .d0(n2313), .sl(n1844), .d1(n1795) );
    mux2i_1 U617 ( .x(n2897), .d0(n2314), .sl(n1844), .d1(n1796) );
    mux2i_1 U618 ( .x(n2898), .d0(n2315), .sl(n1844), .d1(n1797) );
    mux2i_1 U619 ( .x(n2899), .d0(n2316), .sl(n1844), .d1(n1798) );
    and3i_3 U62 ( .x(n1458), .a(n667), .b(n1567), .c(n1566) );
    buf_3 U620 ( .x(n933), .a(n961) );
    or2_2 U621 ( .x(n1754), .a(n3939), .b(n3943) );
    mux2_2 U622 ( .x(n2901), .d0(_RegFile_25__0), .sl(n1843), .d1(WB_data[0])
         );
    mux2_2 U623 ( .x(n2902), .d0(_RegFile_25__1), .sl(n1843), .d1(WB_data[1])
         );
    mux2_2 U624 ( .x(n2903), .d0(_RegFile_25__2), .sl(n1843), .d1(WB_data[2])
         );
    mux2_2 U625 ( .x(n2904), .d0(_RegFile_25__3), .sl(n1843), .d1(WB_data[3])
         );
    mux2_2 U626 ( .x(n2905), .d0(_RegFile_25__4), .sl(n1843), .d1(WB_data[4])
         );
    mux2_2 U627 ( .x(n2906), .d0(_RegFile_25__5), .sl(n1843), .d1(WB_data[5])
         );
    mux2_2 U628 ( .x(n2907), .d0(_RegFile_25__6), .sl(n1843), .d1(WB_data[6])
         );
    mux2_2 U629 ( .x(n2908), .d0(_RegFile_25__7), .sl(n1843), .d1(WB_data[7])
         );
    exnor2_2 U63 ( .x(n1456), .a(n337), .b(n634) );
    mux2i_1 U630 ( .x(n2910), .d0(n2295), .sl(n1843), .d1(n1801) );
    mux2i_1 U631 ( .x(n2911), .d0(n2272), .sl(n1843), .d1(n1778) );
    mux2i_1 U632 ( .x(n2912), .d0(n2273), .sl(n1843), .d1(n1779) );
    mux2i_1 U633 ( .x(n2913), .d0(n2274), .sl(n1843), .d1(n1780) );
    mux2i_1 U634 ( .x(n2914), .d0(n2275), .sl(n1843), .d1(n1781) );
    mux2i_1 U635 ( .x(n2915), .d0(n2276), .sl(n1843), .d1(n1782) );
    mux2i_1 U636 ( .x(n2916), .d0(n2277), .sl(n1843), .d1(n1783) );
    mux2i_1 U637 ( .x(n2917), .d0(n2278), .sl(n1843), .d1(n1784) );
    mux2i_1 U638 ( .x(n2918), .d0(n2279), .sl(n1843), .d1(n1785) );
    mux2i_1 U639 ( .x(n2919), .d0(n2280), .sl(n1843), .d1(n1786) );
    nand2i_2 U64 ( .x(n1723), .a(n3888), .b(WB_data[7]) );
    mux2i_1 U640 ( .x(n2920), .d0(n2281), .sl(n1843), .d1(n1787) );
    mux2i_1 U641 ( .x(n2921), .d0(n2282), .sl(n1843), .d1(n1788) );
    mux2i_1 U642 ( .x(n2922), .d0(n2283), .sl(n1843), .d1(n1789) );
    mux2i_1 U643 ( .x(n2923), .d0(n2284), .sl(n1843), .d1(n1790) );
    mux2i_1 U644 ( .x(n2924), .d0(n2285), .sl(n1843), .d1(n1791) );
    mux2i_1 U645 ( .x(n2925), .d0(n2286), .sl(n1843), .d1(n1792) );
    mux2i_1 U646 ( .x(n2926), .d0(n2287), .sl(n1843), .d1(n1793) );
    mux2i_1 U647 ( .x(n2927), .d0(n2288), .sl(n1843), .d1(n1794) );
    mux2i_1 U648 ( .x(n2928), .d0(n2289), .sl(n1843), .d1(n1795) );
    mux2i_1 U649 ( .x(n2929), .d0(n2290), .sl(n1843), .d1(n1796) );
    nand2i_2 U65 ( .x(n1305), .a(n3888), .b(N13832) );
    mux2i_1 U650 ( .x(n2930), .d0(n2291), .sl(n1843), .d1(n1797) );
    mux2i_1 U651 ( .x(n2931), .d0(n2292), .sl(n1843), .d1(n1798) );
    or2_2 U652 ( .x(n1755), .a(n3939), .b(n3942) );
    mux2_2 U653 ( .x(n2933), .d0(_RegFile_24__0), .sl(n1842), .d1(WB_data[0])
         );
    mux2_2 U654 ( .x(n2934), .d0(_RegFile_24__1), .sl(n1842), .d1(WB_data[1])
         );
    mux2_2 U655 ( .x(n2935), .d0(_RegFile_24__2), .sl(n1842), .d1(WB_data[2])
         );
    mux2_2 U656 ( .x(n2936), .d0(_RegFile_24__3), .sl(n1842), .d1(WB_data[3])
         );
    mux2_2 U657 ( .x(n2937), .d0(_RegFile_24__4), .sl(n1842), .d1(WB_data[4])
         );
    mux2_2 U658 ( .x(n2938), .d0(_RegFile_24__5), .sl(n1842), .d1(WB_data[5])
         );
    mux2_2 U659 ( .x(n2939), .d0(_RegFile_24__6), .sl(n1842), .d1(WB_data[6])
         );
    inv_4 U66 ( .x(n881), .a(n1434) );
    mux2_2 U660 ( .x(n2940), .d0(_RegFile_24__7), .sl(n1842), .d1(WB_data[7])
         );
    mux2i_1 U661 ( .x(n2942), .d0(n2271), .sl(n1842), .d1(n1801) );
    mux2i_1 U662 ( .x(n2943), .d0(n2248), .sl(n1842), .d1(n1778) );
    mux2i_1 U663 ( .x(n2944), .d0(n2249), .sl(n1842), .d1(n1779) );
    mux2i_1 U664 ( .x(n2945), .d0(n2250), .sl(n1842), .d1(n1780) );
    mux2i_1 U665 ( .x(n2946), .d0(n2251), .sl(n1842), .d1(n1781) );
    mux2i_1 U666 ( .x(n2947), .d0(n2252), .sl(n1842), .d1(n1782) );
    mux2i_1 U667 ( .x(n2948), .d0(n2253), .sl(n1842), .d1(n1783) );
    mux2i_1 U668 ( .x(n2949), .d0(n2254), .sl(n1842), .d1(n1784) );
    mux2i_1 U669 ( .x(n2950), .d0(n2255), .sl(n1842), .d1(n1785) );
    nand2i_2 U67 ( .x(n1470), .a(n724), .b(n1517) );
    mux2i_1 U670 ( .x(n2951), .d0(n2256), .sl(n1842), .d1(n1786) );
    mux2i_1 U671 ( .x(n2952), .d0(n2257), .sl(n1842), .d1(n1787) );
    mux2i_1 U672 ( .x(n2953), .d0(n2258), .sl(n1842), .d1(n1788) );
    mux2i_1 U673 ( .x(n2954), .d0(n2259), .sl(n1842), .d1(n1789) );
    mux2i_1 U674 ( .x(n2955), .d0(n2260), .sl(n1842), .d1(n1790) );
    mux2i_1 U675 ( .x(n2956), .d0(n2261), .sl(n1842), .d1(n1791) );
    mux2i_1 U676 ( .x(n2957), .d0(n2262), .sl(n1842), .d1(n1792) );
    mux2i_1 U677 ( .x(n2958), .d0(n2263), .sl(n1842), .d1(n1793) );
    mux2i_1 U678 ( .x(n2959), .d0(n2264), .sl(n1842), .d1(n1794) );
    mux2i_1 U679 ( .x(n2960), .d0(n2265), .sl(n1842), .d1(n1795) );
    mux2i_1 U68 ( .x(n1460), .d0(FREEZE), .sl(delay_slot), .d1(n1576) );
    mux2i_1 U680 ( .x(n2961), .d0(n2266), .sl(n1842), .d1(n1796) );
    mux2i_1 U681 ( .x(n2962), .d0(n2267), .sl(n1842), .d1(n1797) );
    mux2i_1 U682 ( .x(n2963), .d0(n2268), .sl(n1842), .d1(n1798) );
    or2_2 U683 ( .x(n1756), .a(n3939), .b(n3941) );
    mux2_2 U684 ( .x(n2965), .d0(_RegFile_23__0), .sl(n1841), .d1(WB_data[0])
         );
    mux2_2 U685 ( .x(n2966), .d0(_RegFile_23__1), .sl(n1841), .d1(WB_data[1])
         );
    mux2_2 U686 ( .x(n2967), .d0(_RegFile_23__2), .sl(n1841), .d1(n686) );
    mux2_2 U687 ( .x(n2968), .d0(_RegFile_23__3), .sl(n1841), .d1(n685) );
    mux2_2 U688 ( .x(n2969), .d0(_RegFile_23__4), .sl(n1841), .d1(WB_data[4])
         );
    mux2_2 U689 ( .x(n2970), .d0(_RegFile_23__5), .sl(n1841), .d1(WB_data[5])
         );
    nand2_0 U69 ( .x(n1715), .a(n807), .b(n1462) );
    mux2_2 U690 ( .x(n2971), .d0(_RegFile_23__6), .sl(n1841), .d1(WB_data[6])
         );
    mux2_2 U691 ( .x(n2972), .d0(_RegFile_23__7), .sl(n1841), .d1(WB_data[7])
         );
    mux2i_1 U692 ( .x(n2974), .d0(n2247), .sl(n1841), .d1(n1801) );
    mux2i_1 U693 ( .x(n2975), .d0(n2224), .sl(n1841), .d1(n1778) );
    mux2i_1 U694 ( .x(n2976), .d0(n2225), .sl(n1841), .d1(n1779) );
    mux2i_1 U695 ( .x(n2977), .d0(n2226), .sl(n1841), .d1(n1780) );
    mux2i_1 U696 ( .x(n2978), .d0(n2227), .sl(n1841), .d1(n1781) );
    mux2i_1 U697 ( .x(n2979), .d0(n2228), .sl(n1841), .d1(n1782) );
    mux2i_1 U698 ( .x(n2980), .d0(n2229), .sl(n1841), .d1(n1783) );
    mux2i_1 U699 ( .x(n2981), .d0(n2230), .sl(n1841), .d1(n1784) );
    mux2i_1 U70 ( .x(n1265), .d0(n1312), .sl(n1454), .d1(n1591) );
    mux2i_1 U700 ( .x(n2982), .d0(n2231), .sl(n1841), .d1(n1785) );
    mux2i_1 U701 ( .x(n2983), .d0(n2232), .sl(n1841), .d1(n1786) );
    mux2i_1 U702 ( .x(n2984), .d0(n2233), .sl(n1841), .d1(n1787) );
    mux2i_1 U703 ( .x(n2985), .d0(n2234), .sl(n1841), .d1(n1788) );
    mux2i_1 U704 ( .x(n2986), .d0(n2235), .sl(n1841), .d1(n1789) );
    mux2i_1 U705 ( .x(n2987), .d0(n2236), .sl(n1841), .d1(n1790) );
    mux2i_1 U706 ( .x(n2988), .d0(n2237), .sl(n1841), .d1(n1791) );
    mux2i_1 U707 ( .x(n2989), .d0(n2238), .sl(n1841), .d1(n1792) );
    mux2i_1 U708 ( .x(n2990), .d0(n2239), .sl(n1841), .d1(n1793) );
    mux2i_1 U709 ( .x(n2991), .d0(n2240), .sl(n1841), .d1(n1794) );
    inv_5 U71 ( .x(n1454), .a(n1440) );
    mux2i_1 U710 ( .x(n2992), .d0(n2241), .sl(n1841), .d1(n1795) );
    mux2i_1 U711 ( .x(n2993), .d0(n2242), .sl(n1841), .d1(n1796) );
    mux2i_1 U712 ( .x(n2994), .d0(n2243), .sl(n1841), .d1(n1797) );
    mux2i_1 U713 ( .x(n2995), .d0(n2244), .sl(n1841), .d1(n1798) );
    or2_2 U714 ( .x(n1757), .a(n3938), .b(n3944) );
    mux2_2 U715 ( .x(n2997), .d0(_RegFile_22__0), .sl(n1840), .d1(WB_data[0])
         );
    mux2_2 U716 ( .x(n2998), .d0(_RegFile_22__1), .sl(n1840), .d1(WB_data[1])
         );
    mux2_2 U717 ( .x(n2999), .d0(_RegFile_22__2), .sl(n1840), .d1(WB_data[2])
         );
    mux2_2 U718 ( .x(n3000), .d0(_RegFile_22__3), .sl(n1840), .d1(WB_data[3])
         );
    mux2_2 U719 ( .x(n3001), .d0(_RegFile_22__4), .sl(n1840), .d1(WB_data[4])
         );
    nor2_1 U72 ( .x(n1720), .a(n1492), .b(n1484) );
    mux2_2 U720 ( .x(n3002), .d0(_RegFile_22__5), .sl(n1840), .d1(WB_data[5])
         );
    mux2_2 U721 ( .x(n3003), .d0(_RegFile_22__6), .sl(n1840), .d1(WB_data[6])
         );
    mux2_2 U722 ( .x(n3004), .d0(_RegFile_22__7), .sl(n1840), .d1(WB_data[7])
         );
    mux2i_1 U723 ( .x(n3006), .d0(n2223), .sl(n1840), .d1(n1801) );
    mux2i_1 U724 ( .x(n3007), .d0(n2200), .sl(n1840), .d1(n1778) );
    mux2i_1 U725 ( .x(n3008), .d0(n2201), .sl(n1840), .d1(n1779) );
    mux2i_1 U726 ( .x(n3009), .d0(n2202), .sl(n1840), .d1(n1780) );
    mux2i_1 U727 ( .x(n3010), .d0(n2203), .sl(n1840), .d1(n1781) );
    mux2i_1 U728 ( .x(n3011), .d0(n2204), .sl(n1840), .d1(n1782) );
    mux2i_1 U729 ( .x(n3012), .d0(n2205), .sl(n1840), .d1(n1783) );
    nand2i_2 U73 ( .x(n1721), .a(___cell__36997_net125928), .b(n1720) );
    mux2i_1 U730 ( .x(n3013), .d0(n2206), .sl(n1840), .d1(n1784) );
    mux2i_1 U731 ( .x(n3014), .d0(n2207), .sl(n1840), .d1(n1785) );
    mux2i_1 U732 ( .x(n3015), .d0(n2208), .sl(n1840), .d1(n1786) );
    mux2i_1 U733 ( .x(n3016), .d0(n2209), .sl(n1840), .d1(n1787) );
    mux2i_1 U734 ( .x(n3017), .d0(n2210), .sl(n1840), .d1(n1788) );
    mux2i_1 U735 ( .x(n3018), .d0(n2211), .sl(n1840), .d1(n1789) );
    mux2i_1 U736 ( .x(n3019), .d0(n2212), .sl(n1840), .d1(n1790) );
    mux2i_1 U737 ( .x(n3020), .d0(n2213), .sl(n1840), .d1(n1791) );
    mux2i_1 U738 ( .x(n3021), .d0(n2214), .sl(n1840), .d1(n1792) );
    mux2i_1 U739 ( .x(n3022), .d0(n2215), .sl(n1840), .d1(n1793) );
    inv_2 U74 ( .x(n1057), .a(IR_latched_12) );
    mux2i_1 U740 ( .x(n3023), .d0(n2216), .sl(n1840), .d1(n1794) );
    mux2i_1 U741 ( .x(n3024), .d0(n2217), .sl(n1840), .d1(n1795) );
    mux2i_1 U742 ( .x(n3025), .d0(n2218), .sl(n1840), .d1(n1796) );
    mux2i_1 U743 ( .x(n3026), .d0(n2219), .sl(n1840), .d1(n1797) );
    mux2i_1 U744 ( .x(n3027), .d0(n2220), .sl(n1840), .d1(n1798) );
    or2_2 U745 ( .x(n1758), .a(n3938), .b(n3943) );
    mux2_2 U746 ( .x(n3029), .d0(_RegFile_21__0), .sl(n1839), .d1(WB_data[0])
         );
    mux2_2 U747 ( .x(n3030), .d0(_RegFile_21__1), .sl(n1839), .d1(WB_data[1])
         );
    mux2_2 U748 ( .x(n3031), .d0(_RegFile_21__2), .sl(n1839), .d1(WB_data[2])
         );
    mux2_2 U749 ( .x(n3032), .d0(_RegFile_21__3), .sl(n1839), .d1(WB_data[3])
         );
    inv_2 U75 ( .x(n1498), .a(N5379) );
    mux2_2 U750 ( .x(n3033), .d0(_RegFile_21__4), .sl(n1839), .d1(WB_data[4])
         );
    mux2_2 U751 ( .x(n3034), .d0(_RegFile_21__5), .sl(n1839), .d1(WB_data[5])
         );
    mux2_2 U752 ( .x(n3035), .d0(_RegFile_21__6), .sl(n1839), .d1(WB_data[6])
         );
    mux2_2 U753 ( .x(n3036), .d0(_RegFile_21__7), .sl(n1839), .d1(WB_data[7])
         );
    mux2i_1 U754 ( .x(n3038), .d0(n2199), .sl(n1839), .d1(n1801) );
    mux2i_1 U755 ( .x(n3039), .d0(n2176), .sl(n1839), .d1(n1778) );
    mux2i_1 U756 ( .x(n3040), .d0(n2177), .sl(n1839), .d1(n1779) );
    mux2i_1 U757 ( .x(n3041), .d0(n2178), .sl(n1839), .d1(n1780) );
    mux2i_1 U758 ( .x(n3042), .d0(n2179), .sl(n1839), .d1(n1781) );
    mux2i_1 U759 ( .x(n3043), .d0(n2180), .sl(n1839), .d1(n1782) );
    nand2i_2 U76 ( .x(n1587), .a(n557), .b(n1738) );
    mux2i_1 U760 ( .x(n3044), .d0(n2181), .sl(n1839), .d1(n1783) );
    mux2i_1 U761 ( .x(n3045), .d0(n2182), .sl(n1839), .d1(n1784) );
    mux2i_1 U762 ( .x(n3046), .d0(n2183), .sl(n1839), .d1(n1785) );
    mux2i_1 U763 ( .x(n3047), .d0(n2184), .sl(n1839), .d1(n1786) );
    mux2i_1 U764 ( .x(n3048), .d0(n2185), .sl(n1839), .d1(n1787) );
    mux2i_1 U765 ( .x(n3049), .d0(n2186), .sl(n1839), .d1(n1788) );
    mux2i_1 U766 ( .x(n3050), .d0(n2187), .sl(n1839), .d1(n1789) );
    mux2i_1 U767 ( .x(n3051), .d0(n2188), .sl(n1839), .d1(n1790) );
    mux2i_1 U768 ( .x(n3052), .d0(n2189), .sl(n1839), .d1(n1791) );
    mux2i_1 U769 ( .x(n3053), .d0(n2190), .sl(n1839), .d1(n1792) );
    nand2i_2 U77 ( .x(n1589), .a(___cell__36997_net130681), .b(n1738) );
    mux2i_1 U770 ( .x(n3054), .d0(n2191), .sl(n1839), .d1(n1793) );
    mux2i_1 U771 ( .x(n3055), .d0(n2192), .sl(n1839), .d1(n1794) );
    mux2i_1 U772 ( .x(n3056), .d0(n2193), .sl(n1839), .d1(n1795) );
    mux2i_1 U773 ( .x(n3057), .d0(n2194), .sl(n1839), .d1(n1796) );
    mux2i_1 U774 ( .x(n3058), .d0(n2195), .sl(n1839), .d1(n1797) );
    buf_3 U775 ( .x(n965), .a(n952) );
    mux2i_1 U776 ( .x(n3059), .d0(n2196), .sl(n1839), .d1(n1798) );
    or2_2 U777 ( .x(n1759), .a(n3938), .b(n3942) );
    mux2_2 U778 ( .x(n3061), .d0(_RegFile_20__0), .sl(n1838), .d1(WB_data[0])
         );
    mux2_2 U779 ( .x(n3062), .d0(_RegFile_20__1), .sl(n1838), .d1(WB_data[1])
         );
    nand2i_2 U78 ( .x(n1588), .a(n557), .b(n1472) );
    mux2_2 U780 ( .x(n3063), .d0(_RegFile_20__2), .sl(n1838), .d1(WB_data[2])
         );
    mux2_2 U781 ( .x(n3064), .d0(_RegFile_20__3), .sl(n1838), .d1(WB_data[3])
         );
    mux2_2 U782 ( .x(n3065), .d0(_RegFile_20__4), .sl(n1838), .d1(WB_data[4])
         );
    mux2_2 U783 ( .x(n3066), .d0(_RegFile_20__5), .sl(n1838), .d1(WB_data[5])
         );
    mux2_2 U784 ( .x(n3067), .d0(_RegFile_20__6), .sl(n1838), .d1(WB_data[6])
         );
    mux2_2 U785 ( .x(n3068), .d0(_RegFile_20__7), .sl(n1838), .d1(WB_data[7])
         );
    mux2i_1 U786 ( .x(n3070), .d0(n2175), .sl(n1838), .d1(n1801) );
    mux2i_1 U787 ( .x(n3071), .d0(n2152), .sl(n1838), .d1(n1778) );
    mux2i_1 U788 ( .x(n3072), .d0(n2153), .sl(n1838), .d1(n1779) );
    mux2i_1 U789 ( .x(n3073), .d0(n2154), .sl(n1838), .d1(n1780) );
    or2_2 U79 ( .x(n1472), .a(intr_slot), .b(delay_slot) );
    mux2i_1 U790 ( .x(n3074), .d0(n2155), .sl(n1838), .d1(n1781) );
    mux2i_1 U791 ( .x(n3075), .d0(n2156), .sl(n1838), .d1(n1782) );
    mux2i_1 U792 ( .x(n3076), .d0(n2157), .sl(n1838), .d1(n1783) );
    mux2i_1 U793 ( .x(n3077), .d0(n2158), .sl(n1838), .d1(n1784) );
    mux2i_1 U794 ( .x(n3078), .d0(n2159), .sl(n1838), .d1(n1785) );
    mux2i_1 U795 ( .x(n3079), .d0(n2160), .sl(n1838), .d1(n1786) );
    mux2i_1 U796 ( .x(n3080), .d0(n2161), .sl(n1838), .d1(n1787) );
    mux2i_1 U797 ( .x(n3081), .d0(n2162), .sl(n1838), .d1(n1788) );
    mux2i_1 U798 ( .x(n3082), .d0(n2163), .sl(n1838), .d1(n1789) );
    mux2i_1 U799 ( .x(n3083), .d0(n2164), .sl(n1838), .d1(n1790) );
    inv_2 U80 ( .x(n1738), .a(n1472) );
    mux2i_1 U800 ( .x(n3084), .d0(n2165), .sl(n1838), .d1(n1791) );
    mux2i_1 U801 ( .x(n3085), .d0(n2166), .sl(n1838), .d1(n1792) );
    mux2i_1 U802 ( .x(n3086), .d0(n2167), .sl(n1838), .d1(n1793) );
    mux2i_1 U803 ( .x(n3087), .d0(n2168), .sl(n1838), .d1(n1794) );
    mux2i_1 U804 ( .x(n3088), .d0(n2169), .sl(n1838), .d1(n1795) );
    mux2i_1 U805 ( .x(n3089), .d0(n2170), .sl(n1838), .d1(n1796) );
    mux2i_1 U806 ( .x(n3090), .d0(n2171), .sl(n1838), .d1(n1797) );
    mux2i_1 U807 ( .x(n3091), .d0(n2172), .sl(n1838), .d1(n1798) );
    or2_2 U808 ( .x(n1760), .a(n3938), .b(n3941) );
    mux2_2 U809 ( .x(n3093), .d0(_RegFile_19__0), .sl(n1836), .d1(WB_data[0])
         );
    inv_2 U81 ( .x(n1298), .a(N6035) );
    mux2_2 U810 ( .x(n3094), .d0(_RegFile_19__1), .sl(n1836), .d1(WB_data[1])
         );
    mux2_2 U811 ( .x(n3095), .d0(_RegFile_19__2), .sl(n1836), .d1(WB_data[2])
         );
    mux2_2 U812 ( .x(n3096), .d0(_RegFile_19__3), .sl(n1836), .d1(WB_data[3])
         );
    mux2_2 U813 ( .x(n3097), .d0(_RegFile_19__4), .sl(n1836), .d1(WB_data[4])
         );
    mux2_2 U814 ( .x(n3098), .d0(_RegFile_19__5), .sl(n1836), .d1(WB_data[5])
         );
    mux2_2 U815 ( .x(n3099), .d0(_RegFile_19__6), .sl(n1836), .d1(WB_data[6])
         );
    mux2_2 U816 ( .x(n3100), .d0(_RegFile_19__7), .sl(n1836), .d1(WB_data[7])
         );
    mux2i_1 U817 ( .x(n3102), .d0(n2127), .sl(n1836), .d1(n1801) );
    mux2i_1 U818 ( .x(n3103), .d0(n2104), .sl(n1836), .d1(n1778) );
    mux2i_1 U819 ( .x(n3104), .d0(n2105), .sl(n1836), .d1(n1779) );
    nor2_1 U82 ( .x(n1297), .a(___cell__36997_net129239), .b(n1298) );
    mux2i_1 U820 ( .x(n3105), .d0(n2106), .sl(n1836), .d1(n1780) );
    mux2i_1 U821 ( .x(n3106), .d0(n2107), .sl(n1836), .d1(n1781) );
    mux2i_1 U822 ( .x(n3107), .d0(n2108), .sl(n1836), .d1(n1782) );
    mux2i_1 U823 ( .x(n3108), .d0(n2109), .sl(n1836), .d1(n1783) );
    mux2i_1 U824 ( .x(n3109), .d0(n2110), .sl(n1836), .d1(n1784) );
    mux2i_1 U825 ( .x(n3110), .d0(n2111), .sl(n1836), .d1(n1785) );
    mux2i_1 U826 ( .x(n3111), .d0(n2112), .sl(n1836), .d1(n1786) );
    mux2i_1 U827 ( .x(n3112), .d0(n2113), .sl(n1836), .d1(n1787) );
    mux2i_1 U828 ( .x(n3113), .d0(n2114), .sl(n1836), .d1(n1788) );
    mux2i_1 U829 ( .x(n3114), .d0(n2115), .sl(n1836), .d1(n1789) );
    nor2i_1 U83 ( .x(n1301), .a(N6018), .b(___cell__36997_net129239) );
    mux2i_1 U830 ( .x(n3115), .d0(n2116), .sl(n1836), .d1(n1790) );
    mux2i_1 U831 ( .x(n3116), .d0(n2117), .sl(n1836), .d1(n1791) );
    mux2i_1 U832 ( .x(n3117), .d0(n2118), .sl(n1836), .d1(n1792) );
    mux2i_1 U833 ( .x(n3118), .d0(n2119), .sl(n1836), .d1(n1793) );
    mux2i_1 U834 ( .x(n3119), .d0(n2120), .sl(n1836), .d1(n1794) );
    mux2i_1 U835 ( .x(n3120), .d0(n2121), .sl(n1836), .d1(n1795) );
    mux2i_1 U836 ( .x(n3121), .d0(n2122), .sl(n1836), .d1(n1796) );
    mux2i_1 U837 ( .x(n3122), .d0(n2123), .sl(n1836), .d1(n1797) );
    mux2i_1 U838 ( .x(n3123), .d0(n2124), .sl(n1836), .d1(n1798) );
    buf_3 U839 ( .x(n940), .a(n961) );
    inv_2 U84 ( .x(n1508), .a(N5373) );
    or2_2 U840 ( .x(n1762), .a(n3934), .b(n3944) );
    mux2_2 U841 ( .x(n3125), .d0(_RegFile_18__0), .sl(n1835), .d1(WB_data[0])
         );
    mux2_2 U842 ( .x(n3126), .d0(_RegFile_18__1), .sl(n1835), .d1(WB_data[1])
         );
    mux2_2 U843 ( .x(n3127), .d0(_RegFile_18__2), .sl(n1835), .d1(WB_data[2])
         );
    mux2_2 U844 ( .x(n3128), .d0(_RegFile_18__3), .sl(n1835), .d1(WB_data[3])
         );
    mux2_2 U845 ( .x(n3129), .d0(_RegFile_18__4), .sl(n1835), .d1(WB_data[4])
         );
    mux2_2 U846 ( .x(n3130), .d0(_RegFile_18__5), .sl(n1835), .d1(WB_data[5])
         );
    mux2_2 U847 ( .x(n3131), .d0(_RegFile_18__6), .sl(n1835), .d1(WB_data[6])
         );
    mux2_2 U848 ( .x(n3132), .d0(_RegFile_18__7), .sl(n1835), .d1(WB_data[7])
         );
    mux2i_1 U849 ( .x(n3134), .d0(n2103), .sl(n1835), .d1(n1801) );
    mux2i_1 U850 ( .x(n3135), .d0(n2080), .sl(n1835), .d1(n1778) );
    mux2i_1 U851 ( .x(n3136), .d0(n2081), .sl(n1835), .d1(n1779) );
    mux2i_1 U852 ( .x(n3137), .d0(n2082), .sl(n1835), .d1(n1780) );
    mux2i_1 U853 ( .x(n3138), .d0(n2083), .sl(n1835), .d1(n1781) );
    mux2i_1 U854 ( .x(n3139), .d0(n2084), .sl(n1835), .d1(n1782) );
    mux2i_1 U855 ( .x(n3140), .d0(n2085), .sl(n1835), .d1(n1783) );
    mux2i_1 U856 ( .x(n3141), .d0(n2086), .sl(n1835), .d1(n1784) );
    mux2i_1 U857 ( .x(n3142), .d0(n2087), .sl(n1835), .d1(n1785) );
    mux2i_1 U858 ( .x(n3143), .d0(n2088), .sl(n1835), .d1(n1786) );
    mux2i_1 U859 ( .x(n3144), .d0(n2089), .sl(n1835), .d1(n1787) );
    mux2i_1 U860 ( .x(n3145), .d0(n2090), .sl(n1835), .d1(n1788) );
    mux2i_1 U861 ( .x(n3146), .d0(n2091), .sl(n1835), .d1(n1789) );
    mux2i_1 U862 ( .x(n3147), .d0(n2092), .sl(n1835), .d1(n1790) );
    mux2i_1 U863 ( .x(n3148), .d0(n2093), .sl(n1835), .d1(n1791) );
    mux2i_1 U864 ( .x(n3149), .d0(n2094), .sl(n1835), .d1(n1792) );
    mux2i_1 U865 ( .x(n3150), .d0(n2095), .sl(n1835), .d1(n1793) );
    mux2i_1 U866 ( .x(n3151), .d0(n2096), .sl(n1835), .d1(n1794) );
    mux2i_1 U867 ( .x(n3152), .d0(n2097), .sl(n1835), .d1(n1795) );
    mux2i_1 U868 ( .x(n3153), .d0(n2098), .sl(n1835), .d1(n1796) );
    mux2i_1 U869 ( .x(n3154), .d0(n2099), .sl(n1835), .d1(n1797) );
    mux2i_1 U870 ( .x(n3155), .d0(n2100), .sl(n1835), .d1(n1798) );
    buf_3 U871 ( .x(n941), .a(n961) );
    or2_2 U872 ( .x(n1763), .a(n3934), .b(n3943) );
    mux2_2 U873 ( .x(n3157), .d0(_RegFile_17__0), .sl(n1834), .d1(WB_data[0])
         );
    mux2_2 U874 ( .x(n3158), .d0(_RegFile_17__1), .sl(n1834), .d1(WB_data[1])
         );
    mux2_2 U875 ( .x(n3159), .d0(_RegFile_17__2), .sl(n1834), .d1(WB_data[2])
         );
    mux2_2 U876 ( .x(n3160), .d0(_RegFile_17__3), .sl(n1834), .d1(WB_data[3])
         );
    mux2_2 U877 ( .x(n3161), .d0(_RegFile_17__4), .sl(n1834), .d1(WB_data[4])
         );
    mux2_2 U878 ( .x(n3162), .d0(_RegFile_17__5), .sl(n1834), .d1(WB_data[5])
         );
    mux2_2 U879 ( .x(n3163), .d0(_RegFile_17__6), .sl(n1834), .d1(WB_data[6])
         );
    inv_2 U88 ( .x(___cell__36997_net129388), .a(N437) );
    mux2_2 U880 ( .x(n3164), .d0(_RegFile_17__7), .sl(n1834), .d1(WB_data[7])
         );
    mux2i_1 U881 ( .x(n3166), .d0(n2079), .sl(n1834), .d1(n1801) );
    mux2i_1 U882 ( .x(n3167), .d0(n2056), .sl(n1834), .d1(n1778) );
    mux2i_1 U883 ( .x(n3168), .d0(n2057), .sl(n1834), .d1(n1779) );
    mux2i_1 U884 ( .x(n3169), .d0(n2058), .sl(n1834), .d1(n1780) );
    mux2i_1 U885 ( .x(n3170), .d0(n2059), .sl(n1834), .d1(n1781) );
    mux2i_1 U886 ( .x(n3171), .d0(n2060), .sl(n1834), .d1(n1782) );
    mux2i_1 U887 ( .x(n3172), .d0(n2061), .sl(n1834), .d1(n1783) );
    mux2i_1 U888 ( .x(n3173), .d0(n2062), .sl(n1834), .d1(n1784) );
    mux2i_1 U889 ( .x(n3174), .d0(n2063), .sl(n1834), .d1(n1785) );
    mux2i_1 U890 ( .x(n3175), .d0(n2064), .sl(n1834), .d1(n1786) );
    mux2i_1 U891 ( .x(n3176), .d0(n2065), .sl(n1834), .d1(n1787) );
    mux2i_1 U892 ( .x(n3177), .d0(n2066), .sl(n1834), .d1(n1788) );
    mux2i_1 U893 ( .x(n3178), .d0(n2067), .sl(n1834), .d1(n1789) );
    mux2i_1 U894 ( .x(n3179), .d0(n2068), .sl(n1834), .d1(n1790) );
    mux2i_1 U895 ( .x(n3180), .d0(n2069), .sl(n1834), .d1(n1791) );
    mux2i_1 U896 ( .x(n3181), .d0(n2070), .sl(n1834), .d1(n1792) );
    mux2i_1 U897 ( .x(n3182), .d0(n2071), .sl(n1834), .d1(n1793) );
    mux2i_1 U898 ( .x(n3183), .d0(n2072), .sl(n1834), .d1(n1794) );
    mux2i_1 U899 ( .x(n3184), .d0(n2073), .sl(n1834), .d1(n1795) );
    nand2i_2 U90 ( .x(n793), .a(n578), .b(n799) );
    mux2i_1 U900 ( .x(n3185), .d0(n2074), .sl(n1834), .d1(n1796) );
    mux2i_1 U901 ( .x(n3186), .d0(n2075), .sl(n1834), .d1(n1797) );
    mux2i_1 U902 ( .x(n3187), .d0(n2076), .sl(n1834), .d1(n1798) );
    buf_3 U903 ( .x(n942), .a(n934) );
    or2_2 U904 ( .x(n1764), .a(n3934), .b(n3942) );
    mux2_2 U905 ( .x(n3189), .d0(_RegFile_16__0), .sl(n1833), .d1(WB_data[0])
         );
    mux2_2 U906 ( .x(n3190), .d0(_RegFile_16__1), .sl(n1833), .d1(WB_data[1])
         );
    mux2_2 U907 ( .x(n3191), .d0(_RegFile_16__2), .sl(n1833), .d1(WB_data[2])
         );
    mux2_2 U908 ( .x(n3192), .d0(_RegFile_16__3), .sl(n1833), .d1(WB_data[3])
         );
    mux2_2 U909 ( .x(n3193), .d0(_RegFile_16__4), .sl(n1833), .d1(WB_data[4])
         );
    mux2_2 U910 ( .x(n3194), .d0(_RegFile_16__5), .sl(n1833), .d1(WB_data[5])
         );
    mux2_2 U911 ( .x(n3195), .d0(_RegFile_16__6), .sl(n1833), .d1(WB_data[6])
         );
    mux2_2 U912 ( .x(n3196), .d0(_RegFile_16__7), .sl(n1833), .d1(WB_data[7])
         );
    mux2i_1 U913 ( .x(n3198), .d0(n2055), .sl(n1833), .d1(n1801) );
    mux2i_1 U914 ( .x(n3199), .d0(n2032), .sl(n1833), .d1(n1778) );
    mux2i_1 U915 ( .x(n3200), .d0(n2033), .sl(n1833), .d1(n1779) );
    mux2i_1 U916 ( .x(n3201), .d0(n2034), .sl(n1833), .d1(n1780) );
    mux2i_1 U917 ( .x(n3202), .d0(n2035), .sl(n1833), .d1(n1781) );
    mux2i_1 U918 ( .x(n3203), .d0(n2036), .sl(n1833), .d1(n1782) );
    mux2i_1 U919 ( .x(n3204), .d0(n2037), .sl(n1833), .d1(n1783) );
    nor2_1 U92 ( .x(n1259), .a(delay_slot), .b(n2639) );
    mux2i_1 U920 ( .x(n3205), .d0(n2038), .sl(n1833), .d1(n1784) );
    mux2i_1 U921 ( .x(n3206), .d0(n2039), .sl(n1833), .d1(n1785) );
    mux2i_1 U922 ( .x(n3207), .d0(n2040), .sl(n1833), .d1(n1786) );
    mux2i_1 U923 ( .x(n3208), .d0(n2041), .sl(n1833), .d1(n1787) );
    mux2i_1 U924 ( .x(n3209), .d0(n2042), .sl(n1833), .d1(n1788) );
    mux2i_1 U925 ( .x(n3210), .d0(n2043), .sl(n1833), .d1(n1789) );
    mux2i_1 U926 ( .x(n3211), .d0(n2044), .sl(n1833), .d1(n1790) );
    mux2i_1 U927 ( .x(n3212), .d0(n2045), .sl(n1833), .d1(n1791) );
    mux2i_1 U928 ( .x(n3213), .d0(n2046), .sl(n1833), .d1(n1792) );
    mux2i_1 U929 ( .x(n3214), .d0(n2047), .sl(n1833), .d1(n1793) );
    ao21_3 U93 ( .x(n1590), .a(n1448), .b(n861), .c(n755) );
    mux2i_1 U930 ( .x(n3215), .d0(n2048), .sl(n1833), .d1(n1794) );
    mux2i_1 U931 ( .x(n3216), .d0(n2049), .sl(n1833), .d1(n1795) );
    mux2i_1 U932 ( .x(n3217), .d0(n2050), .sl(n1833), .d1(n1796) );
    mux2i_1 U933 ( .x(n3218), .d0(n2051), .sl(n1833), .d1(n1797) );
    mux2i_1 U934 ( .x(n3219), .d0(n2052), .sl(n1833), .d1(n1798) );
    buf_3 U935 ( .x(n943), .a(n934) );
    or2_2 U936 ( .x(n1765), .a(n3934), .b(n3941) );
    mux2_2 U937 ( .x(n3221), .d0(_RegFile_15__0), .sl(n1832), .d1(WB_data[0])
         );
    mux2_2 U938 ( .x(n3222), .d0(_RegFile_15__1), .sl(n1832), .d1(WB_data[1])
         );
    mux2_2 U939 ( .x(n3223), .d0(_RegFile_15__2), .sl(n1832), .d1(WB_data[2])
         );
    inv_4 U94 ( .x(n1356), .a(N440) );
    mux2_2 U940 ( .x(n3224), .d0(_RegFile_15__3), .sl(n1832), .d1(WB_data[3])
         );
    mux2_2 U941 ( .x(n3225), .d0(_RegFile_15__4), .sl(n1832), .d1(WB_data[4])
         );
    mux2_2 U942 ( .x(n3226), .d0(_RegFile_15__5), .sl(n1832), .d1(WB_data[5])
         );
    mux2_2 U943 ( .x(n3227), .d0(_RegFile_15__6), .sl(n1832), .d1(WB_data[6])
         );
    mux2_2 U944 ( .x(n3228), .d0(_RegFile_15__7), .sl(n1832), .d1(WB_data[7])
         );
    buf_3 U945 ( .x(n960), .a(n985) );
    mux2i_1 U946 ( .x(n3230), .d0(n2031), .sl(n1832), .d1(n1801) );
    mux2i_1 U947 ( .x(n3231), .d0(n2008), .sl(n1832), .d1(n1778) );
    mux2i_1 U948 ( .x(n3232), .d0(n2009), .sl(n1832), .d1(n1779) );
    mux2i_1 U949 ( .x(n3233), .d0(n2010), .sl(n1832), .d1(n1780) );
    inv_2 U95 ( .x(n1402), .a(N445) );
    mux2i_1 U950 ( .x(n3234), .d0(n2011), .sl(n1832), .d1(n1781) );
    mux2i_1 U951 ( .x(n3235), .d0(n2012), .sl(n1832), .d1(n1782) );
    mux2i_1 U952 ( .x(n3236), .d0(n2013), .sl(n1832), .d1(n1783) );
    mux2i_1 U953 ( .x(n3237), .d0(n2014), .sl(n1832), .d1(n1784) );
    mux2i_1 U954 ( .x(n3238), .d0(n2015), .sl(n1832), .d1(n1785) );
    mux2i_1 U955 ( .x(n3239), .d0(n2016), .sl(n1832), .d1(n1786) );
    mux2i_1 U956 ( .x(n3240), .d0(n2017), .sl(n1832), .d1(n1787) );
    mux2i_1 U957 ( .x(n3241), .d0(n2018), .sl(n1832), .d1(n1788) );
    mux2i_1 U958 ( .x(n3242), .d0(n2019), .sl(n1832), .d1(n1789) );
    mux2i_1 U959 ( .x(n3243), .d0(n2020), .sl(n1832), .d1(n1790) );
    inv_2 U96 ( .x(n1380), .a(N448) );
    mux2i_1 U960 ( .x(n3244), .d0(n2021), .sl(n1832), .d1(n1791) );
    mux2i_1 U961 ( .x(n3245), .d0(n2022), .sl(n1832), .d1(n1792) );
    mux2i_1 U962 ( .x(n3246), .d0(n2023), .sl(n1832), .d1(n1793) );
    mux2i_1 U963 ( .x(n3247), .d0(n2024), .sl(n1832), .d1(n1794) );
    mux2i_1 U964 ( .x(n3248), .d0(n2025), .sl(n1832), .d1(n1795) );
    mux2i_1 U965 ( .x(n3249), .d0(n2026), .sl(n1832), .d1(n1796) );
    mux2i_1 U966 ( .x(n3250), .d0(n2027), .sl(n1832), .d1(n1797) );
    mux2i_1 U967 ( .x(n3251), .d0(n2028), .sl(n1832), .d1(n1798) );
    buf_3 U968 ( .x(n944), .a(n934) );
    or2_2 U969 ( .x(n1766), .a(n3937), .b(n3940) );
    inv_5 U97 ( .x(n1719), .a(n1307) );
    mux2_2 U970 ( .x(n3253), .d0(_RegFile_14__0), .sl(n1831), .d1(WB_data[0])
         );
    mux2_2 U971 ( .x(n3254), .d0(_RegFile_14__1), .sl(n1831), .d1(WB_data[1])
         );
    mux2_2 U972 ( .x(n3255), .d0(_RegFile_14__2), .sl(n1831), .d1(WB_data[2])
         );
    mux2_2 U973 ( .x(n3256), .d0(_RegFile_14__3), .sl(n1831), .d1(WB_data[3])
         );
    mux2_2 U974 ( .x(n3257), .d0(_RegFile_14__4), .sl(n1831), .d1(WB_data[4])
         );
    mux2_2 U975 ( .x(n3258), .d0(_RegFile_14__5), .sl(n1831), .d1(WB_data[5])
         );
    mux2_2 U976 ( .x(n3259), .d0(_RegFile_14__6), .sl(n1831), .d1(WB_data[6])
         );
    mux2_2 U977 ( .x(n3260), .d0(_RegFile_14__7), .sl(n1831), .d1(WB_data[7])
         );
    mux2i_1 U978 ( .x(n3262), .d0(n2007), .sl(n1831), .d1(n1801) );
    mux2i_1 U979 ( .x(n3263), .d0(n1984), .sl(n1831), .d1(n1778) );
    nand2_1 U98 ( .x(n1307), .a(n1468), .b(___cell__36997_net126612) );
    mux2i_1 U980 ( .x(n3264), .d0(n1985), .sl(n1831), .d1(n1779) );
    mux2i_1 U981 ( .x(n3265), .d0(n1986), .sl(n1831), .d1(n1780) );
    mux2i_1 U982 ( .x(n3266), .d0(n1987), .sl(n1831), .d1(n1781) );
    mux2i_1 U983 ( .x(n3267), .d0(n1988), .sl(n1831), .d1(n1782) );
    mux2i_1 U984 ( .x(n3268), .d0(n1989), .sl(n1831), .d1(n1783) );
    mux2i_1 U985 ( .x(n3269), .d0(n1990), .sl(n1831), .d1(n1784) );
    mux2i_1 U986 ( .x(n3270), .d0(n1991), .sl(n1831), .d1(n1785) );
    mux2i_1 U987 ( .x(n3271), .d0(n1992), .sl(n1831), .d1(n1786) );
    mux2i_1 U988 ( .x(n3272), .d0(n1993), .sl(n1831), .d1(n1787) );
    mux2i_1 U989 ( .x(n3273), .d0(n1994), .sl(n1831), .d1(n1788) );
    nor2_1 U99 ( .x(n1306), .a(n1307), .b(n1308) );
    mux2i_1 U990 ( .x(n3274), .d0(n1995), .sl(n1831), .d1(n1789) );
    mux2i_1 U991 ( .x(n3275), .d0(n1996), .sl(n1831), .d1(n1790) );
    mux2i_1 U992 ( .x(n3276), .d0(n1997), .sl(n1831), .d1(n1791) );
    mux2i_1 U993 ( .x(n3277), .d0(n1998), .sl(n1831), .d1(n1792) );
    mux2i_1 U994 ( .x(n3278), .d0(n1999), .sl(n1831), .d1(n1793) );
    mux2i_1 U995 ( .x(n3279), .d0(n2000), .sl(n1831), .d1(n1794) );
    mux2i_1 U996 ( .x(n3280), .d0(n2001), .sl(n1831), .d1(n1795) );
    mux2i_1 U997 ( .x(n3281), .d0(n2002), .sl(n1831), .d1(n1796) );
    mux2i_1 U998 ( .x(n3282), .d0(n2003), .sl(n1831), .d1(n1797) );
    mux2i_1 U999 ( .x(n3283), .d0(n2004), .sl(n1831), .d1(n1798) );
    smlatnr_1 WB_index_reg_0__master ( .q(WB_index_reg_0__m2s), .d(
        reg_dst_of_MEM_0), .sdi(n2461), .se(test_se), .g(Ctrl__Regs_1__en1), 
        .rb(n913), .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 WB_index_reg_0__slave ( .q(WB_index_0), .qb(n3928), .d(
        WB_index_reg_0__m2s), .g(Ctrl__Regs_1__en2), .rb(n913), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 WB_index_reg_1__master ( .q(WB_index_reg_1__m2s), .d(
        reg_dst_of_MEM_1), .sdi(n3928), .se(test_se), .g(Ctrl__Regs_1__en1), 
        .rb(n912), .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 WB_index_reg_1__slave ( .q(WB_index_1), .qb(n3929), .d(
        WB_index_reg_1__m2s), .g(Ctrl__Regs_1__en2), .rb(n912), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 WB_index_reg_2__master ( .q(WB_index_reg_2__m2s), .d(
        reg_dst_of_MEM_2), .sdi(n3929), .se(test_se), .g(Ctrl__Regs_1__en1), 
        .rb(n913), .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 WB_index_reg_2__slave ( .q(WB_index_2), .qb(n3925), .d(
        WB_index_reg_2__m2s), .g(Ctrl__Regs_1__en2), .rb(n913), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 WB_index_reg_3__master ( .q(WB_index_reg_3__m2s), .d(
        reg_dst_of_MEM_3), .sdi(n3925), .se(test_se), .g(Ctrl__Regs_1__en1), 
        .rb(n913), .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 WB_index_reg_3__slave ( .q(WB_index_3), .qb(n3926), .d(
        WB_index_reg_3__m2s), .g(Ctrl__Regs_1__en2), .rb(n913), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 WB_index_reg_4__master ( .q(WB_index_reg_4__m2s), .d(
        reg_dst_of_MEM_4), .sdi(WB_index_3), .se(test_se), .g(
        Ctrl__Regs_1__en1), .rb(n913), .glob_g(global_g1), .sync_sel(sync_sel)
         );
    mlatnr_2 WB_index_reg_4__slave ( .q(WB_index_4), .qb(
        ___cell__6171_net27367), .d(WB_index_reg_4__m2s), .g(Ctrl__Regs_1__en2
        ), .rb(n913), .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_0__0__master ( .q(_RegFile_reg_0__0__m2s), .d(n3701
        ), .sdi(n4369), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n955), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_0__0__slave ( .q(_RegFile_0__0), .qb(n4368), .d(
        _RegFile_reg_0__0__m2s), .g(Ctrl__Regs_1__en2), .rb(n955), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_0__10__master ( .q(_RegFile_reg_0__10__m2s), .d(
        n3711), .sdi(n1887), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n955), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_0__10__slave ( .q(_RegFile_0__10), .qb(n1864), .d(
        _RegFile_reg_0__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n955), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_0__11__master ( .q(_RegFile_reg_0__11__m2s), .d(
        n3712), .sdi(n1864), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_0__11__slave ( .q(_RegFile_0__11), .qb(n1865), .d(
        _RegFile_reg_0__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_0__12__master ( .q(_RegFile_reg_0__12__m2s), .d(
        n3713), .sdi(n1865), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n955), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_0__12__slave ( .q(_RegFile_0__12), .qb(n1866), .d(
        _RegFile_reg_0__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n955), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_0__13__master ( .q(_RegFile_reg_0__13__m2s), .d(
        n3714), .sdi(n1866), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_0__13__slave ( .q(_RegFile_0__13), .qb(n1867), .d(
        _RegFile_reg_0__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_0__14__master ( .q(_RegFile_reg_0__14__m2s), .d(
        n3715), .sdi(n1867), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n955), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_0__14__slave ( .q(_RegFile_0__14), .qb(n1868), .d(
        _RegFile_reg_0__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n955), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_0__15__master ( .q(_RegFile_reg_0__15__m2s), .d(
        n3716), .sdi(n1868), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_0__15__slave ( .q(_RegFile_0__15), .qb(n1869), .d(
        _RegFile_reg_0__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_0__16__master ( .q(_RegFile_reg_0__16__m2s), .d(
        n3717), .sdi(n1869), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n956), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_0__16__slave ( .q(_RegFile_0__16), .qb(n1870), .d(
        _RegFile_reg_0__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n956), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_0__17__master ( .q(_RegFile_reg_0__17__m2s), .d(
        n3718), .sdi(n1870), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_0__17__slave ( .q(_RegFile_0__17), .qb(n1871), .d(
        _RegFile_reg_0__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_0__18__master ( .q(_RegFile_reg_0__18__m2s), .d(
        n3719), .sdi(n1871), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n956), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_0__18__slave ( .q(_RegFile_0__18), .qb(n1872), .d(
        _RegFile_reg_0__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n956), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_0__19__master ( .q(_RegFile_reg_0__19__m2s), .d(
        n3720), .sdi(n1872), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_0__19__slave ( .q(_RegFile_0__19), .qb(n1873), .d(
        _RegFile_reg_0__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_0__1__master ( .q(_RegFile_reg_0__1__m2s), .d(n3702
        ), .sdi(n4368), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_0__1__slave ( .q(_RegFile_0__1), .qb(n4367), .d(
        _RegFile_reg_0__1__m2s), .g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_0__20__master ( .q(_RegFile_reg_0__20__m2s), .d(
        n3721), .sdi(n1873), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_0__20__slave ( .q(_RegFile_0__20), .qb(n1874), .d(
        _RegFile_reg_0__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_0__21__master ( .q(_RegFile_reg_0__21__m2s), .d(
        n3722), .sdi(n1874), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n956), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_0__21__slave ( .q(_RegFile_0__21), .qb(n1875), .d(
        _RegFile_reg_0__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n956), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_0__22__master ( .q(_RegFile_reg_0__22__m2s), .d(
        n3723), .sdi(n1875), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_0__22__slave ( .q(_RegFile_0__22), .qb(n1876), .d(
        _RegFile_reg_0__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_0__23__master ( .q(_RegFile_reg_0__23__m2s), .d(
        n3724), .sdi(n1876), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n956), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_0__23__slave ( .q(_RegFile_0__23), .qb(n1877), .d(
        _RegFile_reg_0__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n956), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_0__24__master ( .q(_RegFile_reg_0__24__m2s), .d(
        n3725), .sdi(n1877), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_0__24__slave ( .q(_RegFile_0__24), .qb(n1878), .d(
        _RegFile_reg_0__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_0__25__master ( .q(_RegFile_reg_0__25__m2s), .d(
        n3726), .sdi(n1878), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n956), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_0__25__slave ( .q(_RegFile_0__25), .qb(n1879), .d(
        _RegFile_reg_0__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n956), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_0__26__master ( .q(_RegFile_reg_0__26__m2s), .d(
        n3727), .sdi(n1879), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_0__26__slave ( .q(_RegFile_0__26), .qb(n1880), .d(
        _RegFile_reg_0__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_0__27__master ( .q(_RegFile_reg_0__27__m2s), .d(
        n3728), .sdi(n1880), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n956), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_0__27__slave ( .q(_RegFile_0__27), .qb(n1881), .d(
        _RegFile_reg_0__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n956), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_0__28__master ( .q(_RegFile_reg_0__28__m2s), .d(
        n3729), .sdi(n1881), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_0__28__slave ( .q(_RegFile_0__28), .qb(n1882), .d(
        _RegFile_reg_0__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_0__29__master ( .q(_RegFile_reg_0__29__m2s), .d(
        n3730), .sdi(n1882), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n956), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_0__29__slave ( .q(_RegFile_0__29), .qb(n1883), .d(
        _RegFile_reg_0__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n956), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_0__2__master ( .q(_RegFile_reg_0__2__m2s), .d(n3703
        ), .sdi(n4367), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n956), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_0__2__slave ( .q(_RegFile_0__2), .qb(n4366), .d(
        _RegFile_reg_0__2__m2s), .g(Ctrl__Regs_1__en2), .rb(n956), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_0__30__master ( .q(_RegFile_reg_0__30__m2s), .d(
        n3731), .sdi(n1883), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n956), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_0__30__slave ( .q(_RegFile_0__30), .qb(n1884), .d(
        _RegFile_reg_0__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n956), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_0__31__master ( .q(_RegFile_reg_0__31__m2s), .d(
        n3732), .sdi(n1884), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_0__31__slave ( .q(_RegFile_0__31), .qb(n1885), .d(
        _RegFile_reg_0__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_0__3__master ( .q(_RegFile_reg_0__3__m2s), .d(n3704
        ), .sdi(n4366), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_0__3__slave ( .q(_RegFile_0__3), .qb(n4365), .d(
        _RegFile_reg_0__3__m2s), .g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_0__4__master ( .q(_RegFile_reg_0__4__m2s), .d(n3705
        ), .sdi(n4365), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n956), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_0__4__slave ( .q(_RegFile_0__4), .qb(n4364), .d(
        _RegFile_reg_0__4__m2s), .g(Ctrl__Regs_1__en2), .rb(n956), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_0__5__master ( .q(_RegFile_reg_0__5__m2s), .d(n3706
        ), .sdi(n4364), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_0__5__slave ( .q(_RegFile_0__5), .qb(n4363), .d(
        _RegFile_reg_0__5__m2s), .g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_0__6__master ( .q(_RegFile_reg_0__6__m2s), .d(n3707
        ), .sdi(n4363), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n956), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_0__6__slave ( .q(_RegFile_0__6), .qb(n4362), .d(
        _RegFile_reg_0__6__m2s), .g(Ctrl__Regs_1__en2), .rb(n956), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_0__7__master ( .q(_RegFile_reg_0__7__m2s), .d(n3708
        ), .sdi(n4362), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_0__7__slave ( .q(_RegFile_0__7), .qb(n4361), .d(
        _RegFile_reg_0__7__m2s), .g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_0__8__master ( .q(_RegFile_reg_0__8__m2s), .d(n3709
        ), .sdi(n4361), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n956), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_0__8__slave ( .q(_RegFile_0__8), .qb(n1886), .d(
        _RegFile_reg_0__8__m2s), .g(Ctrl__Regs_1__en2), .rb(n956), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_0__9__master ( .q(_RegFile_reg_0__9__m2s), .d(n3710
        ), .sdi(n1886), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_0__9__slave ( .q(_RegFile_0__9), .qb(n1887), .d(
        _RegFile_reg_0__9__m2s), .g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_10__0__master ( .q(_RegFile_reg_10__0__m2s), .d(
        n3381), .sdi(n2629), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n956), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_10__0__slave ( .q(_RegFile_10__0), .qb(n4288), .d(
        _RegFile_reg_10__0__m2s), .g(Ctrl__Regs_1__en2), .rb(n956), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_10__10__master ( .q(_RegFile_reg_10__10__m2s), .d(
        n3391), .sdi(n1911), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n956), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_10__10__slave ( .q(_RegFile_10__10), .qb(n1888), .d(
        _RegFile_reg_10__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n956), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_10__11__master ( .q(_RegFile_reg_10__11__m2s), .d(
        n3392), .sdi(n1888), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_10__11__slave ( .q(_RegFile_10__11), .qb(n1889), .d(
        _RegFile_reg_10__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_10__12__master ( .q(_RegFile_reg_10__12__m2s), .d(
        n3393), .sdi(n1889), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n956), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_10__12__slave ( .q(_RegFile_10__12), .qb(n1890), .d(
        _RegFile_reg_10__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n956), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_10__13__master ( .q(_RegFile_reg_10__13__m2s), .d(
        n3394), .sdi(n1890), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_10__13__slave ( .q(_RegFile_10__13), .qb(n1891), .d(
        _RegFile_reg_10__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_10__14__master ( .q(_RegFile_reg_10__14__m2s), .d(
        n3395), .sdi(n1891), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n957), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_10__14__slave ( .q(_RegFile_10__14), .qb(n1892), .d(
        _RegFile_reg_10__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n957), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_10__15__master ( .q(_RegFile_reg_10__15__m2s), .d(
        n3396), .sdi(n1892), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_10__15__slave ( .q(_RegFile_10__15), .qb(n1893), .d(
        _RegFile_reg_10__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_10__16__master ( .q(_RegFile_reg_10__16__m2s), .d(
        n3397), .sdi(n1893), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n957), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_10__16__slave ( .q(_RegFile_10__16), .qb(n1894), .d(
        _RegFile_reg_10__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n957), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_10__17__master ( .q(_RegFile_reg_10__17__m2s), .d(
        n3398), .sdi(n1894), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_10__17__slave ( .q(_RegFile_10__17), .qb(n1895), .d(
        _RegFile_reg_10__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_10__18__master ( .q(_RegFile_reg_10__18__m2s), .d(
        n3399), .sdi(n1895), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n957), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_10__18__slave ( .q(_RegFile_10__18), .qb(n1896), .d(
        _RegFile_reg_10__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n957), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_10__19__master ( .q(_RegFile_reg_10__19__m2s), .d(
        n3400), .sdi(n1896), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_10__19__slave ( .q(_RegFile_10__19), .qb(n1897), .d(
        _RegFile_reg_10__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_10__1__master ( .q(_RegFile_reg_10__1__m2s), .d(
        n3382), .sdi(n4288), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_10__1__slave ( .q(_RegFile_10__1), .qb(n4287), .d(
        _RegFile_reg_10__1__m2s), .g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_10__20__master ( .q(_RegFile_reg_10__20__m2s), .d(
        n3401), .sdi(n1897), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_10__20__slave ( .q(_RegFile_10__20), .qb(n1898), .d(
        _RegFile_reg_10__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_10__21__master ( .q(_RegFile_reg_10__21__m2s), .d(
        n3402), .sdi(n1898), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n957), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_10__21__slave ( .q(_RegFile_10__21), .qb(n1899), .d(
        _RegFile_reg_10__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n957), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_10__22__master ( .q(_RegFile_reg_10__22__m2s), .d(
        n3403), .sdi(n1899), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_10__22__slave ( .q(_RegFile_10__22), .qb(n1900), .d(
        _RegFile_reg_10__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_10__23__master ( .q(_RegFile_reg_10__23__m2s), .d(
        n3404), .sdi(n1900), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n957), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_10__23__slave ( .q(_RegFile_10__23), .qb(n1901), .d(
        _RegFile_reg_10__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n957), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_10__24__master ( .q(_RegFile_reg_10__24__m2s), .d(
        n3405), .sdi(n1901), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_10__24__slave ( .q(_RegFile_10__24), .qb(n1902), .d(
        _RegFile_reg_10__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_10__25__master ( .q(_RegFile_reg_10__25__m2s), .d(
        n3406), .sdi(n1902), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n957), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_10__25__slave ( .q(_RegFile_10__25), .qb(n1903), .d(
        _RegFile_reg_10__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n957), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_10__26__master ( .q(_RegFile_reg_10__26__m2s), .d(
        n3407), .sdi(n1903), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_10__26__slave ( .q(_RegFile_10__26), .qb(n1904), .d(
        _RegFile_reg_10__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_10__27__master ( .q(_RegFile_reg_10__27__m2s), .d(
        n3408), .sdi(n1904), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n957), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_10__27__slave ( .q(_RegFile_10__27), .qb(n1905), .d(
        _RegFile_reg_10__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n957), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_10__28__master ( .q(_RegFile_reg_10__28__m2s), .d(
        n3409), .sdi(n1905), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n948), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_10__28__slave ( .q(_RegFile_10__28), .qb(n1906), .d(
        _RegFile_reg_10__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n948), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_10__29__master ( .q(_RegFile_reg_10__29__m2s), .d(
        n3410), .sdi(n1906), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n957), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_10__29__slave ( .q(_RegFile_10__29), .qb(n1907), .d(
        _RegFile_reg_10__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n957), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_10__2__master ( .q(_RegFile_reg_10__2__m2s), .d(
        n3383), .sdi(n4287), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n957), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_10__2__slave ( .q(_RegFile_10__2), .qb(n4286), .d(
        _RegFile_reg_10__2__m2s), .g(Ctrl__Regs_1__en2), .rb(n957), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_10__30__master ( .q(_RegFile_reg_10__30__m2s), .d(
        n3411), .sdi(n1907), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n957), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_10__30__slave ( .q(_RegFile_10__30), .qb(n1908), .d(
        _RegFile_reg_10__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n957), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_10__31__master ( .q(_RegFile_reg_10__31__m2s), .d(
        n3412), .sdi(n1908), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n948), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_10__31__slave ( .q(_RegFile_10__31), .qb(n1909), .d(
        _RegFile_reg_10__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n948), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_10__3__master ( .q(_RegFile_reg_10__3__m2s), .d(
        n3384), .sdi(n4286), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n948), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_10__3__slave ( .q(_RegFile_10__3), .qb(n4285), .d(
        _RegFile_reg_10__3__m2s), .g(Ctrl__Regs_1__en2), .rb(n948), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_10__4__master ( .q(_RegFile_reg_10__4__m2s), .d(
        n3385), .sdi(n4285), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n957), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_10__4__slave ( .q(_RegFile_10__4), .qb(n4284), .d(
        _RegFile_reg_10__4__m2s), .g(Ctrl__Regs_1__en2), .rb(n957), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_10__5__master ( .q(_RegFile_reg_10__5__m2s), .d(
        n3386), .sdi(n4284), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n948), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_10__5__slave ( .q(_RegFile_10__5), .qb(n4283), .d(
        _RegFile_reg_10__5__m2s), .g(Ctrl__Regs_1__en2), .rb(n948), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_10__6__master ( .q(_RegFile_reg_10__6__m2s), .d(
        n3387), .sdi(n4283), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n957), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_10__6__slave ( .q(_RegFile_10__6), .qb(n4282), .d(
        _RegFile_reg_10__6__m2s), .g(Ctrl__Regs_1__en2), .rb(n957), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_10__7__master ( .q(_RegFile_reg_10__7__m2s), .d(
        n3388), .sdi(n4282), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n948), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_10__7__slave ( .q(_RegFile_10__7), .qb(n4281), .d(
        _RegFile_reg_10__7__m2s), .g(Ctrl__Regs_1__en2), .rb(n948), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_10__8__master ( .q(_RegFile_reg_10__8__m2s), .d(
        n3389), .sdi(n4281), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n957), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_10__8__slave ( .q(_RegFile_10__8), .qb(n1910), .d(
        _RegFile_reg_10__8__m2s), .g(Ctrl__Regs_1__en2), .rb(n957), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_10__9__master ( .q(_RegFile_reg_10__9__m2s), .d(
        n3390), .sdi(n1910), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n948), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_10__9__slave ( .q(_RegFile_10__9), .qb(n1911), .d(
        _RegFile_reg_10__9__m2s), .g(Ctrl__Regs_1__en2), .rb(n948), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_11__0__master ( .q(_RegFile_reg_11__0__m2s), .d(
        n3349), .sdi(n1909), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n957), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_11__0__slave ( .q(_RegFile_11__0), .qb(n4280), .d(
        _RegFile_reg_11__0__m2s), .g(Ctrl__Regs_1__en2), .rb(n957), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_11__10__master ( .q(_RegFile_reg_11__10__m2s), .d(
        n3359), .sdi(n1935), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n957), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_11__10__slave ( .q(_RegFile_11__10), .qb(n1912), .d(
        _RegFile_reg_11__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n957), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_11__11__master ( .q(_RegFile_reg_11__11__m2s), .d(
        n3360), .sdi(n1912), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n948), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_11__11__slave ( .q(_RegFile_11__11), .qb(n1913), .d(
        _RegFile_reg_11__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n948), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_11__12__master ( .q(_RegFile_reg_11__12__m2s), .d(
        n3361), .sdi(n1913), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n958), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_11__12__slave ( .q(_RegFile_11__12), .qb(n1914), .d(
        _RegFile_reg_11__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n958), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_11__13__master ( .q(_RegFile_reg_11__13__m2s), .d(
        n3362), .sdi(n1914), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n948), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_11__13__slave ( .q(_RegFile_11__13), .qb(n1915), .d(
        _RegFile_reg_11__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n948), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_11__14__master ( .q(_RegFile_reg_11__14__m2s), .d(
        n3363), .sdi(n1915), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n958), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_11__14__slave ( .q(_RegFile_11__14), .qb(n1916), .d(
        _RegFile_reg_11__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n958), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_11__15__master ( .q(_RegFile_reg_11__15__m2s), .d(
        n3364), .sdi(n1916), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n948), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_11__15__slave ( .q(_RegFile_11__15), .qb(n1917), .d(
        _RegFile_reg_11__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n948), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_11__16__master ( .q(_RegFile_reg_11__16__m2s), .d(
        n3365), .sdi(n1917), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n958), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_11__16__slave ( .q(_RegFile_11__16), .qb(n1918), .d(
        _RegFile_reg_11__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n958), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_11__17__master ( .q(_RegFile_reg_11__17__m2s), .d(
        n3366), .sdi(n1918), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n948), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_11__17__slave ( .q(_RegFile_11__17), .qb(n1919), .d(
        _RegFile_reg_11__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n948), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_11__18__master ( .q(_RegFile_reg_11__18__m2s), .d(
        n3367), .sdi(n1919), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n958), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_11__18__slave ( .q(_RegFile_11__18), .qb(n1920), .d(
        _RegFile_reg_11__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n958), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_11__19__master ( .q(_RegFile_reg_11__19__m2s), .d(
        n3368), .sdi(n1920), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n948), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_11__19__slave ( .q(_RegFile_11__19), .qb(n1921), .d(
        _RegFile_reg_11__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n948), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_11__1__master ( .q(_RegFile_reg_11__1__m2s), .d(
        n3350), .sdi(n4280), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n948), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_11__1__slave ( .q(_RegFile_11__1), .qb(n4279), .d(
        _RegFile_reg_11__1__m2s), .g(Ctrl__Regs_1__en2), .rb(n948), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_11__20__master ( .q(_RegFile_reg_11__20__m2s), .d(
        n3369), .sdi(n1921), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n948), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_11__20__slave ( .q(_RegFile_11__20), .qb(n1922), .d(
        _RegFile_reg_11__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n948), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_11__21__master ( .q(_RegFile_reg_11__21__m2s), .d(
        n3370), .sdi(n1922), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n958), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_11__21__slave ( .q(_RegFile_11__21), .qb(n1923), .d(
        _RegFile_reg_11__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n958), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_11__22__master ( .q(_RegFile_reg_11__22__m2s), .d(
        n3371), .sdi(n1923), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n948), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_11__22__slave ( .q(_RegFile_11__22), .qb(n1924), .d(
        _RegFile_reg_11__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n948), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_11__23__master ( .q(_RegFile_reg_11__23__m2s), .d(
        n3372), .sdi(n1924), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n958), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_11__23__slave ( .q(_RegFile_11__23), .qb(n1925), .d(
        _RegFile_reg_11__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n958), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_11__24__master ( .q(_RegFile_reg_11__24__m2s), .d(
        n3373), .sdi(n1925), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n948), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_11__24__slave ( .q(_RegFile_11__24), .qb(n1926), .d(
        _RegFile_reg_11__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n948), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_11__25__master ( .q(_RegFile_reg_11__25__m2s), .d(
        n3374), .sdi(n1926), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n958), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_11__25__slave ( .q(_RegFile_11__25), .qb(n1927), .d(
        _RegFile_reg_11__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n958), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_11__26__master ( .q(_RegFile_reg_11__26__m2s), .d(
        n3375), .sdi(n1927), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_11__26__slave ( .q(_RegFile_11__26), .qb(n1928), .d(
        _RegFile_reg_11__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_11__27__master ( .q(_RegFile_reg_11__27__m2s), .d(
        n3376), .sdi(n1928), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n958), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_11__27__slave ( .q(_RegFile_11__27), .qb(n1929), .d(
        _RegFile_reg_11__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n958), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_11__28__master ( .q(_RegFile_reg_11__28__m2s), .d(
        n3377), .sdi(n1929), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_11__28__slave ( .q(_RegFile_11__28), .qb(n1930), .d(
        _RegFile_reg_11__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_11__29__master ( .q(_RegFile_reg_11__29__m2s), .d(
        n3378), .sdi(n1930), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n958), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_11__29__slave ( .q(_RegFile_11__29), .qb(n1931), .d(
        _RegFile_reg_11__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n958), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_11__2__master ( .q(_RegFile_reg_11__2__m2s), .d(
        n3351), .sdi(n4279), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n958), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_11__2__slave ( .q(_RegFile_11__2), .qb(n4278), .d(
        _RegFile_reg_11__2__m2s), .g(Ctrl__Regs_1__en2), .rb(n958), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_11__30__master ( .q(_RegFile_reg_11__30__m2s), .d(
        n3379), .sdi(n1931), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n958), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_11__30__slave ( .q(_RegFile_11__30), .qb(n1932), .d(
        _RegFile_reg_11__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n958), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_11__31__master ( .q(_RegFile_reg_11__31__m2s), .d(
        n3380), .sdi(n1932), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_11__31__slave ( .q(_RegFile_11__31), .qb(n1933), .d(
        _RegFile_reg_11__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_11__3__master ( .q(_RegFile_reg_11__3__m2s), .d(
        n3352), .sdi(n4278), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_11__3__slave ( .q(_RegFile_11__3), .qb(n4277), .d(
        _RegFile_reg_11__3__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_11__4__master ( .q(_RegFile_reg_11__4__m2s), .d(
        n3353), .sdi(n4277), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n958), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_11__4__slave ( .q(_RegFile_11__4), .qb(n4276), .d(
        _RegFile_reg_11__4__m2s), .g(Ctrl__Regs_1__en2), .rb(n958), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_11__5__master ( .q(_RegFile_reg_11__5__m2s), .d(
        n3354), .sdi(n4276), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_11__5__slave ( .q(_RegFile_11__5), .qb(n4275), .d(
        _RegFile_reg_11__5__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_11__6__master ( .q(_RegFile_reg_11__6__m2s), .d(
        n3355), .sdi(n4275), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n958), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_11__6__slave ( .q(_RegFile_11__6), .qb(n4274), .d(
        _RegFile_reg_11__6__m2s), .g(Ctrl__Regs_1__en2), .rb(n958), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_11__7__master ( .q(_RegFile_reg_11__7__m2s), .d(
        n3356), .sdi(n4274), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_11__7__slave ( .q(_RegFile_11__7), .qb(n4273), .d(
        _RegFile_reg_11__7__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_11__8__master ( .q(_RegFile_reg_11__8__m2s), .d(
        n3357), .sdi(n4273), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n958), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_11__8__slave ( .q(_RegFile_11__8), .qb(n1934), .d(
        _RegFile_reg_11__8__m2s), .g(Ctrl__Regs_1__en2), .rb(n958), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_11__9__master ( .q(_RegFile_reg_11__9__m2s), .d(
        n3358), .sdi(n1934), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_11__9__slave ( .q(_RegFile_11__9), .qb(n1935), .d(
        _RegFile_reg_11__9__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_12__0__master ( .q(_RegFile_reg_12__0__m2s), .d(
        n3317), .sdi(n1933), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n958), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_12__0__slave ( .q(_RegFile_12__0), .qb(n4272), .d(
        _RegFile_reg_12__0__m2s), .g(Ctrl__Regs_1__en2), .rb(n958), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_12__10__master ( .q(_RegFile_reg_12__10__m2s), .d(
        n3327), .sdi(n1959), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n959), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_12__10__slave ( .q(_RegFile_12__10), .qb(n1936), .d(
        _RegFile_reg_12__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n959), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_12__11__master ( .q(_RegFile_reg_12__11__m2s), .d(
        n3328), .sdi(n1936), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_12__11__slave ( .q(_RegFile_12__11), .qb(n1937), .d(
        _RegFile_reg_12__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_12__12__master ( .q(_RegFile_reg_12__12__m2s), .d(
        n3329), .sdi(n1937), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n959), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_12__12__slave ( .q(_RegFile_12__12), .qb(n1938), .d(
        _RegFile_reg_12__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n959), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_12__13__master ( .q(_RegFile_reg_12__13__m2s), .d(
        n3330), .sdi(n1938), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_12__13__slave ( .q(_RegFile_12__13), .qb(n1939), .d(
        _RegFile_reg_12__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_12__14__master ( .q(_RegFile_reg_12__14__m2s), .d(
        n3331), .sdi(n1939), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n959), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_12__14__slave ( .q(_RegFile_12__14), .qb(n1940), .d(
        _RegFile_reg_12__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n959), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_12__15__master ( .q(_RegFile_reg_12__15__m2s), .d(
        n3332), .sdi(n1940), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_12__15__slave ( .q(_RegFile_12__15), .qb(n1941), .d(
        _RegFile_reg_12__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_12__16__master ( .q(_RegFile_reg_12__16__m2s), .d(
        n3333), .sdi(n1941), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n959), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_12__16__slave ( .q(_RegFile_12__16), .qb(n1942), .d(
        _RegFile_reg_12__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n959), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_12__17__master ( .q(_RegFile_reg_12__17__m2s), .d(
        n3334), .sdi(n1942), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_12__17__slave ( .q(_RegFile_12__17), .qb(n1943), .d(
        _RegFile_reg_12__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_12__18__master ( .q(_RegFile_reg_12__18__m2s), .d(
        n3335), .sdi(n1943), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n959), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_12__18__slave ( .q(_RegFile_12__18), .qb(n1944), .d(
        _RegFile_reg_12__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n959), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_12__19__master ( .q(_RegFile_reg_12__19__m2s), .d(
        n3336), .sdi(n1944), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_12__19__slave ( .q(_RegFile_12__19), .qb(n1945), .d(
        _RegFile_reg_12__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_12__1__master ( .q(_RegFile_reg_12__1__m2s), .d(
        n3318), .sdi(n4272), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_12__1__slave ( .q(_RegFile_12__1), .qb(n4271), .d(
        _RegFile_reg_12__1__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_12__20__master ( .q(_RegFile_reg_12__20__m2s), .d(
        n3337), .sdi(n1945), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_12__20__slave ( .q(_RegFile_12__20), .qb(n1946), .d(
        _RegFile_reg_12__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_12__21__master ( .q(_RegFile_reg_12__21__m2s), .d(
        n3338), .sdi(n1946), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n959), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_12__21__slave ( .q(_RegFile_12__21), .qb(n1947), .d(
        _RegFile_reg_12__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n959), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_12__22__master ( .q(_RegFile_reg_12__22__m2s), .d(
        n3339), .sdi(n1947), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_12__22__slave ( .q(_RegFile_12__22), .qb(n1948), .d(
        _RegFile_reg_12__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_12__23__master ( .q(_RegFile_reg_12__23__m2s), .d(
        n3340), .sdi(n1948), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n959), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_12__23__slave ( .q(_RegFile_12__23), .qb(n1949), .d(
        _RegFile_reg_12__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n959), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_12__24__master ( .q(_RegFile_reg_12__24__m2s), .d(
        n3341), .sdi(n1949), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n946), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_12__24__slave ( .q(_RegFile_12__24), .qb(n1950), .d(
        _RegFile_reg_12__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n946), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_12__25__master ( .q(_RegFile_reg_12__25__m2s), .d(
        n3342), .sdi(n1950), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n959), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_12__25__slave ( .q(_RegFile_12__25), .qb(n1951), .d(
        _RegFile_reg_12__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n959), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_12__26__master ( .q(_RegFile_reg_12__26__m2s), .d(
        n3343), .sdi(n1951), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n946), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_12__26__slave ( .q(_RegFile_12__26), .qb(n1952), .d(
        _RegFile_reg_12__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n946), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_12__27__master ( .q(_RegFile_reg_12__27__m2s), .d(
        n3344), .sdi(n1952), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n959), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_12__27__slave ( .q(_RegFile_12__27), .qb(n1953), .d(
        _RegFile_reg_12__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n959), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_12__28__master ( .q(_RegFile_reg_12__28__m2s), .d(
        n3345), .sdi(n1953), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n946), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_12__28__slave ( .q(_RegFile_12__28), .qb(n1954), .d(
        _RegFile_reg_12__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n946), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_12__29__master ( .q(_RegFile_reg_12__29__m2s), .d(
        n3346), .sdi(n1954), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n959), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_12__29__slave ( .q(_RegFile_12__29), .qb(n1955), .d(
        _RegFile_reg_12__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n959), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_12__2__master ( .q(_RegFile_reg_12__2__m2s), .d(
        n3319), .sdi(n4271), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n959), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_12__2__slave ( .q(_RegFile_12__2), .qb(n4270), .d(
        _RegFile_reg_12__2__m2s), .g(Ctrl__Regs_1__en2), .rb(n959), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_12__30__master ( .q(_RegFile_reg_12__30__m2s), .d(
        n3347), .sdi(n1955), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n959), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_12__30__slave ( .q(_RegFile_12__30), .qb(n1956), .d(
        _RegFile_reg_12__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n959), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_12__31__master ( .q(_RegFile_reg_12__31__m2s), .d(
        n3348), .sdi(n1956), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n946), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_12__31__slave ( .q(_RegFile_12__31), .qb(n1957), .d(
        _RegFile_reg_12__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n946), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_12__3__master ( .q(_RegFile_reg_12__3__m2s), .d(
        n3320), .sdi(n4270), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n946), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_12__3__slave ( .q(_RegFile_12__3), .qb(n4269), .d(
        _RegFile_reg_12__3__m2s), .g(Ctrl__Regs_1__en2), .rb(n946), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_12__4__master ( .q(_RegFile_reg_12__4__m2s), .d(
        n3321), .sdi(n4269), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n959), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_12__4__slave ( .q(_RegFile_12__4), .qb(n4268), .d(
        _RegFile_reg_12__4__m2s), .g(Ctrl__Regs_1__en2), .rb(n959), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_12__5__master ( .q(_RegFile_reg_12__5__m2s), .d(
        n3322), .sdi(n4268), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n946), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_12__5__slave ( .q(_RegFile_12__5), .qb(n4267), .d(
        _RegFile_reg_12__5__m2s), .g(Ctrl__Regs_1__en2), .rb(n946), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_12__6__master ( .q(_RegFile_reg_12__6__m2s), .d(
        n3323), .sdi(n4267), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n959), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_12__6__slave ( .q(_RegFile_12__6), .qb(n4266), .d(
        _RegFile_reg_12__6__m2s), .g(Ctrl__Regs_1__en2), .rb(n959), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_12__7__master ( .q(_RegFile_reg_12__7__m2s), .d(
        n3324), .sdi(n4266), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n946), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_12__7__slave ( .q(_RegFile_12__7), .qb(n4265), .d(
        _RegFile_reg_12__7__m2s), .g(Ctrl__Regs_1__en2), .rb(n946), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_12__8__master ( .q(_RegFile_reg_12__8__m2s), .d(
        n3325), .sdi(n4265), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n959), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_12__8__slave ( .q(_RegFile_12__8), .qb(n1958), .d(
        _RegFile_reg_12__8__m2s), .g(Ctrl__Regs_1__en2), .rb(n959), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_12__9__master ( .q(_RegFile_reg_12__9__m2s), .d(
        n3326), .sdi(n1958), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n946), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_12__9__slave ( .q(_RegFile_12__9), .qb(n1959), .d(
        _RegFile_reg_12__9__m2s), .g(Ctrl__Regs_1__en2), .rb(n946), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_13__0__master ( .q(_RegFile_reg_13__0__m2s), .d(
        n3285), .sdi(n1957), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_13__0__slave ( .q(_RegFile_13__0), .qb(n4264), .d(
        _RegFile_reg_13__0__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_13__10__master ( .q(_RegFile_reg_13__10__m2s), .d(
        n3295), .sdi(n1983), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_13__10__slave ( .q(_RegFile_13__10), .qb(n1960), .d(
        _RegFile_reg_13__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_13__11__master ( .q(_RegFile_reg_13__11__m2s), .d(
        n3296), .sdi(n1960), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n946), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_13__11__slave ( .q(_RegFile_13__11), .qb(n1961), .d(
        _RegFile_reg_13__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n946), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_13__12__master ( .q(_RegFile_reg_13__12__m2s), .d(
        n3297), .sdi(n1961), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_13__12__slave ( .q(_RegFile_13__12), .qb(n1962), .d(
        _RegFile_reg_13__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_13__13__master ( .q(_RegFile_reg_13__13__m2s), .d(
        n3298), .sdi(n1962), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n946), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_13__13__slave ( .q(_RegFile_13__13), .qb(n1963), .d(
        _RegFile_reg_13__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n946), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_13__14__master ( .q(_RegFile_reg_13__14__m2s), .d(
        n3299), .sdi(n1963), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_13__14__slave ( .q(_RegFile_13__14), .qb(n1964), .d(
        _RegFile_reg_13__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_13__15__master ( .q(_RegFile_reg_13__15__m2s), .d(
        n3300), .sdi(n1964), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n946), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_13__15__slave ( .q(_RegFile_13__15), .qb(n1965), .d(
        _RegFile_reg_13__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n946), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_13__16__master ( .q(_RegFile_reg_13__16__m2s), .d(
        n3301), .sdi(n1965), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_13__16__slave ( .q(_RegFile_13__16), .qb(n1966), .d(
        _RegFile_reg_13__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_13__17__master ( .q(_RegFile_reg_13__17__m2s), .d(
        n3302), .sdi(n1966), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n946), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_13__17__slave ( .q(_RegFile_13__17), .qb(n1967), .d(
        _RegFile_reg_13__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n946), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_13__18__master ( .q(_RegFile_reg_13__18__m2s), .d(
        n3303), .sdi(n1967), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_13__18__slave ( .q(_RegFile_13__18), .qb(n1968), .d(
        _RegFile_reg_13__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_13__19__master ( .q(_RegFile_reg_13__19__m2s), .d(
        n3304), .sdi(n1968), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n946), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_13__19__slave ( .q(_RegFile_13__19), .qb(n1969), .d(
        _RegFile_reg_13__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n946), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_13__1__master ( .q(_RegFile_reg_13__1__m2s), .d(
        n3286), .sdi(n4264), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n946), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_13__1__slave ( .q(_RegFile_13__1), .qb(n4263), .d(
        _RegFile_reg_13__1__m2s), .g(Ctrl__Regs_1__en2), .rb(n946), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_13__20__master ( .q(_RegFile_reg_13__20__m2s), .d(
        n3305), .sdi(n1969), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n946), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_13__20__slave ( .q(_RegFile_13__20), .qb(n1970), .d(
        _RegFile_reg_13__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n946), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_13__21__master ( .q(_RegFile_reg_13__21__m2s), .d(
        n3306), .sdi(n1970), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_13__21__slave ( .q(_RegFile_13__21), .qb(n1971), .d(
        _RegFile_reg_13__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_13__22__master ( .q(_RegFile_reg_13__22__m2s), .d(
        n3307), .sdi(n1971), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n945), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_13__22__slave ( .q(_RegFile_13__22), .qb(n1972), .d(
        _RegFile_reg_13__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n945), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_13__23__master ( .q(_RegFile_reg_13__23__m2s), .d(
        n3308), .sdi(n1972), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_13__23__slave ( .q(_RegFile_13__23), .qb(n1973), .d(
        _RegFile_reg_13__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_13__24__master ( .q(_RegFile_reg_13__24__m2s), .d(
        n3309), .sdi(n1973), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n945), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_13__24__slave ( .q(_RegFile_13__24), .qb(n1974), .d(
        _RegFile_reg_13__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n945), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_13__25__master ( .q(_RegFile_reg_13__25__m2s), .d(
        n3310), .sdi(n1974), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_13__25__slave ( .q(_RegFile_13__25), .qb(n1975), .d(
        _RegFile_reg_13__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_13__26__master ( .q(_RegFile_reg_13__26__m2s), .d(
        n3311), .sdi(n1975), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n945), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_13__26__slave ( .q(_RegFile_13__26), .qb(n1976), .d(
        _RegFile_reg_13__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n945), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_13__27__master ( .q(_RegFile_reg_13__27__m2s), .d(
        n3312), .sdi(n1976), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_13__27__slave ( .q(_RegFile_13__27), .qb(n1977), .d(
        _RegFile_reg_13__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_13__28__master ( .q(_RegFile_reg_13__28__m2s), .d(
        n3313), .sdi(n1977), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n945), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_13__28__slave ( .q(_RegFile_13__28), .qb(n1978), .d(
        _RegFile_reg_13__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n945), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_13__29__master ( .q(_RegFile_reg_13__29__m2s), .d(
        n3314), .sdi(n1978), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_13__29__slave ( .q(_RegFile_13__29), .qb(n1979), .d(
        _RegFile_reg_13__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_13__2__master ( .q(_RegFile_reg_13__2__m2s), .d(
        n3287), .sdi(n4263), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_13__2__slave ( .q(_RegFile_13__2), .qb(n4262), .d(
        _RegFile_reg_13__2__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_13__30__master ( .q(_RegFile_reg_13__30__m2s), .d(
        n3315), .sdi(n1979), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_13__30__slave ( .q(_RegFile_13__30), .qb(n1980), .d(
        _RegFile_reg_13__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_13__31__master ( .q(_RegFile_reg_13__31__m2s), .d(
        n3316), .sdi(n1980), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n945), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_13__31__slave ( .q(_RegFile_13__31), .qb(n1981), .d(
        _RegFile_reg_13__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n945), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_13__3__master ( .q(_RegFile_reg_13__3__m2s), .d(
        n3288), .sdi(n4262), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n945), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_13__3__slave ( .q(_RegFile_13__3), .qb(n4261), .d(
        _RegFile_reg_13__3__m2s), .g(Ctrl__Regs_1__en2), .rb(n945), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_13__4__master ( .q(_RegFile_reg_13__4__m2s), .d(
        n3289), .sdi(n4261), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_13__4__slave ( .q(_RegFile_13__4), .qb(n4260), .d(
        _RegFile_reg_13__4__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_13__5__master ( .q(_RegFile_reg_13__5__m2s), .d(
        n3290), .sdi(n4260), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n945), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_13__5__slave ( .q(_RegFile_13__5), .qb(n4259), .d(
        _RegFile_reg_13__5__m2s), .g(Ctrl__Regs_1__en2), .rb(n945), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_13__6__master ( .q(_RegFile_reg_13__6__m2s), .d(
        n3291), .sdi(n4259), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_13__6__slave ( .q(_RegFile_13__6), .qb(n4258), .d(
        _RegFile_reg_13__6__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_13__7__master ( .q(_RegFile_reg_13__7__m2s), .d(
        n3292), .sdi(n4258), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n945), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_13__7__slave ( .q(_RegFile_13__7), .qb(n4257), .d(
        _RegFile_reg_13__7__m2s), .g(Ctrl__Regs_1__en2), .rb(n945), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_13__8__master ( .q(_RegFile_reg_13__8__m2s), .d(
        n3293), .sdi(n4257), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_13__8__slave ( .q(_RegFile_13__8), .qb(n1982), .d(
        _RegFile_reg_13__8__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_13__9__master ( .q(_RegFile_reg_13__9__m2s), .d(
        n3294), .sdi(n1982), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n945), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_13__9__slave ( .q(_RegFile_13__9), .qb(n1983), .d(
        _RegFile_reg_13__9__m2s), .g(Ctrl__Regs_1__en2), .rb(n945), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_14__0__master ( .q(_RegFile_reg_14__0__m2s), .d(
        n3253), .sdi(n1981), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_14__0__slave ( .q(_RegFile_14__0), .qb(n4256), .d(
        _RegFile_reg_14__0__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_14__10__master ( .q(_RegFile_reg_14__10__m2s), .d(
        n3263), .sdi(n2007), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_14__10__slave ( .q(_RegFile_14__10), .qb(n1984), .d(
        _RegFile_reg_14__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_14__11__master ( .q(_RegFile_reg_14__11__m2s), .d(
        n3264), .sdi(n1984), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n945), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_14__11__slave ( .q(_RegFile_14__11), .qb(n1985), .d(
        _RegFile_reg_14__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n945), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_14__12__master ( .q(_RegFile_reg_14__12__m2s), .d(
        n3265), .sdi(n1985), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_14__12__slave ( .q(_RegFile_14__12), .qb(n1986), .d(
        _RegFile_reg_14__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_14__13__master ( .q(_RegFile_reg_14__13__m2s), .d(
        n3266), .sdi(n1986), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n945), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_14__13__slave ( .q(_RegFile_14__13), .qb(n1987), .d(
        _RegFile_reg_14__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n945), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_14__14__master ( .q(_RegFile_reg_14__14__m2s), .d(
        n3267), .sdi(n1987), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_14__14__slave ( .q(_RegFile_14__14), .qb(n1988), .d(
        _RegFile_reg_14__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_14__15__master ( .q(_RegFile_reg_14__15__m2s), .d(
        n3268), .sdi(n1988), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n945), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_14__15__slave ( .q(_RegFile_14__15), .qb(n1989), .d(
        _RegFile_reg_14__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n945), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_14__16__master ( .q(_RegFile_reg_14__16__m2s), .d(
        n3269), .sdi(n1989), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_14__16__slave ( .q(_RegFile_14__16), .qb(n1990), .d(
        _RegFile_reg_14__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_14__17__master ( .q(_RegFile_reg_14__17__m2s), .d(
        n3270), .sdi(n1990), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n945), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_14__17__slave ( .q(_RegFile_14__17), .qb(n1991), .d(
        _RegFile_reg_14__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n945), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_14__18__master ( .q(_RegFile_reg_14__18__m2s), .d(
        n3271), .sdi(n1991), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_14__18__slave ( .q(_RegFile_14__18), .qb(n1992), .d(
        _RegFile_reg_14__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_14__19__master ( .q(_RegFile_reg_14__19__m2s), .d(
        n3272), .sdi(n1992), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n945), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_14__19__slave ( .q(_RegFile_14__19), .qb(n1993), .d(
        _RegFile_reg_14__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n945), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_14__1__master ( .q(_RegFile_reg_14__1__m2s), .d(
        n3254), .sdi(n4256), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n945), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_14__1__slave ( .q(_RegFile_14__1), .qb(n4255), .d(
        _RegFile_reg_14__1__m2s), .g(Ctrl__Regs_1__en2), .rb(n945), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_14__20__master ( .q(_RegFile_reg_14__20__m2s), .d(
        n3273), .sdi(n1993), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_14__20__slave ( .q(_RegFile_14__20), .qb(n1994), .d(
        _RegFile_reg_14__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_14__21__master ( .q(_RegFile_reg_14__21__m2s), .d(
        n3274), .sdi(n1994), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_14__21__slave ( .q(_RegFile_14__21), .qb(n1995), .d(
        _RegFile_reg_14__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_14__22__master ( .q(_RegFile_reg_14__22__m2s), .d(
        n3275), .sdi(n1995), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_14__22__slave ( .q(_RegFile_14__22), .qb(n1996), .d(
        _RegFile_reg_14__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_14__23__master ( .q(_RegFile_reg_14__23__m2s), .d(
        n3276), .sdi(n1996), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_14__23__slave ( .q(_RegFile_14__23), .qb(n1997), .d(
        _RegFile_reg_14__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_14__24__master ( .q(_RegFile_reg_14__24__m2s), .d(
        n3277), .sdi(n1997), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_14__24__slave ( .q(_RegFile_14__24), .qb(n1998), .d(
        _RegFile_reg_14__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_14__25__master ( .q(_RegFile_reg_14__25__m2s), .d(
        n3278), .sdi(n1998), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_14__25__slave ( .q(_RegFile_14__25), .qb(n1999), .d(
        _RegFile_reg_14__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_14__26__master ( .q(_RegFile_reg_14__26__m2s), .d(
        n3279), .sdi(n1999), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_14__26__slave ( .q(_RegFile_14__26), .qb(n2000), .d(
        _RegFile_reg_14__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_14__27__master ( .q(_RegFile_reg_14__27__m2s), .d(
        n3280), .sdi(n2000), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_14__27__slave ( .q(_RegFile_14__27), .qb(n2001), .d(
        _RegFile_reg_14__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_14__28__master ( .q(_RegFile_reg_14__28__m2s), .d(
        n3281), .sdi(n2001), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_14__28__slave ( .q(_RegFile_14__28), .qb(n2002), .d(
        _RegFile_reg_14__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_14__29__master ( .q(_RegFile_reg_14__29__m2s), .d(
        n3282), .sdi(n2002), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_14__29__slave ( .q(_RegFile_14__29), .qb(n2003), .d(
        _RegFile_reg_14__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_14__2__master ( .q(_RegFile_reg_14__2__m2s), .d(
        n3255), .sdi(n4255), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_14__2__slave ( .q(_RegFile_14__2), .qb(n4254), .d(
        _RegFile_reg_14__2__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_14__30__master ( .q(_RegFile_reg_14__30__m2s), .d(
        n3283), .sdi(n2003), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_14__30__slave ( .q(_RegFile_14__30), .qb(n2004), .d(
        _RegFile_reg_14__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_14__31__master ( .q(_RegFile_reg_14__31__m2s), .d(
        n3284), .sdi(n2004), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_14__31__slave ( .q(_RegFile_14__31), .qb(n2005), .d(
        _RegFile_reg_14__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_14__3__master ( .q(_RegFile_reg_14__3__m2s), .d(
        n3256), .sdi(n4254), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_14__3__slave ( .q(_RegFile_14__3), .qb(n4253), .d(
        _RegFile_reg_14__3__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_14__4__master ( .q(_RegFile_reg_14__4__m2s), .d(
        n3257), .sdi(n4253), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_14__4__slave ( .q(_RegFile_14__4), .qb(n4252), .d(
        _RegFile_reg_14__4__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_14__5__master ( .q(_RegFile_reg_14__5__m2s), .d(
        n3258), .sdi(n4252), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_14__5__slave ( .q(_RegFile_14__5), .qb(n4251), .d(
        _RegFile_reg_14__5__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_14__6__master ( .q(_RegFile_reg_14__6__m2s), .d(
        n3259), .sdi(n4251), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_14__6__slave ( .q(_RegFile_14__6), .qb(n4250), .d(
        _RegFile_reg_14__6__m2s), .g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_14__7__master ( .q(_RegFile_reg_14__7__m2s), .d(
        n3260), .sdi(n4250), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_14__7__slave ( .q(_RegFile_14__7), .qb(n4249), .d(
        _RegFile_reg_14__7__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_14__8__master ( .q(_RegFile_reg_14__8__m2s), .d(
        n3261), .sdi(n4249), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_14__8__slave ( .q(_RegFile_14__8), .qb(n2006), .d(
        _RegFile_reg_14__8__m2s), .g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_14__9__master ( .q(_RegFile_reg_14__9__m2s), .d(
        n3262), .sdi(n2006), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_14__9__slave ( .q(_RegFile_14__9), .qb(n2007), .d(
        _RegFile_reg_14__9__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_15__0__master ( .q(_RegFile_reg_15__0__m2s), .d(
        n3221), .sdi(n2005), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_15__0__slave ( .q(_RegFile_15__0), .qb(n4248), .d(
        _RegFile_reg_15__0__m2s), .g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_15__10__master ( .q(_RegFile_reg_15__10__m2s), .d(
        n3231), .sdi(n2031), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_15__10__slave ( .q(_RegFile_15__10), .qb(n2008), .d(
        _RegFile_reg_15__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_15__11__master ( .q(_RegFile_reg_15__11__m2s), .d(
        n3232), .sdi(n2008), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_15__11__slave ( .q(_RegFile_15__11), .qb(n2009), .d(
        _RegFile_reg_15__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_15__12__master ( .q(_RegFile_reg_15__12__m2s), .d(
        n3233), .sdi(n2009), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_15__12__slave ( .q(_RegFile_15__12), .qb(n2010), .d(
        _RegFile_reg_15__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_15__13__master ( .q(_RegFile_reg_15__13__m2s), .d(
        n3234), .sdi(n2010), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_15__13__slave ( .q(_RegFile_15__13), .qb(n2011), .d(
        _RegFile_reg_15__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_15__14__master ( .q(_RegFile_reg_15__14__m2s), .d(
        n3235), .sdi(n2011), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_15__14__slave ( .q(_RegFile_15__14), .qb(n2012), .d(
        _RegFile_reg_15__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_15__15__master ( .q(_RegFile_reg_15__15__m2s), .d(
        n3236), .sdi(n2012), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_15__15__slave ( .q(_RegFile_15__15), .qb(n2013), .d(
        _RegFile_reg_15__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_15__16__master ( .q(_RegFile_reg_15__16__m2s), .d(
        n3237), .sdi(n2013), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_15__16__slave ( .q(_RegFile_15__16), .qb(n2014), .d(
        _RegFile_reg_15__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_15__17__master ( .q(_RegFile_reg_15__17__m2s), .d(
        n3238), .sdi(n2014), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_15__17__slave ( .q(_RegFile_15__17), .qb(n2015), .d(
        _RegFile_reg_15__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_15__18__master ( .q(_RegFile_reg_15__18__m2s), .d(
        n3239), .sdi(n2015), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_15__18__slave ( .q(_RegFile_15__18), .qb(n2016), .d(
        _RegFile_reg_15__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_15__19__master ( .q(_RegFile_reg_15__19__m2s), .d(
        n3240), .sdi(n2016), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n944), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_15__19__slave ( .q(_RegFile_15__19), .qb(n2017), .d(
        _RegFile_reg_15__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n944), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_15__1__master ( .q(_RegFile_reg_15__1__m2s), .d(
        n3222), .sdi(n4248), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_15__1__slave ( .q(_RegFile_15__1), .qb(n4247), .d(
        _RegFile_reg_15__1__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_15__20__master ( .q(_RegFile_reg_15__20__m2s), .d(
        n3241), .sdi(n2017), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n944), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_15__20__slave ( .q(_RegFile_15__20), .qb(n2018), .d(
        _RegFile_reg_15__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n944), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_15__21__master ( .q(_RegFile_reg_15__21__m2s), .d(
        n3242), .sdi(n2018), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_15__21__slave ( .q(_RegFile_15__21), .qb(n2019), .d(
        _RegFile_reg_15__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_15__22__master ( .q(_RegFile_reg_15__22__m2s), .d(
        n3243), .sdi(n2019), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n944), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_15__22__slave ( .q(_RegFile_15__22), .qb(n2020), .d(
        _RegFile_reg_15__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n944), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_15__23__master ( .q(_RegFile_reg_15__23__m2s), .d(
        n3244), .sdi(n2020), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_15__23__slave ( .q(_RegFile_15__23), .qb(n2021), .d(
        _RegFile_reg_15__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_15__24__master ( .q(_RegFile_reg_15__24__m2s), .d(
        n3245), .sdi(n2021), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n944), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_15__24__slave ( .q(_RegFile_15__24), .qb(n2022), .d(
        _RegFile_reg_15__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n944), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_15__25__master ( .q(_RegFile_reg_15__25__m2s), .d(
        n3246), .sdi(n2022), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_15__25__slave ( .q(_RegFile_15__25), .qb(n2023), .d(
        _RegFile_reg_15__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_15__26__master ( .q(_RegFile_reg_15__26__m2s), .d(
        n3247), .sdi(n2023), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n944), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_15__26__slave ( .q(_RegFile_15__26), .qb(n2024), .d(
        _RegFile_reg_15__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n944), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_15__27__master ( .q(_RegFile_reg_15__27__m2s), .d(
        n3248), .sdi(n2024), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_15__27__slave ( .q(_RegFile_15__27), .qb(n2025), .d(
        _RegFile_reg_15__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_15__28__master ( .q(_RegFile_reg_15__28__m2s), .d(
        n3249), .sdi(n2025), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n944), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_15__28__slave ( .q(_RegFile_15__28), .qb(n2026), .d(
        _RegFile_reg_15__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n944), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_15__29__master ( .q(_RegFile_reg_15__29__m2s), .d(
        n3250), .sdi(n2026), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_15__29__slave ( .q(_RegFile_15__29), .qb(n2027), .d(
        _RegFile_reg_15__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_15__2__master ( .q(_RegFile_reg_15__2__m2s), .d(
        n3223), .sdi(n4247), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_15__2__slave ( .q(_RegFile_15__2), .qb(n4246), .d(
        _RegFile_reg_15__2__m2s), .g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_15__30__master ( .q(_RegFile_reg_15__30__m2s), .d(
        n3251), .sdi(n2027), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_15__30__slave ( .q(_RegFile_15__30), .qb(n2028), .d(
        _RegFile_reg_15__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_15__31__master ( .q(_RegFile_reg_15__31__m2s), .d(
        n3252), .sdi(n2028), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n944), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_15__31__slave ( .q(_RegFile_15__31), .qb(n2029), .d(
        _RegFile_reg_15__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n944), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_15__3__master ( .q(_RegFile_reg_15__3__m2s), .d(
        n3224), .sdi(n4246), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n944), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_15__3__slave ( .q(_RegFile_15__3), .qb(n4245), .d(
        _RegFile_reg_15__3__m2s), .g(Ctrl__Regs_1__en2), .rb(n944), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_15__4__master ( .q(_RegFile_reg_15__4__m2s), .d(
        n3225), .sdi(n4245), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n960), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_15__4__slave ( .q(_RegFile_15__4), .qb(n4244), .d(
        _RegFile_reg_15__4__m2s), .g(Ctrl__Regs_1__en2), .rb(n960), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_15__5__master ( .q(_RegFile_reg_15__5__m2s), .d(
        n3226), .sdi(n4244), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n944), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_15__5__slave ( .q(_RegFile_15__5), .qb(n4243), .d(
        _RegFile_reg_15__5__m2s), .g(Ctrl__Regs_1__en2), .rb(n944), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_15__6__master ( .q(_RegFile_reg_15__6__m2s), .d(
        n3227), .sdi(n4243), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n960), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_15__6__slave ( .q(_RegFile_15__6), .qb(n4242), .d(
        _RegFile_reg_15__6__m2s), .g(Ctrl__Regs_1__en2), .rb(n960), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_15__7__master ( .q(_RegFile_reg_15__7__m2s), .d(
        n3228), .sdi(n4242), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n944), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_15__7__slave ( .q(_RegFile_15__7), .qb(n4241), .d(
        _RegFile_reg_15__7__m2s), .g(Ctrl__Regs_1__en2), .rb(n944), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_15__8__master ( .q(_RegFile_reg_15__8__m2s), .d(
        n3229), .sdi(n4241), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n960), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_15__8__slave ( .q(_RegFile_15__8), .qb(n2030), .d(
        _RegFile_reg_15__8__m2s), .g(Ctrl__Regs_1__en2), .rb(n960), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_15__9__master ( .q(_RegFile_reg_15__9__m2s), .d(
        n3230), .sdi(n2030), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n944), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_15__9__slave ( .q(_RegFile_15__9), .qb(n2031), .d(
        _RegFile_reg_15__9__m2s), .g(Ctrl__Regs_1__en2), .rb(n944), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_16__0__master ( .q(_RegFile_reg_16__0__m2s), .d(
        n3189), .sdi(n2029), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n960), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_16__0__slave ( .q(_RegFile_16__0), .qb(n4240), .d(
        _RegFile_reg_16__0__m2s), .g(Ctrl__Regs_1__en2), .rb(n960), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_16__10__master ( .q(_RegFile_reg_16__10__m2s), .d(
        n3199), .sdi(n2055), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n960), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_16__10__slave ( .q(_RegFile_16__10), .qb(n2032), .d(
        _RegFile_reg_16__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n960), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_16__11__master ( .q(_RegFile_reg_16__11__m2s), .d(
        n3200), .sdi(n2032), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n944), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_16__11__slave ( .q(_RegFile_16__11), .qb(n2033), .d(
        _RegFile_reg_16__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n944), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_16__12__master ( .q(_RegFile_reg_16__12__m2s), .d(
        n3201), .sdi(n2033), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n960), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_16__12__slave ( .q(_RegFile_16__12), .qb(n2034), .d(
        _RegFile_reg_16__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n960), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_16__13__master ( .q(_RegFile_reg_16__13__m2s), .d(
        n3202), .sdi(n2034), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n944), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_16__13__slave ( .q(_RegFile_16__13), .qb(n2035), .d(
        _RegFile_reg_16__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n944), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_16__14__master ( .q(_RegFile_reg_16__14__m2s), .d(
        n3203), .sdi(n2035), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n960), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_16__14__slave ( .q(_RegFile_16__14), .qb(n2036), .d(
        _RegFile_reg_16__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n960), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_16__15__master ( .q(_RegFile_reg_16__15__m2s), .d(
        n3204), .sdi(n2036), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n944), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_16__15__slave ( .q(_RegFile_16__15), .qb(n2037), .d(
        _RegFile_reg_16__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n944), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_16__16__master ( .q(_RegFile_reg_16__16__m2s), .d(
        n3205), .sdi(n2037), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n960), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_16__16__slave ( .q(_RegFile_16__16), .qb(n2038), .d(
        _RegFile_reg_16__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n960), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_16__17__master ( .q(_RegFile_reg_16__17__m2s), .d(
        n3206), .sdi(n2038), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n943), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_16__17__slave ( .q(_RegFile_16__17), .qb(n2039), .d(
        _RegFile_reg_16__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n943), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_16__18__master ( .q(_RegFile_reg_16__18__m2s), .d(
        n3207), .sdi(n2039), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n960), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_16__18__slave ( .q(_RegFile_16__18), .qb(n2040), .d(
        _RegFile_reg_16__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n960), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_16__19__master ( .q(_RegFile_reg_16__19__m2s), .d(
        n3208), .sdi(n2040), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n943), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_16__19__slave ( .q(_RegFile_16__19), .qb(n2041), .d(
        _RegFile_reg_16__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n943), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_16__1__master ( .q(_RegFile_reg_16__1__m2s), .d(
        n3190), .sdi(n4240), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n944), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_16__1__slave ( .q(_RegFile_16__1), .qb(n4239), .d(
        _RegFile_reg_16__1__m2s), .g(Ctrl__Regs_1__en2), .rb(n944), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_16__20__master ( .q(_RegFile_reg_16__20__m2s), .d(
        n3209), .sdi(n2041), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n943), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_16__20__slave ( .q(_RegFile_16__20), .qb(n2042), .d(
        _RegFile_reg_16__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n943), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_16__21__master ( .q(_RegFile_reg_16__21__m2s), .d(
        n3210), .sdi(n2042), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n960), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_16__21__slave ( .q(_RegFile_16__21), .qb(n2043), .d(
        _RegFile_reg_16__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n960), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_16__22__master ( .q(_RegFile_reg_16__22__m2s), .d(
        n3211), .sdi(n2043), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n943), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_16__22__slave ( .q(_RegFile_16__22), .qb(n2044), .d(
        _RegFile_reg_16__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n943), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_16__23__master ( .q(_RegFile_reg_16__23__m2s), .d(
        n3212), .sdi(n2044), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n960), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_16__23__slave ( .q(_RegFile_16__23), .qb(n2045), .d(
        _RegFile_reg_16__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n960), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_16__24__master ( .q(_RegFile_reg_16__24__m2s), .d(
        n3213), .sdi(n2045), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n943), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_16__24__slave ( .q(_RegFile_16__24), .qb(n2046), .d(
        _RegFile_reg_16__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n943), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_16__25__master ( .q(_RegFile_reg_16__25__m2s), .d(
        n3214), .sdi(n2046), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n960), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_16__25__slave ( .q(_RegFile_16__25), .qb(n2047), .d(
        _RegFile_reg_16__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n960), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_16__26__master ( .q(_RegFile_reg_16__26__m2s), .d(
        n3215), .sdi(n2047), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n943), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_16__26__slave ( .q(_RegFile_16__26), .qb(n2048), .d(
        _RegFile_reg_16__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n943), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_16__27__master ( .q(_RegFile_reg_16__27__m2s), .d(
        n3216), .sdi(n2048), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n960), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_16__27__slave ( .q(_RegFile_16__27), .qb(n2049), .d(
        _RegFile_reg_16__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n960), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_16__28__master ( .q(_RegFile_reg_16__28__m2s), .d(
        n3217), .sdi(n2049), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n943), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_16__28__slave ( .q(_RegFile_16__28), .qb(n2050), .d(
        _RegFile_reg_16__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n943), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_16__29__master ( .q(_RegFile_reg_16__29__m2s), .d(
        n3218), .sdi(n2050), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n960), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_16__29__slave ( .q(_RegFile_16__29), .qb(n2051), .d(
        _RegFile_reg_16__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n960), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_16__2__master ( .q(_RegFile_reg_16__2__m2s), .d(
        n3191), .sdi(n4239), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n960), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_16__2__slave ( .q(_RegFile_16__2), .qb(n4238), .d(
        _RegFile_reg_16__2__m2s), .g(Ctrl__Regs_1__en2), .rb(n960), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_16__30__master ( .q(_RegFile_reg_16__30__m2s), .d(
        n3219), .sdi(n2051), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_16__30__slave ( .q(_RegFile_16__30), .qb(n2052), .d(
        _RegFile_reg_16__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_16__31__master ( .q(_RegFile_reg_16__31__m2s), .d(
        n3220), .sdi(n2052), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n943), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_16__31__slave ( .q(_RegFile_16__31), .qb(n2053), .d(
        _RegFile_reg_16__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n943), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_16__3__master ( .q(_RegFile_reg_16__3__m2s), .d(
        n3192), .sdi(n4238), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n943), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_16__3__slave ( .q(_RegFile_16__3), .qb(n4237), .d(
        _RegFile_reg_16__3__m2s), .g(Ctrl__Regs_1__en2), .rb(n943), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_16__4__master ( .q(_RegFile_reg_16__4__m2s), .d(
        n3193), .sdi(n4237), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_16__4__slave ( .q(_RegFile_16__4), .qb(n4236), .d(
        _RegFile_reg_16__4__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_16__5__master ( .q(_RegFile_reg_16__5__m2s), .d(
        n3194), .sdi(n4236), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n943), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_16__5__slave ( .q(_RegFile_16__5), .qb(n4235), .d(
        _RegFile_reg_16__5__m2s), .g(Ctrl__Regs_1__en2), .rb(n943), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_16__6__master ( .q(_RegFile_reg_16__6__m2s), .d(
        n3195), .sdi(n4235), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_16__6__slave ( .q(_RegFile_16__6), .qb(n4234), .d(
        _RegFile_reg_16__6__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_16__7__master ( .q(_RegFile_reg_16__7__m2s), .d(
        n3196), .sdi(n4234), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n943), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_16__7__slave ( .q(_RegFile_16__7), .qb(n4233), .d(
        _RegFile_reg_16__7__m2s), .g(Ctrl__Regs_1__en2), .rb(n943), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_16__8__master ( .q(_RegFile_reg_16__8__m2s), .d(
        n3197), .sdi(n4233), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_16__8__slave ( .q(_RegFile_16__8), .qb(n2054), .d(
        _RegFile_reg_16__8__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_16__9__master ( .q(_RegFile_reg_16__9__m2s), .d(
        n3198), .sdi(n2054), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n943), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_16__9__slave ( .q(_RegFile_16__9), .qb(n2055), .d(
        _RegFile_reg_16__9__m2s), .g(Ctrl__Regs_1__en2), .rb(n943), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_17__0__master ( .q(_RegFile_reg_17__0__m2s), .d(
        n3157), .sdi(n2053), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_17__0__slave ( .q(_RegFile_17__0), .qb(n4232), .d(
        _RegFile_reg_17__0__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_17__10__master ( .q(_RegFile_reg_17__10__m2s), .d(
        n3167), .sdi(n2079), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_17__10__slave ( .q(_RegFile_17__10), .qb(n2056), .d(
        _RegFile_reg_17__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_17__11__master ( .q(_RegFile_reg_17__11__m2s), .d(
        n3168), .sdi(n2056), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n943), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_17__11__slave ( .q(_RegFile_17__11), .qb(n2057), .d(
        _RegFile_reg_17__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n943), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_17__12__master ( .q(_RegFile_reg_17__12__m2s), .d(
        n3169), .sdi(n2057), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_17__12__slave ( .q(_RegFile_17__12), .qb(n2058), .d(
        _RegFile_reg_17__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_17__13__master ( .q(_RegFile_reg_17__13__m2s), .d(
        n3170), .sdi(n2058), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n943), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_17__13__slave ( .q(_RegFile_17__13), .qb(n2059), .d(
        _RegFile_reg_17__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n943), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_17__14__master ( .q(_RegFile_reg_17__14__m2s), .d(
        n3171), .sdi(n2059), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_17__14__slave ( .q(_RegFile_17__14), .qb(n2060), .d(
        _RegFile_reg_17__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_17__15__master ( .q(_RegFile_reg_17__15__m2s), .d(
        n3172), .sdi(n2060), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n942), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_17__15__slave ( .q(_RegFile_17__15), .qb(n2061), .d(
        _RegFile_reg_17__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n942), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_17__16__master ( .q(_RegFile_reg_17__16__m2s), .d(
        n3173), .sdi(n2061), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_17__16__slave ( .q(_RegFile_17__16), .qb(n2062), .d(
        _RegFile_reg_17__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_17__17__master ( .q(_RegFile_reg_17__17__m2s), .d(
        n3174), .sdi(n2062), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n942), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_17__17__slave ( .q(_RegFile_17__17), .qb(n2063), .d(
        _RegFile_reg_17__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n942), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_17__18__master ( .q(_RegFile_reg_17__18__m2s), .d(
        n3175), .sdi(n2063), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_17__18__slave ( .q(_RegFile_17__18), .qb(n2064), .d(
        _RegFile_reg_17__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_17__19__master ( .q(_RegFile_reg_17__19__m2s), .d(
        n3176), .sdi(n2064), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n942), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_17__19__slave ( .q(_RegFile_17__19), .qb(n2065), .d(
        _RegFile_reg_17__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n942), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_17__1__master ( .q(_RegFile_reg_17__1__m2s), .d(
        n3158), .sdi(n4232), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n943), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_17__1__slave ( .q(_RegFile_17__1), .qb(n4231), .d(
        _RegFile_reg_17__1__m2s), .g(Ctrl__Regs_1__en2), .rb(n943), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_17__20__master ( .q(_RegFile_reg_17__20__m2s), .d(
        n3177), .sdi(n2065), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n942), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_17__20__slave ( .q(_RegFile_17__20), .qb(n2066), .d(
        _RegFile_reg_17__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n942), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_17__21__master ( .q(_RegFile_reg_17__21__m2s), .d(
        n3178), .sdi(n2066), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_17__21__slave ( .q(_RegFile_17__21), .qb(n2067), .d(
        _RegFile_reg_17__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_17__22__master ( .q(_RegFile_reg_17__22__m2s), .d(
        n3179), .sdi(n2067), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n942), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_17__22__slave ( .q(_RegFile_17__22), .qb(n2068), .d(
        _RegFile_reg_17__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n942), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_17__23__master ( .q(_RegFile_reg_17__23__m2s), .d(
        n3180), .sdi(n2068), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_17__23__slave ( .q(_RegFile_17__23), .qb(n2069), .d(
        _RegFile_reg_17__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_17__24__master ( .q(_RegFile_reg_17__24__m2s), .d(
        n3181), .sdi(n2069), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n942), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_17__24__slave ( .q(_RegFile_17__24), .qb(n2070), .d(
        _RegFile_reg_17__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n942), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_17__25__master ( .q(_RegFile_reg_17__25__m2s), .d(
        n3182), .sdi(n2070), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_17__25__slave ( .q(_RegFile_17__25), .qb(n2071), .d(
        _RegFile_reg_17__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_17__26__master ( .q(_RegFile_reg_17__26__m2s), .d(
        n3183), .sdi(n2071), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n942), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_17__26__slave ( .q(_RegFile_17__26), .qb(n2072), .d(
        _RegFile_reg_17__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n942), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_17__27__master ( .q(_RegFile_reg_17__27__m2s), .d(
        n3184), .sdi(n2072), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_17__27__slave ( .q(_RegFile_17__27), .qb(n2073), .d(
        _RegFile_reg_17__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_17__28__master ( .q(_RegFile_reg_17__28__m2s), .d(
        n3185), .sdi(n2073), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n942), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_17__28__slave ( .q(_RegFile_17__28), .qb(n2074), .d(
        _RegFile_reg_17__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n942), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_17__29__master ( .q(_RegFile_reg_17__29__m2s), .d(
        n3186), .sdi(n2074), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n961), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_17__29__slave ( .q(_RegFile_17__29), .qb(n2075), .d(
        _RegFile_reg_17__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n961), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_17__2__master ( .q(_RegFile_reg_17__2__m2s), .d(
        n3159), .sdi(n4231), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_17__2__slave ( .q(_RegFile_17__2), .qb(n4230), .d(
        _RegFile_reg_17__2__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_17__30__master ( .q(_RegFile_reg_17__30__m2s), .d(
        n3187), .sdi(n2075), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n961), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_17__30__slave ( .q(_RegFile_17__30), .qb(n2076), .d(
        _RegFile_reg_17__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n961), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_17__31__master ( .q(_RegFile_reg_17__31__m2s), .d(
        n3188), .sdi(n2076), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n942), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_17__31__slave ( .q(_RegFile_17__31), .qb(n2077), .d(
        _RegFile_reg_17__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n942), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_17__3__master ( .q(_RegFile_reg_17__3__m2s), .d(
        n3160), .sdi(n4230), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n942), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_17__3__slave ( .q(_RegFile_17__3), .qb(n4229), .d(
        _RegFile_reg_17__3__m2s), .g(Ctrl__Regs_1__en2), .rb(n942), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_17__4__master ( .q(_RegFile_reg_17__4__m2s), .d(
        n3161), .sdi(n4229), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n961), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_17__4__slave ( .q(_RegFile_17__4), .qb(n4228), .d(
        _RegFile_reg_17__4__m2s), .g(Ctrl__Regs_1__en2), .rb(n961), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_17__5__master ( .q(_RegFile_reg_17__5__m2s), .d(
        n3162), .sdi(n4228), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n942), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_17__5__slave ( .q(_RegFile_17__5), .qb(n4227), .d(
        _RegFile_reg_17__5__m2s), .g(Ctrl__Regs_1__en2), .rb(n942), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_17__6__master ( .q(_RegFile_reg_17__6__m2s), .d(
        n3163), .sdi(n4227), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n961), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_17__6__slave ( .q(_RegFile_17__6), .qb(n4226), .d(
        _RegFile_reg_17__6__m2s), .g(Ctrl__Regs_1__en2), .rb(n961), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_17__7__master ( .q(_RegFile_reg_17__7__m2s), .d(
        n3164), .sdi(n4226), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n942), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_17__7__slave ( .q(_RegFile_17__7), .qb(n4225), .d(
        _RegFile_reg_17__7__m2s), .g(Ctrl__Regs_1__en2), .rb(n942), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_17__8__master ( .q(_RegFile_reg_17__8__m2s), .d(
        n3165), .sdi(n4225), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n961), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_17__8__slave ( .q(_RegFile_17__8), .qb(n2078), .d(
        _RegFile_reg_17__8__m2s), .g(Ctrl__Regs_1__en2), .rb(n961), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_17__9__master ( .q(_RegFile_reg_17__9__m2s), .d(
        n3166), .sdi(n2078), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n942), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_17__9__slave ( .q(_RegFile_17__9), .qb(n2079), .d(
        _RegFile_reg_17__9__m2s), .g(Ctrl__Regs_1__en2), .rb(n942), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_18__0__master ( .q(_RegFile_reg_18__0__m2s), .d(
        n3125), .sdi(n2077), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n961), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_18__0__slave ( .q(_RegFile_18__0), .qb(n4224), .d(
        _RegFile_reg_18__0__m2s), .g(Ctrl__Regs_1__en2), .rb(n961), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_18__10__master ( .q(_RegFile_reg_18__10__m2s), .d(
        n3135), .sdi(n2103), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n961), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_18__10__slave ( .q(_RegFile_18__10), .qb(n2080), .d(
        _RegFile_reg_18__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n961), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_18__11__master ( .q(_RegFile_reg_18__11__m2s), .d(
        n3136), .sdi(n2080), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n942), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_18__11__slave ( .q(_RegFile_18__11), .qb(n2081), .d(
        _RegFile_reg_18__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n942), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_18__12__master ( .q(_RegFile_reg_18__12__m2s), .d(
        n3137), .sdi(n2081), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n961), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_18__12__slave ( .q(_RegFile_18__12), .qb(n2082), .d(
        _RegFile_reg_18__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n961), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_18__13__master ( .q(_RegFile_reg_18__13__m2s), .d(
        n3138), .sdi(n2082), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n941), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_18__13__slave ( .q(_RegFile_18__13), .qb(n2083), .d(
        _RegFile_reg_18__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n941), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_18__14__master ( .q(_RegFile_reg_18__14__m2s), .d(
        n3139), .sdi(n2083), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n961), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_18__14__slave ( .q(_RegFile_18__14), .qb(n2084), .d(
        _RegFile_reg_18__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n961), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_18__15__master ( .q(_RegFile_reg_18__15__m2s), .d(
        n3140), .sdi(n2084), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n941), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_18__15__slave ( .q(_RegFile_18__15), .qb(n2085), .d(
        _RegFile_reg_18__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n941), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_18__16__master ( .q(_RegFile_reg_18__16__m2s), .d(
        n3141), .sdi(n2085), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n961), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_18__16__slave ( .q(_RegFile_18__16), .qb(n2086), .d(
        _RegFile_reg_18__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n961), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_18__17__master ( .q(_RegFile_reg_18__17__m2s), .d(
        n3142), .sdi(n2086), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n941), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_18__17__slave ( .q(_RegFile_18__17), .qb(n2087), .d(
        _RegFile_reg_18__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n941), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_18__18__master ( .q(_RegFile_reg_18__18__m2s), .d(
        n3143), .sdi(n2087), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n961), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_18__18__slave ( .q(_RegFile_18__18), .qb(n2088), .d(
        _RegFile_reg_18__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n961), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_18__19__master ( .q(_RegFile_reg_18__19__m2s), .d(
        n3144), .sdi(n2088), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n941), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_18__19__slave ( .q(_RegFile_18__19), .qb(n2089), .d(
        _RegFile_reg_18__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n941), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_18__1__master ( .q(_RegFile_reg_18__1__m2s), .d(
        n3126), .sdi(n4224), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n942), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_18__1__slave ( .q(_RegFile_18__1), .qb(n4223), .d(
        _RegFile_reg_18__1__m2s), .g(Ctrl__Regs_1__en2), .rb(n942), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_18__20__master ( .q(_RegFile_reg_18__20__m2s), .d(
        n3145), .sdi(n2089), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n941), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_18__20__slave ( .q(_RegFile_18__20), .qb(n2090), .d(
        _RegFile_reg_18__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n941), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_18__21__master ( .q(_RegFile_reg_18__21__m2s), .d(
        n3146), .sdi(n2090), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n961), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_18__21__slave ( .q(_RegFile_18__21), .qb(n2091), .d(
        _RegFile_reg_18__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n961), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_18__22__master ( .q(_RegFile_reg_18__22__m2s), .d(
        n3147), .sdi(n2091), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n941), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_18__22__slave ( .q(_RegFile_18__22), .qb(n2092), .d(
        _RegFile_reg_18__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n941), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_18__23__master ( .q(_RegFile_reg_18__23__m2s), .d(
        n3148), .sdi(n2092), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n961), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_18__23__slave ( .q(_RegFile_18__23), .qb(n2093), .d(
        _RegFile_reg_18__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n961), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_18__24__master ( .q(_RegFile_reg_18__24__m2s), .d(
        n3149), .sdi(n2093), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n941), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_18__24__slave ( .q(_RegFile_18__24), .qb(n2094), .d(
        _RegFile_reg_18__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n941), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_18__25__master ( .q(_RegFile_reg_18__25__m2s), .d(
        n3150), .sdi(n2094), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n961), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_18__25__slave ( .q(_RegFile_18__25), .qb(n2095), .d(
        _RegFile_reg_18__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n961), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_18__26__master ( .q(_RegFile_reg_18__26__m2s), .d(
        n3151), .sdi(n2095), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n941), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_18__26__slave ( .q(_RegFile_18__26), .qb(n2096), .d(
        _RegFile_reg_18__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n941), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_18__27__master ( .q(_RegFile_reg_18__27__m2s), .d(
        n3152), .sdi(n2096), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_18__27__slave ( .q(_RegFile_18__27), .qb(n2097), .d(
        _RegFile_reg_18__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_18__28__master ( .q(_RegFile_reg_18__28__m2s), .d(
        n3153), .sdi(n2097), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n941), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_18__28__slave ( .q(_RegFile_18__28), .qb(n2098), .d(
        _RegFile_reg_18__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n941), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_18__29__master ( .q(_RegFile_reg_18__29__m2s), .d(
        n3154), .sdi(n2098), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_18__29__slave ( .q(_RegFile_18__29), .qb(n2099), .d(
        _RegFile_reg_18__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_18__2__master ( .q(_RegFile_reg_18__2__m2s), .d(
        n3127), .sdi(n4223), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n961), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_18__2__slave ( .q(_RegFile_18__2), .qb(n4222), .d(
        _RegFile_reg_18__2__m2s), .g(Ctrl__Regs_1__en2), .rb(n961), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_18__30__master ( .q(_RegFile_reg_18__30__m2s), .d(
        n3155), .sdi(n2099), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_18__30__slave ( .q(_RegFile_18__30), .qb(n2100), .d(
        _RegFile_reg_18__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_18__31__master ( .q(_RegFile_reg_18__31__m2s), .d(
        n3156), .sdi(n2100), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n941), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_18__31__slave ( .q(_RegFile_18__31), .qb(n2101), .d(
        _RegFile_reg_18__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n941), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_18__3__master ( .q(_RegFile_reg_18__3__m2s), .d(
        n3128), .sdi(n4222), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n941), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_18__3__slave ( .q(_RegFile_18__3), .qb(n4221), .d(
        _RegFile_reg_18__3__m2s), .g(Ctrl__Regs_1__en2), .rb(n941), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_18__4__master ( .q(_RegFile_reg_18__4__m2s), .d(
        n3129), .sdi(n4221), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_18__4__slave ( .q(_RegFile_18__4), .qb(n4220), .d(
        _RegFile_reg_18__4__m2s), .g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_18__5__master ( .q(_RegFile_reg_18__5__m2s), .d(
        n3130), .sdi(n4220), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n941), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_18__5__slave ( .q(_RegFile_18__5), .qb(n4219), .d(
        _RegFile_reg_18__5__m2s), .g(Ctrl__Regs_1__en2), .rb(n941), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_18__6__master ( .q(_RegFile_reg_18__6__m2s), .d(
        n3131), .sdi(n4219), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_18__6__slave ( .q(_RegFile_18__6), .qb(n4218), .d(
        _RegFile_reg_18__6__m2s), .g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_18__7__master ( .q(_RegFile_reg_18__7__m2s), .d(
        n3132), .sdi(n4218), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n941), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_18__7__slave ( .q(_RegFile_18__7), .qb(n4217), .d(
        _RegFile_reg_18__7__m2s), .g(Ctrl__Regs_1__en2), .rb(n941), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_18__8__master ( .q(_RegFile_reg_18__8__m2s), .d(
        n3133), .sdi(n4217), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_18__8__slave ( .q(_RegFile_18__8), .qb(n2102), .d(
        _RegFile_reg_18__8__m2s), .g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_18__9__master ( .q(_RegFile_reg_18__9__m2s), .d(
        n3134), .sdi(n2102), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n941), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_18__9__slave ( .q(_RegFile_18__9), .qb(n2103), .d(
        _RegFile_reg_18__9__m2s), .g(Ctrl__Regs_1__en2), .rb(n941), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_19__0__master ( .q(_RegFile_reg_19__0__m2s), .d(
        n3093), .sdi(n2101), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_19__0__slave ( .q(_RegFile_19__0), .qb(n4216), .d(
        _RegFile_reg_19__0__m2s), .g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_19__10__master ( .q(_RegFile_reg_19__10__m2s), .d(
        n3103), .sdi(n2127), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_19__10__slave ( .q(_RegFile_19__10), .qb(n2104), .d(
        _RegFile_reg_19__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_19__11__master ( .q(_RegFile_reg_19__11__m2s), .d(
        n3104), .sdi(n2104), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n940), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_19__11__slave ( .q(_RegFile_19__11), .qb(n2105), .d(
        _RegFile_reg_19__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n940), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_19__12__master ( .q(_RegFile_reg_19__12__m2s), .d(
        n3105), .sdi(n2105), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_19__12__slave ( .q(_RegFile_19__12), .qb(n2106), .d(
        _RegFile_reg_19__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_19__13__master ( .q(_RegFile_reg_19__13__m2s), .d(
        n3106), .sdi(n2106), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n940), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_19__13__slave ( .q(_RegFile_19__13), .qb(n2107), .d(
        _RegFile_reg_19__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n940), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_19__14__master ( .q(_RegFile_reg_19__14__m2s), .d(
        n3107), .sdi(n2107), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_19__14__slave ( .q(_RegFile_19__14), .qb(n2108), .d(
        _RegFile_reg_19__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_19__15__master ( .q(_RegFile_reg_19__15__m2s), .d(
        n3108), .sdi(n2108), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n940), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_19__15__slave ( .q(_RegFile_19__15), .qb(n2109), .d(
        _RegFile_reg_19__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n940), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_19__16__master ( .q(_RegFile_reg_19__16__m2s), .d(
        n3109), .sdi(n2109), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_19__16__slave ( .q(_RegFile_19__16), .qb(n2110), .d(
        _RegFile_reg_19__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_19__17__master ( .q(_RegFile_reg_19__17__m2s), .d(
        n3110), .sdi(n2110), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n940), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_19__17__slave ( .q(_RegFile_19__17), .qb(n2111), .d(
        _RegFile_reg_19__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n940), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_19__18__master ( .q(_RegFile_reg_19__18__m2s), .d(
        n3111), .sdi(n2111), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_19__18__slave ( .q(_RegFile_19__18), .qb(n2112), .d(
        _RegFile_reg_19__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_19__19__master ( .q(_RegFile_reg_19__19__m2s), .d(
        n3112), .sdi(n2112), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n940), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_19__19__slave ( .q(_RegFile_19__19), .qb(n2113), .d(
        _RegFile_reg_19__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n940), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_19__1__master ( .q(_RegFile_reg_19__1__m2s), .d(
        n3094), .sdi(n4216), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n941), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_19__1__slave ( .q(_RegFile_19__1), .qb(n4215), .d(
        _RegFile_reg_19__1__m2s), .g(Ctrl__Regs_1__en2), .rb(n941), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_19__20__master ( .q(_RegFile_reg_19__20__m2s), .d(
        n3113), .sdi(n2113), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n940), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_19__20__slave ( .q(_RegFile_19__20), .qb(n2114), .d(
        _RegFile_reg_19__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n940), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_19__21__master ( .q(_RegFile_reg_19__21__m2s), .d(
        n3114), .sdi(n2114), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_19__21__slave ( .q(_RegFile_19__21), .qb(n2115), .d(
        _RegFile_reg_19__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_19__22__master ( .q(_RegFile_reg_19__22__m2s), .d(
        n3115), .sdi(n2115), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n940), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_19__22__slave ( .q(_RegFile_19__22), .qb(n2116), .d(
        _RegFile_reg_19__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n940), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_19__23__master ( .q(_RegFile_reg_19__23__m2s), .d(
        n3116), .sdi(n2116), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_19__23__slave ( .q(_RegFile_19__23), .qb(n2117), .d(
        _RegFile_reg_19__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_19__24__master ( .q(_RegFile_reg_19__24__m2s), .d(
        n3117), .sdi(n2117), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n940), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_19__24__slave ( .q(_RegFile_19__24), .qb(n2118), .d(
        _RegFile_reg_19__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n940), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_19__25__master ( .q(_RegFile_reg_19__25__m2s), .d(
        n3118), .sdi(n2118), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n962), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_19__25__slave ( .q(_RegFile_19__25), .qb(n2119), .d(
        _RegFile_reg_19__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n962), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_19__26__master ( .q(_RegFile_reg_19__26__m2s), .d(
        n3119), .sdi(n2119), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n940), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_19__26__slave ( .q(_RegFile_19__26), .qb(n2120), .d(
        _RegFile_reg_19__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n940), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_19__27__master ( .q(_RegFile_reg_19__27__m2s), .d(
        n3120), .sdi(n2120), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n962), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_19__27__slave ( .q(_RegFile_19__27), .qb(n2121), .d(
        _RegFile_reg_19__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n962), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_19__28__master ( .q(_RegFile_reg_19__28__m2s), .d(
        n3121), .sdi(n2121), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n940), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_19__28__slave ( .q(_RegFile_19__28), .qb(n2122), .d(
        _RegFile_reg_19__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n940), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_19__29__master ( .q(_RegFile_reg_19__29__m2s), .d(
        n3122), .sdi(n2122), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n962), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_19__29__slave ( .q(_RegFile_19__29), .qb(n2123), .d(
        _RegFile_reg_19__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n962), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_19__2__master ( .q(_RegFile_reg_19__2__m2s), .d(
        n3095), .sdi(n4215), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_19__2__slave ( .q(_RegFile_19__2), .qb(n4214), .d(
        _RegFile_reg_19__2__m2s), .g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_19__30__master ( .q(_RegFile_reg_19__30__m2s), .d(
        n3123), .sdi(n2123), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n962), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_19__30__slave ( .q(_RegFile_19__30), .qb(n2124), .d(
        _RegFile_reg_19__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n962), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_19__31__master ( .q(_RegFile_reg_19__31__m2s), .d(
        n3124), .sdi(n2124), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n940), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_19__31__slave ( .q(_RegFile_19__31), .qb(n2125), .d(
        _RegFile_reg_19__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n940), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_19__3__master ( .q(_RegFile_reg_19__3__m2s), .d(
        n3096), .sdi(n4214), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n940), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_19__3__slave ( .q(_RegFile_19__3), .qb(n4213), .d(
        _RegFile_reg_19__3__m2s), .g(Ctrl__Regs_1__en2), .rb(n940), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_19__4__master ( .q(_RegFile_reg_19__4__m2s), .d(
        n3097), .sdi(n4213), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n962), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_19__4__slave ( .q(_RegFile_19__4), .qb(n4212), .d(
        _RegFile_reg_19__4__m2s), .g(Ctrl__Regs_1__en2), .rb(n962), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_19__5__master ( .q(_RegFile_reg_19__5__m2s), .d(
        n3098), .sdi(n4212), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n940), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_19__5__slave ( .q(_RegFile_19__5), .qb(n4211), .d(
        _RegFile_reg_19__5__m2s), .g(Ctrl__Regs_1__en2), .rb(n940), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_19__6__master ( .q(_RegFile_reg_19__6__m2s), .d(
        n3099), .sdi(n4211), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n962), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_19__6__slave ( .q(_RegFile_19__6), .qb(n4210), .d(
        _RegFile_reg_19__6__m2s), .g(Ctrl__Regs_1__en2), .rb(n962), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_19__7__master ( .q(_RegFile_reg_19__7__m2s), .d(
        n3100), .sdi(n4210), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n940), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_19__7__slave ( .q(_RegFile_19__7), .qb(n4209), .d(
        _RegFile_reg_19__7__m2s), .g(Ctrl__Regs_1__en2), .rb(n940), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_19__8__master ( .q(_RegFile_reg_19__8__m2s), .d(
        n3101), .sdi(n4209), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n962), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_19__8__slave ( .q(_RegFile_19__8), .qb(n2126), .d(
        _RegFile_reg_19__8__m2s), .g(Ctrl__Regs_1__en2), .rb(n962), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_19__9__master ( .q(_RegFile_reg_19__9__m2s), .d(
        n3102), .sdi(n2126), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n940), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_19__9__slave ( .q(_RegFile_19__9), .qb(n2127), .d(
        _RegFile_reg_19__9__m2s), .g(Ctrl__Regs_1__en2), .rb(n940), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_1__0__master ( .q(_RegFile_reg_1__0__m2s), .d(n3669
        ), .sdi(n1885), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n962), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_1__0__slave ( .q(_RegFile_1__0), .qb(n4360), .d(
        _RegFile_reg_1__0__m2s), .g(Ctrl__Regs_1__en2), .rb(n962), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_1__10__master ( .q(_RegFile_reg_1__10__m2s), .d(
        n3679), .sdi(n2151), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n962), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_1__10__slave ( .q(_RegFile_1__10), .qb(n2128), .d(
        _RegFile_reg_1__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n962), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_1__11__master ( .q(_RegFile_reg_1__11__m2s), .d(
        n3680), .sdi(n2128), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n939), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_1__11__slave ( .q(_RegFile_1__11), .qb(n2129), .d(
        _RegFile_reg_1__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n939), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_1__12__master ( .q(_RegFile_reg_1__12__m2s), .d(
        n3681), .sdi(n2129), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n962), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_1__12__slave ( .q(_RegFile_1__12), .qb(n2130), .d(
        _RegFile_reg_1__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n962), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_1__13__master ( .q(_RegFile_reg_1__13__m2s), .d(
        n3682), .sdi(n2130), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n939), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_1__13__slave ( .q(_RegFile_1__13), .qb(n2131), .d(
        _RegFile_reg_1__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n939), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_1__14__master ( .q(_RegFile_reg_1__14__m2s), .d(
        n3683), .sdi(n2131), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n962), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_1__14__slave ( .q(_RegFile_1__14), .qb(n2132), .d(
        _RegFile_reg_1__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n962), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_1__15__master ( .q(_RegFile_reg_1__15__m2s), .d(
        n3684), .sdi(n2132), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n939), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_1__15__slave ( .q(_RegFile_1__15), .qb(n2133), .d(
        _RegFile_reg_1__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n939), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_1__16__master ( .q(_RegFile_reg_1__16__m2s), .d(
        n3685), .sdi(n2133), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n962), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_1__16__slave ( .q(_RegFile_1__16), .qb(n2134), .d(
        _RegFile_reg_1__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n962), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_1__17__master ( .q(_RegFile_reg_1__17__m2s), .d(
        n3686), .sdi(n2134), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n939), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_1__17__slave ( .q(_RegFile_1__17), .qb(n2135), .d(
        _RegFile_reg_1__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n939), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_1__18__master ( .q(_RegFile_reg_1__18__m2s), .d(
        n3687), .sdi(n2135), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n962), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_1__18__slave ( .q(_RegFile_1__18), .qb(n2136), .d(
        _RegFile_reg_1__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n962), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_1__19__master ( .q(_RegFile_reg_1__19__m2s), .d(
        n3688), .sdi(n2136), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n939), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_1__19__slave ( .q(_RegFile_1__19), .qb(n2137), .d(
        _RegFile_reg_1__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n939), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_1__1__master ( .q(_RegFile_reg_1__1__m2s), .d(n3670
        ), .sdi(n4360), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n939), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_1__1__slave ( .q(_RegFile_1__1), .qb(n4359), .d(
        _RegFile_reg_1__1__m2s), .g(Ctrl__Regs_1__en2), .rb(n939), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_1__20__master ( .q(_RegFile_reg_1__20__m2s), .d(
        n3689), .sdi(n2137), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n939), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_1__20__slave ( .q(_RegFile_1__20), .qb(n2138), .d(
        _RegFile_reg_1__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n939), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_1__21__master ( .q(_RegFile_reg_1__21__m2s), .d(
        n3690), .sdi(n2138), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n962), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_1__21__slave ( .q(_RegFile_1__21), .qb(n2139), .d(
        _RegFile_reg_1__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n962), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_1__22__master ( .q(_RegFile_reg_1__22__m2s), .d(
        n3691), .sdi(n2139), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n939), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_1__22__slave ( .q(_RegFile_1__22), .qb(n2140), .d(
        _RegFile_reg_1__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n939), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_1__23__master ( .q(_RegFile_reg_1__23__m2s), .d(
        n3692), .sdi(n2140), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n963), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_1__23__slave ( .q(_RegFile_1__23), .qb(n2141), .d(
        _RegFile_reg_1__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n963), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_1__24__master ( .q(_RegFile_reg_1__24__m2s), .d(
        n3693), .sdi(n2141), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n939), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_1__24__slave ( .q(_RegFile_1__24), .qb(n2142), .d(
        _RegFile_reg_1__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n939), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_1__25__master ( .q(_RegFile_reg_1__25__m2s), .d(
        n3694), .sdi(n2142), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n963), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_1__25__slave ( .q(_RegFile_1__25), .qb(n2143), .d(
        _RegFile_reg_1__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n963), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_1__26__master ( .q(_RegFile_reg_1__26__m2s), .d(
        n3695), .sdi(n2143), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n939), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_1__26__slave ( .q(_RegFile_1__26), .qb(n2144), .d(
        _RegFile_reg_1__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n939), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_1__27__master ( .q(_RegFile_reg_1__27__m2s), .d(
        n3696), .sdi(n2144), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n963), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_1__27__slave ( .q(_RegFile_1__27), .qb(n2145), .d(
        _RegFile_reg_1__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n963), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_1__28__master ( .q(_RegFile_reg_1__28__m2s), .d(
        n3697), .sdi(n2145), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n939), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_1__28__slave ( .q(_RegFile_1__28), .qb(n2146), .d(
        _RegFile_reg_1__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n939), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_1__29__master ( .q(_RegFile_reg_1__29__m2s), .d(
        n3698), .sdi(n2146), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n963), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_1__29__slave ( .q(_RegFile_1__29), .qb(n2147), .d(
        _RegFile_reg_1__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n963), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_1__2__master ( .q(_RegFile_reg_1__2__m2s), .d(n3671
        ), .sdi(n4359), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n962), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_1__2__slave ( .q(_RegFile_1__2), .qb(n4358), .d(
        _RegFile_reg_1__2__m2s), .g(Ctrl__Regs_1__en2), .rb(n962), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_1__30__master ( .q(_RegFile_reg_1__30__m2s), .d(
        n3699), .sdi(n2147), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n963), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_1__30__slave ( .q(_RegFile_1__30), .qb(n2148), .d(
        _RegFile_reg_1__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n963), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_1__31__master ( .q(_RegFile_reg_1__31__m2s), .d(
        n3700), .sdi(n2148), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n939), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_1__31__slave ( .q(_RegFile_1__31), .qb(n2149), .d(
        _RegFile_reg_1__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n939), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_1__3__master ( .q(_RegFile_reg_1__3__m2s), .d(n3672
        ), .sdi(n4358), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n939), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_1__3__slave ( .q(_RegFile_1__3), .qb(n4357), .d(
        _RegFile_reg_1__3__m2s), .g(Ctrl__Regs_1__en2), .rb(n939), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_1__4__master ( .q(_RegFile_reg_1__4__m2s), .d(n3673
        ), .sdi(n4357), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n963), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_1__4__slave ( .q(_RegFile_1__4), .qb(n4356), .d(
        _RegFile_reg_1__4__m2s), .g(Ctrl__Regs_1__en2), .rb(n963), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_1__5__master ( .q(_RegFile_reg_1__5__m2s), .d(n3674
        ), .sdi(n4356), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n939), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_1__5__slave ( .q(_RegFile_1__5), .qb(n4355), .d(
        _RegFile_reg_1__5__m2s), .g(Ctrl__Regs_1__en2), .rb(n939), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_1__6__master ( .q(_RegFile_reg_1__6__m2s), .d(n3675
        ), .sdi(n4355), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n963), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_1__6__slave ( .q(_RegFile_1__6), .qb(n4354), .d(
        _RegFile_reg_1__6__m2s), .g(Ctrl__Regs_1__en2), .rb(n963), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_1__7__master ( .q(_RegFile_reg_1__7__m2s), .d(n3676
        ), .sdi(n4354), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n939), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_1__7__slave ( .q(_RegFile_1__7), .qb(n4353), .d(
        _RegFile_reg_1__7__m2s), .g(Ctrl__Regs_1__en2), .rb(n939), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_1__8__master ( .q(_RegFile_reg_1__8__m2s), .d(n3677
        ), .sdi(n4353), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n963), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_1__8__slave ( .q(_RegFile_1__8), .qb(n2150), .d(
        _RegFile_reg_1__8__m2s), .g(Ctrl__Regs_1__en2), .rb(n963), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_1__9__master ( .q(_RegFile_reg_1__9__m2s), .d(n3678
        ), .sdi(n2150), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_1__9__slave ( .q(_RegFile_1__9), .qb(n2151), .d(
        _RegFile_reg_1__9__m2s), .g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_20__0__master ( .q(_RegFile_reg_20__0__m2s), .d(
        n3061), .sdi(n2125), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n963), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_20__0__slave ( .q(_RegFile_20__0), .qb(n4208), .d(
        _RegFile_reg_20__0__m2s), .g(Ctrl__Regs_1__en2), .rb(n963), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_20__10__master ( .q(_RegFile_reg_20__10__m2s), .d(
        n3071), .sdi(n2175), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n963), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_20__10__slave ( .q(_RegFile_20__10), .qb(n2152), .d(
        _RegFile_reg_20__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n963), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_20__11__master ( .q(_RegFile_reg_20__11__m2s), .d(
        n3072), .sdi(n2152), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_20__11__slave ( .q(_RegFile_20__11), .qb(n2153), .d(
        _RegFile_reg_20__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_20__12__master ( .q(_RegFile_reg_20__12__m2s), .d(
        n3073), .sdi(n2153), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n963), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_20__12__slave ( .q(_RegFile_20__12), .qb(n2154), .d(
        _RegFile_reg_20__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n963), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_20__13__master ( .q(_RegFile_reg_20__13__m2s), .d(
        n3074), .sdi(n2154), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_20__13__slave ( .q(_RegFile_20__13), .qb(n2155), .d(
        _RegFile_reg_20__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_20__14__master ( .q(_RegFile_reg_20__14__m2s), .d(
        n3075), .sdi(n2155), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n963), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_20__14__slave ( .q(_RegFile_20__14), .qb(n2156), .d(
        _RegFile_reg_20__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n963), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_20__15__master ( .q(_RegFile_reg_20__15__m2s), .d(
        n3076), .sdi(n2156), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_20__15__slave ( .q(_RegFile_20__15), .qb(n2157), .d(
        _RegFile_reg_20__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_20__16__master ( .q(_RegFile_reg_20__16__m2s), .d(
        n3077), .sdi(n2157), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n963), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_20__16__slave ( .q(_RegFile_20__16), .qb(n2158), .d(
        _RegFile_reg_20__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n963), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_20__17__master ( .q(_RegFile_reg_20__17__m2s), .d(
        n3078), .sdi(n2158), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_20__17__slave ( .q(_RegFile_20__17), .qb(n2159), .d(
        _RegFile_reg_20__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_20__18__master ( .q(_RegFile_reg_20__18__m2s), .d(
        n3079), .sdi(n2159), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n963), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_20__18__slave ( .q(_RegFile_20__18), .qb(n2160), .d(
        _RegFile_reg_20__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n963), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_20__19__master ( .q(_RegFile_reg_20__19__m2s), .d(
        n3080), .sdi(n2160), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_20__19__slave ( .q(_RegFile_20__19), .qb(n2161), .d(
        _RegFile_reg_20__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_20__1__master ( .q(_RegFile_reg_20__1__m2s), .d(
        n3062), .sdi(n4208), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_20__1__slave ( .q(_RegFile_20__1), .qb(n4207), .d(
        _RegFile_reg_20__1__m2s), .g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_20__20__master ( .q(_RegFile_reg_20__20__m2s), .d(
        n3081), .sdi(n2161), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_20__20__slave ( .q(_RegFile_20__20), .qb(n2162), .d(
        _RegFile_reg_20__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_20__21__master ( .q(_RegFile_reg_20__21__m2s), .d(
        n3082), .sdi(n2162), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n964), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_20__21__slave ( .q(_RegFile_20__21), .qb(n2163), .d(
        _RegFile_reg_20__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n964), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_20__22__master ( .q(_RegFile_reg_20__22__m2s), .d(
        n3083), .sdi(n2163), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_20__22__slave ( .q(_RegFile_20__22), .qb(n2164), .d(
        _RegFile_reg_20__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_20__23__master ( .q(_RegFile_reg_20__23__m2s), .d(
        n3084), .sdi(n2164), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n964), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_20__23__slave ( .q(_RegFile_20__23), .qb(n2165), .d(
        _RegFile_reg_20__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n964), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_20__24__master ( .q(_RegFile_reg_20__24__m2s), .d(
        n3085), .sdi(n2165), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_20__24__slave ( .q(_RegFile_20__24), .qb(n2166), .d(
        _RegFile_reg_20__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_20__25__master ( .q(_RegFile_reg_20__25__m2s), .d(
        n3086), .sdi(n2166), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n964), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_20__25__slave ( .q(_RegFile_20__25), .qb(n2167), .d(
        _RegFile_reg_20__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n964), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_20__26__master ( .q(_RegFile_reg_20__26__m2s), .d(
        n3087), .sdi(n2167), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_20__26__slave ( .q(_RegFile_20__26), .qb(n2168), .d(
        _RegFile_reg_20__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_20__27__master ( .q(_RegFile_reg_20__27__m2s), .d(
        n3088), .sdi(n2168), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n964), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_20__27__slave ( .q(_RegFile_20__27), .qb(n2169), .d(
        _RegFile_reg_20__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n964), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_20__28__master ( .q(_RegFile_reg_20__28__m2s), .d(
        n3089), .sdi(n2169), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_20__28__slave ( .q(_RegFile_20__28), .qb(n2170), .d(
        _RegFile_reg_20__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_20__29__master ( .q(_RegFile_reg_20__29__m2s), .d(
        n3090), .sdi(n2170), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n964), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_20__29__slave ( .q(_RegFile_20__29), .qb(n2171), .d(
        _RegFile_reg_20__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n964), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_20__2__master ( .q(_RegFile_reg_20__2__m2s), .d(
        n3063), .sdi(n4207), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n963), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_20__2__slave ( .q(_RegFile_20__2), .qb(n4206), .d(
        _RegFile_reg_20__2__m2s), .g(Ctrl__Regs_1__en2), .rb(n963), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_20__30__master ( .q(_RegFile_reg_20__30__m2s), .d(
        n3091), .sdi(n2171), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n964), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_20__30__slave ( .q(_RegFile_20__30), .qb(n2172), .d(
        _RegFile_reg_20__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n964), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_20__31__master ( .q(_RegFile_reg_20__31__m2s), .d(
        n3092), .sdi(n2172), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_20__31__slave ( .q(_RegFile_20__31), .qb(n2173), .d(
        _RegFile_reg_20__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_20__3__master ( .q(_RegFile_reg_20__3__m2s), .d(
        n3064), .sdi(n4206), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_20__3__slave ( .q(_RegFile_20__3), .qb(n4205), .d(
        _RegFile_reg_20__3__m2s), .g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_20__4__master ( .q(_RegFile_reg_20__4__m2s), .d(
        n3065), .sdi(n4205), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n964), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_20__4__slave ( .q(_RegFile_20__4), .qb(n4204), .d(
        _RegFile_reg_20__4__m2s), .g(Ctrl__Regs_1__en2), .rb(n964), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_20__5__master ( .q(_RegFile_reg_20__5__m2s), .d(
        n3066), .sdi(n4204), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_20__5__slave ( .q(_RegFile_20__5), .qb(n4203), .d(
        _RegFile_reg_20__5__m2s), .g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_20__6__master ( .q(_RegFile_reg_20__6__m2s), .d(
        n3067), .sdi(n4203), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n964), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_20__6__slave ( .q(_RegFile_20__6), .qb(n4202), .d(
        _RegFile_reg_20__6__m2s), .g(Ctrl__Regs_1__en2), .rb(n964), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_20__7__master ( .q(_RegFile_reg_20__7__m2s), .d(
        n3068), .sdi(n4202), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n937), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_20__7__slave ( .q(_RegFile_20__7), .qb(n4201), .d(
        _RegFile_reg_20__7__m2s), .g(Ctrl__Regs_1__en2), .rb(n937), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_20__8__master ( .q(_RegFile_reg_20__8__m2s), .d(
        n3069), .sdi(n4201), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n964), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_20__8__slave ( .q(_RegFile_20__8), .qb(n2174), .d(
        _RegFile_reg_20__8__m2s), .g(Ctrl__Regs_1__en2), .rb(n964), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_20__9__master ( .q(_RegFile_reg_20__9__m2s), .d(
        n3070), .sdi(n2174), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n937), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_20__9__slave ( .q(_RegFile_20__9), .qb(n2175), .d(
        _RegFile_reg_20__9__m2s), .g(Ctrl__Regs_1__en2), .rb(n937), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_21__0__master ( .q(_RegFile_reg_21__0__m2s), .d(
        n3029), .sdi(n2173), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n964), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_21__0__slave ( .q(_RegFile_21__0), .qb(n4200), .d(
        _RegFile_reg_21__0__m2s), .g(Ctrl__Regs_1__en2), .rb(n964), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_21__10__master ( .q(_RegFile_reg_21__10__m2s), .d(
        n3039), .sdi(n2199), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n964), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_21__10__slave ( .q(_RegFile_21__10), .qb(n2176), .d(
        _RegFile_reg_21__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n964), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_21__11__master ( .q(_RegFile_reg_21__11__m2s), .d(
        n3040), .sdi(n2176), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n937), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_21__11__slave ( .q(_RegFile_21__11), .qb(n2177), .d(
        _RegFile_reg_21__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n937), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_21__12__master ( .q(_RegFile_reg_21__12__m2s), .d(
        n3041), .sdi(n2177), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n964), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_21__12__slave ( .q(_RegFile_21__12), .qb(n2178), .d(
        _RegFile_reg_21__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n964), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_21__13__master ( .q(_RegFile_reg_21__13__m2s), .d(
        n3042), .sdi(n2178), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n937), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_21__13__slave ( .q(_RegFile_21__13), .qb(n2179), .d(
        _RegFile_reg_21__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n937), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_21__14__master ( .q(_RegFile_reg_21__14__m2s), .d(
        n3043), .sdi(n2179), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n964), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_21__14__slave ( .q(_RegFile_21__14), .qb(n2180), .d(
        _RegFile_reg_21__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n964), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_21__15__master ( .q(_RegFile_reg_21__15__m2s), .d(
        n3044), .sdi(n2180), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n937), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_21__15__slave ( .q(_RegFile_21__15), .qb(n2181), .d(
        _RegFile_reg_21__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n937), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_21__16__master ( .q(_RegFile_reg_21__16__m2s), .d(
        n3045), .sdi(n2181), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n964), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_21__16__slave ( .q(_RegFile_21__16), .qb(n2182), .d(
        _RegFile_reg_21__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n964), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_21__17__master ( .q(_RegFile_reg_21__17__m2s), .d(
        n3046), .sdi(n2182), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n937), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_21__17__slave ( .q(_RegFile_21__17), .qb(n2183), .d(
        _RegFile_reg_21__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n937), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_21__18__master ( .q(_RegFile_reg_21__18__m2s), .d(
        n3047), .sdi(n2183), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n964), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_21__18__slave ( .q(_RegFile_21__18), .qb(n2184), .d(
        _RegFile_reg_21__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n964), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_21__19__master ( .q(_RegFile_reg_21__19__m2s), .d(
        n3048), .sdi(n2184), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n937), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_21__19__slave ( .q(_RegFile_21__19), .qb(n2185), .d(
        _RegFile_reg_21__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n937), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_21__1__master ( .q(_RegFile_reg_21__1__m2s), .d(
        n3030), .sdi(n4200), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n937), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_21__1__slave ( .q(_RegFile_21__1), .qb(n4199), .d(
        _RegFile_reg_21__1__m2s), .g(Ctrl__Regs_1__en2), .rb(n937), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_21__20__master ( .q(_RegFile_reg_21__20__m2s), .d(
        n3049), .sdi(n2185), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n937), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_21__20__slave ( .q(_RegFile_21__20), .qb(n2186), .d(
        _RegFile_reg_21__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n937), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_21__21__master ( .q(_RegFile_reg_21__21__m2s), .d(
        n3050), .sdi(n2186), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n965), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_21__21__slave ( .q(_RegFile_21__21), .qb(n2187), .d(
        _RegFile_reg_21__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n965), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_21__22__master ( .q(_RegFile_reg_21__22__m2s), .d(
        n3051), .sdi(n2187), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n937), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_21__22__slave ( .q(_RegFile_21__22), .qb(n2188), .d(
        _RegFile_reg_21__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n937), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_21__23__master ( .q(_RegFile_reg_21__23__m2s), .d(
        n3052), .sdi(n2188), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n965), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_21__23__slave ( .q(_RegFile_21__23), .qb(n2189), .d(
        _RegFile_reg_21__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n965), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_21__24__master ( .q(_RegFile_reg_21__24__m2s), .d(
        n3053), .sdi(n2189), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n937), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_21__24__slave ( .q(_RegFile_21__24), .qb(n2190), .d(
        _RegFile_reg_21__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n937), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_21__25__master ( .q(_RegFile_reg_21__25__m2s), .d(
        n3054), .sdi(n2190), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n965), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_21__25__slave ( .q(_RegFile_21__25), .qb(n2191), .d(
        _RegFile_reg_21__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n965), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_21__26__master ( .q(_RegFile_reg_21__26__m2s), .d(
        n3055), .sdi(n2191), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n937), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_21__26__slave ( .q(_RegFile_21__26), .qb(n2192), .d(
        _RegFile_reg_21__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n937), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_21__27__master ( .q(_RegFile_reg_21__27__m2s), .d(
        n3056), .sdi(n2192), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n965), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_21__27__slave ( .q(_RegFile_21__27), .qb(n2193), .d(
        _RegFile_reg_21__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n965), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_21__28__master ( .q(_RegFile_reg_21__28__m2s), .d(
        n3057), .sdi(n2193), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n937), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_21__28__slave ( .q(_RegFile_21__28), .qb(n2194), .d(
        _RegFile_reg_21__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n937), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_21__29__master ( .q(_RegFile_reg_21__29__m2s), .d(
        n3058), .sdi(n2194), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n965), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_21__29__slave ( .q(_RegFile_21__29), .qb(n2195), .d(
        _RegFile_reg_21__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n965), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_21__2__master ( .q(_RegFile_reg_21__2__m2s), .d(
        n3031), .sdi(n4199), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n965), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_21__2__slave ( .q(_RegFile_21__2), .qb(n4198), .d(
        _RegFile_reg_21__2__m2s), .g(Ctrl__Regs_1__en2), .rb(n965), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_21__30__master ( .q(_RegFile_reg_21__30__m2s), .d(
        n3059), .sdi(n2195), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n965), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_21__30__slave ( .q(_RegFile_21__30), .qb(n2196), .d(
        _RegFile_reg_21__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n965), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_21__31__master ( .q(_RegFile_reg_21__31__m2s), .d(
        n3060), .sdi(n2196), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n937), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_21__31__slave ( .q(_RegFile_21__31), .qb(n2197), .d(
        _RegFile_reg_21__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n937), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_21__3__master ( .q(_RegFile_reg_21__3__m2s), .d(
        n3032), .sdi(n4198), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n937), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_21__3__slave ( .q(_RegFile_21__3), .qb(n4197), .d(
        _RegFile_reg_21__3__m2s), .g(Ctrl__Regs_1__en2), .rb(n937), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_21__4__master ( .q(_RegFile_reg_21__4__m2s), .d(
        n3033), .sdi(n4197), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n965), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_21__4__slave ( .q(_RegFile_21__4), .qb(n4196), .d(
        _RegFile_reg_21__4__m2s), .g(Ctrl__Regs_1__en2), .rb(n965), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_21__5__master ( .q(_RegFile_reg_21__5__m2s), .d(
        n3034), .sdi(n4196), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n936), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_21__5__slave ( .q(_RegFile_21__5), .qb(n4195), .d(
        _RegFile_reg_21__5__m2s), .g(Ctrl__Regs_1__en2), .rb(n936), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_21__6__master ( .q(_RegFile_reg_21__6__m2s), .d(
        n3035), .sdi(n4195), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n965), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_21__6__slave ( .q(_RegFile_21__6), .qb(n4194), .d(
        _RegFile_reg_21__6__m2s), .g(Ctrl__Regs_1__en2), .rb(n965), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_21__7__master ( .q(_RegFile_reg_21__7__m2s), .d(
        n3036), .sdi(n4194), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n936), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_21__7__slave ( .q(_RegFile_21__7), .qb(n4193), .d(
        _RegFile_reg_21__7__m2s), .g(Ctrl__Regs_1__en2), .rb(n936), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_21__8__master ( .q(_RegFile_reg_21__8__m2s), .d(
        n3037), .sdi(n4193), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n965), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_21__8__slave ( .q(_RegFile_21__8), .qb(n2198), .d(
        _RegFile_reg_21__8__m2s), .g(Ctrl__Regs_1__en2), .rb(n965), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_21__9__master ( .q(_RegFile_reg_21__9__m2s), .d(
        n3038), .sdi(n2198), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n936), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_21__9__slave ( .q(_RegFile_21__9), .qb(n2199), .d(
        _RegFile_reg_21__9__m2s), .g(Ctrl__Regs_1__en2), .rb(n936), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_22__0__master ( .q(_RegFile_reg_22__0__m2s), .d(
        n2997), .sdi(n2197), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n965), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_22__0__slave ( .q(_RegFile_22__0), .qb(n4192), .d(
        _RegFile_reg_22__0__m2s), .g(Ctrl__Regs_1__en2), .rb(n965), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_22__10__master ( .q(_RegFile_reg_22__10__m2s), .d(
        n3007), .sdi(n2223), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n965), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_22__10__slave ( .q(_RegFile_22__10), .qb(n2200), .d(
        _RegFile_reg_22__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n965), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_22__11__master ( .q(_RegFile_reg_22__11__m2s), .d(
        n3008), .sdi(n2200), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n936), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_22__11__slave ( .q(_RegFile_22__11), .qb(n2201), .d(
        _RegFile_reg_22__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n936), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_22__12__master ( .q(_RegFile_reg_22__12__m2s), .d(
        n3009), .sdi(n2201), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n965), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_22__12__slave ( .q(_RegFile_22__12), .qb(n2202), .d(
        _RegFile_reg_22__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n965), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_22__13__master ( .q(_RegFile_reg_22__13__m2s), .d(
        n3010), .sdi(n2202), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n936), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_22__13__slave ( .q(_RegFile_22__13), .qb(n2203), .d(
        _RegFile_reg_22__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n936), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_22__14__master ( .q(_RegFile_reg_22__14__m2s), .d(
        n3011), .sdi(n2203), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n965), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_22__14__slave ( .q(_RegFile_22__14), .qb(n2204), .d(
        _RegFile_reg_22__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n965), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_22__15__master ( .q(_RegFile_reg_22__15__m2s), .d(
        n3012), .sdi(n2204), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n936), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_22__15__slave ( .q(_RegFile_22__15), .qb(n2205), .d(
        _RegFile_reg_22__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n936), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_22__16__master ( .q(_RegFile_reg_22__16__m2s), .d(
        n3013), .sdi(n2205), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n965), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_22__16__slave ( .q(_RegFile_22__16), .qb(n2206), .d(
        _RegFile_reg_22__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n965), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_22__17__master ( .q(_RegFile_reg_22__17__m2s), .d(
        n3014), .sdi(n2206), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n936), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_22__17__slave ( .q(_RegFile_22__17), .qb(n2207), .d(
        _RegFile_reg_22__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n936), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_22__18__master ( .q(_RegFile_reg_22__18__m2s), .d(
        n3015), .sdi(n2207), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_22__18__slave ( .q(_RegFile_22__18), .qb(n2208), .d(
        _RegFile_reg_22__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_22__19__master ( .q(_RegFile_reg_22__19__m2s), .d(
        n3016), .sdi(n2208), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n936), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_22__19__slave ( .q(_RegFile_22__19), .qb(n2209), .d(
        _RegFile_reg_22__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n936), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_22__1__master ( .q(_RegFile_reg_22__1__m2s), .d(
        n2998), .sdi(n4192), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n936), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_22__1__slave ( .q(_RegFile_22__1), .qb(n4191), .d(
        _RegFile_reg_22__1__m2s), .g(Ctrl__Regs_1__en2), .rb(n936), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_22__20__master ( .q(_RegFile_reg_22__20__m2s), .d(
        n3017), .sdi(n2209), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n936), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_22__20__slave ( .q(_RegFile_22__20), .qb(n2210), .d(
        _RegFile_reg_22__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n936), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_22__21__master ( .q(_RegFile_reg_22__21__m2s), .d(
        n3018), .sdi(n2210), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_22__21__slave ( .q(_RegFile_22__21), .qb(n2211), .d(
        _RegFile_reg_22__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_22__22__master ( .q(_RegFile_reg_22__22__m2s), .d(
        n3019), .sdi(n2211), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n936), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_22__22__slave ( .q(_RegFile_22__22), .qb(n2212), .d(
        _RegFile_reg_22__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n936), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_22__23__master ( .q(_RegFile_reg_22__23__m2s), .d(
        n3020), .sdi(n2212), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_22__23__slave ( .q(_RegFile_22__23), .qb(n2213), .d(
        _RegFile_reg_22__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_22__24__master ( .q(_RegFile_reg_22__24__m2s), .d(
        n3021), .sdi(n2213), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n936), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_22__24__slave ( .q(_RegFile_22__24), .qb(n2214), .d(
        _RegFile_reg_22__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n936), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_22__25__master ( .q(_RegFile_reg_22__25__m2s), .d(
        n3022), .sdi(n2214), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_22__25__slave ( .q(_RegFile_22__25), .qb(n2215), .d(
        _RegFile_reg_22__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_22__26__master ( .q(_RegFile_reg_22__26__m2s), .d(
        n3023), .sdi(n2215), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n936), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_22__26__slave ( .q(_RegFile_22__26), .qb(n2216), .d(
        _RegFile_reg_22__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n936), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_22__27__master ( .q(_RegFile_reg_22__27__m2s), .d(
        n3024), .sdi(n2216), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_22__27__slave ( .q(_RegFile_22__27), .qb(n2217), .d(
        _RegFile_reg_22__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_22__28__master ( .q(_RegFile_reg_22__28__m2s), .d(
        n3025), .sdi(n2217), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n936), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_22__28__slave ( .q(_RegFile_22__28), .qb(n2218), .d(
        _RegFile_reg_22__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n936), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_22__29__master ( .q(_RegFile_reg_22__29__m2s), .d(
        n3026), .sdi(n2218), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_22__29__slave ( .q(_RegFile_22__29), .qb(n2219), .d(
        _RegFile_reg_22__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_22__2__master ( .q(_RegFile_reg_22__2__m2s), .d(
        n2999), .sdi(n4191), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_22__2__slave ( .q(_RegFile_22__2), .qb(n4190), .d(
        _RegFile_reg_22__2__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_22__30__master ( .q(_RegFile_reg_22__30__m2s), .d(
        n3027), .sdi(n2219), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_22__30__slave ( .q(_RegFile_22__30), .qb(n2220), .d(
        _RegFile_reg_22__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_22__31__master ( .q(_RegFile_reg_22__31__m2s), .d(
        n3028), .sdi(n2220), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_22__31__slave ( .q(_RegFile_22__31), .qb(n2221), .d(
        _RegFile_reg_22__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_22__3__master ( .q(_RegFile_reg_22__3__m2s), .d(
        n3000), .sdi(n4190), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n936), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_22__3__slave ( .q(_RegFile_22__3), .qb(n4189), .d(
        _RegFile_reg_22__3__m2s), .g(Ctrl__Regs_1__en2), .rb(n936), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_22__4__master ( .q(_RegFile_reg_22__4__m2s), .d(
        n3001), .sdi(n4189), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_22__4__slave ( .q(_RegFile_22__4), .qb(n4188), .d(
        _RegFile_reg_22__4__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_22__5__master ( .q(_RegFile_reg_22__5__m2s), .d(
        n3002), .sdi(n4188), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_22__5__slave ( .q(_RegFile_22__5), .qb(n4187), .d(
        _RegFile_reg_22__5__m2s), .g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_22__6__master ( .q(_RegFile_reg_22__6__m2s), .d(
        n3003), .sdi(n4187), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_22__6__slave ( .q(_RegFile_22__6), .qb(n4186), .d(
        _RegFile_reg_22__6__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_22__7__master ( .q(_RegFile_reg_22__7__m2s), .d(
        n3004), .sdi(n4186), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_22__7__slave ( .q(_RegFile_22__7), .qb(n4185), .d(
        _RegFile_reg_22__7__m2s), .g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_22__8__master ( .q(_RegFile_reg_22__8__m2s), .d(
        n3005), .sdi(n4185), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_22__8__slave ( .q(_RegFile_22__8), .qb(n2222), .d(
        _RegFile_reg_22__8__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_22__9__master ( .q(_RegFile_reg_22__9__m2s), .d(
        n3006), .sdi(n2222), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_22__9__slave ( .q(_RegFile_22__9), .qb(n2223), .d(
        _RegFile_reg_22__9__m2s), .g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_23__0__master ( .q(_RegFile_reg_23__0__m2s), .d(
        n2965), .sdi(n2221), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_23__0__slave ( .q(_RegFile_23__0), .qb(n4184), .d(
        _RegFile_reg_23__0__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_23__10__master ( .q(_RegFile_reg_23__10__m2s), .d(
        n2975), .sdi(n2247), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_23__10__slave ( .q(_RegFile_23__10), .qb(n2224), .d(
        _RegFile_reg_23__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_23__11__master ( .q(_RegFile_reg_23__11__m2s), .d(
        n2976), .sdi(n2224), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_23__11__slave ( .q(_RegFile_23__11), .qb(n2225), .d(
        _RegFile_reg_23__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_23__12__master ( .q(_RegFile_reg_23__12__m2s), .d(
        n2977), .sdi(n2225), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_23__12__slave ( .q(_RegFile_23__12), .qb(n2226), .d(
        _RegFile_reg_23__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_23__13__master ( .q(_RegFile_reg_23__13__m2s), .d(
        n2978), .sdi(n2226), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_23__13__slave ( .q(_RegFile_23__13), .qb(n2227), .d(
        _RegFile_reg_23__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_23__14__master ( .q(_RegFile_reg_23__14__m2s), .d(
        n2979), .sdi(n2227), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_23__14__slave ( .q(_RegFile_23__14), .qb(n2228), .d(
        _RegFile_reg_23__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_23__15__master ( .q(_RegFile_reg_23__15__m2s), .d(
        n2980), .sdi(n2228), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_23__15__slave ( .q(_RegFile_23__15), .qb(n2229), .d(
        _RegFile_reg_23__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_23__16__master ( .q(_RegFile_reg_23__16__m2s), .d(
        n2981), .sdi(n2229), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_23__16__slave ( .q(_RegFile_23__16), .qb(n2230), .d(
        _RegFile_reg_23__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_23__17__master ( .q(_RegFile_reg_23__17__m2s), .d(
        n2982), .sdi(n2230), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_23__17__slave ( .q(_RegFile_23__17), .qb(n2231), .d(
        _RegFile_reg_23__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_23__18__master ( .q(_RegFile_reg_23__18__m2s), .d(
        n2983), .sdi(n2231), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_23__18__slave ( .q(_RegFile_23__18), .qb(n2232), .d(
        _RegFile_reg_23__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_23__19__master ( .q(_RegFile_reg_23__19__m2s), .d(
        n2984), .sdi(n2232), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_23__19__slave ( .q(_RegFile_23__19), .qb(n2233), .d(
        _RegFile_reg_23__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_23__1__master ( .q(_RegFile_reg_23__1__m2s), .d(
        n2966), .sdi(n4184), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_23__1__slave ( .q(_RegFile_23__1), .qb(n4183), .d(
        _RegFile_reg_23__1__m2s), .g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_23__20__master ( .q(_RegFile_reg_23__20__m2s), .d(
        n2985), .sdi(n2233), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_23__20__slave ( .q(_RegFile_23__20), .qb(n2234), .d(
        _RegFile_reg_23__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_23__21__master ( .q(_RegFile_reg_23__21__m2s), .d(
        n2986), .sdi(n2234), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_23__21__slave ( .q(_RegFile_23__21), .qb(n2235), .d(
        _RegFile_reg_23__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_23__22__master ( .q(_RegFile_reg_23__22__m2s), .d(
        n2987), .sdi(n2235), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_23__22__slave ( .q(_RegFile_23__22), .qb(n2236), .d(
        _RegFile_reg_23__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_23__23__master ( .q(_RegFile_reg_23__23__m2s), .d(
        n2988), .sdi(n2236), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_23__23__slave ( .q(_RegFile_23__23), .qb(n2237), .d(
        _RegFile_reg_23__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_23__24__master ( .q(_RegFile_reg_23__24__m2s), .d(
        n2989), .sdi(n2237), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_23__24__slave ( .q(_RegFile_23__24), .qb(n2238), .d(
        _RegFile_reg_23__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_23__25__master ( .q(_RegFile_reg_23__25__m2s), .d(
        n2990), .sdi(n2238), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_23__25__slave ( .q(_RegFile_23__25), .qb(n2239), .d(
        _RegFile_reg_23__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_23__26__master ( .q(_RegFile_reg_23__26__m2s), .d(
        n2991), .sdi(n2239), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_23__26__slave ( .q(_RegFile_23__26), .qb(n2240), .d(
        _RegFile_reg_23__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_23__27__master ( .q(_RegFile_reg_23__27__m2s), .d(
        n2992), .sdi(n2240), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_23__27__slave ( .q(_RegFile_23__27), .qb(n2241), .d(
        _RegFile_reg_23__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_23__28__master ( .q(_RegFile_reg_23__28__m2s), .d(
        n2993), .sdi(n2241), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_23__28__slave ( .q(_RegFile_23__28), .qb(n2242), .d(
        _RegFile_reg_23__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_23__29__master ( .q(_RegFile_reg_23__29__m2s), .d(
        n2994), .sdi(n2242), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_23__29__slave ( .q(_RegFile_23__29), .qb(n2243), .d(
        _RegFile_reg_23__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_23__2__master ( .q(_RegFile_reg_23__2__m2s), .d(
        n2967), .sdi(n4183), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_23__2__slave ( .q(_RegFile_23__2), .qb(n4182), .d(
        _RegFile_reg_23__2__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_23__30__master ( .q(_RegFile_reg_23__30__m2s), .d(
        n2995), .sdi(n2243), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_23__30__slave ( .q(_RegFile_23__30), .qb(n2244), .d(
        _RegFile_reg_23__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_23__31__master ( .q(_RegFile_reg_23__31__m2s), .d(
        n2996), .sdi(n2244), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n935), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_23__31__slave ( .q(_RegFile_23__31), .qb(n2245), .d(
        _RegFile_reg_23__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n935), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_23__3__master ( .q(_RegFile_reg_23__3__m2s), .d(
        n2968), .sdi(n4182), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n935), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_23__3__slave ( .q(_RegFile_23__3), .qb(n4181), .d(
        _RegFile_reg_23__3__m2s), .g(Ctrl__Regs_1__en2), .rb(n935), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_23__4__master ( .q(_RegFile_reg_23__4__m2s), .d(
        n2969), .sdi(n4181), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_23__4__slave ( .q(_RegFile_23__4), .qb(n4180), .d(
        _RegFile_reg_23__4__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_23__5__master ( .q(_RegFile_reg_23__5__m2s), .d(
        n2970), .sdi(n4180), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n935), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_23__5__slave ( .q(_RegFile_23__5), .qb(n4179), .d(
        _RegFile_reg_23__5__m2s), .g(Ctrl__Regs_1__en2), .rb(n935), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_23__6__master ( .q(_RegFile_reg_23__6__m2s), .d(
        n2971), .sdi(n4179), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_23__6__slave ( .q(_RegFile_23__6), .qb(n4178), .d(
        _RegFile_reg_23__6__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_23__7__master ( .q(_RegFile_reg_23__7__m2s), .d(
        n2972), .sdi(n4178), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n935), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_23__7__slave ( .q(_RegFile_23__7), .qb(n4177), .d(
        _RegFile_reg_23__7__m2s), .g(Ctrl__Regs_1__en2), .rb(n935), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_23__8__master ( .q(_RegFile_reg_23__8__m2s), .d(
        n2973), .sdi(n4177), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_23__8__slave ( .q(_RegFile_23__8), .qb(n2246), .d(
        _RegFile_reg_23__8__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_23__9__master ( .q(_RegFile_reg_23__9__m2s), .d(
        n2974), .sdi(n2246), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n935), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_23__9__slave ( .q(_RegFile_23__9), .qb(n2247), .d(
        _RegFile_reg_23__9__m2s), .g(Ctrl__Regs_1__en2), .rb(n935), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_24__0__master ( .q(_RegFile_reg_24__0__m2s), .d(
        n2933), .sdi(n2245), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_24__0__slave ( .q(_RegFile_24__0), .qb(n4176), .d(
        _RegFile_reg_24__0__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_24__10__master ( .q(_RegFile_reg_24__10__m2s), .d(
        n2943), .sdi(n2271), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_24__10__slave ( .q(_RegFile_24__10), .qb(n2248), .d(
        _RegFile_reg_24__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_24__11__master ( .q(_RegFile_reg_24__11__m2s), .d(
        n2944), .sdi(n2248), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n935), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_24__11__slave ( .q(_RegFile_24__11), .qb(n2249), .d(
        _RegFile_reg_24__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n935), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_24__12__master ( .q(_RegFile_reg_24__12__m2s), .d(
        n2945), .sdi(n2249), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_24__12__slave ( .q(_RegFile_24__12), .qb(n2250), .d(
        _RegFile_reg_24__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_24__13__master ( .q(_RegFile_reg_24__13__m2s), .d(
        n2946), .sdi(n2250), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n935), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_24__13__slave ( .q(_RegFile_24__13), .qb(n2251), .d(
        _RegFile_reg_24__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n935), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_24__14__master ( .q(_RegFile_reg_24__14__m2s), .d(
        n2947), .sdi(n2251), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_24__14__slave ( .q(_RegFile_24__14), .qb(n2252), .d(
        _RegFile_reg_24__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_24__15__master ( .q(_RegFile_reg_24__15__m2s), .d(
        n2948), .sdi(n2252), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n935), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_24__15__slave ( .q(_RegFile_24__15), .qb(n2253), .d(
        _RegFile_reg_24__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n935), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_24__16__master ( .q(_RegFile_reg_24__16__m2s), .d(
        n2949), .sdi(n2253), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_24__16__slave ( .q(_RegFile_24__16), .qb(n2254), .d(
        _RegFile_reg_24__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_24__17__master ( .q(_RegFile_reg_24__17__m2s), .d(
        n2950), .sdi(n2254), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n935), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_24__17__slave ( .q(_RegFile_24__17), .qb(n2255), .d(
        _RegFile_reg_24__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n935), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_24__18__master ( .q(_RegFile_reg_24__18__m2s), .d(
        n2951), .sdi(n2255), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_24__18__slave ( .q(_RegFile_24__18), .qb(n2256), .d(
        _RegFile_reg_24__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_24__19__master ( .q(_RegFile_reg_24__19__m2s), .d(
        n2952), .sdi(n2256), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n935), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_24__19__slave ( .q(_RegFile_24__19), .qb(n2257), .d(
        _RegFile_reg_24__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n935), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_24__1__master ( .q(_RegFile_reg_24__1__m2s), .d(
        n2934), .sdi(n4176), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n935), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_24__1__slave ( .q(_RegFile_24__1), .qb(n4175), .d(
        _RegFile_reg_24__1__m2s), .g(Ctrl__Regs_1__en2), .rb(n935), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_24__20__master ( .q(_RegFile_reg_24__20__m2s), .d(
        n2953), .sdi(n2257), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n935), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_24__20__slave ( .q(_RegFile_24__20), .qb(n2258), .d(
        _RegFile_reg_24__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n935), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_24__21__master ( .q(_RegFile_reg_24__21__m2s), .d(
        n2954), .sdi(n2258), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_24__21__slave ( .q(_RegFile_24__21), .qb(n2259), .d(
        _RegFile_reg_24__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_24__22__master ( .q(_RegFile_reg_24__22__m2s), .d(
        n2955), .sdi(n2259), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n935), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_24__22__slave ( .q(_RegFile_24__22), .qb(n2260), .d(
        _RegFile_reg_24__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n935), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_24__23__master ( .q(_RegFile_reg_24__23__m2s), .d(
        n2956), .sdi(n2260), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_24__23__slave ( .q(_RegFile_24__23), .qb(n2261), .d(
        _RegFile_reg_24__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_24__24__master ( .q(_RegFile_reg_24__24__m2s), .d(
        n2957), .sdi(n2261), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n935), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_24__24__slave ( .q(_RegFile_24__24), .qb(n2262), .d(
        _RegFile_reg_24__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n935), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_24__25__master ( .q(_RegFile_reg_24__25__m2s), .d(
        n2958), .sdi(n2262), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_24__25__slave ( .q(_RegFile_24__25), .qb(n2263), .d(
        _RegFile_reg_24__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_24__26__master ( .q(_RegFile_reg_24__26__m2s), .d(
        n2959), .sdi(n2263), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n935), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_24__26__slave ( .q(_RegFile_24__26), .qb(n2264), .d(
        _RegFile_reg_24__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n935), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_24__27__master ( .q(_RegFile_reg_24__27__m2s), .d(
        n2960), .sdi(n2264), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_24__27__slave ( .q(_RegFile_24__27), .qb(n2265), .d(
        _RegFile_reg_24__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_24__28__master ( .q(_RegFile_reg_24__28__m2s), .d(
        n2961), .sdi(n2265), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_24__28__slave ( .q(_RegFile_24__28), .qb(n2266), .d(
        _RegFile_reg_24__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_24__29__master ( .q(_RegFile_reg_24__29__m2s), .d(
        n2962), .sdi(n2266), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_24__29__slave ( .q(_RegFile_24__29), .qb(n2267), .d(
        _RegFile_reg_24__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_24__2__master ( .q(_RegFile_reg_24__2__m2s), .d(
        n2935), .sdi(n4175), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_24__2__slave ( .q(_RegFile_24__2), .qb(n4174), .d(
        _RegFile_reg_24__2__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_24__30__master ( .q(_RegFile_reg_24__30__m2s), .d(
        n2963), .sdi(n2267), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_24__30__slave ( .q(_RegFile_24__30), .qb(n2268), .d(
        _RegFile_reg_24__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_24__31__master ( .q(_RegFile_reg_24__31__m2s), .d(
        n2964), .sdi(n2268), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_24__31__slave ( .q(_RegFile_24__31), .qb(n2269), .d(
        _RegFile_reg_24__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_24__3__master ( .q(_RegFile_reg_24__3__m2s), .d(
        n2936), .sdi(n4174), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_24__3__slave ( .q(_RegFile_24__3), .qb(n4173), .d(
        _RegFile_reg_24__3__m2s), .g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_24__4__master ( .q(_RegFile_reg_24__4__m2s), .d(
        n2937), .sdi(n4173), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_24__4__slave ( .q(_RegFile_24__4), .qb(n4172), .d(
        _RegFile_reg_24__4__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_24__5__master ( .q(_RegFile_reg_24__5__m2s), .d(
        n2938), .sdi(n4172), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_24__5__slave ( .q(_RegFile_24__5), .qb(n4171), .d(
        _RegFile_reg_24__5__m2s), .g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_24__6__master ( .q(_RegFile_reg_24__6__m2s), .d(
        n2939), .sdi(n4171), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_24__6__slave ( .q(_RegFile_24__6), .qb(n4170), .d(
        _RegFile_reg_24__6__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_24__7__master ( .q(_RegFile_reg_24__7__m2s), .d(
        n2940), .sdi(n4170), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_24__7__slave ( .q(_RegFile_24__7), .qb(n4169), .d(
        _RegFile_reg_24__7__m2s), .g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_24__8__master ( .q(_RegFile_reg_24__8__m2s), .d(
        n2941), .sdi(n4169), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_24__8__slave ( .q(_RegFile_24__8), .qb(n2270), .d(
        _RegFile_reg_24__8__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_24__9__master ( .q(_RegFile_reg_24__9__m2s), .d(
        n2942), .sdi(n2270), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_24__9__slave ( .q(_RegFile_24__9), .qb(n2271), .d(
        _RegFile_reg_24__9__m2s), .g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_25__0__master ( .q(_RegFile_reg_25__0__m2s), .d(
        n2901), .sdi(n2269), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_25__0__slave ( .q(_RegFile_25__0), .qb(n4168), .d(
        _RegFile_reg_25__0__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_25__10__master ( .q(_RegFile_reg_25__10__m2s), .d(
        n2911), .sdi(n2295), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_25__10__slave ( .q(_RegFile_25__10), .qb(n2272), .d(
        _RegFile_reg_25__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_25__11__master ( .q(_RegFile_reg_25__11__m2s), .d(
        n2912), .sdi(n2272), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_25__11__slave ( .q(_RegFile_25__11), .qb(n2273), .d(
        _RegFile_reg_25__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_25__12__master ( .q(_RegFile_reg_25__12__m2s), .d(
        n2913), .sdi(n2273), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_25__12__slave ( .q(_RegFile_25__12), .qb(n2274), .d(
        _RegFile_reg_25__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_25__13__master ( .q(_RegFile_reg_25__13__m2s), .d(
        n2914), .sdi(n2274), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_25__13__slave ( .q(_RegFile_25__13), .qb(n2275), .d(
        _RegFile_reg_25__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_25__14__master ( .q(_RegFile_reg_25__14__m2s), .d(
        n2915), .sdi(n2275), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_25__14__slave ( .q(_RegFile_25__14), .qb(n2276), .d(
        _RegFile_reg_25__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_25__15__master ( .q(_RegFile_reg_25__15__m2s), .d(
        n2916), .sdi(n2276), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_25__15__slave ( .q(_RegFile_25__15), .qb(n2277), .d(
        _RegFile_reg_25__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_25__16__master ( .q(_RegFile_reg_25__16__m2s), .d(
        n2917), .sdi(n2277), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_25__16__slave ( .q(_RegFile_25__16), .qb(n2278), .d(
        _RegFile_reg_25__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_25__17__master ( .q(_RegFile_reg_25__17__m2s), .d(
        n2918), .sdi(n2278), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_25__17__slave ( .q(_RegFile_25__17), .qb(n2279), .d(
        _RegFile_reg_25__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_25__18__master ( .q(_RegFile_reg_25__18__m2s), .d(
        n2919), .sdi(n2279), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_25__18__slave ( .q(_RegFile_25__18), .qb(n2280), .d(
        _RegFile_reg_25__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_25__19__master ( .q(_RegFile_reg_25__19__m2s), .d(
        n2920), .sdi(n2280), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_25__19__slave ( .q(_RegFile_25__19), .qb(n2281), .d(
        _RegFile_reg_25__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_25__1__master ( .q(_RegFile_reg_25__1__m2s), .d(
        n2902), .sdi(n4168), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_25__1__slave ( .q(_RegFile_25__1), .qb(n4167), .d(
        _RegFile_reg_25__1__m2s), .g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_25__20__master ( .q(_RegFile_reg_25__20__m2s), .d(
        n2921), .sdi(n2281), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_25__20__slave ( .q(_RegFile_25__20), .qb(n2282), .d(
        _RegFile_reg_25__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_25__21__master ( .q(_RegFile_reg_25__21__m2s), .d(
        n2922), .sdi(n2282), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_25__21__slave ( .q(_RegFile_25__21), .qb(n2283), .d(
        _RegFile_reg_25__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_25__22__master ( .q(_RegFile_reg_25__22__m2s), .d(
        n2923), .sdi(n2283), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_25__22__slave ( .q(_RegFile_25__22), .qb(n2284), .d(
        _RegFile_reg_25__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_25__23__master ( .q(_RegFile_reg_25__23__m2s), .d(
        n2924), .sdi(n2284), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_25__23__slave ( .q(_RegFile_25__23), .qb(n2285), .d(
        _RegFile_reg_25__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_25__24__master ( .q(_RegFile_reg_25__24__m2s), .d(
        n2925), .sdi(n2285), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_25__24__slave ( .q(_RegFile_25__24), .qb(n2286), .d(
        _RegFile_reg_25__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_25__25__master ( .q(_RegFile_reg_25__25__m2s), .d(
        n2926), .sdi(n2286), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_25__25__slave ( .q(_RegFile_25__25), .qb(n2287), .d(
        _RegFile_reg_25__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_25__26__master ( .q(_RegFile_reg_25__26__m2s), .d(
        n2927), .sdi(n2287), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n934), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_25__26__slave ( .q(_RegFile_25__26), .qb(n2288), .d(
        _RegFile_reg_25__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n934), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_25__27__master ( .q(_RegFile_reg_25__27__m2s), .d(
        n2928), .sdi(n2288), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_25__27__slave ( .q(_RegFile_25__27), .qb(n2289), .d(
        _RegFile_reg_25__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_25__28__master ( .q(_RegFile_reg_25__28__m2s), .d(
        n2929), .sdi(n2289), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n934), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_25__28__slave ( .q(_RegFile_25__28), .qb(n2290), .d(
        _RegFile_reg_25__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n934), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_25__29__master ( .q(_RegFile_reg_25__29__m2s), .d(
        n2930), .sdi(n2290), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_25__29__slave ( .q(_RegFile_25__29), .qb(n2291), .d(
        _RegFile_reg_25__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_25__2__master ( .q(_RegFile_reg_25__2__m2s), .d(
        n2903), .sdi(n4167), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_25__2__slave ( .q(_RegFile_25__2), .qb(n4166), .d(
        _RegFile_reg_25__2__m2s), .g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_25__30__master ( .q(_RegFile_reg_25__30__m2s), .d(
        n2931), .sdi(n2291), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_25__30__slave ( .q(_RegFile_25__30), .qb(n2292), .d(
        _RegFile_reg_25__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_25__31__master ( .q(_RegFile_reg_25__31__m2s), .d(
        n2932), .sdi(n2292), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n934), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_25__31__slave ( .q(_RegFile_25__31), .qb(n2293), .d(
        _RegFile_reg_25__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n934), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_25__3__master ( .q(_RegFile_reg_25__3__m2s), .d(
        n2904), .sdi(n4166), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n934), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_25__3__slave ( .q(_RegFile_25__3), .qb(n4165), .d(
        _RegFile_reg_25__3__m2s), .g(Ctrl__Regs_1__en2), .rb(n934), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_25__4__master ( .q(_RegFile_reg_25__4__m2s), .d(
        n2905), .sdi(n4165), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_25__4__slave ( .q(_RegFile_25__4), .qb(n4164), .d(
        _RegFile_reg_25__4__m2s), .g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_25__5__master ( .q(_RegFile_reg_25__5__m2s), .d(
        n2906), .sdi(n4164), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n934), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_25__5__slave ( .q(_RegFile_25__5), .qb(n4163), .d(
        _RegFile_reg_25__5__m2s), .g(Ctrl__Regs_1__en2), .rb(n934), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_25__6__master ( .q(_RegFile_reg_25__6__m2s), .d(
        n2907), .sdi(n4163), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_25__6__slave ( .q(_RegFile_25__6), .qb(n4162), .d(
        _RegFile_reg_25__6__m2s), .g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_25__7__master ( .q(_RegFile_reg_25__7__m2s), .d(
        n2908), .sdi(n4162), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n934), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_25__7__slave ( .q(_RegFile_25__7), .qb(n4161), .d(
        _RegFile_reg_25__7__m2s), .g(Ctrl__Regs_1__en2), .rb(n934), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_25__8__master ( .q(_RegFile_reg_25__8__m2s), .d(
        n2909), .sdi(n4161), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_25__8__slave ( .q(_RegFile_25__8), .qb(n2294), .d(
        _RegFile_reg_25__8__m2s), .g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_25__9__master ( .q(_RegFile_reg_25__9__m2s), .d(
        n2910), .sdi(n2294), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n934), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_25__9__slave ( .q(_RegFile_25__9), .qb(n2295), .d(
        _RegFile_reg_25__9__m2s), .g(Ctrl__Regs_1__en2), .rb(n934), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_26__0__master ( .q(_RegFile_reg_26__0__m2s), .d(
        n2869), .sdi(n2293), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_26__0__slave ( .q(_RegFile_26__0), .qb(n4160), .d(
        _RegFile_reg_26__0__m2s), .g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_26__10__master ( .q(_RegFile_reg_26__10__m2s), .d(
        n2879), .sdi(n2319), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n970), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_26__10__slave ( .q(_RegFile_26__10), .qb(n2296), .d(
        _RegFile_reg_26__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n970), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_26__11__master ( .q(_RegFile_reg_26__11__m2s), .d(
        n2880), .sdi(n2296), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n934), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_26__11__slave ( .q(_RegFile_26__11), .qb(n2297), .d(
        _RegFile_reg_26__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n934), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_26__12__master ( .q(_RegFile_reg_26__12__m2s), .d(
        n2881), .sdi(n2297), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n970), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_26__12__slave ( .q(_RegFile_26__12), .qb(n2298), .d(
        _RegFile_reg_26__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n970), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_26__13__master ( .q(_RegFile_reg_26__13__m2s), .d(
        n2882), .sdi(n2298), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n934), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_26__13__slave ( .q(_RegFile_26__13), .qb(n2299), .d(
        _RegFile_reg_26__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n934), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_26__14__master ( .q(_RegFile_reg_26__14__m2s), .d(
        n2883), .sdi(n2299), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n970), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_26__14__slave ( .q(_RegFile_26__14), .qb(n2300), .d(
        _RegFile_reg_26__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n970), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_26__15__master ( .q(_RegFile_reg_26__15__m2s), .d(
        n2884), .sdi(n2300), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n934), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_26__15__slave ( .q(_RegFile_26__15), .qb(n2301), .d(
        _RegFile_reg_26__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n934), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_26__16__master ( .q(_RegFile_reg_26__16__m2s), .d(
        n2885), .sdi(n2301), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n970), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_26__16__slave ( .q(_RegFile_26__16), .qb(n2302), .d(
        _RegFile_reg_26__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n970), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_26__17__master ( .q(_RegFile_reg_26__17__m2s), .d(
        n2886), .sdi(n2302), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n934), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_26__17__slave ( .q(_RegFile_26__17), .qb(n2303), .d(
        _RegFile_reg_26__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n934), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_26__18__master ( .q(_RegFile_reg_26__18__m2s), .d(
        n2887), .sdi(n2303), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n970), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_26__18__slave ( .q(_RegFile_26__18), .qb(n2304), .d(
        _RegFile_reg_26__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n970), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_26__19__master ( .q(_RegFile_reg_26__19__m2s), .d(
        n2888), .sdi(n2304), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n934), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_26__19__slave ( .q(_RegFile_26__19), .qb(n2305), .d(
        _RegFile_reg_26__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n934), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_26__1__master ( .q(_RegFile_reg_26__1__m2s), .d(
        n2870), .sdi(n4160), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n934), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_26__1__slave ( .q(_RegFile_26__1), .qb(n4159), .d(
        _RegFile_reg_26__1__m2s), .g(Ctrl__Regs_1__en2), .rb(n934), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_26__20__master ( .q(_RegFile_reg_26__20__m2s), .d(
        n2889), .sdi(n2305), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n934), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_26__20__slave ( .q(_RegFile_26__20), .qb(n2306), .d(
        _RegFile_reg_26__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n934), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_26__21__master ( .q(_RegFile_reg_26__21__m2s), .d(
        n2890), .sdi(n2306), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n970), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_26__21__slave ( .q(_RegFile_26__21), .qb(n2307), .d(
        _RegFile_reg_26__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n970), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_26__22__master ( .q(_RegFile_reg_26__22__m2s), .d(
        n2891), .sdi(n2307), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n934), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_26__22__slave ( .q(_RegFile_26__22), .qb(n2308), .d(
        _RegFile_reg_26__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n934), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_26__23__master ( .q(_RegFile_reg_26__23__m2s), .d(
        n2892), .sdi(n2308), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n970), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_26__23__slave ( .q(_RegFile_26__23), .qb(n2309), .d(
        _RegFile_reg_26__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n970), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_26__24__master ( .q(_RegFile_reg_26__24__m2s), .d(
        n2893), .sdi(n2309), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n933), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_26__24__slave ( .q(_RegFile_26__24), .qb(n2310), .d(
        _RegFile_reg_26__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n933), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_26__25__master ( .q(_RegFile_reg_26__25__m2s), .d(
        n2894), .sdi(n2310), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n970), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_26__25__slave ( .q(_RegFile_26__25), .qb(n2311), .d(
        _RegFile_reg_26__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n970), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_26__26__master ( .q(_RegFile_reg_26__26__m2s), .d(
        n2895), .sdi(n2311), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n933), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_26__26__slave ( .q(_RegFile_26__26), .qb(n2312), .d(
        _RegFile_reg_26__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n933), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_26__27__master ( .q(_RegFile_reg_26__27__m2s), .d(
        n2896), .sdi(n2312), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n970), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_26__27__slave ( .q(_RegFile_26__27), .qb(n2313), .d(
        _RegFile_reg_26__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n970), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_26__28__master ( .q(_RegFile_reg_26__28__m2s), .d(
        n2897), .sdi(n2313), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n933), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_26__28__slave ( .q(_RegFile_26__28), .qb(n2314), .d(
        _RegFile_reg_26__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n933), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_26__29__master ( .q(_RegFile_reg_26__29__m2s), .d(
        n2898), .sdi(n2314), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n970), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_26__29__slave ( .q(_RegFile_26__29), .qb(n2315), .d(
        _RegFile_reg_26__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n970), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_26__2__master ( .q(_RegFile_reg_26__2__m2s), .d(
        n2871), .sdi(n4159), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n970), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_26__2__slave ( .q(_RegFile_26__2), .qb(n4158), .d(
        _RegFile_reg_26__2__m2s), .g(Ctrl__Regs_1__en2), .rb(n970), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_26__30__master ( .q(_RegFile_reg_26__30__m2s), .d(
        n2899), .sdi(n2315), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n970), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_26__30__slave ( .q(_RegFile_26__30), .qb(n2316), .d(
        _RegFile_reg_26__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n970), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_26__31__master ( .q(_RegFile_reg_26__31__m2s), .d(
        n2900), .sdi(n2316), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n933), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_26__31__slave ( .q(_RegFile_26__31), .qb(n2317), .d(
        _RegFile_reg_26__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n933), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_26__3__master ( .q(_RegFile_reg_26__3__m2s), .d(
        n2872), .sdi(n4158), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n933), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_26__3__slave ( .q(_RegFile_26__3), .qb(n4157), .d(
        _RegFile_reg_26__3__m2s), .g(Ctrl__Regs_1__en2), .rb(n933), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_26__4__master ( .q(_RegFile_reg_26__4__m2s), .d(
        n2873), .sdi(n4157), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n970), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_26__4__slave ( .q(_RegFile_26__4), .qb(n4156), .d(
        _RegFile_reg_26__4__m2s), .g(Ctrl__Regs_1__en2), .rb(n970), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_26__5__master ( .q(_RegFile_reg_26__5__m2s), .d(
        n2874), .sdi(n4156), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n933), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_26__5__slave ( .q(_RegFile_26__5), .qb(n4155), .d(
        _RegFile_reg_26__5__m2s), .g(Ctrl__Regs_1__en2), .rb(n933), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_26__6__master ( .q(_RegFile_reg_26__6__m2s), .d(
        n2875), .sdi(n4155), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n970), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_26__6__slave ( .q(_RegFile_26__6), .qb(n4154), .d(
        _RegFile_reg_26__6__m2s), .g(Ctrl__Regs_1__en2), .rb(n970), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_26__7__master ( .q(_RegFile_reg_26__7__m2s), .d(
        n2876), .sdi(n4154), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n933), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_26__7__slave ( .q(_RegFile_26__7), .qb(n4153), .d(
        _RegFile_reg_26__7__m2s), .g(Ctrl__Regs_1__en2), .rb(n933), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_26__8__master ( .q(_RegFile_reg_26__8__m2s), .d(
        n2877), .sdi(n4153), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n970), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_26__8__slave ( .q(_RegFile_26__8), .qb(n2318), .d(
        _RegFile_reg_26__8__m2s), .g(Ctrl__Regs_1__en2), .rb(n970), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_26__9__master ( .q(_RegFile_reg_26__9__m2s), .d(
        n2878), .sdi(n2318), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n933), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_26__9__slave ( .q(_RegFile_26__9), .qb(n2319), .d(
        _RegFile_reg_26__9__m2s), .g(Ctrl__Regs_1__en2), .rb(n933), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_27__0__master ( .q(_RegFile_reg_27__0__m2s), .d(
        n2837), .sdi(n2317), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n971), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_27__0__slave ( .q(_RegFile_27__0), .qb(n4152), .d(
        _RegFile_reg_27__0__m2s), .g(Ctrl__Regs_1__en2), .rb(n971), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_27__10__master ( .q(_RegFile_reg_27__10__m2s), .d(
        n2847), .sdi(n2343), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n971), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_27__10__slave ( .q(_RegFile_27__10), .qb(n2320), .d(
        _RegFile_reg_27__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n971), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_27__11__master ( .q(_RegFile_reg_27__11__m2s), .d(
        n2848), .sdi(n2320), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n933), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_27__11__slave ( .q(_RegFile_27__11), .qb(n2321), .d(
        _RegFile_reg_27__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n933), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_27__12__master ( .q(_RegFile_reg_27__12__m2s), .d(
        n2849), .sdi(n2321), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n971), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_27__12__slave ( .q(_RegFile_27__12), .qb(n2322), .d(
        _RegFile_reg_27__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n971), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_27__13__master ( .q(_RegFile_reg_27__13__m2s), .d(
        n2850), .sdi(n2322), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n933), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_27__13__slave ( .q(_RegFile_27__13), .qb(n2323), .d(
        _RegFile_reg_27__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n933), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_27__14__master ( .q(_RegFile_reg_27__14__m2s), .d(
        n2851), .sdi(n2323), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n971), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_27__14__slave ( .q(_RegFile_27__14), .qb(n2324), .d(
        _RegFile_reg_27__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n971), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_27__15__master ( .q(_RegFile_reg_27__15__m2s), .d(
        n2852), .sdi(n2324), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n933), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_27__15__slave ( .q(_RegFile_27__15), .qb(n2325), .d(
        _RegFile_reg_27__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n933), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_27__16__master ( .q(_RegFile_reg_27__16__m2s), .d(
        n2853), .sdi(n2325), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n971), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_27__16__slave ( .q(_RegFile_27__16), .qb(n2326), .d(
        _RegFile_reg_27__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n971), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_27__17__master ( .q(_RegFile_reg_27__17__m2s), .d(
        n2854), .sdi(n2326), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n933), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_27__17__slave ( .q(_RegFile_27__17), .qb(n2327), .d(
        _RegFile_reg_27__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n933), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_27__18__master ( .q(_RegFile_reg_27__18__m2s), .d(
        n2855), .sdi(n2327), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n971), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_27__18__slave ( .q(_RegFile_27__18), .qb(n2328), .d(
        _RegFile_reg_27__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n971), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_27__19__master ( .q(_RegFile_reg_27__19__m2s), .d(
        n2856), .sdi(n2328), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n933), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_27__19__slave ( .q(_RegFile_27__19), .qb(n2329), .d(
        _RegFile_reg_27__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n933), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_27__1__master ( .q(_RegFile_reg_27__1__m2s), .d(
        n2838), .sdi(n4152), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n933), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_27__1__slave ( .q(_RegFile_27__1), .qb(n4151), .d(
        _RegFile_reg_27__1__m2s), .g(Ctrl__Regs_1__en2), .rb(n933), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_27__20__master ( .q(_RegFile_reg_27__20__m2s), .d(
        n2857), .sdi(n2329), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n933), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_27__20__slave ( .q(_RegFile_27__20), .qb(n2330), .d(
        _RegFile_reg_27__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n933), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_27__21__master ( .q(_RegFile_reg_27__21__m2s), .d(
        n2858), .sdi(n2330), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n971), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_27__21__slave ( .q(_RegFile_27__21), .qb(n2331), .d(
        _RegFile_reg_27__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n971), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_27__22__master ( .q(_RegFile_reg_27__22__m2s), .d(
        n2859), .sdi(n2331), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_27__22__slave ( .q(_RegFile_27__22), .qb(n2332), .d(
        _RegFile_reg_27__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_27__23__master ( .q(_RegFile_reg_27__23__m2s), .d(
        n2860), .sdi(n2332), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n971), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_27__23__slave ( .q(_RegFile_27__23), .qb(n2333), .d(
        _RegFile_reg_27__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n971), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_27__24__master ( .q(_RegFile_reg_27__24__m2s), .d(
        n2861), .sdi(n2333), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_27__24__slave ( .q(_RegFile_27__24), .qb(n2334), .d(
        _RegFile_reg_27__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_27__25__master ( .q(_RegFile_reg_27__25__m2s), .d(
        n2862), .sdi(n2334), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n971), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_27__25__slave ( .q(_RegFile_27__25), .qb(n2335), .d(
        _RegFile_reg_27__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n971), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_27__26__master ( .q(_RegFile_reg_27__26__m2s), .d(
        n2863), .sdi(n2335), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_27__26__slave ( .q(_RegFile_27__26), .qb(n2336), .d(
        _RegFile_reg_27__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_27__27__master ( .q(_RegFile_reg_27__27__m2s), .d(
        n2864), .sdi(n2336), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n971), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_27__27__slave ( .q(_RegFile_27__27), .qb(n2337), .d(
        _RegFile_reg_27__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n971), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_27__28__master ( .q(_RegFile_reg_27__28__m2s), .d(
        n2865), .sdi(n2337), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_27__28__slave ( .q(_RegFile_27__28), .qb(n2338), .d(
        _RegFile_reg_27__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_27__29__master ( .q(_RegFile_reg_27__29__m2s), .d(
        n2866), .sdi(n2338), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n971), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_27__29__slave ( .q(_RegFile_27__29), .qb(n2339), .d(
        _RegFile_reg_27__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n971), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_27__2__master ( .q(_RegFile_reg_27__2__m2s), .d(
        n2839), .sdi(n4151), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n971), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_27__2__slave ( .q(_RegFile_27__2), .qb(n4150), .d(
        _RegFile_reg_27__2__m2s), .g(Ctrl__Regs_1__en2), .rb(n971), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_27__30__master ( .q(_RegFile_reg_27__30__m2s), .d(
        n2867), .sdi(n2339), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n971), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_27__30__slave ( .q(_RegFile_27__30), .qb(n2340), .d(
        _RegFile_reg_27__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n971), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_27__31__master ( .q(_RegFile_reg_27__31__m2s), .d(
        n2868), .sdi(n2340), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_27__31__slave ( .q(_RegFile_27__31), .qb(n2341), .d(
        _RegFile_reg_27__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_27__3__master ( .q(_RegFile_reg_27__3__m2s), .d(
        n2840), .sdi(n4150), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_27__3__slave ( .q(_RegFile_27__3), .qb(n4149), .d(
        _RegFile_reg_27__3__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_27__4__master ( .q(_RegFile_reg_27__4__m2s), .d(
        n2841), .sdi(n4149), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n971), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_27__4__slave ( .q(_RegFile_27__4), .qb(n4148), .d(
        _RegFile_reg_27__4__m2s), .g(Ctrl__Regs_1__en2), .rb(n971), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_27__5__master ( .q(_RegFile_reg_27__5__m2s), .d(
        n2842), .sdi(n4148), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_27__5__slave ( .q(_RegFile_27__5), .qb(n4147), .d(
        _RegFile_reg_27__5__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_27__6__master ( .q(_RegFile_reg_27__6__m2s), .d(
        n2843), .sdi(n4147), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n971), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_27__6__slave ( .q(_RegFile_27__6), .qb(n4146), .d(
        _RegFile_reg_27__6__m2s), .g(Ctrl__Regs_1__en2), .rb(n971), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_27__7__master ( .q(_RegFile_reg_27__7__m2s), .d(
        n2844), .sdi(n4146), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_27__7__slave ( .q(_RegFile_27__7), .qb(n4145), .d(
        _RegFile_reg_27__7__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_27__8__master ( .q(_RegFile_reg_27__8__m2s), .d(
        n2845), .sdi(n4145), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_27__8__slave ( .q(_RegFile_27__8), .qb(n2342), .d(
        _RegFile_reg_27__8__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_27__9__master ( .q(_RegFile_reg_27__9__m2s), .d(
        n2846), .sdi(n2342), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_27__9__slave ( .q(_RegFile_27__9), .qb(n2343), .d(
        _RegFile_reg_27__9__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_28__0__master ( .q(_RegFile_reg_28__0__m2s), .d(
        n2805), .sdi(n2341), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_28__0__slave ( .q(_RegFile_28__0), .qb(n4144), .d(
        _RegFile_reg_28__0__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_28__10__master ( .q(_RegFile_reg_28__10__m2s), .d(
        n2815), .sdi(n2367), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_28__10__slave ( .q(_RegFile_28__10), .qb(n2344), .d(
        _RegFile_reg_28__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_28__11__master ( .q(_RegFile_reg_28__11__m2s), .d(
        n2816), .sdi(n2344), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_28__11__slave ( .q(_RegFile_28__11), .qb(n2345), .d(
        _RegFile_reg_28__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_28__12__master ( .q(_RegFile_reg_28__12__m2s), .d(
        n2817), .sdi(n2345), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_28__12__slave ( .q(_RegFile_28__12), .qb(n2346), .d(
        _RegFile_reg_28__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_28__13__master ( .q(_RegFile_reg_28__13__m2s), .d(
        n2818), .sdi(n2346), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_28__13__slave ( .q(_RegFile_28__13), .qb(n2347), .d(
        _RegFile_reg_28__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_28__14__master ( .q(_RegFile_reg_28__14__m2s), .d(
        n2819), .sdi(n2347), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_28__14__slave ( .q(_RegFile_28__14), .qb(n2348), .d(
        _RegFile_reg_28__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_28__15__master ( .q(_RegFile_reg_28__15__m2s), .d(
        n2820), .sdi(n2348), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_28__15__slave ( .q(_RegFile_28__15), .qb(n2349), .d(
        _RegFile_reg_28__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_28__16__master ( .q(_RegFile_reg_28__16__m2s), .d(
        n2821), .sdi(n2349), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_28__16__slave ( .q(_RegFile_28__16), .qb(n2350), .d(
        _RegFile_reg_28__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_28__17__master ( .q(_RegFile_reg_28__17__m2s), .d(
        n2822), .sdi(n2350), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_28__17__slave ( .q(_RegFile_28__17), .qb(n2351), .d(
        _RegFile_reg_28__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_28__18__master ( .q(_RegFile_reg_28__18__m2s), .d(
        n2823), .sdi(n2351), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_28__18__slave ( .q(_RegFile_28__18), .qb(n2352), .d(
        _RegFile_reg_28__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_28__19__master ( .q(_RegFile_reg_28__19__m2s), .d(
        n2824), .sdi(n2352), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_28__19__slave ( .q(_RegFile_28__19), .qb(n2353), .d(
        _RegFile_reg_28__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_28__1__master ( .q(_RegFile_reg_28__1__m2s), .d(
        n2806), .sdi(n4144), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_28__1__slave ( .q(_RegFile_28__1), .qb(n4143), .d(
        _RegFile_reg_28__1__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_28__20__master ( .q(_RegFile_reg_28__20__m2s), .d(
        n2825), .sdi(n2353), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n931), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_28__20__slave ( .q(_RegFile_28__20), .qb(n2354), .d(
        _RegFile_reg_28__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n931), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_28__21__master ( .q(_RegFile_reg_28__21__m2s), .d(
        n2826), .sdi(n2354), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_28__21__slave ( .q(_RegFile_28__21), .qb(n2355), .d(
        _RegFile_reg_28__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_28__22__master ( .q(_RegFile_reg_28__22__m2s), .d(
        n2827), .sdi(n2355), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n931), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_28__22__slave ( .q(_RegFile_28__22), .qb(n2356), .d(
        _RegFile_reg_28__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n931), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_28__23__master ( .q(_RegFile_reg_28__23__m2s), .d(
        n2828), .sdi(n2356), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_28__23__slave ( .q(_RegFile_28__23), .qb(n2357), .d(
        _RegFile_reg_28__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_28__24__master ( .q(_RegFile_reg_28__24__m2s), .d(
        n2829), .sdi(n2357), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n931), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_28__24__slave ( .q(_RegFile_28__24), .qb(n2358), .d(
        _RegFile_reg_28__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n931), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_28__25__master ( .q(_RegFile_reg_28__25__m2s), .d(
        n2830), .sdi(n2358), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_28__25__slave ( .q(_RegFile_28__25), .qb(n2359), .d(
        _RegFile_reg_28__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_28__26__master ( .q(_RegFile_reg_28__26__m2s), .d(
        n2831), .sdi(n2359), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n931), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_28__26__slave ( .q(_RegFile_28__26), .qb(n2360), .d(
        _RegFile_reg_28__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n931), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_28__27__master ( .q(_RegFile_reg_28__27__m2s), .d(
        n2832), .sdi(n2360), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_28__27__slave ( .q(_RegFile_28__27), .qb(n2361), .d(
        _RegFile_reg_28__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_28__28__master ( .q(_RegFile_reg_28__28__m2s), .d(
        n2833), .sdi(n2361), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n931), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_28__28__slave ( .q(_RegFile_28__28), .qb(n2362), .d(
        _RegFile_reg_28__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n931), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_28__29__master ( .q(_RegFile_reg_28__29__m2s), .d(
        n2834), .sdi(n2362), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_28__29__slave ( .q(_RegFile_28__29), .qb(n2363), .d(
        _RegFile_reg_28__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_28__2__master ( .q(_RegFile_reg_28__2__m2s), .d(
        n2807), .sdi(n4143), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_28__2__slave ( .q(_RegFile_28__2), .qb(n4142), .d(
        _RegFile_reg_28__2__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_28__30__master ( .q(_RegFile_reg_28__30__m2s), .d(
        n2835), .sdi(n2363), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_28__30__slave ( .q(_RegFile_28__30), .qb(n2364), .d(
        _RegFile_reg_28__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_28__31__master ( .q(_RegFile_reg_28__31__m2s), .d(
        n2836), .sdi(n2364), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n931), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_28__31__slave ( .q(_RegFile_28__31), .qb(n2365), .d(
        _RegFile_reg_28__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n931), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_28__3__master ( .q(_RegFile_reg_28__3__m2s), .d(
        n2808), .sdi(n4142), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n931), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_28__3__slave ( .q(_RegFile_28__3), .qb(n4141), .d(
        _RegFile_reg_28__3__m2s), .g(Ctrl__Regs_1__en2), .rb(n931), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_28__4__master ( .q(_RegFile_reg_28__4__m2s), .d(
        n2809), .sdi(n4141), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_28__4__slave ( .q(_RegFile_28__4), .qb(n4140), .d(
        _RegFile_reg_28__4__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_28__5__master ( .q(_RegFile_reg_28__5__m2s), .d(
        n2810), .sdi(n4140), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n931), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_28__5__slave ( .q(_RegFile_28__5), .qb(n4139), .d(
        _RegFile_reg_28__5__m2s), .g(Ctrl__Regs_1__en2), .rb(n931), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_28__6__master ( .q(_RegFile_reg_28__6__m2s), .d(
        n2811), .sdi(n4139), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n972), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_28__6__slave ( .q(_RegFile_28__6), .qb(n4138), .d(
        _RegFile_reg_28__6__m2s), .g(Ctrl__Regs_1__en2), .rb(n972), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_28__7__master ( .q(_RegFile_reg_28__7__m2s), .d(
        n2812), .sdi(n4138), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n931), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_28__7__slave ( .q(_RegFile_28__7), .qb(n4137), .d(
        _RegFile_reg_28__7__m2s), .g(Ctrl__Regs_1__en2), .rb(n931), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_28__8__master ( .q(_RegFile_reg_28__8__m2s), .d(
        n2813), .sdi(n4137), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n972), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_28__8__slave ( .q(_RegFile_28__8), .qb(n2366), .d(
        _RegFile_reg_28__8__m2s), .g(Ctrl__Regs_1__en2), .rb(n972), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_28__9__master ( .q(_RegFile_reg_28__9__m2s), .d(
        n2814), .sdi(n2366), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n931), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_28__9__slave ( .q(_RegFile_28__9), .qb(n2367), .d(
        _RegFile_reg_28__9__m2s), .g(Ctrl__Regs_1__en2), .rb(n931), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_29__0__master ( .q(_RegFile_reg_29__0__m2s), .d(
        n2773), .sdi(n2365), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n972), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_29__0__slave ( .q(_RegFile_29__0), .qb(n4136), .d(
        _RegFile_reg_29__0__m2s), .g(Ctrl__Regs_1__en2), .rb(n972), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_29__10__master ( .q(_RegFile_reg_29__10__m2s), .d(
        n2783), .sdi(n2391), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n972), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_29__10__slave ( .q(_RegFile_29__10), .qb(n2368), .d(
        _RegFile_reg_29__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n972), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_29__11__master ( .q(_RegFile_reg_29__11__m2s), .d(
        n2784), .sdi(n2368), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n931), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_29__11__slave ( .q(_RegFile_29__11), .qb(n2369), .d(
        _RegFile_reg_29__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n931), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_29__12__master ( .q(_RegFile_reg_29__12__m2s), .d(
        n2785), .sdi(n2369), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n972), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_29__12__slave ( .q(_RegFile_29__12), .qb(n2370), .d(
        _RegFile_reg_29__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n972), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_29__13__master ( .q(_RegFile_reg_29__13__m2s), .d(
        n2786), .sdi(n2370), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n931), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_29__13__slave ( .q(_RegFile_29__13), .qb(n2371), .d(
        _RegFile_reg_29__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n931), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_29__14__master ( .q(_RegFile_reg_29__14__m2s), .d(
        n2787), .sdi(n2371), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n972), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_29__14__slave ( .q(_RegFile_29__14), .qb(n2372), .d(
        _RegFile_reg_29__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n972), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_29__15__master ( .q(_RegFile_reg_29__15__m2s), .d(
        n2788), .sdi(n2372), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n931), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_29__15__slave ( .q(_RegFile_29__15), .qb(n2373), .d(
        _RegFile_reg_29__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n931), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_29__16__master ( .q(_RegFile_reg_29__16__m2s), .d(
        n2789), .sdi(n2373), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n972), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_29__16__slave ( .q(_RegFile_29__16), .qb(n2374), .d(
        _RegFile_reg_29__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n972), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_29__17__master ( .q(_RegFile_reg_29__17__m2s), .d(
        n2790), .sdi(n2374), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n931), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_29__17__slave ( .q(_RegFile_29__17), .qb(n2375), .d(
        _RegFile_reg_29__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n931), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_29__18__master ( .q(_RegFile_reg_29__18__m2s), .d(
        n2791), .sdi(n2375), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n972), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_29__18__slave ( .q(_RegFile_29__18), .qb(n2376), .d(
        _RegFile_reg_29__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n972), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_29__19__master ( .q(_RegFile_reg_29__19__m2s), .d(
        n2792), .sdi(n2376), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n930), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_29__19__slave ( .q(_RegFile_29__19), .qb(n2377), .d(
        _RegFile_reg_29__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n930), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_29__1__master ( .q(_RegFile_reg_29__1__m2s), .d(
        n2774), .sdi(n4136), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n931), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_29__1__slave ( .q(_RegFile_29__1), .qb(n4135), .d(
        _RegFile_reg_29__1__m2s), .g(Ctrl__Regs_1__en2), .rb(n931), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_29__20__master ( .q(_RegFile_reg_29__20__m2s), .d(
        n2793), .sdi(n2377), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n930), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_29__20__slave ( .q(_RegFile_29__20), .qb(n2378), .d(
        _RegFile_reg_29__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n930), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_29__21__master ( .q(_RegFile_reg_29__21__m2s), .d(
        n2794), .sdi(n2378), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n972), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_29__21__slave ( .q(_RegFile_29__21), .qb(n2379), .d(
        _RegFile_reg_29__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n972), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_29__22__master ( .q(_RegFile_reg_29__22__m2s), .d(
        n2795), .sdi(n2379), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n930), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_29__22__slave ( .q(_RegFile_29__22), .qb(n2380), .d(
        _RegFile_reg_29__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n930), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_29__23__master ( .q(_RegFile_reg_29__23__m2s), .d(
        n2796), .sdi(n2380), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n972), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_29__23__slave ( .q(_RegFile_29__23), .qb(n2381), .d(
        _RegFile_reg_29__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n972), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_29__24__master ( .q(_RegFile_reg_29__24__m2s), .d(
        n2797), .sdi(n2381), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n930), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_29__24__slave ( .q(_RegFile_29__24), .qb(n2382), .d(
        _RegFile_reg_29__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n930), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_29__25__master ( .q(_RegFile_reg_29__25__m2s), .d(
        n2798), .sdi(n2382), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n972), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_29__25__slave ( .q(_RegFile_29__25), .qb(n2383), .d(
        _RegFile_reg_29__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n972), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_29__26__master ( .q(_RegFile_reg_29__26__m2s), .d(
        n2799), .sdi(n2383), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n930), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_29__26__slave ( .q(_RegFile_29__26), .qb(n2384), .d(
        _RegFile_reg_29__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n930), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_29__27__master ( .q(_RegFile_reg_29__27__m2s), .d(
        n2800), .sdi(n2384), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n972), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_29__27__slave ( .q(_RegFile_29__27), .qb(n2385), .d(
        _RegFile_reg_29__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n972), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_29__28__master ( .q(_RegFile_reg_29__28__m2s), .d(
        n2801), .sdi(n2385), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n930), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_29__28__slave ( .q(_RegFile_29__28), .qb(n2386), .d(
        _RegFile_reg_29__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n930), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_29__29__master ( .q(_RegFile_reg_29__29__m2s), .d(
        n2802), .sdi(n2386), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n972), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_29__29__slave ( .q(_RegFile_29__29), .qb(n2387), .d(
        _RegFile_reg_29__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n972), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_29__2__master ( .q(_RegFile_reg_29__2__m2s), .d(
        n2775), .sdi(n4135), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n972), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_29__2__slave ( .q(_RegFile_29__2), .qb(n4134), .d(
        _RegFile_reg_29__2__m2s), .g(Ctrl__Regs_1__en2), .rb(n972), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_29__30__master ( .q(_RegFile_reg_29__30__m2s), .d(
        n2803), .sdi(n2387), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n972), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_29__30__slave ( .q(_RegFile_29__30), .qb(n2388), .d(
        _RegFile_reg_29__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n972), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_29__31__master ( .q(_RegFile_reg_29__31__m2s), .d(
        n2804), .sdi(n2388), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n930), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_29__31__slave ( .q(_RegFile_29__31), .qb(n2389), .d(
        _RegFile_reg_29__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n930), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_29__3__master ( .q(_RegFile_reg_29__3__m2s), .d(
        n2776), .sdi(n4134), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n930), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_29__3__slave ( .q(_RegFile_29__3), .qb(n4133), .d(
        _RegFile_reg_29__3__m2s), .g(Ctrl__Regs_1__en2), .rb(n930), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_29__4__master ( .q(_RegFile_reg_29__4__m2s), .d(
        n2777), .sdi(n4133), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n973), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_29__4__slave ( .q(_RegFile_29__4), .qb(n4132), .d(
        _RegFile_reg_29__4__m2s), .g(Ctrl__Regs_1__en2), .rb(n973), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_29__5__master ( .q(_RegFile_reg_29__5__m2s), .d(
        n2778), .sdi(n4132), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n930), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_29__5__slave ( .q(_RegFile_29__5), .qb(n4131), .d(
        _RegFile_reg_29__5__m2s), .g(Ctrl__Regs_1__en2), .rb(n930), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_29__6__master ( .q(_RegFile_reg_29__6__m2s), .d(
        n2779), .sdi(n4131), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n973), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_29__6__slave ( .q(_RegFile_29__6), .qb(n4130), .d(
        _RegFile_reg_29__6__m2s), .g(Ctrl__Regs_1__en2), .rb(n973), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_29__7__master ( .q(_RegFile_reg_29__7__m2s), .d(
        n2780), .sdi(n4130), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n930), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_29__7__slave ( .q(_RegFile_29__7), .qb(n4129), .d(
        _RegFile_reg_29__7__m2s), .g(Ctrl__Regs_1__en2), .rb(n930), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_29__8__master ( .q(_RegFile_reg_29__8__m2s), .d(
        n2781), .sdi(n4129), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n973), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_29__8__slave ( .q(_RegFile_29__8), .qb(n2390), .d(
        _RegFile_reg_29__8__m2s), .g(Ctrl__Regs_1__en2), .rb(n973), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_29__9__master ( .q(_RegFile_reg_29__9__m2s), .d(
        n2782), .sdi(n2390), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n930), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_29__9__slave ( .q(_RegFile_29__9), .qb(n2391), .d(
        _RegFile_reg_29__9__m2s), .g(Ctrl__Regs_1__en2), .rb(n930), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_2__0__master ( .q(_RegFile_reg_2__0__m2s), .d(n3637
        ), .sdi(n2149), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n973), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_2__0__slave ( .q(_RegFile_2__0), .qb(n4352), .d(
        _RegFile_reg_2__0__m2s), .g(Ctrl__Regs_1__en2), .rb(n973), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_2__10__master ( .q(_RegFile_reg_2__10__m2s), .d(
        n3647), .sdi(n2415), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n973), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_2__10__slave ( .q(_RegFile_2__10), .qb(n2392), .d(
        _RegFile_reg_2__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n973), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_2__11__master ( .q(_RegFile_reg_2__11__m2s), .d(
        n3648), .sdi(n2392), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n930), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_2__11__slave ( .q(_RegFile_2__11), .qb(n2393), .d(
        _RegFile_reg_2__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n930), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_2__12__master ( .q(_RegFile_reg_2__12__m2s), .d(
        n3649), .sdi(n2393), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n973), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_2__12__slave ( .q(_RegFile_2__12), .qb(n2394), .d(
        _RegFile_reg_2__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n973), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_2__13__master ( .q(_RegFile_reg_2__13__m2s), .d(
        n3650), .sdi(n2394), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n930), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_2__13__slave ( .q(_RegFile_2__13), .qb(n2395), .d(
        _RegFile_reg_2__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n930), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_2__14__master ( .q(_RegFile_reg_2__14__m2s), .d(
        n3651), .sdi(n2395), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n973), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_2__14__slave ( .q(_RegFile_2__14), .qb(n2396), .d(
        _RegFile_reg_2__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n973), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_2__15__master ( .q(_RegFile_reg_2__15__m2s), .d(
        n3652), .sdi(n2396), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n930), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_2__15__slave ( .q(_RegFile_2__15), .qb(n2397), .d(
        _RegFile_reg_2__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n930), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_2__16__master ( .q(_RegFile_reg_2__16__m2s), .d(
        n3653), .sdi(n2397), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n973), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_2__16__slave ( .q(_RegFile_2__16), .qb(n2398), .d(
        _RegFile_reg_2__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n973), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_2__17__master ( .q(_RegFile_reg_2__17__m2s), .d(
        n3654), .sdi(n2398), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n929), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_2__17__slave ( .q(_RegFile_2__17), .qb(n2399), .d(
        _RegFile_reg_2__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n929), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_2__18__master ( .q(_RegFile_reg_2__18__m2s), .d(
        n3655), .sdi(n2399), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n973), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_2__18__slave ( .q(_RegFile_2__18), .qb(n2400), .d(
        _RegFile_reg_2__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n973), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_2__19__master ( .q(_RegFile_reg_2__19__m2s), .d(
        n3656), .sdi(n2400), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n929), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_2__19__slave ( .q(_RegFile_2__19), .qb(n2401), .d(
        _RegFile_reg_2__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n929), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_2__1__master ( .q(_RegFile_reg_2__1__m2s), .d(n3638
        ), .sdi(n4352), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n930), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_2__1__slave ( .q(_RegFile_2__1), .qb(n4351), .d(
        _RegFile_reg_2__1__m2s), .g(Ctrl__Regs_1__en2), .rb(n930), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_2__20__master ( .q(_RegFile_reg_2__20__m2s), .d(
        n3657), .sdi(n2401), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n929), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_2__20__slave ( .q(_RegFile_2__20), .qb(n2402), .d(
        _RegFile_reg_2__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n929), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_2__21__master ( .q(_RegFile_reg_2__21__m2s), .d(
        n3658), .sdi(n2402), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n973), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_2__21__slave ( .q(_RegFile_2__21), .qb(n2403), .d(
        _RegFile_reg_2__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n973), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_2__22__master ( .q(_RegFile_reg_2__22__m2s), .d(
        n3659), .sdi(n2403), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n929), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_2__22__slave ( .q(_RegFile_2__22), .qb(n2404), .d(
        _RegFile_reg_2__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n929), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_2__23__master ( .q(_RegFile_reg_2__23__m2s), .d(
        n3660), .sdi(n2404), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n973), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_2__23__slave ( .q(_RegFile_2__23), .qb(n2405), .d(
        _RegFile_reg_2__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n973), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_2__24__master ( .q(_RegFile_reg_2__24__m2s), .d(
        n3661), .sdi(n2405), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n929), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_2__24__slave ( .q(_RegFile_2__24), .qb(n2406), .d(
        _RegFile_reg_2__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n929), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_2__25__master ( .q(_RegFile_reg_2__25__m2s), .d(
        n3662), .sdi(n2406), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n973), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_2__25__slave ( .q(_RegFile_2__25), .qb(n2407), .d(
        _RegFile_reg_2__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n973), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_2__26__master ( .q(_RegFile_reg_2__26__m2s), .d(
        n3663), .sdi(n2407), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n929), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_2__26__slave ( .q(_RegFile_2__26), .qb(n2408), .d(
        _RegFile_reg_2__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n929), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_2__27__master ( .q(_RegFile_reg_2__27__m2s), .d(
        n3664), .sdi(n2408), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n973), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_2__27__slave ( .q(_RegFile_2__27), .qb(n2409), .d(
        _RegFile_reg_2__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n973), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_2__28__master ( .q(_RegFile_reg_2__28__m2s), .d(
        n3665), .sdi(n2409), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n929), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_2__28__slave ( .q(_RegFile_2__28), .qb(n2410), .d(
        _RegFile_reg_2__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n929), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_2__29__master ( .q(_RegFile_reg_2__29__m2s), .d(
        n3666), .sdi(n2410), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n973), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_2__29__slave ( .q(_RegFile_2__29), .qb(n2411), .d(
        _RegFile_reg_2__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n973), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_2__2__master ( .q(_RegFile_reg_2__2__m2s), .d(n3639
        ), .sdi(n4351), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n973), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_2__2__slave ( .q(_RegFile_2__2), .qb(n4350), .d(
        _RegFile_reg_2__2__m2s), .g(Ctrl__Regs_1__en2), .rb(n973), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_2__30__master ( .q(_RegFile_reg_2__30__m2s), .d(
        n3667), .sdi(n2411), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_2__30__slave ( .q(_RegFile_2__30), .qb(n2412), .d(
        _RegFile_reg_2__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_2__31__master ( .q(_RegFile_reg_2__31__m2s), .d(
        n3668), .sdi(n2412), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n929), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_2__31__slave ( .q(_RegFile_2__31), .qb(n2413), .d(
        _RegFile_reg_2__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n929), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_2__3__master ( .q(_RegFile_reg_2__3__m2s), .d(n3640
        ), .sdi(n4350), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n929), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_2__3__slave ( .q(_RegFile_2__3), .qb(n4349), .d(
        _RegFile_reg_2__3__m2s), .g(Ctrl__Regs_1__en2), .rb(n929), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_2__4__master ( .q(_RegFile_reg_2__4__m2s), .d(n3641
        ), .sdi(n4349), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_2__4__slave ( .q(_RegFile_2__4), .qb(n4348), .d(
        _RegFile_reg_2__4__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_2__5__master ( .q(_RegFile_reg_2__5__m2s), .d(n3642
        ), .sdi(n4348), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n929), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_2__5__slave ( .q(_RegFile_2__5), .qb(n4347), .d(
        _RegFile_reg_2__5__m2s), .g(Ctrl__Regs_1__en2), .rb(n929), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_2__6__master ( .q(_RegFile_reg_2__6__m2s), .d(n3643
        ), .sdi(n4347), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_2__6__slave ( .q(_RegFile_2__6), .qb(n4346), .d(
        _RegFile_reg_2__6__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_2__7__master ( .q(_RegFile_reg_2__7__m2s), .d(n3644
        ), .sdi(n4346), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n929), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_2__7__slave ( .q(_RegFile_2__7), .qb(n4345), .d(
        _RegFile_reg_2__7__m2s), .g(Ctrl__Regs_1__en2), .rb(n929), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_2__8__master ( .q(_RegFile_reg_2__8__m2s), .d(n3645
        ), .sdi(n4345), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_2__8__slave ( .q(_RegFile_2__8), .qb(n2414), .d(
        _RegFile_reg_2__8__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_2__9__master ( .q(_RegFile_reg_2__9__m2s), .d(n3646
        ), .sdi(n2414), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n929), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_2__9__slave ( .q(_RegFile_2__9), .qb(n2415), .d(
        _RegFile_reg_2__9__m2s), .g(Ctrl__Regs_1__en2), .rb(n929), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_30__0__master ( .q(_RegFile_reg_30__0__m2s), .d(
        n2741), .sdi(n2389), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_30__0__slave ( .q(_RegFile_30__0), .qb(n4128), .d(
        _RegFile_reg_30__0__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_30__10__master ( .q(_RegFile_reg_30__10__m2s), .d(
        n2751), .sdi(n2439), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_30__10__slave ( .q(_RegFile_30__10), .qb(n2416), .d(
        _RegFile_reg_30__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_30__11__master ( .q(_RegFile_reg_30__11__m2s), .d(
        n2752), .sdi(n2416), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n929), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_30__11__slave ( .q(_RegFile_30__11), .qb(n2417), .d(
        _RegFile_reg_30__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n929), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_30__12__master ( .q(_RegFile_reg_30__12__m2s), .d(
        n2753), .sdi(n2417), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_30__12__slave ( .q(_RegFile_30__12), .qb(n2418), .d(
        _RegFile_reg_30__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_30__13__master ( .q(_RegFile_reg_30__13__m2s), .d(
        n2754), .sdi(n2418), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n929), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_30__13__slave ( .q(_RegFile_30__13), .qb(n2419), .d(
        _RegFile_reg_30__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n929), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_30__14__master ( .q(_RegFile_reg_30__14__m2s), .d(
        n2755), .sdi(n2419), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_30__14__slave ( .q(_RegFile_30__14), .qb(n2420), .d(
        _RegFile_reg_30__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_30__15__master ( .q(_RegFile_reg_30__15__m2s), .d(
        n2756), .sdi(n2420), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n928), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_30__15__slave ( .q(_RegFile_30__15), .qb(n2421), .d(
        _RegFile_reg_30__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n928), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_30__16__master ( .q(_RegFile_reg_30__16__m2s), .d(
        n2757), .sdi(n2421), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_30__16__slave ( .q(_RegFile_30__16), .qb(n2422), .d(
        _RegFile_reg_30__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_30__17__master ( .q(_RegFile_reg_30__17__m2s), .d(
        n2758), .sdi(n2422), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n928), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_30__17__slave ( .q(_RegFile_30__17), .qb(n2423), .d(
        _RegFile_reg_30__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n928), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_30__18__master ( .q(_RegFile_reg_30__18__m2s), .d(
        n2759), .sdi(n2423), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_30__18__slave ( .q(_RegFile_30__18), .qb(n2424), .d(
        _RegFile_reg_30__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_30__19__master ( .q(_RegFile_reg_30__19__m2s), .d(
        n2760), .sdi(n2424), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n928), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_30__19__slave ( .q(_RegFile_30__19), .qb(n2425), .d(
        _RegFile_reg_30__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n928), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_30__1__master ( .q(_RegFile_reg_30__1__m2s), .d(
        n2742), .sdi(n4128), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n929), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_30__1__slave ( .q(_RegFile_30__1), .qb(n4127), .d(
        _RegFile_reg_30__1__m2s), .g(Ctrl__Regs_1__en2), .rb(n929), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_30__20__master ( .q(_RegFile_reg_30__20__m2s), .d(
        n2761), .sdi(n2425), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n928), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_30__20__slave ( .q(_RegFile_30__20), .qb(n2426), .d(
        _RegFile_reg_30__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n928), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_30__21__master ( .q(_RegFile_reg_30__21__m2s), .d(
        n2762), .sdi(n2426), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_30__21__slave ( .q(_RegFile_30__21), .qb(n2427), .d(
        _RegFile_reg_30__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_30__22__master ( .q(_RegFile_reg_30__22__m2s), .d(
        n2763), .sdi(n2427), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n928), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_30__22__slave ( .q(_RegFile_30__22), .qb(n2428), .d(
        _RegFile_reg_30__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n928), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_30__23__master ( .q(_RegFile_reg_30__23__m2s), .d(
        n2764), .sdi(n2428), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_30__23__slave ( .q(_RegFile_30__23), .qb(n2429), .d(
        _RegFile_reg_30__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_30__24__master ( .q(_RegFile_reg_30__24__m2s), .d(
        n2765), .sdi(n2429), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n928), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_30__24__slave ( .q(_RegFile_30__24), .qb(n2430), .d(
        _RegFile_reg_30__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n928), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_30__25__master ( .q(_RegFile_reg_30__25__m2s), .d(
        n2766), .sdi(n2430), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_30__25__slave ( .q(_RegFile_30__25), .qb(n2431), .d(
        _RegFile_reg_30__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_30__26__master ( .q(_RegFile_reg_30__26__m2s), .d(
        n2767), .sdi(n2431), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n928), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_30__26__slave ( .q(_RegFile_30__26), .qb(n2432), .d(
        _RegFile_reg_30__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n928), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_30__27__master ( .q(_RegFile_reg_30__27__m2s), .d(
        n2768), .sdi(n2432), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_30__27__slave ( .q(_RegFile_30__27), .qb(n2433), .d(
        _RegFile_reg_30__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_30__28__master ( .q(_RegFile_reg_30__28__m2s), .d(
        n2769), .sdi(n2433), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n928), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_30__28__slave ( .q(_RegFile_30__28), .qb(n2434), .d(
        _RegFile_reg_30__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n928), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_30__29__master ( .q(_RegFile_reg_30__29__m2s), .d(
        n2770), .sdi(n2434), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_30__29__slave ( .q(_RegFile_30__29), .qb(n2435), .d(
        _RegFile_reg_30__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_30__2__master ( .q(_RegFile_reg_30__2__m2s), .d(
        n2743), .sdi(n4127), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_30__2__slave ( .q(_RegFile_30__2), .qb(n4126), .d(
        _RegFile_reg_30__2__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_30__30__master ( .q(_RegFile_reg_30__30__m2s), .d(
        n2771), .sdi(n2435), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_30__30__slave ( .q(_RegFile_30__30), .qb(n2436), .d(
        _RegFile_reg_30__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_30__31__master ( .q(_RegFile_reg_30__31__m2s), .d(
        n2772), .sdi(n2436), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n928), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_30__31__slave ( .q(_RegFile_30__31), .qb(n2437), .d(
        _RegFile_reg_30__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n928), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_30__3__master ( .q(_RegFile_reg_30__3__m2s), .d(
        n2744), .sdi(n4126), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n928), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_30__3__slave ( .q(_RegFile_30__3), .qb(n4125), .d(
        _RegFile_reg_30__3__m2s), .g(Ctrl__Regs_1__en2), .rb(n928), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_30__4__master ( .q(_RegFile_reg_30__4__m2s), .d(
        n2745), .sdi(n4125), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_30__4__slave ( .q(_RegFile_30__4), .qb(n4124), .d(
        _RegFile_reg_30__4__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_30__5__master ( .q(_RegFile_reg_30__5__m2s), .d(
        n2746), .sdi(n4124), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n928), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_30__5__slave ( .q(_RegFile_30__5), .qb(n4123), .d(
        _RegFile_reg_30__5__m2s), .g(Ctrl__Regs_1__en2), .rb(n928), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_30__6__master ( .q(_RegFile_reg_30__6__m2s), .d(
        n2747), .sdi(n4123), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_30__6__slave ( .q(_RegFile_30__6), .qb(n4122), .d(
        _RegFile_reg_30__6__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_30__7__master ( .q(_RegFile_reg_30__7__m2s), .d(
        n2748), .sdi(n4122), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n928), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_30__7__slave ( .q(_RegFile_30__7), .qb(n4121), .d(
        _RegFile_reg_30__7__m2s), .g(Ctrl__Regs_1__en2), .rb(n928), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_30__8__master ( .q(_RegFile_reg_30__8__m2s), .d(
        n2749), .sdi(n4121), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_30__8__slave ( .q(_RegFile_30__8), .qb(n2438), .d(
        _RegFile_reg_30__8__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_30__9__master ( .q(_RegFile_reg_30__9__m2s), .d(
        n2750), .sdi(n2438), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n928), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_30__9__slave ( .q(_RegFile_30__9), .qb(n2439), .d(
        _RegFile_reg_30__9__m2s), .g(Ctrl__Regs_1__en2), .rb(n928), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_31__0__master ( .q(_RegFile_reg_31__0__m2s), .d(
        n2709), .sdi(n2437), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_31__0__slave ( .q(_RegFile_31__0), .qb(n4120), .d(
        _RegFile_reg_31__0__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_31__10__master ( .q(_RegFile_reg_31__10__m2s), .d(
        n2719), .sdi(n2463), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_31__10__slave ( .q(_RegFile_31__10), .qb(n2440), .d(
        _RegFile_reg_31__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_31__11__master ( .q(_RegFile_reg_31__11__m2s), .d(
        n2720), .sdi(n2440), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n928), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_31__11__slave ( .q(_RegFile_31__11), .qb(n2441), .d(
        _RegFile_reg_31__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n928), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_31__12__master ( .q(_RegFile_reg_31__12__m2s), .d(
        n2721), .sdi(n2441), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_31__12__slave ( .q(_RegFile_31__12), .qb(n2442), .d(
        _RegFile_reg_31__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_31__13__master ( .q(_RegFile_reg_31__13__m2s), .d(
        n2722), .sdi(n2442), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n927), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_31__13__slave ( .q(_RegFile_31__13), .qb(n2443), .d(
        _RegFile_reg_31__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n927), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_31__14__master ( .q(_RegFile_reg_31__14__m2s), .d(
        n2723), .sdi(n2443), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_31__14__slave ( .q(_RegFile_31__14), .qb(n2444), .d(
        _RegFile_reg_31__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_31__15__master ( .q(_RegFile_reg_31__15__m2s), .d(
        n2724), .sdi(n2444), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n927), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_31__15__slave ( .q(_RegFile_31__15), .qb(n2445), .d(
        _RegFile_reg_31__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n927), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_31__16__master ( .q(_RegFile_reg_31__16__m2s), .d(
        n2725), .sdi(n2445), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_31__16__slave ( .q(_RegFile_31__16), .qb(n2446), .d(
        _RegFile_reg_31__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_31__17__master ( .q(_RegFile_reg_31__17__m2s), .d(
        n2726), .sdi(n2446), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n927), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_31__17__slave ( .q(_RegFile_31__17), .qb(n2447), .d(
        _RegFile_reg_31__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n927), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_31__18__master ( .q(_RegFile_reg_31__18__m2s), .d(
        n2727), .sdi(n2447), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_31__18__slave ( .q(_RegFile_31__18), .qb(n2448), .d(
        _RegFile_reg_31__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_31__19__master ( .q(_RegFile_reg_31__19__m2s), .d(
        n2728), .sdi(n2448), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n927), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_31__19__slave ( .q(_RegFile_31__19), .qb(n2449), .d(
        _RegFile_reg_31__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n927), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_31__1__master ( .q(_RegFile_reg_31__1__m2s), .d(
        n2710), .sdi(n4120), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n928), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_31__1__slave ( .q(_RegFile_31__1), .qb(n4119), .d(
        _RegFile_reg_31__1__m2s), .g(Ctrl__Regs_1__en2), .rb(n928), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_31__20__master ( .q(_RegFile_reg_31__20__m2s), .d(
        n2729), .sdi(n2449), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n927), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_31__20__slave ( .q(_RegFile_31__20), .qb(n2450), .d(
        _RegFile_reg_31__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n927), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_31__21__master ( .q(_RegFile_reg_31__21__m2s), .d(
        n2730), .sdi(n2450), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_31__21__slave ( .q(_RegFile_31__21), .qb(n2451), .d(
        _RegFile_reg_31__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_31__22__master ( .q(_RegFile_reg_31__22__m2s), .d(
        n2731), .sdi(n2451), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n927), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_31__22__slave ( .q(_RegFile_31__22), .qb(n2452), .d(
        _RegFile_reg_31__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n927), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_31__23__master ( .q(_RegFile_reg_31__23__m2s), .d(
        n2732), .sdi(n2452), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_31__23__slave ( .q(_RegFile_31__23), .qb(n2453), .d(
        _RegFile_reg_31__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_31__24__master ( .q(_RegFile_reg_31__24__m2s), .d(
        n2733), .sdi(n2453), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n927), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_31__24__slave ( .q(_RegFile_31__24), .qb(n2454), .d(
        _RegFile_reg_31__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n927), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_31__25__master ( .q(_RegFile_reg_31__25__m2s), .d(
        n2734), .sdi(n2454), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_31__25__slave ( .q(_RegFile_31__25), .qb(n2455), .d(
        _RegFile_reg_31__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_31__26__master ( .q(_RegFile_reg_31__26__m2s), .d(
        n2735), .sdi(n2455), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n927), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_31__26__slave ( .q(_RegFile_31__26), .qb(n2456), .d(
        _RegFile_reg_31__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n927), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_31__27__master ( .q(_RegFile_reg_31__27__m2s), .d(
        n2736), .sdi(n2456), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_31__27__slave ( .q(_RegFile_31__27), .qb(n2457), .d(
        _RegFile_reg_31__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_31__28__master ( .q(_RegFile_reg_31__28__m2s), .d(
        n2737), .sdi(n2457), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n927), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_31__28__slave ( .q(_RegFile_31__28), .qb(n2458), .d(
        _RegFile_reg_31__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n927), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_31__29__master ( .q(_RegFile_reg_31__29__m2s), .d(
        n2738), .sdi(n2458), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_31__29__slave ( .q(_RegFile_31__29), .qb(n2459), .d(
        _RegFile_reg_31__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_31__2__master ( .q(_RegFile_reg_31__2__m2s), .d(
        n2711), .sdi(n4119), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_31__2__slave ( .q(_RegFile_31__2), .qb(n4118), .d(
        _RegFile_reg_31__2__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_31__30__master ( .q(_RegFile_reg_31__30__m2s), .d(
        n2739), .sdi(n2459), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_31__30__slave ( .q(_RegFile_31__30), .qb(n2460), .d(
        _RegFile_reg_31__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_31__31__master ( .q(_RegFile_reg_31__31__m2s), .d(
        n2740), .sdi(n2460), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n927), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_31__31__slave ( .q(_RegFile_31__31), .qb(n2461), .d(
        _RegFile_reg_31__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n927), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_31__3__master ( .q(_RegFile_reg_31__3__m2s), .d(
        n2712), .sdi(n4118), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n927), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_31__3__slave ( .q(_RegFile_31__3), .qb(n4117), .d(
        _RegFile_reg_31__3__m2s), .g(Ctrl__Regs_1__en2), .rb(n927), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_31__4__master ( .q(_RegFile_reg_31__4__m2s), .d(
        n2713), .sdi(n4117), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_31__4__slave ( .q(_RegFile_31__4), .qb(n4116), .d(
        _RegFile_reg_31__4__m2s), .g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_31__5__master ( .q(_RegFile_reg_31__5__m2s), .d(
        n2714), .sdi(n4116), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n927), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_31__5__slave ( .q(_RegFile_31__5), .qb(n4115), .d(
        _RegFile_reg_31__5__m2s), .g(Ctrl__Regs_1__en2), .rb(n927), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_31__6__master ( .q(_RegFile_reg_31__6__m2s), .d(
        n2715), .sdi(n4115), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_31__6__slave ( .q(_RegFile_31__6), .qb(n4114), .d(
        _RegFile_reg_31__6__m2s), .g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_31__7__master ( .q(_RegFile_reg_31__7__m2s), .d(
        n2716), .sdi(n4114), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n927), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_31__7__slave ( .q(_RegFile_31__7), .qb(n4113), .d(
        _RegFile_reg_31__7__m2s), .g(Ctrl__Regs_1__en2), .rb(n927), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_31__8__master ( .q(_RegFile_reg_31__8__m2s), .d(
        n2717), .sdi(n4113), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_31__8__slave ( .q(_RegFile_31__8), .qb(n2462), .d(
        _RegFile_reg_31__8__m2s), .g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_31__9__master ( .q(_RegFile_reg_31__9__m2s), .d(
        n2718), .sdi(n2462), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n927), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_31__9__slave ( .q(_RegFile_31__9), .qb(n2463), .d(
        _RegFile_reg_31__9__m2s), .g(Ctrl__Regs_1__en2), .rb(n927), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_3__0__master ( .q(_RegFile_reg_3__0__m2s), .d(n3605
        ), .sdi(n2413), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_3__0__slave ( .q(_RegFile_3__0), .qb(n4344), .d(
        _RegFile_reg_3__0__m2s), .g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_3__10__master ( .q(_RegFile_reg_3__10__m2s), .d(
        n3615), .sdi(n2487), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_3__10__slave ( .q(_RegFile_3__10), .qb(n2464), .d(
        _RegFile_reg_3__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_3__11__master ( .q(_RegFile_reg_3__11__m2s), .d(
        n3616), .sdi(n2464), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n926), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_3__11__slave ( .q(_RegFile_3__11), .qb(n2465), .d(
        _RegFile_reg_3__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n926), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_3__12__master ( .q(_RegFile_reg_3__12__m2s), .d(
        n3617), .sdi(n2465), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_3__12__slave ( .q(_RegFile_3__12), .qb(n2466), .d(
        _RegFile_reg_3__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_3__13__master ( .q(_RegFile_reg_3__13__m2s), .d(
        n3618), .sdi(n2466), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n926), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_3__13__slave ( .q(_RegFile_3__13), .qb(n2467), .d(
        _RegFile_reg_3__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n926), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_3__14__master ( .q(_RegFile_reg_3__14__m2s), .d(
        n3619), .sdi(n2467), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_3__14__slave ( .q(_RegFile_3__14), .qb(n2468), .d(
        _RegFile_reg_3__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_3__15__master ( .q(_RegFile_reg_3__15__m2s), .d(
        n3620), .sdi(n2468), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n926), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_3__15__slave ( .q(_RegFile_3__15), .qb(n2469), .d(
        _RegFile_reg_3__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n926), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_3__16__master ( .q(_RegFile_reg_3__16__m2s), .d(
        n3621), .sdi(n2469), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_3__16__slave ( .q(_RegFile_3__16), .qb(n2470), .d(
        _RegFile_reg_3__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_3__17__master ( .q(_RegFile_reg_3__17__m2s), .d(
        n3622), .sdi(n2470), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n926), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_3__17__slave ( .q(_RegFile_3__17), .qb(n2471), .d(
        _RegFile_reg_3__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n926), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_3__18__master ( .q(_RegFile_reg_3__18__m2s), .d(
        n3623), .sdi(n2471), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_3__18__slave ( .q(_RegFile_3__18), .qb(n2472), .d(
        _RegFile_reg_3__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_3__19__master ( .q(_RegFile_reg_3__19__m2s), .d(
        n3624), .sdi(n2472), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n926), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_3__19__slave ( .q(_RegFile_3__19), .qb(n2473), .d(
        _RegFile_reg_3__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n926), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_3__1__master ( .q(_RegFile_reg_3__1__m2s), .d(n3606
        ), .sdi(n4344), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n927), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_3__1__slave ( .q(_RegFile_3__1), .qb(n4343), .d(
        _RegFile_reg_3__1__m2s), .g(Ctrl__Regs_1__en2), .rb(n927), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_3__20__master ( .q(_RegFile_reg_3__20__m2s), .d(
        n3625), .sdi(n2473), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n926), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_3__20__slave ( .q(_RegFile_3__20), .qb(n2474), .d(
        _RegFile_reg_3__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n926), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_3__21__master ( .q(_RegFile_reg_3__21__m2s), .d(
        n3626), .sdi(n2474), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_3__21__slave ( .q(_RegFile_3__21), .qb(n2475), .d(
        _RegFile_reg_3__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_3__22__master ( .q(_RegFile_reg_3__22__m2s), .d(
        n3627), .sdi(n2475), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n926), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_3__22__slave ( .q(_RegFile_3__22), .qb(n2476), .d(
        _RegFile_reg_3__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n926), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_3__23__master ( .q(_RegFile_reg_3__23__m2s), .d(
        n3628), .sdi(n2476), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_3__23__slave ( .q(_RegFile_3__23), .qb(n2477), .d(
        _RegFile_reg_3__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_3__24__master ( .q(_RegFile_reg_3__24__m2s), .d(
        n3629), .sdi(n2477), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n926), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_3__24__slave ( .q(_RegFile_3__24), .qb(n2478), .d(
        _RegFile_reg_3__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n926), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_3__25__master ( .q(_RegFile_reg_3__25__m2s), .d(
        n3630), .sdi(n2478), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_3__25__slave ( .q(_RegFile_3__25), .qb(n2479), .d(
        _RegFile_reg_3__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_3__26__master ( .q(_RegFile_reg_3__26__m2s), .d(
        n3631), .sdi(n2479), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n926), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_3__26__slave ( .q(_RegFile_3__26), .qb(n2480), .d(
        _RegFile_reg_3__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n926), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_3__27__master ( .q(_RegFile_reg_3__27__m2s), .d(
        n3632), .sdi(n2480), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_3__27__slave ( .q(_RegFile_3__27), .qb(n2481), .d(
        _RegFile_reg_3__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_3__28__master ( .q(_RegFile_reg_3__28__m2s), .d(
        n3633), .sdi(n2481), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n926), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_3__28__slave ( .q(_RegFile_3__28), .qb(n2482), .d(
        _RegFile_reg_3__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n926), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_3__29__master ( .q(_RegFile_reg_3__29__m2s), .d(
        n3634), .sdi(n2482), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_3__29__slave ( .q(_RegFile_3__29), .qb(n2483), .d(
        _RegFile_reg_3__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_3__2__master ( .q(_RegFile_reg_3__2__m2s), .d(n3607
        ), .sdi(n4343), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_3__2__slave ( .q(_RegFile_3__2), .qb(n4342), .d(
        _RegFile_reg_3__2__m2s), .g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_3__30__master ( .q(_RegFile_reg_3__30__m2s), .d(
        n3635), .sdi(n2483), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_3__30__slave ( .q(_RegFile_3__30), .qb(n2484), .d(
        _RegFile_reg_3__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_3__31__master ( .q(_RegFile_reg_3__31__m2s), .d(
        n3636), .sdi(n2484), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n926), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_3__31__slave ( .q(_RegFile_3__31), .qb(n2485), .d(
        _RegFile_reg_3__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n926), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_3__3__master ( .q(_RegFile_reg_3__3__m2s), .d(n3608
        ), .sdi(n4342), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n926), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_3__3__slave ( .q(_RegFile_3__3), .qb(n4341), .d(
        _RegFile_reg_3__3__m2s), .g(Ctrl__Regs_1__en2), .rb(n926), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_3__4__master ( .q(_RegFile_reg_3__4__m2s), .d(n3609
        ), .sdi(n4341), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_3__4__slave ( .q(_RegFile_3__4), .qb(n4340), .d(
        _RegFile_reg_3__4__m2s), .g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_3__5__master ( .q(_RegFile_reg_3__5__m2s), .d(n3610
        ), .sdi(n4340), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n926), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_3__5__slave ( .q(_RegFile_3__5), .qb(n4339), .d(
        _RegFile_reg_3__5__m2s), .g(Ctrl__Regs_1__en2), .rb(n926), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_3__6__master ( .q(_RegFile_reg_3__6__m2s), .d(n3611
        ), .sdi(n4339), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_3__6__slave ( .q(_RegFile_3__6), .qb(n4338), .d(
        _RegFile_reg_3__6__m2s), .g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_3__7__master ( .q(_RegFile_reg_3__7__m2s), .d(n3612
        ), .sdi(n4338), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n926), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_3__7__slave ( .q(_RegFile_3__7), .qb(n4337), .d(
        _RegFile_reg_3__7__m2s), .g(Ctrl__Regs_1__en2), .rb(n926), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_3__8__master ( .q(_RegFile_reg_3__8__m2s), .d(n3613
        ), .sdi(n4337), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_3__8__slave ( .q(_RegFile_3__8), .qb(n2486), .d(
        _RegFile_reg_3__8__m2s), .g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_3__9__master ( .q(_RegFile_reg_3__9__m2s), .d(n3614
        ), .sdi(n2486), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n926), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_3__9__slave ( .q(_RegFile_3__9), .qb(n2487), .d(
        _RegFile_reg_3__9__m2s), .g(Ctrl__Regs_1__en2), .rb(n926), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_4__0__master ( .q(_RegFile_reg_4__0__m2s), .d(n3573
        ), .sdi(n2485), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_4__0__slave ( .q(_RegFile_4__0), .qb(n4336), .d(
        _RegFile_reg_4__0__m2s), .g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_4__10__master ( .q(_RegFile_reg_4__10__m2s), .d(
        n3583), .sdi(n2511), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_4__10__slave ( .q(_RegFile_4__10), .qb(n2488), .d(
        _RegFile_reg_4__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_4__11__master ( .q(_RegFile_reg_4__11__m2s), .d(
        n3584), .sdi(n2488), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n925), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_4__11__slave ( .q(_RegFile_4__11), .qb(n2489), .d(
        _RegFile_reg_4__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n925), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_4__12__master ( .q(_RegFile_reg_4__12__m2s), .d(
        n3585), .sdi(n2489), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_4__12__slave ( .q(_RegFile_4__12), .qb(n2490), .d(
        _RegFile_reg_4__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_4__13__master ( .q(_RegFile_reg_4__13__m2s), .d(
        n3586), .sdi(n2490), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n925), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_4__13__slave ( .q(_RegFile_4__13), .qb(n2491), .d(
        _RegFile_reg_4__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n925), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_4__14__master ( .q(_RegFile_reg_4__14__m2s), .d(
        n3587), .sdi(n2491), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_4__14__slave ( .q(_RegFile_4__14), .qb(n2492), .d(
        _RegFile_reg_4__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_4__15__master ( .q(_RegFile_reg_4__15__m2s), .d(
        n3588), .sdi(n2492), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n925), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_4__15__slave ( .q(_RegFile_4__15), .qb(n2493), .d(
        _RegFile_reg_4__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n925), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_4__16__master ( .q(_RegFile_reg_4__16__m2s), .d(
        n3589), .sdi(n2493), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_4__16__slave ( .q(_RegFile_4__16), .qb(n2494), .d(
        _RegFile_reg_4__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_4__17__master ( .q(_RegFile_reg_4__17__m2s), .d(
        n3590), .sdi(n2494), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n925), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_4__17__slave ( .q(_RegFile_4__17), .qb(n2495), .d(
        _RegFile_reg_4__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n925), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_4__18__master ( .q(_RegFile_reg_4__18__m2s), .d(
        n3591), .sdi(n2495), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_4__18__slave ( .q(_RegFile_4__18), .qb(n2496), .d(
        _RegFile_reg_4__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_4__19__master ( .q(_RegFile_reg_4__19__m2s), .d(
        n3592), .sdi(n2496), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n925), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_4__19__slave ( .q(_RegFile_4__19), .qb(n2497), .d(
        _RegFile_reg_4__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n925), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_4__1__master ( .q(_RegFile_reg_4__1__m2s), .d(n3574
        ), .sdi(n4336), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n925), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_4__1__slave ( .q(_RegFile_4__1), .qb(n4335), .d(
        _RegFile_reg_4__1__m2s), .g(Ctrl__Regs_1__en2), .rb(n925), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_4__20__master ( .q(_RegFile_reg_4__20__m2s), .d(
        n3593), .sdi(n2497), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n925), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_4__20__slave ( .q(_RegFile_4__20), .qb(n2498), .d(
        _RegFile_reg_4__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n925), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_4__21__master ( .q(_RegFile_reg_4__21__m2s), .d(
        n3594), .sdi(n2498), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_4__21__slave ( .q(_RegFile_4__21), .qb(n2499), .d(
        _RegFile_reg_4__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_4__22__master ( .q(_RegFile_reg_4__22__m2s), .d(
        n3595), .sdi(n2499), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n925), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_4__22__slave ( .q(_RegFile_4__22), .qb(n2500), .d(
        _RegFile_reg_4__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n925), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_4__23__master ( .q(_RegFile_reg_4__23__m2s), .d(
        n3596), .sdi(n2500), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n977), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_4__23__slave ( .q(_RegFile_4__23), .qb(n2501), .d(
        _RegFile_reg_4__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n977), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_4__24__master ( .q(_RegFile_reg_4__24__m2s), .d(
        n3597), .sdi(n2501), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n925), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_4__24__slave ( .q(_RegFile_4__24), .qb(n2502), .d(
        _RegFile_reg_4__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n925), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_4__25__master ( .q(_RegFile_reg_4__25__m2s), .d(
        n3598), .sdi(n2502), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n977), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_4__25__slave ( .q(_RegFile_4__25), .qb(n2503), .d(
        _RegFile_reg_4__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n977), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_4__26__master ( .q(_RegFile_reg_4__26__m2s), .d(
        n3599), .sdi(n2503), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n925), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_4__26__slave ( .q(_RegFile_4__26), .qb(n2504), .d(
        _RegFile_reg_4__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n925), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_4__27__master ( .q(_RegFile_reg_4__27__m2s), .d(
        n3600), .sdi(n2504), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n977), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_4__27__slave ( .q(_RegFile_4__27), .qb(n2505), .d(
        _RegFile_reg_4__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n977), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_4__28__master ( .q(_RegFile_reg_4__28__m2s), .d(
        n3601), .sdi(n2505), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n925), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_4__28__slave ( .q(_RegFile_4__28), .qb(n2506), .d(
        _RegFile_reg_4__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n925), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_4__29__master ( .q(_RegFile_reg_4__29__m2s), .d(
        n3602), .sdi(n2506), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n977), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_4__29__slave ( .q(_RegFile_4__29), .qb(n2507), .d(
        _RegFile_reg_4__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n977), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_4__2__master ( .q(_RegFile_reg_4__2__m2s), .d(n3575
        ), .sdi(n4335), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_4__2__slave ( .q(_RegFile_4__2), .qb(n4334), .d(
        _RegFile_reg_4__2__m2s), .g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_4__30__master ( .q(_RegFile_reg_4__30__m2s), .d(
        n3603), .sdi(n2507), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n977), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_4__30__slave ( .q(_RegFile_4__30), .qb(n2508), .d(
        _RegFile_reg_4__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n977), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_4__31__master ( .q(_RegFile_reg_4__31__m2s), .d(
        n3604), .sdi(n2508), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n925), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_4__31__slave ( .q(_RegFile_4__31), .qb(n2509), .d(
        _RegFile_reg_4__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n925), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_4__3__master ( .q(_RegFile_reg_4__3__m2s), .d(n3576
        ), .sdi(n4334), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n925), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_4__3__slave ( .q(_RegFile_4__3), .qb(n4333), .d(
        _RegFile_reg_4__3__m2s), .g(Ctrl__Regs_1__en2), .rb(n925), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_4__4__master ( .q(_RegFile_reg_4__4__m2s), .d(n3577
        ), .sdi(n4333), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n977), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_4__4__slave ( .q(_RegFile_4__4), .qb(n4332), .d(
        _RegFile_reg_4__4__m2s), .g(Ctrl__Regs_1__en2), .rb(n977), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_4__5__master ( .q(_RegFile_reg_4__5__m2s), .d(n3578
        ), .sdi(n4332), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n925), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_4__5__slave ( .q(_RegFile_4__5), .qb(n4331), .d(
        _RegFile_reg_4__5__m2s), .g(Ctrl__Regs_1__en2), .rb(n925), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_4__6__master ( .q(_RegFile_reg_4__6__m2s), .d(n3579
        ), .sdi(n4331), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n977), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_4__6__slave ( .q(_RegFile_4__6), .qb(n4330), .d(
        _RegFile_reg_4__6__m2s), .g(Ctrl__Regs_1__en2), .rb(n977), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_4__7__master ( .q(_RegFile_reg_4__7__m2s), .d(n3580
        ), .sdi(n4330), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n925), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_4__7__slave ( .q(_RegFile_4__7), .qb(n4329), .d(
        _RegFile_reg_4__7__m2s), .g(Ctrl__Regs_1__en2), .rb(n925), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_4__8__master ( .q(_RegFile_reg_4__8__m2s), .d(n3581
        ), .sdi(n4329), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n977), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_4__8__slave ( .q(_RegFile_4__8), .qb(n2510), .d(
        _RegFile_reg_4__8__m2s), .g(Ctrl__Regs_1__en2), .rb(n977), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_4__9__master ( .q(_RegFile_reg_4__9__m2s), .d(n3582
        ), .sdi(n2510), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n924), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_4__9__slave ( .q(_RegFile_4__9), .qb(n2511), .d(
        _RegFile_reg_4__9__m2s), .g(Ctrl__Regs_1__en2), .rb(n924), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_5__0__master ( .q(_RegFile_reg_5__0__m2s), .d(n3541
        ), .sdi(n2509), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n977), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_5__0__slave ( .q(_RegFile_5__0), .qb(n4328), .d(
        _RegFile_reg_5__0__m2s), .g(Ctrl__Regs_1__en2), .rb(n977), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_5__10__master ( .q(_RegFile_reg_5__10__m2s), .d(
        n3551), .sdi(n2535), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n977), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_5__10__slave ( .q(_RegFile_5__10), .qb(n2512), .d(
        _RegFile_reg_5__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n977), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_5__11__master ( .q(_RegFile_reg_5__11__m2s), .d(
        n3552), .sdi(n2512), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n924), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_5__11__slave ( .q(_RegFile_5__11), .qb(n2513), .d(
        _RegFile_reg_5__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n924), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_5__12__master ( .q(_RegFile_reg_5__12__m2s), .d(
        n3553), .sdi(n2513), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n977), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_5__12__slave ( .q(_RegFile_5__12), .qb(n2514), .d(
        _RegFile_reg_5__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n977), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_5__13__master ( .q(_RegFile_reg_5__13__m2s), .d(
        n3554), .sdi(n2514), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n924), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_5__13__slave ( .q(_RegFile_5__13), .qb(n2515), .d(
        _RegFile_reg_5__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n924), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_5__14__master ( .q(_RegFile_reg_5__14__m2s), .d(
        n3555), .sdi(n2515), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n977), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_5__14__slave ( .q(_RegFile_5__14), .qb(n2516), .d(
        _RegFile_reg_5__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n977), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_5__15__master ( .q(_RegFile_reg_5__15__m2s), .d(
        n3556), .sdi(n2516), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n924), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_5__15__slave ( .q(_RegFile_5__15), .qb(n2517), .d(
        _RegFile_reg_5__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n924), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_5__16__master ( .q(_RegFile_reg_5__16__m2s), .d(
        n3557), .sdi(n2517), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n977), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_5__16__slave ( .q(_RegFile_5__16), .qb(n2518), .d(
        _RegFile_reg_5__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n977), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_5__17__master ( .q(_RegFile_reg_5__17__m2s), .d(
        n3558), .sdi(n2518), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n924), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_5__17__slave ( .q(_RegFile_5__17), .qb(n2519), .d(
        _RegFile_reg_5__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n924), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_5__18__master ( .q(_RegFile_reg_5__18__m2s), .d(
        n3559), .sdi(n2519), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n977), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_5__18__slave ( .q(_RegFile_5__18), .qb(n2520), .d(
        _RegFile_reg_5__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n977), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_5__19__master ( .q(_RegFile_reg_5__19__m2s), .d(
        n3560), .sdi(n2520), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n924), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_5__19__slave ( .q(_RegFile_5__19), .qb(n2521), .d(
        _RegFile_reg_5__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n924), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_5__1__master ( .q(_RegFile_reg_5__1__m2s), .d(n3542
        ), .sdi(n4328), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n924), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_5__1__slave ( .q(_RegFile_5__1), .qb(n4327), .d(
        _RegFile_reg_5__1__m2s), .g(Ctrl__Regs_1__en2), .rb(n924), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_5__20__master ( .q(_RegFile_reg_5__20__m2s), .d(
        n3561), .sdi(n2521), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n924), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_5__20__slave ( .q(_RegFile_5__20), .qb(n2522), .d(
        _RegFile_reg_5__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n924), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_5__21__master ( .q(_RegFile_reg_5__21__m2s), .d(
        n3562), .sdi(n2522), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n978), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_5__21__slave ( .q(_RegFile_5__21), .qb(n2523), .d(
        _RegFile_reg_5__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n978), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_5__22__master ( .q(_RegFile_reg_5__22__m2s), .d(
        n3563), .sdi(n2523), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n924), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_5__22__slave ( .q(_RegFile_5__22), .qb(n2524), .d(
        _RegFile_reg_5__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n924), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_5__23__master ( .q(_RegFile_reg_5__23__m2s), .d(
        n3564), .sdi(n2524), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n978), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_5__23__slave ( .q(_RegFile_5__23), .qb(n2525), .d(
        _RegFile_reg_5__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n978), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_5__24__master ( .q(_RegFile_reg_5__24__m2s), .d(
        n3565), .sdi(n2525), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n924), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_5__24__slave ( .q(_RegFile_5__24), .qb(n2526), .d(
        _RegFile_reg_5__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n924), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_5__25__master ( .q(_RegFile_reg_5__25__m2s), .d(
        n3566), .sdi(n2526), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n978), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_5__25__slave ( .q(_RegFile_5__25), .qb(n2527), .d(
        _RegFile_reg_5__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n978), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_5__26__master ( .q(_RegFile_reg_5__26__m2s), .d(
        n3567), .sdi(n2527), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n924), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_5__26__slave ( .q(_RegFile_5__26), .qb(n2528), .d(
        _RegFile_reg_5__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n924), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_5__27__master ( .q(_RegFile_reg_5__27__m2s), .d(
        n3568), .sdi(n2528), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n978), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_5__27__slave ( .q(_RegFile_5__27), .qb(n2529), .d(
        _RegFile_reg_5__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n978), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_5__28__master ( .q(_RegFile_reg_5__28__m2s), .d(
        n3569), .sdi(n2529), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n924), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_5__28__slave ( .q(_RegFile_5__28), .qb(n2530), .d(
        _RegFile_reg_5__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n924), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_5__29__master ( .q(_RegFile_reg_5__29__m2s), .d(
        n3570), .sdi(n2530), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n978), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_5__29__slave ( .q(_RegFile_5__29), .qb(n2531), .d(
        _RegFile_reg_5__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n978), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_5__2__master ( .q(_RegFile_reg_5__2__m2s), .d(n3543
        ), .sdi(n4327), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n977), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_5__2__slave ( .q(_RegFile_5__2), .qb(n4326), .d(
        _RegFile_reg_5__2__m2s), .g(Ctrl__Regs_1__en2), .rb(n977), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_5__30__master ( .q(_RegFile_reg_5__30__m2s), .d(
        n3571), .sdi(n2531), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n978), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_5__30__slave ( .q(_RegFile_5__30), .qb(n2532), .d(
        _RegFile_reg_5__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n978), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_5__31__master ( .q(_RegFile_reg_5__31__m2s), .d(
        n3572), .sdi(n2532), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n924), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_5__31__slave ( .q(_RegFile_5__31), .qb(n2533), .d(
        _RegFile_reg_5__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n924), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_5__3__master ( .q(_RegFile_reg_5__3__m2s), .d(n3544
        ), .sdi(n4326), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n924), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_5__3__slave ( .q(_RegFile_5__3), .qb(n4325), .d(
        _RegFile_reg_5__3__m2s), .g(Ctrl__Regs_1__en2), .rb(n924), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_5__4__master ( .q(_RegFile_reg_5__4__m2s), .d(n3545
        ), .sdi(n4325), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n978), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_5__4__slave ( .q(_RegFile_5__4), .qb(n4324), .d(
        _RegFile_reg_5__4__m2s), .g(Ctrl__Regs_1__en2), .rb(n978), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_5__5__master ( .q(_RegFile_reg_5__5__m2s), .d(n3546
        ), .sdi(n4324), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n924), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_5__5__slave ( .q(_RegFile_5__5), .qb(n4323), .d(
        _RegFile_reg_5__5__m2s), .g(Ctrl__Regs_1__en2), .rb(n924), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_5__6__master ( .q(_RegFile_reg_5__6__m2s), .d(n3547
        ), .sdi(n4323), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n978), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_5__6__slave ( .q(_RegFile_5__6), .qb(n4322), .d(
        _RegFile_reg_5__6__m2s), .g(Ctrl__Regs_1__en2), .rb(n978), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_5__7__master ( .q(_RegFile_reg_5__7__m2s), .d(n3548
        ), .sdi(n4322), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_5__7__slave ( .q(_RegFile_5__7), .qb(n4321), .d(
        _RegFile_reg_5__7__m2s), .g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_5__8__master ( .q(_RegFile_reg_5__8__m2s), .d(n3549
        ), .sdi(n4321), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n978), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_5__8__slave ( .q(_RegFile_5__8), .qb(n2534), .d(
        _RegFile_reg_5__8__m2s), .g(Ctrl__Regs_1__en2), .rb(n978), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_5__9__master ( .q(_RegFile_reg_5__9__m2s), .d(n3550
        ), .sdi(n2534), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_5__9__slave ( .q(_RegFile_5__9), .qb(n2535), .d(
        _RegFile_reg_5__9__m2s), .g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_6__0__master ( .q(_RegFile_reg_6__0__m2s), .d(n3509
        ), .sdi(n2533), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n978), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_6__0__slave ( .q(_RegFile_6__0), .qb(n4320), .d(
        _RegFile_reg_6__0__m2s), .g(Ctrl__Regs_1__en2), .rb(n978), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_6__10__master ( .q(_RegFile_reg_6__10__m2s), .d(
        n3519), .sdi(n2559), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n978), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_6__10__slave ( .q(_RegFile_6__10), .qb(n2536), .d(
        _RegFile_reg_6__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n978), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_6__11__master ( .q(_RegFile_reg_6__11__m2s), .d(
        n3520), .sdi(n2536), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_6__11__slave ( .q(_RegFile_6__11), .qb(n2537), .d(
        _RegFile_reg_6__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_6__12__master ( .q(_RegFile_reg_6__12__m2s), .d(
        n3521), .sdi(n2537), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n978), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_6__12__slave ( .q(_RegFile_6__12), .qb(n2538), .d(
        _RegFile_reg_6__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n978), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_6__13__master ( .q(_RegFile_reg_6__13__m2s), .d(
        n3522), .sdi(n2538), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_6__13__slave ( .q(_RegFile_6__13), .qb(n2539), .d(
        _RegFile_reg_6__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_6__14__master ( .q(_RegFile_reg_6__14__m2s), .d(
        n3523), .sdi(n2539), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n978), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_6__14__slave ( .q(_RegFile_6__14), .qb(n2540), .d(
        _RegFile_reg_6__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n978), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_6__15__master ( .q(_RegFile_reg_6__15__m2s), .d(
        n3524), .sdi(n2540), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_6__15__slave ( .q(_RegFile_6__15), .qb(n2541), .d(
        _RegFile_reg_6__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_6__16__master ( .q(_RegFile_reg_6__16__m2s), .d(
        n3525), .sdi(n2541), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n978), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_6__16__slave ( .q(_RegFile_6__16), .qb(n2542), .d(
        _RegFile_reg_6__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n978), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_6__17__master ( .q(_RegFile_reg_6__17__m2s), .d(
        n3526), .sdi(n2542), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_6__17__slave ( .q(_RegFile_6__17), .qb(n2543), .d(
        _RegFile_reg_6__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_6__18__master ( .q(_RegFile_reg_6__18__m2s), .d(
        n3527), .sdi(n2543), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n978), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_6__18__slave ( .q(_RegFile_6__18), .qb(n2544), .d(
        _RegFile_reg_6__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n978), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_6__19__master ( .q(_RegFile_reg_6__19__m2s), .d(
        n3528), .sdi(n2544), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_6__19__slave ( .q(_RegFile_6__19), .qb(n2545), .d(
        _RegFile_reg_6__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_6__1__master ( .q(_RegFile_reg_6__1__m2s), .d(n3510
        ), .sdi(n4320), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_6__1__slave ( .q(_RegFile_6__1), .qb(n4319), .d(
        _RegFile_reg_6__1__m2s), .g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_6__20__master ( .q(_RegFile_reg_6__20__m2s), .d(
        n3529), .sdi(n2545), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_6__20__slave ( .q(_RegFile_6__20), .qb(n2546), .d(
        _RegFile_reg_6__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_6__21__master ( .q(_RegFile_reg_6__21__m2s), .d(
        n3530), .sdi(n2546), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n979), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_6__21__slave ( .q(_RegFile_6__21), .qb(n2547), .d(
        _RegFile_reg_6__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n979), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_6__22__master ( .q(_RegFile_reg_6__22__m2s), .d(
        n3531), .sdi(n2547), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_6__22__slave ( .q(_RegFile_6__22), .qb(n2548), .d(
        _RegFile_reg_6__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_6__23__master ( .q(_RegFile_reg_6__23__m2s), .d(
        n3532), .sdi(n2548), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n979), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_6__23__slave ( .q(_RegFile_6__23), .qb(n2549), .d(
        _RegFile_reg_6__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n979), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_6__24__master ( .q(_RegFile_reg_6__24__m2s), .d(
        n3533), .sdi(n2549), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_6__24__slave ( .q(_RegFile_6__24), .qb(n2550), .d(
        _RegFile_reg_6__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_6__25__master ( .q(_RegFile_reg_6__25__m2s), .d(
        n3534), .sdi(n2550), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n979), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_6__25__slave ( .q(_RegFile_6__25), .qb(n2551), .d(
        _RegFile_reg_6__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n979), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_6__26__master ( .q(_RegFile_reg_6__26__m2s), .d(
        n3535), .sdi(n2551), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_6__26__slave ( .q(_RegFile_6__26), .qb(n2552), .d(
        _RegFile_reg_6__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_6__27__master ( .q(_RegFile_reg_6__27__m2s), .d(
        n3536), .sdi(n2552), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n979), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_6__27__slave ( .q(_RegFile_6__27), .qb(n2553), .d(
        _RegFile_reg_6__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n979), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_6__28__master ( .q(_RegFile_reg_6__28__m2s), .d(
        n3537), .sdi(n2553), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_6__28__slave ( .q(_RegFile_6__28), .qb(n2554), .d(
        _RegFile_reg_6__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_6__29__master ( .q(_RegFile_reg_6__29__m2s), .d(
        n3538), .sdi(n2554), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n979), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_6__29__slave ( .q(_RegFile_6__29), .qb(n2555), .d(
        _RegFile_reg_6__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n979), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_6__2__master ( .q(_RegFile_reg_6__2__m2s), .d(n3511
        ), .sdi(n4319), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n979), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_6__2__slave ( .q(_RegFile_6__2), .qb(n4318), .d(
        _RegFile_reg_6__2__m2s), .g(Ctrl__Regs_1__en2), .rb(n979), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_6__30__master ( .q(_RegFile_reg_6__30__m2s), .d(
        n3539), .sdi(n2555), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n979), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_6__30__slave ( .q(_RegFile_6__30), .qb(n2556), .d(
        _RegFile_reg_6__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n979), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_6__31__master ( .q(_RegFile_reg_6__31__m2s), .d(
        n3540), .sdi(n2556), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_6__31__slave ( .q(_RegFile_6__31), .qb(n2557), .d(
        _RegFile_reg_6__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_6__3__master ( .q(_RegFile_reg_6__3__m2s), .d(n3512
        ), .sdi(n4318), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_6__3__slave ( .q(_RegFile_6__3), .qb(n4317), .d(
        _RegFile_reg_6__3__m2s), .g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_6__4__master ( .q(_RegFile_reg_6__4__m2s), .d(n3513
        ), .sdi(n4317), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n979), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_6__4__slave ( .q(_RegFile_6__4), .qb(n4316), .d(
        _RegFile_reg_6__4__m2s), .g(Ctrl__Regs_1__en2), .rb(n979), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_6__5__master ( .q(_RegFile_reg_6__5__m2s), .d(n3514
        ), .sdi(n4316), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n922), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_6__5__slave ( .q(_RegFile_6__5), .qb(n4315), .d(
        _RegFile_reg_6__5__m2s), .g(Ctrl__Regs_1__en2), .rb(n922), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_6__6__master ( .q(_RegFile_reg_6__6__m2s), .d(n3515
        ), .sdi(n4315), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n979), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_6__6__slave ( .q(_RegFile_6__6), .qb(n4314), .d(
        _RegFile_reg_6__6__m2s), .g(Ctrl__Regs_1__en2), .rb(n979), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_6__7__master ( .q(_RegFile_reg_6__7__m2s), .d(n3516
        ), .sdi(n4314), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n922), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_6__7__slave ( .q(_RegFile_6__7), .qb(n4313), .d(
        _RegFile_reg_6__7__m2s), .g(Ctrl__Regs_1__en2), .rb(n922), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_6__8__master ( .q(_RegFile_reg_6__8__m2s), .d(n3517
        ), .sdi(n4313), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n979), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_6__8__slave ( .q(_RegFile_6__8), .qb(n2558), .d(
        _RegFile_reg_6__8__m2s), .g(Ctrl__Regs_1__en2), .rb(n979), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_6__9__master ( .q(_RegFile_reg_6__9__m2s), .d(n3518
        ), .sdi(n2558), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n922), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_6__9__slave ( .q(_RegFile_6__9), .qb(n2559), .d(
        _RegFile_reg_6__9__m2s), .g(Ctrl__Regs_1__en2), .rb(n922), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_7__0__master ( .q(_RegFile_reg_7__0__m2s), .d(n3477
        ), .sdi(n2557), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n979), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_7__0__slave ( .q(_RegFile_7__0), .qb(n4312), .d(
        _RegFile_reg_7__0__m2s), .g(Ctrl__Regs_1__en2), .rb(n979), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_7__10__master ( .q(_RegFile_reg_7__10__m2s), .d(
        n3487), .sdi(n2583), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n979), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_7__10__slave ( .q(_RegFile_7__10), .qb(n2560), .d(
        _RegFile_reg_7__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n979), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_7__11__master ( .q(_RegFile_reg_7__11__m2s), .d(
        n3488), .sdi(n2560), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n922), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_7__11__slave ( .q(_RegFile_7__11), .qb(n2561), .d(
        _RegFile_reg_7__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n922), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_7__12__master ( .q(_RegFile_reg_7__12__m2s), .d(
        n3489), .sdi(n2561), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n979), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_7__12__slave ( .q(_RegFile_7__12), .qb(n2562), .d(
        _RegFile_reg_7__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n979), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_7__13__master ( .q(_RegFile_reg_7__13__m2s), .d(
        n3490), .sdi(n2562), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n922), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_7__13__slave ( .q(_RegFile_7__13), .qb(n2563), .d(
        _RegFile_reg_7__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n922), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_7__14__master ( .q(_RegFile_reg_7__14__m2s), .d(
        n3491), .sdi(n2563), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n979), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_7__14__slave ( .q(_RegFile_7__14), .qb(n2564), .d(
        _RegFile_reg_7__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n979), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_7__15__master ( .q(_RegFile_reg_7__15__m2s), .d(
        n3492), .sdi(n2564), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n922), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_7__15__slave ( .q(_RegFile_7__15), .qb(n2565), .d(
        _RegFile_reg_7__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n922), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_7__16__master ( .q(_RegFile_reg_7__16__m2s), .d(
        n3493), .sdi(n2565), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n979), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_7__16__slave ( .q(_RegFile_7__16), .qb(n2566), .d(
        _RegFile_reg_7__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n979), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_7__17__master ( .q(_RegFile_reg_7__17__m2s), .d(
        n3494), .sdi(n2566), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n922), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_7__17__slave ( .q(_RegFile_7__17), .qb(n2567), .d(
        _RegFile_reg_7__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n922), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_7__18__master ( .q(_RegFile_reg_7__18__m2s), .d(
        n3495), .sdi(n2567), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_7__18__slave ( .q(_RegFile_7__18), .qb(n2568), .d(
        _RegFile_reg_7__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_7__19__master ( .q(_RegFile_reg_7__19__m2s), .d(
        n3496), .sdi(n2568), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n922), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_7__19__slave ( .q(_RegFile_7__19), .qb(n2569), .d(
        _RegFile_reg_7__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n922), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_7__1__master ( .q(_RegFile_reg_7__1__m2s), .d(n3478
        ), .sdi(n4312), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n922), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_7__1__slave ( .q(_RegFile_7__1), .qb(n4311), .d(
        _RegFile_reg_7__1__m2s), .g(Ctrl__Regs_1__en2), .rb(n922), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_7__20__master ( .q(_RegFile_reg_7__20__m2s), .d(
        n3497), .sdi(n2569), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n922), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_7__20__slave ( .q(_RegFile_7__20), .qb(n2570), .d(
        _RegFile_reg_7__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n922), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_7__21__master ( .q(_RegFile_reg_7__21__m2s), .d(
        n3498), .sdi(n2570), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_7__21__slave ( .q(_RegFile_7__21), .qb(n2571), .d(
        _RegFile_reg_7__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_7__22__master ( .q(_RegFile_reg_7__22__m2s), .d(
        n3499), .sdi(n2571), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n922), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_7__22__slave ( .q(_RegFile_7__22), .qb(n2572), .d(
        _RegFile_reg_7__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n922), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_7__23__master ( .q(_RegFile_reg_7__23__m2s), .d(
        n3500), .sdi(n2572), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_7__23__slave ( .q(_RegFile_7__23), .qb(n2573), .d(
        _RegFile_reg_7__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_7__24__master ( .q(_RegFile_reg_7__24__m2s), .d(
        n3501), .sdi(n2573), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n922), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_7__24__slave ( .q(_RegFile_7__24), .qb(n2574), .d(
        _RegFile_reg_7__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n922), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_7__25__master ( .q(_RegFile_reg_7__25__m2s), .d(
        n3502), .sdi(n2574), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_7__25__slave ( .q(_RegFile_7__25), .qb(n2575), .d(
        _RegFile_reg_7__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_7__26__master ( .q(_RegFile_reg_7__26__m2s), .d(
        n3503), .sdi(n2575), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n922), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_7__26__slave ( .q(_RegFile_7__26), .qb(n2576), .d(
        _RegFile_reg_7__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n922), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_7__27__master ( .q(_RegFile_reg_7__27__m2s), .d(
        n3504), .sdi(n2576), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_7__27__slave ( .q(_RegFile_7__27), .qb(n2577), .d(
        _RegFile_reg_7__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_7__28__master ( .q(_RegFile_reg_7__28__m2s), .d(
        n3505), .sdi(n2577), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n922), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_7__28__slave ( .q(_RegFile_7__28), .qb(n2578), .d(
        _RegFile_reg_7__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n922), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_7__29__master ( .q(_RegFile_reg_7__29__m2s), .d(
        n3506), .sdi(n2578), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_7__29__slave ( .q(_RegFile_7__29), .qb(n2579), .d(
        _RegFile_reg_7__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_7__2__master ( .q(_RegFile_reg_7__2__m2s), .d(n3479
        ), .sdi(n4311), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_7__2__slave ( .q(_RegFile_7__2), .qb(n4310), .d(
        _RegFile_reg_7__2__m2s), .g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_7__30__master ( .q(_RegFile_reg_7__30__m2s), .d(
        n3507), .sdi(n2579), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_7__30__slave ( .q(_RegFile_7__30), .qb(n2580), .d(
        _RegFile_reg_7__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_7__31__master ( .q(_RegFile_reg_7__31__m2s), .d(
        n3508), .sdi(n2580), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n921), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_7__31__slave ( .q(_RegFile_7__31), .qb(n2581), .d(
        _RegFile_reg_7__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n921), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_7__3__master ( .q(_RegFile_reg_7__3__m2s), .d(n3480
        ), .sdi(n4310), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n922), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_7__3__slave ( .q(_RegFile_7__3), .qb(n4309), .d(
        _RegFile_reg_7__3__m2s), .g(Ctrl__Regs_1__en2), .rb(n922), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_7__4__master ( .q(_RegFile_reg_7__4__m2s), .d(n3481
        ), .sdi(n4309), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_7__4__slave ( .q(_RegFile_7__4), .qb(n4308), .d(
        _RegFile_reg_7__4__m2s), .g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_7__5__master ( .q(_RegFile_reg_7__5__m2s), .d(n3482
        ), .sdi(n4308), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n921), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_7__5__slave ( .q(_RegFile_7__5), .qb(n4307), .d(
        _RegFile_reg_7__5__m2s), .g(Ctrl__Regs_1__en2), .rb(n921), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_7__6__master ( .q(_RegFile_reg_7__6__m2s), .d(n3483
        ), .sdi(n4307), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_7__6__slave ( .q(_RegFile_7__6), .qb(n4306), .d(
        _RegFile_reg_7__6__m2s), .g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_7__7__master ( .q(_RegFile_reg_7__7__m2s), .d(n3484
        ), .sdi(n4306), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n921), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_7__7__slave ( .q(_RegFile_7__7), .qb(n4305), .d(
        _RegFile_reg_7__7__m2s), .g(Ctrl__Regs_1__en2), .rb(n921), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_7__8__master ( .q(_RegFile_reg_7__8__m2s), .d(n3485
        ), .sdi(n4305), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_7__8__slave ( .q(_RegFile_7__8), .qb(n2582), .d(
        _RegFile_reg_7__8__m2s), .g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_7__9__master ( .q(_RegFile_reg_7__9__m2s), .d(n3486
        ), .sdi(n2582), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n921), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_7__9__slave ( .q(_RegFile_7__9), .qb(n2583), .d(
        _RegFile_reg_7__9__m2s), .g(Ctrl__Regs_1__en2), .rb(n921), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_8__0__master ( .q(_RegFile_reg_8__0__m2s), .d(n3445
        ), .sdi(n2581), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_8__0__slave ( .q(_RegFile_8__0), .qb(n4304), .d(
        _RegFile_reg_8__0__m2s), .g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_8__10__master ( .q(_RegFile_reg_8__10__m2s), .d(
        n3455), .sdi(n2607), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_8__10__slave ( .q(_RegFile_8__10), .qb(n2584), .d(
        _RegFile_reg_8__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_8__11__master ( .q(_RegFile_reg_8__11__m2s), .d(
        n3456), .sdi(n2584), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n921), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_8__11__slave ( .q(_RegFile_8__11), .qb(n2585), .d(
        _RegFile_reg_8__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n921), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_8__12__master ( .q(_RegFile_reg_8__12__m2s), .d(
        n3457), .sdi(n2585), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_8__12__slave ( .q(_RegFile_8__12), .qb(n2586), .d(
        _RegFile_reg_8__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_8__13__master ( .q(_RegFile_reg_8__13__m2s), .d(
        n3458), .sdi(n2586), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n921), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_8__13__slave ( .q(_RegFile_8__13), .qb(n2587), .d(
        _RegFile_reg_8__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n921), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_8__14__master ( .q(_RegFile_reg_8__14__m2s), .d(
        n3459), .sdi(n2587), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_8__14__slave ( .q(_RegFile_8__14), .qb(n2588), .d(
        _RegFile_reg_8__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_8__15__master ( .q(_RegFile_reg_8__15__m2s), .d(
        n3460), .sdi(n2588), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n921), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_8__15__slave ( .q(_RegFile_8__15), .qb(n2589), .d(
        _RegFile_reg_8__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n921), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_8__16__master ( .q(_RegFile_reg_8__16__m2s), .d(
        n3461), .sdi(n2589), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n980), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_8__16__slave ( .q(_RegFile_8__16), .qb(n2590), .d(
        _RegFile_reg_8__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n980), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_8__17__master ( .q(_RegFile_reg_8__17__m2s), .d(
        n3462), .sdi(n2590), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n921), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_8__17__slave ( .q(_RegFile_8__17), .qb(n2591), .d(
        _RegFile_reg_8__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n921), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_8__18__master ( .q(_RegFile_reg_8__18__m2s), .d(
        n3463), .sdi(n2591), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n980), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_8__18__slave ( .q(_RegFile_8__18), .qb(n2592), .d(
        _RegFile_reg_8__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n980), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_8__19__master ( .q(_RegFile_reg_8__19__m2s), .d(
        n3464), .sdi(n2592), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n921), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_8__19__slave ( .q(_RegFile_8__19), .qb(n2593), .d(
        _RegFile_reg_8__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n921), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_8__1__master ( .q(_RegFile_reg_8__1__m2s), .d(n3446
        ), .sdi(n4304), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n921), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_8__1__slave ( .q(_RegFile_8__1), .qb(n4303), .d(
        _RegFile_reg_8__1__m2s), .g(Ctrl__Regs_1__en2), .rb(n921), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_8__20__master ( .q(_RegFile_reg_8__20__m2s), .d(
        n3465), .sdi(n2593), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n921), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_8__20__slave ( .q(_RegFile_8__20), .qb(n2594), .d(
        _RegFile_reg_8__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n921), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_8__21__master ( .q(_RegFile_reg_8__21__m2s), .d(
        n3466), .sdi(n2594), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n980), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_8__21__slave ( .q(_RegFile_8__21), .qb(n2595), .d(
        _RegFile_reg_8__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n980), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_8__22__master ( .q(_RegFile_reg_8__22__m2s), .d(
        n3467), .sdi(n2595), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n921), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_8__22__slave ( .q(_RegFile_8__22), .qb(n2596), .d(
        _RegFile_reg_8__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n921), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_8__23__master ( .q(_RegFile_reg_8__23__m2s), .d(
        n3468), .sdi(n2596), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n980), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_8__23__slave ( .q(_RegFile_8__23), .qb(n2597), .d(
        _RegFile_reg_8__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n980), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_8__24__master ( .q(_RegFile_reg_8__24__m2s), .d(
        n3469), .sdi(n2597), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n921), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_8__24__slave ( .q(_RegFile_8__24), .qb(n2598), .d(
        _RegFile_reg_8__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n921), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_8__25__master ( .q(_RegFile_reg_8__25__m2s), .d(
        n3470), .sdi(n2598), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n980), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_8__25__slave ( .q(_RegFile_8__25), .qb(n2599), .d(
        _RegFile_reg_8__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n980), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_8__26__master ( .q(_RegFile_reg_8__26__m2s), .d(
        n3471), .sdi(n2599), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n921), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_8__26__slave ( .q(_RegFile_8__26), .qb(n2600), .d(
        _RegFile_reg_8__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n921), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_8__27__master ( .q(_RegFile_reg_8__27__m2s), .d(
        n3472), .sdi(n2600), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n980), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_8__27__slave ( .q(_RegFile_8__27), .qb(n2601), .d(
        _RegFile_reg_8__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n980), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_8__28__master ( .q(_RegFile_reg_8__28__m2s), .d(
        n3473), .sdi(n2601), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n921), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_8__28__slave ( .q(_RegFile_8__28), .qb(n2602), .d(
        _RegFile_reg_8__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n921), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_8__29__master ( .q(_RegFile_reg_8__29__m2s), .d(
        n3474), .sdi(n2602), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n980), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_8__29__slave ( .q(_RegFile_8__29), .qb(n2603), .d(
        _RegFile_reg_8__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n980), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_8__2__master ( .q(_RegFile_reg_8__2__m2s), .d(n3447
        ), .sdi(n4303), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n980), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_8__2__slave ( .q(_RegFile_8__2), .qb(n4302), .d(
        _RegFile_reg_8__2__m2s), .g(Ctrl__Regs_1__en2), .rb(n980), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_8__30__master ( .q(_RegFile_reg_8__30__m2s), .d(
        n3475), .sdi(n2603), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n980), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_8__30__slave ( .q(_RegFile_8__30), .qb(n2604), .d(
        _RegFile_reg_8__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n980), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_8__31__master ( .q(_RegFile_reg_8__31__m2s), .d(
        n3476), .sdi(n2604), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n920), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_8__31__slave ( .q(_RegFile_8__31), .qb(n2605), .d(
        _RegFile_reg_8__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n920), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_8__3__master ( .q(_RegFile_reg_8__3__m2s), .d(n3448
        ), .sdi(n4302), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n920), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_8__3__slave ( .q(_RegFile_8__3), .qb(n4301), .d(
        _RegFile_reg_8__3__m2s), .g(Ctrl__Regs_1__en2), .rb(n920), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_8__4__master ( .q(_RegFile_reg_8__4__m2s), .d(n3449
        ), .sdi(n4301), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n980), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_8__4__slave ( .q(_RegFile_8__4), .qb(n4300), .d(
        _RegFile_reg_8__4__m2s), .g(Ctrl__Regs_1__en2), .rb(n980), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_8__5__master ( .q(_RegFile_reg_8__5__m2s), .d(n3450
        ), .sdi(n4300), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n920), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_8__5__slave ( .q(_RegFile_8__5), .qb(n4299), .d(
        _RegFile_reg_8__5__m2s), .g(Ctrl__Regs_1__en2), .rb(n920), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_8__6__master ( .q(_RegFile_reg_8__6__m2s), .d(n3451
        ), .sdi(n4299), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n980), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_8__6__slave ( .q(_RegFile_8__6), .qb(n4298), .d(
        _RegFile_reg_8__6__m2s), .g(Ctrl__Regs_1__en2), .rb(n980), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_8__7__master ( .q(_RegFile_reg_8__7__m2s), .d(n3452
        ), .sdi(n4298), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n920), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_8__7__slave ( .q(_RegFile_8__7), .qb(n4297), .d(
        _RegFile_reg_8__7__m2s), .g(Ctrl__Regs_1__en2), .rb(n920), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_8__8__master ( .q(_RegFile_reg_8__8__m2s), .d(n3453
        ), .sdi(n4297), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n980), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_8__8__slave ( .q(_RegFile_8__8), .qb(n2606), .d(
        _RegFile_reg_8__8__m2s), .g(Ctrl__Regs_1__en2), .rb(n980), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_8__9__master ( .q(_RegFile_reg_8__9__m2s), .d(n3454
        ), .sdi(n2606), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n920), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_8__9__slave ( .q(_RegFile_8__9), .qb(n2607), .d(
        _RegFile_reg_8__9__m2s), .g(Ctrl__Regs_1__en2), .rb(n920), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_9__0__master ( .q(_RegFile_reg_9__0__m2s), .d(n3413
        ), .sdi(n2605), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n980), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_9__0__slave ( .q(_RegFile_9__0), .qb(n4296), .d(
        _RegFile_reg_9__0__m2s), .g(Ctrl__Regs_1__en2), .rb(n980), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_9__10__master ( .q(_RegFile_reg_9__10__m2s), .d(
        n3423), .sdi(n2631), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n980), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_9__10__slave ( .q(_RegFile_9__10), .qb(n2608), .d(
        _RegFile_reg_9__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n980), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_9__11__master ( .q(_RegFile_reg_9__11__m2s), .d(
        n3424), .sdi(n2608), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n920), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_9__11__slave ( .q(_RegFile_9__11), .qb(n2609), .d(
        _RegFile_reg_9__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n920), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_9__12__master ( .q(_RegFile_reg_9__12__m2s), .d(
        n3425), .sdi(n2609), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n980), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_9__12__slave ( .q(_RegFile_9__12), .qb(n2610), .d(
        _RegFile_reg_9__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n980), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_9__13__master ( .q(_RegFile_reg_9__13__m2s), .d(
        n3426), .sdi(n2610), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n920), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_9__13__slave ( .q(_RegFile_9__13), .qb(n2611), .d(
        _RegFile_reg_9__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n920), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_9__14__master ( .q(_RegFile_reg_9__14__m2s), .d(
        n3427), .sdi(n2611), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_9__14__slave ( .q(_RegFile_9__14), .qb(n2612), .d(
        _RegFile_reg_9__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_9__15__master ( .q(_RegFile_reg_9__15__m2s), .d(
        n3428), .sdi(n2612), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n920), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_9__15__slave ( .q(_RegFile_9__15), .qb(n2613), .d(
        _RegFile_reg_9__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n920), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_9__16__master ( .q(_RegFile_reg_9__16__m2s), .d(
        n3429), .sdi(n2613), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_9__16__slave ( .q(_RegFile_9__16), .qb(n2614), .d(
        _RegFile_reg_9__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_9__17__master ( .q(_RegFile_reg_9__17__m2s), .d(
        n3430), .sdi(n2614), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n920), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_9__17__slave ( .q(_RegFile_9__17), .qb(n2615), .d(
        _RegFile_reg_9__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n920), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_9__18__master ( .q(_RegFile_reg_9__18__m2s), .d(
        n3431), .sdi(n2615), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_9__18__slave ( .q(_RegFile_9__18), .qb(n2616), .d(
        _RegFile_reg_9__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_9__19__master ( .q(_RegFile_reg_9__19__m2s), .d(
        n3432), .sdi(n2616), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n920), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_9__19__slave ( .q(_RegFile_9__19), .qb(n2617), .d(
        _RegFile_reg_9__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n920), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_9__1__master ( .q(_RegFile_reg_9__1__m2s), .d(n3414
        ), .sdi(n4296), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n920), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_9__1__slave ( .q(_RegFile_9__1), .qb(n4295), .d(
        _RegFile_reg_9__1__m2s), .g(Ctrl__Regs_1__en2), .rb(n920), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_9__20__master ( .q(_RegFile_reg_9__20__m2s), .d(
        n3433), .sdi(n2617), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n920), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_9__20__slave ( .q(_RegFile_9__20), .qb(n2618), .d(
        _RegFile_reg_9__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n920), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_9__21__master ( .q(_RegFile_reg_9__21__m2s), .d(
        n3434), .sdi(n2618), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_9__21__slave ( .q(_RegFile_9__21), .qb(n2619), .d(
        _RegFile_reg_9__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_9__22__master ( .q(_RegFile_reg_9__22__m2s), .d(
        n3435), .sdi(n2619), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n920), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_9__22__slave ( .q(_RegFile_9__22), .qb(n2620), .d(
        _RegFile_reg_9__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n920), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_9__23__master ( .q(_RegFile_reg_9__23__m2s), .d(
        n3436), .sdi(n2620), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_9__23__slave ( .q(_RegFile_9__23), .qb(n2621), .d(
        _RegFile_reg_9__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_9__24__master ( .q(_RegFile_reg_9__24__m2s), .d(
        n3437), .sdi(n2621), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n920), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_9__24__slave ( .q(_RegFile_9__24), .qb(n2622), .d(
        _RegFile_reg_9__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n920), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_9__25__master ( .q(_RegFile_reg_9__25__m2s), .d(
        n3438), .sdi(n2622), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_9__25__slave ( .q(_RegFile_9__25), .qb(n2623), .d(
        _RegFile_reg_9__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_9__26__master ( .q(_RegFile_reg_9__26__m2s), .d(
        n3439), .sdi(n2623), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n920), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_9__26__slave ( .q(_RegFile_9__26), .qb(n2624), .d(
        _RegFile_reg_9__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n920), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_9__27__master ( .q(_RegFile_reg_9__27__m2s), .d(
        n3440), .sdi(n2624), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_9__27__slave ( .q(_RegFile_9__27), .qb(n2625), .d(
        _RegFile_reg_9__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_9__28__master ( .q(_RegFile_reg_9__28__m2s), .d(
        n3441), .sdi(n2625), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n919), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_9__28__slave ( .q(_RegFile_9__28), .qb(n2626), .d(
        _RegFile_reg_9__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n919), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_9__29__master ( .q(_RegFile_reg_9__29__m2s), .d(
        n3442), .sdi(n2626), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_9__29__slave ( .q(_RegFile_9__29), .qb(n2627), .d(
        _RegFile_reg_9__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_9__2__master ( .q(_RegFile_reg_9__2__m2s), .d(n3415
        ), .sdi(n4295), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_9__2__slave ( .q(_RegFile_9__2), .qb(n4294), .d(
        _RegFile_reg_9__2__m2s), .g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_9__30__master ( .q(_RegFile_reg_9__30__m2s), .d(
        n3443), .sdi(n2627), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_9__30__slave ( .q(_RegFile_9__30), .qb(n2628), .d(
        _RegFile_reg_9__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_9__31__master ( .q(_RegFile_reg_9__31__m2s), .d(
        n3444), .sdi(n2628), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n919), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_9__31__slave ( .q(_RegFile_9__31), .qb(n2629), .d(
        _RegFile_reg_9__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n919), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_9__3__master ( .q(_RegFile_reg_9__3__m2s), .d(n3416
        ), .sdi(n4294), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n919), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_9__3__slave ( .q(_RegFile_9__3), .qb(n4293), .d(
        _RegFile_reg_9__3__m2s), .g(Ctrl__Regs_1__en2), .rb(n919), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_9__4__master ( .q(_RegFile_reg_9__4__m2s), .d(n3417
        ), .sdi(n4293), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_9__4__slave ( .q(_RegFile_9__4), .qb(n4292), .d(
        _RegFile_reg_9__4__m2s), .g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_9__5__master ( .q(_RegFile_reg_9__5__m2s), .d(n3418
        ), .sdi(n4292), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n919), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_9__5__slave ( .q(_RegFile_9__5), .qb(n4291), .d(
        _RegFile_reg_9__5__m2s), .g(Ctrl__Regs_1__en2), .rb(n919), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_9__6__master ( .q(_RegFile_reg_9__6__m2s), .d(n3419
        ), .sdi(n4291), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_9__6__slave ( .q(_RegFile_9__6), .qb(n4290), .d(
        _RegFile_reg_9__6__m2s), .g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_9__7__master ( .q(_RegFile_reg_9__7__m2s), .d(n3420
        ), .sdi(n4290), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n919), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_9__7__slave ( .q(_RegFile_9__7), .qb(n4289), .d(
        _RegFile_reg_9__7__m2s), .g(Ctrl__Regs_1__en2), .rb(n919), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_9__8__master ( .q(_RegFile_reg_9__8__m2s), .d(n3421
        ), .sdi(n4289), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_9__8__slave ( .q(_RegFile_9__8), .qb(n2630), .d(
        _RegFile_reg_9__8__m2s), .g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 _RegFile_reg_9__9__master ( .q(_RegFile_reg_9__9__m2s), .d(n3422
        ), .sdi(n2630), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n919), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 _RegFile_reg_9__9__slave ( .q(_RegFile_9__9), .qb(n2631), .d(
        _RegFile_reg_9__9__m2s), .g(Ctrl__Regs_1__en2), .rb(n919), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    ID_DW01_sub_32_2_test_1 add_489 ( .A({NPC[31], NPC[30], NPC[29], NPC[28], 
        NPC[27], NPC[26], NPC[25], NPC[24], NPC[23], NPC[22], NPC[21], NPC[20], 
        NPC[19], NPC[18], NPC[17], NPC[16], NPC[15], NPC[14], NPC[13], NPC[12], 
        NPC[11], NPC[10], NPC[9], NPC[8], NPC[7], NPC[6], NPC[5], NPC[4], 
        NPC[3], n737, NPC[1], NPC[0]}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 
        1'b0, 1'b0}), .CI(1'b0), .DIFF({N5350, N5349, N5348, N5347, N5346, 
        N5345, N5344, N5343, N5342, N5341, N5340, N5339, N5338, N5337, N5336, 
        N5335, N5334, N5333, N5332, N5331, N5330, N5329, N5328, N5327, N5326, 
        N5325, N5324, N5323, N5322, N5321, N5320, N5319}) );
    ID_DW01_sub_32_0_test_1 add_609 ( .A(NPC), .B({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b1, 1'b0, 1'b0}), .CI(1'b0), .DIFF({N5418, N5417, N5416, N5415, 
        N5414, N5413, N5412, N5411, N5410, N5409, N5408, N5407, N5406, N5405, 
        N5404, N5403, N5402, N5401, N5400, N5399, N5398, N5397, N5396, N5395, 
        N5394, N5393, N5392, N5391, N5390, N5389, N5388, N5387}) );
    ID_DW01_sub_32_1_test_1 add_779 ( .A({NPC[31], NPC[30], NPC[29], NPC[28], 
        NPC[27], NPC[26], NPC[25], NPC[24], NPC[23], NPC[22], NPC[21], NPC[20], 
        NPC[19], NPC[18], NPC[17], NPC[16], NPC[15], NPC[14], NPC[13], NPC[12], 
        NPC[11], NPC[10], NPC[9], NPC[8], NPC[7], NPC[6], NPC[5], NPC[4], n811, 
        n866, NPC[1], NPC[0]}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 
        1'b0}), .CI(1'b0), .DIFF({N6017, N6016, N6015, N6014, N6013, N6012, 
        N6011, N6010, N6009, N6008, N6007, N6006, N6005, N6004, N6003, N6002, 
        N6001, N6000, N5999, N5998, N5997, N5996, N5995, N5994, N5993, N5992, 
        N5991, N5990, N5989, N5988, N5987, N5986}) );
    smlatnr_2 branch_address_reg_0__master ( .q(branch_address_reg_0__m2s), 
        .d(n3824), .sdi(WB_index_4), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(
        n969), .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_8 branch_address_reg_0__slave ( .q(branch_address[0]), .qb(n4112), 
        .d(branch_address_reg_0__m2s), .g(Ctrl__Regs_1__en2), .rb(n969), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_2 branch_address_reg_10__master ( .q(branch_address_reg_10__m2s), 
        .d(n3834), .sdi(n4104), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_8 branch_address_reg_10__slave ( .q(branch_address[10]), .qb(n4103), 
        .d(branch_address_reg_10__m2s), .g(Ctrl__Regs_1__en2), .rb(n969), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_2 branch_address_reg_11__master ( .q(branch_address_reg_11__m2s), 
        .d(n3835), .sdi(n4103), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n919), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_8 branch_address_reg_11__slave ( .q(branch_address[11]), .qb(n4102), 
        .d(branch_address_reg_11__m2s), .g(Ctrl__Regs_1__en2), .rb(n919), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_2 branch_address_reg_12__master ( .q(branch_address_reg_12__m2s), 
        .d(n3836), .sdi(n4102), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n981), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_8 branch_address_reg_12__slave ( .q(branch_address[12]), .qb(n4101), 
        .d(branch_address_reg_12__m2s), .g(Ctrl__Regs_1__en2), .rb(n981), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_2 branch_address_reg_13__master ( .q(branch_address_reg_13__m2s), 
        .d(n3837), .sdi(n4101), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n919), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_8 branch_address_reg_13__slave ( .q(branch_address[13]), .qb(n4100), 
        .d(branch_address_reg_13__m2s), .g(Ctrl__Regs_1__en2), .rb(n919), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_2 branch_address_reg_14__master ( .q(branch_address_reg_14__m2s), 
        .d(n3838), .sdi(n4100), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n981), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_8 branch_address_reg_14__slave ( .q(branch_address[14]), .qb(n4099), 
        .d(branch_address_reg_14__m2s), .g(Ctrl__Regs_1__en2), .rb(n981), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_1 branch_address_reg_15__master ( .q(branch_address_reg_15__m2s), 
        .d(n3839), .sdi(n4099), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n919), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 branch_address_reg_15__slave ( .q(branch_address[15]), .qb(n4098), 
        .d(branch_address_reg_15__m2s), .g(Ctrl__Regs_1__en2), .rb(n919), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_2 branch_address_reg_16__master ( .q(branch_address_reg_16__m2s), 
        .d(n3840), .sdi(n4098), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n981), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_8 branch_address_reg_16__slave ( .q(branch_address[16]), .qb(n4097), 
        .d(branch_address_reg_16__m2s), .g(Ctrl__Regs_1__en2), .rb(n981), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_2 branch_address_reg_17__master ( .q(branch_address_reg_17__m2s), 
        .d(n3841), .sdi(n4097), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n919), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_8 branch_address_reg_17__slave ( .q(branch_address[17]), .qb(n4096), 
        .d(branch_address_reg_17__m2s), .g(Ctrl__Regs_1__en2), .rb(n919), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_2 branch_address_reg_18__master ( .q(branch_address_reg_18__m2s), 
        .d(n3842), .sdi(n4096), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n981), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_8 branch_address_reg_18__slave ( .q(branch_address[18]), .qb(n4095), 
        .d(branch_address_reg_18__m2s), .g(Ctrl__Regs_1__en2), .rb(n981), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_2 branch_address_reg_19__master ( .q(branch_address_reg_19__m2s), 
        .d(n3843), .sdi(n4095), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n919), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_8 branch_address_reg_19__slave ( .q(branch_address[19]), .qb(n4094), 
        .d(branch_address_reg_19__m2s), .g(Ctrl__Regs_1__en2), .rb(n919), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_1 branch_address_reg_1__master ( .q(branch_address_reg_1__m2s), 
        .d(n3825), .sdi(n4112), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n919), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 branch_address_reg_1__slave ( .q(branch_address[1]), .qb(n4111), 
        .d(branch_address_reg_1__m2s), .g(Ctrl__Regs_1__en2), .rb(n919), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_2 branch_address_reg_20__master ( .q(branch_address_reg_20__m2s), 
        .d(n3844), .sdi(n4094), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n919), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_8 branch_address_reg_20__slave ( .q(branch_address[20]), .qb(n4093), 
        .d(branch_address_reg_20__m2s), .g(Ctrl__Regs_1__en2), .rb(n919), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_2 branch_address_reg_21__master ( .q(branch_address_reg_21__m2s), 
        .d(n3845), .sdi(n4093), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n981), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_8 branch_address_reg_21__slave ( .q(branch_address[21]), .qb(n4092), 
        .d(branch_address_reg_21__m2s), .g(Ctrl__Regs_1__en2), .rb(n981), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_2 branch_address_reg_22__master ( .q(branch_address_reg_22__m2s), 
        .d(n3846), .sdi(n4092), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n919), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_8 branch_address_reg_22__slave ( .q(branch_address[22]), .qb(n4091), 
        .d(branch_address_reg_22__m2s), .g(Ctrl__Regs_1__en2), .rb(n919), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_2 branch_address_reg_23__master ( .q(branch_address_reg_23__m2s), 
        .d(n3847), .sdi(n4091), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n981), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_8 branch_address_reg_23__slave ( .q(branch_address[23]), .qb(n4090), 
        .d(branch_address_reg_23__m2s), .g(Ctrl__Regs_1__en2), .rb(n981), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_2 branch_address_reg_24__master ( .q(branch_address_reg_24__m2s), 
        .d(n3848), .sdi(n4090), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n919), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_8 branch_address_reg_24__slave ( .q(branch_address[24]), .qb(n4089), 
        .d(branch_address_reg_24__m2s), .g(Ctrl__Regs_1__en2), .rb(n919), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_2 branch_address_reg_25__master ( .q(branch_address_reg_25__m2s), 
        .d(n3849), .sdi(n4089), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n981), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_8 branch_address_reg_25__slave ( .q(branch_address[25]), .qb(n4088), 
        .d(branch_address_reg_25__m2s), .g(Ctrl__Regs_1__en2), .rb(n981), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_2 branch_address_reg_26__master ( .q(branch_address_reg_26__m2s), 
        .d(n3850), .sdi(n4088), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n918), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_8 branch_address_reg_26__slave ( .q(branch_address[26]), .qb(n4087), 
        .d(branch_address_reg_26__m2s), .g(Ctrl__Regs_1__en2), .rb(n918), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_1 branch_address_reg_27__master ( .q(branch_address_reg_27__m2s), 
        .d(n3851), .sdi(n4087), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n981), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 branch_address_reg_27__slave ( .q(branch_address[27]), .qb(n4086), 
        .d(branch_address_reg_27__m2s), .g(Ctrl__Regs_1__en2), .rb(n981), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_2 branch_address_reg_28__master ( .q(branch_address_reg_28__m2s), 
        .d(n3852), .sdi(n4086), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n918), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_8 branch_address_reg_28__slave ( .q(branch_address[28]), .qb(n4085), 
        .d(branch_address_reg_28__m2s), .g(Ctrl__Regs_1__en2), .rb(n918), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_2 branch_address_reg_29__master ( .q(branch_address_reg_29__m2s), 
        .d(n3853), .sdi(n4085), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n981), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_8 branch_address_reg_29__slave ( .q(branch_address[29]), .qb(n4084), 
        .d(branch_address_reg_29__m2s), .g(Ctrl__Regs_1__en2), .rb(n981), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_2 branch_address_reg_2__master ( .q(branch_address_reg_2__m2s), 
        .d(n3826), .sdi(n4111), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n981), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_8 branch_address_reg_2__slave ( .q(branch_address[2]), .qb(n4110), 
        .d(branch_address_reg_2__m2s), .g(Ctrl__Regs_1__en2), .rb(n981), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_2 branch_address_reg_30__master ( .q(branch_address_reg_30__m2s), 
        .d(n3854), .sdi(n4084), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n981), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_8 branch_address_reg_30__slave ( .q(branch_address[30]), .qb(n4083), 
        .d(branch_address_reg_30__m2s), .g(Ctrl__Regs_1__en2), .rb(n981), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_2 branch_address_reg_31__master ( .q(branch_address_reg_31__m2s), 
        .d(_branch_address_reg_31_net46811), .sdi(n4083), .se(test_se), .g(
        Ctrl__Regs_1__en1), .rb(n918), .glob_g(global_g1), .sync_sel(sync_sel)
         );
    mlatnr_8 branch_address_reg_31__slave ( .q(branch_address[31]), .qb(n2632), 
        .d(branch_address_reg_31__m2s), .g(Ctrl__Regs_1__en2), .rb(n918), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_2 branch_address_reg_3__master ( .q(branch_address_reg_3__m2s), 
        .d(n3827), .sdi(n4110), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n918), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_8 branch_address_reg_3__slave ( .q(branch_address[3]), .qb(n4109), 
        .d(branch_address_reg_3__m2s), .g(Ctrl__Regs_1__en2), .rb(n918), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_2 branch_address_reg_4__master ( .q(branch_address_reg_4__m2s), 
        .d(n3828), .sdi(n4109), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n981), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_8 branch_address_reg_4__slave ( .q(branch_address[4]), .qb(n4108), 
        .d(branch_address_reg_4__m2s), .g(Ctrl__Regs_1__en2), .rb(n981), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_2 branch_address_reg_5__master ( .q(branch_address_reg_5__m2s), 
        .d(n3829), .sdi(n4108), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n918), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_8 branch_address_reg_5__slave ( .q(branch_address[5]), .qb(n4107), 
        .d(branch_address_reg_5__m2s), .g(Ctrl__Regs_1__en2), .rb(n918), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_2 branch_address_reg_6__master ( .q(branch_address_reg_6__m2s), 
        .d(n3830), .sdi(n4107), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n981), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_8 branch_address_reg_6__slave ( .q(branch_address[6]), .qb(n4106), 
        .d(branch_address_reg_6__m2s), .g(Ctrl__Regs_1__en2), .rb(n981), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_2 branch_address_reg_7__master ( .q(branch_address_reg_7__m2s), 
        .d(n3831), .sdi(n4106), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n918), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_8 branch_address_reg_7__slave ( .q(branch_address[7]), .qb(n2633), 
        .d(branch_address_reg_7__m2s), .g(Ctrl__Regs_1__en2), .rb(n918), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_2 branch_address_reg_8__master ( .q(branch_address_reg_8__m2s), 
        .d(n3832), .sdi(branch_address[7]), .se(test_se), .g(Ctrl__Regs_1__en1
        ), .rb(n981), .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_8 branch_address_reg_8__slave ( .q(branch_address[8]), .qb(n4105), 
        .d(branch_address_reg_8__m2s), .g(Ctrl__Regs_1__en2), .rb(n981), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_2 branch_address_reg_9__master ( .q(branch_address_reg_9__m2s), 
        .d(n3833), .sdi(n4105), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n918), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_8 branch_address_reg_9__slave ( .q(branch_address[9]), .qb(n4104), 
        .d(branch_address_reg_9__m2s), .g(Ctrl__Regs_1__en2), .rb(n918), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_2 branch_sig_reg__master ( .q(branch_sig_reg__m2s), .d(n3823), 
        .sdi(branch_address[31]), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(
        n912), .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_8 branch_sig_reg__slave ( .q(branch_sig), .qb(n2634), .d(
        branch_sig_reg__m2s), .g(Ctrl__Regs_1__en2), .rb(n912), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 counter_reg_0__master ( .q(counter_reg_0__m2s), .d(
        _counter_reg_0_net48671), .sdi(n2634), .se(test_se), .g(
        Ctrl__Regs_1__en1), .rb(n916), .glob_g(global_g1), .sync_sel(sync_sel)
         );
    mlatnr_4 counter_reg_0__slave ( .q(n3950), .qb(n787), .d(
        counter_reg_0__m2s), .g(Ctrl__Regs_1__en2), .rb(n916), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 counter_reg_1__master ( .q(counter_reg_1__m2s), .d(
        _counter_reg_1_net48651), .sdi(counter[0]), .se(test_se), .g(
        Ctrl__Regs_1__en1), .rb(n916), .glob_g(global_g1), .sync_sel(sync_sel)
         );
    mlatnr_2 counter_reg_1__slave ( .q(n3949), .qb(n780), .d(
        counter_reg_1__m2s), .g(Ctrl__Regs_1__en2), .rb(n916), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 current_IR_reg_0__master ( .q(current_IR_reg_0__m2s), .d(n3733), 
        .sdi(n790), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n918), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 current_IR_reg_0__slave ( .q(current_IR_0), .qb(n4082), .d(
        current_IR_reg_0__m2s), .g(Ctrl__Regs_1__en2), .rb(n918), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 current_IR_reg_10__master ( .q(current_IR_reg_10__m2s), .d(n3742
        ), .sdi(n629), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n918), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 current_IR_reg_10__slave ( .q(current_IR_10), .qb(n632), .d(
        current_IR_reg_10__m2s), .g(Ctrl__Regs_1__en2), .rb(n918), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 current_IR_reg_11__master ( .q(current_IR_reg_11__m2s), .d(n3743
        ), .sdi(n632), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 current_IR_reg_11__slave ( .q(n4076), .qb(n571), .d(
        current_IR_reg_11__m2s), .g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 current_IR_reg_12__master ( .q(current_IR_reg_12__m2s), .d(n3744
        ), .sdi(n4076), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n918), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 current_IR_reg_12__slave ( .q(n4075), .qb(n652), .d(
        current_IR_reg_12__m2s), .g(Ctrl__Regs_1__en2), .rb(n918), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 current_IR_reg_13__master ( .q(current_IR_reg_13__m2s), .d(n3745
        ), .sdi(n4075), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 current_IR_reg_13__slave ( .q(n4074), .qb(n570), .d(
        current_IR_reg_13__m2s), .g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 current_IR_reg_14__master ( .q(current_IR_reg_14__m2s), .d(n3746
        ), .sdi(n4074), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n918), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 current_IR_reg_14__slave ( .q(n4073), .qb(n569), .d(
        current_IR_reg_14__m2s), .g(Ctrl__Regs_1__en2), .rb(n918), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 current_IR_reg_15__master ( .q(current_IR_reg_15__m2s), .d(n3747
        ), .sdi(n4073), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 current_IR_reg_15__slave ( .q(n4072), .qb(n568), .d(
        current_IR_reg_15__m2s), .g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 current_IR_reg_16__master ( .q(current_IR_reg_16__m2s), .d(n3748
        ), .sdi(n4072), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n918), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 current_IR_reg_16__slave ( .q(n644), .qb(n645), .d(
        current_IR_reg_16__m2s), .g(Ctrl__Regs_1__en2), .rb(n918), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 current_IR_reg_17__master ( .q(current_IR_reg_17__m2s), .d(n3749
        ), .sdi(n645), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 current_IR_reg_17__slave ( .q(current_IR_17), .qb(n4071), .d(
        current_IR_reg_17__m2s), .g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 current_IR_reg_18__master ( .q(current_IR_reg_18__m2s), .d(n3750
        ), .sdi(n4071), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n918), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 current_IR_reg_18__slave ( .q(current_IR_18), .qb(n4070), .d(
        current_IR_reg_18__m2s), .g(Ctrl__Regs_1__en2), .rb(n918), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 current_IR_reg_19__master ( .q(current_IR_reg_19__m2s), .d(n3751
        ), .sdi(n4070), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 current_IR_reg_19__slave ( .q(current_IR_19), .qb(n657), .d(
        current_IR_reg_19__m2s), .g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 current_IR_reg_1__master ( .q(current_IR_reg_1__m2s), .d(
        _current_IR_reg_1_net49291), .sdi(n4082), .se(test_se), .g(
        Ctrl__Regs_1__en1), .rb(n981), .glob_g(global_g1), .sync_sel(sync_sel)
         );
    mlatnr_2 current_IR_reg_1__slave ( .q(current_IR_1), .qb(n4081), .d(
        current_IR_reg_1__m2s), .g(Ctrl__Regs_1__en2), .rb(n981), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 current_IR_reg_20__master ( .q(current_IR_reg_20__m2s), .d(n3752
        ), .sdi(n657), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 current_IR_reg_20__slave ( .q(n4069), .qb(n567), .d(
        current_IR_reg_20__m2s), .g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 current_IR_reg_21__master ( .q(current_IR_reg_21__m2s), .d(n3753
        ), .sdi(n4069), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n918), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 current_IR_reg_21__slave ( .q(current_IR_21), .qb(n646), .d(
        current_IR_reg_21__m2s), .g(Ctrl__Regs_1__en2), .rb(n918), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 current_IR_reg_22__master ( .q(current_IR_reg_22__m2s), .d(n3754
        ), .sdi(n646), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n948), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 current_IR_reg_22__slave ( .q(n660), .qb(n661), .d(
        current_IR_reg_22__m2s), .g(Ctrl__Regs_1__en2), .rb(n948), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 current_IR_reg_23__master ( .q(current_IR_reg_23__m2s), .d(n3755
        ), .sdi(n661), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n917), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 current_IR_reg_23__slave ( .q(current_IR_23), .qb(n659), .d(
        current_IR_reg_23__m2s), .g(Ctrl__Regs_1__en2), .rb(n917), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 current_IR_reg_24__master ( .q(current_IR_reg_24__m2s), .d(n3756
        ), .sdi(n659), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 current_IR_reg_24__slave ( .q(current_IR_24), .qb(n4068), .d(
        current_IR_reg_24__m2s), .g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 current_IR_reg_25__master ( .q(current_IR_reg_25__m2s), .d(n3757
        ), .sdi(n4068), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n916), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 current_IR_reg_25__slave ( .q(n4067), .qb(n666), .d(
        current_IR_reg_25__m2s), .g(Ctrl__Regs_1__en2), .rb(n916), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 current_IR_reg_26__master ( .q(current_IR_reg_26__m2s), .d(n3758
        ), .sdi(n4067), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 current_IR_reg_26__slave ( .q(n4066), .qb(n852), .d(
        current_IR_reg_26__m2s), .g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 current_IR_reg_27__master ( .q(current_IR_reg_27__m2s), .d(n3759
        ), .sdi(n4066), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n917), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 current_IR_reg_27__slave ( .q(current_IR_27), .qb(n4065), .d(
        current_IR_reg_27__m2s), .g(Ctrl__Regs_1__en2), .rb(n917), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 current_IR_reg_28__master ( .q(current_IR_reg_28__m2s), .d(n3760
        ), .sdi(n4065), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 current_IR_reg_28__slave ( .q(n4064), .qb(n566), .d(
        current_IR_reg_28__m2s), .g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 current_IR_reg_29__master ( .q(current_IR_reg_29__m2s), .d(n3761
        ), .sdi(n4064), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n917), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 current_IR_reg_29__slave ( .q(current_IR_29), .qb(n656), .d(
        current_IR_reg_29__m2s), .g(Ctrl__Regs_1__en2), .rb(n917), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 current_IR_reg_2__master ( .q(current_IR_reg_2__m2s), .d(n3734), 
        .sdi(n4081), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n918), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 current_IR_reg_2__slave ( .q(current_IR_2), .qb(n4080), .d(
        current_IR_reg_2__m2s), .g(Ctrl__Regs_1__en2), .rb(n918), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 current_IR_reg_30__master ( .q(current_IR_reg_30__m2s), .d(n3762
        ), .sdi(n656), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n917), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 current_IR_reg_30__slave ( .q(current_IR_30), .qb(n658), .d(
        current_IR_reg_30__m2s), .g(Ctrl__Regs_1__en2), .rb(n917), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 current_IR_reg_31__master ( .q(current_IR_reg_31__m2s), .d(n3763
        ), .sdi(n658), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n948), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 current_IR_reg_31__slave ( .q(current_IR_31), .qb(n633), .d(
        current_IR_reg_31__m2s), .g(Ctrl__Regs_1__en2), .rb(n948), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 current_IR_reg_3__master ( .q(current_IR_reg_3__m2s), .d(n3735), 
        .sdi(n4080), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n948), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 current_IR_reg_3__slave ( .q(current_IR_3), .qb(n651), .d(
        current_IR_reg_3__m2s), .g(Ctrl__Regs_1__en2), .rb(n948), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 current_IR_reg_4__master ( .q(current_IR_reg_4__m2s), .d(n3736), 
        .sdi(n651), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n917), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 current_IR_reg_4__slave ( .q(current_IR_4), .qb(n4079), .d(
        current_IR_reg_4__m2s), .g(Ctrl__Regs_1__en2), .rb(n917), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 current_IR_reg_5__master ( .q(current_IR_reg_5__m2s), .d(n3737), 
        .sdi(n4079), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 current_IR_reg_5__slave ( .q(n4078), .qb(n565), .d(
        current_IR_reg_5__m2s), .g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 current_IR_reg_6__master ( .q(current_IR_reg_6__m2s), .d(n3738), 
        .sdi(n4078), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n917), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 current_IR_reg_6__slave ( .q(current_IR_6), .qb(n631), .d(
        current_IR_reg_6__m2s), .g(Ctrl__Regs_1__en2), .rb(n917), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 current_IR_reg_7__master ( .q(current_IR_reg_7__m2s), .d(n3739), 
        .sdi(n631), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 current_IR_reg_7__slave ( .q(current_IR_7), .qb(n4077), .d(
        current_IR_reg_7__m2s), .g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 current_IR_reg_8__master ( .q(current_IR_reg_8__m2s), .d(n3740), 
        .sdi(n4077), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n917), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 current_IR_reg_8__slave ( .q(current_IR_8), .qb(n630), .d(
        current_IR_reg_8__m2s), .g(Ctrl__Regs_1__en2), .rb(n917), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 current_IR_reg_9__master ( .q(current_IR_reg_9__m2s), .d(n3741), 
        .sdi(n630), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 current_IR_reg_9__slave ( .q(current_IR_9), .qb(n629), .d(
        current_IR_reg_9__m2s), .g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 delay_slot_reg__master ( .q(delay_slot_reg__m2s), .d(n2707), 
        .sdi(n633), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n917), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_4 delay_slot_reg__slave ( .q(delay_slot), .qb(n883), .d(
        delay_slot_reg__m2s), .g(Ctrl__Regs_1__en2), .rb(n917), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 intr_slot_reg__master ( .q(intr_slot_reg__m2s), .d(n2640), .sdi(
        n883), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 intr_slot_reg__slave ( .q(intr_slot), .qb(n564), .d(
        intr_slot_reg__m2s), .g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 mem_read_reg__master ( .q(mem_read_reg__m2s), .d(n3777), .sdi(
        intr_slot), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n917), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 mem_read_reg__slave ( .q(mem_read), .qb(n2635), .d(
        mem_read_reg__m2s), .g(Ctrl__Regs_1__en2), .rb(n917), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 mem_to_reg_reg__master ( .q(mem_to_reg_reg__m2s), .d(n3778), 
        .sdi(mem_read), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 mem_to_reg_reg__slave ( .q(mem_to_reg), .qb(n2636), .d(
        mem_to_reg_reg__m2s), .g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 mem_write_reg__master ( .q(mem_write_reg__m2s), .d(n3776), .sdi(
        mem_to_reg), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n917), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 mem_write_reg__slave ( .q(mem_write), .qb(n2637), .d(
        mem_write_reg__m2s), .g(Ctrl__Regs_1__en2), .rb(n917), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 opcode_of_MEM_reg_0__master ( .q(opcode_of_MEM_reg_0__m2s), .d(
        IR_opcode_field[0]), .sdi(mem_write), .se(test_se), .g(
        Ctrl__Regs_1__en1), .rb(n913), .glob_g(global_g1), .sync_sel(sync_sel)
         );
    mlatnr_2 opcode_of_MEM_reg_0__slave ( .q(opcode_of_MEM_0), .qb(n3924), .d(
        opcode_of_MEM_reg_0__m2s), .g(Ctrl__Regs_1__en2), .rb(n913), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 opcode_of_MEM_reg_1__master ( .q(opcode_of_MEM_reg_1__m2s), .d(
        IR_opcode_field[1]), .sdi(opcode_of_MEM_0), .se(test_se), .g(
        Ctrl__Regs_1__en1), .rb(n913), .glob_g(global_g1), .sync_sel(sync_sel)
         );
    mlatnr_2 opcode_of_MEM_reg_1__slave ( .q(opcode_of_MEM_1), .qb(n4063), .d(
        opcode_of_MEM_reg_1__m2s), .g(Ctrl__Regs_1__en2), .rb(n913), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 opcode_of_MEM_reg_2__master ( .q(opcode_of_MEM_reg_2__m2s), .d(
        IR_opcode_field[2]), .sdi(n4063), .se(test_se), .g(Ctrl__Regs_1__en1), 
        .rb(n913), .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 opcode_of_MEM_reg_2__slave ( .q(opcode_of_MEM_2), .qb(n3933), .d(
        opcode_of_MEM_reg_2__m2s), .g(Ctrl__Regs_1__en2), .rb(n913), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 opcode_of_MEM_reg_3__master ( .q(opcode_of_MEM_reg_3__m2s), .d(
        IR_opcode_field[3]), .sdi(n3933), .se(test_se), .g(Ctrl__Regs_1__en1), 
        .rb(n913), .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 opcode_of_MEM_reg_3__slave ( .q(opcode_of_MEM_3), .qb(n3932), .d(
        opcode_of_MEM_reg_3__m2s), .g(Ctrl__Regs_1__en2), .rb(n913), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 opcode_of_MEM_reg_4__master ( .q(opcode_of_MEM_reg_4__m2s), .d(
        IR_opcode_field[4]), .sdi(opcode_of_MEM_3), .se(test_se), .g(
        Ctrl__Regs_1__en1), .rb(n911), .glob_g(global_g1), .sync_sel(sync_sel)
         );
    mlatnr_4 opcode_of_MEM_reg_4__slave ( .q(opcode_of_MEM_4), .qb(n4062), .d(
        opcode_of_MEM_reg_4__m2s), .g(Ctrl__Regs_1__en2), .rb(n911), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 opcode_of_MEM_reg_5__master ( .q(opcode_of_MEM_reg_5__m2s), .d(
        IR_opcode_field[5]), .sdi(n4062), .se(test_se), .g(Ctrl__Regs_1__en1), 
        .rb(n913), .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 opcode_of_MEM_reg_5__slave ( .q(opcode_of_MEM_5), .qb(n4061), .d(
        opcode_of_MEM_reg_5__m2s), .g(Ctrl__Regs_1__en2), .rb(n913), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 opcode_of_WB_reg_0__master ( .q(opcode_of_WB_reg_0__m2s), .d(
        opcode_of_MEM_0), .sdi(n4061), .se(test_se), .g(Ctrl__Regs_1__en1), 
        .rb(n912), .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 opcode_of_WB_reg_0__slave ( .q(N13832), .qb(n4060), .d(
        opcode_of_WB_reg_0__m2s), .g(Ctrl__Regs_1__en2), .rb(n912), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 opcode_of_WB_reg_1__master ( .q(opcode_of_WB_reg_1__m2s), .d(
        opcode_of_MEM_1), .sdi(n4060), .se(test_se), .g(Ctrl__Regs_1__en1), 
        .rb(n912), .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 opcode_of_WB_reg_1__slave ( .q(n4059), .qb(n3887), .d(
        opcode_of_WB_reg_1__m2s), .g(Ctrl__Regs_1__en2), .rb(n912), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 opcode_of_WB_reg_2__master ( .q(opcode_of_WB_reg_2__m2s), .d(
        opcode_of_MEM_2), .sdi(n4059), .se(test_se), .g(Ctrl__Regs_1__en1), 
        .rb(n912), .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 opcode_of_WB_reg_2__slave ( .q(n3888), .qb(n4058), .d(
        opcode_of_WB_reg_2__m2s), .g(Ctrl__Regs_1__en2), .rb(n912), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 opcode_of_WB_reg_3__master ( .q(opcode_of_WB_reg_3__m2s), .d(
        opcode_of_MEM_3), .sdi(n4058), .se(test_se), .g(Ctrl__Regs_1__en1), 
        .rb(n912), .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 opcode_of_WB_reg_3__slave ( .q(n4057), .qb(n3889), .d(
        opcode_of_WB_reg_3__m2s), .g(Ctrl__Regs_1__en2), .rb(n912), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 opcode_of_WB_reg_4__master ( .q(opcode_of_WB_reg_4__m2s), .d(
        opcode_of_MEM_4), .sdi(n4057), .se(test_se), .g(Ctrl__Regs_1__en1), 
        .rb(n912), .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 opcode_of_WB_reg_4__slave ( .q(n4056), .qb(n3890), .d(
        opcode_of_WB_reg_4__m2s), .g(Ctrl__Regs_1__en2), .rb(n912), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 opcode_of_WB_reg_5__master ( .q(opcode_of_WB_reg_5__m2s), .d(
        opcode_of_MEM_5), .sdi(n4056), .se(test_se), .g(Ctrl__Regs_1__en1), 
        .rb(n913), .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 opcode_of_WB_reg_5__slave ( .q(opcode_of_WB_5), .qb(n4055), .d(
        opcode_of_WB_reg_5__m2s), .g(Ctrl__Regs_1__en2), .rb(n913), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 rd_addr_reg_0__master ( .q(rd_addr_reg_0__m2s), .d(n3781), .sdi(
        n4055), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 rd_addr_reg_0__slave ( .q(rd_addr[0]), .qb(n669), .d(
        rd_addr_reg_0__m2s), .g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 rd_addr_reg_1__master ( .q(rd_addr_reg_1__m2s), .d(n3782), .sdi(
        rd_addr[0]), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n917), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 rd_addr_reg_1__slave ( .q(rd_addr[1]), .qb(n563), .d(
        rd_addr_reg_1__m2s), .g(Ctrl__Regs_1__en2), .rb(n917), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 rd_addr_reg_2__master ( .q(rd_addr_reg_2__m2s), .d(n3783), .sdi(
        rd_addr[1]), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 rd_addr_reg_2__slave ( .q(rd_addr[2]), .qb(n670), .d(
        rd_addr_reg_2__m2s), .g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 rd_addr_reg_3__master ( .q(rd_addr_reg_3__m2s), .d(n3784), .sdi(
        rd_addr[2]), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n917), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 rd_addr_reg_3__slave ( .q(rd_addr[3]), .qb(n4054), .d(
        rd_addr_reg_3__m2s), .g(Ctrl__Regs_1__en2), .rb(n917), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 rd_addr_reg_4__master ( .q(rd_addr_reg_4__m2s), .d(n3785), .sdi(
        n4054), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 rd_addr_reg_4__slave ( .q(rd_addr[4]), .qb(n562), .d(
        rd_addr_reg_4__m2s), .g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_dst_of_MEM_reg_0__master ( .q(reg_dst_of_MEM_reg_0__m2s), 
        .d(reg_dst_of_EX_0), .sdi(rd_addr[4]), .se(test_se), .g(
        Ctrl__Regs_1__en1), .rb(n913), .glob_g(global_g1), .sync_sel(sync_sel)
         );
    mlatnr_2 reg_dst_of_MEM_reg_0__slave ( .q(reg_dst_of_MEM_0), .qb(n4053), 
        .d(reg_dst_of_MEM_reg_0__m2s), .g(Ctrl__Regs_1__en2), .rb(n913), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_dst_of_MEM_reg_1__master ( .q(reg_dst_of_MEM_reg_1__m2s), 
        .d(reg_dst_of_EX_1), .sdi(n4053), .se(test_se), .g(Ctrl__Regs_1__en1), 
        .rb(n913), .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_1 reg_dst_of_MEM_reg_1__slave ( .q(reg_dst_of_MEM_1), .qb(n4052), 
        .d(reg_dst_of_MEM_reg_1__m2s), .g(Ctrl__Regs_1__en2), .rb(n913), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_dst_of_MEM_reg_2__master ( .q(reg_dst_of_MEM_reg_2__m2s), 
        .d(reg_dst_of_EX_2), .sdi(n4052), .se(test_se), .g(Ctrl__Regs_1__en1), 
        .rb(n913), .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 reg_dst_of_MEM_reg_2__slave ( .q(reg_dst_of_MEM_2), .qb(n655), 
        .d(reg_dst_of_MEM_reg_2__m2s), .g(Ctrl__Regs_1__en2), .rb(n913), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_dst_of_MEM_reg_3__master ( .q(reg_dst_of_MEM_reg_3__m2s), 
        .d(reg_dst_of_EX_3), .sdi(reg_dst_of_MEM_2), .se(test_se), .g(
        Ctrl__Regs_1__en1), .rb(n914), .glob_g(global_g1), .sync_sel(sync_sel)
         );
    mlatnr_2 reg_dst_of_MEM_reg_3__slave ( .q(reg_dst_of_MEM_3), .qb(n634), 
        .d(reg_dst_of_MEM_reg_3__m2s), .g(Ctrl__Regs_1__en2), .rb(n914), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_dst_of_MEM_reg_4__master ( .q(reg_dst_of_MEM_reg_4__m2s), 
        .d(reg_dst_of_EX_4), .sdi(reg_dst_of_MEM_3), .se(test_se), .g(
        Ctrl__Regs_1__en1), .rb(n914), .glob_g(global_g1), .sync_sel(sync_sel)
         );
    mlatnr_2 reg_dst_of_MEM_reg_4__slave ( .q(reg_dst_of_MEM_4), .qb(n635), 
        .d(reg_dst_of_MEM_reg_4__m2s), .g(Ctrl__Regs_1__en2), .rb(n914), 
        .glob_g(global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_dst_reg__master ( .q(reg_dst_reg__m2s), .d(n3780), .sdi(
        reg_dst_of_MEM_4), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n917), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_4 reg_dst_reg__slave ( .q(reg_dst), .qb(n703), .d(reg_dst_reg__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n917), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 reg_out_A_reg_0__master ( .q(reg_out_A_reg_0__m2s), .d(N6718), 
        .sdi(n703), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n914), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_4 reg_out_A_reg_0__slave ( .q(reg_out_A[0]), .qb(n4051), .d(
        reg_out_A_reg_0__m2s), .g(Ctrl__Regs_1__en2), .rb(n914), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_A_reg_10__master ( .q(reg_out_A_reg_10__m2s), .d(N6728), 
        .sdi(n4042), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n915), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 reg_out_A_reg_10__slave ( .q(n3968), .qb(n4041), .d(
        reg_out_A_reg_10__m2s), .g(Ctrl__Regs_1__en2), .rb(n915), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_A_reg_11__master ( .q(reg_out_A_reg_11__m2s), .d(N6729), 
        .sdi(n4041), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n915), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_4 reg_out_A_reg_11__slave ( .q(n3967), .qb(n4040), .d(
        reg_out_A_reg_11__m2s), .g(Ctrl__Regs_1__en2), .rb(n915), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_A_reg_12__master ( .q(reg_out_A_reg_12__m2s), .d(N6730), 
        .sdi(n4040), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n915), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 reg_out_A_reg_12__slave ( .q(n3966), .qb(n4039), .d(
        reg_out_A_reg_12__m2s), .g(Ctrl__Regs_1__en2), .rb(n915), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_A_reg_13__master ( .q(reg_out_A_reg_13__m2s), .d(N6731), 
        .sdi(n4039), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n915), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_4 reg_out_A_reg_13__slave ( .q(reg_out_A[13]), .qb(n4038), .d(
        reg_out_A_reg_13__m2s), .g(Ctrl__Regs_1__en2), .rb(n915), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_A_reg_14__master ( .q(reg_out_A_reg_14__m2s), .d(N6732), 
        .sdi(n4038), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n915), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_4 reg_out_A_reg_14__slave ( .q(reg_out_A[14]), .qb(n4037), .d(
        reg_out_A_reg_14__m2s), .g(Ctrl__Regs_1__en2), .rb(n915), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_A_reg_15__master ( .q(reg_out_A_reg_15__m2s), .d(N6733), 
        .sdi(n4037), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n915), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_4 reg_out_A_reg_15__slave ( .q(reg_out_A[15]), .qb(n4036), .d(
        reg_out_A_reg_15__m2s), .g(Ctrl__Regs_1__en2), .rb(n915), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_A_reg_16__master ( .q(reg_out_A_reg_16__m2s), .d(N6734), 
        .sdi(n4036), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n915), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 reg_out_A_reg_16__slave ( .q(n3965), .qb(n4035), .d(
        reg_out_A_reg_16__m2s), .g(Ctrl__Regs_1__en2), .rb(n915), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_A_reg_17__master ( .q(reg_out_A_reg_17__m2s), .d(N6735), 
        .sdi(n4035), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n915), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_4 reg_out_A_reg_17__slave ( .q(n3964), .qb(n4034), .d(
        reg_out_A_reg_17__m2s), .g(Ctrl__Regs_1__en2), .rb(n915), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_A_reg_18__master ( .q(reg_out_A_reg_18__m2s), .d(N6736), 
        .sdi(n4034), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n916), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_4 reg_out_A_reg_18__slave ( .q(n3963), .qb(n4033), .d(
        reg_out_A_reg_18__m2s), .g(Ctrl__Regs_1__en2), .rb(n916), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_A_reg_19__master ( .q(reg_out_A_reg_19__m2s), .d(N6737), 
        .sdi(n4033), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n915), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 reg_out_A_reg_19__slave ( .q(n3962), .qb(n4032), .d(
        reg_out_A_reg_19__m2s), .g(Ctrl__Regs_1__en2), .rb(n915), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_A_reg_1__master ( .q(reg_out_A_reg_1__m2s), .d(N6719), 
        .sdi(n4051), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_4 reg_out_A_reg_1__slave ( .q(reg_out_A[1]), .qb(n4050), .d(
        reg_out_A_reg_1__m2s), .g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_A_reg_20__master ( .q(reg_out_A_reg_20__m2s), .d(N6738), 
        .sdi(n4032), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n916), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 reg_out_A_reg_20__slave ( .q(n3961), .qb(n4031), .d(
        reg_out_A_reg_20__m2s), .g(Ctrl__Regs_1__en2), .rb(n916), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_A_reg_21__master ( .q(reg_out_A_reg_21__m2s), .d(N6739), 
        .sdi(n4031), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n916), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 reg_out_A_reg_21__slave ( .q(n3960), .qb(n4030), .d(
        reg_out_A_reg_21__m2s), .g(Ctrl__Regs_1__en2), .rb(n916), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_A_reg_22__master ( .q(reg_out_A_reg_22__m2s), .d(N6740), 
        .sdi(n4030), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n916), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 reg_out_A_reg_22__slave ( .q(n3959), .qb(n4029), .d(
        reg_out_A_reg_22__m2s), .g(Ctrl__Regs_1__en2), .rb(n916), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_A_reg_23__master ( .q(reg_out_A_reg_23__m2s), .d(N6741), 
        .sdi(n4029), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n916), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 reg_out_A_reg_23__slave ( .q(n3958), .qb(n4028), .d(
        reg_out_A_reg_23__m2s), .g(Ctrl__Regs_1__en2), .rb(n916), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_A_reg_24__master ( .q(reg_out_A_reg_24__m2s), .d(N6742), 
        .sdi(n4028), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n913), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 reg_out_A_reg_24__slave ( .q(n3957), .qb(n4027), .d(
        reg_out_A_reg_24__m2s), .g(Ctrl__Regs_1__en2), .rb(n913), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_A_reg_25__master ( .q(reg_out_A_reg_25__m2s), .d(N6743), 
        .sdi(n4027), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n914), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 reg_out_A_reg_25__slave ( .q(n3956), .qb(n4026), .d(
        reg_out_A_reg_25__m2s), .g(Ctrl__Regs_1__en2), .rb(n914), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_A_reg_26__master ( .q(reg_out_A_reg_26__m2s), .d(N6744), 
        .sdi(n4026), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n914), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 reg_out_A_reg_26__slave ( .q(n3955), .qb(n4025), .d(
        reg_out_A_reg_26__m2s), .g(Ctrl__Regs_1__en2), .rb(n914), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_A_reg_27__master ( .q(reg_out_A_reg_27__m2s), .d(N6745), 
        .sdi(n4025), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n912), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 reg_out_A_reg_27__slave ( .q(n3954), .qb(n4024), .d(
        reg_out_A_reg_27__m2s), .g(Ctrl__Regs_1__en2), .rb(n912), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_A_reg_28__master ( .q(reg_out_A_reg_28__m2s), .d(N6746), 
        .sdi(n4024), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n916), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 reg_out_A_reg_28__slave ( .q(n3953), .qb(n4023), .d(
        reg_out_A_reg_28__m2s), .g(Ctrl__Regs_1__en2), .rb(n916), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_A_reg_29__master ( .q(reg_out_A_reg_29__m2s), .d(N6747), 
        .sdi(n4023), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n916), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 reg_out_A_reg_29__slave ( .q(n3952), .qb(n4022), .d(
        reg_out_A_reg_29__m2s), .g(Ctrl__Regs_1__en2), .rb(n916), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_A_reg_2__master ( .q(reg_out_A_reg_2__m2s), .d(N6720), 
        .sdi(n4050), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 reg_out_A_reg_2__slave ( .q(reg_out_A[2]), .qb(n4049), .d(
        reg_out_A_reg_2__m2s), .g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_A_reg_30__master ( .q(reg_out_A_reg_30__m2s), .d(N6748), 
        .sdi(n4022), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n916), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 reg_out_A_reg_30__slave ( .q(n3951), .qb(n4021), .d(
        reg_out_A_reg_30__m2s), .g(Ctrl__Regs_1__en2), .rb(n916), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_2 reg_out_A_reg_31__master ( .q(reg_out_A_reg_31__m2s), .d(N6749), 
        .sdi(n4021), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n912), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_8 reg_out_A_reg_31__slave ( .q(reg_out_A[31]), .qb(n4020), .d(
        reg_out_A_reg_31__m2s), .g(Ctrl__Regs_1__en2), .rb(n912), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_A_reg_3__master ( .q(reg_out_A_reg_3__m2s), .d(N6721), 
        .sdi(n4049), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n915), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_4 reg_out_A_reg_3__slave ( .q(n3974), .qb(n4048), .d(
        reg_out_A_reg_3__m2s), .g(Ctrl__Regs_1__en2), .rb(n915), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_A_reg_4__master ( .q(reg_out_A_reg_4__m2s), .d(N6722), 
        .sdi(n4048), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n915), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_4 reg_out_A_reg_4__slave ( .q(n3973), .qb(n4047), .d(
        reg_out_A_reg_4__m2s), .g(Ctrl__Regs_1__en2), .rb(n915), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_A_reg_5__master ( .q(reg_out_A_reg_5__m2s), .d(N6723), 
        .sdi(n4047), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n915), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_4 reg_out_A_reg_5__slave ( .q(n3972), .qb(n4046), .d(
        reg_out_A_reg_5__m2s), .g(Ctrl__Regs_1__en2), .rb(n915), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_A_reg_6__master ( .q(reg_out_A_reg_6__m2s), .d(N6724), 
        .sdi(n4046), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n916), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_4 reg_out_A_reg_6__slave ( .q(reg_out_A[6]), .qb(n4045), .d(
        reg_out_A_reg_6__m2s), .g(Ctrl__Regs_1__en2), .rb(n916), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_A_reg_7__master ( .q(reg_out_A_reg_7__m2s), .d(N6725), 
        .sdi(n4045), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n915), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_4 reg_out_A_reg_7__slave ( .q(n3971), .qb(n4044), .d(
        reg_out_A_reg_7__m2s), .g(Ctrl__Regs_1__en2), .rb(n915), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_A_reg_8__master ( .q(reg_out_A_reg_8__m2s), .d(N6726), 
        .sdi(n4044), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_4 reg_out_A_reg_8__slave ( .q(n3970), .qb(n4043), .d(
        reg_out_A_reg_8__m2s), .g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_A_reg_9__master ( .q(reg_out_A_reg_9__m2s), .d(N6727), 
        .sdi(n4043), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n915), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 reg_out_A_reg_9__slave ( .q(n3969), .qb(n4042), .d(
        reg_out_A_reg_9__m2s), .g(Ctrl__Regs_1__en2), .rb(n915), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_reg_0__master ( .q(reg_out_B_reg_0__m2s), .d(n4392), 
        .sdi(n4020), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n910), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_4 reg_out_B_reg_0__slave ( .q(n4458), .qb(n4393), .d(
        reg_out_B_reg_0__m2s), .g(Ctrl__Regs_1__en2), .rb(n910), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_2 reg_out_B_reg_10__master ( .q(reg_out_B_reg_10__m2s), .d(n4412), 
        .sdi(n4389), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n909), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_8 reg_out_B_reg_10__slave ( .q(reg_out_B[10]), .qb(n4413), .d(
        reg_out_B_reg_10__m2s), .g(Ctrl__Regs_1__en2), .rb(n909), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_2 reg_out_B_reg_11__master ( .q(reg_out_B_reg_11__m2s), .d(n4394), 
        .sdi(n4413), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n909), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_8 reg_out_B_reg_11__slave ( .q(reg_out_B[11]), .qb(n4395), .d(
        reg_out_B_reg_11__m2s), .g(Ctrl__Regs_1__en2), .rb(n909), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_reg_12__master ( .q(reg_out_B_reg_12__m2s), .d(n4432), 
        .sdi(n4395), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n909), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_4 reg_out_B_reg_12__slave ( .q(n3979), .qb(n4433), .d(
        reg_out_B_reg_12__m2s), .g(Ctrl__Regs_1__en2), .rb(n909), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_2 reg_out_B_reg_13__master ( .q(reg_out_B_reg_13__m2s), .d(n4424), 
        .sdi(n4433), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n909), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_8 reg_out_B_reg_13__slave ( .q(reg_out_B[13]), .qb(n4425), .d(
        reg_out_B_reg_13__m2s), .g(Ctrl__Regs_1__en2), .rb(n909), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_2 reg_out_B_reg_14__master ( .q(reg_out_B_reg_14__m2s), .d(n4420), 
        .sdi(n4425), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n910), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_8 reg_out_B_reg_14__slave ( .q(reg_out_B[14]), .qb(n4421), .d(
        reg_out_B_reg_14__m2s), .g(Ctrl__Regs_1__en2), .rb(n910), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_2 reg_out_B_reg_15__master ( .q(reg_out_B_reg_15__m2s), .d(n4402), 
        .sdi(n4421), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n909), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_8 reg_out_B_reg_15__slave ( .q(reg_out_B[15]), .qb(n4403), .d(
        reg_out_B_reg_15__m2s), .g(Ctrl__Regs_1__en2), .rb(n909), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_2 reg_out_B_reg_16__master ( .q(reg_out_B_reg_16__m2s), .d(n4410), 
        .sdi(n4403), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n910), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_8 reg_out_B_reg_16__slave ( .q(reg_out_B[16]), .qb(n4411), .d(
        reg_out_B_reg_16__m2s), .g(Ctrl__Regs_1__en2), .rb(n910), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_reg_17__master ( .q(reg_out_B_reg_17__m2s), .d(n4442), 
        .sdi(n4411), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n910), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_4 reg_out_B_reg_17__slave ( .q(n3978), .qb(n4443), .d(
        reg_out_B_reg_17__m2s), .g(Ctrl__Regs_1__en2), .rb(n910), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_2 reg_out_B_reg_18__master ( .q(reg_out_B_reg_18__m2s), .d(n4426), 
        .sdi(n4443), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n910), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_8 reg_out_B_reg_18__slave ( .q(reg_out_B[18]), .qb(n4427), .d(
        reg_out_B_reg_18__m2s), .g(Ctrl__Regs_1__en2), .rb(n910), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_reg_19__master ( .q(reg_out_B_reg_19__m2s), .d(n4422), 
        .sdi(n4427), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n910), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_4 reg_out_B_reg_19__slave ( .q(n4456), .qb(n4423), .d(
        reg_out_B_reg_19__m2s), .g(Ctrl__Regs_1__en2), .rb(n910), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_reg_1__master ( .q(reg_out_B_reg_1__m2s), .d(n4444), 
        .sdi(n4393), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n909), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_1 reg_out_B_reg_1__slave ( .q(n3983), .qb(n4445), .d(
        reg_out_B_reg_1__m2s), .g(Ctrl__Regs_1__en2), .rb(n909), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_2 reg_out_B_reg_20__master ( .q(reg_out_B_reg_20__m2s), .d(n4390), 
        .sdi(n4423), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n910), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_8 reg_out_B_reg_20__slave ( .q(reg_out_B[20]), .qb(n4391), .d(
        reg_out_B_reg_20__m2s), .g(Ctrl__Regs_1__en2), .rb(n910), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_reg_21__master ( .q(reg_out_B_reg_21__m2s), .d(n4436), 
        .sdi(n4391), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n909), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_4 reg_out_B_reg_21__slave ( .q(reg_out_B[21]), .qb(n4437), .d(
        reg_out_B_reg_21__m2s), .g(Ctrl__Regs_1__en2), .rb(n909), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_reg_22__master ( .q(reg_out_B_reg_22__m2s), .d(n4446), 
        .sdi(n4437), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n910), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_4 reg_out_B_reg_22__slave ( .q(n3977), .qb(n4447), .d(
        reg_out_B_reg_22__m2s), .g(Ctrl__Regs_1__en2), .rb(n910), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_2 reg_out_B_reg_23__master ( .q(reg_out_B_reg_23__m2s), .d(n4414), 
        .sdi(n4447), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n910), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_8 reg_out_B_reg_23__slave ( .q(reg_out_B[23]), .qb(n4415), .d(
        reg_out_B_reg_23__m2s), .g(Ctrl__Regs_1__en2), .rb(n910), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_2 reg_out_B_reg_24__master ( .q(reg_out_B_reg_24__m2s), .d(n4416), 
        .sdi(n4415), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n910), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_8 reg_out_B_reg_24__slave ( .q(reg_out_B[24]), .qb(n4417), .d(
        reg_out_B_reg_24__m2s), .g(Ctrl__Regs_1__en2), .rb(n910), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_reg_25__master ( .q(reg_out_B_reg_25__m2s), .d(n4434), 
        .sdi(n4417), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n911), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_4 reg_out_B_reg_25__slave ( .q(n4455), .qb(n4435), .d(
        reg_out_B_reg_25__m2s), .g(Ctrl__Regs_1__en2), .rb(n911), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_2 reg_out_B_reg_26__master ( .q(reg_out_B_reg_26__m2s), .d(n4406), 
        .sdi(n4435), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n910), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_8 reg_out_B_reg_26__slave ( .q(reg_out_B[26]), .qb(n4407), .d(
        reg_out_B_reg_26__m2s), .g(Ctrl__Regs_1__en2), .rb(n910), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_2 reg_out_B_reg_27__master ( .q(reg_out_B_reg_27__m2s), .d(n4430), 
        .sdi(n4407), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n910), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_8 reg_out_B_reg_27__slave ( .q(reg_out_B[27]), .qb(n4431), .d(
        reg_out_B_reg_27__m2s), .g(Ctrl__Regs_1__en2), .rb(n910), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_2 reg_out_B_reg_28__master ( .q(reg_out_B_reg_28__m2s), .d(n4400), 
        .sdi(n4431), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n909), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_8 reg_out_B_reg_28__slave ( .q(reg_out_B[28]), .qb(n4401), .d(
        reg_out_B_reg_28__m2s), .g(Ctrl__Regs_1__en2), .rb(n909), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_2 reg_out_B_reg_29__master ( .q(reg_out_B_reg_29__m2s), .d(n4396), 
        .sdi(n4401), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n910), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_8 reg_out_B_reg_29__slave ( .q(reg_out_B[29]), .qb(n4397), .d(
        reg_out_B_reg_29__m2s), .g(Ctrl__Regs_1__en2), .rb(n910), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_reg_2__master ( .q(reg_out_B_reg_2__m2s), .d(n4438), 
        .sdi(n4445), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n912), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_4 reg_out_B_reg_2__slave ( .q(n3982), .qb(n4439), .d(
        reg_out_B_reg_2__m2s), .g(Ctrl__Regs_1__en2), .rb(n912), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_2 reg_out_B_reg_30__master ( .q(reg_out_B_reg_30__m2s), .d(n4448), 
        .sdi(n4397), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n911), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_8 reg_out_B_reg_30__slave ( .q(reg_out_B[30]), .qb(n4449), .d(
        reg_out_B_reg_30__m2s), .g(Ctrl__Regs_1__en2), .rb(n911), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_reg_31__master ( .q(reg_out_B_reg_31__m2s), .d(n4450), 
        .sdi(n4449), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n911), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_4 reg_out_B_reg_31__slave ( .q(reg_out_B[31]), .qb(n4451), .d(
        reg_out_B_reg_31__m2s), .g(Ctrl__Regs_1__en2), .rb(n911), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_reg_3__master ( .q(reg_out_B_reg_3__m2s), .d(n4440), 
        .sdi(n4439), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n912), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_1 reg_out_B_reg_3__slave ( .q(n3981), .qb(n4441), .d(
        reg_out_B_reg_3__m2s), .g(Ctrl__Regs_1__en2), .rb(n912), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_reg_4__master ( .q(reg_out_B_reg_4__m2s), .d(n4398), 
        .sdi(n4441), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n912), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_1 reg_out_B_reg_4__slave ( .q(n3980), .qb(n4399), .d(
        reg_out_B_reg_4__m2s), .g(Ctrl__Regs_1__en2), .rb(n912), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_2 reg_out_B_reg_5__master ( .q(reg_out_B_reg_5__m2s), .d(n4418), 
        .sdi(n4399), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n909), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_8 reg_out_B_reg_5__slave ( .q(reg_out_B[5]), .qb(n4419), .d(
        reg_out_B_reg_5__m2s), .g(Ctrl__Regs_1__en2), .rb(n909), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_reg_6__master ( .q(reg_out_B_reg_6__m2s), .d(n4404), 
        .sdi(n4419), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n909), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 reg_out_B_reg_6__slave ( .q(n4457), .qb(n4405), .d(
        reg_out_B_reg_6__m2s), .g(Ctrl__Regs_1__en2), .rb(n909), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_reg_7__master ( .q(reg_out_B_reg_7__m2s), .d(n4428), 
        .sdi(n4405), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n909), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_4 reg_out_B_reg_7__slave ( .q(reg_out_B[7]), .qb(n4429), .d(
        reg_out_B_reg_7__m2s), .g(Ctrl__Regs_1__en2), .rb(n909), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_2 reg_out_B_reg_8__master ( .q(reg_out_B_reg_8__m2s), .d(n4408), 
        .sdi(n4429), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n909), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_8 reg_out_B_reg_8__slave ( .q(reg_out_B[8]), .qb(n4409), .d(
        reg_out_B_reg_8__m2s), .g(Ctrl__Regs_1__en2), .rb(n909), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_2 reg_out_B_reg_9__master ( .q(reg_out_B_reg_9__m2s), .d(n4388), 
        .sdi(n4409), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n909), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_8 reg_out_B_reg_9__slave ( .q(reg_out_B[9]), .qb(n4389), .d(
        reg_out_B_reg_9__m2s), .g(Ctrl__Regs_1__en2), .rb(n909), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_write_reg__master ( .q(reg_write_reg__m2s), .d(n3779), .sdi(
        n4451), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 reg_write_reg__slave ( .q(reg_write), .qb(n2638), .d(
        reg_write_reg__m2s), .g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 rt_addr_reg_0__master ( .q(rt_addr_reg_0__m2s), .d(n3786), .sdi(
        reg_write), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n917), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 rt_addr_reg_0__slave ( .q(rt_addr[0]), .qb(n561), .d(
        rt_addr_reg_0__m2s), .g(Ctrl__Regs_1__en2), .rb(n917), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 rt_addr_reg_1__master ( .q(rt_addr_reg_1__m2s), .d(n3787), .sdi(
        rt_addr[0]), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 rt_addr_reg_1__slave ( .q(rt_addr[1]), .qb(n560), .d(
        rt_addr_reg_1__m2s), .g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 rt_addr_reg_2__master ( .q(rt_addr_reg_2__m2s), .d(n3788), .sdi(
        rt_addr[1]), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n917), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 rt_addr_reg_2__slave ( .q(rt_addr[2]), .qb(n559), .d(
        rt_addr_reg_2__m2s), .g(Ctrl__Regs_1__en2), .rb(n917), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 rt_addr_reg_3__master ( .q(rt_addr_reg_3__m2s), .d(n3789), .sdi(
        rt_addr[2]), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 rt_addr_reg_3__slave ( .q(rt_addr[3]), .qb(n671), .d(
        rt_addr_reg_3__m2s), .g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 rt_addr_reg_4__master ( .q(rt_addr_reg_4__m2s), .d(n3790), .sdi(
        n671), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n916), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 rt_addr_reg_4__slave ( .q(rt_addr[4]), .qb(n558), .d(
        rt_addr_reg_4__m2s), .g(Ctrl__Regs_1__en2), .rb(n916), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 slot_num_reg_0__master ( .q(slot_num_reg_0__m2s), .d(n2705), 
        .sdi(rt_addr[4]), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_4 slot_num_reg_0__slave ( .q(slot_num_0), .qb(n4019), .d(
        slot_num_reg_0__m2s), .g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 slot_num_reg_1__master ( .q(slot_num_reg_1__m2s), .d(n2706), 
        .sdi(n4019), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n916), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_4 slot_num_reg_1__slave ( .q(slot_num_1), .qb(n557), .d(
        slot_num_reg_1__m2s), .g(Ctrl__Regs_1__en2), .rb(n916), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 stall_reg__master ( .q(stall_reg__m2s), .d(n2708), .sdi(n557), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 stall_reg__slave ( .q(stall), .qb(n2639), .d(stall_reg__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n982), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    ID_DW01_add_32_0_test_1 sub_489 ( .A({n331, n331, n331, n331, n331, n331, 
        n331, n824, n695, n3990, n3998, n802, n337, n878, n892, n340, n887, 
        IR_latched_14, IR_latched_13, IR_latched_12, IR_latched_11, 
        IR_latched_10, n809, IR_latched_8, n817, n3999, n888, n832, 
        IR_latched_3, IR_latched_2, IR_latched_1, IR_latched_0}), .B({N5350, 
        N5349, N5348, N5347, N5346, N5345, N5344, N5343, N5342, N5341, N5340, 
        N5339, N5338, N5337, N5336, N5335, N5334, N5333, N5332, N5331, N5330, 
        N5329, N5328, N5327, N5326, N5325, N5324, N5323, N5322, N5321, N5320, 
        N5319}), .CI(1'b0), .SUM({N5382, N5381, N5380, N5379, N5378, N5377, 
        N5376, N5375, N5374, N5373, N5372, N5371, N5370, N5369, N5368, N5367, 
        N5366, N5365, N5364, N5363, N5362, N5361, N5360, N5359, N5358, N5357, 
        N5356, N5355, N5354, N5353, N5352, N5351}) );
    ID_DW01_add_32_2_test_1 sub_609 ( .A({n331, n331, n331, n331, n331, n331, 
        n331, n719, n695, n3990, n335, n336, n337, n878, n833, n340, 
        IR_latched_15, IR_latched_14, IR_latched_13, IR_latched_12, 
        IR_latched_11, IR_latched_10, IR_latched_9, IR_latched_8, n817, n3999, 
        n888, IR_latched_4, IR_latched_3, IR_latched_2, IR_latched_1, 
        IR_latched_0}), .B({N5418, N5417, N5416, N5415, N5414, N5413, N5412, 
        N5411, N5410, N5409, N5408, N5407, N5406, N5405, N5404, N5403, N5402, 
        N5401, N5400, N5399, N5398, N5397, N5396, N5395, N5394, N5393, N5392, 
        N5391, N5390, N5389, N5388, N5387}), .CI(1'b0), .SUM({N5450, N5449, 
        N5448, N5447, N5446, N5445, N5444, N5443, N5442, N5441, N5440, N5439, 
        N5438, N5437, N5436, N5435, N5434, N5433, N5432, N5431, N5430, N5429, 
        N5428, N5427, N5426, N5425, N5424, N5423, N5422, N5421, N5420, N5419})
         );
    ID_DW01_add_32_1_test_1 sub_779 ( .A({n887, n887, n887, n887, n887, n887, 
        n887, n887, n887, n887, n887, n887, n887, n887, n887, n887, n887, 
        IR_latched_14, IR_latched_13, IR_latched_12, IR_latched_11, 
        IR_latched_10, n809, IR_latched_8, n817, n3999, n888, n831, 
        IR_latched_3, IR_latched_2, IR_latched_1, IR_latched_0}), .B({N6017, 
        N6016, N6015, N6014, N6013, N6012, N6011, N6010, N6009, N6008, N6007, 
        N6006, N6005, N6004, N6003, N6002, N6001, N6000, N5999, N5998, N5997, 
        N5996, N5995, N5994, N5993, N5992, N5991, N5990, N5989, N5988, N5987, 
        N5986}), .CI(1'b0), .SUM({N6049, N6048, N6047, N6046, N6045, N6044, 
        N6043, N6042, N6041, N6040, N6039, N6038, N6037, N6036, N6035, N6034, 
        N6033, N6032, N6031, N6030, N6029, N6028, N6027, N6026, N6025, N6024, 
        N6023, N6022, N6021, N6020, N6019, N6018}) );
endmodule


module IF_DW01_add_32_0_test_1 ( A, B, CI, SUM, CO );
input  [31:0] A;
input  [31:0] B;
output [31:0] SUM;
input  CI;
output CO;
    wire A_1, A_0, n72, n106, n107, n80, n114, n115, n82, n121, n79, n116, 
        n122, n81, n94, n111, n83, n131, n62, n71, n130, n67, n129, n102, n64, 
        n69, n112, n74, n77, n132, n59, n99, n104, n109, n128, n68, n70, n105, 
        n92, n58, n125, n57, n123, n96, n124, n49, n101, n66, n63, n65, n97, 
        n61, n126, n60, n117, n118, n53, n87, n88, n52, n54, n56, n91, n73, 
        n75, n76, n78, n108, n95, n50, n86, n84, n120, n51, n103, n100, n98, 
        n127, n119, n90, n89, n55, n93, n110, n113, n85;
    assign A_1 = A[1];
    assign A_0 = A[0];
    assign SUM[1] = A_1;
    assign SUM[0] = A_0;
    nand2i_2 U10 ( .x(n72), .a(n106), .b(n107) );
    nand2i_4 U100 ( .x(n80), .a(n114), .b(n115) );
    exnor2_5 U101 ( .x(SUM[31]), .a(n82), .b(n121) );
    exnor2_5 U102 ( .x(SUM[30]), .a(n79), .b(n116) );
    exnor2_3 U103 ( .x(SUM[29]), .a(n122), .b(n81) );
    nand4_1 U104 ( .x(n94), .a(A[7]), .b(A[8]), .c(A[10]), .d(A[9]) );
    nand2_2 U106 ( .x(n111), .a(A[26]), .b(A[25]) );
    nand2_2 U107 ( .x(n114), .a(A[27]), .b(A[28]) );
    nand2_2 U108 ( .x(n83), .a(A[30]), .b(A[29]) );
    inv_5 U109 ( .x(n131), .a(n62) );
    nor2i_1 U11 ( .x(n71), .a(A[23]), .b(n72) );
    inv_5 U110 ( .x(n130), .a(n67) );
    inv_5 U111 ( .x(n129), .a(n72) );
    inv_5 U112 ( .x(n102), .a(n64) );
    inv_5 U113 ( .x(n107), .a(n69) );
    inv_5 U114 ( .x(n112), .a(n74) );
    inv_5 U115 ( .x(n115), .a(n77) );
    inv_6 U116 ( .x(n132), .a(n59) );
    nand2i_6 U117 ( .x(n64), .a(n99), .b(n131) );
    nand2i_6 U118 ( .x(n69), .a(n104), .b(n130) );
    nand2i_0 U119 ( .x(n109), .a(n128), .b(A[24]) );
    nor2_1 U12 ( .x(n68), .a(n69), .b(n70) );
    nand2_0 U120 ( .x(n106), .a(A[21]), .b(A[22]) );
    inv_0 U121 ( .x(n105), .a(A[22]) );
    nand2i_2 U13 ( .x(n59), .a(n94), .b(n92) );
    inv_2 U14 ( .x(n58), .a(n125) );
    nor2i_1 U15 ( .x(n57), .a(n58), .b(n59) );
    nand2i_2 U16 ( .x(n123), .a(n96), .b(n124) );
    nor2i_1 U17 ( .x(n49), .a(A[3]), .b(SUM[2]) );
    nand2i_2 U18 ( .x(n67), .a(n101), .b(n102) );
    nor2i_1 U19 ( .x(n66), .a(A[19]), .b(n67) );
    nor2_1 U20 ( .x(n63), .a(n64), .b(n65) );
    nand2i_2 U21 ( .x(n62), .a(n97), .b(n132) );
    inv_2 U22 ( .x(n61), .a(n126) );
    nor2i_1 U23 ( .x(n60), .a(n61), .b(n62) );
    inv_0 U24 ( .x(n125), .a(A[11]) );
    nand2i_2 U25 ( .x(n117), .a(n118), .b(n132) );
    inv_2 U26 ( .x(n92), .a(n53) );
    nand3i_1 U27 ( .x(n53), .a(SUM[2]), .b(n87), .c(n88) );
    nor2_1 U28 ( .x(n52), .a(n53), .b(n54) );
    nand2i_2 U29 ( .x(n56), .a(n91), .b(n92) );
    nand2i_2 U30 ( .x(n74), .a(n109), .b(n129) );
    nor2_1 U31 ( .x(n73), .a(n74), .b(n75) );
    nand2i_2 U32 ( .x(n77), .a(n111), .b(n112) );
    nor2_1 U33 ( .x(n76), .a(n77), .b(n78) );
    exnor2_1 U34 ( .x(SUM[24]), .a(n71), .b(n108) );
    exnor2_1 U35 ( .x(SUM[22]), .a(n68), .b(n105) );
    exnor2_1 U36 ( .x(SUM[12]), .a(n57), .b(n95) );
    exnor2_2 U37 ( .x(SUM[21]), .a(n107), .b(n70) );
    exnor2_2 U38 ( .x(SUM[25]), .a(n112), .b(n75) );
    exnor2_1 U39 ( .x(SUM[6]), .a(n50), .b(n86) );
    exnor2_1 U40 ( .x(SUM[4]), .a(n49), .b(n84) );
    inv_2 U41 ( .x(n120), .a(n51) );
    exnor2_1 U42 ( .x(SUM[11]), .a(n132), .b(n125) );
    exnor2_1 U43 ( .x(SUM[20]), .a(n66), .b(n103) );
    exnor2_3 U44 ( .x(SUM[23]), .a(n129), .b(n128) );
    exnor2_1 U45 ( .x(SUM[18]), .a(n63), .b(n100) );
    exnor2_1 U46 ( .x(SUM[17]), .a(n102), .b(n65) );
    exnor2_1 U47 ( .x(SUM[15]), .a(n131), .b(n126) );
    exnor2_1 U48 ( .x(SUM[16]), .a(n60), .b(n98) );
    exnor2_1 U49 ( .x(SUM[13]), .a(n124), .b(n96) );
    nand2i_2 U5 ( .x(n104), .a(n127), .b(A[20]) );
    inv_2 U50 ( .x(n124), .a(n117) );
    exnor2_2 U51 ( .x(SUM[19]), .a(n130), .b(n127) );
    exnor2_2 U52 ( .x(SUM[7]), .a(n92), .b(n54) );
    inv_2 U53 ( .x(n54), .a(A[7]) );
    exnor2_1 U54 ( .x(SUM[9]), .a(n119), .b(n90) );
    inv_2 U55 ( .x(n119), .a(n56) );
    exnor2_1 U56 ( .x(SUM[8]), .a(n52), .b(n89) );
    exnor2_1 U57 ( .x(SUM[10]), .a(n55), .b(n93) );
    exor2_1 U58 ( .x(SUM[3]), .a(A[3]), .b(A[2]) );
    inv_2 U59 ( .x(SUM[2]), .a(A[2]) );
    nand2i_0 U6 ( .x(n99), .a(n126), .b(A[16]) );
    inv_1 U60 ( .x(n103), .a(A[20]) );
    inv_0 U61 ( .x(n75), .a(A[25]) );
    inv_2 U62 ( .x(n81), .a(A[29]) );
    exnor2_1 U63 ( .x(SUM[26]), .a(n73), .b(n110) );
    exnor2_1 U64 ( .x(SUM[27]), .a(n115), .b(n78) );
    exnor2_1 U65 ( .x(SUM[28]), .a(n76), .b(n113) );
    inv_2 U66 ( .x(n122), .a(n80) );
    inv_0 U67 ( .x(n108), .a(A[24]) );
    inv_0 U69 ( .x(n70), .a(A[21]) );
    nor2i_1 U7 ( .x(n88), .a(A[3]), .b(n84) );
    inv_0 U70 ( .x(n127), .a(A[19]) );
    inv_2 U71 ( .x(n78), .a(A[27]) );
    inv_2 U72 ( .x(n113), .a(A[28]) );
    inv_2 U73 ( .x(n116), .a(A[30]) );
    inv_2 U74 ( .x(n121), .a(A[31]) );
    inv_2 U75 ( .x(n128), .a(A[23]) );
    exnor2_1 U76 ( .x(SUM[5]), .a(n120), .b(n85) );
    inv_0 U77 ( .x(n98), .a(A[16]) );
    inv_0 U78 ( .x(n126), .a(A[15]) );
    inv_0 U79 ( .x(n65), .a(A[17]) );
    inv_0 U80 ( .x(n89), .a(A[8]) );
    nor2i_0 U81 ( .x(n87), .a(A[6]), .b(n85) );
    inv_0 U82 ( .x(n86), .a(A[6]) );
    inv_0 U83 ( .x(n96), .a(A[13]) );
    nand2_0 U84 ( .x(n101), .a(A[17]), .b(A[18]) );
    inv_0 U85 ( .x(n100), .a(A[18]) );
    nand3i_0 U86 ( .x(n51), .a(SUM[2]), .b(A[4]), .c(A[3]) );
    inv_1 U87 ( .x(n84), .a(A[4]) );
    exnor2_1 U88 ( .x(SUM[14]), .a(A[14]), .b(n123) );
    inv_0 U89 ( .x(n93), .a(A[10]) );
    inv_0 U9 ( .x(n110), .a(A[26]) );
    inv_0 U90 ( .x(n90), .a(A[9]) );
    nor2i_0 U91 ( .x(n55), .a(A[9]), .b(n56) );
    nand2_0 U92 ( .x(n91), .a(A[7]), .b(A[8]) );
    inv_0 U93 ( .x(n95), .a(A[12]) );
    nand2i_0 U94 ( .x(n118), .a(n125), .b(A[12]) );
    nand4i_1 U95 ( .x(n97), .a(n125), .b(A[13]), .c(A[12]), .d(A[14]) );
    nor2i_0 U96 ( .x(n50), .a(A[5]), .b(n51) );
    inv_0 U97 ( .x(n85), .a(A[5]) );
    nor2_5 U98 ( .x(n79), .a(n80), .b(n81) );
    nor2_5 U99 ( .x(n82), .a(n80), .b(n83) );
endmodule


module IF_test_1_desync ( NPC, PC, IR_latched, reset, branch_sig, 
    branch_address, IR, stall, counter, test_si1, test_so1, test_si2, test_se, 
    sync_sel, global_g1, global_g2, Ctrl__Regs_1__en1, Ctrl__Regs_1__en2 );
output [31:0] NPC;
output [31:0] PC;
output [31:0] IR_latched;
input  [31:0] branch_address;
input  [31:0] IR;
input  [1:0] counter;
input  reset, branch_sig, stall, test_si1, test_si2, test_se, sync_sel, 
    global_g1, global_g2, Ctrl__Regs_1__en1, Ctrl__Regs_1__en2;
output test_so1;
    wire IR_curr_reg_0__m2s, n136, n41, IR_curr_0, n358, IR_curr_reg_10__m2s, 
        n146, n349, IR_curr_10, n348, IR_curr_reg_11__m2s, n147, IR_curr_11, 
        n347, IR_curr_reg_12__m2s, n148, IR_curr_12, n346, IR_curr_reg_13__m2s, 
        n149, IR_curr_13, n345, IR_curr_reg_14__m2s, n150, n42, IR_curr_14, 
        n344, IR_curr_reg_15__m2s, n151, IR_curr_15, n343, IR_curr_reg_16__m2s, 
        n152, IR_curr_16, n342, IR_curr_reg_17__m2s, n153, IR_curr_17, n341, 
        IR_curr_reg_18__m2s, n154, IR_curr_18, n340, IR_curr_reg_19__m2s, n155, 
        IR_curr_19, n339, IR_curr_reg_1__m2s, n137, IR_curr_1, n357, 
        IR_curr_reg_20__m2s, n156, IR_curr_20, n338, IR_curr_reg_21__m2s, n157, 
        IR_curr_21, n337, IR_curr_reg_22__m2s, n158, IR_curr_22, n336, 
        IR_curr_reg_23__m2s, n159, IR_curr_23, n335, IR_curr_reg_24__m2s, n160, 
        IR_curr_24, n334, IR_curr_reg_25__m2s, n161, IR_curr_25, n333, 
        IR_curr_reg_26__m2s, n162, IR_curr_26, n332, IR_curr_reg_27__m2s, n163, 
        IR_curr_27, n331, IR_curr_reg_28__m2s, n164, IR_curr_28, n330, 
        IR_curr_reg_29__m2s, n165, IR_curr_29, n329, IR_curr_reg_2__m2s, n138, 
        IR_curr_2, n356, IR_curr_reg_30__m2s, n166, IR_curr_30, n328, 
        IR_curr_reg_31__m2s, n167, IR_curr_31, n327, IR_curr_reg_3__m2s, n139, 
        IR_curr_3, n355, IR_curr_reg_4__m2s, n140, IR_curr_4, n354, 
        IR_curr_reg_5__m2s, n141, IR_curr_5, n353, IR_curr_reg_6__m2s, n142, 
        IR_curr_6, n352, IR_curr_reg_7__m2s, n143, n40, IR_curr_7, n351, 
        IR_curr_reg_8__m2s, n144, IR_curr_8, n350, IR_curr_reg_9__m2s, n145, 
        IR_curr_9, IR_latched_reg_0__m2s, N119, n38, n326, 
        IR_latched_reg_10__m2s, N129, n317, n316, IR_latched_reg_11__m2s, N130, 
        n315, IR_latched_reg_12__m2s, N131, n314, IR_latched_reg_13__m2s, N132, 
        n313, IR_latched_reg_14__m2s, N133, n312, IR_latched_reg_15__m2s, N134, 
        n311, IR_latched_reg_16__m2s, N135, n37, n310, IR_latched_reg_17__m2s, 
        N136, n309, IR_latched_reg_18__m2s, N137, n308, IR_latched_reg_19__m2s, 
        N138, n307, IR_latched_reg_1__m2s, N120, n325, IR_latched_reg_20__m2s, 
        N139, n306, IR_latched_reg_21__m2s, N140, n305, IR_latched_reg_22__m2s, 
        N141, n304, IR_latched_reg_23__m2s, N142, n303, IR_latched_reg_24__m2s, 
        N143, n302, IR_latched_reg_25__m2s, N144, n301, IR_latched_reg_26__m2s, 
        N145, n300, IR_latched_reg_27__m2s, N146, n299, IR_latched_reg_28__m2s, 
        N147, n298, IR_latched_reg_29__m2s, N148, n297, IR_latched_reg_2__m2s, 
        N121, n324, IR_latched_reg_30__m2s, N149, n296, IR_latched_reg_31__m2s, 
        N150, n295, IR_latched_reg_3__m2s, N122, n323, IR_latched_reg_4__m2s, 
        N123, n322, IR_latched_reg_5__m2s, N124, n321, IR_latched_reg_6__m2s, 
        N125, n320, IR_latched_reg_7__m2s, N126, n319, IR_latched_reg_8__m2s, 
        N127, n318, IR_latched_reg_9__m2s, N128, IR_previous_reg_0__m2s, n104, 
        IR_previous_0, n294, IR_previous_reg_10__m2s, n114, n285, 
        IR_previous_10, n284, IR_previous_reg_11__m2s, n115, IR_previous_11, 
        n283, IR_previous_reg_12__m2s, n116, IR_previous_12, n282, 
        IR_previous_reg_13__m2s, n117, IR_previous_13, n281, 
        IR_previous_reg_14__m2s, n118, IR_previous_14, n280, 
        IR_previous_reg_15__m2s, n119, IR_previous_15, n279, 
        IR_previous_reg_16__m2s, n120, n43, IR_previous_16, n278, 
        IR_previous_reg_17__m2s, n121, IR_previous_17, n277, 
        IR_previous_reg_18__m2s, n122, IR_previous_18, n276, 
        IR_previous_reg_19__m2s, n123, IR_previous_19, n275, 
        IR_previous_reg_1__m2s, n105, IR_previous_1, n293, 
        IR_previous_reg_20__m2s, n124, IR_previous_20, n274, 
        IR_previous_reg_21__m2s, n125, IR_previous_21, n273, 
        IR_previous_reg_22__m2s, n126, IR_previous_22, n272, 
        IR_previous_reg_23__m2s, n127, IR_previous_23, n271, 
        IR_previous_reg_24__m2s, n128, IR_previous_24, n270, 
        IR_previous_reg_25__m2s, n129, IR_previous_25, n269, 
        IR_previous_reg_26__m2s, n130, IR_previous_26, n268, 
        IR_previous_reg_27__m2s, n131, IR_previous_27, n267, 
        IR_previous_reg_28__m2s, n132, IR_previous_28, n266, 
        IR_previous_reg_29__m2s, n133, IR_previous_29, n265, 
        IR_previous_reg_2__m2s, n106, IR_previous_2, n292, 
        IR_previous_reg_30__m2s, n134, IR_previous_30, n264, 
        IR_previous_reg_31__m2s, n135, IR_previous_31, n263, 
        IR_previous_reg_3__m2s, n107, IR_previous_3, n291, 
        IR_previous_reg_4__m2s, n108, IR_previous_4, n290, 
        IR_previous_reg_5__m2s, n109, IR_previous_5, n289, 
        IR_previous_reg_6__m2s, n110, IR_previous_6, n288, 
        IR_previous_reg_7__m2s, n111, IR_previous_7, n287, 
        IR_previous_reg_8__m2s, n112, IR_previous_8, n286, 
        IR_previous_reg_9__m2s, n113, n39, IR_previous_9, NPC_reg_0__m2s, N87, 
        n36, n262, NPC_reg_10__m2s, N97, n22, n24, NPC_reg_11__m2s, N98, n205, 
        n257, NPC_reg_12__m2s, N99, n28, NPC_reg_13__m2s, N100, n14, 
        NPC_reg_14__m2s, N101, n360, n12, NPC_reg_15__m2s, N102, n204, n256, 
        NPC_reg_16__m2s, N103, n255, NPC_reg_17__m2s, N104, n10, 
        NPC_reg_18__m2s, N105, n254, NPC_reg_19__m2s, N106, n253, 
        NPC_reg_1__m2s, N88, n261, NPC_reg_20__m2s, N107, n252, 
        NPC_reg_21__m2s, N108, n251, NPC_reg_22__m2s, N109, n250, 
        NPC_reg_23__m2s, N110, n249, NPC_reg_24__m2s, N111, n91, n248, 
        NPC_reg_25__m2s, N112, n247, NPC_reg_26__m2s, N113, n246, 
        NPC_reg_27__m2s, N114, n245, NPC_reg_28__m2s, N115, n244, 
        NPC_reg_29__m2s, N116, n243, NPC_reg_2__m2s, N89, n210, n32, 
        NPC_reg_30__m2s, N117, n242, NPC_reg_31__m2s, N118, NPC_reg_3__m2s, 
        N90, n209, n30, NPC_reg_4__m2s, N91, n208, n260, NPC_reg_5__m2s, N92, 
        n207, n259, NPC_reg_6__m2s, N93, n206, n258, NPC_reg_7__m2s, N94, n26, 
        NPC_reg_8__m2s, N95, n16, NPC_reg_9__m2s, N96, PC_reg_0__m2s, n168, 
        n241, PC_reg_10__m2s, n178, n232, n231, PC_reg_11__m2s, n179, n230, 
        PC_reg_12__m2s, n180, n229, PC_reg_13__m2s, n181, n228, PC_reg_14__m2s, 
        n182, n227, PC_reg_15__m2s, n183, n226, PC_reg_16__m2s, n184, n225, 
        PC_reg_17__m2s, n185, n224, PC_reg_18__m2s, n186, n223, PC_reg_19__m2s, 
        n187, n222, PC_reg_1__m2s, n169, n240, PC_reg_20__m2s, n188, n221, 
        PC_reg_21__m2s, n189, n92, PC_reg_22__m2s, n190, n93, PC_reg_23__m2s, 
        n191, n94, PC_reg_24__m2s, n192, n95, PC_reg_25__m2s, n193, n96, 
        PC_reg_26__m2s, n194, n97, PC_reg_27__m2s, n195, n98, PC_reg_28__m2s, 
        n196, n99, PC_reg_29__m2s, n197, n100, PC_reg_2__m2s, n170, n239, 
        PC_reg_30__m2s, n198, n101, PC_reg_31__m2s, n199, n102, PC_reg_3__m2s, 
        n171, n238, PC_reg_4__m2s, n172, n237, PC_reg_5__m2s, n173, n236, 
        PC_reg_6__m2s, n174, n235, PC_reg_7__m2s, n175, n234, PC_reg_8__m2s, 
        n176, n233, PC_reg_9__m2s, n177, n48, n87, n81, n83, n89, n218, n49, 
        N152, n33, n90, n31, n214, n4, n202, n200, n88, n5, n6, N18, N215, 
        n201, n44, n45, n46, N50, n203, n61, n59, N43, N38, n60, n64, n63, n62, 
        N44, n67, n66, n65, N45, n86, n69, n70, n68, n85, n78, n79, n77, n76, 
        N48, n84, n74, n75, n73, n82, n72, N34, N28, n8, n7, n56, n57, n58, 
        N22, N31, n11, n13, n15, N17, N21, N42, N27, N23, n17, n23, n211, n25, 
        n27, N20, n29, n212, n71, N46, n80, N47, N29, N37, n213, n215, N33, 
        n217, N30, n50, n51, n52, N36, N40, n53, n54, n55, N35, N32, N24, N26, 
        N25, N19, N41, n47, N39, stalled_reg__m2s;
    smlatnr_1 IR_curr_reg_0__master ( .q(IR_curr_reg_0__m2s), .d(n136), .sdi(
        test_si1), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n41), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_curr_reg_0__slave ( .q(IR_curr_0), .qb(n358), .d(
        IR_curr_reg_0__m2s), .g(Ctrl__Regs_1__en2), .rb(n41), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_curr_reg_10__master ( .q(IR_curr_reg_10__m2s), .d(n146), 
        .sdi(n349), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n41), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_curr_reg_10__slave ( .q(IR_curr_10), .qb(n348), .d(
        IR_curr_reg_10__m2s), .g(Ctrl__Regs_1__en2), .rb(n41), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_curr_reg_11__master ( .q(IR_curr_reg_11__m2s), .d(n147), 
        .sdi(n348), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n41), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_curr_reg_11__slave ( .q(IR_curr_11), .qb(n347), .d(
        IR_curr_reg_11__m2s), .g(Ctrl__Regs_1__en2), .rb(n41), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_curr_reg_12__master ( .q(IR_curr_reg_12__m2s), .d(n148), 
        .sdi(n347), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n41), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_curr_reg_12__slave ( .q(IR_curr_12), .qb(n346), .d(
        IR_curr_reg_12__m2s), .g(Ctrl__Regs_1__en2), .rb(n41), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_curr_reg_13__master ( .q(IR_curr_reg_13__m2s), .d(n149), 
        .sdi(n346), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n41), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_curr_reg_13__slave ( .q(IR_curr_13), .qb(n345), .d(
        IR_curr_reg_13__m2s), .g(Ctrl__Regs_1__en2), .rb(n41), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_curr_reg_14__master ( .q(IR_curr_reg_14__m2s), .d(n150), 
        .sdi(n345), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n42), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_curr_reg_14__slave ( .q(IR_curr_14), .qb(n344), .d(
        IR_curr_reg_14__m2s), .g(Ctrl__Regs_1__en2), .rb(n42), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_curr_reg_15__master ( .q(IR_curr_reg_15__m2s), .d(n151), 
        .sdi(n344), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n41), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_curr_reg_15__slave ( .q(IR_curr_15), .qb(n343), .d(
        IR_curr_reg_15__m2s), .g(Ctrl__Regs_1__en2), .rb(n41), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_curr_reg_16__master ( .q(IR_curr_reg_16__m2s), .d(n152), 
        .sdi(n343), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n42), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_curr_reg_16__slave ( .q(IR_curr_16), .qb(n342), .d(
        IR_curr_reg_16__m2s), .g(Ctrl__Regs_1__en2), .rb(n42), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_curr_reg_17__master ( .q(IR_curr_reg_17__m2s), .d(n153), 
        .sdi(n342), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n41), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_curr_reg_17__slave ( .q(IR_curr_17), .qb(n341), .d(
        IR_curr_reg_17__m2s), .g(Ctrl__Regs_1__en2), .rb(n41), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_curr_reg_18__master ( .q(IR_curr_reg_18__m2s), .d(n154), 
        .sdi(n341), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n42), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_curr_reg_18__slave ( .q(IR_curr_18), .qb(n340), .d(
        IR_curr_reg_18__m2s), .g(Ctrl__Regs_1__en2), .rb(n42), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_curr_reg_19__master ( .q(IR_curr_reg_19__m2s), .d(n155), 
        .sdi(n340), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n41), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_curr_reg_19__slave ( .q(IR_curr_19), .qb(n339), .d(
        IR_curr_reg_19__m2s), .g(Ctrl__Regs_1__en2), .rb(n41), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_curr_reg_1__master ( .q(IR_curr_reg_1__m2s), .d(n137), .sdi(
        n358), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n41), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_curr_reg_1__slave ( .q(IR_curr_1), .qb(n357), .d(
        IR_curr_reg_1__m2s), .g(Ctrl__Regs_1__en2), .rb(n41), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_curr_reg_20__master ( .q(IR_curr_reg_20__m2s), .d(n156), 
        .sdi(n339), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n41), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_curr_reg_20__slave ( .q(IR_curr_20), .qb(n338), .d(
        IR_curr_reg_20__m2s), .g(Ctrl__Regs_1__en2), .rb(n41), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_curr_reg_21__master ( .q(IR_curr_reg_21__m2s), .d(n157), 
        .sdi(n338), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n42), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_curr_reg_21__slave ( .q(IR_curr_21), .qb(n337), .d(
        IR_curr_reg_21__m2s), .g(Ctrl__Regs_1__en2), .rb(n42), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_curr_reg_22__master ( .q(IR_curr_reg_22__m2s), .d(n158), 
        .sdi(n337), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n41), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_curr_reg_22__slave ( .q(IR_curr_22), .qb(n336), .d(
        IR_curr_reg_22__m2s), .g(Ctrl__Regs_1__en2), .rb(n41), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_curr_reg_23__master ( .q(IR_curr_reg_23__m2s), .d(n159), 
        .sdi(n336), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n42), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_curr_reg_23__slave ( .q(IR_curr_23), .qb(n335), .d(
        IR_curr_reg_23__m2s), .g(Ctrl__Regs_1__en2), .rb(n42), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_curr_reg_24__master ( .q(IR_curr_reg_24__m2s), .d(n160), 
        .sdi(n335), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n41), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_curr_reg_24__slave ( .q(IR_curr_24), .qb(n334), .d(
        IR_curr_reg_24__m2s), .g(Ctrl__Regs_1__en2), .rb(n41), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_curr_reg_25__master ( .q(IR_curr_reg_25__m2s), .d(n161), 
        .sdi(n334), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n42), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_curr_reg_25__slave ( .q(IR_curr_25), .qb(n333), .d(
        IR_curr_reg_25__m2s), .g(Ctrl__Regs_1__en2), .rb(n42), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_curr_reg_26__master ( .q(IR_curr_reg_26__m2s), .d(n162), 
        .sdi(n333), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n41), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_curr_reg_26__slave ( .q(IR_curr_26), .qb(n332), .d(
        IR_curr_reg_26__m2s), .g(Ctrl__Regs_1__en2), .rb(n41), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_curr_reg_27__master ( .q(IR_curr_reg_27__m2s), .d(n163), 
        .sdi(n332), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n42), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_curr_reg_27__slave ( .q(IR_curr_27), .qb(n331), .d(
        IR_curr_reg_27__m2s), .g(Ctrl__Regs_1__en2), .rb(n42), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_curr_reg_28__master ( .q(IR_curr_reg_28__m2s), .d(n164), 
        .sdi(n331), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n41), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_curr_reg_28__slave ( .q(IR_curr_28), .qb(n330), .d(
        IR_curr_reg_28__m2s), .g(Ctrl__Regs_1__en2), .rb(n41), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_curr_reg_29__master ( .q(IR_curr_reg_29__m2s), .d(n165), 
        .sdi(n330), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n42), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_curr_reg_29__slave ( .q(IR_curr_29), .qb(n329), .d(
        IR_curr_reg_29__m2s), .g(Ctrl__Regs_1__en2), .rb(n42), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_curr_reg_2__master ( .q(IR_curr_reg_2__m2s), .d(n138), .sdi(
        n357), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n42), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_curr_reg_2__slave ( .q(IR_curr_2), .qb(n356), .d(
        IR_curr_reg_2__m2s), .g(Ctrl__Regs_1__en2), .rb(n42), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_curr_reg_30__master ( .q(IR_curr_reg_30__m2s), .d(n166), 
        .sdi(n329), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n42), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_curr_reg_30__slave ( .q(IR_curr_30), .qb(n328), .d(
        IR_curr_reg_30__m2s), .g(Ctrl__Regs_1__en2), .rb(n42), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_curr_reg_31__master ( .q(IR_curr_reg_31__m2s), .d(n167), 
        .sdi(n328), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n41), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_curr_reg_31__slave ( .q(IR_curr_31), .qb(n327), .d(
        IR_curr_reg_31__m2s), .g(Ctrl__Regs_1__en2), .rb(n41), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_curr_reg_3__master ( .q(IR_curr_reg_3__m2s), .d(n139), .sdi(
        n356), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n41), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_curr_reg_3__slave ( .q(IR_curr_3), .qb(n355), .d(
        IR_curr_reg_3__m2s), .g(Ctrl__Regs_1__en2), .rb(n41), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_curr_reg_4__master ( .q(IR_curr_reg_4__m2s), .d(n140), .sdi(
        n355), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n42), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_curr_reg_4__slave ( .q(IR_curr_4), .qb(n354), .d(
        IR_curr_reg_4__m2s), .g(Ctrl__Regs_1__en2), .rb(n42), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_curr_reg_5__master ( .q(IR_curr_reg_5__m2s), .d(n141), .sdi(
        n354), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n41), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_curr_reg_5__slave ( .q(IR_curr_5), .qb(n353), .d(
        IR_curr_reg_5__m2s), .g(Ctrl__Regs_1__en2), .rb(n41), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_curr_reg_6__master ( .q(IR_curr_reg_6__m2s), .d(n142), .sdi(
        n353), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n42), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_curr_reg_6__slave ( .q(IR_curr_6), .qb(n352), .d(
        IR_curr_reg_6__m2s), .g(Ctrl__Regs_1__en2), .rb(n42), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_curr_reg_7__master ( .q(IR_curr_reg_7__m2s), .d(n143), .sdi(
        n352), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_curr_reg_7__slave ( .q(IR_curr_7), .qb(n351), .d(
        IR_curr_reg_7__m2s), .g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_curr_reg_8__master ( .q(IR_curr_reg_8__m2s), .d(n144), .sdi(
        n351), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n42), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_curr_reg_8__slave ( .q(IR_curr_8), .qb(n350), .d(
        IR_curr_reg_8__m2s), .g(Ctrl__Regs_1__en2), .rb(n42), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_curr_reg_9__master ( .q(IR_curr_reg_9__m2s), .d(n145), .sdi(
        n350), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_curr_reg_9__slave ( .q(IR_curr_9), .qb(n349), .d(
        IR_curr_reg_9__m2s), .g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_latched_reg_0__master ( .q(IR_latched_reg_0__m2s), .d(N119), 
        .sdi(n327), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_latched_reg_0__slave ( .q(IR_latched[0]), .qb(n326), .d(
        IR_latched_reg_0__m2s), .g(Ctrl__Regs_1__en2), .rb(n38), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_latched_reg_10__master ( .q(IR_latched_reg_10__m2s), .d(N129), 
        .sdi(n317), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_latched_reg_10__slave ( .q(IR_latched[10]), .qb(n316), .d(
        IR_latched_reg_10__m2s), .g(Ctrl__Regs_1__en2), .rb(n38), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_latched_reg_11__master ( .q(IR_latched_reg_11__m2s), .d(N130), 
        .sdi(n316), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_latched_reg_11__slave ( .q(IR_latched[11]), .qb(n315), .d(
        IR_latched_reg_11__m2s), .g(Ctrl__Regs_1__en2), .rb(n38), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_latched_reg_12__master ( .q(IR_latched_reg_12__m2s), .d(N131), 
        .sdi(n315), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_latched_reg_12__slave ( .q(IR_latched[12]), .qb(n314), .d(
        IR_latched_reg_12__m2s), .g(Ctrl__Regs_1__en2), .rb(n38), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_latched_reg_13__master ( .q(IR_latched_reg_13__m2s), .d(N132), 
        .sdi(n314), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_latched_reg_13__slave ( .q(IR_latched[13]), .qb(n313), .d(
        IR_latched_reg_13__m2s), .g(Ctrl__Regs_1__en2), .rb(n38), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_latched_reg_14__master ( .q(IR_latched_reg_14__m2s), .d(N133), 
        .sdi(n313), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_latched_reg_14__slave ( .q(IR_latched[14]), .qb(n312), .d(
        IR_latched_reg_14__m2s), .g(Ctrl__Regs_1__en2), .rb(n38), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_latched_reg_15__master ( .q(IR_latched_reg_15__m2s), .d(N134), 
        .sdi(n312), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_latched_reg_15__slave ( .q(IR_latched[15]), .qb(n311), .d(
        IR_latched_reg_15__m2s), .g(Ctrl__Regs_1__en2), .rb(n38), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_latched_reg_16__master ( .q(IR_latched_reg_16__m2s), .d(N135), 
        .sdi(n311), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n37), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_latched_reg_16__slave ( .q(IR_latched[16]), .qb(n310), .d(
        IR_latched_reg_16__m2s), .g(Ctrl__Regs_1__en2), .rb(n37), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_latched_reg_17__master ( .q(IR_latched_reg_17__m2s), .d(N136), 
        .sdi(n310), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n37), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_latched_reg_17__slave ( .q(IR_latched[17]), .qb(n309), .d(
        IR_latched_reg_17__m2s), .g(Ctrl__Regs_1__en2), .rb(n37), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_latched_reg_18__master ( .q(IR_latched_reg_18__m2s), .d(N137), 
        .sdi(n309), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n37), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_latched_reg_18__slave ( .q(IR_latched[18]), .qb(n308), .d(
        IR_latched_reg_18__m2s), .g(Ctrl__Regs_1__en2), .rb(n37), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_latched_reg_19__master ( .q(IR_latched_reg_19__m2s), .d(N138), 
        .sdi(n308), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n37), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_latched_reg_19__slave ( .q(IR_latched[19]), .qb(n307), .d(
        IR_latched_reg_19__m2s), .g(Ctrl__Regs_1__en2), .rb(n37), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_latched_reg_1__master ( .q(IR_latched_reg_1__m2s), .d(N120), 
        .sdi(n326), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_latched_reg_1__slave ( .q(IR_latched[1]), .qb(n325), .d(
        IR_latched_reg_1__m2s), .g(Ctrl__Regs_1__en2), .rb(n38), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_latched_reg_20__master ( .q(IR_latched_reg_20__m2s), .d(N139), 
        .sdi(n307), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n37), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_latched_reg_20__slave ( .q(IR_latched[20]), .qb(n306), .d(
        IR_latched_reg_20__m2s), .g(Ctrl__Regs_1__en2), .rb(n37), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_latched_reg_21__master ( .q(IR_latched_reg_21__m2s), .d(N140), 
        .sdi(n306), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n37), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_latched_reg_21__slave ( .q(IR_latched[21]), .qb(n305), .d(
        IR_latched_reg_21__m2s), .g(Ctrl__Regs_1__en2), .rb(n37), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_latched_reg_22__master ( .q(IR_latched_reg_22__m2s), .d(N141), 
        .sdi(n305), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n37), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_latched_reg_22__slave ( .q(IR_latched[22]), .qb(n304), .d(
        IR_latched_reg_22__m2s), .g(Ctrl__Regs_1__en2), .rb(n37), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_latched_reg_23__master ( .q(IR_latched_reg_23__m2s), .d(N142), 
        .sdi(n304), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n37), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_latched_reg_23__slave ( .q(IR_latched[23]), .qb(n303), .d(
        IR_latched_reg_23__m2s), .g(Ctrl__Regs_1__en2), .rb(n37), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_latched_reg_24__master ( .q(IR_latched_reg_24__m2s), .d(N143), 
        .sdi(n303), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n37), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_latched_reg_24__slave ( .q(IR_latched[24]), .qb(n302), .d(
        IR_latched_reg_24__m2s), .g(Ctrl__Regs_1__en2), .rb(n37), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_latched_reg_25__master ( .q(IR_latched_reg_25__m2s), .d(N144), 
        .sdi(n302), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n37), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_latched_reg_25__slave ( .q(IR_latched[25]), .qb(n301), .d(
        IR_latched_reg_25__m2s), .g(Ctrl__Regs_1__en2), .rb(n37), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_latched_reg_26__master ( .q(IR_latched_reg_26__m2s), .d(N145), 
        .sdi(n301), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n37), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_latched_reg_26__slave ( .q(IR_latched[26]), .qb(n300), .d(
        IR_latched_reg_26__m2s), .g(Ctrl__Regs_1__en2), .rb(n37), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_latched_reg_27__master ( .q(IR_latched_reg_27__m2s), .d(N146), 
        .sdi(n300), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n37), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_latched_reg_27__slave ( .q(IR_latched[27]), .qb(n299), .d(
        IR_latched_reg_27__m2s), .g(Ctrl__Regs_1__en2), .rb(n37), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_latched_reg_28__master ( .q(IR_latched_reg_28__m2s), .d(N147), 
        .sdi(n299), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n37), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_latched_reg_28__slave ( .q(IR_latched[28]), .qb(n298), .d(
        IR_latched_reg_28__m2s), .g(Ctrl__Regs_1__en2), .rb(n37), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_latched_reg_29__master ( .q(IR_latched_reg_29__m2s), .d(N148), 
        .sdi(n298), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n37), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_latched_reg_29__slave ( .q(IR_latched[29]), .qb(n297), .d(
        IR_latched_reg_29__m2s), .g(Ctrl__Regs_1__en2), .rb(n37), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_latched_reg_2__master ( .q(IR_latched_reg_2__m2s), .d(N121), 
        .sdi(n325), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_latched_reg_2__slave ( .q(IR_latched[2]), .qb(n324), .d(
        IR_latched_reg_2__m2s), .g(Ctrl__Regs_1__en2), .rb(n38), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_latched_reg_30__master ( .q(IR_latched_reg_30__m2s), .d(N149), 
        .sdi(n297), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n37), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_latched_reg_30__slave ( .q(IR_latched[30]), .qb(n296), .d(
        IR_latched_reg_30__m2s), .g(Ctrl__Regs_1__en2), .rb(n37), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_latched_reg_31__master ( .q(IR_latched_reg_31__m2s), .d(N150), 
        .sdi(n296), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n37), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_latched_reg_31__slave ( .q(IR_latched[31]), .qb(n295), .d(
        IR_latched_reg_31__m2s), .g(Ctrl__Regs_1__en2), .rb(n37), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_latched_reg_3__master ( .q(IR_latched_reg_3__m2s), .d(N122), 
        .sdi(n324), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_latched_reg_3__slave ( .q(IR_latched[3]), .qb(n323), .d(
        IR_latched_reg_3__m2s), .g(Ctrl__Regs_1__en2), .rb(n38), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_latched_reg_4__master ( .q(IR_latched_reg_4__m2s), .d(N123), 
        .sdi(n323), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_latched_reg_4__slave ( .q(IR_latched[4]), .qb(n322), .d(
        IR_latched_reg_4__m2s), .g(Ctrl__Regs_1__en2), .rb(n38), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_latched_reg_5__master ( .q(IR_latched_reg_5__m2s), .d(N124), 
        .sdi(n322), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_latched_reg_5__slave ( .q(IR_latched[5]), .qb(n321), .d(
        IR_latched_reg_5__m2s), .g(Ctrl__Regs_1__en2), .rb(n38), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_latched_reg_6__master ( .q(IR_latched_reg_6__m2s), .d(N125), 
        .sdi(n321), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_latched_reg_6__slave ( .q(IR_latched[6]), .qb(n320), .d(
        IR_latched_reg_6__m2s), .g(Ctrl__Regs_1__en2), .rb(n38), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_latched_reg_7__master ( .q(IR_latched_reg_7__m2s), .d(N126), 
        .sdi(n320), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_latched_reg_7__slave ( .q(IR_latched[7]), .qb(n319), .d(
        IR_latched_reg_7__m2s), .g(Ctrl__Regs_1__en2), .rb(n38), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_latched_reg_8__master ( .q(IR_latched_reg_8__m2s), .d(N127), 
        .sdi(n319), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_latched_reg_8__slave ( .q(IR_latched[8]), .qb(n318), .d(
        IR_latched_reg_8__m2s), .g(Ctrl__Regs_1__en2), .rb(n38), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_latched_reg_9__master ( .q(IR_latched_reg_9__m2s), .d(N128), 
        .sdi(n318), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_latched_reg_9__slave ( .q(IR_latched[9]), .qb(n317), .d(
        IR_latched_reg_9__m2s), .g(Ctrl__Regs_1__en2), .rb(n38), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_previous_reg_0__master ( .q(IR_previous_reg_0__m2s), .d(n104), 
        .sdi(n295), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n42), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_previous_reg_0__slave ( .q(IR_previous_0), .qb(n294), .d(
        IR_previous_reg_0__m2s), .g(Ctrl__Regs_1__en2), .rb(n42), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_previous_reg_10__master ( .q(IR_previous_reg_10__m2s), .d(
        n114), .sdi(n285), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n42), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_previous_reg_10__slave ( .q(IR_previous_10), .qb(n284), .d(
        IR_previous_reg_10__m2s), .g(Ctrl__Regs_1__en2), .rb(n42), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_previous_reg_11__master ( .q(IR_previous_reg_11__m2s), .d(
        n115), .sdi(n284), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_previous_reg_11__slave ( .q(IR_previous_11), .qb(n283), .d(
        IR_previous_reg_11__m2s), .g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_previous_reg_12__master ( .q(IR_previous_reg_12__m2s), .d(
        n116), .sdi(n283), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n42), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_previous_reg_12__slave ( .q(IR_previous_12), .qb(n282), .d(
        IR_previous_reg_12__m2s), .g(Ctrl__Regs_1__en2), .rb(n42), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_previous_reg_13__master ( .q(IR_previous_reg_13__m2s), .d(
        n117), .sdi(n282), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_previous_reg_13__slave ( .q(IR_previous_13), .qb(n281), .d(
        IR_previous_reg_13__m2s), .g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_previous_reg_14__master ( .q(IR_previous_reg_14__m2s), .d(
        n118), .sdi(n281), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n42), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_previous_reg_14__slave ( .q(IR_previous_14), .qb(n280), .d(
        IR_previous_reg_14__m2s), .g(Ctrl__Regs_1__en2), .rb(n42), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_previous_reg_15__master ( .q(IR_previous_reg_15__m2s), .d(
        n119), .sdi(n280), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_previous_reg_15__slave ( .q(IR_previous_15), .qb(n279), .d(
        IR_previous_reg_15__m2s), .g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_previous_reg_16__master ( .q(IR_previous_reg_16__m2s), .d(
        n120), .sdi(n279), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n43), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_previous_reg_16__slave ( .q(IR_previous_16), .qb(n278), .d(
        IR_previous_reg_16__m2s), .g(Ctrl__Regs_1__en2), .rb(n43), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_previous_reg_17__master ( .q(IR_previous_reg_17__m2s), .d(
        n121), .sdi(n278), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_previous_reg_17__slave ( .q(IR_previous_17), .qb(n277), .d(
        IR_previous_reg_17__m2s), .g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_previous_reg_18__master ( .q(IR_previous_reg_18__m2s), .d(
        n122), .sdi(n277), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n43), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_previous_reg_18__slave ( .q(IR_previous_18), .qb(n276), .d(
        IR_previous_reg_18__m2s), .g(Ctrl__Regs_1__en2), .rb(n43), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_previous_reg_19__master ( .q(IR_previous_reg_19__m2s), .d(
        n123), .sdi(n276), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_previous_reg_19__slave ( .q(IR_previous_19), .qb(n275), .d(
        IR_previous_reg_19__m2s), .g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_previous_reg_1__master ( .q(IR_previous_reg_1__m2s), .d(n105), 
        .sdi(n294), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_previous_reg_1__slave ( .q(IR_previous_1), .qb(n293), .d(
        IR_previous_reg_1__m2s), .g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_previous_reg_20__master ( .q(IR_previous_reg_20__m2s), .d(
        n124), .sdi(n275), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_previous_reg_20__slave ( .q(IR_previous_20), .qb(n274), .d(
        IR_previous_reg_20__m2s), .g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_previous_reg_21__master ( .q(IR_previous_reg_21__m2s), .d(
        n125), .sdi(n274), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n43), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_previous_reg_21__slave ( .q(IR_previous_21), .qb(n273), .d(
        IR_previous_reg_21__m2s), .g(Ctrl__Regs_1__en2), .rb(n43), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_previous_reg_22__master ( .q(IR_previous_reg_22__m2s), .d(
        n126), .sdi(n273), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_previous_reg_22__slave ( .q(IR_previous_22), .qb(n272), .d(
        IR_previous_reg_22__m2s), .g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_previous_reg_23__master ( .q(IR_previous_reg_23__m2s), .d(
        n127), .sdi(n272), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n43), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_previous_reg_23__slave ( .q(IR_previous_23), .qb(n271), .d(
        IR_previous_reg_23__m2s), .g(Ctrl__Regs_1__en2), .rb(n43), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_previous_reg_24__master ( .q(IR_previous_reg_24__m2s), .d(
        n128), .sdi(n271), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_previous_reg_24__slave ( .q(IR_previous_24), .qb(n270), .d(
        IR_previous_reg_24__m2s), .g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_previous_reg_25__master ( .q(IR_previous_reg_25__m2s), .d(
        n129), .sdi(n270), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n43), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_previous_reg_25__slave ( .q(IR_previous_25), .qb(n269), .d(
        IR_previous_reg_25__m2s), .g(Ctrl__Regs_1__en2), .rb(n43), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_previous_reg_26__master ( .q(IR_previous_reg_26__m2s), .d(
        n130), .sdi(n269), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_previous_reg_26__slave ( .q(IR_previous_26), .qb(n268), .d(
        IR_previous_reg_26__m2s), .g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_previous_reg_27__master ( .q(IR_previous_reg_27__m2s), .d(
        n131), .sdi(n268), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n43), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_previous_reg_27__slave ( .q(IR_previous_27), .qb(n267), .d(
        IR_previous_reg_27__m2s), .g(Ctrl__Regs_1__en2), .rb(n43), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_previous_reg_28__master ( .q(IR_previous_reg_28__m2s), .d(
        n132), .sdi(n267), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_previous_reg_28__slave ( .q(IR_previous_28), .qb(n266), .d(
        IR_previous_reg_28__m2s), .g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_previous_reg_29__master ( .q(IR_previous_reg_29__m2s), .d(
        n133), .sdi(n266), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n43), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_previous_reg_29__slave ( .q(IR_previous_29), .qb(n265), .d(
        IR_previous_reg_29__m2s), .g(Ctrl__Regs_1__en2), .rb(n43), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_previous_reg_2__master ( .q(IR_previous_reg_2__m2s), .d(n106), 
        .sdi(n293), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n43), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_previous_reg_2__slave ( .q(IR_previous_2), .qb(n292), .d(
        IR_previous_reg_2__m2s), .g(Ctrl__Regs_1__en2), .rb(n43), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_previous_reg_30__master ( .q(IR_previous_reg_30__m2s), .d(
        n134), .sdi(n265), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n43), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_previous_reg_30__slave ( .q(IR_previous_30), .qb(n264), .d(
        IR_previous_reg_30__m2s), .g(Ctrl__Regs_1__en2), .rb(n43), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_previous_reg_31__master ( .q(IR_previous_reg_31__m2s), .d(
        n135), .sdi(n264), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40), 
        .glob_g(global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_previous_reg_31__slave ( .q(IR_previous_31), .qb(n263), .d(
        IR_previous_reg_31__m2s), .g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_previous_reg_3__master ( .q(IR_previous_reg_3__m2s), .d(n107), 
        .sdi(n292), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_previous_reg_3__slave ( .q(IR_previous_3), .qb(n291), .d(
        IR_previous_reg_3__m2s), .g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_previous_reg_4__master ( .q(IR_previous_reg_4__m2s), .d(n108), 
        .sdi(n291), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n43), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_previous_reg_4__slave ( .q(IR_previous_4), .qb(n290), .d(
        IR_previous_reg_4__m2s), .g(Ctrl__Regs_1__en2), .rb(n43), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_previous_reg_5__master ( .q(IR_previous_reg_5__m2s), .d(n109), 
        .sdi(n290), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_previous_reg_5__slave ( .q(IR_previous_5), .qb(n289), .d(
        IR_previous_reg_5__m2s), .g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_previous_reg_6__master ( .q(IR_previous_reg_6__m2s), .d(n110), 
        .sdi(n289), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n43), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_previous_reg_6__slave ( .q(IR_previous_6), .qb(n288), .d(
        IR_previous_reg_6__m2s), .g(Ctrl__Regs_1__en2), .rb(n43), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_previous_reg_7__master ( .q(IR_previous_reg_7__m2s), .d(n111), 
        .sdi(n288), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_previous_reg_7__slave ( .q(IR_previous_7), .qb(n287), .d(
        IR_previous_reg_7__m2s), .g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_previous_reg_8__master ( .q(IR_previous_reg_8__m2s), .d(n112), 
        .sdi(n287), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n43), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_previous_reg_8__slave ( .q(IR_previous_8), .qb(n286), .d(
        IR_previous_reg_8__m2s), .g(Ctrl__Regs_1__en2), .rb(n43), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 IR_previous_reg_9__master ( .q(IR_previous_reg_9__m2s), .d(n113), 
        .sdi(n286), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n39), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 IR_previous_reg_9__slave ( .q(IR_previous_9), .qb(n285), .d(
        IR_previous_reg_9__m2s), .g(Ctrl__Regs_1__en2), .rb(n39), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_2 NPC_reg_0__master ( .q(NPC_reg_0__m2s), .d(N87), .sdi(n263), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n36), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_8 NPC_reg_0__slave ( .q(NPC[0]), .qb(n262), .d(NPC_reg_0__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n36), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 NPC_reg_10__master ( .q(NPC_reg_10__m2s), .d(N97), .sdi(n22), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n36), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_4 NPC_reg_10__slave ( .q(NPC[10]), .qb(n24), .d(NPC_reg_10__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n36), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 NPC_reg_11__master ( .q(NPC_reg_11__m2s), .d(N98), .sdi(n24), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n36), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 NPC_reg_11__slave ( .q(n205), .qb(n257), .d(NPC_reg_11__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n36), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 NPC_reg_12__master ( .q(NPC_reg_12__m2s), .d(N99), .sdi(n257), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n36), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 NPC_reg_12__slave ( .q(NPC[12]), .qb(n28), .d(NPC_reg_12__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n36), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_2 NPC_reg_13__master ( .q(NPC_reg_13__m2s), .d(N100), .sdi(n28), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n36), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_8 NPC_reg_13__slave ( .q(NPC[13]), .qb(n14), .d(NPC_reg_13__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n36), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 NPC_reg_14__master ( .q(NPC_reg_14__m2s), .d(N101), .sdi(n14), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n36), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_4 NPC_reg_14__slave ( .q(n360), .qb(n12), .d(NPC_reg_14__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n36), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 NPC_reg_15__master ( .q(NPC_reg_15__m2s), .d(N102), .sdi(n12), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n36), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 NPC_reg_15__slave ( .q(n204), .qb(n256), .d(NPC_reg_15__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n36), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_2 NPC_reg_16__master ( .q(NPC_reg_16__m2s), .d(N103), .sdi(n256), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n36), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_8 NPC_reg_16__slave ( .q(NPC[16]), .qb(n255), .d(NPC_reg_16__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n36), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_2 NPC_reg_17__master ( .q(NPC_reg_17__m2s), .d(N104), .sdi(n255), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n36), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_8 NPC_reg_17__slave ( .q(NPC[17]), .qb(n10), .d(NPC_reg_17__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n36), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_2 NPC_reg_18__master ( .q(NPC_reg_18__m2s), .d(N105), .sdi(n10), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n36), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_8 NPC_reg_18__slave ( .q(NPC[18]), .qb(n254), .d(NPC_reg_18__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n36), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_2 NPC_reg_19__master ( .q(NPC_reg_19__m2s), .d(N106), .sdi(n254), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_8 NPC_reg_19__slave ( .q(NPC[19]), .qb(n253), .d(NPC_reg_19__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_2 NPC_reg_1__master ( .q(NPC_reg_1__m2s), .d(N88), .sdi(n262), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n36), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_8 NPC_reg_1__slave ( .q(NPC[1]), .qb(n261), .d(NPC_reg_1__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n36), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_2 NPC_reg_20__master ( .q(NPC_reg_20__m2s), .d(N107), .sdi(n253), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_8 NPC_reg_20__slave ( .q(NPC[20]), .qb(n252), .d(NPC_reg_20__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_2 NPC_reg_21__master ( .q(NPC_reg_21__m2s), .d(N108), .sdi(n252), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_8 NPC_reg_21__slave ( .q(NPC[21]), .qb(n251), .d(NPC_reg_21__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_2 NPC_reg_22__master ( .q(NPC_reg_22__m2s), .d(N109), .sdi(n251), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_8 NPC_reg_22__slave ( .q(NPC[22]), .qb(n250), .d(NPC_reg_22__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_2 NPC_reg_23__master ( .q(NPC_reg_23__m2s), .d(N110), .sdi(n250), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_8 NPC_reg_23__slave ( .q(NPC[23]), .qb(n249), .d(NPC_reg_23__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 NPC_reg_24__master ( .q(NPC_reg_24__m2s), .d(N111), .sdi(n249), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n91), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_4 NPC_reg_24__slave ( .q(NPC[24]), .qb(n248), .d(NPC_reg_24__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n91), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 NPC_reg_25__master ( .q(NPC_reg_25__m2s), .d(N112), .sdi(n248), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_4 NPC_reg_25__slave ( .q(NPC[25]), .qb(n247), .d(NPC_reg_25__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 NPC_reg_26__master ( .q(NPC_reg_26__m2s), .d(N113), .sdi(n247), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 NPC_reg_26__slave ( .q(NPC[26]), .qb(n246), .d(NPC_reg_26__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 NPC_reg_27__master ( .q(NPC_reg_27__m2s), .d(N114), .sdi(n246), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 NPC_reg_27__slave ( .q(NPC[27]), .qb(n245), .d(NPC_reg_27__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 NPC_reg_28__master ( .q(NPC_reg_28__m2s), .d(N115), .sdi(n245), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 NPC_reg_28__slave ( .q(NPC[28]), .qb(n244), .d(NPC_reg_28__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 NPC_reg_29__master ( .q(NPC_reg_29__m2s), .d(N116), .sdi(n244), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 NPC_reg_29__slave ( .q(NPC[29]), .qb(n243), .d(NPC_reg_29__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 NPC_reg_2__master ( .q(NPC_reg_2__m2s), .d(N89), .sdi(n261), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_4 NPC_reg_2__slave ( .q(n210), .qb(n32), .d(NPC_reg_2__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n40), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 NPC_reg_30__master ( .q(NPC_reg_30__m2s), .d(N117), .sdi(n243), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 NPC_reg_30__slave ( .q(NPC[30]), .qb(n242), .d(NPC_reg_30__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(global_g2), .sync_sel(
        sync_sel) );
    smlatnr_1 NPC_reg_31__master ( .q(NPC_reg_31__m2s), .d(N118), .sdi(
        test_si2), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 NPC_reg_31__slave ( .q(NPC[31]), .d(NPC_reg_31__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n40), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 NPC_reg_3__master ( .q(NPC_reg_3__m2s), .d(N90), .sdi(n32), .se(
        test_se), .g(Ctrl__Regs_1__en1), .rb(n40), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_4 NPC_reg_3__slave ( .q(n209), .qb(n30), .d(NPC_reg_3__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n40), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 NPC_reg_4__master ( .q(NPC_reg_4__m2s), .d(N91), .sdi(n30), .se(
        test_se), .g(Ctrl__Regs_1__en1), .rb(n40), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 NPC_reg_4__slave ( .q(n208), .qb(n260), .d(NPC_reg_4__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n40), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 NPC_reg_5__master ( .q(NPC_reg_5__m2s), .d(N92), .sdi(n260), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n36), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_4 NPC_reg_5__slave ( .q(n207), .qb(n259), .d(NPC_reg_5__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n36), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 NPC_reg_6__master ( .q(NPC_reg_6__m2s), .d(N93), .sdi(n259), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n36), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_4 NPC_reg_6__slave ( .q(n206), .qb(n258), .d(NPC_reg_6__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n36), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 NPC_reg_7__master ( .q(NPC_reg_7__m2s), .d(N94), .sdi(n258), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n36), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_4 NPC_reg_7__slave ( .q(NPC[7]), .qb(n26), .d(NPC_reg_7__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n36), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_2 NPC_reg_8__master ( .q(NPC_reg_8__m2s), .d(N95), .sdi(n26), .se(
        test_se), .g(Ctrl__Regs_1__en1), .rb(n36), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_8 NPC_reg_8__slave ( .q(NPC[8]), .qb(n16), .d(NPC_reg_8__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n36), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_2 NPC_reg_9__master ( .q(NPC_reg_9__m2s), .d(N96), .sdi(n16), .se(
        test_se), .g(Ctrl__Regs_1__en1), .rb(n36), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_8 NPC_reg_9__slave ( .q(NPC[9]), .qb(n22), .d(NPC_reg_9__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n36), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 PC_reg_0__master ( .q(PC_reg_0__m2s), .d(n168), .sdi(n242), .se(
        test_se), .g(Ctrl__Regs_1__en1), .rb(n43), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 PC_reg_0__slave ( .q(PC[0]), .qb(n241), .d(PC_reg_0__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n43), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 PC_reg_10__master ( .q(PC_reg_10__m2s), .d(n178), .sdi(n232), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n43), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 PC_reg_10__slave ( .q(PC[10]), .qb(n231), .d(PC_reg_10__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n43), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 PC_reg_11__master ( .q(PC_reg_11__m2s), .d(n179), .sdi(n231), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n39), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 PC_reg_11__slave ( .q(PC[11]), .qb(n230), .d(PC_reg_11__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n39), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 PC_reg_12__master ( .q(PC_reg_12__m2s), .d(n180), .sdi(n230), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n43), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 PC_reg_12__slave ( .q(PC[12]), .qb(n229), .d(PC_reg_12__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n43), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 PC_reg_13__master ( .q(PC_reg_13__m2s), .d(n181), .sdi(n229), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n39), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 PC_reg_13__slave ( .q(PC[13]), .qb(n228), .d(PC_reg_13__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n39), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 PC_reg_14__master ( .q(PC_reg_14__m2s), .d(n182), .sdi(n228), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n43), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 PC_reg_14__slave ( .q(PC[14]), .qb(n227), .d(PC_reg_14__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n43), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 PC_reg_15__master ( .q(PC_reg_15__m2s), .d(n183), .sdi(n227), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n39), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 PC_reg_15__slave ( .q(PC[15]), .qb(n226), .d(PC_reg_15__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n39), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 PC_reg_16__master ( .q(PC_reg_16__m2s), .d(n184), .sdi(n226), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n43), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 PC_reg_16__slave ( .q(PC[16]), .qb(n225), .d(PC_reg_16__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n43), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 PC_reg_17__master ( .q(PC_reg_17__m2s), .d(n185), .sdi(n225), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n39), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 PC_reg_17__slave ( .q(PC[17]), .qb(n224), .d(PC_reg_17__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n39), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 PC_reg_18__master ( .q(PC_reg_18__m2s), .d(n186), .sdi(n224), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 PC_reg_18__slave ( .q(PC[18]), .qb(n223), .d(PC_reg_18__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n38), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 PC_reg_19__master ( .q(PC_reg_19__m2s), .d(n187), .sdi(n223), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n39), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 PC_reg_19__slave ( .q(PC[19]), .qb(n222), .d(PC_reg_19__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n39), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 PC_reg_1__master ( .q(PC_reg_1__m2s), .d(n169), .sdi(n241), .se(
        test_se), .g(Ctrl__Regs_1__en1), .rb(n39), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 PC_reg_1__slave ( .q(PC[1]), .qb(n240), .d(PC_reg_1__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n39), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 PC_reg_20__master ( .q(PC_reg_20__m2s), .d(n188), .sdi(n222), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n39), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 PC_reg_20__slave ( .q(PC[20]), .qb(n221), .d(PC_reg_20__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n39), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 PC_reg_21__master ( .q(PC_reg_21__m2s), .d(n189), .sdi(n221), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 PC_reg_21__slave ( .q(PC[21]), .qb(n92), .d(PC_reg_21__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n38), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 PC_reg_22__master ( .q(PC_reg_22__m2s), .d(n190), .sdi(PC[21]), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n39), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 PC_reg_22__slave ( .q(PC[22]), .qb(n93), .d(PC_reg_22__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n39), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 PC_reg_23__master ( .q(PC_reg_23__m2s), .d(n191), .sdi(PC[22]), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 PC_reg_23__slave ( .q(PC[23]), .qb(n94), .d(PC_reg_23__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n38), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 PC_reg_24__master ( .q(PC_reg_24__m2s), .d(n192), .sdi(PC[23]), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n39), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 PC_reg_24__slave ( .q(PC[24]), .qb(n95), .d(PC_reg_24__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n39), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 PC_reg_25__master ( .q(PC_reg_25__m2s), .d(n193), .sdi(PC[24]), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 PC_reg_25__slave ( .q(PC[25]), .qb(n96), .d(PC_reg_25__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n38), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 PC_reg_26__master ( .q(PC_reg_26__m2s), .d(n194), .sdi(PC[25]), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n39), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 PC_reg_26__slave ( .q(PC[26]), .qb(n97), .d(PC_reg_26__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n39), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 PC_reg_27__master ( .q(PC_reg_27__m2s), .d(n195), .sdi(PC[26]), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 PC_reg_27__slave ( .q(PC[27]), .qb(n98), .d(PC_reg_27__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n38), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 PC_reg_28__master ( .q(PC_reg_28__m2s), .d(n196), .sdi(PC[27]), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n39), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 PC_reg_28__slave ( .q(PC[28]), .qb(n99), .d(PC_reg_28__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n39), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 PC_reg_29__master ( .q(PC_reg_29__m2s), .d(n197), .sdi(PC[28]), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 PC_reg_29__slave ( .q(PC[29]), .qb(n100), .d(PC_reg_29__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n38), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 PC_reg_2__master ( .q(PC_reg_2__m2s), .d(n170), .sdi(n240), .se(
        test_se), .g(Ctrl__Regs_1__en1), .rb(n38), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 PC_reg_2__slave ( .q(PC[2]), .qb(n239), .d(PC_reg_2__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n38), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 PC_reg_30__master ( .q(PC_reg_30__m2s), .d(n198), .sdi(PC[29]), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 PC_reg_30__slave ( .q(PC[30]), .qb(n101), .d(PC_reg_30__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n38), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 PC_reg_31__master ( .q(PC_reg_31__m2s), .d(n199), .sdi(PC[30]), 
        .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n39), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 PC_reg_31__slave ( .q(PC[31]), .qb(n102), .d(PC_reg_31__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n39), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 PC_reg_3__master ( .q(PC_reg_3__m2s), .d(n171), .sdi(n239), .se(
        test_se), .g(Ctrl__Regs_1__en1), .rb(n39), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 PC_reg_3__slave ( .q(PC[3]), .qb(n238), .d(PC_reg_3__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n39), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 PC_reg_4__master ( .q(PC_reg_4__m2s), .d(n172), .sdi(n238), .se(
        test_se), .g(Ctrl__Regs_1__en1), .rb(n38), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 PC_reg_4__slave ( .q(PC[4]), .qb(n237), .d(PC_reg_4__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n38), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 PC_reg_5__master ( .q(PC_reg_5__m2s), .d(n173), .sdi(n237), .se(
        test_se), .g(Ctrl__Regs_1__en1), .rb(n39), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 PC_reg_5__slave ( .q(PC[5]), .qb(n236), .d(PC_reg_5__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n39), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 PC_reg_6__master ( .q(PC_reg_6__m2s), .d(n174), .sdi(n236), .se(
        test_se), .g(Ctrl__Regs_1__en1), .rb(n38), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 PC_reg_6__slave ( .q(PC[6]), .qb(n235), .d(PC_reg_6__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n38), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 PC_reg_7__master ( .q(PC_reg_7__m2s), .d(n175), .sdi(n235), .se(
        test_se), .g(Ctrl__Regs_1__en1), .rb(n39), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 PC_reg_7__slave ( .q(PC[7]), .qb(n234), .d(PC_reg_7__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n39), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 PC_reg_8__master ( .q(PC_reg_8__m2s), .d(n176), .sdi(n234), .se(
        test_se), .g(Ctrl__Regs_1__en1), .rb(n38), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 PC_reg_8__slave ( .q(PC[8]), .qb(n233), .d(PC_reg_8__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n38), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    smlatnr_1 PC_reg_9__master ( .q(PC_reg_9__m2s), .d(n177), .sdi(n233), .se(
        test_se), .g(Ctrl__Regs_1__en1), .rb(n39), .glob_g(global_g1), 
        .sync_sel(sync_sel) );
    mlatnr_2 PC_reg_9__slave ( .q(PC[9]), .qb(n232), .d(PC_reg_9__m2s), .g(
        Ctrl__Regs_1__en2), .rb(n39), .glob_g(global_g2), .sync_sel(sync_sel)
         );
    nand2_2 U10 ( .x(n48), .a(branch_address[22]), .b(branch_sig) );
    mux2_2 U100 ( .x(n163), .d0(IR_curr_27), .sl(n87), .d1(IR[27]) );
    mux2_2 U101 ( .x(n164), .d0(IR_curr_28), .sl(n87), .d1(IR[28]) );
    mux2_2 U102 ( .x(n165), .d0(IR_curr_29), .sl(n87), .d1(IR[29]) );
    buf_3 U103 ( .x(n42), .a(n91) );
    mux2_2 U104 ( .x(n166), .d0(IR_curr_30), .sl(n87), .d1(IR[30]) );
    buf_3 U105 ( .x(n41), .a(n91) );
    inv_2 U106 ( .x(n81), .a(counter[0]) );
    inv_2 U107 ( .x(n83), .a(counter[1]) );
    mux2_2 U108 ( .x(n168), .d0(PC[0]), .sl(n89), .d1(n218) );
    mux2_2 U109 ( .x(n169), .d0(PC[1]), .sl(n89), .d1(NPC[1]) );
    nand2i_2 U11 ( .x(n49), .a(n93), .b(N152) );
    mux2_2 U110 ( .x(n170), .d0(PC[2]), .sl(n89), .d1(n33) );
    mux2_2 U111 ( .x(n171), .d0(PC[3]), .sl(n90), .d1(n31) );
    buf_3 U112 ( .x(n43), .a(n91) );
    mux2_3 U113 ( .x(n186), .d0(PC[18]), .sl(n89), .d1(NPC[18]) );
    mux2_3 U114 ( .x(n187), .d0(PC[19]), .sl(n90), .d1(NPC[19]) );
    mux2_3 U115 ( .x(n188), .d0(PC[20]), .sl(n89), .d1(NPC[20]) );
    mux2_2 U116 ( .x(n189), .d0(PC[21]), .sl(n90), .d1(n214) );
    mux2_2 U117 ( .x(n190), .d0(PC[22]), .sl(n90), .d1(NPC[22]) );
    mux2_2 U118 ( .x(n191), .d0(PC[23]), .sl(n89), .d1(NPC[23]) );
    mux2_2 U119 ( .x(n192), .d0(PC[24]), .sl(n90), .d1(NPC[24]) );
    ao222_1 U12 ( .x(N150), .a(IR_previous_31), .b(N152), .c(IR_curr_31), .d(
        n4), .e(IR[31]), .f(n202) );
    mux2_3 U120 ( .x(n193), .d0(PC[25]), .sl(n89), .d1(NPC[25]) );
    mux2_2 U121 ( .x(n194), .d0(PC[26]), .sl(n89), .d1(NPC[26]) );
    mux2_2 U122 ( .x(n195), .d0(PC[27]), .sl(n90), .d1(NPC[27]) );
    mux2_2 U123 ( .x(n196), .d0(PC[28]), .sl(n90), .d1(NPC[28]) );
    mux2_2 U124 ( .x(n197), .d0(PC[29]), .sl(n89), .d1(NPC[29]) );
    mux2_2 U125 ( .x(n198), .d0(PC[30]), .sl(n89), .d1(NPC[30]) );
    buf_3 U126 ( .x(n39), .a(n91) );
    mux2_2 U127 ( .x(n199), .d0(PC[31]), .sl(n89), .d1(NPC[31]) );
    oai21_1 U128 ( .x(n200), .a(n90), .b(test_so1), .c(n88) );
    ao222_1 U129 ( .x(N119), .a(IR_previous_0), .b(n5), .c(IR_curr_0), .d(n4), 
        .e(IR[0]), .f(n202) );
    ao222_1 U13 ( .x(N148), .a(IR_previous_29), .b(N152), .c(IR_curr_29), .d(
        n4), .e(IR[29]), .f(n202) );
    ao222_1 U130 ( .x(N120), .a(IR_previous_1), .b(n5), .c(IR_curr_1), .d(n4), 
        .e(IR[1]), .f(n202) );
    ao222_1 U131 ( .x(N121), .a(IR_previous_2), .b(n5), .c(IR_curr_2), .d(n4), 
        .e(IR[2]), .f(n202) );
    ao222_1 U132 ( .x(N122), .a(IR_previous_3), .b(n5), .c(IR_curr_3), .d(n4), 
        .e(IR[3]), .f(n202) );
    ao222_1 U133 ( .x(N123), .a(IR_previous_4), .b(n5), .c(IR_curr_4), .d(n4), 
        .e(IR[4]), .f(n202) );
    ao222_1 U134 ( .x(N124), .a(IR_previous_5), .b(n5), .c(IR_curr_5), .d(n4), 
        .e(IR[5]), .f(n202) );
    ao222_1 U135 ( .x(N125), .a(IR_previous_6), .b(n5), .c(IR_curr_6), .d(n4), 
        .e(IR[6]), .f(n202) );
    ao222_1 U136 ( .x(N127), .a(IR_previous_8), .b(n5), .c(IR_curr_8), .d(n4), 
        .e(IR[8]), .f(n202) );
    ao222_1 U137 ( .x(N128), .a(IR_previous_9), .b(n5), .c(IR_curr_9), .d(n4), 
        .e(IR[9]), .f(n202) );
    ao222_1 U138 ( .x(N129), .a(IR_previous_10), .b(n5), .c(IR_curr_10), .d(n4
        ), .e(IR[10]), .f(n202) );
    ao222_1 U139 ( .x(N130), .a(IR_previous_11), .b(n5), .c(IR_curr_11), .d(n4
        ), .e(IR[11]), .f(n202) );
    ao222_1 U14 ( .x(N88), .a(PC[1]), .b(n5), .c(branch_address[1]), .d(n6), 
        .e(N18), .f(N215) );
    ao222_1 U140 ( .x(N131), .a(IR_previous_12), .b(n5), .c(IR_curr_12), .d(n4
        ), .e(IR[12]), .f(n202) );
    ao222_1 U141 ( .x(N132), .a(IR_previous_13), .b(n5), .c(IR_curr_13), .d(n4
        ), .e(IR[13]), .f(n202) );
    ao222_1 U142 ( .x(N133), .a(IR_previous_14), .b(n5), .c(IR_curr_14), .d(n4
        ), .e(IR[14]), .f(n202) );
    ao222_1 U143 ( .x(N134), .a(IR_previous_15), .b(n5), .c(IR_curr_15), .d(n4
        ), .e(IR[15]), .f(n202) );
    ao222_1 U144 ( .x(N135), .a(IR_previous_16), .b(n5), .c(IR_curr_16), .d(n4
        ), .e(IR[16]), .f(n202) );
    ao222_1 U145 ( .x(N136), .a(IR_previous_17), .b(n5), .c(IR_curr_17), .d(n4
        ), .e(IR[17]), .f(n202) );
    ao222_1 U146 ( .x(N137), .a(IR_previous_18), .b(n5), .c(IR_curr_18), .d(n4
        ), .e(IR[18]), .f(n202) );
    ao222_1 U147 ( .x(N139), .a(IR_previous_20), .b(n5), .c(IR_curr_20), .d(n4
        ), .e(IR[20]), .f(n202) );
    ao222_1 U148 ( .x(N140), .a(IR_previous_21), .b(n5), .c(IR_curr_21), .d(n4
        ), .e(IR[21]), .f(n202) );
    ao222_1 U149 ( .x(N141), .a(IR_previous_22), .b(n5), .c(IR_curr_22), .d(n4
        ), .e(IR[22]), .f(n202) );
    oai211_1 U15 ( .x(N108), .a(n201), .b(n44), .c(n45), .d(n46) );
    ao222_1 U150 ( .x(N142), .a(IR_previous_23), .b(n5), .c(IR_curr_23), .d(n4
        ), .e(IR[23]), .f(n202) );
    ao222_1 U151 ( .x(N143), .a(IR_previous_24), .b(n5), .c(IR_curr_24), .d(n4
        ), .e(IR[24]), .f(n202) );
    ao222_1 U152 ( .x(N144), .a(IR_previous_25), .b(n5), .c(IR_curr_25), .d(n4
        ), .e(IR[25]), .f(n202) );
    ao222_1 U153 ( .x(N146), .a(IR_previous_27), .b(n5), .c(IR_curr_27), .d(n4
        ), .e(IR[27]), .f(n202) );
    ao222_1 U154 ( .x(N147), .a(IR_previous_28), .b(n5), .c(IR_curr_28), .d(n4
        ), .e(IR[28]), .f(n202) );
    buf_3 U155 ( .x(n37), .a(n91) );
    oai21_2 U156 ( .x(n202), .a(N50), .b(n201), .c(n203) );
    ao222_1 U157 ( .x(N149), .a(IR_previous_30), .b(n5), .c(IR_curr_30), .d(n4
        ), .e(IR[30]), .f(n202) );
    nand2i_2 U158 ( .x(n61), .a(n97), .b(N152) );
    inv_2 U159 ( .x(n59), .a(N43) );
    inv_2 U16 ( .x(n44), .a(N38) );
    oai211_1 U160 ( .x(N113), .a(n201), .b(n59), .c(n60), .d(n61) );
    nand2i_2 U161 ( .x(n64), .a(n98), .b(N152) );
    nand2_2 U162 ( .x(n63), .a(branch_address[27]), .b(branch_sig) );
    inv_2 U163 ( .x(n62), .a(N44) );
    oai211_1 U164 ( .x(N114), .a(n201), .b(n62), .c(n63), .d(n64) );
    nand2i_2 U165 ( .x(n67), .a(n99), .b(N152) );
    nand2_2 U166 ( .x(n66), .a(branch_address[28]), .b(branch_sig) );
    inv_2 U167 ( .x(n65), .a(N45) );
    oai211_1 U168 ( .x(N115), .a(n201), .b(n65), .c(n66), .d(n67) );
    inv_2 U169 ( .x(n86), .a(n69) );
    nand2_2 U17 ( .x(n45), .a(branch_address[21]), .b(branch_sig) );
    nor2i_1 U170 ( .x(n70), .a(n68), .b(n86) );
    nand2i_2 U171 ( .x(n69), .a(n100), .b(N152) );
    nand2_2 U172 ( .x(n68), .a(branch_address[29]), .b(branch_sig) );
    inv_2 U173 ( .x(n85), .a(n78) );
    nor2i_1 U174 ( .x(n79), .a(n77), .b(n85) );
    nand2_2 U175 ( .x(n77), .a(branch_address[30]), .b(branch_sig) );
    inv_2 U176 ( .x(n89), .a(n201) );
    inv_2 U177 ( .x(n90), .a(n201) );
    inv_5 U178 ( .x(n76), .a(N48) );
    inv_2 U179 ( .x(n84), .a(n74) );
    nand2i_2 U18 ( .x(n46), .a(n92), .b(N152) );
    nor2i_1 U180 ( .x(n75), .a(n73), .b(n84) );
    nand2_2 U181 ( .x(n73), .a(branch_address[31]), .b(branch_sig) );
    aoi23_1 U182 ( .x(N118), .a(n75), .b(n76), .c(n73), .d(n201), .e(n74) );
    buf_14 U183 ( .x(NPC[4]), .a(n208) );
    inv_2 U184 ( .x(n82), .a(stall) );
    and2_3 U185 ( .x(n4), .a(N50), .b(N215) );
    buf_3 U186 ( .x(n40), .a(n91) );
    buf_3 U187 ( .x(n38), .a(n91) );
    inv_5 U188 ( .x(N152), .a(n88) );
    inv_2 U189 ( .x(n5), .a(n88) );
    ao222_1 U19 ( .x(N138), .a(IR_previous_19), .b(N152), .c(IR_curr_19), .d(
        n4), .e(IR[19]), .f(n202) );
    nand2i_2 U190 ( .x(n88), .a(branch_sig), .b(n72) );
    ao222_1 U191 ( .x(N104), .a(PC[17]), .b(N152), .c(branch_address[17]), .d(
        n6), .e(N34), .f(N215) );
    ao222_1 U192 ( .x(N98), .a(PC[11]), .b(N152), .c(branch_address[11]), .d(
        branch_sig), .e(N28), .f(N215) );
    inv_2 U193 ( .x(n6), .a(n203) );
    inv_2 U194 ( .x(n203), .a(branch_sig) );
    inv_2 U195 ( .x(n8), .a(n72) );
    inv_2 U196 ( .x(n7), .a(n72) );
    inv_2 U197 ( .x(n87), .a(n72) );
    nand3_1 U198 ( .x(n72), .a(n81), .b(n82), .c(n83) );
    buf_14 U199 ( .x(NPC[15]), .a(n204) );
    oai211_1 U20 ( .x(N112), .a(n201), .b(n56), .c(n57), .d(n58) );
    ao222_1 U201 ( .x(N92), .a(PC[5]), .b(N152), .c(branch_address[5]), .d(
        branch_sig), .e(N22), .f(N215) );
    ao222_1 U202 ( .x(N101), .a(PC[14]), .b(N152), .c(branch_address[14]), .d(
        branch_sig), .e(N31), .f(N215) );
    inv_2 U203 ( .x(n11), .a(n10) );
    buf_10 U204 ( .x(NPC[11]), .a(n205) );
    inv_2 U205 ( .x(n13), .a(n12) );
    inv_2 U206 ( .x(n15), .a(n14) );
    mux2_1 U207 ( .x(n184), .d0(PC[16]), .sl(n90), .d1(NPC[16]) );
    ao222_1 U208 ( .x(N87), .a(PC[0]), .b(N152), .c(branch_address[0]), .d(
        branch_sig), .e(N17), .f(N215) );
    ao222_1 U209 ( .x(N91), .a(PC[4]), .b(N152), .c(branch_address[4]), .d(
        branch_sig), .e(N21), .f(N215) );
    inv_2 U21 ( .x(n56), .a(N42) );
    ao222_1 U210 ( .x(N97), .a(PC[10]), .b(N152), .c(branch_address[10]), .d(
        branch_sig), .e(N27), .f(N215) );
    ao222_1 U211 ( .x(N93), .a(PC[6]), .b(N152), .c(branch_address[6]), .d(
        branch_sig), .e(N23), .f(N215) );
    nand2_2 U212 ( .x(n60), .a(branch_address[26]), .b(branch_sig) );
    inv_2 U214 ( .x(n17), .a(n16) );
    mux2_1 U215 ( .x(n183), .d0(PC[15]), .sl(n89), .d1(NPC[15]) );
    mux2_1 U216 ( .x(n185), .d0(PC[17]), .sl(n90), .d1(n11) );
    mux2_1 U217 ( .x(n176), .d0(PC[8]), .sl(n89), .d1(n17) );
    inv_2 U218 ( .x(n23), .a(n22) );
    mux2_1 U219 ( .x(n174), .d0(PC[6]), .sl(n89), .d1(n211) );
    nand2_2 U22 ( .x(n57), .a(branch_address[25]), .b(branch_sig) );
    inv_2 U220 ( .x(n25), .a(n24) );
    inv_2 U221 ( .x(n27), .a(n26) );
    mux2_1 U222 ( .x(n181), .d0(PC[13]), .sl(n90), .d1(n15) );
    mux2_1 U223 ( .x(n172), .d0(PC[4]), .sl(n90), .d1(NPC[4]) );
    mux2_1 U224 ( .x(n182), .d0(PC[14]), .sl(n89), .d1(n13) );
    ao222_1 U225 ( .x(N90), .a(PC[3]), .b(N152), .c(branch_address[3]), .d(
        branch_sig), .e(N20), .f(N215) );
    mux2_1 U226 ( .x(n178), .d0(PC[10]), .sl(n89), .d1(n25) );
    inv_2 U227 ( .x(n29), .a(n28) );
    inv_2 U228 ( .x(n31), .a(n30) );
    inv_2 U229 ( .x(n33), .a(n32) );
    nand2i_2 U23 ( .x(n58), .a(n96), .b(N152) );
    mux2_1 U230 ( .x(n179), .d0(PC[11]), .sl(n90), .d1(NPC[11]) );
    mux2_1 U231 ( .x(n177), .d0(PC[9]), .sl(n89), .d1(n23) );
    mux2_1 U232 ( .x(n175), .d0(PC[7]), .sl(n90), .d1(n27) );
    mux2_1 U233 ( .x(n180), .d0(PC[12]), .sl(n89), .d1(n29) );
    buf_16 U234 ( .x(NPC[3]), .a(n209) );
    buf_16 U235 ( .x(NPC[2]), .a(n210) );
    mux2_1 U236 ( .x(n173), .d0(PC[5]), .sl(n90), .d1(n212) );
    inv_6 U237 ( .x(n71), .a(N46) );
    inv_6 U238 ( .x(n80), .a(N47) );
    nand2i_4 U239 ( .x(n74), .a(n102), .b(N152) );
    ao222_1 U24 ( .x(N126), .a(IR_previous_7), .b(N152), .c(IR_curr_7), .d(n4), 
        .e(IR[7]), .f(n202) );
    nand2i_4 U240 ( .x(n78), .a(n101), .b(N152) );
    nand2i_6 U241 ( .x(n201), .a(branch_sig), .b(n7) );
    aoi23_4 U242 ( .x(N116), .a(n70), .b(n71), .c(n68), .d(n201), .e(n69) );
    aoi23_4 U243 ( .x(N117), .a(n79), .b(n80), .c(n77), .d(n201), .e(n78) );
    mux2_4 U244 ( .x(n167), .d0(IR_curr_31), .sl(n87), .d1(IR[31]) );
    inv_2 U245 ( .x(n91), .a(reset) );
    ao222_5 U247 ( .x(N99), .a(N152), .b(PC[12]), .c(branch_sig), .d(
        branch_address[12]), .e(N29), .f(N215) );
    inv_2 U248 ( .x(n211), .a(n258) );
    buf_10 U249 ( .x(NPC[6]), .a(n206) );
    ao222_2 U25 ( .x(N107), .a(PC[20]), .b(n5), .c(branch_address[20]), .d(n6), 
        .e(N37), .f(N215) );
    inv_2 U250 ( .x(n212), .a(n259) );
    buf_10 U251 ( .x(NPC[5]), .a(n207) );
    inv_0 U252 ( .x(n213), .a(NPC[21]) );
    inv_2 U253 ( .x(n214), .a(n213) );
    inv_5 U254 ( .x(n215), .a(n360) );
    inv_10 U255 ( .x(NPC[14]), .a(n215) );
    ao222_1 U256 ( .x(N103), .a(PC[16]), .b(n5), .c(branch_address[16]), .d(
        branch_sig), .e(N33), .f(N215) );
    inv_0 U257 ( .x(n217), .a(NPC[0]) );
    inv_2 U258 ( .x(n218), .a(n217) );
    ao222_1 U259 ( .x(N100), .a(PC[13]), .b(N152), .c(branch_address[13]), .d(
        branch_sig), .e(N30), .f(N215) );
    oai211_1 U26 ( .x(N110), .a(n201), .b(n50), .c(n51), .d(n52) );
    ao222_1 U260 ( .x(N106), .a(PC[19]), .b(N152), .c(branch_address[19]), .d(
        branch_sig), .e(N36), .f(N215) );
    inv_5 U27 ( .x(n50), .a(N40) );
    nand2_2 U28 ( .x(n51), .a(branch_address[23]), .b(branch_sig) );
    nand2i_2 U29 ( .x(n52), .a(n94), .b(N152) );
    oai211_1 U3 ( .x(N111), .a(n201), .b(n53), .c(n54), .d(n55) );
    inv_2 U30 ( .x(N215), .a(n201) );
    ao222_1 U31 ( .x(N105), .a(PC[18]), .b(N152), .c(branch_address[18]), .d(
        branch_sig), .e(N35), .f(N215) );
    ao222_1 U32 ( .x(N145), .a(IR_previous_26), .b(N152), .c(IR_curr_26), .d(
        n4), .e(IR[26]), .f(n202) );
    ao222_1 U33 ( .x(N102), .a(PC[15]), .b(n5), .c(branch_address[15]), .d(
        branch_sig), .e(N32), .f(N215) );
    ao222_4 U36 ( .x(N94), .a(PC[7]), .b(N152), .c(branch_address[7]), .d(
        branch_sig), .e(N24), .f(N215) );
    ao222_4 U37 ( .x(N96), .a(PC[9]), .b(n5), .c(branch_address[9]), .d(
        branch_sig), .e(N26), .f(N215) );
    ao222_1 U38 ( .x(N95), .a(PC[8]), .b(N152), .c(branch_address[8]), .d(
        branch_sig), .e(N25), .f(N215) );
    buf_3 U39 ( .x(n36), .a(n91) );
    ao222_1 U40 ( .x(N89), .a(PC[2]), .b(N152), .c(branch_address[2]), .d(
        branch_sig), .e(N19), .f(N215) );
    mux2_2 U41 ( .x(n104), .d0(IR_previous_0), .sl(n8), .d1(IR_latched[0]) );
    mux2_2 U42 ( .x(n105), .d0(IR_previous_1), .sl(n8), .d1(IR_latched[1]) );
    mux2_2 U43 ( .x(n106), .d0(IR_previous_2), .sl(n8), .d1(IR_latched[2]) );
    mux2_2 U44 ( .x(n107), .d0(IR_previous_3), .sl(n87), .d1(IR_latched[3]) );
    mux2_2 U45 ( .x(n108), .d0(IR_previous_4), .sl(n8), .d1(IR_latched[4]) );
    mux2_2 U46 ( .x(n109), .d0(IR_previous_5), .sl(n87), .d1(IR_latched[5]) );
    mux2_2 U47 ( .x(n110), .d0(IR_previous_6), .sl(n8), .d1(IR_latched[6]) );
    mux2_2 U48 ( .x(n111), .d0(IR_previous_7), .sl(n87), .d1(IR_latched[7]) );
    mux2_2 U49 ( .x(n112), .d0(IR_previous_8), .sl(n87), .d1(IR_latched[8]) );
    inv_2 U5 ( .x(n53), .a(N41) );
    mux2_2 U50 ( .x(n113), .d0(IR_previous_9), .sl(n87), .d1(IR_latched[9]) );
    mux2_2 U51 ( .x(n114), .d0(IR_previous_10), .sl(n8), .d1(IR_latched[10])
         );
    mux2_2 U52 ( .x(n115), .d0(IR_previous_11), .sl(n8), .d1(IR_latched[11])
         );
    mux2_2 U53 ( .x(n116), .d0(IR_previous_12), .sl(n8), .d1(IR_latched[12])
         );
    mux2_2 U54 ( .x(n117), .d0(IR_previous_13), .sl(n8), .d1(IR_latched[13])
         );
    mux2_2 U55 ( .x(n118), .d0(IR_previous_14), .sl(n8), .d1(IR_latched[14])
         );
    mux2_2 U56 ( .x(n119), .d0(IR_previous_15), .sl(n87), .d1(IR_latched[15])
         );
    mux2_2 U57 ( .x(n120), .d0(IR_previous_16), .sl(n8), .d1(IR_latched[16])
         );
    mux2_2 U58 ( .x(n121), .d0(IR_previous_17), .sl(n87), .d1(IR_latched[17])
         );
    mux2_2 U59 ( .x(n122), .d0(IR_previous_18), .sl(n8), .d1(IR_latched[18])
         );
    nand2_2 U6 ( .x(n54), .a(branch_address[24]), .b(branch_sig) );
    mux2_2 U60 ( .x(n123), .d0(IR_previous_19), .sl(n87), .d1(IR_latched[19])
         );
    mux2_2 U61 ( .x(n124), .d0(IR_previous_20), .sl(n87), .d1(IR_latched[20])
         );
    mux2_2 U62 ( .x(n125), .d0(IR_previous_21), .sl(n8), .d1(IR_latched[21])
         );
    mux2_2 U63 ( .x(n126), .d0(IR_previous_22), .sl(n87), .d1(IR_latched[22])
         );
    mux2_2 U64 ( .x(n127), .d0(IR_previous_23), .sl(n8), .d1(IR_latched[23])
         );
    mux2_2 U65 ( .x(n128), .d0(IR_previous_24), .sl(n87), .d1(IR_latched[24])
         );
    mux2_2 U66 ( .x(n129), .d0(IR_previous_25), .sl(n8), .d1(IR_latched[25])
         );
    mux2_2 U67 ( .x(n130), .d0(IR_previous_26), .sl(n87), .d1(IR_latched[26])
         );
    mux2_2 U68 ( .x(n131), .d0(IR_previous_27), .sl(n8), .d1(IR_latched[27])
         );
    mux2_2 U69 ( .x(n132), .d0(IR_previous_28), .sl(n87), .d1(IR_latched[28])
         );
    nand2i_2 U7 ( .x(n55), .a(n95), .b(N152) );
    mux2_2 U70 ( .x(n133), .d0(IR_previous_29), .sl(n8), .d1(IR_latched[29])
         );
    mux2_2 U71 ( .x(n134), .d0(IR_previous_30), .sl(n8), .d1(IR_latched[30])
         );
    mux2_2 U72 ( .x(n135), .d0(IR_previous_31), .sl(n87), .d1(IR_latched[31])
         );
    mux2_2 U73 ( .x(n136), .d0(IR_curr_0), .sl(n8), .d1(IR[0]) );
    mux2_2 U74 ( .x(n137), .d0(IR_curr_1), .sl(n8), .d1(IR[1]) );
    mux2_2 U75 ( .x(n138), .d0(IR_curr_2), .sl(n87), .d1(IR[2]) );
    mux2_2 U76 ( .x(n139), .d0(IR_curr_3), .sl(n87), .d1(IR[3]) );
    mux2_2 U77 ( .x(n140), .d0(IR_curr_4), .sl(n87), .d1(IR[4]) );
    mux2_2 U78 ( .x(n141), .d0(IR_curr_5), .sl(n87), .d1(IR[5]) );
    mux2_2 U79 ( .x(n142), .d0(IR_curr_6), .sl(n87), .d1(IR[6]) );
    oai211_1 U8 ( .x(N109), .a(n201), .b(n47), .c(n48), .d(n49) );
    mux2_2 U80 ( .x(n143), .d0(IR_curr_7), .sl(n87), .d1(IR[7]) );
    mux2_2 U81 ( .x(n144), .d0(IR_curr_8), .sl(n87), .d1(IR[8]) );
    mux2_2 U82 ( .x(n145), .d0(IR_curr_9), .sl(n87), .d1(IR[9]) );
    mux2_2 U83 ( .x(n146), .d0(IR_curr_10), .sl(n8), .d1(IR[10]) );
    mux2_2 U84 ( .x(n147), .d0(IR_curr_11), .sl(n8), .d1(IR[11]) );
    mux2_2 U85 ( .x(n148), .d0(IR_curr_12), .sl(n8), .d1(IR[12]) );
    mux2_2 U86 ( .x(n149), .d0(IR_curr_13), .sl(n8), .d1(IR[13]) );
    mux2_2 U87 ( .x(n150), .d0(IR_curr_14), .sl(n8), .d1(IR[14]) );
    mux2_2 U88 ( .x(n151), .d0(IR_curr_15), .sl(n8), .d1(IR[15]) );
    mux2_2 U89 ( .x(n152), .d0(IR_curr_16), .sl(n8), .d1(IR[16]) );
    inv_2 U9 ( .x(n47), .a(N39) );
    mux2_2 U90 ( .x(n153), .d0(IR_curr_17), .sl(n8), .d1(IR[17]) );
    mux2_2 U91 ( .x(n154), .d0(IR_curr_18), .sl(n8), .d1(IR[18]) );
    mux2_2 U92 ( .x(n155), .d0(IR_curr_19), .sl(n87), .d1(IR[19]) );
    mux2_2 U93 ( .x(n156), .d0(IR_curr_20), .sl(n87), .d1(IR[20]) );
    mux2_2 U94 ( .x(n157), .d0(IR_curr_21), .sl(n87), .d1(IR[21]) );
    mux2_2 U95 ( .x(n158), .d0(IR_curr_22), .sl(n8), .d1(IR[22]) );
    mux2_2 U96 ( .x(n159), .d0(IR_curr_23), .sl(n8), .d1(IR[23]) );
    mux2_2 U97 ( .x(n160), .d0(IR_curr_24), .sl(n8), .d1(IR[24]) );
    mux2_2 U98 ( .x(n161), .d0(IR_curr_25), .sl(n87), .d1(IR[25]) );
    mux2_2 U99 ( .x(n162), .d0(IR_curr_26), .sl(n87), .d1(IR[26]) );
    IF_DW01_add_32_0_test_1 add_100 ( .A({NPC[31], NPC[30], NPC[29], NPC[28], 
        NPC[27], NPC[26], NPC[25], NPC[24], NPC[23], NPC[22], n214, NPC[20], 
        NPC[19], NPC[18], n11, NPC[16], NPC[15], n13, n15, n29, NPC[11], n25, 
        n23, n17, n27, n211, n212, NPC[4], n31, n33, NPC[1], n218}), .B({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0}), .CI(1'b0), .SUM({N48, N47, 
        N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, 
        N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, 
        N18, N17}) );
    smlatnr_1 stalled_reg__master ( .q(stalled_reg__m2s), .d(n200), .sdi(PC
        [31]), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 stalled_reg__slave ( .q(N50), .qb(test_so1), .d(stalled_reg__m2s), 
        .g(Ctrl__Regs_1__en2), .rb(n38), .glob_g(global_g2), .sync_sel(
        sync_sel) );
endmodule


module MEM_test_1_desync ( reg_write_MEM, mem_to_reg_EX, reset, ALU_result, 
    reg_write_EX, mem_to_reg_MEM, reg_out_B_EX, reg_out_B_MEM, DM_read_data, 
    RF_data_in, test_si, test_so, test_se, sync_sel, global_g1, global_g2, 
    Ctrl__Regs_1__en1, Ctrl__Regs_1__en2 );
input  [31:0] ALU_result;
input  [31:0] reg_out_B_EX;
output [31:0] reg_out_B_MEM;
input  [31:0] DM_read_data;
output [31:0] RF_data_in;
input  mem_to_reg_EX, reset, reg_write_EX, test_si, test_se, sync_sel, 
    global_g1, global_g2, Ctrl__Regs_1__en1, Ctrl__Regs_1__en2;
output reg_write_MEM, mem_to_reg_MEM, test_so;
    wire RF_data_in_reg_0__m2s, n15, n4, n16, RF_data_in_reg_10__m2s, n69, n18, 
        n6, n70, RF_data_in_reg_11__m2s, n43, n44, RF_data_in_reg_12__m2s, n67, 
        n5, n68, RF_data_in_reg_13__m2s, n65, n66, RF_data_in_reg_14__m2s, n11, 
        n12, RF_data_in_reg_15__m2s, n63, n64, RF_data_in_reg_16__m2s, n61, 
        n62, RF_data_in_reg_17__m2s, n59, n60, RF_data_in_reg_18__m2s, n57, 
        n58, RF_data_in_reg_19__m2s, n35, n36, RF_data_in_reg_1__m2s, n13, n14, 
        RF_data_in_reg_20__m2s, n55, n56, RF_data_in_reg_21__m2s, n53, n54, 
        RF_data_in_reg_22__m2s, n33, n34, RF_data_in_reg_23__m2s, n51, n52, 
        RF_data_in_reg_24__m2s, n49, n50, RF_data_in_reg_25__m2s, n47, n48, 
        RF_data_in_reg_26__m2s, n21, n22, RF_data_in_reg_27__m2s, n31, n32, 
        RF_data_in_reg_28__m2s, n45, n46, RF_data_in_reg_29__m2s, n29, n30, 
        RF_data_in_reg_2__m2s, n39, n40, RF_data_in_reg_30__m2s, n25, n26, 
        RF_data_in_reg_31__m2s, n23, n24, RF_data_in_reg_3__m2s, n41, n42, 
        RF_data_in_reg_4__m2s, n73, n74, RF_data_in_reg_5__m2s, n71, n72, 
        RF_data_in_reg_6__m2s, n37, n38, RF_data_in_reg_7__m2s, n19, n75, n20, 
        RF_data_in_reg_8__m2s, n27, n28, RF_data_in_reg_9__m2s, n17, n3, 
        mem_to_reg_MEM_reg__m2s, reg_out_B_MEM_reg_0__m2s, 
        reg_out_B_MEM_reg_10__m2s, reg_out_B_MEM_reg_11__m2s, 
        reg_out_B_MEM_reg_12__m2s, reg_out_B_MEM_reg_13__m2s, 
        reg_out_B_MEM_reg_14__m2s, reg_out_B_MEM_reg_15__m2s, 
        reg_out_B_MEM_reg_16__m2s, reg_out_B_MEM_reg_17__m2s, 
        reg_out_B_MEM_reg_18__m2s, reg_out_B_MEM_reg_19__m2s, 
        reg_out_B_MEM_reg_1__m2s, reg_out_B_MEM_reg_20__m2s, 
        reg_out_B_MEM_reg_21__m2s, reg_out_B_MEM_reg_22__m2s, 
        reg_out_B_MEM_reg_23__m2s, reg_out_B_MEM_reg_24__m2s, 
        reg_out_B_MEM_reg_25__m2s, reg_out_B_MEM_reg_26__m2s, 
        reg_out_B_MEM_reg_27__m2s, reg_out_B_MEM_reg_28__m2s, 
        reg_out_B_MEM_reg_29__m2s, reg_out_B_MEM_reg_2__m2s, 
        reg_out_B_MEM_reg_30__m2s, reg_out_B_MEM_reg_31__m2s, 
        reg_out_B_MEM_reg_3__m2s, reg_out_B_MEM_reg_4__m2s, 
        reg_out_B_MEM_reg_5__m2s, reg_out_B_MEM_reg_6__m2s, 
        reg_out_B_MEM_reg_7__m2s, reg_out_B_MEM_reg_8__m2s, 
        reg_out_B_MEM_reg_9__m2s, reg_write_MEM_reg__m2s;
    smlatnr_1 RF_data_in_reg_0__master ( .q(RF_data_in_reg_0__m2s), .d(n15), 
        .sdi(test_si), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 RF_data_in_reg_0__slave ( .q(RF_data_in[0]), .qb(n16), .d(
        RF_data_in_reg_0__m2s), .g(Ctrl__Regs_1__en2), .rb(n4), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 RF_data_in_reg_10__master ( .q(RF_data_in_reg_10__m2s), .d(n69), 
        .sdi(n18), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n6), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_1 RF_data_in_reg_10__slave ( .q(RF_data_in[10]), .qb(n70), .d(
        RF_data_in_reg_10__m2s), .g(Ctrl__Regs_1__en2), .rb(n6), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 RF_data_in_reg_11__master ( .q(RF_data_in_reg_11__m2s), .d(n43), 
        .sdi(n70), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_1 RF_data_in_reg_11__slave ( .q(RF_data_in[11]), .qb(n44), .d(
        RF_data_in_reg_11__m2s), .g(Ctrl__Regs_1__en2), .rb(n4), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 RF_data_in_reg_12__master ( .q(RF_data_in_reg_12__m2s), .d(n67), 
        .sdi(n44), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n5), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_1 RF_data_in_reg_12__slave ( .q(RF_data_in[12]), .qb(n68), .d(
        RF_data_in_reg_12__m2s), .g(Ctrl__Regs_1__en2), .rb(n5), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 RF_data_in_reg_13__master ( .q(RF_data_in_reg_13__m2s), .d(n65), 
        .sdi(n68), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n5), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_1 RF_data_in_reg_13__slave ( .q(RF_data_in[13]), .qb(n66), .d(
        RF_data_in_reg_13__m2s), .g(Ctrl__Regs_1__en2), .rb(n5), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 RF_data_in_reg_14__master ( .q(RF_data_in_reg_14__m2s), .d(n11), 
        .sdi(n66), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n5), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_1 RF_data_in_reg_14__slave ( .q(RF_data_in[14]), .qb(n12), .d(
        RF_data_in_reg_14__m2s), .g(Ctrl__Regs_1__en2), .rb(n5), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 RF_data_in_reg_15__master ( .q(RF_data_in_reg_15__m2s), .d(n63), 
        .sdi(n12), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n5), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_1 RF_data_in_reg_15__slave ( .q(RF_data_in[15]), .qb(n64), .d(
        RF_data_in_reg_15__m2s), .g(Ctrl__Regs_1__en2), .rb(n5), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 RF_data_in_reg_16__master ( .q(RF_data_in_reg_16__m2s), .d(n61), 
        .sdi(n64), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_1 RF_data_in_reg_16__slave ( .q(RF_data_in[16]), .qb(n62), .d(
        RF_data_in_reg_16__m2s), .g(Ctrl__Regs_1__en2), .rb(n4), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 RF_data_in_reg_17__master ( .q(RF_data_in_reg_17__m2s), .d(n59), 
        .sdi(n62), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n6), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_1 RF_data_in_reg_17__slave ( .q(RF_data_in[17]), .qb(n60), .d(
        RF_data_in_reg_17__m2s), .g(Ctrl__Regs_1__en2), .rb(n6), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 RF_data_in_reg_18__master ( .q(RF_data_in_reg_18__m2s), .d(n57), 
        .sdi(n60), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_1 RF_data_in_reg_18__slave ( .q(RF_data_in[18]), .qb(n58), .d(
        RF_data_in_reg_18__m2s), .g(Ctrl__Regs_1__en2), .rb(n4), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 RF_data_in_reg_19__master ( .q(RF_data_in_reg_19__m2s), .d(n35), 
        .sdi(n58), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n6), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_1 RF_data_in_reg_19__slave ( .q(RF_data_in[19]), .qb(n36), .d(
        RF_data_in_reg_19__m2s), .g(Ctrl__Regs_1__en2), .rb(n6), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 RF_data_in_reg_1__master ( .q(RF_data_in_reg_1__m2s), .d(n13), 
        .sdi(n16), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n5), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 RF_data_in_reg_1__slave ( .q(RF_data_in[1]), .qb(n14), .d(
        RF_data_in_reg_1__m2s), .g(Ctrl__Regs_1__en2), .rb(n5), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 RF_data_in_reg_20__master ( .q(RF_data_in_reg_20__m2s), .d(n55), 
        .sdi(n36), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n6), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_1 RF_data_in_reg_20__slave ( .q(RF_data_in[20]), .qb(n56), .d(
        RF_data_in_reg_20__m2s), .g(Ctrl__Regs_1__en2), .rb(n6), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 RF_data_in_reg_21__master ( .q(RF_data_in_reg_21__m2s), .d(n53), 
        .sdi(n56), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n6), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_1 RF_data_in_reg_21__slave ( .q(RF_data_in[21]), .qb(n54), .d(
        RF_data_in_reg_21__m2s), .g(Ctrl__Regs_1__en2), .rb(n6), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 RF_data_in_reg_22__master ( .q(RF_data_in_reg_22__m2s), .d(n33), 
        .sdi(n54), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_1 RF_data_in_reg_22__slave ( .q(RF_data_in[22]), .qb(n34), .d(
        RF_data_in_reg_22__m2s), .g(Ctrl__Regs_1__en2), .rb(n4), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 RF_data_in_reg_23__master ( .q(RF_data_in_reg_23__m2s), .d(n51), 
        .sdi(n34), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_1 RF_data_in_reg_23__slave ( .q(RF_data_in[23]), .qb(n52), .d(
        RF_data_in_reg_23__m2s), .g(Ctrl__Regs_1__en2), .rb(n4), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 RF_data_in_reg_24__master ( .q(RF_data_in_reg_24__m2s), .d(n49), 
        .sdi(n52), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n6), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_1 RF_data_in_reg_24__slave ( .q(RF_data_in[24]), .qb(n50), .d(
        RF_data_in_reg_24__m2s), .g(Ctrl__Regs_1__en2), .rb(n6), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 RF_data_in_reg_25__master ( .q(RF_data_in_reg_25__m2s), .d(n47), 
        .sdi(n50), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n5), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_1 RF_data_in_reg_25__slave ( .q(RF_data_in[25]), .qb(n48), .d(
        RF_data_in_reg_25__m2s), .g(Ctrl__Regs_1__en2), .rb(n5), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 RF_data_in_reg_26__master ( .q(RF_data_in_reg_26__m2s), .d(n21), 
        .sdi(n48), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n5), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_1 RF_data_in_reg_26__slave ( .q(RF_data_in[26]), .qb(n22), .d(
        RF_data_in_reg_26__m2s), .g(Ctrl__Regs_1__en2), .rb(n5), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 RF_data_in_reg_27__master ( .q(RF_data_in_reg_27__m2s), .d(n31), 
        .sdi(n22), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n5), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_1 RF_data_in_reg_27__slave ( .q(RF_data_in[27]), .qb(n32), .d(
        RF_data_in_reg_27__m2s), .g(Ctrl__Regs_1__en2), .rb(n5), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 RF_data_in_reg_28__master ( .q(RF_data_in_reg_28__m2s), .d(n45), 
        .sdi(n32), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_1 RF_data_in_reg_28__slave ( .q(RF_data_in[28]), .qb(n46), .d(
        RF_data_in_reg_28__m2s), .g(Ctrl__Regs_1__en2), .rb(n4), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 RF_data_in_reg_29__master ( .q(RF_data_in_reg_29__m2s), .d(n29), 
        .sdi(n46), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n5), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_1 RF_data_in_reg_29__slave ( .q(RF_data_in[29]), .qb(n30), .d(
        RF_data_in_reg_29__m2s), .g(Ctrl__Regs_1__en2), .rb(n5), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 RF_data_in_reg_2__master ( .q(RF_data_in_reg_2__m2s), .d(n39), 
        .sdi(n14), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n6), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 RF_data_in_reg_2__slave ( .q(RF_data_in[2]), .qb(n40), .d(
        RF_data_in_reg_2__m2s), .g(Ctrl__Regs_1__en2), .rb(n6), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 RF_data_in_reg_30__master ( .q(RF_data_in_reg_30__m2s), .d(n25), 
        .sdi(n30), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_1 RF_data_in_reg_30__slave ( .q(RF_data_in[30]), .qb(n26), .d(
        RF_data_in_reg_30__m2s), .g(Ctrl__Regs_1__en2), .rb(n4), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 RF_data_in_reg_31__master ( .q(RF_data_in_reg_31__m2s), .d(n23), 
        .sdi(n26), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n6), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_1 RF_data_in_reg_31__slave ( .q(RF_data_in[31]), .qb(n24), .d(
        RF_data_in_reg_31__m2s), .g(Ctrl__Regs_1__en2), .rb(n6), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 RF_data_in_reg_3__master ( .q(RF_data_in_reg_3__m2s), .d(n41), 
        .sdi(n40), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 RF_data_in_reg_3__slave ( .q(RF_data_in[3]), .qb(n42), .d(
        RF_data_in_reg_3__m2s), .g(Ctrl__Regs_1__en2), .rb(n4), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 RF_data_in_reg_4__master ( .q(RF_data_in_reg_4__m2s), .d(n73), 
        .sdi(n42), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n5), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 RF_data_in_reg_4__slave ( .q(RF_data_in[4]), .qb(n74), .d(
        RF_data_in_reg_4__m2s), .g(Ctrl__Regs_1__en2), .rb(n5), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 RF_data_in_reg_5__master ( .q(RF_data_in_reg_5__m2s), .d(n71), 
        .sdi(n74), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n6), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 RF_data_in_reg_5__slave ( .q(RF_data_in[5]), .qb(n72), .d(
        RF_data_in_reg_5__m2s), .g(Ctrl__Regs_1__en2), .rb(n6), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 RF_data_in_reg_6__master ( .q(RF_data_in_reg_6__m2s), .d(n37), 
        .sdi(n72), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_4 RF_data_in_reg_6__slave ( .q(RF_data_in[6]), .qb(n38), .d(
        RF_data_in_reg_6__m2s), .g(Ctrl__Regs_1__en2), .rb(n4), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 RF_data_in_reg_7__master ( .q(RF_data_in_reg_7__m2s), .d(n19), 
        .sdi(n38), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n6), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_4 RF_data_in_reg_7__slave ( .q(n75), .qb(n20), .d(
        RF_data_in_reg_7__m2s), .g(Ctrl__Regs_1__en2), .rb(n6), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 RF_data_in_reg_8__master ( .q(RF_data_in_reg_8__m2s), .d(n27), 
        .sdi(n20), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n6), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_1 RF_data_in_reg_8__slave ( .q(RF_data_in[8]), .qb(n28), .d(
        RF_data_in_reg_8__m2s), .g(Ctrl__Regs_1__en2), .rb(n6), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 RF_data_in_reg_9__master ( .q(RF_data_in_reg_9__m2s), .d(n17), 
        .sdi(n28), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n5), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_1 RF_data_in_reg_9__slave ( .q(RF_data_in[9]), .qb(n18), .d(
        RF_data_in_reg_9__m2s), .g(Ctrl__Regs_1__en2), .rb(n5), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    mux2_1 U10 ( .x(n23), .d0(ALU_result[31]), .sl(mem_to_reg_EX), .d1(
        DM_read_data[31]) );
    mux2_1 U11 ( .x(n25), .d0(ALU_result[30]), .sl(mem_to_reg_EX), .d1(
        DM_read_data[30]) );
    mux2_1 U12 ( .x(n27), .d0(ALU_result[8]), .sl(mem_to_reg_EX), .d1(
        DM_read_data[8]) );
    mux2_1 U13 ( .x(n29), .d0(ALU_result[29]), .sl(mem_to_reg_EX), .d1(
        DM_read_data[29]) );
    mux2_1 U14 ( .x(n31), .d0(ALU_result[27]), .sl(mem_to_reg_EX), .d1(
        DM_read_data[27]) );
    mux2_1 U15 ( .x(n33), .d0(ALU_result[22]), .sl(mem_to_reg_EX), .d1(
        DM_read_data[22]) );
    mux2_1 U16 ( .x(n35), .d0(ALU_result[19]), .sl(mem_to_reg_EX), .d1(
        DM_read_data[19]) );
    mux2_1 U17 ( .x(n37), .d0(ALU_result[6]), .sl(mem_to_reg_EX), .d1(
        DM_read_data[6]) );
    mux2_1 U18 ( .x(n39), .d0(ALU_result[2]), .sl(mem_to_reg_EX), .d1(
        DM_read_data[2]) );
    mux2_1 U19 ( .x(n41), .d0(ALU_result[3]), .sl(mem_to_reg_EX), .d1(
        DM_read_data[3]) );
    mux2_1 U20 ( .x(n43), .d0(ALU_result[11]), .sl(mem_to_reg_EX), .d1(
        DM_read_data[11]) );
    mux2_1 U21 ( .x(n45), .d0(ALU_result[28]), .sl(mem_to_reg_EX), .d1(
        DM_read_data[28]) );
    mux2_1 U22 ( .x(n47), .d0(ALU_result[25]), .sl(mem_to_reg_EX), .d1(
        DM_read_data[25]) );
    mux2_1 U23 ( .x(n49), .d0(ALU_result[24]), .sl(mem_to_reg_EX), .d1(
        DM_read_data[24]) );
    mux2_1 U24 ( .x(n51), .d0(ALU_result[23]), .sl(mem_to_reg_EX), .d1(
        DM_read_data[23]) );
    mux2_1 U25 ( .x(n53), .d0(ALU_result[21]), .sl(mem_to_reg_EX), .d1(
        DM_read_data[21]) );
    mux2_1 U26 ( .x(n55), .d0(ALU_result[20]), .sl(mem_to_reg_EX), .d1(
        DM_read_data[20]) );
    mux2_1 U27 ( .x(n57), .d0(ALU_result[18]), .sl(mem_to_reg_EX), .d1(
        DM_read_data[18]) );
    mux2_1 U28 ( .x(n59), .d0(ALU_result[17]), .sl(mem_to_reg_EX), .d1(
        DM_read_data[17]) );
    mux2_1 U29 ( .x(n61), .d0(ALU_result[16]), .sl(mem_to_reg_EX), .d1(
        DM_read_data[16]) );
    buf_3 U3 ( .x(n3), .a(mem_to_reg_EX) );
    mux2_1 U30 ( .x(n63), .d0(ALU_result[15]), .sl(mem_to_reg_EX), .d1(
        DM_read_data[15]) );
    mux2_1 U31 ( .x(n65), .d0(ALU_result[13]), .sl(mem_to_reg_EX), .d1(
        DM_read_data[13]) );
    mux2_1 U32 ( .x(n67), .d0(ALU_result[12]), .sl(mem_to_reg_EX), .d1(
        DM_read_data[12]) );
    mux2_1 U33 ( .x(n69), .d0(ALU_result[10]), .sl(mem_to_reg_EX), .d1(
        DM_read_data[10]) );
    mux2_1 U34 ( .x(n71), .d0(ALU_result[5]), .sl(mem_to_reg_EX), .d1(
        DM_read_data[5]) );
    mux2_1 U35 ( .x(n73), .d0(ALU_result[4]), .sl(n3), .d1(DM_read_data[4]) );
    inv_2 U4 ( .x(n5), .a(reset) );
    inv_2 U5 ( .x(n4), .a(reset) );
    inv_2 U6 ( .x(n6), .a(reset) );
    buf_16 U7 ( .x(RF_data_in[7]), .a(n75) );
    mux2_1 U8 ( .x(n19), .d0(ALU_result[7]), .sl(mem_to_reg_EX), .d1(
        DM_read_data[7]) );
    mux2_1 U9 ( .x(n21), .d0(ALU_result[26]), .sl(mem_to_reg_EX), .d1(
        DM_read_data[26]) );
    mux2_1 _RF_data_in_reg_0_U4 ( .x(n15), .d0(ALU_result[0]), .sl(
        mem_to_reg_EX), .d1(DM_read_data[0]) );
    mux2_1 _RF_data_in_reg_14_U4 ( .x(n11), .d0(ALU_result[14]), .sl(
        mem_to_reg_EX), .d1(DM_read_data[14]) );
    mux2_1 _RF_data_in_reg_1_U4 ( .x(n13), .d0(ALU_result[1]), .sl(
        mem_to_reg_EX), .d1(DM_read_data[1]) );
    mux2_1 _RF_data_in_reg_9_U4 ( .x(n17), .d0(ALU_result[9]), .sl(
        mem_to_reg_EX), .d1(DM_read_data[9]) );
    smlatnr_1 mem_to_reg_MEM_reg__master ( .q(mem_to_reg_MEM_reg__m2s), .d(n3), 
        .sdi(n24), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n5), .glob_g(
        global_g1), .sync_sel(sync_sel) );
    mlatnr_2 mem_to_reg_MEM_reg__slave ( .q(mem_to_reg_MEM), .d(
        mem_to_reg_MEM_reg__m2s), .g(Ctrl__Regs_1__en2), .rb(n5), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_MEM_reg_0__master ( .q(reg_out_B_MEM_reg_0__m2s), .d(
        reg_out_B_EX[0]), .sdi(mem_to_reg_MEM), .se(test_se), .g(
        Ctrl__Regs_1__en1), .rb(n4), .glob_g(global_g1), .sync_sel(sync_sel)
         );
    mlatnr_2 reg_out_B_MEM_reg_0__slave ( .q(reg_out_B_MEM[0]), .d(
        reg_out_B_MEM_reg_0__m2s), .g(Ctrl__Regs_1__en2), .rb(n4), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_MEM_reg_10__master ( .q(reg_out_B_MEM_reg_10__m2s), 
        .d(reg_out_B_EX[10]), .sdi(reg_out_B_MEM[9]), .se(test_se), .g(
        Ctrl__Regs_1__en1), .rb(n5), .glob_g(global_g1), .sync_sel(sync_sel)
         );
    mlatnr_2 reg_out_B_MEM_reg_10__slave ( .q(reg_out_B_MEM[10]), .d(
        reg_out_B_MEM_reg_10__m2s), .g(Ctrl__Regs_1__en2), .rb(n5), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_MEM_reg_11__master ( .q(reg_out_B_MEM_reg_11__m2s), 
        .d(reg_out_B_EX[11]), .sdi(reg_out_B_MEM[10]), .se(test_se), .g(
        Ctrl__Regs_1__en1), .rb(n5), .glob_g(global_g1), .sync_sel(sync_sel)
         );
    mlatnr_2 reg_out_B_MEM_reg_11__slave ( .q(reg_out_B_MEM[11]), .d(
        reg_out_B_MEM_reg_11__m2s), .g(Ctrl__Regs_1__en2), .rb(n5), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_MEM_reg_12__master ( .q(reg_out_B_MEM_reg_12__m2s), 
        .d(reg_out_B_EX[12]), .sdi(reg_out_B_MEM[11]), .se(test_se), .g(
        Ctrl__Regs_1__en1), .rb(n4), .glob_g(global_g1), .sync_sel(sync_sel)
         );
    mlatnr_2 reg_out_B_MEM_reg_12__slave ( .q(reg_out_B_MEM[12]), .d(
        reg_out_B_MEM_reg_12__m2s), .g(Ctrl__Regs_1__en2), .rb(n4), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_MEM_reg_13__master ( .q(reg_out_B_MEM_reg_13__m2s), 
        .d(reg_out_B_EX[13]), .sdi(reg_out_B_MEM[12]), .se(test_se), .g(
        Ctrl__Regs_1__en1), .rb(n6), .glob_g(global_g1), .sync_sel(sync_sel)
         );
    mlatnr_2 reg_out_B_MEM_reg_13__slave ( .q(reg_out_B_MEM[13]), .d(
        reg_out_B_MEM_reg_13__m2s), .g(Ctrl__Regs_1__en2), .rb(n6), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_MEM_reg_14__master ( .q(reg_out_B_MEM_reg_14__m2s), 
        .d(reg_out_B_EX[14]), .sdi(reg_out_B_MEM[13]), .se(test_se), .g(
        Ctrl__Regs_1__en1), .rb(n6), .glob_g(global_g1), .sync_sel(sync_sel)
         );
    mlatnr_2 reg_out_B_MEM_reg_14__slave ( .q(reg_out_B_MEM[14]), .d(
        reg_out_B_MEM_reg_14__m2s), .g(Ctrl__Regs_1__en2), .rb(n6), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_MEM_reg_15__master ( .q(reg_out_B_MEM_reg_15__m2s), 
        .d(reg_out_B_EX[15]), .sdi(reg_out_B_MEM[14]), .se(test_se), .g(
        Ctrl__Regs_1__en1), .rb(n4), .glob_g(global_g1), .sync_sel(sync_sel)
         );
    mlatnr_2 reg_out_B_MEM_reg_15__slave ( .q(reg_out_B_MEM[15]), .d(
        reg_out_B_MEM_reg_15__m2s), .g(Ctrl__Regs_1__en2), .rb(n4), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_MEM_reg_16__master ( .q(reg_out_B_MEM_reg_16__m2s), 
        .d(reg_out_B_EX[16]), .sdi(reg_out_B_MEM[15]), .se(test_se), .g(
        Ctrl__Regs_1__en1), .rb(n5), .glob_g(global_g1), .sync_sel(sync_sel)
         );
    mlatnr_2 reg_out_B_MEM_reg_16__slave ( .q(reg_out_B_MEM[16]), .d(
        reg_out_B_MEM_reg_16__m2s), .g(Ctrl__Regs_1__en2), .rb(n5), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_MEM_reg_17__master ( .q(reg_out_B_MEM_reg_17__m2s), 
        .d(reg_out_B_EX[17]), .sdi(reg_out_B_MEM[16]), .se(test_se), .g(
        Ctrl__Regs_1__en1), .rb(n6), .glob_g(global_g1), .sync_sel(sync_sel)
         );
    mlatnr_2 reg_out_B_MEM_reg_17__slave ( .q(reg_out_B_MEM[17]), .d(
        reg_out_B_MEM_reg_17__m2s), .g(Ctrl__Regs_1__en2), .rb(n6), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_MEM_reg_18__master ( .q(reg_out_B_MEM_reg_18__m2s), 
        .d(reg_out_B_EX[18]), .sdi(reg_out_B_MEM[17]), .se(test_se), .g(
        Ctrl__Regs_1__en1), .rb(n4), .glob_g(global_g1), .sync_sel(sync_sel)
         );
    mlatnr_2 reg_out_B_MEM_reg_18__slave ( .q(reg_out_B_MEM[18]), .d(
        reg_out_B_MEM_reg_18__m2s), .g(Ctrl__Regs_1__en2), .rb(n4), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_MEM_reg_19__master ( .q(reg_out_B_MEM_reg_19__m2s), 
        .d(reg_out_B_EX[19]), .sdi(reg_out_B_MEM[18]), .se(test_se), .g(
        Ctrl__Regs_1__en1), .rb(n5), .glob_g(global_g1), .sync_sel(sync_sel)
         );
    mlatnr_2 reg_out_B_MEM_reg_19__slave ( .q(reg_out_B_MEM[19]), .d(
        reg_out_B_MEM_reg_19__m2s), .g(Ctrl__Regs_1__en2), .rb(n5), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_MEM_reg_1__master ( .q(reg_out_B_MEM_reg_1__m2s), .d(
        reg_out_B_EX[1]), .sdi(reg_out_B_MEM[0]), .se(test_se), .g(
        Ctrl__Regs_1__en1), .rb(n4), .glob_g(global_g1), .sync_sel(sync_sel)
         );
    mlatnr_2 reg_out_B_MEM_reg_1__slave ( .q(reg_out_B_MEM[1]), .d(
        reg_out_B_MEM_reg_1__m2s), .g(Ctrl__Regs_1__en2), .rb(n4), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_MEM_reg_20__master ( .q(reg_out_B_MEM_reg_20__m2s), 
        .d(reg_out_B_EX[20]), .sdi(reg_out_B_MEM[19]), .se(test_se), .g(
        Ctrl__Regs_1__en1), .rb(n6), .glob_g(global_g1), .sync_sel(sync_sel)
         );
    mlatnr_2 reg_out_B_MEM_reg_20__slave ( .q(reg_out_B_MEM[20]), .d(
        reg_out_B_MEM_reg_20__m2s), .g(Ctrl__Regs_1__en2), .rb(n6), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_MEM_reg_21__master ( .q(reg_out_B_MEM_reg_21__m2s), 
        .d(reg_out_B_EX[21]), .sdi(reg_out_B_MEM[20]), .se(test_se), .g(
        Ctrl__Regs_1__en1), .rb(n4), .glob_g(global_g1), .sync_sel(sync_sel)
         );
    mlatnr_2 reg_out_B_MEM_reg_21__slave ( .q(reg_out_B_MEM[21]), .d(
        reg_out_B_MEM_reg_21__m2s), .g(Ctrl__Regs_1__en2), .rb(n4), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_MEM_reg_22__master ( .q(reg_out_B_MEM_reg_22__m2s), 
        .d(reg_out_B_EX[22]), .sdi(reg_out_B_MEM[21]), .se(test_se), .g(
        Ctrl__Regs_1__en1), .rb(n5), .glob_g(global_g1), .sync_sel(sync_sel)
         );
    mlatnr_2 reg_out_B_MEM_reg_22__slave ( .q(reg_out_B_MEM[22]), .d(
        reg_out_B_MEM_reg_22__m2s), .g(Ctrl__Regs_1__en2), .rb(n5), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_MEM_reg_23__master ( .q(reg_out_B_MEM_reg_23__m2s), 
        .d(reg_out_B_EX[23]), .sdi(reg_out_B_MEM[22]), .se(test_se), .g(
        Ctrl__Regs_1__en1), .rb(n6), .glob_g(global_g1), .sync_sel(sync_sel)
         );
    mlatnr_2 reg_out_B_MEM_reg_23__slave ( .q(reg_out_B_MEM[23]), .d(
        reg_out_B_MEM_reg_23__m2s), .g(Ctrl__Regs_1__en2), .rb(n6), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_MEM_reg_24__master ( .q(reg_out_B_MEM_reg_24__m2s), 
        .d(reg_out_B_EX[24]), .sdi(reg_out_B_MEM[23]), .se(test_se), .g(
        Ctrl__Regs_1__en1), .rb(n4), .glob_g(global_g1), .sync_sel(sync_sel)
         );
    mlatnr_2 reg_out_B_MEM_reg_24__slave ( .q(reg_out_B_MEM[24]), .d(
        reg_out_B_MEM_reg_24__m2s), .g(Ctrl__Regs_1__en2), .rb(n4), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_MEM_reg_25__master ( .q(reg_out_B_MEM_reg_25__m2s), 
        .d(reg_out_B_EX[25]), .sdi(reg_out_B_MEM[24]), .se(test_se), .g(
        Ctrl__Regs_1__en1), .rb(n5), .glob_g(global_g1), .sync_sel(sync_sel)
         );
    mlatnr_2 reg_out_B_MEM_reg_25__slave ( .q(reg_out_B_MEM[25]), .d(
        reg_out_B_MEM_reg_25__m2s), .g(Ctrl__Regs_1__en2), .rb(n5), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_MEM_reg_26__master ( .q(reg_out_B_MEM_reg_26__m2s), 
        .d(reg_out_B_EX[26]), .sdi(reg_out_B_MEM[25]), .se(test_se), .g(
        Ctrl__Regs_1__en1), .rb(n6), .glob_g(global_g1), .sync_sel(sync_sel)
         );
    mlatnr_2 reg_out_B_MEM_reg_26__slave ( .q(reg_out_B_MEM[26]), .d(
        reg_out_B_MEM_reg_26__m2s), .g(Ctrl__Regs_1__en2), .rb(n6), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_MEM_reg_27__master ( .q(reg_out_B_MEM_reg_27__m2s), 
        .d(reg_out_B_EX[27]), .sdi(reg_out_B_MEM[26]), .se(test_se), .g(
        Ctrl__Regs_1__en1), .rb(n4), .glob_g(global_g1), .sync_sel(sync_sel)
         );
    mlatnr_2 reg_out_B_MEM_reg_27__slave ( .q(reg_out_B_MEM[27]), .d(
        reg_out_B_MEM_reg_27__m2s), .g(Ctrl__Regs_1__en2), .rb(n4), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_MEM_reg_28__master ( .q(reg_out_B_MEM_reg_28__m2s), 
        .d(reg_out_B_EX[28]), .sdi(reg_out_B_MEM[27]), .se(test_se), .g(
        Ctrl__Regs_1__en1), .rb(n5), .glob_g(global_g1), .sync_sel(sync_sel)
         );
    mlatnr_2 reg_out_B_MEM_reg_28__slave ( .q(reg_out_B_MEM[28]), .d(
        reg_out_B_MEM_reg_28__m2s), .g(Ctrl__Regs_1__en2), .rb(n5), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_MEM_reg_29__master ( .q(reg_out_B_MEM_reg_29__m2s), 
        .d(reg_out_B_EX[29]), .sdi(reg_out_B_MEM[28]), .se(test_se), .g(
        Ctrl__Regs_1__en1), .rb(n4), .glob_g(global_g1), .sync_sel(sync_sel)
         );
    mlatnr_2 reg_out_B_MEM_reg_29__slave ( .q(reg_out_B_MEM[29]), .d(
        reg_out_B_MEM_reg_29__m2s), .g(Ctrl__Regs_1__en2), .rb(n4), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_MEM_reg_2__master ( .q(reg_out_B_MEM_reg_2__m2s), .d(
        reg_out_B_EX[2]), .sdi(reg_out_B_MEM[1]), .se(test_se), .g(
        Ctrl__Regs_1__en1), .rb(n5), .glob_g(global_g1), .sync_sel(sync_sel)
         );
    mlatnr_2 reg_out_B_MEM_reg_2__slave ( .q(reg_out_B_MEM[2]), .d(
        reg_out_B_MEM_reg_2__m2s), .g(Ctrl__Regs_1__en2), .rb(n5), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_MEM_reg_30__master ( .q(reg_out_B_MEM_reg_30__m2s), 
        .d(reg_out_B_EX[30]), .sdi(reg_out_B_MEM[29]), .se(test_se), .g(
        Ctrl__Regs_1__en1), .rb(n6), .glob_g(global_g1), .sync_sel(sync_sel)
         );
    mlatnr_2 reg_out_B_MEM_reg_30__slave ( .q(reg_out_B_MEM[30]), .d(
        reg_out_B_MEM_reg_30__m2s), .g(Ctrl__Regs_1__en2), .rb(n6), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_MEM_reg_31__master ( .q(reg_out_B_MEM_reg_31__m2s), 
        .d(reg_out_B_EX[31]), .sdi(reg_out_B_MEM[30]), .se(test_se), .g(
        Ctrl__Regs_1__en1), .rb(n5), .glob_g(global_g1), .sync_sel(sync_sel)
         );
    mlatnr_2 reg_out_B_MEM_reg_31__slave ( .q(reg_out_B_MEM[31]), .d(
        reg_out_B_MEM_reg_31__m2s), .g(Ctrl__Regs_1__en2), .rb(n5), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_MEM_reg_3__master ( .q(reg_out_B_MEM_reg_3__m2s), .d(
        reg_out_B_EX[3]), .sdi(reg_out_B_MEM[2]), .se(test_se), .g(
        Ctrl__Regs_1__en1), .rb(n4), .glob_g(global_g1), .sync_sel(sync_sel)
         );
    mlatnr_2 reg_out_B_MEM_reg_3__slave ( .q(reg_out_B_MEM[3]), .d(
        reg_out_B_MEM_reg_3__m2s), .g(Ctrl__Regs_1__en2), .rb(n4), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_MEM_reg_4__master ( .q(reg_out_B_MEM_reg_4__m2s), .d(
        reg_out_B_EX[4]), .sdi(reg_out_B_MEM[3]), .se(test_se), .g(
        Ctrl__Regs_1__en1), .rb(n4), .glob_g(global_g1), .sync_sel(sync_sel)
         );
    mlatnr_2 reg_out_B_MEM_reg_4__slave ( .q(reg_out_B_MEM[4]), .d(
        reg_out_B_MEM_reg_4__m2s), .g(Ctrl__Regs_1__en2), .rb(n4), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_MEM_reg_5__master ( .q(reg_out_B_MEM_reg_5__m2s), .d(
        reg_out_B_EX[5]), .sdi(reg_out_B_MEM[4]), .se(test_se), .g(
        Ctrl__Regs_1__en1), .rb(n6), .glob_g(global_g1), .sync_sel(sync_sel)
         );
    mlatnr_2 reg_out_B_MEM_reg_5__slave ( .q(reg_out_B_MEM[5]), .d(
        reg_out_B_MEM_reg_5__m2s), .g(Ctrl__Regs_1__en2), .rb(n6), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_MEM_reg_6__master ( .q(reg_out_B_MEM_reg_6__m2s), .d(
        reg_out_B_EX[6]), .sdi(reg_out_B_MEM[5]), .se(test_se), .g(
        Ctrl__Regs_1__en1), .rb(n5), .glob_g(global_g1), .sync_sel(sync_sel)
         );
    mlatnr_2 reg_out_B_MEM_reg_6__slave ( .q(reg_out_B_MEM[6]), .d(
        reg_out_B_MEM_reg_6__m2s), .g(Ctrl__Regs_1__en2), .rb(n5), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_MEM_reg_7__master ( .q(reg_out_B_MEM_reg_7__m2s), .d(
        reg_out_B_EX[7]), .sdi(reg_out_B_MEM[6]), .se(test_se), .g(
        Ctrl__Regs_1__en1), .rb(n4), .glob_g(global_g1), .sync_sel(sync_sel)
         );
    mlatnr_2 reg_out_B_MEM_reg_7__slave ( .q(reg_out_B_MEM[7]), .d(
        reg_out_B_MEM_reg_7__m2s), .g(Ctrl__Regs_1__en2), .rb(n4), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_MEM_reg_8__master ( .q(reg_out_B_MEM_reg_8__m2s), .d(
        reg_out_B_EX[8]), .sdi(reg_out_B_MEM[7]), .se(test_se), .g(
        Ctrl__Regs_1__en1), .rb(n6), .glob_g(global_g1), .sync_sel(sync_sel)
         );
    mlatnr_2 reg_out_B_MEM_reg_8__slave ( .q(reg_out_B_MEM[8]), .d(
        reg_out_B_MEM_reg_8__m2s), .g(Ctrl__Regs_1__en2), .rb(n6), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_out_B_MEM_reg_9__master ( .q(reg_out_B_MEM_reg_9__m2s), .d(
        reg_out_B_EX[9]), .sdi(reg_out_B_MEM[8]), .se(test_se), .g(
        Ctrl__Regs_1__en1), .rb(n6), .glob_g(global_g1), .sync_sel(sync_sel)
         );
    mlatnr_2 reg_out_B_MEM_reg_9__slave ( .q(reg_out_B_MEM[9]), .d(
        reg_out_B_MEM_reg_9__m2s), .g(Ctrl__Regs_1__en2), .rb(n6), .glob_g(
        global_g2), .sync_sel(sync_sel) );
    smlatnr_1 reg_write_MEM_reg__master ( .q(reg_write_MEM_reg__m2s), .d(
        reg_write_EX), .sdi(reg_out_B_MEM[31]), .se(test_se), .g(
        Ctrl__Regs_1__en1), .rb(n6), .glob_g(global_g1), .sync_sel(sync_sel)
         );
    mlatnr_2 reg_write_MEM_reg__slave ( .q(reg_write_MEM), .qb(test_so), .d(
        reg_write_MEM_reg__m2s), .g(Ctrl__Regs_1__en2), .rb(n6), .glob_g(
        global_g2), .sync_sel(sync_sel) );
endmodule


module DLX_sync_desync ( DM_read_data, DM_write_data, DM_addr, DM_write, 
    DM_read, NPC, reset, IR, byte0, word, INT, CLI, PIPEEMPTY, FREEZE, test_si, 
    test_se, sync_sel, global_g1, global_g2, Ctrl__EXinst___Regs_1__en1, 
    Ctrl__EXinst___Regs_1__en2, Ctrl__IDinst___Regs_1__en1, 
    Ctrl__IDinst___Regs_1__en2, Ctrl__IFinst___Regs_1__en1, 
    Ctrl__IFinst___Regs_1__en2, Ctrl__MEMinst___Regs_1__en1, 
    Ctrl__MEMinst___Regs_1__en2 );
input  [31:0] DM_read_data;
output [31:0] DM_write_data;
output [31:0] DM_addr;
output [31:0] NPC;
input  [31:0] IR;
input  reset, INT, FREEZE, test_si, test_se, sync_sel, global_g1, global_g2, 
    Ctrl__EXinst___Regs_1__en1, Ctrl__EXinst___Regs_1__en2, 
    Ctrl__IDinst___Regs_1__en1, Ctrl__IDinst___Regs_1__en2, 
    Ctrl__IFinst___Regs_1__en1, Ctrl__IFinst___Regs_1__en2, 
    Ctrl__MEMinst___Regs_1__en1, Ctrl__MEMinst___Regs_1__en2;
output DM_write, DM_read, byte0, word, CLI, PIPEEMPTY;
    wire mem_to_reg_EX, reg_write_EX, reg_dst, reg_write, mem_to_reg, mem_read, 
        mem_write, n14, counter_1_0, counter_0_0, Imm_31_0, Imm_30_0, Imm_29_0, 
        Imm_28_0, Imm_27_0, Imm_26_0, Imm_25_0, Imm_24_0, Imm_23_0, Imm_22_0, 
        Imm_21_0, Imm_20_0, Imm_19_0, Imm_18_0, Imm_17_0, Imm_16_0, Imm_15_0, 
        Imm_14_0, Imm_13_0, Imm_12_0, Imm_11_0, Imm_10_0, Imm_9_0, Imm_8_0, 
        Imm_7_0, Imm_6_0, Imm_5_0, Imm_4_0, Imm_3_0, Imm_2_0, Imm_1_0, Imm_0_0, 
        reg_out_B_31_0, reg_out_B_30_0, reg_out_B_29_0, reg_out_B_28_0, 
        reg_out_B_27_0, reg_out_B_26_0, reg_out_B_25_0, reg_out_B_24_0, 
        reg_out_B_23_0, reg_out_B_22_0, reg_out_B_21_0, reg_out_B_20_0, 
        reg_out_B_19_0, reg_out_B_18_0, reg_out_B_17_0, reg_out_B_16_0, 
        reg_out_B_15_0, reg_out_B_14_0, reg_out_B_13_0, reg_out_B_12_0, 
        reg_out_B_11_0, reg_out_B_10_0, reg_out_B_9_0, reg_out_B_8_0, 
        reg_out_B_7_0, reg_out_B_6_0, reg_out_B_5_0, reg_out_B_4_0, 
        reg_out_B_3_0, reg_out_B_2_0, reg_out_B_1_0, reg_out_B_0_0, 
        reg_out_A_31_0, reg_out_A_30_0, reg_out_A_29_0, reg_out_A_28_0, 
        reg_out_A_27_0, reg_out_A_26_0, reg_out_A_25_0, reg_out_A_24_0, 
        reg_out_A_23_0, reg_out_A_22_0, reg_out_A_21_0, reg_out_A_20_0, 
        reg_out_A_19_0, reg_out_A_18_0, reg_out_A_17_0, reg_out_A_16_0, 
        reg_out_A_15_0, reg_out_A_14_0, reg_out_A_13_0, reg_out_A_12_0, 
        reg_out_A_11_0, reg_out_A_10_0, reg_out_A_9_0, reg_out_A_8_0, 
        reg_out_A_7_0, reg_out_A_6_0, reg_out_A_5_0, reg_out_A_4_0, 
        reg_out_A_3_0, reg_out_A_2_0, reg_out_A_1_0, reg_out_A_0_0, 
        IR_function_field_5_0, IR_function_field_4_0, IR_function_field_3_0, 
        IR_function_field_2_0, IR_function_field_1_0, IR_function_field_0_0, 
        IR_opcode_field_5_0, IR_opcode_field_4_0, IR_opcode_field_3_0, 
        IR_opcode_field_2_0, IR_opcode_field_1_0, IR_opcode_field_0_0, 
        branch_sig, stall, reg_write_MEM, n13, RF_data_old_31_0, 
        RF_data_old_30_0, RF_data_old_29_0, RF_data_old_28_0, RF_data_old_27_0, 
        RF_data_old_26_0, RF_data_old_25_0, RF_data_old_24_0, RF_data_old_23_0, 
        RF_data_old_22_0, RF_data_old_21_0, RF_data_old_20_0, RF_data_old_19_0, 
        RF_data_old_18_0, RF_data_old_17_0, RF_data_old_16_0, RF_data_old_15_0, 
        RF_data_old_14_0, RF_data_old_13_0, RF_data_old_12_0, RF_data_old_11_0, 
        RF_data_old_10_0, RF_data_old_9_0, RF_data_old_8_0, RF_data_old_7_0, 
        RF_data_old_6_0, RF_data_old_5_0, RF_data_old_4_0, RF_data_old_3_0, 
        RF_data_old_2_0, RF_data_old_1_0, RF_data_old_0_0, RF_data_in_31_0, 
        RF_data_in_30_0, RF_data_in_29_0, RF_data_in_28_0, RF_data_in_27_0, 
        RF_data_in_26_0, RF_data_in_25_0, RF_data_in_24_0, RF_data_in_23_0, 
        RF_data_in_22_0, RF_data_in_21_0, RF_data_in_20_0, RF_data_in_19_0, 
        RF_data_in_18_0, RF_data_in_17_0, RF_data_in_16_0, RF_data_in_15_0, 
        RF_data_in_14_0, RF_data_in_13_0, RF_data_in_12_0, RF_data_in_11_0, 
        RF_data_in_10_0, RF_data_in_9_0, RF_data_in_8_0, RF_data_in_7_0, 
        RF_data_in_6_0, RF_data_in_5_0, RF_data_in_4_0, RF_data_in_3_0, 
        RF_data_in_2_0, RF_data_in_1_0, RF_data_in_0_0, IR_latched_31_0, 
        IR_latched_30_0, IR_latched_29_0, IR_latched_28_0, IR_latched_27_0, 
        IR_latched_26_0, IR_latched_25_0, IR_latched_24_0, IR_latched_23_0, 
        IR_latched_22_0, IR_latched_21_0, IR_latched_20_0, IR_latched_19_0, 
        IR_latched_18_0, IR_latched_17_0, IR_latched_16_0, IR_latched_15_0, 
        IR_latched_14_0, IR_latched_13_0, IR_latched_12_0, IR_latched_11_0, 
        IR_latched_10_0, IR_latched_9_0, IR_latched_8_0, IR_latched_7_0, 
        IR_latched_6_0, IR_latched_5_0, IR_latched_4_0, IR_latched_3_0, 
        IR_latched_2_0, IR_latched_1_0, IR_latched_0_0, n5, 
        branch_address_31_0, branch_address_30_0, branch_address_29_0, 
        branch_address_28_0, branch_address_27_0, branch_address_26_0, 
        branch_address_25_0, branch_address_24_0, branch_address_23_0, 
        branch_address_22_0, branch_address_21_0, branch_address_20_0, 
        branch_address_19_0, branch_address_18_0, branch_address_17_0, 
        branch_address_16_0, branch_address_15_0, branch_address_14_0, 
        branch_address_13_0, branch_address_12_0, branch_address_11_0, 
        branch_address_10_0, branch_address_9_0, branch_address_8_0, 
        branch_address_7_0, branch_address_6_0, branch_address_5_0, 
        branch_address_4_0, branch_address_3_0, branch_address_2_0, 
        branch_address_1_0, branch_address_0_0, n12, n11, n4, n16, n17, n2, n6, 
        n8;
    EX_test_1_desync EXinst ( .ALU_result(DM_addr), .reg_out_B_EX(
        DM_write_data), .mem_write_EX(DM_write), .mem_read_EX(DM_read), 
        .mem_to_reg_EX(mem_to_reg_EX), .reg_write_EX(reg_write_EX), .reset(
        reset), .IR_opcode_field({IR_opcode_field_5_0, IR_opcode_field_4_0, 
        IR_opcode_field_3_0, IR_opcode_field_2_0, IR_opcode_field_1_0, 
        IR_opcode_field_0_0}), .IR_function_field({IR_function_field_5_0, 
        IR_function_field_4_0, IR_function_field_3_0, IR_function_field_2_0, 
        IR_function_field_1_0, IR_function_field_0_0}), .reg_out_A({
        reg_out_A_31_0, reg_out_A_30_0, reg_out_A_29_0, reg_out_A_28_0, 
        reg_out_A_27_0, reg_out_A_26_0, reg_out_A_25_0, reg_out_A_24_0, 
        reg_out_A_23_0, reg_out_A_22_0, reg_out_A_21_0, reg_out_A_20_0, 
        reg_out_A_19_0, reg_out_A_18_0, reg_out_A_17_0, reg_out_A_16_0, 
        reg_out_A_15_0, reg_out_A_14_0, reg_out_A_13_0, reg_out_A_12_0, 
        reg_out_A_11_0, reg_out_A_10_0, reg_out_A_9_0, reg_out_A_8_0, 
        reg_out_A_7_0, reg_out_A_6_0, reg_out_A_5_0, reg_out_A_4_0, 
        reg_out_A_3_0, reg_out_A_2_0, reg_out_A_1_0, reg_out_A_0_0}), 
        .reg_out_B({reg_out_B_31_0, reg_out_B_30_0, reg_out_B_29_0, 
        reg_out_B_28_0, reg_out_B_27_0, reg_out_B_26_0, reg_out_B_25_0, 
        reg_out_B_24_0, reg_out_B_23_0, reg_out_B_22_0, reg_out_B_21_0, 
        reg_out_B_20_0, reg_out_B_19_0, reg_out_B_18_0, reg_out_B_17_0, 
        reg_out_B_16_0, reg_out_B_15_0, reg_out_B_14_0, reg_out_B_13_0, 
        reg_out_B_12_0, reg_out_B_11_0, reg_out_B_10_0, reg_out_B_9_0, 
        reg_out_B_8_0, reg_out_B_7_0, reg_out_B_6_0, reg_out_B_5_0, 
        reg_out_B_4_0, reg_out_B_3_0, reg_out_B_2_0, reg_out_B_1_0, 
        reg_out_B_0_0}), .Imm({Imm_31_0, Imm_30_0, Imm_29_0, Imm_28_0, 
        Imm_27_0, Imm_26_0, Imm_25_0, Imm_24_0, Imm_23_0, Imm_22_0, Imm_21_0, 
        Imm_20_0, Imm_19_0, Imm_18_0, Imm_17_0, Imm_16_0, Imm_15_0, Imm_14_0, 
        Imm_13_0, Imm_12_0, Imm_11_0, Imm_10_0, Imm_9_0, Imm_8_0, Imm_7_0, 
        Imm_6_0, Imm_5_0, Imm_4_0, Imm_3_0, Imm_2_0, Imm_1_0, Imm_0_0}), 
        .reg_dst(reg_dst), .reg_write(reg_write), .mem_to_reg(mem_to_reg), 
        .mem_read(mem_read), .mem_write(mem_write), ._byte(byte0), .word(word), 
        .counter({counter_1_0, counter_0_0}), .test_si(test_si), .test_so(n14), 
        .test_se(test_se), .sync_sel(sync_sel), .global_g1(global_g1), 
        .global_g2(global_g2), .Ctrl__Regs_1__en1(Ctrl__EXinst___Regs_1__en1), 
        .Ctrl__Regs_1__en2(Ctrl__EXinst___Regs_1__en2) );
    ID_test_1_desync IDinst ( .INT(INT), .CLI(CLI), .PIPEEMPTY(PIPEEMPTY), 
        .FREEZE(FREEZE), .branch_address({branch_address_31_0, 
        branch_address_30_0, branch_address_29_0, branch_address_28_0, 
        branch_address_27_0, branch_address_26_0, branch_address_25_0, 
        branch_address_24_0, branch_address_23_0, branch_address_22_0, 
        branch_address_21_0, branch_address_20_0, branch_address_19_0, 
        branch_address_18_0, branch_address_17_0, branch_address_16_0, 
        branch_address_15_0, branch_address_14_0, branch_address_13_0, 
        branch_address_12_0, branch_address_11_0, branch_address_10_0, 
        branch_address_9_0, branch_address_8_0, branch_address_7_0, 
        branch_address_6_0, branch_address_5_0, branch_address_4_0, 
        branch_address_3_0, branch_address_2_0, branch_address_1_0, 
        branch_address_0_0}), .branch_sig(branch_sig), .Imm({Imm_31_0, 
        Imm_30_0, Imm_29_0, Imm_28_0, Imm_27_0, Imm_26_0, Imm_25_0, Imm_24_0, 
        Imm_23_0, Imm_22_0, Imm_21_0, Imm_20_0, Imm_19_0, Imm_18_0, Imm_17_0, 
        Imm_16_0, Imm_15_0, Imm_14_0, Imm_13_0, Imm_12_0, Imm_11_0, Imm_10_0, 
        Imm_9_0, Imm_8_0, Imm_7_0, Imm_6_0, Imm_5_0, Imm_4_0, Imm_3_0, Imm_2_0, 
        Imm_1_0, Imm_0_0}), .reg_dst(reg_dst), .reg_write(reg_write), 
        .mem_to_reg(mem_to_reg), .mem_write(mem_write), .mem_read(mem_read), 
        .IR_opcode_field({IR_opcode_field_5_0, IR_opcode_field_4_0, 
        IR_opcode_field_3_0, IR_opcode_field_2_0, IR_opcode_field_1_0, 
        IR_opcode_field_0_0}), .IR_function_field({IR_function_field_5_0, 
        IR_function_field_4_0, IR_function_field_3_0, IR_function_field_2_0, 
        IR_function_field_1_0, IR_function_field_0_0}), .stall(stall), 
        .counter({counter_1_0, counter_0_0}), .reset(reset), .NPC({NPC[31], 
        NPC[30], NPC[29], NPC[28], NPC[27], NPC[26], NPC[25], NPC[24], NPC[23], 
        NPC[22], NPC[21], NPC[20], NPC[19], NPC[18], NPC[17], NPC[16], NPC[15], 
        NPC[14], NPC[13], NPC[12], NPC[11], NPC[10], NPC[9], NPC[8], NPC[7], 
        NPC[6], NPC[5], NPC[4], NPC[3], n5, NPC[1], NPC[0]}), 
        .IR_latched_input({IR_latched_31_0, IR_latched_30_0, IR_latched_29_0, 
        IR_latched_28_0, IR_latched_27_0, IR_latched_26_0, IR_latched_25_0, 
        IR_latched_24_0, IR_latched_23_0, IR_latched_22_0, IR_latched_21_0, 
        IR_latched_20_0, IR_latched_19_0, IR_latched_18_0, IR_latched_17_0, 
        IR_latched_16_0, IR_latched_15_0, IR_latched_14_0, IR_latched_13_0, 
        IR_latched_12_0, IR_latched_11_0, IR_latched_10_0, IR_latched_9_0, 
        IR_latched_8_0, IR_latched_7_0, IR_latched_6_0, IR_latched_5_0, 
        IR_latched_4_0, IR_latched_3_0, IR_latched_2_0, IR_latched_1_0, 
        IR_latched_0_0}), .reg_out_A({reg_out_A_31_0, reg_out_A_30_0, 
        reg_out_A_29_0, reg_out_A_28_0, reg_out_A_27_0, reg_out_A_26_0, 
        reg_out_A_25_0, reg_out_A_24_0, reg_out_A_23_0, reg_out_A_22_0, 
        reg_out_A_21_0, reg_out_A_20_0, reg_out_A_19_0, reg_out_A_18_0, 
        reg_out_A_17_0, reg_out_A_16_0, reg_out_A_15_0, reg_out_A_14_0, 
        reg_out_A_13_0, reg_out_A_12_0, reg_out_A_11_0, reg_out_A_10_0, 
        reg_out_A_9_0, reg_out_A_8_0, reg_out_A_7_0, reg_out_A_6_0, 
        reg_out_A_5_0, reg_out_A_4_0, reg_out_A_3_0, reg_out_A_2_0, 
        reg_out_A_1_0, reg_out_A_0_0}), .reg_out_B({reg_out_B_31_0, 
        reg_out_B_30_0, reg_out_B_29_0, reg_out_B_28_0, reg_out_B_27_0, 
        reg_out_B_26_0, reg_out_B_25_0, reg_out_B_24_0, reg_out_B_23_0, 
        reg_out_B_22_0, reg_out_B_21_0, reg_out_B_20_0, reg_out_B_19_0, 
        reg_out_B_18_0, reg_out_B_17_0, reg_out_B_16_0, reg_out_B_15_0, 
        reg_out_B_14_0, reg_out_B_13_0, reg_out_B_12_0, reg_out_B_11_0, 
        reg_out_B_10_0, reg_out_B_9_0, reg_out_B_8_0, reg_out_B_7_0, 
        reg_out_B_6_0, reg_out_B_5_0, reg_out_B_4_0, reg_out_B_3_0, 
        reg_out_B_2_0, reg_out_B_1_0, reg_out_B_0_0}), .reg_write_WB(
        reg_write_MEM), .WB_data({RF_data_in_31_0, RF_data_in_30_0, 
        RF_data_in_29_0, RF_data_in_28_0, RF_data_in_27_0, RF_data_in_26_0, 
        RF_data_in_25_0, RF_data_in_24_0, RF_data_in_23_0, RF_data_in_22_0, 
        RF_data_in_21_0, RF_data_in_20_0, RF_data_in_19_0, RF_data_in_18_0, 
        RF_data_in_17_0, RF_data_in_16_0, RF_data_in_15_0, RF_data_in_14_0, 
        RF_data_in_13_0, RF_data_in_12_0, RF_data_in_11_0, RF_data_in_10_0, 
        RF_data_in_9_0, RF_data_in_8_0, RF_data_in_7_0, RF_data_in_6_0, 
        RF_data_in_5_0, RF_data_in_4_0, RF_data_in_3_0, RF_data_in_2_0, 
        RF_data_in_1_0, RF_data_in_0_0}), .WB_data_old({RF_data_old_31_0, 
        RF_data_old_30_0, RF_data_old_29_0, RF_data_old_28_0, RF_data_old_27_0, 
        RF_data_old_26_0, RF_data_old_25_0, RF_data_old_24_0, RF_data_old_23_0, 
        RF_data_old_22_0, RF_data_old_21_0, RF_data_old_20_0, RF_data_old_19_0, 
        RF_data_old_18_0, RF_data_old_17_0, RF_data_old_16_0, RF_data_old_15_0, 
        RF_data_old_14_0, RF_data_old_13_0, RF_data_old_12_0, RF_data_old_11_0, 
        RF_data_old_10_0, RF_data_old_9_0, RF_data_old_8_0, RF_data_old_7_0, 
        RF_data_old_6_0, RF_data_old_5_0, RF_data_old_4_0, RF_data_old_3_0, 
        RF_data_old_2_0, RF_data_old_1_0, RF_data_old_0_0}), .test_si(n14), 
        .test_so(n13), .test_se(test_se), .sync_sel(sync_sel), .global_g1(
        global_g1), .global_g2(global_g2), .Ctrl__Regs_1__en1(
        Ctrl__IDinst___Regs_1__en1), .Ctrl__Regs_1__en2(
        Ctrl__IDinst___Regs_1__en2) );
    IF_test_1_desync IFinst ( .NPC({NPC[31], NPC[30], NPC[29], NPC[28], 
        NPC[27], NPC[26], NPC[25], NPC[24], NPC[23], NPC[22], NPC[21], NPC[20], 
        NPC[19], NPC[18], NPC[17], NPC[16], NPC[15], NPC[14], NPC[13], n4, 
        NPC[11], n16, NPC[9], NPC[8], n17, NPC[6], NPC[5], NPC[4], NPC[3], n5, 
        NPC[1], NPC[0]}), .IR_latched({IR_latched_31_0, IR_latched_30_0, 
        IR_latched_29_0, IR_latched_28_0, IR_latched_27_0, IR_latched_26_0, 
        IR_latched_25_0, IR_latched_24_0, IR_latched_23_0, IR_latched_22_0, 
        IR_latched_21_0, IR_latched_20_0, IR_latched_19_0, IR_latched_18_0, 
        IR_latched_17_0, IR_latched_16_0, IR_latched_15_0, IR_latched_14_0, 
        IR_latched_13_0, IR_latched_12_0, IR_latched_11_0, IR_latched_10_0, 
        IR_latched_9_0, IR_latched_8_0, IR_latched_7_0, IR_latched_6_0, 
        IR_latched_5_0, IR_latched_4_0, IR_latched_3_0, IR_latched_2_0, 
        IR_latched_1_0, IR_latched_0_0}), .reset(reset), .branch_sig(
        branch_sig), .branch_address({branch_address_31_0, branch_address_30_0, 
        branch_address_29_0, branch_address_28_0, branch_address_27_0, 
        branch_address_26_0, branch_address_25_0, branch_address_24_0, 
        branch_address_23_0, branch_address_22_0, branch_address_21_0, 
        branch_address_20_0, branch_address_19_0, branch_address_18_0, 
        branch_address_17_0, branch_address_16_0, branch_address_15_0, 
        branch_address_14_0, branch_address_13_0, branch_address_12_0, 
        branch_address_11_0, branch_address_10_0, branch_address_9_0, 
        branch_address_8_0, branch_address_7_0, branch_address_6_0, 
        branch_address_5_0, branch_address_4_0, branch_address_3_0, 
        branch_address_2_0, branch_address_1_0, branch_address_0_0}), .IR(IR), 
        .stall(stall), .counter({counter_1_0, counter_0_0}), .test_si1(n13), 
        .test_so1(n12), .test_si2(n11), .test_se(test_se), .sync_sel(sync_sel), 
        .global_g1(global_g1), .global_g2(global_g2), .Ctrl__Regs_1__en1(
        Ctrl__IFinst___Regs_1__en1), .Ctrl__Regs_1__en2(
        Ctrl__IFinst___Regs_1__en2) );
    MEM_test_1_desync MEMinst ( .reg_write_MEM(reg_write_MEM), .mem_to_reg_EX(
        mem_to_reg_EX), .reset(reset), .ALU_result(DM_addr), .reg_write_EX(
        reg_write_EX), .reg_out_B_EX(DM_write_data), .reg_out_B_MEM({
        RF_data_old_31_0, RF_data_old_30_0, RF_data_old_29_0, RF_data_old_28_0, 
        RF_data_old_27_0, RF_data_old_26_0, RF_data_old_25_0, RF_data_old_24_0, 
        RF_data_old_23_0, RF_data_old_22_0, RF_data_old_21_0, RF_data_old_20_0, 
        RF_data_old_19_0, RF_data_old_18_0, RF_data_old_17_0, RF_data_old_16_0, 
        RF_data_old_15_0, RF_data_old_14_0, RF_data_old_13_0, RF_data_old_12_0, 
        RF_data_old_11_0, RF_data_old_10_0, RF_data_old_9_0, RF_data_old_8_0, 
        RF_data_old_7_0, RF_data_old_6_0, RF_data_old_5_0, RF_data_old_4_0, 
        RF_data_old_3_0, RF_data_old_2_0, RF_data_old_1_0, RF_data_old_0_0}), 
        .DM_read_data(DM_read_data), .RF_data_in({RF_data_in_31_0, 
        RF_data_in_30_0, RF_data_in_29_0, RF_data_in_28_0, RF_data_in_27_0, 
        RF_data_in_26_0, RF_data_in_25_0, RF_data_in_24_0, RF_data_in_23_0, 
        RF_data_in_22_0, RF_data_in_21_0, RF_data_in_20_0, RF_data_in_19_0, 
        RF_data_in_18_0, RF_data_in_17_0, RF_data_in_16_0, RF_data_in_15_0, 
        RF_data_in_14_0, RF_data_in_13_0, RF_data_in_12_0, RF_data_in_11_0, 
        RF_data_in_10_0, RF_data_in_9_0, RF_data_in_8_0, RF_data_in_7_0, 
        RF_data_in_6_0, RF_data_in_5_0, RF_data_in_4_0, RF_data_in_3_0, 
        RF_data_in_2_0, RF_data_in_1_0, RF_data_in_0_0}), .test_si(n12), 
        .test_so(n11), .test_se(test_se), .sync_sel(sync_sel), .global_g1(
        global_g1), .global_g2(global_g2), .Ctrl__Regs_1__en1(
        Ctrl__MEMinst___Regs_1__en1), .Ctrl__Regs_1__en2(
        Ctrl__MEMinst___Regs_1__en2) );
    buf_10 U1 ( .x(NPC[12]), .a(n4) );
    inv_0 U2 ( .x(n2), .a(n5) );
    inv_2 U3 ( .x(NPC[2]), .a(n2) );
    inv_6 U4 ( .x(n6), .a(n16) );
    inv_10 U5 ( .x(NPC[10]), .a(n6) );
    inv_6 U6 ( .x(n8), .a(n17) );
    inv_10 U7 ( .x(NPC[7]), .a(n8) );
endmodule


module DLX_sync_desync_with_ctrls ( DM_read_data, DM_write_data, DM_addr, 
    DM_write, DM_read, NPC, reset, IR, byte0, word, INT, CLI, PIPEEMPTY, 
    FREEZE, test_si, test_se, sync_sel, global_g1, global_g2, Ctrl__reset, 
    Ctrl__EXinst___Regs_1__ai, Ctrl__IDinst___Regs_1__ai, 
    Ctrl__IDinst___Regs_1__ro, Ctrl__MEMinst___Regs_1__ro, 
    Ctrl__IFinst___Regs_1__ri, Ctrl__IFinst___Regs_1__ai, 
    Ctrl__MEMinst___Regs_1__ri, Ctrl__MEMinst___Regs_1__ai, 
    Ctrl__EXinst___Regs_1__ro, Ctrl__EXinst___Regs_1__ao, 
    Ctrl__IFinst___Regs_1__ro, Ctrl__IFinst___Regs_1__ao, 
    Ctrl__EXinst___Regs_1__delay_mux_sel, Ctrl__IDinst___Regs_1__delay_mux_sel, 
    Ctrl__IFinst___Regs_1__delay_mux_sel, 
    Ctrl__MEMinst___Regs_1__delay_mux_sel, Ctrl__EXinst___Regs_1__en1, 
    Ctrl__EXinst___Regs_1__en2, Ctrl__IDinst___Regs_1__en1, 
    Ctrl__IDinst___Regs_1__en2, Ctrl__IFinst___Regs_1__en1, 
    Ctrl__IFinst___Regs_1__en2, Ctrl__MEMinst___Regs_1__en1, 
    Ctrl__MEMinst___Regs_1__en2 );
input  [31:0] DM_read_data;
output [31:0] DM_write_data;
output [31:0] DM_addr;
output [31:0] NPC;
input  [31:0] IR;
input  [1:0] Ctrl__EXinst___Regs_1__delay_mux_sel;
input  [1:0] Ctrl__IDinst___Regs_1__delay_mux_sel;
input  [1:0] Ctrl__IFinst___Regs_1__delay_mux_sel;
input  [1:0] Ctrl__MEMinst___Regs_1__delay_mux_sel;
input  reset, INT, FREEZE, test_si, test_se, sync_sel, global_g1, global_g2, 
    Ctrl__reset, Ctrl__IFinst___Regs_1__ri, Ctrl__MEMinst___Regs_1__ri, 
    Ctrl__EXinst___Regs_1__ao, Ctrl__IFinst___Regs_1__ao;
output DM_write, DM_read, byte0, word, CLI, PIPEEMPTY, 
    Ctrl__EXinst___Regs_1__ai, Ctrl__IDinst___Regs_1__ai, 
    Ctrl__IDinst___Regs_1__ro, Ctrl__MEMinst___Regs_1__ro, 
    Ctrl__IFinst___Regs_1__ai, Ctrl__MEMinst___Regs_1__ai, 
    Ctrl__EXinst___Regs_1__ro, Ctrl__IFinst___Regs_1__ro, 
    Ctrl__EXinst___Regs_1__en1, Ctrl__EXinst___Regs_1__en2, 
    Ctrl__IDinst___Regs_1__en1, Ctrl__IDinst___Regs_1__en2, 
    Ctrl__IFinst___Regs_1__en1, Ctrl__IFinst___Regs_1__en2, 
    Ctrl__MEMinst___Regs_1__en1, Ctrl__MEMinst___Regs_1__en2;
    controller_d32__0_85__1__1_38__1_77_r1_a2 Ctrl__EXinst___Regs_1 ( .reset(
        Ctrl__reset), .en1(Ctrl__EXinst___Regs_1__en1), .en2(
        Ctrl__EXinst___Regs_1__en2), .ri1(Ctrl__IDinst___Regs_1__ro), .ai(
        Ctrl__EXinst___Regs_1__ai), .ro(Ctrl__EXinst___Regs_1__ro), .ao1(
        Ctrl__EXinst___Regs_1__ao), .ao2(Ctrl__MEMinst___Regs_1__ai), 
        .delay_mux_sel(Ctrl__EXinst___Regs_1__delay_mux_sel) );
    controller_d31__0_85__1__1_47__1_93_r2_a2 Ctrl__IDinst___Regs_1 ( .reset(
        Ctrl__reset), .en1(Ctrl__IDinst___Regs_1__en1), .en2(
        Ctrl__IDinst___Regs_1__en2), .ri1(Ctrl__IFinst___Regs_1__ro), .ri2(
        Ctrl__MEMinst___Regs_1__ro), .ai(Ctrl__IDinst___Regs_1__ai), .ro(
        Ctrl__IDinst___Regs_1__ro), .ao1(Ctrl__EXinst___Regs_1__ai), .ao2(
        Ctrl__IFinst___Regs_1__ai), .delay_mux_sel(
        Ctrl__IDinst___Regs_1__delay_mux_sel) );
    controller_d28__0_85__1__1_48__1_95_r2_a2 Ctrl__IFinst___Regs_1 ( .reset(
        Ctrl__reset), .en1(Ctrl__IFinst___Regs_1__en1), .en2(
        Ctrl__IFinst___Regs_1__en2), .ri1(Ctrl__IFinst___Regs_1__ri), .ri2(
        Ctrl__IDinst___Regs_1__ro), .ai(Ctrl__IFinst___Regs_1__ai), .ro(
        Ctrl__IFinst___Regs_1__ro), .ao1(Ctrl__IFinst___Regs_1__ao), .ao2(
        Ctrl__IDinst___Regs_1__ai), .delay_mux_sel(
        Ctrl__IFinst___Regs_1__delay_mux_sel) );
    controller_d6__0_85__1__1_18__1_36_r2_a1 Ctrl__MEMinst___Regs_1 ( .reset(
        Ctrl__reset), .en1(Ctrl__MEMinst___Regs_1__en1), .en2(
        Ctrl__MEMinst___Regs_1__en2), .ri1(Ctrl__MEMinst___Regs_1__ri), .ri2(
        Ctrl__EXinst___Regs_1__ro), .ai(Ctrl__MEMinst___Regs_1__ai), .ro(
        Ctrl__MEMinst___Regs_1__ro), .ao1(Ctrl__IDinst___Regs_1__ai), 
        .delay_mux_sel(Ctrl__MEMinst___Regs_1__delay_mux_sel) );
    DLX_sync_desync DLX_sync ( .DM_read_data(DM_read_data), .DM_write_data(
        DM_write_data), .DM_addr(DM_addr), .DM_write(DM_write), .DM_read(
        DM_read), .NPC(NPC), .reset(reset), .IR(IR), .byte0(byte0), .word(word
        ), .INT(INT), .CLI(CLI), .PIPEEMPTY(PIPEEMPTY), .FREEZE(FREEZE), 
        .test_si(test_si), .test_se(test_se), .sync_sel(sync_sel), .global_g1(
        global_g1), .global_g2(global_g2), .Ctrl__EXinst___Regs_1__en1(
        Ctrl__EXinst___Regs_1__en1), .Ctrl__EXinst___Regs_1__en2(
        Ctrl__EXinst___Regs_1__en2), .Ctrl__IDinst___Regs_1__en1(
        Ctrl__IDinst___Regs_1__en1), .Ctrl__IDinst___Regs_1__en2(
        Ctrl__IDinst___Regs_1__en2), .Ctrl__IFinst___Regs_1__en1(
        Ctrl__IFinst___Regs_1__en1), .Ctrl__IFinst___Regs_1__en2(
        Ctrl__IFinst___Regs_1__en2), .Ctrl__MEMinst___Regs_1__en1(
        Ctrl__MEMinst___Regs_1__en1), .Ctrl__MEMinst___Regs_1__en2(
        Ctrl__MEMinst___Regs_1__en2) );
endmodule


module mem_if ( DM_addr_CPU, DM_read_data_CPU, DM_write_data_CPU, word, \byte , 
    DM_addr_MEM, DM_read_data_MEM, DM_write_data_MEM, DM_write, mask );
input  [31:0] DM_addr_CPU;
output [31:0] DM_read_data_CPU;
input  [31:0] DM_write_data_CPU;
output [8:0] DM_addr_MEM;
input  [31:0] DM_read_data_MEM;
output [31:0] DM_write_data_MEM;
output [3:0] mask;
input  word, \byte , DM_write;
    wire DM_addr_CPU_10, DM_addr_CPU_9, DM_addr_CPU_8, DM_addr_CPU_7, 
        DM_addr_CPU_6, DM_addr_CPU_5, DM_addr_CPU_4, DM_addr_CPU_3, 
        DM_addr_CPU_2, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, 
        n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, 
        n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, 
        n67, n68, n69, n70, n71, n72, n73, n74, n75, n76;
    assign DM_addr_CPU_10 = DM_addr_CPU[10];
    assign DM_addr_CPU_9 = DM_addr_CPU[9];
    assign DM_addr_CPU_8 = DM_addr_CPU[8];
    assign DM_addr_CPU_7 = DM_addr_CPU[7];
    assign DM_addr_CPU_6 = DM_addr_CPU[6];
    assign DM_addr_CPU_5 = DM_addr_CPU[5];
    assign DM_addr_CPU_4 = DM_addr_CPU[4];
    assign DM_addr_CPU_3 = DM_addr_CPU[3];
    assign DM_addr_CPU_2 = DM_addr_CPU[2];
    assign DM_addr_MEM[8] = DM_addr_CPU_10;
    assign DM_addr_MEM[7] = DM_addr_CPU_9;
    assign DM_addr_MEM[6] = DM_addr_CPU_8;
    assign DM_addr_MEM[5] = DM_addr_CPU_7;
    assign DM_addr_MEM[4] = DM_addr_CPU_6;
    assign DM_addr_MEM[3] = DM_addr_CPU_5;
    assign DM_addr_MEM[2] = DM_addr_CPU_4;
    assign DM_addr_MEM[1] = DM_addr_CPU_3;
    assign DM_addr_MEM[0] = DM_addr_CPU_2;
    mx4_1 U3 ( .x(DM_read_data_CPU[7]), .d0(DM_read_data_MEM[7]), .sl0(mask[0]
        ), .d1(DM_read_data_MEM[23]), .sl1(n32), .d2(DM_read_data_MEM[31]), 
        .sl2(n30), .d3(DM_read_data_MEM[15]), .sl3(n33) );
    mx4_1 U4 ( .x(DM_read_data_CPU[6]), .d0(DM_read_data_MEM[6]), .sl0(mask[0]
        ), .d1(DM_read_data_MEM[22]), .sl1(n32), .d2(DM_read_data_MEM[30]), 
        .sl2(n30), .d3(DM_read_data_MEM[14]), .sl3(n33) );
    mx4_1 U5 ( .x(DM_read_data_CPU[5]), .d0(DM_read_data_MEM[5]), .sl0(mask[0]
        ), .d1(DM_read_data_MEM[21]), .sl1(n32), .d2(DM_read_data_MEM[29]), 
        .sl2(n30), .d3(DM_read_data_MEM[13]), .sl3(n33) );
    mx4_1 U6 ( .x(DM_read_data_CPU[4]), .d0(DM_read_data_MEM[4]), .sl0(mask[0]
        ), .d1(DM_read_data_MEM[20]), .sl1(n32), .d2(DM_read_data_MEM[28]), 
        .sl2(n30), .d3(DM_read_data_MEM[12]), .sl3(n33) );
    mx4_1 U7 ( .x(DM_read_data_CPU[3]), .d0(DM_read_data_MEM[3]), .sl0(mask[0]
        ), .d1(DM_read_data_MEM[19]), .sl1(n32), .d2(DM_read_data_MEM[27]), 
        .sl2(n30), .d3(DM_read_data_MEM[11]), .sl3(n33) );
    and2_1 U8 ( .x(DM_read_data_CPU[31]), .a(DM_read_data_MEM[31]), .b(n29) );
    and2_1 U9 ( .x(DM_read_data_CPU[30]), .a(DM_read_data_MEM[30]), .b(n29) );
    mx4_1 U10 ( .x(DM_read_data_CPU[2]), .d0(DM_read_data_MEM[2]), .sl0(mask
        [0]), .d1(DM_read_data_MEM[18]), .sl1(n32), .d2(DM_read_data_MEM[26]), 
        .sl2(n30), .d3(DM_read_data_MEM[10]), .sl3(n33) );
    and2_1 U11 ( .x(DM_read_data_CPU[29]), .a(DM_read_data_MEM[29]), .b(n29)
         );
    and2_1 U12 ( .x(DM_read_data_CPU[28]), .a(DM_read_data_MEM[28]), .b(n29)
         );
    and2_1 U13 ( .x(DM_read_data_CPU[27]), .a(DM_read_data_MEM[27]), .b(n29)
         );
    and2_1 U14 ( .x(DM_read_data_CPU[26]), .a(DM_read_data_MEM[26]), .b(n29)
         );
    and2_1 U15 ( .x(DM_read_data_CPU[25]), .a(DM_read_data_MEM[25]), .b(n29)
         );
    and2_1 U16 ( .x(DM_read_data_CPU[24]), .a(DM_read_data_MEM[24]), .b(n29)
         );
    and2_1 U17 ( .x(DM_read_data_CPU[23]), .a(DM_read_data_MEM[23]), .b(n29)
         );
    and2_1 U18 ( .x(DM_read_data_CPU[22]), .a(DM_read_data_MEM[22]), .b(n29)
         );
    and2_1 U19 ( .x(DM_read_data_CPU[21]), .a(DM_read_data_MEM[21]), .b(n29)
         );
    and2_1 U20 ( .x(DM_read_data_CPU[20]), .a(DM_read_data_MEM[20]), .b(n29)
         );
    mx4_1 U21 ( .x(DM_read_data_CPU[1]), .d0(DM_read_data_MEM[1]), .sl0(mask
        [0]), .d1(DM_read_data_MEM[17]), .sl1(n32), .d2(DM_read_data_MEM[25]), 
        .sl2(n30), .d3(DM_read_data_MEM[9]), .sl3(n33) );
    and2_1 U22 ( .x(DM_read_data_CPU[19]), .a(DM_read_data_MEM[19]), .b(n29)
         );
    and2_1 U23 ( .x(DM_read_data_CPU[18]), .a(DM_read_data_MEM[18]), .b(n29)
         );
    and2_1 U24 ( .x(DM_read_data_CPU[17]), .a(DM_read_data_MEM[17]), .b(n29)
         );
    and2_1 U25 ( .x(DM_read_data_CPU[16]), .a(DM_read_data_MEM[16]), .b(n29)
         );
    mx4_1 U26 ( .x(DM_read_data_CPU[0]), .d0(DM_read_data_MEM[0]), .sl0(mask
        [0]), .d1(DM_read_data_MEM[16]), .sl1(n32), .d2(DM_read_data_MEM[24]), 
        .sl2(n30), .d3(DM_read_data_MEM[8]), .sl3(n33) );
    inv_2 U27 ( .x(n60), .a(DM_read_data_MEM[8]) );
    inv_2 U28 ( .x(n58), .a(DM_read_data_MEM[9]) );
    inv_2 U29 ( .x(n72), .a(DM_read_data_MEM[10]) );
    inv_2 U30 ( .x(n70), .a(DM_read_data_MEM[11]) );
    inv_2 U31 ( .x(n68), .a(DM_read_data_MEM[12]) );
    inv_2 U32 ( .x(n66), .a(DM_read_data_MEM[13]) );
    inv_2 U33 ( .x(n64), .a(DM_read_data_MEM[14]) );
    inv_2 U34 ( .x(n62), .a(DM_read_data_MEM[15]) );
    inv_2 U35 ( .x(n59), .a(DM_read_data_MEM[24]) );
    inv_2 U36 ( .x(n57), .a(DM_read_data_MEM[25]) );
    inv_2 U37 ( .x(n71), .a(DM_read_data_MEM[26]) );
    inv_2 U38 ( .x(n69), .a(DM_read_data_MEM[27]) );
    inv_2 U39 ( .x(n67), .a(DM_read_data_MEM[28]) );
    inv_2 U40 ( .x(n65), .a(DM_read_data_MEM[29]) );
    inv_2 U41 ( .x(n63), .a(DM_read_data_MEM[30]) );
    inv_2 U42 ( .x(n61), .a(DM_read_data_MEM[31]) );
    nand3_1 U43 ( .x(n34), .a(n39), .b(n40), .c(\byte ) );
    oai31_2 U44 ( .x(n32), .a(n75), .b(DM_addr_CPU[1]), .c(n39), .d(n36) );
    nand2_2 U45 ( .x(n36), .a(n76), .b(n40) );
    nand2_2 U46 ( .x(n74), .a(word), .b(n75) );
    nand2_2 U47 ( .x(n35), .a(n73), .b(n75) );
    inv_2 U48 ( .x(n73), .a(word) );
    inv_2 U49 ( .x(n76), .a(n74) );
    nand3_1 U50 ( .x(n38), .a(\byte ), .b(n39), .c(DM_addr_CPU[1]) );
    inv_2 U51 ( .x(n33), .a(n38) );
    inv_2 U52 ( .x(n75), .a(\byte ) );
    oai21_1 U53 ( .x(mask[0]), .a(n39), .b(n40), .c(n28) );
    inv_2 U54 ( .x(n39), .a(DM_addr_CPU[0]) );
    inv_2 U55 ( .x(n40), .a(DM_addr_CPU[1]) );
    nand2_2 U56 ( .x(mask[1]), .a(n28), .b(n38) );
    nand2_2 U57 ( .x(mask[2]), .a(n37), .b(n35) );
    inv_2 U58 ( .x(n37), .a(n32) );
    nand3_1 U59 ( .x(mask[3]), .a(n34), .b(n35), .c(n36) );
    ao222_1 U60 ( .x(DM_write_data_MEM[31]), .a(n29), .b(DM_write_data_CPU[31]
        ), .c(n30), .d(DM_write_data_CPU[7]), .e(DM_write_data_CPU[15]), .f(
        n31) );
    ao222_1 U61 ( .x(DM_write_data_MEM[30]), .a(DM_write_data_CPU[30]), .b(n29
        ), .c(n30), .d(DM_write_data_CPU[6]), .e(DM_write_data_CPU[14]), .f(
        n31) );
    ao222_1 U62 ( .x(DM_write_data_MEM[29]), .a(DM_write_data_CPU[29]), .b(n29
        ), .c(n30), .d(DM_write_data_CPU[5]), .e(DM_write_data_CPU[13]), .f(
        n31) );
    ao222_1 U63 ( .x(DM_write_data_MEM[28]), .a(DM_write_data_CPU[28]), .b(n29
        ), .c(n30), .d(DM_write_data_CPU[4]), .e(DM_write_data_CPU[12]), .f(
        n31) );
    ao222_1 U64 ( .x(DM_write_data_MEM[27]), .a(DM_write_data_CPU[27]), .b(n29
        ), .c(DM_write_data_CPU[3]), .d(n30), .e(DM_write_data_CPU[11]), .f(
        n31) );
    ao222_1 U65 ( .x(DM_write_data_MEM[26]), .a(DM_write_data_CPU[26]), .b(n29
        ), .c(DM_write_data_CPU[2]), .d(n30), .e(DM_write_data_CPU[10]), .f(
        n31) );
    ao222_1 U66 ( .x(DM_write_data_MEM[25]), .a(DM_write_data_CPU[25]), .b(n29
        ), .c(n30), .d(DM_write_data_CPU[1]), .e(n31), .f(DM_write_data_CPU[9]
        ) );
    ao222_1 U67 ( .x(DM_write_data_MEM[24]), .a(DM_write_data_CPU[24]), .b(n29
        ), .c(n30), .d(DM_write_data_CPU[0]), .e(n31), .f(DM_write_data_CPU[8]
        ) );
    inv_2 U68 ( .x(n30), .a(n34) );
    inv_2 U69 ( .x(n31), .a(n36) );
    ao22_1 U70 ( .x(DM_write_data_MEM[23]), .a(DM_write_data_CPU[23]), .b(n29), 
        .c(DM_write_data_CPU[7]), .d(n32) );
    ao22_1 U71 ( .x(DM_write_data_MEM[22]), .a(DM_write_data_CPU[22]), .b(n29), 
        .c(DM_write_data_CPU[6]), .d(n32) );
    ao22_1 U72 ( .x(DM_write_data_MEM[21]), .a(DM_write_data_CPU[21]), .b(n29), 
        .c(DM_write_data_CPU[5]), .d(n32) );
    ao22_1 U73 ( .x(DM_write_data_MEM[20]), .a(DM_write_data_CPU[20]), .b(n29), 
        .c(DM_write_data_CPU[4]), .d(n32) );
    ao22_1 U74 ( .x(DM_write_data_MEM[19]), .a(DM_write_data_CPU[19]), .b(n29), 
        .c(DM_write_data_CPU[3]), .d(n32) );
    ao22_1 U75 ( .x(DM_write_data_MEM[18]), .a(DM_write_data_CPU[18]), .b(n29), 
        .c(DM_write_data_CPU[2]), .d(n32) );
    ao22_1 U76 ( .x(DM_write_data_MEM[17]), .a(DM_write_data_CPU[17]), .b(n29), 
        .c(DM_write_data_CPU[1]), .d(n32) );
    ao22_1 U77 ( .x(DM_write_data_MEM[16]), .a(DM_write_data_CPU[16]), .b(n29), 
        .c(DM_write_data_CPU[0]), .d(n32) );
    inv_2 U78 ( .x(n29), .a(n35) );
    inv_2 U79 ( .x(n46), .a(DM_write_data_CPU[15]) );
    inv_2 U80 ( .x(n48), .a(DM_write_data_CPU[14]) );
    inv_2 U81 ( .x(n50), .a(DM_write_data_CPU[13]) );
    inv_2 U82 ( .x(n52), .a(DM_write_data_CPU[12]) );
    inv_2 U83 ( .x(n54), .a(DM_write_data_CPU[11]) );
    inv_2 U84 ( .x(n56), .a(DM_write_data_CPU[10]) );
    inv_2 U85 ( .x(n42), .a(DM_write_data_CPU[9]) );
    inv_2 U86 ( .x(n44), .a(DM_write_data_CPU[8]) );
    and2_1 U87 ( .x(DM_write_data_MEM[7]), .a(DM_write_data_CPU[7]), .b(mask
        [0]) );
    inv_2 U88 ( .x(n45), .a(DM_write_data_CPU[7]) );
    and2_1 U89 ( .x(DM_write_data_MEM[6]), .a(DM_write_data_CPU[6]), .b(mask
        [0]) );
    inv_2 U90 ( .x(n47), .a(DM_write_data_CPU[6]) );
    and2_1 U91 ( .x(DM_write_data_MEM[5]), .a(DM_write_data_CPU[5]), .b(mask
        [0]) );
    inv_2 U92 ( .x(n49), .a(DM_write_data_CPU[5]) );
    and2_1 U93 ( .x(DM_write_data_MEM[4]), .a(DM_write_data_CPU[4]), .b(mask
        [0]) );
    inv_2 U94 ( .x(n51), .a(DM_write_data_CPU[4]) );
    and2_1 U95 ( .x(DM_write_data_MEM[3]), .a(DM_write_data_CPU[3]), .b(mask
        [0]) );
    inv_2 U96 ( .x(n53), .a(DM_write_data_CPU[3]) );
    and2_1 U97 ( .x(DM_write_data_MEM[2]), .a(DM_write_data_CPU[2]), .b(mask
        [0]) );
    inv_2 U98 ( .x(n55), .a(DM_write_data_CPU[2]) );
    and2_1 U99 ( .x(DM_write_data_MEM[1]), .a(DM_write_data_CPU[1]), .b(mask
        [0]) );
    inv_2 U100 ( .x(n41), .a(DM_write_data_CPU[1]) );
    and2_1 U101 ( .x(DM_write_data_MEM[0]), .a(DM_write_data_CPU[0]), .b(mask
        [0]) );
    inv_2 U102 ( .x(n43), .a(DM_write_data_CPU[0]) );
    oai22_1 U103 ( .x(DM_write_data_MEM[15]), .a(n38), .b(n45), .c(n28), .d(
        n46) );
    oai22_1 U104 ( .x(DM_write_data_MEM[14]), .a(n38), .b(n47), .c(n28), .d(
        n48) );
    oai22_1 U105 ( .x(DM_write_data_MEM[13]), .a(n38), .b(n49), .c(n28), .d(
        n50) );
    oai22_1 U106 ( .x(DM_write_data_MEM[12]), .a(n38), .b(n51), .c(n28), .d(
        n52) );
    oai22_1 U107 ( .x(DM_write_data_MEM[11]), .a(n38), .b(n53), .c(n28), .d(
        n54) );
    oai22_1 U108 ( .x(DM_write_data_MEM[10]), .a(n38), .b(n55), .c(n28), .d(
        n56) );
    oai22_1 U109 ( .x(DM_write_data_MEM[9]), .a(n38), .b(n41), .c(n28), .d(n42
        ) );
    oai22_1 U110 ( .x(DM_write_data_MEM[8]), .a(n38), .b(n43), .c(n28), .d(n44
        ) );
    oai22_1 U111 ( .x(DM_read_data_CPU[15]), .a(n36), .b(n61), .c(n28), .d(n62
        ) );
    oai22_1 U112 ( .x(DM_read_data_CPU[14]), .a(n36), .b(n63), .c(n28), .d(n64
        ) );
    oai22_1 U113 ( .x(DM_read_data_CPU[13]), .a(n36), .b(n65), .c(n28), .d(n66
        ) );
    oai22_1 U114 ( .x(DM_read_data_CPU[12]), .a(n36), .b(n67), .c(n28), .d(n68
        ) );
    oai22_1 U115 ( .x(DM_read_data_CPU[11]), .a(n36), .b(n69), .c(n28), .d(n70
        ) );
    oai22_1 U116 ( .x(DM_read_data_CPU[10]), .a(n36), .b(n71), .c(n28), .d(n72
        ) );
    oai22_1 U117 ( .x(DM_read_data_CPU[9]), .a(n36), .b(n57), .c(n28), .d(n58)
         );
    oai22_1 U118 ( .x(DM_read_data_CPU[8]), .a(n36), .b(n59), .c(n28), .d(n60)
         );
    oa21_2 U119 ( .x(n28), .a(n74), .b(n40), .c(n35) );
endmodule


module mem_load ( start, scan_in, scan_out, scan_clk, data_out, data_in, 
    data_write, read, addr_out );
output [31:0] data_out;
input  [31:0] data_in;
output [10:0] addr_out;
input  start, scan_in, scan_clk, read;
output scan_out, data_write;
    wire shifter_43, shifter_42, shifter_41, shifter_40, shifter_39, 
        shifter_38, shifter_37, shifter_36, shifter_35, shifter_34, shifter_33, 
        shifter_32, shifter_31, shifter_30, shifter_29, shifter_28, shifter_27, 
        shifter_26, shifter_25, shifter_24, shifter_23, shifter_22, shifter_21, 
        shifter_20, shifter_19, shifter_18, shifter_17, shifter_16, shifter_15, 
        shifter_14, shifter_13, shifter_12, shifter_11, shifter_10, shifter_9, 
        shifter_8, shifter_7, shifter_6, shifter_5, shifter_4, shifter_3, 
        shifter_2, shifter_1, rw, unload_1, unload_0, N26, N28, N30, N32, N34, 
        N36, N38, N40, N42, N44, N46, N48, N50, N52, N54, N56, N58, N60, N62, 
        N64, N66, N68, N70, N72, N74, N76, N78, N80, N82, N84, N86, N88, N112, 
        N206, N90, N92, N94, N96, N98, N100, N102, N104, N106, N108, N110, 
        N116, N118, N111, N117, N139, N205, n5, n6, n7, n8, n9, n10, n11, n12, 
        n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, 
        n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, 
        n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, 
        n55, n56, n57, n58, n59, n60, n61, n62;
    and3i_1 U3 ( .x(n61), .a(unload_0), .b(n54), .c(n55) );
    oa21_2 U4 ( .x(N139), .a(n46), .b(n47), .c(n48) );
    nand2_2 U5 ( .x(n58), .a(scan_out), .b(n57) );
    nand3_1 U6 ( .x(n56), .a(scan_out), .b(rw), .c(n61) );
    oai21_1 U7 ( .x(N116), .a(n52), .b(n54), .c(n45) );
    nand3_1 U8 ( .x(N117), .a(n43), .b(n44), .c(n45) );
    nand2_2 U9 ( .x(n43), .a(n58), .b(n59) );
    oai21_1 U10 ( .x(N118), .a(n52), .b(n53), .c(n45) );
    and2_1 U11 ( .x(N90), .a(shifter_33), .b(n50) );
    and2_1 U12 ( .x(N92), .a(shifter_34), .b(n62) );
    and2_1 U13 ( .x(N94), .a(shifter_35), .b(n50) );
    and2_1 U14 ( .x(N96), .a(shifter_36), .b(n62) );
    and2_1 U15 ( .x(N98), .a(n62), .b(shifter_37) );
    and2_1 U16 ( .x(N100), .a(shifter_38), .b(n50) );
    and2_1 U17 ( .x(N102), .a(shifter_39), .b(n62) );
    and2_1 U18 ( .x(N104), .a(shifter_40), .b(n50) );
    and2_1 U19 ( .x(N106), .a(shifter_41), .b(n62) );
    and2_1 U20 ( .x(N108), .a(shifter_42), .b(n50) );
    and2_1 U21 ( .x(N110), .a(shifter_43), .b(n62) );
    oa21_2 U22 ( .x(n49), .a(n46), .b(n43), .c(n48) );
    inv_2 U23 ( .x(n46), .a(n56) );
    inv_2 U24 ( .x(n51), .a(n45) );
    ao21_1 U25 ( .x(N112), .a(scan_in), .b(n50), .c(start) );
    inv_2 U26 ( .x(n50), .a(n52) );
    nand2_2 U27 ( .x(n52), .a(n44), .b(n60) );
    inv_2 U28 ( .x(n60), .a(n43) );
    inv_2 U29 ( .x(n62), .a(n52) );
    oai21_1 U30 ( .x(N205), .a(n40), .b(n41), .c(n42) );
    inv_2 U31 ( .x(n40), .a(n59) );
    nand3_1 U32 ( .x(n59), .a(n54), .b(n53), .c(unload_1) );
    nand2_2 U33 ( .x(n41), .a(n48), .b(n56) );
    inv_2 U34 ( .x(n48), .a(start) );
    inv_2 U35 ( .x(n47), .a(n58) );
    inv_2 U36 ( .x(n44), .a(n41) );
    dffph_2 data_out_reg_0 ( .q(data_out[0]), .d(shifter_1), .ck(scan_clk), 
        .g(N206) );
    dffph_2 data_out_reg_1 ( .q(data_out[1]), .d(shifter_2), .ck(scan_clk), 
        .g(N206) );
    dffph_2 data_out_reg_2 ( .q(data_out[2]), .d(shifter_3), .ck(scan_clk), 
        .g(N206) );
    dffph_2 data_out_reg_3 ( .q(data_out[3]), .d(shifter_4), .ck(scan_clk), 
        .g(N206) );
    dffph_2 data_out_reg_4 ( .q(data_out[4]), .d(shifter_5), .ck(scan_clk), 
        .g(N206) );
    dffph_2 data_out_reg_5 ( .q(data_out[5]), .d(shifter_6), .ck(scan_clk), 
        .g(N206) );
    dffph_2 data_out_reg_6 ( .q(data_out[6]), .d(shifter_7), .ck(scan_clk), 
        .g(N206) );
    dffph_2 data_out_reg_7 ( .q(data_out[7]), .d(shifter_8), .ck(scan_clk), 
        .g(N206) );
    dffph_2 data_out_reg_8 ( .q(data_out[8]), .d(shifter_9), .ck(scan_clk), 
        .g(N206) );
    dffph_2 data_out_reg_9 ( .q(data_out[9]), .d(shifter_10), .ck(scan_clk), 
        .g(N206) );
    dffph_2 data_out_reg_10 ( .q(data_out[10]), .d(shifter_11), .ck(scan_clk), 
        .g(N206) );
    dffph_2 data_out_reg_11 ( .q(data_out[11]), .d(shifter_12), .ck(scan_clk), 
        .g(N206) );
    dffph_2 data_out_reg_12 ( .q(data_out[12]), .d(shifter_13), .ck(scan_clk), 
        .g(N206) );
    dffph_2 data_out_reg_13 ( .q(data_out[13]), .d(shifter_14), .ck(scan_clk), 
        .g(N206) );
    dffph_2 data_out_reg_14 ( .q(data_out[14]), .d(shifter_15), .ck(scan_clk), 
        .g(N206) );
    dffph_2 data_out_reg_15 ( .q(data_out[15]), .d(shifter_16), .ck(scan_clk), 
        .g(n38) );
    dffph_2 data_out_reg_16 ( .q(data_out[16]), .d(shifter_17), .ck(scan_clk), 
        .g(N206) );
    dffph_2 data_out_reg_17 ( .q(data_out[17]), .d(shifter_18), .ck(scan_clk), 
        .g(N206) );
    dffph_2 data_out_reg_18 ( .q(data_out[18]), .d(shifter_19), .ck(scan_clk), 
        .g(N206) );
    dffph_2 data_out_reg_19 ( .q(data_out[19]), .d(shifter_20), .ck(scan_clk), 
        .g(N206) );
    dffph_2 data_out_reg_20 ( .q(data_out[20]), .d(shifter_21), .ck(scan_clk), 
        .g(N206) );
    dffph_2 data_out_reg_21 ( .q(data_out[21]), .d(shifter_22), .ck(scan_clk), 
        .g(N206) );
    dffph_2 data_out_reg_22 ( .q(data_out[22]), .d(shifter_23), .ck(scan_clk), 
        .g(N206) );
    dffph_2 data_out_reg_23 ( .q(data_out[23]), .d(shifter_24), .ck(scan_clk), 
        .g(N206) );
    dffph_2 data_out_reg_24 ( .q(data_out[24]), .d(shifter_25), .ck(scan_clk), 
        .g(N206) );
    dffph_2 data_out_reg_25 ( .q(data_out[25]), .d(shifter_26), .ck(scan_clk), 
        .g(N206) );
    dffph_2 data_out_reg_26 ( .q(data_out[26]), .d(shifter_27), .ck(scan_clk), 
        .g(N206) );
    dffph_2 data_out_reg_27 ( .q(data_out[27]), .d(shifter_28), .ck(scan_clk), 
        .g(N206) );
    dffph_2 data_out_reg_28 ( .q(data_out[28]), .d(shifter_29), .ck(scan_clk), 
        .g(N206) );
    dffph_2 data_out_reg_29 ( .q(data_out[29]), .d(shifter_30), .ck(scan_clk), 
        .g(N206) );
    dffph_2 data_out_reg_30 ( .q(data_out[30]), .d(shifter_31), .ck(scan_clk), 
        .g(N206) );
    dffph_2 data_out_reg_31 ( .q(data_out[31]), .d(shifter_32), .ck(scan_clk), 
        .g(N206) );
    dffph_2 addr_out_reg_0 ( .q(addr_out[0]), .d(shifter_33), .ck(scan_clk), 
        .g(N139) );
    dffph_2 addr_out_reg_1 ( .q(addr_out[1]), .d(shifter_34), .ck(scan_clk), 
        .g(N139) );
    dffph_2 addr_out_reg_2 ( .q(addr_out[2]), .d(shifter_35), .ck(scan_clk), 
        .g(N139) );
    dffph_2 addr_out_reg_3 ( .q(addr_out[3]), .d(shifter_36), .ck(scan_clk), 
        .g(N139) );
    dffph_2 addr_out_reg_4 ( .q(addr_out[4]), .d(shifter_37), .ck(scan_clk), 
        .g(N139) );
    dffph_2 addr_out_reg_5 ( .q(addr_out[5]), .d(shifter_38), .ck(scan_clk), 
        .g(N139) );
    dffph_2 addr_out_reg_6 ( .q(addr_out[6]), .d(shifter_39), .ck(scan_clk), 
        .g(N139) );
    dffph_2 addr_out_reg_7 ( .q(addr_out[7]), .d(shifter_40), .ck(scan_clk), 
        .g(N139) );
    dffph_2 addr_out_reg_8 ( .q(addr_out[8]), .d(shifter_41), .ck(scan_clk), 
        .g(N139) );
    dffph_2 addr_out_reg_9 ( .q(addr_out[9]), .d(shifter_42), .ck(scan_clk), 
        .g(N139) );
    dffph_2 addr_out_reg_10 ( .q(addr_out[10]), .d(shifter_43), .ck(scan_clk), 
        .g(N139) );
    dffph_2 unload_reg_0 ( .q(unload_0), .qb(n53), .d(n5), .ck(scan_clk), .g(
        N117) );
    dffph_2 unload_reg_1 ( .q(unload_1), .qb(n55), .d(N116), .ck(scan_clk), 
        .g(N117) );
    dffph_2 unload_reg_2 ( .qb(n54), .d(N118), .ck(scan_clk), .g(N117) );
    dffph_2 shifter_reg_0 ( .q(scan_out), .d(N26), .ck(scan_clk), .g(n39) );
    dffph_2 shifter_reg_1 ( .q(shifter_1), .d(N28), .ck(scan_clk), .g(n39) );
    dffph_2 shifter_reg_2 ( .q(shifter_2), .d(N30), .ck(scan_clk), .g(n39) );
    dffph_2 shifter_reg_3 ( .q(shifter_3), .d(N32), .ck(scan_clk), .g(n39) );
    dffph_2 shifter_reg_4 ( .q(shifter_4), .d(N34), .ck(scan_clk), .g(n39) );
    dffph_2 shifter_reg_5 ( .q(shifter_5), .d(N36), .ck(scan_clk), .g(n39) );
    dffph_2 shifter_reg_6 ( .q(shifter_6), .d(N38), .ck(scan_clk), .g(n39) );
    dffph_2 shifter_reg_7 ( .q(shifter_7), .d(N40), .ck(scan_clk), .g(N111) );
    dffph_2 shifter_reg_8 ( .q(shifter_8), .d(N42), .ck(scan_clk), .g(N111) );
    dffph_2 shifter_reg_9 ( .q(shifter_9), .d(N44), .ck(scan_clk), .g(N111) );
    dffph_2 shifter_reg_10 ( .q(shifter_10), .d(N46), .ck(scan_clk), .g(N111)
         );
    dffph_2 shifter_reg_11 ( .q(shifter_11), .d(N48), .ck(scan_clk), .g(N111)
         );
    dffph_2 shifter_reg_12 ( .q(shifter_12), .d(N50), .ck(scan_clk), .g(N111)
         );
    dffph_2 shifter_reg_13 ( .q(shifter_13), .d(N52), .ck(scan_clk), .g(N111)
         );
    dffph_2 shifter_reg_14 ( .q(shifter_14), .d(N54), .ck(scan_clk), .g(N111)
         );
    dffph_2 shifter_reg_15 ( .q(shifter_15), .d(N56), .ck(scan_clk), .g(N111)
         );
    dffph_2 shifter_reg_16 ( .q(shifter_16), .d(N58), .ck(scan_clk), .g(N111)
         );
    dffph_2 shifter_reg_17 ( .q(shifter_17), .d(N60), .ck(scan_clk), .g(N111)
         );
    dffph_2 shifter_reg_18 ( .q(shifter_18), .d(N62), .ck(scan_clk), .g(N111)
         );
    dffph_2 shifter_reg_19 ( .q(shifter_19), .d(N64), .ck(scan_clk), .g(N111)
         );
    dffph_2 shifter_reg_20 ( .q(shifter_20), .d(N66), .ck(scan_clk), .g(N111)
         );
    dffph_2 shifter_reg_21 ( .q(shifter_21), .d(N68), .ck(scan_clk), .g(N111)
         );
    dffph_2 shifter_reg_22 ( .q(shifter_22), .d(N70), .ck(scan_clk), .g(N111)
         );
    dffph_2 shifter_reg_23 ( .q(shifter_23), .d(N72), .ck(scan_clk), .g(n39)
         );
    dffph_2 shifter_reg_24 ( .q(shifter_24), .d(N74), .ck(scan_clk), .g(N111)
         );
    dffph_2 shifter_reg_25 ( .q(shifter_25), .d(N76), .ck(scan_clk), .g(n39)
         );
    dffph_2 shifter_reg_26 ( .q(shifter_26), .d(N78), .ck(scan_clk), .g(N111)
         );
    dffph_2 shifter_reg_27 ( .q(shifter_27), .d(N80), .ck(scan_clk), .g(n39)
         );
    dffph_2 shifter_reg_28 ( .q(shifter_28), .d(N82), .ck(scan_clk), .g(N111)
         );
    dffph_2 shifter_reg_29 ( .q(shifter_29), .d(N84), .ck(scan_clk), .g(n39)
         );
    dffph_2 shifter_reg_30 ( .q(shifter_30), .d(N86), .ck(scan_clk), .g(N111)
         );
    dffph_2 shifter_reg_31 ( .q(shifter_31), .d(N88), .ck(scan_clk), .g(N111)
         );
    dffph_2 shifter_reg_32 ( .q(shifter_32), .d(N90), .ck(scan_clk), .g(N111)
         );
    dffph_2 shifter_reg_33 ( .q(shifter_33), .d(N92), .ck(scan_clk), .g(n39)
         );
    dffph_2 shifter_reg_34 ( .q(shifter_34), .d(N94), .ck(scan_clk), .g(N111)
         );
    dffph_2 shifter_reg_35 ( .q(shifter_35), .d(N96), .ck(scan_clk), .g(N111)
         );
    dffph_2 shifter_reg_36 ( .q(shifter_36), .d(N98), .ck(scan_clk), .g(N111)
         );
    dffph_2 shifter_reg_37 ( .q(shifter_37), .d(N100), .ck(scan_clk), .g(n39)
         );
    dffph_2 shifter_reg_38 ( .q(shifter_38), .d(N102), .ck(scan_clk), .g(N111)
         );
    dffph_2 shifter_reg_39 ( .q(shifter_39), .d(N104), .ck(scan_clk), .g(N111)
         );
    dffph_2 shifter_reg_40 ( .q(shifter_40), .d(N106), .ck(scan_clk), .g(N111)
         );
    dffph_2 shifter_reg_41 ( .q(shifter_41), .d(N108), .ck(scan_clk), .g(n39)
         );
    dffph_2 shifter_reg_42 ( .q(shifter_42), .d(N110), .ck(scan_clk), .g(N111)
         );
    dffph_2 shifter_reg_43 ( .q(shifter_43), .d(N112), .ck(scan_clk), .g(N111)
         );
    dffph_2 rw_reg ( .q(rw), .qb(n57), .d(read), .ck(scan_clk), .g(start) );
    dffph_2 data_write_reg ( .q(data_write), .d(N206), .ck(scan_clk), .g(N205)
         );
    oai221_1 U37 ( .x(n5), .a(n55), .b(n52), .c(start), .d(n56), .e(n45) );
    and2_1 U38 ( .x(n6), .a(shifter_32), .b(n62) );
    and2_1 U39 ( .x(n7), .a(shifter_31), .b(n50) );
    and2_1 U40 ( .x(n8), .a(shifter_30), .b(n62) );
    and2_1 U41 ( .x(n9), .a(shifter_29), .b(n50) );
    and2_1 U42 ( .x(n10), .a(shifter_28), .b(n62) );
    and2_1 U43 ( .x(n11), .a(shifter_27), .b(n50) );
    and2_1 U44 ( .x(n12), .a(shifter_26), .b(n62) );
    and2_1 U45 ( .x(n13), .a(shifter_25), .b(n50) );
    and2_1 U46 ( .x(n14), .a(shifter_24), .b(n62) );
    and2_1 U47 ( .x(n15), .a(shifter_23), .b(n50) );
    and2_1 U48 ( .x(n16), .a(shifter_22), .b(n62) );
    and2_1 U49 ( .x(n17), .a(shifter_21), .b(n50) );
    and2_1 U50 ( .x(n18), .a(shifter_20), .b(n62) );
    and2_1 U51 ( .x(n19), .a(shifter_19), .b(n50) );
    and2_1 U52 ( .x(n20), .a(shifter_18), .b(n62) );
    and2_1 U53 ( .x(n21), .a(shifter_17), .b(n50) );
    and2_1 U54 ( .x(n22), .a(shifter_16), .b(n62) );
    and2_1 U55 ( .x(n23), .a(shifter_15), .b(n50) );
    and2_1 U56 ( .x(n24), .a(shifter_14), .b(n62) );
    and2_1 U57 ( .x(n25), .a(shifter_13), .b(n50) );
    and2_1 U58 ( .x(n26), .a(shifter_12), .b(n62) );
    and2_1 U59 ( .x(n27), .a(shifter_11), .b(n50) );
    and2_1 U60 ( .x(n28), .a(shifter_10), .b(n62) );
    and2_1 U61 ( .x(n29), .a(shifter_9), .b(n50) );
    and2_1 U62 ( .x(n30), .a(shifter_8), .b(n62) );
    and2_1 U63 ( .x(n31), .a(shifter_7), .b(n50) );
    and2_1 U64 ( .x(n32), .a(shifter_6), .b(n62) );
    and2_1 U65 ( .x(n33), .a(shifter_5), .b(n50) );
    and2_1 U66 ( .x(n34), .a(shifter_4), .b(n62) );
    and2_1 U67 ( .x(n35), .a(shifter_3), .b(n50) );
    and2_1 U68 ( .x(n36), .a(shifter_2), .b(n62) );
    and2_1 U69 ( .x(n37), .a(shifter_1), .b(n50) );
    inv_0 U70 ( .x(n38), .a(n42) );
    inv_2 U71 ( .x(N206), .a(n42) );
    nand2_2 U72 ( .x(n42), .a(n47), .b(n44) );
    buf_1 U73 ( .x(n39), .a(N111) );
    nand2_2 U74 ( .x(N111), .a(n49), .b(n45) );
    nand3_1 U75 ( .x(n45), .a(n40), .b(n58), .c(n44) );
    oa22_4 U76 ( .x(N88), .a(data_in[31]), .b(n6), .c(n6), .d(n51) );
    oa22_4 U77 ( .x(N86), .a(n7), .b(n51), .c(data_in[30]), .d(n7) );
    oa22_4 U78 ( .x(N84), .a(n8), .b(n51), .c(data_in[29]), .d(n8) );
    oa22_4 U79 ( .x(N82), .a(n9), .b(n51), .c(data_in[28]), .d(n9) );
    oa22_4 U80 ( .x(N80), .a(n10), .b(n51), .c(data_in[27]), .d(n10) );
    oa22_4 U81 ( .x(N78), .a(n11), .b(n51), .c(data_in[26]), .d(n11) );
    oa22_4 U82 ( .x(N76), .a(n12), .b(n51), .c(data_in[25]), .d(n12) );
    oa22_4 U83 ( .x(N74), .a(n13), .b(n51), .c(data_in[24]), .d(n13) );
    oa22_4 U84 ( .x(N72), .a(n14), .b(n51), .c(data_in[23]), .d(n14) );
    oa22_4 U85 ( .x(N70), .a(n15), .b(n51), .c(data_in[22]), .d(n15) );
    oa22_4 U86 ( .x(N68), .a(n16), .b(n51), .c(data_in[21]), .d(n16) );
    oa22_4 U87 ( .x(N66), .a(n17), .b(n51), .c(data_in[20]), .d(n17) );
    oa22_4 U88 ( .x(N64), .a(n18), .b(n51), .c(data_in[19]), .d(n18) );
    oa22_4 U89 ( .x(N62), .a(n19), .b(n51), .c(data_in[18]), .d(n19) );
    oa22_4 U90 ( .x(N60), .a(n20), .b(n51), .c(data_in[17]), .d(n20) );
    oa22_4 U91 ( .x(N58), .a(n21), .b(n51), .c(data_in[16]), .d(n21) );
    oa22_4 U92 ( .x(N56), .a(n22), .b(n51), .c(data_in[15]), .d(n22) );
    oa22_4 U93 ( .x(N54), .a(n23), .b(n51), .c(data_in[14]), .d(n23) );
    oa22_4 U94 ( .x(N52), .a(n24), .b(n51), .c(data_in[13]), .d(n24) );
    oa22_4 U95 ( .x(N50), .a(n25), .b(n51), .c(data_in[12]), .d(n25) );
    oa22_4 U96 ( .x(N48), .a(n26), .b(n51), .c(data_in[11]), .d(n26) );
    oa22_4 U97 ( .x(N46), .a(n27), .b(n51), .c(data_in[10]), .d(n27) );
    oa22_4 U98 ( .x(N44), .a(n28), .b(n51), .c(data_in[9]), .d(n28) );
    oa22_4 U99 ( .x(N42), .a(n29), .b(n51), .c(data_in[8]), .d(n29) );
    oa22_4 U100 ( .x(N40), .a(n30), .b(n51), .c(data_in[7]), .d(n30) );
    oa22_4 U101 ( .x(N38), .a(n31), .b(n51), .c(data_in[6]), .d(n31) );
    oa22_4 U102 ( .x(N36), .a(n32), .b(n51), .c(data_in[5]), .d(n32) );
    oa22_4 U103 ( .x(N34), .a(n33), .b(n51), .c(data_in[4]), .d(n33) );
    oa22_4 U104 ( .x(N32), .a(n34), .b(n51), .c(data_in[3]), .d(n34) );
    oa22_4 U105 ( .x(N30), .a(n35), .b(n51), .c(data_in[2]), .d(n35) );
    oa22_4 U106 ( .x(N28), .a(n36), .b(n51), .c(data_in[1]), .d(n36) );
    oa22_4 U107 ( .x(N26), .a(n37), .b(n51), .c(data_in[0]), .d(n37) );
endmodule


module matched_delay_m2cp_com_iport ( x, a );
input  a;
output x;
    wire n2;
    buf_1 I1 ( .x(n2), .a(a) );
    buf_16 U1 ( .x(x), .a(n2) );
endmodule


module sr2dr_word_1 ( i, req, h, l );
input  [31:0] i;
output [31:0] h;
output [31:0] l;
input  req;
    wire \U31/ni , \U31/nh , \U31/nl , n9, n1, n2, \U30/ni , \U30/nh , 
        \U30/nl , n8, \U29/ni , \U29/nh , \U29/nl , \U28/ni , \U28/nh , 
        \U28/nl , \U27/ni , \U27/nh , \U27/nl , \U26/ni , \U26/nh , \U26/nl , 
        n7, n4, \U25/ni , \U25/nh , \U25/nl , \U24/ni , \U24/nh , \U24/nl , 
        \U23/ni , \U23/nh , \U23/nl , n3, \U22/ni , \U22/nh , \U22/nl , n6, 
        \U21/ni , \U21/nh , \U21/nl , \U20/ni , \U20/nh , \U20/nl , n5, 
        \U19/ni , \U19/nh , \U19/nl , \U18/ni , \U18/nh , \U18/nl , \U17/ni , 
        \U17/nh , \U17/nl , \U16/ni , \U16/nh , \U16/nl , \U15/ni , \U15/nh , 
        \U15/nl , \U14/ni , \U14/nh , \U14/nl , \U13/ni , \U13/nh , \U13/nl , 
        \U12/ni , \U12/nh , \U12/nl , \U11/ni , \U11/nh , \U11/nl , \U10/ni , 
        \U10/nh , \U10/nl , \U9/ni , \U9/nh , \U9/nl , \U8/ni , \U8/nh , 
        \U8/nl , \U7/ni , \U7/nh , \U7/nl , \U6/ni , \U6/nh , \U6/nl , \U5/ni , 
        \U5/nh , \U5/nl , \U4/ni , \U4/nh , \U4/nl , \U3/ni , \U3/nh , \U3/nl , 
        \U2/ni , \U2/nh , \U2/nl , \U1/ni , \U1/nh , \U1/nl , \U0/ni , \U0/nh , 
        \U0/nl , n12, n11, n10;
    inv_1 \U31/Uii  ( .x(\U31/ni ), .a(i[31]) );
    inv_1 \U31/Uih  ( .x(\U31/nh ), .a(h[31]) );
    inv_1 \U31/Uil  ( .x(\U31/nl ), .a(l[31]) );
    ao23_1 \U31/Ucl/U1/U1  ( .x(l[31]), .a(n9), .b(l[31]), .c(n1), .d(\U31/ni 
        ), .e(\U31/nh ) );
    ao23_1 \U31/Uch/U1/U1  ( .x(h[31]), .a(n9), .b(h[31]), .c(n2), .d(i[31]), 
        .e(\U31/nl ) );
    inv_1 \U30/Uii  ( .x(\U30/ni ), .a(i[30]) );
    inv_1 \U30/Uih  ( .x(\U30/nh ), .a(h[30]) );
    inv_1 \U30/Uil  ( .x(\U30/nl ), .a(l[30]) );
    ao23_1 \U30/Ucl/U1/U1  ( .x(l[30]), .a(n8), .b(l[30]), .c(n1), .d(\U30/ni 
        ), .e(\U30/nh ) );
    ao23_1 \U30/Uch/U1/U1  ( .x(h[30]), .a(n8), .b(h[30]), .c(n1), .d(i[30]), 
        .e(\U30/nl ) );
    inv_1 \U29/Uii  ( .x(\U29/ni ), .a(i[29]) );
    inv_1 \U29/Uih  ( .x(\U29/nh ), .a(h[29]) );
    inv_1 \U29/Uil  ( .x(\U29/nl ), .a(l[29]) );
    ao23_1 \U29/Ucl/U1/U1  ( .x(l[29]), .a(n8), .b(l[29]), .c(n1), .d(\U29/ni 
        ), .e(\U29/nh ) );
    ao23_1 \U29/Uch/U1/U1  ( .x(h[29]), .a(n8), .b(h[29]), .c(n2), .d(i[29]), 
        .e(\U29/nl ) );
    inv_1 \U28/Uii  ( .x(\U28/ni ), .a(i[28]) );
    inv_1 \U28/Uih  ( .x(\U28/nh ), .a(h[28]) );
    inv_1 \U28/Uil  ( .x(\U28/nl ), .a(l[28]) );
    ao23_1 \U28/Ucl/U1/U1  ( .x(l[28]), .a(n8), .b(l[28]), .c(n2), .d(\U28/ni 
        ), .e(\U28/nh ) );
    ao23_1 \U28/Uch/U1/U1  ( .x(h[28]), .a(n8), .b(h[28]), .c(n2), .d(i[28]), 
        .e(\U28/nl ) );
    inv_1 \U27/Uii  ( .x(\U27/ni ), .a(i[27]) );
    inv_1 \U27/Uih  ( .x(\U27/nh ), .a(h[27]) );
    inv_1 \U27/Uil  ( .x(\U27/nl ), .a(l[27]) );
    ao23_1 \U27/Ucl/U1/U1  ( .x(l[27]), .a(n8), .b(l[27]), .c(n2), .d(\U27/ni 
        ), .e(\U27/nh ) );
    ao23_1 \U27/Uch/U1/U1  ( .x(h[27]), .a(n8), .b(h[27]), .c(n2), .d(i[27]), 
        .e(\U27/nl ) );
    inv_1 \U26/Uii  ( .x(\U26/ni ), .a(i[26]) );
    inv_1 \U26/Uih  ( .x(\U26/nh ), .a(h[26]) );
    inv_1 \U26/Uil  ( .x(\U26/nl ), .a(l[26]) );
    ao23_1 \U26/Ucl/U1/U1  ( .x(l[26]), .a(n7), .b(l[26]), .c(n2), .d(\U26/ni 
        ), .e(\U26/nh ) );
    ao23_1 \U26/Uch/U1/U1  ( .x(h[26]), .a(n7), .b(h[26]), .c(n4), .d(i[26]), 
        .e(\U26/nl ) );
    inv_1 \U25/Uii  ( .x(\U25/ni ), .a(i[25]) );
    inv_1 \U25/Uih  ( .x(\U25/nh ), .a(h[25]) );
    inv_1 \U25/Uil  ( .x(\U25/nl ), .a(l[25]) );
    ao23_1 \U25/Ucl/U1/U1  ( .x(l[25]), .a(n7), .b(l[25]), .c(n4), .d(\U25/ni 
        ), .e(\U25/nh ) );
    ao23_1 \U25/Uch/U1/U1  ( .x(h[25]), .a(n7), .b(h[25]), .c(n4), .d(i[25]), 
        .e(\U25/nl ) );
    inv_1 \U24/Uii  ( .x(\U24/ni ), .a(i[24]) );
    inv_1 \U24/Uih  ( .x(\U24/nh ), .a(h[24]) );
    inv_1 \U24/Uil  ( .x(\U24/nl ), .a(l[24]) );
    ao23_1 \U24/Ucl/U1/U1  ( .x(l[24]), .a(n7), .b(l[24]), .c(n4), .d(\U24/ni 
        ), .e(\U24/nh ) );
    ao23_1 \U24/Uch/U1/U1  ( .x(h[24]), .a(n7), .b(h[24]), .c(n4), .d(i[24]), 
        .e(\U24/nl ) );
    inv_1 \U23/Uii  ( .x(\U23/ni ), .a(i[23]) );
    inv_1 \U23/Uih  ( .x(\U23/nh ), .a(h[23]) );
    inv_1 \U23/Uil  ( .x(\U23/nl ), .a(l[23]) );
    ao23_1 \U23/Ucl/U1/U1  ( .x(l[23]), .a(n7), .b(l[23]), .c(n3), .d(\U23/ni 
        ), .e(\U23/nh ) );
    ao23_1 \U23/Uch/U1/U1  ( .x(h[23]), .a(n7), .b(h[23]), .c(n3), .d(i[23]), 
        .e(\U23/nl ) );
    inv_1 \U22/Uii  ( .x(\U22/ni ), .a(i[22]) );
    inv_1 \U22/Uih  ( .x(\U22/nh ), .a(h[22]) );
    inv_1 \U22/Uil  ( .x(\U22/nl ), .a(l[22]) );
    ao23_1 \U22/Ucl/U1/U1  ( .x(l[22]), .a(n6), .b(l[22]), .c(n3), .d(\U22/ni 
        ), .e(\U22/nh ) );
    ao23_1 \U22/Uch/U1/U1  ( .x(h[22]), .a(n6), .b(h[22]), .c(n3), .d(i[22]), 
        .e(\U22/nl ) );
    inv_1 \U21/Uii  ( .x(\U21/ni ), .a(i[21]) );
    inv_1 \U21/Uih  ( .x(\U21/nh ), .a(h[21]) );
    inv_1 \U21/Uil  ( .x(\U21/nl ), .a(l[21]) );
    ao23_1 \U21/Ucl/U1/U1  ( .x(l[21]), .a(n6), .b(l[21]), .c(n3), .d(\U21/ni 
        ), .e(\U21/nh ) );
    ao23_1 \U21/Uch/U1/U1  ( .x(h[21]), .a(n6), .b(h[21]), .c(n3), .d(i[21]), 
        .e(\U21/nl ) );
    inv_1 \U20/Uii  ( .x(\U20/ni ), .a(i[20]) );
    inv_1 \U20/Uih  ( .x(\U20/nh ), .a(h[20]) );
    inv_1 \U20/Uil  ( .x(\U20/nl ), .a(l[20]) );
    ao23_1 \U20/Ucl/U1/U1  ( .x(l[20]), .a(n6), .b(l[20]), .c(n5), .d(\U20/ni 
        ), .e(\U20/nh ) );
    ao23_1 \U20/Uch/U1/U1  ( .x(h[20]), .a(n6), .b(h[20]), .c(n4), .d(i[20]), 
        .e(\U20/nl ) );
    inv_1 \U19/Uii  ( .x(\U19/ni ), .a(i[19]) );
    inv_1 \U19/Uih  ( .x(\U19/nh ), .a(h[19]) );
    inv_1 \U19/Uil  ( .x(\U19/nl ), .a(l[19]) );
    ao23_1 \U19/Ucl/U1/U1  ( .x(l[19]), .a(n6), .b(l[19]), .c(n4), .d(\U19/ni 
        ), .e(\U19/nh ) );
    ao23_1 \U19/Uch/U1/U1  ( .x(h[19]), .a(n6), .b(h[19]), .c(n4), .d(i[19]), 
        .e(\U19/nl ) );
    inv_1 \U18/Uii  ( .x(\U18/ni ), .a(i[18]) );
    inv_1 \U18/Uih  ( .x(\U18/nh ), .a(h[18]) );
    inv_1 \U18/Uil  ( .x(\U18/nl ), .a(l[18]) );
    ao23_1 \U18/Ucl/U1/U1  ( .x(l[18]), .a(n5), .b(l[18]), .c(n5), .d(\U18/ni 
        ), .e(\U18/nh ) );
    ao23_1 \U18/Uch/U1/U1  ( .x(h[18]), .a(n5), .b(h[18]), .c(n5), .d(i[18]), 
        .e(\U18/nl ) );
    inv_1 \U17/Uii  ( .x(\U17/ni ), .a(i[17]) );
    inv_1 \U17/Uih  ( .x(\U17/nh ), .a(h[17]) );
    inv_1 \U17/Uil  ( .x(\U17/nl ), .a(l[17]) );
    ao23_1 \U17/Ucl/U1/U1  ( .x(l[17]), .a(n6), .b(l[17]), .c(n5), .d(\U17/ni 
        ), .e(\U17/nh ) );
    ao23_1 \U17/Uch/U1/U1  ( .x(h[17]), .a(n7), .b(h[17]), .c(n4), .d(i[17]), 
        .e(\U17/nl ) );
    inv_1 \U16/Uii  ( .x(\U16/ni ), .a(i[16]) );
    inv_1 \U16/Uih  ( .x(\U16/nh ), .a(h[16]) );
    inv_1 \U16/Uil  ( .x(\U16/nl ), .a(l[16]) );
    ao23_1 \U16/Ucl/U1/U1  ( .x(l[16]), .a(n9), .b(l[16]), .c(n3), .d(\U16/ni 
        ), .e(\U16/nh ) );
    ao23_1 \U16/Uch/U1/U1  ( .x(h[16]), .a(n9), .b(h[16]), .c(n1), .d(i[16]), 
        .e(\U16/nl ) );
    inv_1 \U15/Uii  ( .x(\U15/ni ), .a(i[15]) );
    inv_1 \U15/Uih  ( .x(\U15/nh ), .a(h[15]) );
    inv_1 \U15/Uil  ( .x(\U15/nl ), .a(l[15]) );
    ao23_1 \U15/Ucl/U1/U1  ( .x(l[15]), .a(n8), .b(l[15]), .c(n1), .d(\U15/ni 
        ), .e(\U15/nh ) );
    ao23_1 \U15/Uch/U1/U1  ( .x(h[15]), .a(n7), .b(h[15]), .c(n1), .d(i[15]), 
        .e(\U15/nl ) );
    inv_1 \U14/Uii  ( .x(\U14/ni ), .a(i[14]) );
    inv_1 \U14/Uih  ( .x(\U14/nh ), .a(h[14]) );
    inv_1 \U14/Uil  ( .x(\U14/nl ), .a(l[14]) );
    ao23_1 \U14/Ucl/U1/U1  ( .x(l[14]), .a(n6), .b(l[14]), .c(n1), .d(\U14/ni 
        ), .e(\U14/nh ) );
    ao23_1 \U14/Uch/U1/U1  ( .x(h[14]), .a(n6), .b(h[14]), .c(n3), .d(i[14]), 
        .e(\U14/nl ) );
    inv_1 \U13/Uii  ( .x(\U13/ni ), .a(i[13]) );
    inv_1 \U13/Uih  ( .x(\U13/nh ), .a(h[13]) );
    inv_1 \U13/Uil  ( .x(\U13/nl ), .a(l[13]) );
    ao23_1 \U13/Ucl/U1/U1  ( .x(l[13]), .a(n6), .b(l[13]), .c(n4), .d(\U13/ni 
        ), .e(\U13/nh ) );
    ao23_1 \U13/Uch/U1/U1  ( .x(h[13]), .a(n6), .b(h[13]), .c(n4), .d(i[13]), 
        .e(\U13/nl ) );
    inv_1 \U12/Uii  ( .x(\U12/ni ), .a(i[12]) );
    inv_1 \U12/Uih  ( .x(\U12/nh ), .a(h[12]) );
    inv_1 \U12/Uil  ( .x(\U12/nl ), .a(l[12]) );
    ao23_1 \U12/Ucl/U1/U1  ( .x(l[12]), .a(n5), .b(l[12]), .c(n4), .d(\U12/ni 
        ), .e(\U12/nh ) );
    ao23_1 \U12/Uch/U1/U1  ( .x(h[12]), .a(n5), .b(h[12]), .c(n4), .d(i[12]), 
        .e(\U12/nl ) );
    inv_1 \U11/Uii  ( .x(\U11/ni ), .a(i[11]) );
    inv_1 \U11/Uih  ( .x(\U11/nh ), .a(h[11]) );
    inv_1 \U11/Uil  ( .x(\U11/nl ), .a(l[11]) );
    ao23_1 \U11/Ucl/U1/U1  ( .x(l[11]), .a(n5), .b(l[11]), .c(n4), .d(\U11/ni 
        ), .e(\U11/nh ) );
    ao23_1 \U11/Uch/U1/U1  ( .x(h[11]), .a(n5), .b(h[11]), .c(n4), .d(i[11]), 
        .e(\U11/nl ) );
    inv_1 \U10/Uii  ( .x(\U10/ni ), .a(i[10]) );
    inv_1 \U10/Uih  ( .x(\U10/nh ), .a(h[10]) );
    inv_1 \U10/Uil  ( .x(\U10/nl ), .a(l[10]) );
    ao23_1 \U10/Ucl/U1/U1  ( .x(l[10]), .a(n5), .b(l[10]), .c(n3), .d(\U10/ni 
        ), .e(\U10/nh ) );
    ao23_1 \U10/Uch/U1/U1  ( .x(h[10]), .a(n5), .b(h[10]), .c(n3), .d(i[10]), 
        .e(\U10/nl ) );
    inv_1 \U9/Uii  ( .x(\U9/ni ), .a(i[9]) );
    inv_1 \U9/Uih  ( .x(\U9/nh ), .a(h[9]) );
    inv_1 \U9/Uil  ( .x(\U9/nl ), .a(l[9]) );
    ao23_1 \U9/Ucl/U1/U1  ( .x(l[9]), .a(n5), .b(l[9]), .c(n3), .d(\U9/ni ), 
        .e(\U9/nh ) );
    ao23_1 \U9/Uch/U1/U1  ( .x(h[9]), .a(n5), .b(h[9]), .c(n3), .d(i[9]), .e(
        \U9/nl ) );
    inv_1 \U8/Uii  ( .x(\U8/ni ), .a(i[8]) );
    inv_1 \U8/Uih  ( .x(\U8/nh ), .a(h[8]) );
    inv_1 \U8/Uil  ( .x(\U8/nl ), .a(l[8]) );
    ao23_1 \U8/Ucl/U1/U1  ( .x(l[8]), .a(n5), .b(l[8]), .c(n3), .d(\U8/ni ), 
        .e(\U8/nh ) );
    ao23_1 \U8/Uch/U1/U1  ( .x(h[8]), .a(n5), .b(h[8]), .c(n3), .d(i[8]), .e(
        \U8/nl ) );
    inv_1 \U7/Uii  ( .x(\U7/ni ), .a(i[7]) );
    inv_1 \U7/Uih  ( .x(\U7/nh ), .a(h[7]) );
    inv_1 \U7/Uil  ( .x(\U7/nl ), .a(l[7]) );
    ao23_1 \U7/Ucl/U1/U1  ( .x(l[7]), .a(n7), .b(l[7]), .c(n3), .d(\U7/ni ), 
        .e(\U7/nh ) );
    ao23_1 \U7/Uch/U1/U1  ( .x(h[7]), .a(n7), .b(h[7]), .c(n2), .d(i[7]), .e(
        \U7/nl ) );
    inv_1 \U6/Uii  ( .x(\U6/ni ), .a(i[6]) );
    inv_1 \U6/Uih  ( .x(\U6/nh ), .a(h[6]) );
    inv_1 \U6/Uil  ( .x(\U6/nl ), .a(l[6]) );
    ao23_1 \U6/Ucl/U1/U1  ( .x(l[6]), .a(n7), .b(l[6]), .c(n2), .d(\U6/ni ), 
        .e(\U6/nh ) );
    ao23_1 \U6/Uch/U1/U1  ( .x(h[6]), .a(n7), .b(h[6]), .c(n2), .d(i[6]), .e(
        \U6/nl ) );
    inv_1 \U5/Uii  ( .x(\U5/ni ), .a(i[5]) );
    inv_1 \U5/Uih  ( .x(\U5/nh ), .a(h[5]) );
    inv_1 \U5/Uil  ( .x(\U5/nl ), .a(l[5]) );
    ao23_1 \U5/Ucl/U1/U1  ( .x(l[5]), .a(n7), .b(l[5]), .c(n2), .d(\U5/ni ), 
        .e(\U5/nh ) );
    ao23_1 \U5/Uch/U1/U1  ( .x(h[5]), .a(n7), .b(h[5]), .c(n2), .d(i[5]), .e(
        \U5/nl ) );
    inv_1 \U4/Uii  ( .x(\U4/ni ), .a(i[4]) );
    inv_1 \U4/Uih  ( .x(\U4/nh ), .a(h[4]) );
    inv_1 \U4/Uil  ( .x(\U4/nl ), .a(l[4]) );
    ao23_1 \U4/Ucl/U1/U1  ( .x(l[4]), .a(n6), .b(l[4]), .c(n2), .d(\U4/ni ), 
        .e(\U4/nh ) );
    ao23_1 \U4/Uch/U1/U1  ( .x(h[4]), .a(n6), .b(h[4]), .c(n2), .d(i[4]), .e(
        \U4/nl ) );
    inv_1 \U3/Uii  ( .x(\U3/ni ), .a(i[3]) );
    inv_1 \U3/Uih  ( .x(\U3/nh ), .a(h[3]) );
    inv_1 \U3/Uil  ( .x(\U3/nl ), .a(l[3]) );
    ao23_1 \U3/Ucl/U1/U1  ( .x(l[3]), .a(n6), .b(l[3]), .c(n2), .d(\U3/ni ), 
        .e(\U3/nh ) );
    ao23_1 \U3/Uch/U1/U1  ( .x(h[3]), .a(n8), .b(h[3]), .c(n1), .d(i[3]), .e(
        \U3/nl ) );
    inv_1 \U2/Uii  ( .x(\U2/ni ), .a(i[2]) );
    inv_1 \U2/Uih  ( .x(\U2/nh ), .a(h[2]) );
    inv_1 \U2/Uil  ( .x(\U2/nl ), .a(l[2]) );
    ao23_1 \U2/Ucl/U1/U1  ( .x(l[2]), .a(n8), .b(l[2]), .c(n1), .d(\U2/ni ), 
        .e(\U2/nh ) );
    ao23_1 \U2/Uch/U1/U1  ( .x(h[2]), .a(n8), .b(h[2]), .c(n1), .d(i[2]), .e(
        \U2/nl ) );
    inv_1 \U1/Uii  ( .x(\U1/ni ), .a(i[1]) );
    inv_1 \U1/Uih  ( .x(\U1/nh ), .a(h[1]) );
    inv_1 \U1/Uil  ( .x(\U1/nl ), .a(l[1]) );
    ao23_1 \U1/Ucl/U1/U1  ( .x(l[1]), .a(n8), .b(l[1]), .c(n1), .d(\U1/ni ), 
        .e(\U1/nh ) );
    ao23_1 \U1/Uch/U1/U1  ( .x(h[1]), .a(n8), .b(h[1]), .c(n1), .d(i[1]), .e(
        \U1/nl ) );
    inv_1 \U0/Uii  ( .x(\U0/ni ), .a(i[0]) );
    inv_1 \U0/Uih  ( .x(\U0/nh ), .a(h[0]) );
    inv_1 \U0/Uil  ( .x(\U0/nl ), .a(l[0]) );
    ao23_1 \U0/Ucl/U1/U1  ( .x(l[0]), .a(n8), .b(l[0]), .c(n1), .d(\U0/ni ), 
        .e(\U0/nh ) );
    ao23_1 \U0/Uch/U1/U1  ( .x(h[0]), .a(n8), .b(h[0]), .c(n1), .d(i[0]), .e(
        \U0/nl ) );
    buf_16 U1 ( .x(n1), .a(n12) );
    buf_16 U2 ( .x(n2), .a(n12) );
    buf_16 U3 ( .x(n3), .a(n12) );
    buf_16 U4 ( .x(n4), .a(n11) );
    buf_16 U5 ( .x(n5), .a(n11) );
    buf_16 U6 ( .x(n6), .a(n11) );
    buf_16 U7 ( .x(n7), .a(n10) );
    buf_16 U8 ( .x(n8), .a(n10) );
    buf_16 U9 ( .x(n9), .a(n10) );
    buf_16 U10 ( .x(n10), .a(req) );
    buf_16 U11 ( .x(n11), .a(req) );
    buf_16 U12 ( .x(n12), .a(req) );
endmodule


module sr2dr_word_0 ( i, req, h, l );
input  [31:0] i;
output [31:0] h;
output [31:0] l;
input  req;
    wire \U31/ni , \U31/nh , \U31/nl , n9, n1, n2, \U30/ni , \U30/nh , 
        \U30/nl , n8, \U29/ni , \U29/nh , \U29/nl , \U28/ni , \U28/nh , 
        \U28/nl , \U27/ni , \U27/nh , \U27/nl , \U26/ni , \U26/nh , \U26/nl , 
        n7, n4, \U25/ni , \U25/nh , \U25/nl , \U24/ni , \U24/nh , \U24/nl , 
        \U23/ni , \U23/nh , \U23/nl , n3, \U22/ni , \U22/nh , \U22/nl , n6, 
        \U21/ni , \U21/nh , \U21/nl , \U20/ni , \U20/nh , \U20/nl , n5, 
        \U19/ni , \U19/nh , \U19/nl , \U18/ni , \U18/nh , \U18/nl , \U17/ni , 
        \U17/nh , \U17/nl , \U16/ni , \U16/nh , \U16/nl , \U15/ni , \U15/nh , 
        \U15/nl , \U14/ni , \U14/nh , \U14/nl , \U13/ni , \U13/nh , \U13/nl , 
        \U12/ni , \U12/nh , \U12/nl , \U11/ni , \U11/nh , \U11/nl , \U10/ni , 
        \U10/nh , \U10/nl , \U9/ni , \U9/nh , \U9/nl , \U8/ni , \U8/nh , 
        \U8/nl , \U7/ni , \U7/nh , \U7/nl , \U6/ni , \U6/nh , \U6/nl , \U5/ni , 
        \U5/nh , \U5/nl , \U4/ni , \U4/nh , \U4/nl , \U3/ni , \U3/nh , \U3/nl , 
        \U2/ni , \U2/nh , \U2/nl , \U1/ni , \U1/nh , \U1/nl , \U0/ni , \U0/nh , 
        \U0/nl , n12, n11, n10;
    inv_1 \U31/Uii  ( .x(\U31/ni ), .a(i[31]) );
    inv_1 \U31/Uih  ( .x(\U31/nh ), .a(h[31]) );
    inv_1 \U31/Uil  ( .x(\U31/nl ), .a(l[31]) );
    ao23_1 \U31/Ucl/U1/U1  ( .x(l[31]), .a(n9), .b(l[31]), .c(n1), .d(\U31/ni 
        ), .e(\U31/nh ) );
    ao23_1 \U31/Uch/U1/U1  ( .x(h[31]), .a(n9), .b(h[31]), .c(n2), .d(i[31]), 
        .e(\U31/nl ) );
    inv_1 \U30/Uii  ( .x(\U30/ni ), .a(i[30]) );
    inv_1 \U30/Uih  ( .x(\U30/nh ), .a(h[30]) );
    inv_1 \U30/Uil  ( .x(\U30/nl ), .a(l[30]) );
    ao23_1 \U30/Ucl/U1/U1  ( .x(l[30]), .a(n8), .b(l[30]), .c(n1), .d(\U30/ni 
        ), .e(\U30/nh ) );
    ao23_1 \U30/Uch/U1/U1  ( .x(h[30]), .a(n8), .b(h[30]), .c(n1), .d(i[30]), 
        .e(\U30/nl ) );
    inv_1 \U29/Uii  ( .x(\U29/ni ), .a(i[29]) );
    inv_1 \U29/Uih  ( .x(\U29/nh ), .a(h[29]) );
    inv_1 \U29/Uil  ( .x(\U29/nl ), .a(l[29]) );
    ao23_1 \U29/Ucl/U1/U1  ( .x(l[29]), .a(n8), .b(l[29]), .c(n1), .d(\U29/ni 
        ), .e(\U29/nh ) );
    ao23_1 \U29/Uch/U1/U1  ( .x(h[29]), .a(n8), .b(h[29]), .c(n2), .d(i[29]), 
        .e(\U29/nl ) );
    inv_1 \U28/Uii  ( .x(\U28/ni ), .a(i[28]) );
    inv_1 \U28/Uih  ( .x(\U28/nh ), .a(h[28]) );
    inv_1 \U28/Uil  ( .x(\U28/nl ), .a(l[28]) );
    ao23_1 \U28/Ucl/U1/U1  ( .x(l[28]), .a(n8), .b(l[28]), .c(n2), .d(\U28/ni 
        ), .e(\U28/nh ) );
    ao23_1 \U28/Uch/U1/U1  ( .x(h[28]), .a(n8), .b(h[28]), .c(n2), .d(i[28]), 
        .e(\U28/nl ) );
    inv_1 \U27/Uii  ( .x(\U27/ni ), .a(i[27]) );
    inv_1 \U27/Uih  ( .x(\U27/nh ), .a(h[27]) );
    inv_1 \U27/Uil  ( .x(\U27/nl ), .a(l[27]) );
    ao23_1 \U27/Ucl/U1/U1  ( .x(l[27]), .a(n8), .b(l[27]), .c(n2), .d(\U27/ni 
        ), .e(\U27/nh ) );
    ao23_1 \U27/Uch/U1/U1  ( .x(h[27]), .a(n8), .b(h[27]), .c(n2), .d(i[27]), 
        .e(\U27/nl ) );
    inv_1 \U26/Uii  ( .x(\U26/ni ), .a(i[26]) );
    inv_1 \U26/Uih  ( .x(\U26/nh ), .a(h[26]) );
    inv_1 \U26/Uil  ( .x(\U26/nl ), .a(l[26]) );
    ao23_1 \U26/Ucl/U1/U1  ( .x(l[26]), .a(n7), .b(l[26]), .c(n2), .d(\U26/ni 
        ), .e(\U26/nh ) );
    ao23_1 \U26/Uch/U1/U1  ( .x(h[26]), .a(n7), .b(h[26]), .c(n4), .d(i[26]), 
        .e(\U26/nl ) );
    inv_1 \U25/Uii  ( .x(\U25/ni ), .a(i[25]) );
    inv_1 \U25/Uih  ( .x(\U25/nh ), .a(h[25]) );
    inv_1 \U25/Uil  ( .x(\U25/nl ), .a(l[25]) );
    ao23_1 \U25/Ucl/U1/U1  ( .x(l[25]), .a(n7), .b(l[25]), .c(n4), .d(\U25/ni 
        ), .e(\U25/nh ) );
    ao23_1 \U25/Uch/U1/U1  ( .x(h[25]), .a(n7), .b(h[25]), .c(n4), .d(i[25]), 
        .e(\U25/nl ) );
    inv_1 \U24/Uii  ( .x(\U24/ni ), .a(i[24]) );
    inv_1 \U24/Uih  ( .x(\U24/nh ), .a(h[24]) );
    inv_1 \U24/Uil  ( .x(\U24/nl ), .a(l[24]) );
    ao23_1 \U24/Ucl/U1/U1  ( .x(l[24]), .a(n7), .b(l[24]), .c(n4), .d(\U24/ni 
        ), .e(\U24/nh ) );
    ao23_1 \U24/Uch/U1/U1  ( .x(h[24]), .a(n7), .b(h[24]), .c(n4), .d(i[24]), 
        .e(\U24/nl ) );
    inv_1 \U23/Uii  ( .x(\U23/ni ), .a(i[23]) );
    inv_1 \U23/Uih  ( .x(\U23/nh ), .a(h[23]) );
    inv_1 \U23/Uil  ( .x(\U23/nl ), .a(l[23]) );
    ao23_1 \U23/Ucl/U1/U1  ( .x(l[23]), .a(n7), .b(l[23]), .c(n3), .d(\U23/ni 
        ), .e(\U23/nh ) );
    ao23_1 \U23/Uch/U1/U1  ( .x(h[23]), .a(n7), .b(h[23]), .c(n3), .d(i[23]), 
        .e(\U23/nl ) );
    inv_1 \U22/Uii  ( .x(\U22/ni ), .a(i[22]) );
    inv_1 \U22/Uih  ( .x(\U22/nh ), .a(h[22]) );
    inv_1 \U22/Uil  ( .x(\U22/nl ), .a(l[22]) );
    ao23_1 \U22/Ucl/U1/U1  ( .x(l[22]), .a(n6), .b(l[22]), .c(n3), .d(\U22/ni 
        ), .e(\U22/nh ) );
    ao23_1 \U22/Uch/U1/U1  ( .x(h[22]), .a(n6), .b(h[22]), .c(n3), .d(i[22]), 
        .e(\U22/nl ) );
    inv_1 \U21/Uii  ( .x(\U21/ni ), .a(i[21]) );
    inv_1 \U21/Uih  ( .x(\U21/nh ), .a(h[21]) );
    inv_1 \U21/Uil  ( .x(\U21/nl ), .a(l[21]) );
    ao23_1 \U21/Ucl/U1/U1  ( .x(l[21]), .a(n6), .b(l[21]), .c(n3), .d(\U21/ni 
        ), .e(\U21/nh ) );
    ao23_1 \U21/Uch/U1/U1  ( .x(h[21]), .a(n6), .b(h[21]), .c(n3), .d(i[21]), 
        .e(\U21/nl ) );
    inv_1 \U20/Uii  ( .x(\U20/ni ), .a(i[20]) );
    inv_1 \U20/Uih  ( .x(\U20/nh ), .a(h[20]) );
    inv_1 \U20/Uil  ( .x(\U20/nl ), .a(l[20]) );
    ao23_1 \U20/Ucl/U1/U1  ( .x(l[20]), .a(n6), .b(l[20]), .c(n5), .d(\U20/ni 
        ), .e(\U20/nh ) );
    ao23_1 \U20/Uch/U1/U1  ( .x(h[20]), .a(n6), .b(h[20]), .c(n4), .d(i[20]), 
        .e(\U20/nl ) );
    inv_1 \U19/Uii  ( .x(\U19/ni ), .a(i[19]) );
    inv_1 \U19/Uih  ( .x(\U19/nh ), .a(h[19]) );
    inv_1 \U19/Uil  ( .x(\U19/nl ), .a(l[19]) );
    ao23_1 \U19/Ucl/U1/U1  ( .x(l[19]), .a(n6), .b(l[19]), .c(n4), .d(\U19/ni 
        ), .e(\U19/nh ) );
    ao23_1 \U19/Uch/U1/U1  ( .x(h[19]), .a(n6), .b(h[19]), .c(n4), .d(i[19]), 
        .e(\U19/nl ) );
    inv_1 \U18/Uii  ( .x(\U18/ni ), .a(i[18]) );
    inv_1 \U18/Uih  ( .x(\U18/nh ), .a(h[18]) );
    inv_1 \U18/Uil  ( .x(\U18/nl ), .a(l[18]) );
    ao23_1 \U18/Ucl/U1/U1  ( .x(l[18]), .a(n5), .b(l[18]), .c(n5), .d(\U18/ni 
        ), .e(\U18/nh ) );
    ao23_1 \U18/Uch/U1/U1  ( .x(h[18]), .a(n5), .b(h[18]), .c(n5), .d(i[18]), 
        .e(\U18/nl ) );
    inv_1 \U17/Uii  ( .x(\U17/ni ), .a(i[17]) );
    inv_1 \U17/Uih  ( .x(\U17/nh ), .a(h[17]) );
    inv_1 \U17/Uil  ( .x(\U17/nl ), .a(l[17]) );
    ao23_1 \U17/Ucl/U1/U1  ( .x(l[17]), .a(n6), .b(l[17]), .c(n5), .d(\U17/ni 
        ), .e(\U17/nh ) );
    ao23_1 \U17/Uch/U1/U1  ( .x(h[17]), .a(n7), .b(h[17]), .c(n4), .d(i[17]), 
        .e(\U17/nl ) );
    inv_1 \U16/Uii  ( .x(\U16/ni ), .a(i[16]) );
    inv_1 \U16/Uih  ( .x(\U16/nh ), .a(h[16]) );
    inv_1 \U16/Uil  ( .x(\U16/nl ), .a(l[16]) );
    ao23_1 \U16/Ucl/U1/U1  ( .x(l[16]), .a(n9), .b(l[16]), .c(n3), .d(\U16/ni 
        ), .e(\U16/nh ) );
    ao23_1 \U16/Uch/U1/U1  ( .x(h[16]), .a(n9), .b(h[16]), .c(n1), .d(i[16]), 
        .e(\U16/nl ) );
    inv_1 \U15/Uii  ( .x(\U15/ni ), .a(i[15]) );
    inv_1 \U15/Uih  ( .x(\U15/nh ), .a(h[15]) );
    inv_1 \U15/Uil  ( .x(\U15/nl ), .a(l[15]) );
    ao23_1 \U15/Ucl/U1/U1  ( .x(l[15]), .a(n8), .b(l[15]), .c(n1), .d(\U15/ni 
        ), .e(\U15/nh ) );
    ao23_1 \U15/Uch/U1/U1  ( .x(h[15]), .a(n7), .b(h[15]), .c(n1), .d(i[15]), 
        .e(\U15/nl ) );
    inv_1 \U14/Uii  ( .x(\U14/ni ), .a(i[14]) );
    inv_1 \U14/Uih  ( .x(\U14/nh ), .a(h[14]) );
    inv_1 \U14/Uil  ( .x(\U14/nl ), .a(l[14]) );
    ao23_1 \U14/Ucl/U1/U1  ( .x(l[14]), .a(n6), .b(l[14]), .c(n1), .d(\U14/ni 
        ), .e(\U14/nh ) );
    ao23_1 \U14/Uch/U1/U1  ( .x(h[14]), .a(n6), .b(h[14]), .c(n3), .d(i[14]), 
        .e(\U14/nl ) );
    inv_1 \U13/Uii  ( .x(\U13/ni ), .a(i[13]) );
    inv_1 \U13/Uih  ( .x(\U13/nh ), .a(h[13]) );
    inv_1 \U13/Uil  ( .x(\U13/nl ), .a(l[13]) );
    ao23_1 \U13/Ucl/U1/U1  ( .x(l[13]), .a(n6), .b(l[13]), .c(n4), .d(\U13/ni 
        ), .e(\U13/nh ) );
    ao23_1 \U13/Uch/U1/U1  ( .x(h[13]), .a(n6), .b(h[13]), .c(n4), .d(i[13]), 
        .e(\U13/nl ) );
    inv_1 \U12/Uii  ( .x(\U12/ni ), .a(i[12]) );
    inv_1 \U12/Uih  ( .x(\U12/nh ), .a(h[12]) );
    inv_1 \U12/Uil  ( .x(\U12/nl ), .a(l[12]) );
    ao23_1 \U12/Ucl/U1/U1  ( .x(l[12]), .a(n5), .b(l[12]), .c(n4), .d(\U12/ni 
        ), .e(\U12/nh ) );
    ao23_1 \U12/Uch/U1/U1  ( .x(h[12]), .a(n5), .b(h[12]), .c(n4), .d(i[12]), 
        .e(\U12/nl ) );
    inv_1 \U11/Uii  ( .x(\U11/ni ), .a(i[11]) );
    inv_1 \U11/Uih  ( .x(\U11/nh ), .a(h[11]) );
    inv_1 \U11/Uil  ( .x(\U11/nl ), .a(l[11]) );
    ao23_1 \U11/Ucl/U1/U1  ( .x(l[11]), .a(n5), .b(l[11]), .c(n4), .d(\U11/ni 
        ), .e(\U11/nh ) );
    ao23_1 \U11/Uch/U1/U1  ( .x(h[11]), .a(n5), .b(h[11]), .c(n4), .d(i[11]), 
        .e(\U11/nl ) );
    inv_1 \U10/Uii  ( .x(\U10/ni ), .a(i[10]) );
    inv_1 \U10/Uih  ( .x(\U10/nh ), .a(h[10]) );
    inv_1 \U10/Uil  ( .x(\U10/nl ), .a(l[10]) );
    ao23_1 \U10/Ucl/U1/U1  ( .x(l[10]), .a(n5), .b(l[10]), .c(n3), .d(\U10/ni 
        ), .e(\U10/nh ) );
    ao23_1 \U10/Uch/U1/U1  ( .x(h[10]), .a(n5), .b(h[10]), .c(n3), .d(i[10]), 
        .e(\U10/nl ) );
    inv_1 \U9/Uii  ( .x(\U9/ni ), .a(i[9]) );
    inv_1 \U9/Uih  ( .x(\U9/nh ), .a(h[9]) );
    inv_1 \U9/Uil  ( .x(\U9/nl ), .a(l[9]) );
    ao23_1 \U9/Ucl/U1/U1  ( .x(l[9]), .a(n5), .b(l[9]), .c(n3), .d(\U9/ni ), 
        .e(\U9/nh ) );
    ao23_1 \U9/Uch/U1/U1  ( .x(h[9]), .a(n5), .b(h[9]), .c(n3), .d(i[9]), .e(
        \U9/nl ) );
    inv_1 \U8/Uii  ( .x(\U8/ni ), .a(i[8]) );
    inv_1 \U8/Uih  ( .x(\U8/nh ), .a(h[8]) );
    inv_1 \U8/Uil  ( .x(\U8/nl ), .a(l[8]) );
    ao23_1 \U8/Ucl/U1/U1  ( .x(l[8]), .a(n5), .b(l[8]), .c(n3), .d(\U8/ni ), 
        .e(\U8/nh ) );
    ao23_1 \U8/Uch/U1/U1  ( .x(h[8]), .a(n5), .b(h[8]), .c(n3), .d(i[8]), .e(
        \U8/nl ) );
    inv_1 \U7/Uii  ( .x(\U7/ni ), .a(i[7]) );
    inv_1 \U7/Uih  ( .x(\U7/nh ), .a(h[7]) );
    inv_1 \U7/Uil  ( .x(\U7/nl ), .a(l[7]) );
    ao23_1 \U7/Ucl/U1/U1  ( .x(l[7]), .a(n7), .b(l[7]), .c(n3), .d(\U7/ni ), 
        .e(\U7/nh ) );
    ao23_1 \U7/Uch/U1/U1  ( .x(h[7]), .a(n7), .b(h[7]), .c(n2), .d(i[7]), .e(
        \U7/nl ) );
    inv_1 \U6/Uii  ( .x(\U6/ni ), .a(i[6]) );
    inv_1 \U6/Uih  ( .x(\U6/nh ), .a(h[6]) );
    inv_1 \U6/Uil  ( .x(\U6/nl ), .a(l[6]) );
    ao23_1 \U6/Ucl/U1/U1  ( .x(l[6]), .a(n7), .b(l[6]), .c(n2), .d(\U6/ni ), 
        .e(\U6/nh ) );
    ao23_1 \U6/Uch/U1/U1  ( .x(h[6]), .a(n7), .b(h[6]), .c(n2), .d(i[6]), .e(
        \U6/nl ) );
    inv_1 \U5/Uii  ( .x(\U5/ni ), .a(i[5]) );
    inv_1 \U5/Uih  ( .x(\U5/nh ), .a(h[5]) );
    inv_1 \U5/Uil  ( .x(\U5/nl ), .a(l[5]) );
    ao23_1 \U5/Ucl/U1/U1  ( .x(l[5]), .a(n7), .b(l[5]), .c(n2), .d(\U5/ni ), 
        .e(\U5/nh ) );
    ao23_1 \U5/Uch/U1/U1  ( .x(h[5]), .a(n7), .b(h[5]), .c(n2), .d(i[5]), .e(
        \U5/nl ) );
    inv_1 \U4/Uii  ( .x(\U4/ni ), .a(i[4]) );
    inv_1 \U4/Uih  ( .x(\U4/nh ), .a(h[4]) );
    inv_1 \U4/Uil  ( .x(\U4/nl ), .a(l[4]) );
    ao23_1 \U4/Ucl/U1/U1  ( .x(l[4]), .a(n6), .b(l[4]), .c(n2), .d(\U4/ni ), 
        .e(\U4/nh ) );
    ao23_1 \U4/Uch/U1/U1  ( .x(h[4]), .a(n6), .b(h[4]), .c(n2), .d(i[4]), .e(
        \U4/nl ) );
    inv_1 \U3/Uii  ( .x(\U3/ni ), .a(i[3]) );
    inv_1 \U3/Uih  ( .x(\U3/nh ), .a(h[3]) );
    inv_1 \U3/Uil  ( .x(\U3/nl ), .a(l[3]) );
    ao23_1 \U3/Ucl/U1/U1  ( .x(l[3]), .a(n6), .b(l[3]), .c(n2), .d(\U3/ni ), 
        .e(\U3/nh ) );
    ao23_1 \U3/Uch/U1/U1  ( .x(h[3]), .a(n8), .b(h[3]), .c(n1), .d(i[3]), .e(
        \U3/nl ) );
    inv_1 \U2/Uii  ( .x(\U2/ni ), .a(i[2]) );
    inv_1 \U2/Uih  ( .x(\U2/nh ), .a(h[2]) );
    inv_1 \U2/Uil  ( .x(\U2/nl ), .a(l[2]) );
    ao23_1 \U2/Ucl/U1/U1  ( .x(l[2]), .a(n8), .b(l[2]), .c(n1), .d(\U2/ni ), 
        .e(\U2/nh ) );
    ao23_1 \U2/Uch/U1/U1  ( .x(h[2]), .a(n8), .b(h[2]), .c(n1), .d(i[2]), .e(
        \U2/nl ) );
    inv_1 \U1/Uii  ( .x(\U1/ni ), .a(i[1]) );
    inv_1 \U1/Uih  ( .x(\U1/nh ), .a(h[1]) );
    inv_1 \U1/Uil  ( .x(\U1/nl ), .a(l[1]) );
    ao23_1 \U1/Ucl/U1/U1  ( .x(l[1]), .a(n8), .b(l[1]), .c(n1), .d(\U1/ni ), 
        .e(\U1/nh ) );
    ao23_1 \U1/Uch/U1/U1  ( .x(h[1]), .a(n8), .b(h[1]), .c(n1), .d(i[1]), .e(
        \U1/nl ) );
    inv_1 \U0/Uii  ( .x(\U0/ni ), .a(i[0]) );
    inv_1 \U0/Uih  ( .x(\U0/nh ), .a(h[0]) );
    inv_1 \U0/Uil  ( .x(\U0/nl ), .a(l[0]) );
    ao23_1 \U0/Ucl/U1/U1  ( .x(l[0]), .a(n8), .b(l[0]), .c(n1), .d(\U0/ni ), 
        .e(\U0/nh ) );
    ao23_1 \U0/Uch/U1/U1  ( .x(h[0]), .a(n8), .b(h[0]), .c(n1), .d(i[0]), .e(
        \U0/nl ) );
    buf_16 U1 ( .x(n1), .a(n12) );
    buf_16 U2 ( .x(n2), .a(n12) );
    buf_16 U3 ( .x(n3), .a(n12) );
    buf_16 U4 ( .x(n4), .a(n11) );
    buf_16 U5 ( .x(n5), .a(n11) );
    buf_16 U6 ( .x(n6), .a(n11) );
    buf_16 U7 ( .x(n7), .a(n10) );
    buf_16 U8 ( .x(n8), .a(n10) );
    buf_16 U9 ( .x(n9), .a(n10) );
    buf_16 U10 ( .x(n10), .a(req) );
    buf_16 U11 ( .x(n11), .a(req) );
    buf_16 U12 ( .x(n12), .a(req) );
endmodule


module latch_ctrl_0 ( rin, ain, rout, aout, en, reset );
input  rin, aout, reset;
output ain, rout, en;
    wire nreset, na, n1, a, N6, N5, n_rout, n3, \c_rout/ob ;
    inv_1 U0 ( .x(nreset), .a(reset) );
    nor2_1 U1 ( .x(ain), .a(na), .b(n1) );
    inv_1 U2 ( .x(na), .a(a) );
    inv_1 U3 ( .x(N6), .a(N5) );
    inv_1 U4 ( .x(rout), .a(n_rout) );
    and2_1 C9 ( .x(n3), .a(na), .b(N6) );
    or2_1 C11 ( .x(N5), .a(rout), .b(aout) );
    oa21_1 \c_na/__tmp99/U1  ( .x(a), .a(n1), .b(a), .c(rin) );
    oai21_1 \c_rout/U1  ( .x(\c_rout/ob ), .a(aout), .b(n_rout), .c(na) );
    nand2_1 \c_rout/U2  ( .x(n_rout), .a(nreset), .b(\c_rout/ob ) );
    buf_1 U5 ( .x(en), .a(n3) );
    buf_1 U6 ( .x(n1), .a(n3) );
endmodule


module matched_delay_m2cp_resp_iport ( x, a );
input  a;
output x;
    assign x = a;
endmodule


module m2cp_iport ( req_in, ts_o, sel_o, mult_o, we_o, prd_o, seq_o, adr_o, 
    dat_o, ain, ic_seq, ic_pred, ic_size, ic_itag, ic_wd, ic_lock, ic_a, 
    ic_rnw, ic_col, ic_ack, req_out, ts_i, we_i, err_i, rty_i, acc_i, dat_i, 
    aout, ir_rd, ir_err, ir_rnw, ir_ack, tag_id, reset );
input  [2:0] ts_o;
input  [3:0] sel_o;
input  [31:0] adr_o;
input  [31:0] dat_o;
output [1:0] ic_seq;
output [1:0] ic_pred;
output [3:0] ic_size;
output [9:0] ic_itag;
output [63:0] ic_wd;
output [1:0] ic_lock;
output [63:0] ic_a;
output [1:0] ic_rnw;
output [5:0] ic_col;
output [2:0] ts_i;
output [31:0] dat_i;
input  [63:0] ir_rd;
input  [1:0] ir_err;
input  [1:0] ir_rnw;
input  [4:0] tag_id;
input  req_in, mult_o, we_o, prd_o, seq_o, ic_ack, aout, reset;
output ain, req_out, we_i, err_i, rty_i, acc_i, ir_ack;
    wire req_in_delayed, n8, \data[15] , \data[14] , \data[13] , \data[12] , 
        \data[11] , \data[10] , \data[9] , \data[8] , \data[7] , \data[6] , 
        \data[5] , \data[4] , \data[3] , \data[2] , \data[1] , \data[0] , 
        complete_delayed, en, _26_net_, n72, n77, _27_net_, _24_net_, n112, 
        n124, n118, n206, n208, n210, n197, n199, n202, n201, n203, n204, 
        \size[1] , n83, n84, n89, n205, n64, n2, n90, n97, n198, n3, n98, n87, 
        n63, n4, n88, n85, n5, n86, n290, n289, n288, n79, n277, n270, n273, 
        n276, n266, n269, n283, n282, n281, n298, n70, n68, n213, n223, n80, 
        n291, n284, n287, n280, n99, n100, n95, n96, n93, n94, n91, n92, n81, 
        all_r, n69, n300, n294, n302, n296, n306, n292, n304, low_ir_rd, n73, 
        n74, n75, n76, complete, n82, n200, n207, n209, n211, n224, n225, n226, 
        n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, 
        n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, 
        n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, 
        n263, n265, n264, n268, n267, n272, n271, n275, n274, n279, n278, n286, 
        n285, n293, n295, n297, n299, n301, n303, n305, n307, n222, n221, n220, 
        n219, n218, n217, n216, n215, all_w, n65, n214, high_ir_rd, \size[0] , 
        n212, n308, n182, n179, n176, n173, n194, n191, n188, n185, n158, n155, 
        n152, n149, n170, n167, n164, n161, n134, n131, n128, n125, n146, n143, 
        n140, n137, n110, n107, n104, n101, n122, n119, n116, n113, n183, n184, 
        n180, n181, n177, n178, n174, n175, n195, n196, n192, n193, n189, n190, 
        n186, n187, n159, n160, n156, n157, n153, n154, n150, n151, n171, n172, 
        n168, n169, n165, n166, n162, n163, n135, n136, n132, n133, n129, n130, 
        n126, n127, n147, n148, n144, n145, n141, n142, n138, n139, n111, n108, 
        n109, n105, n106, n102, n103, n123, n120, n121, n117, n114, n115, n7, 
        n6, n1, _28_net_, comp_basic, \all_read/__tmp99/loop , comp_rd, 
        _25_net_, \Ucol2/ni , \Ucol2/nh , \Ucol2/nl , n11, \Ucol1/ni , 
        \Ucol1/nh , \Ucol1/nl , n9, \Ucol0/ni , \Ucol0/nh , \Ucol0/nl , n10, 
        \Utag4/ni , \Utag4/nh , \Utag4/nl , \Utag3/ni , \Utag3/nh , \Utag3/nl , 
        \Utag2/ni , \Utag2/nh , \Utag2/nl , \Utag1/ni , \Utag1/nh , \Utag1/nl , 
        \Utag0/ni , \Utag0/nh , \Utag0/nl , \Usze1/ni , \Usze1/nh , \Usze1/nl , 
        \Usze0/ni , \Usze0/nh , \Usze0/nl , \Urnw/ni , \Urnw/nh , \Urnw/nl , 
        \Ulock/ni , \Ulock/nh , \Ulock/nl , \Upred/ni , \Upred/nh , \Upred/nl , 
        \Useq/ni , \Useq/nh , \Useq/nl , n78;
    assign ain = ic_ack;
    assign ts_i[2] = 1'b0;
    assign ts_i[1] = 1'b0;
    assign ts_i[0] = 1'b0;
    assign rty_i = 1'b0;
    assign acc_i = 1'b0;
    matched_delay_m2cp_com_iport U130 ( .x(req_in_delayed), .a(req_in) );
    sr2dr_word_1 Uwd ( .i({dat_o[31], dat_o[30], dat_o[29], dat_o[28], 
        dat_o[27], dat_o[26], dat_o[25], dat_o[24], dat_o[23], dat_o[22], 
        dat_o[21], dat_o[20], dat_o[19], dat_o[18], dat_o[17], dat_o[16], 
        \data[15] , \data[14] , \data[13] , \data[12] , \data[11] , \data[10] , 
        \data[9] , \data[8] , \data[7] , \data[6] , \data[5] , \data[4] , 
        \data[3] , \data[2] , \data[1] , \data[0] }), .req(n8), .h(ic_wd
        [63:32]), .l(ic_wd[31:0]) );
    sr2dr_word_0 Ua ( .i(adr_o), .req(n8), .h(ic_a[63:32]), .l(ic_a[31:0]) );
    latch_ctrl_0 lc ( .rin(complete_delayed), .ain(ir_ack), .rout(req_out), 
        .aout(aout), .en(en), .reset(reset) );
    nand2_1 U61 ( .x(_26_net_), .a(n72), .b(n77) );
    and2_1 U274 ( .x(_27_net_), .a(ir_rnw[1]), .b(ir_err[0]) );
    inv_1 U275 ( .x(_24_net_), .a(we_o) );
    inv_1 U2 ( .x(n112), .a(ir_rd[4]) );
    inv_1 U3 ( .x(n124), .a(ir_rd[0]) );
    inv_1 U4 ( .x(n118), .a(ir_rd[2]) );
    inv_1 U5 ( .x(n206), .a(dat_o[28]) );
    inv_1 U6 ( .x(n208), .a(dat_o[27]) );
    inv_1 U7 ( .x(n210), .a(dat_o[26]) );
    inv_1 U8 ( .x(n197), .a(dat_o[25]) );
    inv_1 U9 ( .x(n199), .a(dat_o[24]) );
    inv_1 U10 ( .x(n202), .a(dat_o[15]) );
    inv_1 U11 ( .x(n201), .a(dat_o[31]) );
    inv_1 U12 ( .x(n203), .a(dat_o[30]) );
    inv_1 U13 ( .x(n204), .a(dat_o[29]) );
    nor2_1 U14 ( .x(\size[1] ), .a(n83), .b(n84) );
    inv_1 U15 ( .x(n72), .a(ir_rnw[0]) );
    oa21_1 U16 ( .x(n89), .a(n205), .b(n64), .c(n2) );
    inv_1 U24 ( .x(n2), .a(n90) );
    inv_1 U17 ( .x(n205), .a(dat_o[13]) );
    inv_1 U18 ( .x(n64), .a(sel_o[1]) );
    oa21_1 U19 ( .x(n97), .a(n198), .b(n64), .c(n3) );
    inv_1 U276 ( .x(n3), .a(n98) );
    inv_1 U20 ( .x(n198), .a(dat_o[9]) );
    oa21_1 U21 ( .x(n87), .a(n63), .b(n64), .c(n4) );
    inv_1 U277 ( .x(n4), .a(n88) );
    inv_1 U22 ( .x(n63), .a(dat_o[14]) );
    oa21_1 U23 ( .x(n85), .a(n202), .b(n64), .c(n5) );
    inv_1 U278 ( .x(n5), .a(n86) );
    nand2_1 U25 ( .x(n290), .a(n289), .b(n288) );
    nand2_1 U26 ( .x(n79), .a(n277), .b(n270) );
    nor2_1 U27 ( .x(n277), .a(n273), .b(n276) );
    nor2_1 U28 ( .x(n270), .a(n266), .b(n269) );
    nand2_1 U29 ( .x(n283), .a(n282), .b(n281) );
    nand2_1 U30 ( .x(n298), .a(dat_o[20]), .b(n70) );
    inv_1 U31 ( .x(n70), .a(n68) );
    nand2_1 U32 ( .x(n213), .a(n223), .b(sel_o[1]) );
    nand2_1 U33 ( .x(n80), .a(n291), .b(n284) );
    nor2_1 U34 ( .x(n291), .a(n287), .b(n290) );
    nor2_1 U35 ( .x(n284), .a(n280), .b(n283) );
    aoi21_1 U36 ( .x(n99), .a(dat_o[8]), .b(sel_o[1]), .c(n100) );
    aoi21_1 U37 ( .x(n95), .a(dat_o[10]), .b(sel_o[1]), .c(n96) );
    aoi21_1 U38 ( .x(n93), .a(dat_o[11]), .b(sel_o[1]), .c(n94) );
    aoi21_1 U39 ( .x(n91), .a(dat_o[12]), .b(sel_o[1]), .c(n92) );
    inv_1 U40 ( .x(n81), .a(all_r) );
    nand2_1 U42 ( .x(n84), .a(sel_o[0]), .b(sel_o[1]) );
    inv_1 U45 ( .x(n68), .a(sel_o[2]) );
    inv_1 U46 ( .x(n69), .a(n68) );
    nand2_1 U51 ( .x(n300), .a(dat_o[19]), .b(n69) );
    nand2_1 U52 ( .x(n294), .a(dat_o[22]), .b(n69) );
    nand2_1 U53 ( .x(n302), .a(dat_o[18]), .b(n69) );
    nand2_1 U54 ( .x(n296), .a(dat_o[21]), .b(n69) );
    nand2_1 U55 ( .x(n306), .a(dat_o[16]), .b(n69) );
    nand2_1 U56 ( .x(n292), .a(dat_o[23]), .b(n69) );
    nand2_1 U57 ( .x(n304), .a(dat_o[17]), .b(n69) );
    nand4_1 U60 ( .x(low_ir_rd), .a(n73), .b(n74), .c(n75), .d(n76) );
    nand2_1 U62 ( .x(complete), .a(n81), .b(n82) );
    matched_delay_m2cp_resp_iport mdel ( .x(complete_delayed), .a(complete) );
    inv_1 U63 ( .x(n200), .a(dat_o[8]) );
    inv_1 U64 ( .x(n207), .a(dat_o[12]) );
    inv_1 U65 ( .x(n209), .a(dat_o[11]) );
    inv_1 U66 ( .x(n211), .a(dat_o[10]) );
    nand4_1 U67 ( .x(n224), .a(n225), .b(n226), .c(n227), .d(n228) );
    nand4_1 U68 ( .x(n229), .a(n230), .b(n231), .c(n232), .d(n233) );
    nor2_1 U69 ( .x(n76), .a(n224), .b(n229) );
    nand4_1 U70 ( .x(n234), .a(n235), .b(n236), .c(n237), .d(n238) );
    nand4_1 U71 ( .x(n239), .a(n240), .b(n241), .c(n242), .d(n243) );
    nor2_1 U72 ( .x(n75), .a(n234), .b(n239) );
    nand4_1 U73 ( .x(n244), .a(n245), .b(n246), .c(n247), .d(n248) );
    nand4_1 U74 ( .x(n249), .a(n250), .b(n251), .c(n252), .d(n253) );
    nor2_1 U75 ( .x(n74), .a(n244), .b(n249) );
    nand4_1 U76 ( .x(n254), .a(n255), .b(n256), .c(n257), .d(n258) );
    nand4_1 U77 ( .x(n259), .a(n260), .b(n261), .c(n262), .d(n263) );
    nor2_1 U78 ( .x(n73), .a(n254), .b(n259) );
    nand2_1 U79 ( .x(n266), .a(n265), .b(n264) );
    nand2_1 U80 ( .x(n269), .a(n268), .b(n267) );
    nand2_1 U81 ( .x(n273), .a(n272), .b(n271) );
    nand2_1 U82 ( .x(n276), .a(n275), .b(n274) );
    nand2_1 U83 ( .x(n280), .a(n279), .b(n278) );
    nand2_1 U84 ( .x(n287), .a(n286), .b(n285) );
    nand2_1 U85 ( .x(n86), .a(n292), .b(n293) );
    nand2_1 U86 ( .x(n88), .a(n294), .b(n295) );
    nand2_1 U87 ( .x(n90), .a(n296), .b(n297) );
    nand2_1 U88 ( .x(n92), .a(n298), .b(n299) );
    nand2_1 U89 ( .x(n94), .a(n300), .b(n301) );
    nand2_1 U90 ( .x(n96), .a(n302), .b(n303) );
    nand2_1 U91 ( .x(n98), .a(n304), .b(n305) );
    nand2_1 U92 ( .x(n100), .a(n306), .b(n307) );
    inv_1 U93 ( .x(n222), .a(dat_o[0]) );
    inv_1 U94 ( .x(n221), .a(dat_o[1]) );
    inv_1 U95 ( .x(n220), .a(dat_o[2]) );
    inv_1 U96 ( .x(n219), .a(dat_o[3]) );
    inv_1 U97 ( .x(n218), .a(dat_o[4]) );
    inv_1 U98 ( .x(n217), .a(dat_o[5]) );
    inv_1 U99 ( .x(n216), .a(dat_o[6]) );
    inv_1 U100 ( .x(n215), .a(dat_o[7]) );
    inv_1 U101 ( .x(n77), .a(ir_rnw[1]) );
    inv_1 U103 ( .x(n82), .a(all_w) );
    nand2_1 U104 ( .x(n293), .a(dat_o[31]), .b(sel_o[3]) );
    nand2_1 U105 ( .x(n295), .a(dat_o[30]), .b(sel_o[3]) );
    nand2_1 U109 ( .x(n303), .a(dat_o[26]), .b(sel_o[3]) );
    nand2_1 U110 ( .x(n305), .a(dat_o[25]), .b(sel_o[3]) );
    nand2_1 U111 ( .x(n307), .a(dat_o[24]), .b(sel_o[3]) );
    mux2i_1 U113 ( .x(\data[0] ), .d0(n99), .sl(n65), .d1(n222) );
    mux2i_1 U114 ( .x(\data[10] ), .d0(n211), .sl(n214), .d1(n210) );
    mux2i_1 U115 ( .x(\data[11] ), .d0(n209), .sl(n214), .d1(n208) );
    mux2i_1 U116 ( .x(\data[12] ), .d0(n207), .sl(n214), .d1(n206) );
    mux2i_1 U117 ( .x(\data[13] ), .d0(n205), .sl(n214), .d1(n204) );
    mux2i_1 U118 ( .x(\data[14] ), .d0(n63), .sl(n214), .d1(n203) );
    mux2i_1 U119 ( .x(\data[15] ), .d0(n202), .sl(n214), .d1(n201) );
    mux2i_1 U120 ( .x(\data[1] ), .d0(n97), .sl(n65), .d1(n221) );
    mux2i_1 U121 ( .x(\data[2] ), .d0(n95), .sl(n65), .d1(n220) );
    mux2i_1 U122 ( .x(\data[3] ), .d0(n93), .sl(n65), .d1(n219) );
    mux2i_1 U123 ( .x(\data[4] ), .d0(n91), .sl(n65), .d1(n218) );
    mux2i_1 U124 ( .x(\data[5] ), .d0(n89), .sl(n65), .d1(n217) );
    mux2i_1 U125 ( .x(\data[6] ), .d0(n87), .sl(n65), .d1(n216) );
    mux2i_1 U126 ( .x(\data[7] ), .d0(n85), .sl(n65), .d1(n215) );
    mux2i_1 U127 ( .x(\data[8] ), .d0(n200), .sl(n214), .d1(n199) );
    mux2i_1 U128 ( .x(\data[9] ), .d0(n198), .sl(n214), .d1(n197) );
    nor2_1 U129 ( .x(high_ir_rd), .a(n79), .b(n80) );
    mux2i_1 U131 ( .x(\size[0] ), .d0(n212), .sl(n65), .d1(n213) );
    nand2i_1 U132 ( .x(n308), .a(sel_o[1]), .b(n70) );
    inv_1 U133 ( .x(n255), .a(n182) );
    inv_1 U134 ( .x(n256), .a(n179) );
    inv_1 U135 ( .x(n257), .a(n176) );
    inv_1 U136 ( .x(n258), .a(n173) );
    inv_1 U137 ( .x(n260), .a(n194) );
    inv_1 U138 ( .x(n261), .a(n191) );
    inv_1 U139 ( .x(n262), .a(n188) );
    inv_1 U140 ( .x(n263), .a(n185) );
    inv_1 U141 ( .x(n245), .a(n158) );
    inv_1 U142 ( .x(n246), .a(n155) );
    inv_1 U143 ( .x(n247), .a(n152) );
    inv_1 U144 ( .x(n248), .a(n149) );
    inv_1 U145 ( .x(n250), .a(n170) );
    inv_1 U146 ( .x(n251), .a(n167) );
    inv_1 U147 ( .x(n252), .a(n164) );
    inv_1 U148 ( .x(n253), .a(n161) );
    inv_1 U149 ( .x(n235), .a(n134) );
    inv_1 U150 ( .x(n236), .a(n131) );
    inv_1 U151 ( .x(n237), .a(n128) );
    inv_1 U152 ( .x(n238), .a(n125) );
    inv_1 U153 ( .x(n240), .a(n146) );
    inv_1 U154 ( .x(n241), .a(n143) );
    inv_1 U155 ( .x(n242), .a(n140) );
    inv_1 U156 ( .x(n243), .a(n137) );
    inv_1 U157 ( .x(n225), .a(n110) );
    inv_1 U158 ( .x(n226), .a(n107) );
    inv_1 U159 ( .x(n227), .a(n104) );
    inv_1 U160 ( .x(n228), .a(n101) );
    inv_1 U161 ( .x(n230), .a(n122) );
    inv_1 U162 ( .x(n231), .a(n119) );
    inv_1 U163 ( .x(n232), .a(n116) );
    inv_1 U164 ( .x(n233), .a(n113) );
    nor2_1 U165 ( .x(n272), .a(n252), .b(n253) );
    nor2_1 U166 ( .x(n271), .a(n250), .b(n251) );
    nor2_1 U167 ( .x(n275), .a(n247), .b(n248) );
    nor2_1 U168 ( .x(n274), .a(n245), .b(n246) );
    nor2_1 U169 ( .x(n265), .a(n262), .b(n263) );
    nor2_1 U170 ( .x(n264), .a(n260), .b(n261) );
    nor2_1 U171 ( .x(n268), .a(n257), .b(n258) );
    nor2_1 U172 ( .x(n267), .a(n255), .b(n256) );
    nor2_1 U173 ( .x(n286), .a(n232), .b(n233) );
    nor2_1 U174 ( .x(n285), .a(n230), .b(n231) );
    nor2_1 U175 ( .x(n289), .a(n227), .b(n228) );
    nor2_1 U176 ( .x(n288), .a(n225), .b(n226) );
    nor2_1 U177 ( .x(n279), .a(n242), .b(n243) );
    nor2_1 U178 ( .x(n278), .a(n240), .b(n241) );
    nor2_1 U179 ( .x(n282), .a(n237), .b(n238) );
    nor2_1 U180 ( .x(n281), .a(n235), .b(n236) );
    nand2_1 U181 ( .x(n182), .a(n183), .b(n184) );
    nand2_1 U182 ( .x(n179), .a(n180), .b(n181) );
    nand2_1 U183 ( .x(n176), .a(n177), .b(n178) );
    nand2_1 U184 ( .x(n173), .a(n174), .b(n175) );
    nand2_1 U185 ( .x(n194), .a(n195), .b(n196) );
    nand2_1 U186 ( .x(n191), .a(n192), .b(n193) );
    nand2_1 U187 ( .x(n188), .a(n189), .b(n190) );
    nand2_1 U188 ( .x(n185), .a(n186), .b(n187) );
    nand2_1 U189 ( .x(n158), .a(n159), .b(n160) );
    nand2_1 U190 ( .x(n155), .a(n156), .b(n157) );
    nand2_1 U191 ( .x(n152), .a(n153), .b(n154) );
    nand2_1 U192 ( .x(n149), .a(n150), .b(n151) );
    nand2_1 U193 ( .x(n170), .a(n171), .b(n172) );
    nand2_1 U194 ( .x(n167), .a(n168), .b(n169) );
    nand2_1 U195 ( .x(n164), .a(n165), .b(n166) );
    nand2_1 U196 ( .x(n161), .a(n162), .b(n163) );
    nand2_1 U197 ( .x(n134), .a(n135), .b(n136) );
    nand2_1 U198 ( .x(n131), .a(n132), .b(n133) );
    nand2_1 U199 ( .x(n128), .a(n129), .b(n130) );
    nand2_1 U200 ( .x(n125), .a(n126), .b(n127) );
    nand2_1 U201 ( .x(n146), .a(n147), .b(n148) );
    nand2_1 U202 ( .x(n143), .a(n144), .b(n145) );
    nand2_1 U203 ( .x(n140), .a(n141), .b(n142) );
    nand2_1 U204 ( .x(n137), .a(n138), .b(n139) );
    nand2_1 U205 ( .x(n110), .a(n111), .b(n112) );
    nand2_1 U206 ( .x(n107), .a(n108), .b(n109) );
    nand2_1 U207 ( .x(n104), .a(n105), .b(n106) );
    nand2_1 U208 ( .x(n101), .a(n102), .b(n103) );
    nand2_1 U209 ( .x(n122), .a(n123), .b(n124) );
    nand2_1 U210 ( .x(n119), .a(n120), .b(n121) );
    nand2_1 U211 ( .x(n116), .a(n117), .b(n118) );
    nand2_1 U212 ( .x(n113), .a(n114), .b(n115) );
    inv_1 U213 ( .x(n183), .a(ir_rd[60]) );
    inv_1 U214 ( .x(n184), .a(ir_rd[28]) );
    inv_1 U215 ( .x(n180), .a(ir_rd[61]) );
    inv_1 U216 ( .x(n181), .a(ir_rd[29]) );
    inv_1 U217 ( .x(n177), .a(ir_rd[62]) );
    inv_1 U218 ( .x(n178), .a(ir_rd[30]) );
    inv_1 U219 ( .x(n174), .a(ir_rd[63]) );
    inv_1 U220 ( .x(n175), .a(ir_rd[31]) );
    inv_1 U221 ( .x(n195), .a(ir_rd[56]) );
    inv_1 U222 ( .x(n196), .a(ir_rd[24]) );
    inv_1 U223 ( .x(n192), .a(ir_rd[57]) );
    inv_1 U224 ( .x(n193), .a(ir_rd[25]) );
    inv_1 U225 ( .x(n189), .a(ir_rd[58]) );
    inv_1 U226 ( .x(n190), .a(ir_rd[26]) );
    inv_1 U227 ( .x(n186), .a(ir_rd[59]) );
    inv_1 U228 ( .x(n187), .a(ir_rd[27]) );
    inv_1 U229 ( .x(n159), .a(ir_rd[52]) );
    inv_1 U230 ( .x(n160), .a(ir_rd[20]) );
    inv_1 U231 ( .x(n156), .a(ir_rd[53]) );
    inv_1 U232 ( .x(n157), .a(ir_rd[21]) );
    inv_1 U233 ( .x(n153), .a(ir_rd[54]) );
    inv_1 U234 ( .x(n154), .a(ir_rd[22]) );
    inv_1 U235 ( .x(n150), .a(ir_rd[55]) );
    inv_1 U236 ( .x(n151), .a(ir_rd[23]) );
    inv_1 U237 ( .x(n171), .a(ir_rd[48]) );
    inv_1 U238 ( .x(n172), .a(ir_rd[16]) );
    inv_1 U239 ( .x(n168), .a(ir_rd[49]) );
    inv_1 U240 ( .x(n169), .a(ir_rd[17]) );
    inv_1 U241 ( .x(n165), .a(ir_rd[50]) );
    inv_1 U242 ( .x(n166), .a(ir_rd[18]) );
    inv_1 U243 ( .x(n162), .a(ir_rd[51]) );
    inv_1 U244 ( .x(n163), .a(ir_rd[19]) );
    inv_1 U245 ( .x(n135), .a(ir_rd[44]) );
    inv_1 U246 ( .x(n136), .a(ir_rd[12]) );
    inv_1 U247 ( .x(n132), .a(ir_rd[45]) );
    inv_1 U248 ( .x(n133), .a(ir_rd[13]) );
    inv_1 U249 ( .x(n129), .a(ir_rd[46]) );
    inv_1 U250 ( .x(n130), .a(ir_rd[14]) );
    inv_1 U251 ( .x(n126), .a(ir_rd[47]) );
    inv_1 U252 ( .x(n127), .a(ir_rd[15]) );
    inv_1 U253 ( .x(n147), .a(ir_rd[40]) );
    inv_1 U254 ( .x(n148), .a(ir_rd[8]) );
    inv_1 U255 ( .x(n144), .a(ir_rd[41]) );
    inv_1 U256 ( .x(n145), .a(ir_rd[9]) );
    inv_1 U257 ( .x(n141), .a(ir_rd[42]) );
    inv_1 U258 ( .x(n142), .a(ir_rd[10]) );
    inv_1 U259 ( .x(n138), .a(ir_rd[43]) );
    inv_1 U260 ( .x(n139), .a(ir_rd[11]) );
    inv_1 U261 ( .x(n111), .a(ir_rd[36]) );
    inv_1 U262 ( .x(n108), .a(ir_rd[37]) );
    inv_1 U263 ( .x(n109), .a(ir_rd[5]) );
    inv_1 U264 ( .x(n105), .a(ir_rd[38]) );
    inv_1 U265 ( .x(n106), .a(ir_rd[6]) );
    inv_1 U266 ( .x(n102), .a(ir_rd[39]) );
    inv_1 U267 ( .x(n103), .a(ir_rd[7]) );
    inv_1 U268 ( .x(n123), .a(ir_rd[32]) );
    inv_1 U269 ( .x(n120), .a(ir_rd[33]) );
    inv_1 U270 ( .x(n121), .a(ir_rd[1]) );
    inv_1 U271 ( .x(n117), .a(ir_rd[34]) );
    inv_1 U272 ( .x(n114), .a(ir_rd[35]) );
    inv_1 U273 ( .x(n115), .a(ir_rd[3]) );
    latn_1 \dat_i_reg[30]  ( .q(dat_i[30]), .d(ir_rd[62]), .g(n7) );
    latn_1 \dat_i_reg[28]  ( .q(dat_i[28]), .d(ir_rd[60]), .g(n7) );
    latn_1 \dat_i_reg[27]  ( .q(dat_i[27]), .d(ir_rd[59]), .g(n7) );
    latn_1 \dat_i_reg[26]  ( .q(dat_i[26]), .d(ir_rd[58]), .g(n7) );
    latn_1 \dat_i_reg[25]  ( .q(dat_i[25]), .d(ir_rd[57]), .g(n7) );
    latn_1 \dat_i_reg[24]  ( .q(dat_i[24]), .d(ir_rd[56]), .g(n7) );
    latn_1 \dat_i_reg[22]  ( .q(dat_i[22]), .d(ir_rd[54]), .g(n7) );
    latn_1 \dat_i_reg[20]  ( .q(dat_i[20]), .d(ir_rd[52]), .g(n7) );
    latn_1 \dat_i_reg[19]  ( .q(dat_i[19]), .d(ir_rd[51]), .g(n7) );
    latn_1 \dat_i_reg[18]  ( .q(dat_i[18]), .d(ir_rd[50]), .g(n7) );
    latn_1 \dat_i_reg[17]  ( .q(dat_i[17]), .d(ir_rd[49]), .g(n7) );
    latn_1 \dat_i_reg[16]  ( .q(dat_i[16]), .d(ir_rd[48]), .g(n6) );
    latn_1 \dat_i_reg[14]  ( .q(dat_i[14]), .d(ir_rd[46]), .g(n6) );
    latn_1 \dat_i_reg[12]  ( .q(dat_i[12]), .d(ir_rd[44]), .g(n6) );
    latn_1 \dat_i_reg[10]  ( .q(dat_i[10]), .d(ir_rd[42]), .g(n6) );
    latn_1 \dat_i_reg[8]  ( .q(dat_i[8]), .d(ir_rd[40]), .g(n6) );
    latn_1 \dat_i_reg[6]  ( .q(dat_i[6]), .d(ir_rd[38]), .g(n6) );
    latn_1 \dat_i_reg[4]  ( .q(dat_i[4]), .d(ir_rd[36]), .g(n6) );
    latn_1 \dat_i_reg[3]  ( .q(dat_i[3]), .d(ir_rd[35]), .g(n1) );
    latn_1 \dat_i_reg[2]  ( .q(dat_i[2]), .d(ir_rd[34]), .g(n1) );
    latn_1 \dat_i_reg[1]  ( .q(dat_i[1]), .d(ir_rd[33]), .g(n1) );
    latn_1 \dat_i_reg[0]  ( .q(dat_i[0]), .d(ir_rd[32]), .g(n1) );
    latn_1 we_i_reg ( .q(we_i), .d(ir_rnw[0]), .g(n1) );
    latn_1 err_i_reg ( .q(err_i), .d(ir_err[1]), .g(n1) );
    latn_1 \dat_i_reg[13]  ( .q(dat_i[13]), .d(ir_rd[45]), .g(n6) );
    latn_1 \dat_i_reg[5]  ( .q(dat_i[5]), .d(ir_rd[37]), .g(n1) );
    latn_1 \dat_i_reg[15]  ( .q(dat_i[15]), .d(ir_rd[47]), .g(n6) );
    latn_1 \dat_i_reg[7]  ( .q(dat_i[7]), .d(ir_rd[39]), .g(n1) );
    latn_1 \dat_i_reg[29]  ( .q(dat_i[29]), .d(ir_rd[61]), .g(n6) );
    latn_1 \dat_i_reg[21]  ( .q(dat_i[21]), .d(ir_rd[53]), .g(n1) );
    latn_1 \dat_i_reg[31]  ( .q(dat_i[31]), .d(ir_rd[63]), .g(n6) );
    latn_1 \dat_i_reg[23]  ( .q(dat_i[23]), .d(ir_rd[55]), .g(n1) );
    latn_1 \dat_i_reg[9]  ( .q(dat_i[9]), .d(ir_rd[41]), .g(n6) );
    latn_1 \dat_i_reg[11]  ( .q(dat_i[11]), .d(ir_rd[43]), .g(n1) );
    oa21_1 \all_write/__tmp99/U1  ( .x(all_w), .a(_28_net_), .b(all_w), .c(
        comp_basic) );
    ao31_1 \all_read/__tmp99/aoi  ( .x(\all_read/__tmp99/loop ), .a(comp_basic
        ), .b(comp_rd), .c(_27_net_), .d(all_r) );
    oa21_1 \all_read/__tmp99/outGate  ( .x(all_r), .a(comp_basic), .b(comp_rd), 
        .c(\all_read/__tmp99/loop ) );
    ao222_1 \rd/__tmp99/U1  ( .x(comp_rd), .a(high_ir_rd), .b(low_ir_rd), .c(
        high_ir_rd), .d(comp_rd), .e(low_ir_rd), .f(comp_rd) );
    ao222_1 \basic/__tmp99/U1  ( .x(comp_basic), .a(_25_net_), .b(_26_net_), 
        .c(_25_net_), .d(comp_basic), .e(_26_net_), .f(comp_basic) );
    inv_1 \Ucol2/Uii  ( .x(\Ucol2/ni ), .a(ts_o[2]) );
    inv_1 \Ucol2/Uih  ( .x(\Ucol2/nh ), .a(ic_col[5]) );
    inv_1 \Ucol2/Uil  ( .x(\Ucol2/nl ), .a(ic_col[2]) );
    ao23_1 \Ucol2/Ucl/U1/U1  ( .x(ic_col[2]), .a(n11), .b(ic_col[2]), .c(n8), 
        .d(\Ucol2/ni ), .e(\Ucol2/nh ) );
    ao23_1 \Ucol2/Uch/U1/U1  ( .x(ic_col[5]), .a(n11), .b(ic_col[5]), .c(n8), 
        .d(ts_o[2]), .e(\Ucol2/nl ) );
    inv_1 \Ucol1/Uii  ( .x(\Ucol1/ni ), .a(ts_o[1]) );
    inv_1 \Ucol1/Uih  ( .x(\Ucol1/nh ), .a(ic_col[4]) );
    inv_1 \Ucol1/Uil  ( .x(\Ucol1/nl ), .a(ic_col[1]) );
    ao23_1 \Ucol1/Ucl/U1/U1  ( .x(ic_col[1]), .a(n11), .b(ic_col[1]), .c(n8), 
        .d(\Ucol1/ni ), .e(\Ucol1/nh ) );
    ao23_1 \Ucol1/Uch/U1/U1  ( .x(ic_col[4]), .a(n11), .b(ic_col[4]), .c(n9), 
        .d(ts_o[1]), .e(\Ucol1/nl ) );
    inv_1 \Ucol0/Uii  ( .x(\Ucol0/ni ), .a(ts_o[0]) );
    inv_1 \Ucol0/Uih  ( .x(\Ucol0/nh ), .a(ic_col[3]) );
    inv_1 \Ucol0/Uil  ( .x(\Ucol0/nl ), .a(ic_col[0]) );
    ao23_1 \Ucol0/Ucl/U1/U1  ( .x(ic_col[0]), .a(n11), .b(ic_col[0]), .c(n10), 
        .d(\Ucol0/ni ), .e(\Ucol0/nh ) );
    ao23_1 \Ucol0/Uch/U1/U1  ( .x(ic_col[3]), .a(n11), .b(ic_col[3]), .c(n9), 
        .d(ts_o[0]), .e(\Ucol0/nl ) );
    inv_1 \Utag4/Uii  ( .x(\Utag4/ni ), .a(tag_id[4]) );
    inv_1 \Utag4/Uih  ( .x(\Utag4/nh ), .a(ic_itag[9]) );
    inv_1 \Utag4/Uil  ( .x(\Utag4/nl ), .a(ic_itag[4]) );
    ao23_1 \Utag4/Ucl/U1/U1  ( .x(ic_itag[4]), .a(n11), .b(ic_itag[4]), .c(n9), 
        .d(\Utag4/ni ), .e(\Utag4/nh ) );
    ao23_1 \Utag4/Uch/U1/U1  ( .x(ic_itag[9]), .a(n10), .b(ic_itag[9]), .c(n9), 
        .d(tag_id[4]), .e(\Utag4/nl ) );
    inv_1 \Utag3/Uii  ( .x(\Utag3/ni ), .a(tag_id[3]) );
    inv_1 \Utag3/Uih  ( .x(\Utag3/nh ), .a(ic_itag[8]) );
    inv_1 \Utag3/Uil  ( .x(\Utag3/nl ), .a(ic_itag[3]) );
    ao23_1 \Utag3/Ucl/U1/U1  ( .x(ic_itag[3]), .a(n10), .b(ic_itag[3]), .c(n9), 
        .d(\Utag3/ni ), .e(\Utag3/nh ) );
    ao23_1 \Utag3/Uch/U1/U1  ( .x(ic_itag[8]), .a(n10), .b(ic_itag[8]), .c(n9), 
        .d(tag_id[3]), .e(\Utag3/nl ) );
    inv_1 \Utag2/Uii  ( .x(\Utag2/ni ), .a(tag_id[2]) );
    inv_1 \Utag2/Uih  ( .x(\Utag2/nh ), .a(ic_itag[7]) );
    inv_1 \Utag2/Uil  ( .x(\Utag2/nl ), .a(ic_itag[2]) );
    ao23_1 \Utag2/Ucl/U1/U1  ( .x(ic_itag[2]), .a(n10), .b(ic_itag[2]), .c(n9), 
        .d(\Utag2/ni ), .e(\Utag2/nh ) );
    ao23_1 \Utag2/Uch/U1/U1  ( .x(ic_itag[7]), .a(n10), .b(ic_itag[7]), .c(n10
        ), .d(tag_id[2]), .e(\Utag2/nl ) );
    inv_1 \Utag1/Uii  ( .x(\Utag1/ni ), .a(tag_id[1]) );
    inv_1 \Utag1/Uih  ( .x(\Utag1/nh ), .a(ic_itag[6]) );
    inv_1 \Utag1/Uil  ( .x(\Utag1/nl ), .a(ic_itag[1]) );
    ao23_1 \Utag1/Ucl/U1/U1  ( .x(ic_itag[1]), .a(n11), .b(ic_itag[1]), .c(n9), 
        .d(\Utag1/ni ), .e(\Utag1/nh ) );
    ao23_1 \Utag1/Uch/U1/U1  ( .x(ic_itag[6]), .a(n11), .b(ic_itag[6]), .c(n9), 
        .d(tag_id[1]), .e(\Utag1/nl ) );
    inv_1 \Utag0/Uii  ( .x(\Utag0/ni ), .a(tag_id[0]) );
    inv_1 \Utag0/Uih  ( .x(\Utag0/nh ), .a(ic_itag[5]) );
    inv_1 \Utag0/Uil  ( .x(\Utag0/nl ), .a(ic_itag[0]) );
    ao23_1 \Utag0/Ucl/U1/U1  ( .x(ic_itag[0]), .a(n11), .b(ic_itag[0]), .c(n8), 
        .d(\Utag0/ni ), .e(\Utag0/nh ) );
    ao23_1 \Utag0/Uch/U1/U1  ( .x(ic_itag[5]), .a(n10), .b(ic_itag[5]), .c(n8), 
        .d(tag_id[0]), .e(\Utag0/nl ) );
    inv_1 \Usze1/Uii  ( .x(\Usze1/ni ), .a(\size[1] ) );
    inv_1 \Usze1/Uih  ( .x(\Usze1/nh ), .a(ic_size[3]) );
    inv_1 \Usze1/Uil  ( .x(\Usze1/nl ), .a(ic_size[1]) );
    ao23_1 \Usze1/Ucl/U1/U1  ( .x(ic_size[1]), .a(n10), .b(ic_size[1]), .c(n9), 
        .d(\Usze1/ni ), .e(\Usze1/nh ) );
    ao23_1 \Usze1/Uch/U1/U1  ( .x(ic_size[3]), .a(n10), .b(ic_size[3]), .c(n9), 
        .d(\size[1] ), .e(\Usze1/nl ) );
    inv_1 \Usze0/Uii  ( .x(\Usze0/ni ), .a(\size[0] ) );
    inv_1 \Usze0/Uih  ( .x(\Usze0/nh ), .a(ic_size[2]) );
    inv_1 \Usze0/Uil  ( .x(\Usze0/nl ), .a(ic_size[0]) );
    ao23_1 \Usze0/Ucl/U1/U1  ( .x(ic_size[0]), .a(n10), .b(ic_size[0]), .c(n9), 
        .d(\Usze0/ni ), .e(\Usze0/nh ) );
    ao23_1 \Usze0/Uch/U1/U1  ( .x(ic_size[2]), .a(n10), .b(ic_size[2]), .c(n9), 
        .d(\size[0] ), .e(\Usze0/nl ) );
    inv_1 \Urnw/Uii  ( .x(\Urnw/ni ), .a(_24_net_) );
    inv_1 \Urnw/Uih  ( .x(\Urnw/nh ), .a(ic_rnw[1]) );
    inv_1 \Urnw/Uil  ( .x(\Urnw/nl ), .a(ic_rnw[0]) );
    ao23_1 \Urnw/Ucl/U1/U1  ( .x(ic_rnw[0]), .a(n10), .b(ic_rnw[0]), .c(n9), 
        .d(\Urnw/ni ), .e(\Urnw/nh ) );
    ao23_1 \Urnw/Uch/U1/U1  ( .x(ic_rnw[1]), .a(n10), .b(ic_rnw[1]), .c(n9), 
        .d(_24_net_), .e(\Urnw/nl ) );
    inv_1 \Ulock/Uii  ( .x(\Ulock/ni ), .a(mult_o) );
    inv_1 \Ulock/Uih  ( .x(\Ulock/nh ), .a(ic_lock[1]) );
    inv_1 \Ulock/Uil  ( .x(\Ulock/nl ), .a(ic_lock[0]) );
    ao23_1 \Ulock/Ucl/U1/U1  ( .x(ic_lock[0]), .a(n11), .b(ic_lock[0]), .c(n9), 
        .d(\Ulock/ni ), .e(\Ulock/nh ) );
    ao23_1 \Ulock/Uch/U1/U1  ( .x(ic_lock[1]), .a(n11), .b(ic_lock[1]), .c(n8), 
        .d(mult_o), .e(\Ulock/nl ) );
    inv_1 \Upred/Uii  ( .x(\Upred/ni ), .a(prd_o) );
    inv_1 \Upred/Uih  ( .x(\Upred/nh ), .a(ic_pred[1]) );
    inv_1 \Upred/Uil  ( .x(\Upred/nl ), .a(ic_pred[0]) );
    ao23_1 \Upred/Ucl/U1/U1  ( .x(ic_pred[0]), .a(n11), .b(ic_pred[0]), .c(n8), 
        .d(\Upred/ni ), .e(\Upred/nh ) );
    ao23_1 \Upred/Uch/U1/U1  ( .x(ic_pred[1]), .a(n10), .b(ic_pred[1]), .c(n8), 
        .d(prd_o), .e(\Upred/nl ) );
    inv_1 \Useq/Uii  ( .x(\Useq/ni ), .a(seq_o) );
    inv_1 \Useq/Uih  ( .x(\Useq/nh ), .a(ic_seq[1]) );
    inv_1 \Useq/Uil  ( .x(\Useq/nl ), .a(ic_seq[0]) );
    ao23_1 \Useq/Ucl/U1/U1  ( .x(ic_seq[0]), .a(n10), .b(ic_seq[0]), .c(n8), 
        .d(\Useq/ni ), .e(\Useq/nh ) );
    ao23_1 \Useq/Uch/U1/U1  ( .x(ic_seq[1]), .a(n11), .b(ic_seq[1]), .c(n8), 
        .d(seq_o), .e(\Useq/nl ) );
    buf_3 U1 ( .x(n1), .a(en) );
    buf_3 U41 ( .x(n7), .a(en) );
    buf_3 U43 ( .x(n6), .a(en) );
    inv_2 U44 ( .x(n214), .a(n308) );
    buf_3 U47 ( .x(n65), .a(sel_o[0]) );
    nand3i_0 U48 ( .x(n212), .a(sel_o[1]), .b(sel_o[3]), .c(n70) );
    nor2_0 U49 ( .x(n223), .a(n70), .b(sel_o[3]) );
    nand2_0 U50 ( .x(n297), .a(dat_o[29]), .b(sel_o[3]) );
    nand2_0 U58 ( .x(n301), .a(dat_o[27]), .b(sel_o[3]) );
    nand2_0 U59 ( .x(n299), .a(dat_o[28]), .b(sel_o[3]) );
    nand2_0 U102 ( .x(n83), .a(n70), .b(sel_o[3]) );
    inv_0 U106 ( .x(n78), .a(ir_err[0]) );
    nand2i_0 U107 ( .x(_28_net_), .a(ir_err[1]), .b(n72) );
    nand2i_0 U108 ( .x(_25_net_), .a(ir_err[1]), .b(n78) );
    buf_16 U112 ( .x(n8), .a(req_in_delayed) );
    buf_16 U279 ( .x(n9), .a(req_in_delayed) );
    buf_16 U280 ( .x(n10), .a(req_in_delayed) );
    buf_16 U281 ( .x(n11), .a(req_in_delayed) );
endmodule


module i_adec_iport ( e_h, e_l, r_h, r_l, ah, al, e_bare, e_dm, e_im, e_wish, 
    r_bare, r_dm, r_im, r_wish, force_bare );
output [3:0] e_h;
output [3:0] e_l;
output [3:0] r_h;
output [3:0] r_l;
input  [31:0] ah;
input  [31:0] al;
input  [3:0] e_bare;
input  [3:0] e_dm;
input  [3:0] e_im;
input  [3:0] e_wish;
input  [3:0] r_bare;
input  [3:0] r_dm;
input  [3:0] r_im;
input  [3:0] r_wish;
input  force_bare;
    wire e_h_0, e_l_3, e_l_2, e_l_0, wish_i, n6, bare_i, im_i, n7, dm_i, 
        \r_l[2] , \r_l[0] , n1, n2, n3, n15, n14, n12;
    assign e_h[3] = 1'b0;
    assign e_h[0] = e_h_0;
    assign e_l[3] = e_l_3;
    assign e_l[2] = e_l_2;
    assign e_l[0] = e_l_0;
    assign r_h[3] = e_l_2;
    assign r_h[2] = e_h_0;
    assign r_h[0] = 1'b0;
    assign r_l[2] = e_l_0;
    assign r_l[0] = e_l_3;
    ao222_1 \U1632/U18/U1/U1  ( .x(wish_i), .a(n6), .b(al[30]), .c(n6), .d(
        wish_i), .e(al[30]), .f(wish_i) );
    ao222_1 \U1633/U18/U1/U1  ( .x(bare_i), .a(n6), .b(ah[30]), .c(n6), .d(
        bare_i), .e(ah[30]), .f(bare_i) );
    ao222_1 \U1634/U18/U1/U1  ( .x(im_i), .a(al[11]), .b(n7), .c(al[11]), .d(
        im_i), .e(n7), .f(im_i) );
    ao222_1 \U1635/U18/U1/U1  ( .x(dm_i), .a(ah[11]), .b(n7), .c(ah[11]), .d(
        dm_i), .e(n7), .f(dm_i) );
    or3_1 U1 ( .x(\r_l[2] ), .a(wish_i), .b(bare_i), .c(force_bare) );
    or2_1 U2 ( .x(r_l[1]), .a(e_l_0), .b(im_i) );
    or2_1 U3 ( .x(\r_l[0] ), .a(dm_i), .b(r_l[1]) );
    nor2_0 U4 ( .x(n1), .a(bare_i), .b(force_bare) );
    aoi21_1 U6 ( .x(n2), .a(n3), .b(im_i), .c(r_h[1]) );
    inv_0 U8 ( .x(n3), .a(force_bare) );
    nor2i_0 U9 ( .x(n15), .a(wish_i), .b(force_bare) );
    nor2i_0 U10 ( .x(n14), .a(dm_i), .b(force_bare) );
    inv_0 U11 ( .x(e_h[1]), .a(n1) );
    buf_1 U15 ( .x(n6), .a(ah[31]) );
    buf_1 U16 ( .x(n7), .a(al[31]) );
    nand2_2 U17 ( .x(e_l_2), .a(n2), .b(n1) );
    buf_1 U18 ( .x(r_h[1]), .a(n14) );
    inv_2 U19 ( .x(e_h_0), .a(n2) );
    buf_3 U20 ( .x(e_l_3), .a(\r_l[0] ) );
    buf_3 U21 ( .x(e_l_0), .a(\r_l[2] ) );
    nand2i_2 U22 ( .x(e_l[1]), .a(n12), .b(n2) );
    buf_1 U23 ( .x(e_h[2]), .a(n15) );
    buf_1 U24 ( .x(r_l[3]), .a(n15) );
    buf_1 U25 ( .x(n12), .a(n15) );
endmodule


module chain_selement_ga_4 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_symbol_0 ( o, txack, txack_last, e, oa, r, txreq );
output [2:0] o;
input  [1:0] e;
input  [1:0] r;
input  oa, txreq;
output txack, txack_last;
    wire ack, net10, \c[0] , \c[1] ;
    chain_selement_ga_4 U1239 ( .Aa(ack), .Br(net10), .Ar(txreq), .Ba(oa) );
    and2_1 \U1229_0_/U8  ( .x(o[0]), .a(\c[0] ), .b(net10) );
    and2_1 \U1229_1_/U8  ( .x(o[1]), .a(\c[1] ), .b(net10) );
    and2_1 \U1229_2_/U8  ( .x(o[2]), .a(e[1]), .b(net10) );
    ao23_1 \U1251/U19/U21/U1/U1  ( .x(txack_last), .a(ack), .b(txack_last), 
        .c(ack), .d(e[1]), .e(e[1]) );
    ao23_1 \U1250/U19/U21/U1/U1  ( .x(txack), .a(ack), .b(txack), .c(ack), .d(
        e[0]), .e(e[0]) );
    ao222_1 \U1210/U18/U1/U1  ( .x(\c[0] ), .a(e[0]), .b(r[0]), .c(e[0]), .d(
        \c[0] ), .e(r[0]), .f(\c[0] ) );
    ao222_1 \U1209/U18/U1/U1  ( .x(\c[1] ), .a(e[0]), .b(r[1]), .c(e[0]), .d(
        \c[1] ), .e(r[1]), .f(\c[1] ) );
endmodule


module chain_selement_ga_5 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_symbol_1 ( o, txack, txack_last, e, oa, r, txreq );
output [2:0] o;
input  [1:0] e;
input  [1:0] r;
input  oa, txreq;
output txack, txack_last;
    wire ack, net10, \c[0] , \c[1] ;
    chain_selement_ga_5 U1239 ( .Aa(ack), .Br(net10), .Ar(txreq), .Ba(oa) );
    and2_1 \U1229_0_/U8  ( .x(o[0]), .a(\c[0] ), .b(net10) );
    and2_1 \U1229_1_/U8  ( .x(o[1]), .a(\c[1] ), .b(net10) );
    and2_1 \U1229_2_/U8  ( .x(o[2]), .a(e[1]), .b(net10) );
    ao23_1 \U1251/U19/U21/U1/U1  ( .x(txack_last), .a(ack), .b(txack_last), 
        .c(ack), .d(e[1]), .e(e[1]) );
    ao23_1 \U1250/U19/U21/U1/U1  ( .x(txack), .a(ack), .b(txack), .c(ack), .d(
        e[0]), .e(e[0]) );
    ao222_1 \U1210/U18/U1/U1  ( .x(\c[0] ), .a(e[0]), .b(r[0]), .c(e[0]), .d(
        \c[0] ), .e(r[0]), .f(\c[0] ) );
    ao222_1 \U1209/U18/U1/U1  ( .x(\c[1] ), .a(e[0]), .b(r[1]), .c(e[0]), .d(
        \c[1] ), .e(r[1]), .f(\c[1] ) );
endmodule


module chain_selement_ga_6 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_symbol_2 ( o, txack, txack_last, e, oa, r, txreq );
output [2:0] o;
input  [1:0] e;
input  [1:0] r;
input  oa, txreq;
output txack, txack_last;
    wire ack, net10, \c[0] , \c[1] ;
    chain_selement_ga_6 U1239 ( .Aa(ack), .Br(net10), .Ar(txreq), .Ba(oa) );
    and2_1 \U1229_0_/U8  ( .x(o[0]), .a(\c[0] ), .b(net10) );
    and2_1 \U1229_1_/U8  ( .x(o[1]), .a(\c[1] ), .b(net10) );
    and2_1 \U1229_2_/U8  ( .x(o[2]), .a(e[1]), .b(net10) );
    ao23_1 \U1251/U19/U21/U1/U1  ( .x(txack_last), .a(ack), .b(txack_last), 
        .c(ack), .d(e[1]), .e(e[1]) );
    ao23_1 \U1250/U19/U21/U1/U1  ( .x(txack), .a(ack), .b(txack), .c(ack), .d(
        e[0]), .e(e[0]) );
    ao222_1 \U1210/U18/U1/U1  ( .x(\c[0] ), .a(e[0]), .b(r[0]), .c(e[0]), .d(
        \c[0] ), .e(r[0]), .f(\c[0] ) );
    ao222_1 \U1209/U18/U1/U1  ( .x(\c[1] ), .a(e[0]), .b(r[1]), .c(e[0]), .d(
        \c[1] ), .e(r[1]), .f(\c[1] ) );
endmodule


module chain_selement_ga_7 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_symbol_3 ( o, txack, txack_last, e, oa, r, txreq );
output [2:0] o;
input  [1:0] e;
input  [1:0] r;
input  oa, txreq;
output txack, txack_last;
    wire ack, net10, \c[0] , \c[1] ;
    chain_selement_ga_7 U1239 ( .Aa(ack), .Br(net10), .Ar(txreq), .Ba(oa) );
    and2_1 \U1229_0_/U8  ( .x(o[0]), .a(\c[0] ), .b(net10) );
    and2_1 \U1229_1_/U8  ( .x(o[1]), .a(\c[1] ), .b(net10) );
    and2_1 \U1229_2_/U8  ( .x(o[2]), .a(e[1]), .b(net10) );
    ao23_1 \U1251/U19/U21/U1/U1  ( .x(txack_last), .a(ack), .b(txack_last), 
        .c(ack), .d(e[1]), .e(e[1]) );
    ao23_1 \U1250/U19/U21/U1/U1  ( .x(txack), .a(ack), .b(txack), .c(ack), .d(
        e[0]), .e(e[0]) );
    ao222_1 \U1210/U18/U1/U1  ( .x(\c[0] ), .a(e[0]), .b(r[0]), .c(e[0]), .d(
        \c[0] ), .e(r[0]), .f(\c[0] ) );
    ao222_1 \U1209/U18/U1/U1  ( .x(\c[1] ), .a(e[0]), .b(r[1]), .c(e[0]), .d(
        \c[1] ), .e(r[1]), .f(\c[1] ) );
endmodule


module chain_selement_ga_77 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_tx_iport ( o, rtxack, e_h, e_l, noa, r_h, r_l, rtxreq );
output [4:0] o;
input  [3:0] e_h;
input  [3:0] e_l;
input  [3:0] r_h;
input  [3:0] r_l;
input  noa, rtxreq;
output rtxack;
    wire net33, \last[4] , net60, \r3[2] , \r3[1] , \r3[0] , net40, \last[3] , 
        \r2[2] , \r2[1] , \r2[0] , net47, \last[2] , \r1[2] , \r1[1] , \r1[0] , 
        net50, \last[1] , \r0[2] , \r0[1] , \r0[0] , \last[0] , eopsym, 
        \I8/nb , \I8/na , \net55[1] , \net55[0] , \net52[1] , \net52[0] , 
        \I11/nc , \I11/nb , \I11/na , net16, net11, net9, net6, 
        \I7_0_/U25/U1/clr , \I7_0_/U25/U1/ob , \I7_1_/U25/U1/clr , 
        \I7_1_/U25/U1/ob ;
    assign o[3] = 1'b0;
    assign o[2] = 1'b0;
    route_symbol_0 I0 ( .o({\r3[2] , \r3[1] , \r3[0] }), .txack(net33), 
        .txack_last(\last[4] ), .e({e_h[3], e_l[3]}), .oa(net60), .r({r_h[3], 
        r_l[3]}), .txreq(rtxreq) );
    route_symbol_1 I1 ( .o({\r2[2] , \r2[1] , \r2[0] }), .txack(net40), 
        .txack_last(\last[3] ), .e({e_h[2], e_l[2]}), .oa(net60), .r({r_h[2], 
        r_l[2]}), .txreq(net33) );
    route_symbol_2 I2 ( .o({\r1[2] , \r1[1] , \r1[0] }), .txack(net47), 
        .txack_last(\last[2] ), .e({e_h[1], e_l[1]}), .oa(net60), .r({r_h[1], 
        r_l[1]}), .txreq(net40) );
    route_symbol_3 I3 ( .o({\r0[2] , \r0[1] , \r0[0] }), .txack(net50), 
        .txack_last(\last[1] ), .e({e_h[0], e_l[0]}), .oa(net60), .r({r_h[0], 
        r_l[0]}), .txreq(net47) );
    chain_selement_ga_77 I9 ( .Aa(\last[0] ), .Br(eopsym), .Ar(net50), .Ba(
        net60) );
    nor3_1 \I8/U27  ( .x(\I8/nb ), .a(o[4]), .b(1'b0), .c(1'b0) );
    nor2_1 \I8/U26  ( .x(\I8/na ), .a(o[1]), .b(o[0]) );
    nand2_2 \I8/U29  ( .x(net60), .a(\I8/nb ), .b(\I8/na ) );
    or2_1 \I13_0_/U12  ( .x(\net55[1] ), .a(\r1[0] ), .b(\r0[0] ) );
    or2_1 \I13_1_/U12  ( .x(\net55[0] ), .a(\r1[1] ), .b(\r0[1] ) );
    or2_1 \I14_0_/U12  ( .x(\net52[1] ), .a(\r3[0] ), .b(\r2[0] ) );
    or2_1 \I14_1_/U12  ( .x(\net52[0] ), .a(\r3[1] ), .b(\r2[1] ) );
    nand3_1 \I11/U31  ( .x(rtxack), .a(\I11/nc ), .b(\I11/nb ), .c(\I11/na )
         );
    inv_1 \I11/U33  ( .x(\I11/nc ), .a(\last[0] ) );
    nor2_1 \I11/U26  ( .x(\I11/na ), .a(\last[3] ), .b(\last[4] ) );
    nor2_1 \I11/U32  ( .x(\I11/nb ), .a(\last[1] ), .b(\last[2] ) );
    nor2_1 \I16/U5  ( .x(net16), .a(\r1[2] ), .b(\r0[2] ) );
    nor2_1 \I5/U5  ( .x(net11), .a(\r3[2] ), .b(\r2[2] ) );
    nand3_1 \I17/U9  ( .x(net9), .a(net6), .b(net11), .c(net16) );
    inv_1 \I18/U3  ( .x(net6), .a(eopsym) );
    oa31_1 \I7_0_/U25/U1/Uclr  ( .x(\I7_0_/U25/U1/clr ), .a(noa), .b(
        \net55[1] ), .c(\net52[1] ), .d(o[0]) );
    oaoi211_1 \I7_0_/U25/U1/Uaoi  ( .x(\I7_0_/U25/U1/ob ), .a(\net55[1] ), .b(
        \net52[1] ), .c(noa), .d(\I7_0_/U25/U1/clr ) );
    inv_2 \I7_0_/U25/U1/Ui  ( .x(o[0]), .a(\I7_0_/U25/U1/ob ) );
    oa31_1 \I7_1_/U25/U1/Uclr  ( .x(\I7_1_/U25/U1/clr ), .a(noa), .b(
        \net55[0] ), .c(\net52[0] ), .d(o[1]) );
    oaoi211_1 \I7_1_/U25/U1/Uaoi  ( .x(\I7_1_/U25/U1/ob ), .a(\net55[0] ), .b(
        \net52[0] ), .c(noa), .d(\I7_1_/U25/U1/clr ) );
    inv_2 \I7_1_/U25/U1/Ui  ( .x(o[1]), .a(\I7_1_/U25/U1/ob ) );
    ao222_1 \I15/U18/U1/U1  ( .x(o[4]), .a(noa), .b(net9), .c(noa), .d(o[4]), 
        .e(net9), .f(o[4]) );
endmodule


module chain_irdemuxNew_0 ( err, ncback, rd, rnw, status, cbh, cbl, nReset, 
    nack, statusack );
output [1:0] err;
output [63:0] rd;
output [1:0] rnw;
output [1:0] status;
input  [7:0] cbh;
input  [7:0] cbl;
input  nReset, nack, statusack;
output ncback;
    wire bpullcd, pullcd, net162, reset, pkt_normal, \opc_l[2] , \opc_l[1] , 
        net150, \opc_h[1] , pkt_done, write, net193, \ncd[0] , \ncd[1] , 
        \ncd[2] , \ncd[3] , \ncd[4] , \ncd[5] , \ncd[6] , \ncd[7] , 
        start_receiving, notify, net176, net86, net172, net173, net171, net169, 
        net170, net168, net166, net167, \U1664/x[3] , \U1664/U28/Z , 
        \U1664/x[0] , \U1664/U32/Z , \U1664/x[2] , \U1664/U29/Z , \U1664/y[0] , 
        \U1664/x[1] , \U1664/U33/Z , \U1664/y[1] , \U1664/U30/Z , 
        \U1664/U31/Z , \U1664/U37/Z , \U1697/U21/nr , net149, \U1697/U21/nd , 
        \U1697/U21/n2 , \U307/U21/nr , \U307/U21/nd , \U307/U21/n2 , 
        \U1698/nr , \U1698/nd , \U1698/n2 , read, n17, \opc_h[0] , n18, 
        \opc_l[0] , net0187, net0208, \I6/latch , \I6/nlocalcd , \I6/localcd , 
        \I6/ncd[0] , \I6/ncd[1] , \I6/ncd[2] , \I6/oh[2] , \I6/ncd[3] , 
        \I6/ol[3] , \I6/oh[3] , \I6/ncd[4] , \I6/ol[4] , \I6/oh[4] , 
        \I6/ncd[5] , \I6/ncd[6] , \I6/ol[6] , \I6/oh[6] , \I6/ncd[7] , 
        \I6/ol[7] , \I6/oh[7] , \I6/ctrlack_internal , \I6/acb , \I6/ba , 
        \I6/driveh , net139, \I6/drivel , n12, n13, \I6/U4/U28/U1/clr , 
        \I6/U4/U28/U1/set , \I6/U1/Z , n14, \I6/U1664/x[3] , \I6/U1664/U28/Z , 
        \I6/U1664/x[0] , \I6/U1664/U32/Z , \I6/U1664/x[2] , \I6/U1664/U29/Z , 
        \I6/U1664/y[0] , \I6/U1664/x[1] , \I6/U1664/U33/Z , \I6/U1664/y[1] , 
        \I6/U1664/U30/Z , \I6/U1664/U31/Z , \I6/U1664/U37/Z , \I6/U1669/nr , 
        \I6/U1669/nd , \I6/U1669/n2 , \U1667/latch , \U1667/nlocalcd , 
        \U1667/localcd , \U1667/ncd[0] , \U1667/ncd[1] , \U1667/ncd[2] , 
        \U1667/ncd[3] , \U1667/ncd[4] , \U1667/ncd[5] , \U1667/ncd[6] , 
        \U1667/ncd[7] , \U1667/ctrlack_internal , \U1667/acb , \U1667/ba , 
        \U1667/driveh , read_lhw, \U1667/drivel , n11, n10, 
        \U1667/U4/U28/U1/clr , \U1667/U4/U28/U1/set , \U1667/U1/Z , 
        \U1667/U1664/x[3] , \U1667/U1664/U28/Z , \U1667/U1664/x[0] , 
        \U1667/U1664/U32/Z , \U1667/U1664/x[2] , \U1667/U1664/U29/Z , 
        \U1667/U1664/y[0] , \U1667/U1664/x[1] , \U1667/U1664/U33/Z , 
        \U1667/U1664/y[1] , \U1667/U1664/U30/Z , \U1667/U1664/U31/Z , 
        \U1667/U1664/U37/Z , \U1667/U1669/nr , \U1667/U1669/nd , 
        \U1667/U1669/n2 , \U1650/latch , \U1650/nlocalcd , \U1650/localcd , 
        \U1650/ncd[0] , \U1650/ol[0] , \U1650/oh[0] , \U1650/ncd[1] , 
        \U1650/ol[1] , \U1650/oh[1] , \U1650/ncd[2] , \U1650/ol[2] , 
        \U1650/oh[2] , \U1650/ncd[3] , \U1650/ol[3] , \U1650/oh[3] , 
        \U1650/ncd[4] , \U1650/ol[4] , \U1650/oh[4] , \U1650/ncd[5] , 
        \col_l[0] , \col_h[0] , \U1650/ncd[6] , \col_l[1] , \col_h[1] , 
        \U1650/ncd[7] , \col_l[2] , \col_h[2] , \U1650/ctrlack_internal , 
        \U1650/acb , \U1650/ba , \U1650/driveh , \U1650/drivel , n7, n9, n8, 
        \U1650/U4/U28/U1/clr , \U1650/U4/U28/U1/set , \U1650/U1/Z , 
        \U1650/U1664/x[3] , \U1650/U1664/U28/Z , \U1650/U1664/x[0] , 
        \U1650/U1664/U32/Z , \U1650/U1664/x[2] , \U1650/U1664/U29/Z , 
        \U1650/U1664/y[0] , \U1650/U1664/x[1] , \U1650/U1664/U33/Z , 
        \U1650/U1664/y[1] , \U1650/U1664/U30/Z , \U1650/U1664/U31/Z , 
        \U1650/U1664/U37/Z , \U1650/U1669/nr , \U1650/U1669/nd , 
        \U1650/U1669/n2 , \U1666/latch , \U1666/nlocalcd , \U1666/localcd , 
        \U1666/ncd[0] , \U1666/ncd[1] , \U1666/ncd[2] , \U1666/ncd[3] , 
        \U1666/ncd[4] , \U1666/ncd[5] , \U1666/ncd[6] , \U1666/ncd[7] , 
        \U1666/ctrlack_internal , \U1666/acb , \U1666/ba , \U1666/driveh , 
        \U1666/drivel , n6, n5, \U1666/U4/U28/U1/clr , \U1666/U4/U28/U1/set , 
        \U1666/U1/Z , \U1666/U1664/x[3] , \U1666/U1664/U28/Z , 
        \U1666/U1664/x[0] , \U1666/U1664/U32/Z , \U1666/U1664/x[2] , 
        \U1666/U1664/U29/Z , \U1666/U1664/y[0] , \U1666/U1664/x[1] , 
        \U1666/U1664/U33/Z , \U1666/U1664/y[1] , \U1666/U1664/U30/Z , 
        \U1666/U1664/U31/Z , \U1666/U1664/U37/Z , \U1666/U1669/nr , 
        \U1666/U1669/nd , \U1666/U1669/n2 , net94, \I1/latch , \I1/nlocalcd , 
        \I1/localcd , \I1/ncd[0] , \I1/ncd[1] , \I1/ncd[2] , \I1/ncd[3] , 
        \I1/ncd[4] , \I1/ncd[5] , \I1/ncd[6] , \I1/ncd[7] , 
        \I1/ctrlack_internal , \I1/acb , \I1/ba , \I1/driveh , net103, 
        \I1/drivel , n4, n3, \I1/U4/U28/U1/clr , \I1/U4/U28/U1/set , \I1/U1/Z , 
        \I1/U1664/x[3] , \I1/U1664/U28/Z , \I1/U1664/x[0] , \I1/U1664/U32/Z , 
        \I1/U1664/x[2] , \I1/U1664/U29/Z , \I1/U1664/y[0] , \I1/U1664/x[1] , 
        \I1/U1664/U33/Z , \I1/U1664/y[1] , \I1/U1664/U30/Z , \I1/U1664/U31/Z , 
        \I1/U1664/U37/Z , \I1/U1669/nr , \I1/U1669/nd , \I1/U1669/n2 , 
        \I2/latch , \I2/nlocalcd , \I2/localcd , \I2/ncd[0] , \I2/ncd[1] , 
        \I2/ncd[2] , \I2/ncd[3] , \I2/ncd[4] , \I2/ncd[5] , \I2/ncd[6] , 
        \I2/ncd[7] , \I2/ctrlack_internal , \I2/acb , \I2/ba , \I2/driveh , 
        \I2/drivel , n2, n1, \I2/U4/U28/U1/clr , \I2/U4/U28/U1/set , \I2/U1/Z , 
        \I2/U1664/x[3] , \I2/U1664/U28/Z , \I2/U1664/x[0] , \I2/U1664/U32/Z , 
        \I2/U1664/x[2] , \I2/U1664/U29/Z , \I2/U1664/y[0] , \I2/U1664/x[1] , 
        \I2/U1664/U33/Z , \I2/U1664/y[1] , \I2/U1664/U30/Z , \I2/U1664/U31/Z , 
        \I2/U1664/U37/Z , \I2/U1669/nr , \I2/U1669/nd , \I2/U1669/n2 ;
    buf_1 U262 ( .x(bpullcd), .a(pullcd) );
    or2_4 \U1674/U12  ( .x(net162), .a(nack), .b(reset) );
    and2_4 \U1785/U8  ( .x(pkt_normal), .a(\opc_l[2] ), .b(\opc_l[1] ) );
    and2_4 \U1777/U8  ( .x(net150), .a(\opc_l[2] ), .b(\opc_h[1] ) );
    or3_1 \U1813/U12  ( .x(pkt_done), .a(write), .b(reset), .c(net193) );
    nor2_1 \U1651_0_/U5  ( .x(\ncd[0] ), .a(cbh[0]), .b(cbl[0]) );
    nor2_1 \U1651_1_/U5  ( .x(\ncd[1] ), .a(cbh[1]), .b(cbl[1]) );
    nor2_1 \U1651_2_/U5  ( .x(\ncd[2] ), .a(cbh[2]), .b(cbl[2]) );
    nor2_1 \U1651_3_/U5  ( .x(\ncd[3] ), .a(cbh[3]), .b(cbl[3]) );
    nor2_1 \U1651_4_/U5  ( .x(\ncd[4] ), .a(cbh[4]), .b(cbl[4]) );
    nor2_1 \U1651_5_/U5  ( .x(\ncd[5] ), .a(cbh[5]), .b(cbl[5]) );
    nor2_1 \U1651_6_/U5  ( .x(\ncd[6] ), .a(cbh[6]), .b(cbl[6]) );
    nor2_1 \U1651_7_/U5  ( .x(\ncd[7] ), .a(cbh[7]), .b(cbl[7]) );
    nor2_1 \U1812/U5  ( .x(start_receiving), .a(notify), .b(net176) );
    nor2_1 \I7/U5  ( .x(net86), .a(net172), .b(net173) );
    nor2_1 \I4/U5  ( .x(net171), .a(net169), .b(net170) );
    nor2_1 \I3/U5  ( .x(net168), .a(net166), .b(net167) );
    inv_2 \U1675/U3  ( .x(reset), .a(nReset) );
    nand3_2 \U193/U16  ( .x(ncback), .a(net86), .b(net171), .c(net168) );
    ao222_1 \U1811/U18/U1/U1  ( .x(net176), .a(net162), .b(pkt_done), .c(
        net162), .d(net176), .e(pkt_done), .f(net176) );
    aoi222_1 \U1664/U28/U30/U1  ( .x(\U1664/x[3] ), .a(\ncd[7] ), .b(\ncd[6] ), 
        .c(\ncd[7] ), .d(\U1664/U28/Z ), .e(\ncd[6] ), .f(\U1664/U28/Z ) );
    inv_1 \U1664/U28/U30/Uinv  ( .x(\U1664/U28/Z ), .a(\U1664/x[3] ) );
    aoi222_1 \U1664/U32/U30/U1  ( .x(\U1664/x[0] ), .a(\ncd[1] ), .b(\ncd[0] ), 
        .c(\ncd[1] ), .d(\U1664/U32/Z ), .e(\ncd[0] ), .f(\U1664/U32/Z ) );
    inv_1 \U1664/U32/U30/Uinv  ( .x(\U1664/U32/Z ), .a(\U1664/x[0] ) );
    aoi222_1 \U1664/U29/U30/U1  ( .x(\U1664/x[2] ), .a(\ncd[5] ), .b(\ncd[4] ), 
        .c(\ncd[5] ), .d(\U1664/U29/Z ), .e(\ncd[4] ), .f(\U1664/U29/Z ) );
    inv_1 \U1664/U29/U30/Uinv  ( .x(\U1664/U29/Z ), .a(\U1664/x[2] ) );
    aoi222_1 \U1664/U33/U30/U1  ( .x(\U1664/y[0] ), .a(\U1664/x[1] ), .b(
        \U1664/x[0] ), .c(\U1664/x[1] ), .d(\U1664/U33/Z ), .e(\U1664/x[0] ), 
        .f(\U1664/U33/Z ) );
    inv_1 \U1664/U33/U30/Uinv  ( .x(\U1664/U33/Z ), .a(\U1664/y[0] ) );
    aoi222_1 \U1664/U30/U30/U1  ( .x(\U1664/y[1] ), .a(\U1664/x[3] ), .b(
        \U1664/x[2] ), .c(\U1664/x[3] ), .d(\U1664/U30/Z ), .e(\U1664/x[2] ), 
        .f(\U1664/U30/Z ) );
    inv_1 \U1664/U30/U30/Uinv  ( .x(\U1664/U30/Z ), .a(\U1664/y[1] ) );
    aoi222_1 \U1664/U31/U30/U1  ( .x(\U1664/x[1] ), .a(\ncd[3] ), .b(\ncd[2] ), 
        .c(\ncd[3] ), .d(\U1664/U31/Z ), .e(\ncd[2] ), .f(\U1664/U31/Z ) );
    inv_1 \U1664/U31/U30/Uinv  ( .x(\U1664/U31/Z ), .a(\U1664/x[1] ) );
    aoi222_1 \U1664/U37/U30/U1  ( .x(pullcd), .a(\U1664/y[0] ), .b(
        \U1664/y[1] ), .c(\U1664/y[0] ), .d(\U1664/U37/Z ), .e(\U1664/y[1] ), 
        .f(\U1664/U37/Z ) );
    inv_1 \U1664/U37/U30/Uinv  ( .x(\U1664/U37/Z ), .a(pullcd) );
    nor3_1 \U1697/U21/Unr  ( .x(\U1697/U21/nr ), .a(rnw[0]), .b(pkt_normal), 
        .c(net149) );
    nand3_1 \U1697/U21/Und  ( .x(\U1697/U21/nd ), .a(rnw[0]), .b(pkt_normal), 
        .c(net149) );
    oa21_1 \U1697/U21/U1  ( .x(\U1697/U21/n2 ), .a(\U1697/U21/n2 ), .b(
        \U1697/U21/nr ), .c(\U1697/U21/nd ) );
    inv_1 \U1697/U21/U3  ( .x(write), .a(\U1697/U21/n2 ) );
    nor3_1 \U307/U21/Unr  ( .x(\U307/U21/nr ), .a(net149), .b(net150), .c(
        statusack) );
    nand3_1 \U307/U21/Und  ( .x(\U307/U21/nd ), .a(net149), .b(net150), .c(
        statusack) );
    oa21_1 \U307/U21/U1  ( .x(\U307/U21/n2 ), .a(\U307/U21/n2 ), .b(
        \U307/U21/nr ), .c(\U307/U21/nd ) );
    inv_1 \U307/U21/U3  ( .x(notify), .a(\U307/U21/n2 ) );
    nor3_1 \U1698/Unr  ( .x(\U1698/nr ), .a(rnw[1]), .b(pkt_normal), .c(net149
        ) );
    nand3_1 \U1698/Und  ( .x(\U1698/nd ), .a(rnw[1]), .b(pkt_normal), .c(
        net149) );
    oa21_1 \U1698/U1  ( .x(\U1698/n2 ), .a(\U1698/n2 ), .b(\U1698/nr ), .c(
        \U1698/nd ) );
    inv_2 \U1698/U3  ( .x(read), .a(\U1698/n2 ) );
    and2_1 \U1756/U1754/U8  ( .x(n17), .a(\opc_h[0] ), .b(pkt_normal) );
    and2_1 \U1756/U1755/U8  ( .x(n18), .a(\opc_l[0] ), .b(pkt_normal) );
    and2_1 \U1800/U1754/U8  ( .x(rnw[1]), .a(net0187), .b(pkt_normal) );
    and2_1 \U1800/U1755/U8  ( .x(rnw[0]), .a(net0208), .b(pkt_normal) );
    and2_1 \U1758/U1754/U8  ( .x(status[1]), .a(\opc_h[0] ), .b(net150) );
    and2_1 \U1758/U1755/U8  ( .x(status[0]), .a(\opc_l[0] ), .b(net150) );
    buf_2 \I6/U1653  ( .x(\I6/latch ), .a(net173) );
    nor2_1 \I6/U264/U5  ( .x(\I6/nlocalcd ), .a(reset), .b(\I6/localcd ) );
    nor2_1 \I6/U1659_0_/U5  ( .x(\I6/ncd[0] ), .a(\opc_l[0] ), .b(\opc_h[0] )
         );
    nor2_1 \I6/U1659_1_/U5  ( .x(\I6/ncd[1] ), .a(\opc_l[1] ), .b(\opc_h[1] )
         );
    nor2_1 \I6/U1659_2_/U5  ( .x(\I6/ncd[2] ), .a(\opc_l[2] ), .b(\I6/oh[2] )
         );
    nor2_1 \I6/U1659_3_/U5  ( .x(\I6/ncd[3] ), .a(\I6/ol[3] ), .b(\I6/oh[3] )
         );
    nor2_1 \I6/U1659_4_/U5  ( .x(\I6/ncd[4] ), .a(\I6/ol[4] ), .b(\I6/oh[4] )
         );
    nor2_1 \I6/U1659_5_/U5  ( .x(\I6/ncd[5] ), .a(net0208), .b(net0187) );
    nor2_1 \I6/U1659_6_/U5  ( .x(\I6/ncd[6] ), .a(\I6/ol[6] ), .b(\I6/oh[6] )
         );
    nor2_1 \I6/U1659_7_/U5  ( .x(\I6/ncd[7] ), .a(\I6/ol[7] ), .b(\I6/oh[7] )
         );
    nor2_1 \I6/U3/U5  ( .x(\I6/ctrlack_internal ), .a(\I6/acb ), .b(\I6/ba )
         );
    buf_2 \I6/U1665/U7  ( .x(\I6/driveh ), .a(net139) );
    buf_2 \I6/U1666/U7  ( .x(\I6/drivel ), .a(net139) );
    ao23_1 \I6/U1658_0_/U21/U1/U1  ( .x(\opc_l[0] ), .a(\I6/driveh ), .b(
        \opc_l[0] ), .c(\I6/driveh ), .d(cbl[0]), .e(n12) );
    ao23_1 \I6/U1658_1_/U21/U1/U1  ( .x(\opc_l[1] ), .a(\I6/driveh ), .b(
        \opc_l[1] ), .c(\I6/drivel ), .d(cbl[1]), .e(n12) );
    ao23_1 \I6/U1658_2_/U21/U1/U1  ( .x(\opc_l[2] ), .a(\I6/drivel ), .b(
        \opc_l[2] ), .c(n13), .d(cbl[2]), .e(n12) );
    ao23_1 \I6/U1658_3_/U21/U1/U1  ( .x(\I6/ol[3] ), .a(\I6/drivel ), .b(
        \I6/ol[3] ), .c(\I6/drivel ), .d(cbl[3]), .e(\I6/latch ) );
    ao23_1 \I6/U1658_4_/U21/U1/U1  ( .x(\I6/ol[4] ), .a(n13), .b(\I6/ol[4] ), 
        .c(n13), .d(cbl[4]), .e(\I6/latch ) );
    ao23_1 \I6/U1658_5_/U21/U1/U1  ( .x(net0208), .a(\I6/driveh ), .b(net0208), 
        .c(\I6/driveh ), .d(cbl[5]), .e(\I6/latch ) );
    ao23_1 \I6/U1658_6_/U21/U1/U1  ( .x(\I6/ol[6] ), .a(n13), .b(\I6/ol[6] ), 
        .c(n13), .d(cbl[6]), .e(\I6/latch ) );
    ao23_1 \I6/U1658_7_/U21/U1/U1  ( .x(\I6/ol[7] ), .a(n13), .b(\I6/ol[7] ), 
        .c(\I6/driveh ), .d(cbl[7]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_0_/U21/U1/U1  ( .x(\opc_h[0] ), .a(n13), .b(\opc_h[0] ), 
        .c(\I6/drivel ), .d(cbh[0]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_1_/U21/U1/U1  ( .x(\opc_h[1] ), .a(\I6/driveh ), .b(
        \opc_h[1] ), .c(n13), .d(cbh[1]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_2_/U21/U1/U1  ( .x(\I6/oh[2] ), .a(\I6/driveh ), .b(
        \I6/oh[2] ), .c(n13), .d(cbh[2]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_3_/U21/U1/U1  ( .x(\I6/oh[3] ), .a(\I6/drivel ), .b(
        \I6/oh[3] ), .c(\I6/drivel ), .d(cbh[3]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_4_/U21/U1/U1  ( .x(\I6/oh[4] ), .a(n13), .b(\I6/oh[4] ), 
        .c(\I6/driveh ), .d(cbh[4]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_5_/U21/U1/U1  ( .x(net0187), .a(\I6/driveh ), .b(net0187), 
        .c(\I6/driveh ), .d(cbh[5]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_6_/U21/U1/U1  ( .x(\I6/oh[6] ), .a(\I6/drivel ), .b(
        \I6/oh[6] ), .c(\I6/drivel ), .d(cbh[6]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_7_/U21/U1/U1  ( .x(\I6/oh[7] ), .a(\I6/drivel ), .b(
        \I6/oh[7] ), .c(n13), .d(cbh[7]), .e(\I6/latch ) );
    aoai211_1 \I6/U4/U28/U1/U1  ( .x(\I6/U4/U28/U1/clr ), .a(net139), .b(
        \I6/acb ), .c(\I6/nlocalcd ), .d(net173) );
    nand3_1 \I6/U4/U28/U1/U2  ( .x(\I6/U4/U28/U1/set ), .a(\I6/nlocalcd ), .b(
        net139), .c(\I6/acb ) );
    nand2_2 \I6/U4/U28/U1/U3  ( .x(net173), .a(\I6/U4/U28/U1/clr ), .b(
        \I6/U4/U28/U1/set ) );
    oai21_1 \I6/U1/U30/U1/U1  ( .x(\I6/acb ), .a(\I6/U1/Z ), .b(\I6/ba ), .c(
        net139) );
    inv_1 \I6/U1/U30/U1/U2  ( .x(\I6/U1/Z ), .a(\I6/acb ) );
    ao222_1 \I6/U5/U18/U1/U1  ( .x(\I6/ba ), .a(\I6/latch ), .b(n14), .c(
        \I6/latch ), .d(\I6/ba ), .e(n14), .f(\I6/ba ) );
    aoi222_1 \I6/U1664/U28/U30/U1  ( .x(\I6/U1664/x[3] ), .a(\I6/ncd[7] ), .b(
        \I6/ncd[6] ), .c(\I6/ncd[7] ), .d(\I6/U1664/U28/Z ), .e(\I6/ncd[6] ), 
        .f(\I6/U1664/U28/Z ) );
    inv_1 \I6/U1664/U28/U30/Uinv  ( .x(\I6/U1664/U28/Z ), .a(\I6/U1664/x[3] )
         );
    aoi222_1 \I6/U1664/U32/U30/U1  ( .x(\I6/U1664/x[0] ), .a(\I6/ncd[1] ), .b(
        \I6/ncd[0] ), .c(\I6/ncd[1] ), .d(\I6/U1664/U32/Z ), .e(\I6/ncd[0] ), 
        .f(\I6/U1664/U32/Z ) );
    inv_1 \I6/U1664/U32/U30/Uinv  ( .x(\I6/U1664/U32/Z ), .a(\I6/U1664/x[0] )
         );
    aoi222_1 \I6/U1664/U29/U30/U1  ( .x(\I6/U1664/x[2] ), .a(\I6/ncd[5] ), .b(
        \I6/ncd[4] ), .c(\I6/ncd[5] ), .d(\I6/U1664/U29/Z ), .e(\I6/ncd[4] ), 
        .f(\I6/U1664/U29/Z ) );
    inv_1 \I6/U1664/U29/U30/Uinv  ( .x(\I6/U1664/U29/Z ), .a(\I6/U1664/x[2] )
         );
    aoi222_1 \I6/U1664/U33/U30/U1  ( .x(\I6/U1664/y[0] ), .a(\I6/U1664/x[1] ), 
        .b(\I6/U1664/x[0] ), .c(\I6/U1664/x[1] ), .d(\I6/U1664/U33/Z ), .e(
        \I6/U1664/x[0] ), .f(\I6/U1664/U33/Z ) );
    inv_1 \I6/U1664/U33/U30/Uinv  ( .x(\I6/U1664/U33/Z ), .a(\I6/U1664/y[0] )
         );
    aoi222_1 \I6/U1664/U30/U30/U1  ( .x(\I6/U1664/y[1] ), .a(\I6/U1664/x[3] ), 
        .b(\I6/U1664/x[2] ), .c(\I6/U1664/x[3] ), .d(\I6/U1664/U30/Z ), .e(
        \I6/U1664/x[2] ), .f(\I6/U1664/U30/Z ) );
    inv_1 \I6/U1664/U30/U30/Uinv  ( .x(\I6/U1664/U30/Z ), .a(\I6/U1664/y[1] )
         );
    aoi222_1 \I6/U1664/U31/U30/U1  ( .x(\I6/U1664/x[1] ), .a(\I6/ncd[3] ), .b(
        \I6/ncd[2] ), .c(\I6/ncd[3] ), .d(\I6/U1664/U31/Z ), .e(\I6/ncd[2] ), 
        .f(\I6/U1664/U31/Z ) );
    inv_1 \I6/U1664/U31/U30/Uinv  ( .x(\I6/U1664/U31/Z ), .a(\I6/U1664/x[1] )
         );
    aoi222_1 \I6/U1664/U37/U30/U1  ( .x(\I6/localcd ), .a(\I6/U1664/y[0] ), 
        .b(\I6/U1664/y[1] ), .c(\I6/U1664/y[0] ), .d(\I6/U1664/U37/Z ), .e(
        \I6/U1664/y[1] ), .f(\I6/U1664/U37/Z ) );
    inv_1 \I6/U1664/U37/U30/Uinv  ( .x(\I6/U1664/U37/Z ), .a(\I6/localcd ) );
    nor3_1 \I6/U1669/Unr  ( .x(\I6/U1669/nr ), .a(\I6/ctrlack_internal ), .b(
        n13), .c(\I6/drivel ) );
    nand3_1 \I6/U1669/Und  ( .x(\I6/U1669/nd ), .a(\I6/ctrlack_internal ), .b(
        \I6/driveh ), .c(\I6/drivel ) );
    oa21_1 \I6/U1669/U1  ( .x(\I6/U1669/n2 ), .a(\I6/U1669/n2 ), .b(
        \I6/U1669/nr ), .c(\I6/U1669/nd ) );
    inv_2 \I6/U1669/U3  ( .x(net149), .a(\I6/U1669/n2 ) );
    buf_2 \U1667/U1653  ( .x(\U1667/latch ), .a(net167) );
    nor2_1 \U1667/U264/U5  ( .x(\U1667/nlocalcd ), .a(reset), .b(
        \U1667/localcd ) );
    nor2_1 \U1667/U1659_0_/U5  ( .x(\U1667/ncd[0] ), .a(rd[0]), .b(rd[32]) );
    nor2_1 \U1667/U1659_1_/U5  ( .x(\U1667/ncd[1] ), .a(rd[1]), .b(rd[33]) );
    nor2_1 \U1667/U1659_2_/U5  ( .x(\U1667/ncd[2] ), .a(rd[2]), .b(rd[34]) );
    nor2_1 \U1667/U1659_3_/U5  ( .x(\U1667/ncd[3] ), .a(rd[3]), .b(rd[35]) );
    nor2_1 \U1667/U1659_4_/U5  ( .x(\U1667/ncd[4] ), .a(rd[4]), .b(rd[36]) );
    nor2_1 \U1667/U1659_5_/U5  ( .x(\U1667/ncd[5] ), .a(rd[5]), .b(rd[37]) );
    nor2_1 \U1667/U1659_6_/U5  ( .x(\U1667/ncd[6] ), .a(rd[6]), .b(rd[38]) );
    nor2_1 \U1667/U1659_7_/U5  ( .x(\U1667/ncd[7] ), .a(rd[7]), .b(rd[39]) );
    nor2_1 \U1667/U3/U5  ( .x(\U1667/ctrlack_internal ), .a(\U1667/acb ), .b(
        \U1667/ba ) );
    buf_2 \U1667/U1665/U7  ( .x(\U1667/driveh ), .a(read_lhw) );
    buf_2 \U1667/U1666/U7  ( .x(\U1667/drivel ), .a(read_lhw) );
    ao23_1 \U1667/U1658_0_/U21/U1/U1  ( .x(rd[0]), .a(n11), .b(rd[0]), .c(
        \U1667/drivel ), .d(cbl[0]), .e(n10) );
    ao23_1 \U1667/U1658_1_/U21/U1/U1  ( .x(rd[1]), .a(n11), .b(rd[1]), .c(
        \U1667/driveh ), .d(cbl[1]), .e(n10) );
    ao23_1 \U1667/U1658_2_/U21/U1/U1  ( .x(rd[2]), .a(\U1667/driveh ), .b(rd
        [2]), .c(n11), .d(cbl[2]), .e(n10) );
    ao23_1 \U1667/U1658_3_/U21/U1/U1  ( .x(rd[3]), .a(n11), .b(rd[3]), .c(
        \U1667/driveh ), .d(cbl[3]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1658_4_/U21/U1/U1  ( .x(rd[4]), .a(\U1667/drivel ), .b(rd
        [4]), .c(n11), .d(cbl[4]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1658_5_/U21/U1/U1  ( .x(rd[5]), .a(\U1667/drivel ), .b(rd
        [5]), .c(n11), .d(cbl[5]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1658_6_/U21/U1/U1  ( .x(rd[6]), .a(\U1667/driveh ), .b(rd
        [6]), .c(\U1667/drivel ), .d(cbl[6]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1658_7_/U21/U1/U1  ( .x(rd[7]), .a(\U1667/driveh ), .b(rd
        [7]), .c(\U1667/driveh ), .d(cbl[7]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_0_/U21/U1/U1  ( .x(rd[32]), .a(\U1667/drivel ), .b(rd
        [32]), .c(n11), .d(cbh[0]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_1_/U21/U1/U1  ( .x(rd[33]), .a(\U1667/driveh ), .b(rd
        [33]), .c(\U1667/drivel ), .d(cbh[1]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_2_/U21/U1/U1  ( .x(rd[34]), .a(\U1667/drivel ), .b(rd
        [34]), .c(\U1667/drivel ), .d(cbh[2]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_3_/U21/U1/U1  ( .x(rd[35]), .a(\U1667/driveh ), .b(rd
        [35]), .c(\U1667/driveh ), .d(cbh[3]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_4_/U21/U1/U1  ( .x(rd[36]), .a(\U1667/drivel ), .b(rd
        [36]), .c(\U1667/driveh ), .d(cbh[4]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_5_/U21/U1/U1  ( .x(rd[37]), .a(\U1667/driveh ), .b(rd
        [37]), .c(n11), .d(cbh[5]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_6_/U21/U1/U1  ( .x(rd[38]), .a(n11), .b(rd[38]), .c(
        \U1667/drivel ), .d(cbh[6]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_7_/U21/U1/U1  ( .x(rd[39]), .a(n11), .b(rd[39]), .c(
        n11), .d(cbh[7]), .e(\U1667/latch ) );
    aoai211_1 \U1667/U4/U28/U1/U1  ( .x(\U1667/U4/U28/U1/clr ), .a(read_lhw), 
        .b(\U1667/acb ), .c(\U1667/nlocalcd ), .d(net167) );
    nand3_1 \U1667/U4/U28/U1/U2  ( .x(\U1667/U4/U28/U1/set ), .a(
        \U1667/nlocalcd ), .b(read_lhw), .c(\U1667/acb ) );
    nand2_2 \U1667/U4/U28/U1/U3  ( .x(net167), .a(\U1667/U4/U28/U1/clr ), .b(
        \U1667/U4/U28/U1/set ) );
    oai21_1 \U1667/U1/U30/U1/U1  ( .x(\U1667/acb ), .a(\U1667/U1/Z ), .b(
        \U1667/ba ), .c(read_lhw) );
    inv_1 \U1667/U1/U30/U1/U2  ( .x(\U1667/U1/Z ), .a(\U1667/acb ) );
    ao222_1 \U1667/U5/U18/U1/U1  ( .x(\U1667/ba ), .a(\U1667/latch ), .b(n14), 
        .c(\U1667/latch ), .d(\U1667/ba ), .e(n14), .f(\U1667/ba ) );
    aoi222_1 \U1667/U1664/U28/U30/U1  ( .x(\U1667/U1664/x[3] ), .a(
        \U1667/ncd[7] ), .b(\U1667/ncd[6] ), .c(\U1667/ncd[7] ), .d(
        \U1667/U1664/U28/Z ), .e(\U1667/ncd[6] ), .f(\U1667/U1664/U28/Z ) );
    inv_1 \U1667/U1664/U28/U30/Uinv  ( .x(\U1667/U1664/U28/Z ), .a(
        \U1667/U1664/x[3] ) );
    aoi222_1 \U1667/U1664/U32/U30/U1  ( .x(\U1667/U1664/x[0] ), .a(
        \U1667/ncd[1] ), .b(\U1667/ncd[0] ), .c(\U1667/ncd[1] ), .d(
        \U1667/U1664/U32/Z ), .e(\U1667/ncd[0] ), .f(\U1667/U1664/U32/Z ) );
    inv_1 \U1667/U1664/U32/U30/Uinv  ( .x(\U1667/U1664/U32/Z ), .a(
        \U1667/U1664/x[0] ) );
    aoi222_1 \U1667/U1664/U29/U30/U1  ( .x(\U1667/U1664/x[2] ), .a(
        \U1667/ncd[5] ), .b(\U1667/ncd[4] ), .c(\U1667/ncd[5] ), .d(
        \U1667/U1664/U29/Z ), .e(\U1667/ncd[4] ), .f(\U1667/U1664/U29/Z ) );
    inv_1 \U1667/U1664/U29/U30/Uinv  ( .x(\U1667/U1664/U29/Z ), .a(
        \U1667/U1664/x[2] ) );
    aoi222_1 \U1667/U1664/U33/U30/U1  ( .x(\U1667/U1664/y[0] ), .a(
        \U1667/U1664/x[1] ), .b(\U1667/U1664/x[0] ), .c(\U1667/U1664/x[1] ), 
        .d(\U1667/U1664/U33/Z ), .e(\U1667/U1664/x[0] ), .f(
        \U1667/U1664/U33/Z ) );
    inv_1 \U1667/U1664/U33/U30/Uinv  ( .x(\U1667/U1664/U33/Z ), .a(
        \U1667/U1664/y[0] ) );
    aoi222_1 \U1667/U1664/U30/U30/U1  ( .x(\U1667/U1664/y[1] ), .a(
        \U1667/U1664/x[3] ), .b(\U1667/U1664/x[2] ), .c(\U1667/U1664/x[3] ), 
        .d(\U1667/U1664/U30/Z ), .e(\U1667/U1664/x[2] ), .f(
        \U1667/U1664/U30/Z ) );
    inv_1 \U1667/U1664/U30/U30/Uinv  ( .x(\U1667/U1664/U30/Z ), .a(
        \U1667/U1664/y[1] ) );
    aoi222_1 \U1667/U1664/U31/U30/U1  ( .x(\U1667/U1664/x[1] ), .a(
        \U1667/ncd[3] ), .b(\U1667/ncd[2] ), .c(\U1667/ncd[3] ), .d(
        \U1667/U1664/U31/Z ), .e(\U1667/ncd[2] ), .f(\U1667/U1664/U31/Z ) );
    inv_1 \U1667/U1664/U31/U30/Uinv  ( .x(\U1667/U1664/U31/Z ), .a(
        \U1667/U1664/x[1] ) );
    aoi222_1 \U1667/U1664/U37/U30/U1  ( .x(\U1667/localcd ), .a(
        \U1667/U1664/y[0] ), .b(\U1667/U1664/y[1] ), .c(\U1667/U1664/y[0] ), 
        .d(\U1667/U1664/U37/Z ), .e(\U1667/U1664/y[1] ), .f(
        \U1667/U1664/U37/Z ) );
    inv_1 \U1667/U1664/U37/U30/Uinv  ( .x(\U1667/U1664/U37/Z ), .a(
        \U1667/localcd ) );
    nor3_1 \U1667/U1669/Unr  ( .x(\U1667/U1669/nr ), .a(
        \U1667/ctrlack_internal ), .b(n11), .c(\U1667/drivel ) );
    nand3_1 \U1667/U1669/Und  ( .x(\U1667/U1669/nd ), .a(
        \U1667/ctrlack_internal ), .b(\U1667/driveh ), .c(\U1667/drivel ) );
    oa21_1 \U1667/U1669/U1  ( .x(\U1667/U1669/n2 ), .a(\U1667/U1669/n2 ), .b(
        \U1667/U1669/nr ), .c(\U1667/U1669/nd ) );
    inv_2 \U1667/U1669/U3  ( .x(net193), .a(\U1667/U1669/n2 ) );
    buf_2 \U1650/U1653  ( .x(\U1650/latch ), .a(net172) );
    nor2_1 \U1650/U264/U5  ( .x(\U1650/nlocalcd ), .a(reset), .b(
        \U1650/localcd ) );
    nor2_1 \U1650/U1659_0_/U5  ( .x(\U1650/ncd[0] ), .a(\U1650/ol[0] ), .b(
        \U1650/oh[0] ) );
    nor2_1 \U1650/U1659_1_/U5  ( .x(\U1650/ncd[1] ), .a(\U1650/ol[1] ), .b(
        \U1650/oh[1] ) );
    nor2_1 \U1650/U1659_2_/U5  ( .x(\U1650/ncd[2] ), .a(\U1650/ol[2] ), .b(
        \U1650/oh[2] ) );
    nor2_1 \U1650/U1659_3_/U5  ( .x(\U1650/ncd[3] ), .a(\U1650/ol[3] ), .b(
        \U1650/oh[3] ) );
    nor2_1 \U1650/U1659_4_/U5  ( .x(\U1650/ncd[4] ), .a(\U1650/ol[4] ), .b(
        \U1650/oh[4] ) );
    nor2_1 \U1650/U1659_5_/U5  ( .x(\U1650/ncd[5] ), .a(\col_l[0] ), .b(
        \col_h[0] ) );
    nor2_1 \U1650/U1659_6_/U5  ( .x(\U1650/ncd[6] ), .a(\col_l[1] ), .b(
        \col_h[1] ) );
    nor2_1 \U1650/U1659_7_/U5  ( .x(\U1650/ncd[7] ), .a(\col_l[2] ), .b(
        \col_h[2] ) );
    nor2_1 \U1650/U3/U5  ( .x(\U1650/ctrlack_internal ), .a(\U1650/acb ), .b(
        \U1650/ba ) );
    buf_2 \U1650/U1665/U7  ( .x(\U1650/driveh ), .a(start_receiving) );
    buf_2 \U1650/U1666/U7  ( .x(\U1650/drivel ), .a(start_receiving) );
    ao23_1 \U1650/U1658_0_/U21/U1/U1  ( .x(\U1650/ol[0] ), .a(\U1650/drivel ), 
        .b(\U1650/ol[0] ), .c(\U1650/drivel ), .d(cbl[0]), .e(n7) );
    ao23_1 \U1650/U1658_1_/U21/U1/U1  ( .x(\U1650/ol[1] ), .a(\U1650/drivel ), 
        .b(\U1650/ol[1] ), .c(\U1650/drivel ), .d(cbl[1]), .e(n7) );
    ao23_1 \U1650/U1658_2_/U21/U1/U1  ( .x(\U1650/ol[2] ), .a(\U1650/drivel ), 
        .b(\U1650/ol[2] ), .c(\U1650/drivel ), .d(cbl[2]), .e(n7) );
    ao23_1 \U1650/U1658_3_/U21/U1/U1  ( .x(\U1650/ol[3] ), .a(n9), .b(
        \U1650/ol[3] ), .c(\U1650/drivel ), .d(cbl[3]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1658_4_/U21/U1/U1  ( .x(\U1650/ol[4] ), .a(\U1650/drivel ), 
        .b(\U1650/ol[4] ), .c(\U1650/drivel ), .d(cbl[4]), .e(\U1650/latch )
         );
    ao23_1 \U1650/U1658_5_/U21/U1/U1  ( .x(\col_l[0] ), .a(\U1650/drivel ), 
        .b(\col_l[0] ), .c(\U1650/drivel ), .d(cbl[5]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1658_6_/U21/U1/U1  ( .x(\col_l[1] ), .a(n9), .b(\col_l[1] ), 
        .c(\U1650/drivel ), .d(cbl[6]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1658_7_/U21/U1/U1  ( .x(\col_l[2] ), .a(n9), .b(\col_l[2] ), 
        .c(\U1650/drivel ), .d(cbl[7]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1651_0_/U21/U1/U1  ( .x(\U1650/oh[0] ), .a(\U1650/driveh ), 
        .b(\U1650/oh[0] ), .c(\U1650/driveh ), .d(cbh[0]), .e(\U1650/latch )
         );
    ao23_1 \U1650/U1651_1_/U21/U1/U1  ( .x(\U1650/oh[1] ), .a(\U1650/driveh ), 
        .b(\U1650/oh[1] ), .c(\U1650/driveh ), .d(cbh[1]), .e(\U1650/latch )
         );
    ao23_1 \U1650/U1651_2_/U21/U1/U1  ( .x(\U1650/oh[2] ), .a(\U1650/driveh ), 
        .b(\U1650/oh[2] ), .c(\U1650/driveh ), .d(cbh[2]), .e(\U1650/latch )
         );
    ao23_1 \U1650/U1651_3_/U21/U1/U1  ( .x(\U1650/oh[3] ), .a(n8), .b(
        \U1650/oh[3] ), .c(\U1650/driveh ), .d(cbh[3]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1651_4_/U21/U1/U1  ( .x(\U1650/oh[4] ), .a(n8), .b(
        \U1650/oh[4] ), .c(\U1650/driveh ), .d(cbh[4]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1651_5_/U21/U1/U1  ( .x(\col_h[0] ), .a(\U1650/driveh ), 
        .b(\col_h[0] ), .c(\U1650/driveh ), .d(cbh[5]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1651_6_/U21/U1/U1  ( .x(\col_h[1] ), .a(n8), .b(\col_h[1] ), 
        .c(\U1650/driveh ), .d(cbh[6]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1651_7_/U21/U1/U1  ( .x(\col_h[2] ), .a(\U1650/driveh ), 
        .b(\col_h[2] ), .c(\U1650/driveh ), .d(cbh[7]), .e(\U1650/latch ) );
    aoai211_1 \U1650/U4/U28/U1/U1  ( .x(\U1650/U4/U28/U1/clr ), .a(
        start_receiving), .b(\U1650/acb ), .c(\U1650/nlocalcd ), .d(net172) );
    nand3_1 \U1650/U4/U28/U1/U2  ( .x(\U1650/U4/U28/U1/set ), .a(
        \U1650/nlocalcd ), .b(start_receiving), .c(\U1650/acb ) );
    nand2_2 \U1650/U4/U28/U1/U3  ( .x(net172), .a(\U1650/U4/U28/U1/clr ), .b(
        \U1650/U4/U28/U1/set ) );
    oai21_1 \U1650/U1/U30/U1/U1  ( .x(\U1650/acb ), .a(\U1650/U1/Z ), .b(
        \U1650/ba ), .c(start_receiving) );
    inv_1 \U1650/U1/U30/U1/U2  ( .x(\U1650/U1/Z ), .a(\U1650/acb ) );
    ao222_1 \U1650/U5/U18/U1/U1  ( .x(\U1650/ba ), .a(\U1650/latch ), .b(n14), 
        .c(\U1650/latch ), .d(\U1650/ba ), .e(n14), .f(\U1650/ba ) );
    aoi222_1 \U1650/U1664/U28/U30/U1  ( .x(\U1650/U1664/x[3] ), .a(
        \U1650/ncd[7] ), .b(\U1650/ncd[6] ), .c(\U1650/ncd[7] ), .d(
        \U1650/U1664/U28/Z ), .e(\U1650/ncd[6] ), .f(\U1650/U1664/U28/Z ) );
    inv_1 \U1650/U1664/U28/U30/Uinv  ( .x(\U1650/U1664/U28/Z ), .a(
        \U1650/U1664/x[3] ) );
    aoi222_1 \U1650/U1664/U32/U30/U1  ( .x(\U1650/U1664/x[0] ), .a(
        \U1650/ncd[1] ), .b(\U1650/ncd[0] ), .c(\U1650/ncd[1] ), .d(
        \U1650/U1664/U32/Z ), .e(\U1650/ncd[0] ), .f(\U1650/U1664/U32/Z ) );
    inv_1 \U1650/U1664/U32/U30/Uinv  ( .x(\U1650/U1664/U32/Z ), .a(
        \U1650/U1664/x[0] ) );
    aoi222_1 \U1650/U1664/U29/U30/U1  ( .x(\U1650/U1664/x[2] ), .a(
        \U1650/ncd[5] ), .b(\U1650/ncd[4] ), .c(\U1650/ncd[5] ), .d(
        \U1650/U1664/U29/Z ), .e(\U1650/ncd[4] ), .f(\U1650/U1664/U29/Z ) );
    inv_1 \U1650/U1664/U29/U30/Uinv  ( .x(\U1650/U1664/U29/Z ), .a(
        \U1650/U1664/x[2] ) );
    aoi222_1 \U1650/U1664/U33/U30/U1  ( .x(\U1650/U1664/y[0] ), .a(
        \U1650/U1664/x[1] ), .b(\U1650/U1664/x[0] ), .c(\U1650/U1664/x[1] ), 
        .d(\U1650/U1664/U33/Z ), .e(\U1650/U1664/x[0] ), .f(
        \U1650/U1664/U33/Z ) );
    inv_1 \U1650/U1664/U33/U30/Uinv  ( .x(\U1650/U1664/U33/Z ), .a(
        \U1650/U1664/y[0] ) );
    aoi222_1 \U1650/U1664/U30/U30/U1  ( .x(\U1650/U1664/y[1] ), .a(
        \U1650/U1664/x[3] ), .b(\U1650/U1664/x[2] ), .c(\U1650/U1664/x[3] ), 
        .d(\U1650/U1664/U30/Z ), .e(\U1650/U1664/x[2] ), .f(
        \U1650/U1664/U30/Z ) );
    inv_1 \U1650/U1664/U30/U30/Uinv  ( .x(\U1650/U1664/U30/Z ), .a(
        \U1650/U1664/y[1] ) );
    aoi222_1 \U1650/U1664/U31/U30/U1  ( .x(\U1650/U1664/x[1] ), .a(
        \U1650/ncd[3] ), .b(\U1650/ncd[2] ), .c(\U1650/ncd[3] ), .d(
        \U1650/U1664/U31/Z ), .e(\U1650/ncd[2] ), .f(\U1650/U1664/U31/Z ) );
    inv_1 \U1650/U1664/U31/U30/Uinv  ( .x(\U1650/U1664/U31/Z ), .a(
        \U1650/U1664/x[1] ) );
    aoi222_1 \U1650/U1664/U37/U30/U1  ( .x(\U1650/localcd ), .a(
        \U1650/U1664/y[0] ), .b(\U1650/U1664/y[1] ), .c(\U1650/U1664/y[0] ), 
        .d(\U1650/U1664/U37/Z ), .e(\U1650/U1664/y[1] ), .f(
        \U1650/U1664/U37/Z ) );
    inv_1 \U1650/U1664/U37/U30/Uinv  ( .x(\U1650/U1664/U37/Z ), .a(
        \U1650/localcd ) );
    nor3_1 \U1650/U1669/Unr  ( .x(\U1650/U1669/nr ), .a(
        \U1650/ctrlack_internal ), .b(\U1650/drivel ), .c(\U1650/driveh ) );
    nand3_1 \U1650/U1669/Und  ( .x(\U1650/U1669/nd ), .a(
        \U1650/ctrlack_internal ), .b(\U1650/drivel ), .c(\U1650/driveh ) );
    oa21_1 \U1650/U1669/U1  ( .x(\U1650/U1669/n2 ), .a(\U1650/U1669/n2 ), .b(
        \U1650/U1669/nr ), .c(\U1650/U1669/nd ) );
    inv_2 \U1650/U1669/U3  ( .x(net139), .a(\U1650/U1669/n2 ) );
    buf_2 \U1666/U1653  ( .x(\U1666/latch ), .a(net169) );
    nor2_1 \U1666/U264/U5  ( .x(\U1666/nlocalcd ), .a(reset), .b(
        \U1666/localcd ) );
    nor2_1 \U1666/U1659_0_/U5  ( .x(\U1666/ncd[0] ), .a(rd[24]), .b(rd[56]) );
    nor2_1 \U1666/U1659_1_/U5  ( .x(\U1666/ncd[1] ), .a(rd[25]), .b(rd[57]) );
    nor2_1 \U1666/U1659_2_/U5  ( .x(\U1666/ncd[2] ), .a(rd[26]), .b(rd[58]) );
    nor2_1 \U1666/U1659_3_/U5  ( .x(\U1666/ncd[3] ), .a(rd[27]), .b(rd[59]) );
    nor2_1 \U1666/U1659_4_/U5  ( .x(\U1666/ncd[4] ), .a(rd[28]), .b(rd[60]) );
    nor2_1 \U1666/U1659_5_/U5  ( .x(\U1666/ncd[5] ), .a(rd[29]), .b(rd[61]) );
    nor2_1 \U1666/U1659_6_/U5  ( .x(\U1666/ncd[6] ), .a(rd[30]), .b(rd[62]) );
    nor2_1 \U1666/U1659_7_/U5  ( .x(\U1666/ncd[7] ), .a(rd[31]), .b(rd[63]) );
    nor2_1 \U1666/U3/U5  ( .x(\U1666/ctrlack_internal ), .a(\U1666/acb ), .b(
        \U1666/ba ) );
    buf_2 \U1666/U1665/U7  ( .x(\U1666/driveh ), .a(read) );
    buf_2 \U1666/U1666/U7  ( .x(\U1666/drivel ), .a(read) );
    ao23_1 \U1666/U1658_0_/U21/U1/U1  ( .x(rd[24]), .a(n6), .b(rd[24]), .c(
        \U1666/drivel ), .d(cbl[0]), .e(n5) );
    ao23_1 \U1666/U1658_1_/U21/U1/U1  ( .x(rd[25]), .a(n6), .b(rd[25]), .c(
        \U1666/driveh ), .d(cbl[1]), .e(n5) );
    ao23_1 \U1666/U1658_2_/U21/U1/U1  ( .x(rd[26]), .a(\U1666/driveh ), .b(rd
        [26]), .c(n6), .d(cbl[2]), .e(n5) );
    ao23_1 \U1666/U1658_3_/U21/U1/U1  ( .x(rd[27]), .a(n6), .b(rd[27]), .c(
        \U1666/driveh ), .d(cbl[3]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1658_4_/U21/U1/U1  ( .x(rd[28]), .a(\U1666/drivel ), .b(rd
        [28]), .c(n6), .d(cbl[4]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1658_5_/U21/U1/U1  ( .x(rd[29]), .a(\U1666/drivel ), .b(rd
        [29]), .c(n6), .d(cbl[5]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1658_6_/U21/U1/U1  ( .x(rd[30]), .a(\U1666/driveh ), .b(rd
        [30]), .c(\U1666/drivel ), .d(cbl[6]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1658_7_/U21/U1/U1  ( .x(rd[31]), .a(\U1666/driveh ), .b(rd
        [31]), .c(\U1666/driveh ), .d(cbl[7]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_0_/U21/U1/U1  ( .x(rd[56]), .a(\U1666/drivel ), .b(rd
        [56]), .c(n6), .d(cbh[0]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_1_/U21/U1/U1  ( .x(rd[57]), .a(\U1666/driveh ), .b(rd
        [57]), .c(\U1666/drivel ), .d(cbh[1]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_2_/U21/U1/U1  ( .x(rd[58]), .a(\U1666/drivel ), .b(rd
        [58]), .c(\U1666/drivel ), .d(cbh[2]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_3_/U21/U1/U1  ( .x(rd[59]), .a(\U1666/driveh ), .b(rd
        [59]), .c(\U1666/driveh ), .d(cbh[3]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_4_/U21/U1/U1  ( .x(rd[60]), .a(\U1666/drivel ), .b(rd
        [60]), .c(\U1666/driveh ), .d(cbh[4]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_5_/U21/U1/U1  ( .x(rd[61]), .a(\U1666/driveh ), .b(rd
        [61]), .c(n6), .d(cbh[5]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_6_/U21/U1/U1  ( .x(rd[62]), .a(n6), .b(rd[62]), .c(
        \U1666/drivel ), .d(cbh[6]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_7_/U21/U1/U1  ( .x(rd[63]), .a(n6), .b(rd[63]), .c(n6), 
        .d(cbh[7]), .e(\U1666/latch ) );
    aoai211_1 \U1666/U4/U28/U1/U1  ( .x(\U1666/U4/U28/U1/clr ), .a(read), .b(
        \U1666/acb ), .c(\U1666/nlocalcd ), .d(net169) );
    nand3_1 \U1666/U4/U28/U1/U2  ( .x(\U1666/U4/U28/U1/set ), .a(
        \U1666/nlocalcd ), .b(read), .c(\U1666/acb ) );
    nand2_2 \U1666/U4/U28/U1/U3  ( .x(net169), .a(\U1666/U4/U28/U1/clr ), .b(
        \U1666/U4/U28/U1/set ) );
    oai21_1 \U1666/U1/U30/U1/U1  ( .x(\U1666/acb ), .a(\U1666/U1/Z ), .b(
        \U1666/ba ), .c(read) );
    inv_1 \U1666/U1/U30/U1/U2  ( .x(\U1666/U1/Z ), .a(\U1666/acb ) );
    ao222_1 \U1666/U5/U18/U1/U1  ( .x(\U1666/ba ), .a(\U1666/latch ), .b(n14), 
        .c(\U1666/latch ), .d(\U1666/ba ), .e(n14), .f(\U1666/ba ) );
    aoi222_1 \U1666/U1664/U28/U30/U1  ( .x(\U1666/U1664/x[3] ), .a(
        \U1666/ncd[7] ), .b(\U1666/ncd[6] ), .c(\U1666/ncd[7] ), .d(
        \U1666/U1664/U28/Z ), .e(\U1666/ncd[6] ), .f(\U1666/U1664/U28/Z ) );
    inv_1 \U1666/U1664/U28/U30/Uinv  ( .x(\U1666/U1664/U28/Z ), .a(
        \U1666/U1664/x[3] ) );
    aoi222_1 \U1666/U1664/U32/U30/U1  ( .x(\U1666/U1664/x[0] ), .a(
        \U1666/ncd[1] ), .b(\U1666/ncd[0] ), .c(\U1666/ncd[1] ), .d(
        \U1666/U1664/U32/Z ), .e(\U1666/ncd[0] ), .f(\U1666/U1664/U32/Z ) );
    inv_1 \U1666/U1664/U32/U30/Uinv  ( .x(\U1666/U1664/U32/Z ), .a(
        \U1666/U1664/x[0] ) );
    aoi222_1 \U1666/U1664/U29/U30/U1  ( .x(\U1666/U1664/x[2] ), .a(
        \U1666/ncd[5] ), .b(\U1666/ncd[4] ), .c(\U1666/ncd[5] ), .d(
        \U1666/U1664/U29/Z ), .e(\U1666/ncd[4] ), .f(\U1666/U1664/U29/Z ) );
    inv_1 \U1666/U1664/U29/U30/Uinv  ( .x(\U1666/U1664/U29/Z ), .a(
        \U1666/U1664/x[2] ) );
    aoi222_1 \U1666/U1664/U33/U30/U1  ( .x(\U1666/U1664/y[0] ), .a(
        \U1666/U1664/x[1] ), .b(\U1666/U1664/x[0] ), .c(\U1666/U1664/x[1] ), 
        .d(\U1666/U1664/U33/Z ), .e(\U1666/U1664/x[0] ), .f(
        \U1666/U1664/U33/Z ) );
    inv_1 \U1666/U1664/U33/U30/Uinv  ( .x(\U1666/U1664/U33/Z ), .a(
        \U1666/U1664/y[0] ) );
    aoi222_1 \U1666/U1664/U30/U30/U1  ( .x(\U1666/U1664/y[1] ), .a(
        \U1666/U1664/x[3] ), .b(\U1666/U1664/x[2] ), .c(\U1666/U1664/x[3] ), 
        .d(\U1666/U1664/U30/Z ), .e(\U1666/U1664/x[2] ), .f(
        \U1666/U1664/U30/Z ) );
    inv_1 \U1666/U1664/U30/U30/Uinv  ( .x(\U1666/U1664/U30/Z ), .a(
        \U1666/U1664/y[1] ) );
    aoi222_1 \U1666/U1664/U31/U30/U1  ( .x(\U1666/U1664/x[1] ), .a(
        \U1666/ncd[3] ), .b(\U1666/ncd[2] ), .c(\U1666/ncd[3] ), .d(
        \U1666/U1664/U31/Z ), .e(\U1666/ncd[2] ), .f(\U1666/U1664/U31/Z ) );
    inv_1 \U1666/U1664/U31/U30/Uinv  ( .x(\U1666/U1664/U31/Z ), .a(
        \U1666/U1664/x[1] ) );
    aoi222_1 \U1666/U1664/U37/U30/U1  ( .x(\U1666/localcd ), .a(
        \U1666/U1664/y[0] ), .b(\U1666/U1664/y[1] ), .c(\U1666/U1664/y[0] ), 
        .d(\U1666/U1664/U37/Z ), .e(\U1666/U1664/y[1] ), .f(
        \U1666/U1664/U37/Z ) );
    inv_1 \U1666/U1664/U37/U30/Uinv  ( .x(\U1666/U1664/U37/Z ), .a(
        \U1666/localcd ) );
    nor3_1 \U1666/U1669/Unr  ( .x(\U1666/U1669/nr ), .a(
        \U1666/ctrlack_internal ), .b(n6), .c(\U1666/drivel ) );
    nand3_1 \U1666/U1669/Und  ( .x(\U1666/U1669/nd ), .a(
        \U1666/ctrlack_internal ), .b(\U1666/driveh ), .c(\U1666/drivel ) );
    oa21_1 \U1666/U1669/U1  ( .x(\U1666/U1669/n2 ), .a(\U1666/U1669/n2 ), .b(
        \U1666/U1669/nr ), .c(\U1666/U1669/nd ) );
    inv_2 \U1666/U1669/U3  ( .x(net94), .a(\U1666/U1669/n2 ) );
    buf_2 \I1/U1653  ( .x(\I1/latch ), .a(net166) );
    nor2_1 \I1/U264/U5  ( .x(\I1/nlocalcd ), .a(reset), .b(\I1/localcd ) );
    nor2_1 \I1/U1659_0_/U5  ( .x(\I1/ncd[0] ), .a(rd[8]), .b(rd[40]) );
    nor2_1 \I1/U1659_1_/U5  ( .x(\I1/ncd[1] ), .a(rd[9]), .b(rd[41]) );
    nor2_1 \I1/U1659_2_/U5  ( .x(\I1/ncd[2] ), .a(rd[10]), .b(rd[42]) );
    nor2_1 \I1/U1659_3_/U5  ( .x(\I1/ncd[3] ), .a(rd[11]), .b(rd[43]) );
    nor2_1 \I1/U1659_4_/U5  ( .x(\I1/ncd[4] ), .a(rd[12]), .b(rd[44]) );
    nor2_1 \I1/U1659_5_/U5  ( .x(\I1/ncd[5] ), .a(rd[13]), .b(rd[45]) );
    nor2_1 \I1/U1659_6_/U5  ( .x(\I1/ncd[6] ), .a(rd[14]), .b(rd[46]) );
    nor2_1 \I1/U1659_7_/U5  ( .x(\I1/ncd[7] ), .a(rd[15]), .b(rd[47]) );
    nor2_1 \I1/U3/U5  ( .x(\I1/ctrlack_internal ), .a(\I1/acb ), .b(\I1/ba )
         );
    buf_2 \I1/U1665/U7  ( .x(\I1/driveh ), .a(net103) );
    buf_2 \I1/U1666/U7  ( .x(\I1/drivel ), .a(net103) );
    ao23_1 \I1/U1658_0_/U21/U1/U1  ( .x(rd[8]), .a(n4), .b(rd[8]), .c(
        \I1/drivel ), .d(cbl[0]), .e(n3) );
    ao23_1 \I1/U1658_1_/U21/U1/U1  ( .x(rd[9]), .a(n4), .b(rd[9]), .c(
        \I1/driveh ), .d(cbl[1]), .e(n3) );
    ao23_1 \I1/U1658_2_/U21/U1/U1  ( .x(rd[10]), .a(\I1/driveh ), .b(rd[10]), 
        .c(n4), .d(cbl[2]), .e(n3) );
    ao23_1 \I1/U1658_3_/U21/U1/U1  ( .x(rd[11]), .a(n4), .b(rd[11]), .c(
        \I1/driveh ), .d(cbl[3]), .e(\I1/latch ) );
    ao23_1 \I1/U1658_4_/U21/U1/U1  ( .x(rd[12]), .a(\I1/drivel ), .b(rd[12]), 
        .c(n4), .d(cbl[4]), .e(\I1/latch ) );
    ao23_1 \I1/U1658_5_/U21/U1/U1  ( .x(rd[13]), .a(\I1/drivel ), .b(rd[13]), 
        .c(n4), .d(cbl[5]), .e(\I1/latch ) );
    ao23_1 \I1/U1658_6_/U21/U1/U1  ( .x(rd[14]), .a(\I1/driveh ), .b(rd[14]), 
        .c(\I1/drivel ), .d(cbl[6]), .e(\I1/latch ) );
    ao23_1 \I1/U1658_7_/U21/U1/U1  ( .x(rd[15]), .a(\I1/driveh ), .b(rd[15]), 
        .c(\I1/driveh ), .d(cbl[7]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_0_/U21/U1/U1  ( .x(rd[40]), .a(\I1/drivel ), .b(rd[40]), 
        .c(n4), .d(cbh[0]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_1_/U21/U1/U1  ( .x(rd[41]), .a(\I1/driveh ), .b(rd[41]), 
        .c(\I1/drivel ), .d(cbh[1]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_2_/U21/U1/U1  ( .x(rd[42]), .a(\I1/drivel ), .b(rd[42]), 
        .c(\I1/drivel ), .d(cbh[2]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_3_/U21/U1/U1  ( .x(rd[43]), .a(\I1/driveh ), .b(rd[43]), 
        .c(\I1/driveh ), .d(cbh[3]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_4_/U21/U1/U1  ( .x(rd[44]), .a(\I1/drivel ), .b(rd[44]), 
        .c(\I1/driveh ), .d(cbh[4]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_5_/U21/U1/U1  ( .x(rd[45]), .a(\I1/driveh ), .b(rd[45]), 
        .c(n4), .d(cbh[5]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_6_/U21/U1/U1  ( .x(rd[46]), .a(n4), .b(rd[46]), .c(
        \I1/drivel ), .d(cbh[6]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_7_/U21/U1/U1  ( .x(rd[47]), .a(n4), .b(rd[47]), .c(n4), 
        .d(cbh[7]), .e(\I1/latch ) );
    aoai211_1 \I1/U4/U28/U1/U1  ( .x(\I1/U4/U28/U1/clr ), .a(net103), .b(
        \I1/acb ), .c(\I1/nlocalcd ), .d(net166) );
    nand3_1 \I1/U4/U28/U1/U2  ( .x(\I1/U4/U28/U1/set ), .a(\I1/nlocalcd ), .b(
        net103), .c(\I1/acb ) );
    nand2_2 \I1/U4/U28/U1/U3  ( .x(net166), .a(\I1/U4/U28/U1/clr ), .b(
        \I1/U4/U28/U1/set ) );
    oai21_1 \I1/U1/U30/U1/U1  ( .x(\I1/acb ), .a(\I1/U1/Z ), .b(\I1/ba ), .c(
        net103) );
    inv_1 \I1/U1/U30/U1/U2  ( .x(\I1/U1/Z ), .a(\I1/acb ) );
    ao222_1 \I1/U5/U18/U1/U1  ( .x(\I1/ba ), .a(\I1/latch ), .b(n14), .c(
        \I1/latch ), .d(\I1/ba ), .e(n14), .f(\I1/ba ) );
    aoi222_1 \I1/U1664/U28/U30/U1  ( .x(\I1/U1664/x[3] ), .a(\I1/ncd[7] ), .b(
        \I1/ncd[6] ), .c(\I1/ncd[7] ), .d(\I1/U1664/U28/Z ), .e(\I1/ncd[6] ), 
        .f(\I1/U1664/U28/Z ) );
    inv_1 \I1/U1664/U28/U30/Uinv  ( .x(\I1/U1664/U28/Z ), .a(\I1/U1664/x[3] )
         );
    aoi222_1 \I1/U1664/U32/U30/U1  ( .x(\I1/U1664/x[0] ), .a(\I1/ncd[1] ), .b(
        \I1/ncd[0] ), .c(\I1/ncd[1] ), .d(\I1/U1664/U32/Z ), .e(\I1/ncd[0] ), 
        .f(\I1/U1664/U32/Z ) );
    inv_1 \I1/U1664/U32/U30/Uinv  ( .x(\I1/U1664/U32/Z ), .a(\I1/U1664/x[0] )
         );
    aoi222_1 \I1/U1664/U29/U30/U1  ( .x(\I1/U1664/x[2] ), .a(\I1/ncd[5] ), .b(
        \I1/ncd[4] ), .c(\I1/ncd[5] ), .d(\I1/U1664/U29/Z ), .e(\I1/ncd[4] ), 
        .f(\I1/U1664/U29/Z ) );
    inv_1 \I1/U1664/U29/U30/Uinv  ( .x(\I1/U1664/U29/Z ), .a(\I1/U1664/x[2] )
         );
    aoi222_1 \I1/U1664/U33/U30/U1  ( .x(\I1/U1664/y[0] ), .a(\I1/U1664/x[1] ), 
        .b(\I1/U1664/x[0] ), .c(\I1/U1664/x[1] ), .d(\I1/U1664/U33/Z ), .e(
        \I1/U1664/x[0] ), .f(\I1/U1664/U33/Z ) );
    inv_1 \I1/U1664/U33/U30/Uinv  ( .x(\I1/U1664/U33/Z ), .a(\I1/U1664/y[0] )
         );
    aoi222_1 \I1/U1664/U30/U30/U1  ( .x(\I1/U1664/y[1] ), .a(\I1/U1664/x[3] ), 
        .b(\I1/U1664/x[2] ), .c(\I1/U1664/x[3] ), .d(\I1/U1664/U30/Z ), .e(
        \I1/U1664/x[2] ), .f(\I1/U1664/U30/Z ) );
    inv_1 \I1/U1664/U30/U30/Uinv  ( .x(\I1/U1664/U30/Z ), .a(\I1/U1664/y[1] )
         );
    aoi222_1 \I1/U1664/U31/U30/U1  ( .x(\I1/U1664/x[1] ), .a(\I1/ncd[3] ), .b(
        \I1/ncd[2] ), .c(\I1/ncd[3] ), .d(\I1/U1664/U31/Z ), .e(\I1/ncd[2] ), 
        .f(\I1/U1664/U31/Z ) );
    inv_1 \I1/U1664/U31/U30/Uinv  ( .x(\I1/U1664/U31/Z ), .a(\I1/U1664/x[1] )
         );
    aoi222_1 \I1/U1664/U37/U30/U1  ( .x(\I1/localcd ), .a(\I1/U1664/y[0] ), 
        .b(\I1/U1664/y[1] ), .c(\I1/U1664/y[0] ), .d(\I1/U1664/U37/Z ), .e(
        \I1/U1664/y[1] ), .f(\I1/U1664/U37/Z ) );
    inv_1 \I1/U1664/U37/U30/Uinv  ( .x(\I1/U1664/U37/Z ), .a(\I1/localcd ) );
    nor3_1 \I1/U1669/Unr  ( .x(\I1/U1669/nr ), .a(\I1/ctrlack_internal ), .b(
        n4), .c(\I1/drivel ) );
    nand3_1 \I1/U1669/Und  ( .x(\I1/U1669/nd ), .a(\I1/ctrlack_internal ), .b(
        \I1/driveh ), .c(\I1/drivel ) );
    oa21_1 \I1/U1669/U1  ( .x(\I1/U1669/n2 ), .a(\I1/U1669/n2 ), .b(
        \I1/U1669/nr ), .c(\I1/U1669/nd ) );
    inv_2 \I1/U1669/U3  ( .x(read_lhw), .a(\I1/U1669/n2 ) );
    buf_2 \I2/U1653  ( .x(\I2/latch ), .a(net170) );
    nor2_1 \I2/U264/U5  ( .x(\I2/nlocalcd ), .a(reset), .b(\I2/localcd ) );
    nor2_1 \I2/U1659_0_/U5  ( .x(\I2/ncd[0] ), .a(rd[16]), .b(rd[48]) );
    nor2_1 \I2/U1659_1_/U5  ( .x(\I2/ncd[1] ), .a(rd[17]), .b(rd[49]) );
    nor2_1 \I2/U1659_2_/U5  ( .x(\I2/ncd[2] ), .a(rd[18]), .b(rd[50]) );
    nor2_1 \I2/U1659_3_/U5  ( .x(\I2/ncd[3] ), .a(rd[19]), .b(rd[51]) );
    nor2_1 \I2/U1659_4_/U5  ( .x(\I2/ncd[4] ), .a(rd[20]), .b(rd[52]) );
    nor2_1 \I2/U1659_5_/U5  ( .x(\I2/ncd[5] ), .a(rd[21]), .b(rd[53]) );
    nor2_1 \I2/U1659_6_/U5  ( .x(\I2/ncd[6] ), .a(rd[22]), .b(rd[54]) );
    nor2_1 \I2/U1659_7_/U5  ( .x(\I2/ncd[7] ), .a(rd[23]), .b(rd[55]) );
    nor2_1 \I2/U3/U5  ( .x(\I2/ctrlack_internal ), .a(\I2/acb ), .b(\I2/ba )
         );
    buf_2 \I2/U1665/U7  ( .x(\I2/driveh ), .a(net94) );
    buf_2 \I2/U1666/U7  ( .x(\I2/drivel ), .a(net94) );
    ao23_1 \I2/U1658_0_/U21/U1/U1  ( .x(rd[16]), .a(n2), .b(rd[16]), .c(
        \I2/drivel ), .d(cbl[0]), .e(n1) );
    ao23_1 \I2/U1658_1_/U21/U1/U1  ( .x(rd[17]), .a(n2), .b(rd[17]), .c(
        \I2/driveh ), .d(cbl[1]), .e(n1) );
    ao23_1 \I2/U1658_2_/U21/U1/U1  ( .x(rd[18]), .a(\I2/driveh ), .b(rd[18]), 
        .c(n2), .d(cbl[2]), .e(n1) );
    ao23_1 \I2/U1658_3_/U21/U1/U1  ( .x(rd[19]), .a(n2), .b(rd[19]), .c(
        \I2/driveh ), .d(cbl[3]), .e(\I2/latch ) );
    ao23_1 \I2/U1658_4_/U21/U1/U1  ( .x(rd[20]), .a(\I2/drivel ), .b(rd[20]), 
        .c(n2), .d(cbl[4]), .e(\I2/latch ) );
    ao23_1 \I2/U1658_5_/U21/U1/U1  ( .x(rd[21]), .a(\I2/drivel ), .b(rd[21]), 
        .c(n2), .d(cbl[5]), .e(\I2/latch ) );
    ao23_1 \I2/U1658_6_/U21/U1/U1  ( .x(rd[22]), .a(\I2/driveh ), .b(rd[22]), 
        .c(\I2/drivel ), .d(cbl[6]), .e(\I2/latch ) );
    ao23_1 \I2/U1658_7_/U21/U1/U1  ( .x(rd[23]), .a(\I2/driveh ), .b(rd[23]), 
        .c(\I2/driveh ), .d(cbl[7]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_0_/U21/U1/U1  ( .x(rd[48]), .a(\I2/drivel ), .b(rd[48]), 
        .c(n2), .d(cbh[0]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_1_/U21/U1/U1  ( .x(rd[49]), .a(\I2/driveh ), .b(rd[49]), 
        .c(\I2/drivel ), .d(cbh[1]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_2_/U21/U1/U1  ( .x(rd[50]), .a(\I2/drivel ), .b(rd[50]), 
        .c(\I2/drivel ), .d(cbh[2]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_3_/U21/U1/U1  ( .x(rd[51]), .a(\I2/driveh ), .b(rd[51]), 
        .c(\I2/driveh ), .d(cbh[3]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_4_/U21/U1/U1  ( .x(rd[52]), .a(\I2/drivel ), .b(rd[52]), 
        .c(\I2/driveh ), .d(cbh[4]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_5_/U21/U1/U1  ( .x(rd[53]), .a(\I2/driveh ), .b(rd[53]), 
        .c(n2), .d(cbh[5]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_6_/U21/U1/U1  ( .x(rd[54]), .a(n2), .b(rd[54]), .c(
        \I2/drivel ), .d(cbh[6]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_7_/U21/U1/U1  ( .x(rd[55]), .a(n2), .b(rd[55]), .c(n2), 
        .d(cbh[7]), .e(\I2/latch ) );
    aoai211_1 \I2/U4/U28/U1/U1  ( .x(\I2/U4/U28/U1/clr ), .a(net94), .b(
        \I2/acb ), .c(\I2/nlocalcd ), .d(net170) );
    nand3_1 \I2/U4/U28/U1/U2  ( .x(\I2/U4/U28/U1/set ), .a(\I2/nlocalcd ), .b(
        net94), .c(\I2/acb ) );
    nand2_2 \I2/U4/U28/U1/U3  ( .x(net170), .a(\I2/U4/U28/U1/clr ), .b(
        \I2/U4/U28/U1/set ) );
    oai21_1 \I2/U1/U30/U1/U1  ( .x(\I2/acb ), .a(\I2/U1/Z ), .b(\I2/ba ), .c(
        net94) );
    inv_1 \I2/U1/U30/U1/U2  ( .x(\I2/U1/Z ), .a(\I2/acb ) );
    ao222_1 \I2/U5/U18/U1/U1  ( .x(\I2/ba ), .a(\I2/latch ), .b(n14), .c(
        \I2/latch ), .d(\I2/ba ), .e(n14), .f(\I2/ba ) );
    aoi222_1 \I2/U1664/U28/U30/U1  ( .x(\I2/U1664/x[3] ), .a(\I2/ncd[7] ), .b(
        \I2/ncd[6] ), .c(\I2/ncd[7] ), .d(\I2/U1664/U28/Z ), .e(\I2/ncd[6] ), 
        .f(\I2/U1664/U28/Z ) );
    inv_1 \I2/U1664/U28/U30/Uinv  ( .x(\I2/U1664/U28/Z ), .a(\I2/U1664/x[3] )
         );
    aoi222_1 \I2/U1664/U32/U30/U1  ( .x(\I2/U1664/x[0] ), .a(\I2/ncd[1] ), .b(
        \I2/ncd[0] ), .c(\I2/ncd[1] ), .d(\I2/U1664/U32/Z ), .e(\I2/ncd[0] ), 
        .f(\I2/U1664/U32/Z ) );
    inv_1 \I2/U1664/U32/U30/Uinv  ( .x(\I2/U1664/U32/Z ), .a(\I2/U1664/x[0] )
         );
    aoi222_1 \I2/U1664/U29/U30/U1  ( .x(\I2/U1664/x[2] ), .a(\I2/ncd[5] ), .b(
        \I2/ncd[4] ), .c(\I2/ncd[5] ), .d(\I2/U1664/U29/Z ), .e(\I2/ncd[4] ), 
        .f(\I2/U1664/U29/Z ) );
    inv_1 \I2/U1664/U29/U30/Uinv  ( .x(\I2/U1664/U29/Z ), .a(\I2/U1664/x[2] )
         );
    aoi222_1 \I2/U1664/U33/U30/U1  ( .x(\I2/U1664/y[0] ), .a(\I2/U1664/x[1] ), 
        .b(\I2/U1664/x[0] ), .c(\I2/U1664/x[1] ), .d(\I2/U1664/U33/Z ), .e(
        \I2/U1664/x[0] ), .f(\I2/U1664/U33/Z ) );
    inv_1 \I2/U1664/U33/U30/Uinv  ( .x(\I2/U1664/U33/Z ), .a(\I2/U1664/y[0] )
         );
    aoi222_1 \I2/U1664/U30/U30/U1  ( .x(\I2/U1664/y[1] ), .a(\I2/U1664/x[3] ), 
        .b(\I2/U1664/x[2] ), .c(\I2/U1664/x[3] ), .d(\I2/U1664/U30/Z ), .e(
        \I2/U1664/x[2] ), .f(\I2/U1664/U30/Z ) );
    inv_1 \I2/U1664/U30/U30/Uinv  ( .x(\I2/U1664/U30/Z ), .a(\I2/U1664/y[1] )
         );
    aoi222_1 \I2/U1664/U31/U30/U1  ( .x(\I2/U1664/x[1] ), .a(\I2/ncd[3] ), .b(
        \I2/ncd[2] ), .c(\I2/ncd[3] ), .d(\I2/U1664/U31/Z ), .e(\I2/ncd[2] ), 
        .f(\I2/U1664/U31/Z ) );
    inv_1 \I2/U1664/U31/U30/Uinv  ( .x(\I2/U1664/U31/Z ), .a(\I2/U1664/x[1] )
         );
    aoi222_1 \I2/U1664/U37/U30/U1  ( .x(\I2/localcd ), .a(\I2/U1664/y[0] ), 
        .b(\I2/U1664/y[1] ), .c(\I2/U1664/y[0] ), .d(\I2/U1664/U37/Z ), .e(
        \I2/U1664/y[1] ), .f(\I2/U1664/U37/Z ) );
    inv_1 \I2/U1664/U37/U30/Uinv  ( .x(\I2/U1664/U37/Z ), .a(\I2/localcd ) );
    nor3_1 \I2/U1669/Unr  ( .x(\I2/U1669/nr ), .a(\I2/ctrlack_internal ), .b(
        n2), .c(\I2/drivel ) );
    nand3_1 \I2/U1669/Und  ( .x(\I2/U1669/nd ), .a(\I2/ctrlack_internal ), .b(
        \I2/driveh ), .c(\I2/drivel ) );
    oa21_1 \I2/U1669/U1  ( .x(\I2/U1669/n2 ), .a(\I2/U1669/n2 ), .b(
        \I2/U1669/nr ), .c(\I2/U1669/nd ) );
    inv_2 \I2/U1669/U3  ( .x(net103), .a(\I2/U1669/n2 ) );
    buf_1 U1 ( .x(n1), .a(\I2/latch ) );
    buf_2 U2 ( .x(n2), .a(net94) );
    buf_1 U3 ( .x(n3), .a(\I1/latch ) );
    buf_2 U4 ( .x(n4), .a(net103) );
    buf_1 U5 ( .x(n5), .a(\U1666/latch ) );
    buf_2 U6 ( .x(n6), .a(read) );
    buf_1 U7 ( .x(n7), .a(\U1650/latch ) );
    buf_1 U8 ( .x(n8), .a(\U1650/driveh ) );
    buf_1 U9 ( .x(n9), .a(\U1650/drivel ) );
    buf_1 U10 ( .x(n10), .a(\U1667/latch ) );
    buf_2 U11 ( .x(n11), .a(read_lhw) );
    buf_1 U12 ( .x(n12), .a(\I6/latch ) );
    buf_2 U13 ( .x(n13), .a(net139) );
    buf_3 U14 ( .x(n14), .a(bpullcd) );
    buf_3 U15 ( .x(err[0]), .a(n18) );
    buf_3 U16 ( .x(err[1]), .a(n17) );
endmodule


module chain_fr2dr_byte_3 ( nia, oh, ol, i, nReset, noa );
output [7:0] oh;
output [7:0] ol;
input  [4:0] i;
input  nReset, noa;
output nia;
    wire nbReset, eop, ncla, csela, asela, \U891/reset , \U891/neopack , 
        \U891/iay , \U891/naack[0] , \U891/naack[1] , \U891/U1128/nb , \b[3] , 
        \b[2] , \U891/U1128/na , \b[1] , \b[0] , \U891/ackb , \a[3] , \a[2] , 
        \U891/nack , \U891/acka , \a[1] , \a[0] , bsela, bsel, asel, 
        \U891/U1118_0_/nr , naa, \U891/U1118_0_/nd , \U891/U1118_0_/n2 , 
        \U891/U1118_1_/nr , \U891/U1118_1_/nd , \U891/U1118_1_/n2 , 
        \U891/U1118_2_/nr , \U891/U1118_2_/nd , \U891/U1118_2_/n2 , 
        \U891/U1118_3_/nr , \U891/U1118_3_/nd , \U891/U1118_3_/n2 , 
        \U891/U1117_0_/nr , nba, \U891/U1117_0_/nd , \U891/U1117_0_/n2 , 
        \U891/U1117_1_/nr , \U891/U1117_1_/nd , \U891/U1117_1_/n2 , 
        \U891/U1117_2_/nr , \U891/U1117_2_/nd , \U891/U1117_2_/n2 , 
        \U891/U1117_3_/nr , \U891/U1117_3_/nd , \U891/U1117_3_/n2 , 
        \U886/reset , \U886/U1128/nb , \f[3] , \f[2] , \U886/U1128/na , \f[1] , 
        \f[0] , \U886/ackb , \U886/nack , \U886/acka , \U886/U1127/n5 , 
        \U886/U1127/n1 , \U886/U1127/n2 , \U886/U1127/n3 , \U886/U1127/n4 , 
        \e[3] , \e[2] , \e[1] , \e[0] , fsela, fsel, esela, esel, 
        \U886/U1118_0_/nr , nea, \U886/U1118_0_/nd , \U886/U1118_0_/n2 , 
        \U886/U1118_1_/nr , \U886/U1118_1_/nd , \U886/U1118_1_/n2 , 
        \U886/U1118_2_/nr , \U886/U1118_2_/nd , \U886/U1118_2_/n2 , 
        \U886/U1118_3_/nr , \U886/U1118_3_/nd , \U886/U1118_3_/n2 , 
        \U886/U1117_0_/nr , nfa, \U886/U1117_0_/nd , \U886/U1117_0_/n2 , 
        \U886/U1117_1_/nr , \U886/U1117_1_/nd , \U886/U1117_1_/n2 , 
        \U886/U1117_2_/nr , \U886/U1117_2_/nd , \U886/U1117_2_/n2 , 
        \U886/U1117_3_/nr , \U886/U1117_3_/nd , \U886/U1117_3_/n2 , 
        \U884/reset , \U884/U1128/nb , \d[3] , \d[2] , \U884/U1128/na , \d[1] , 
        \d[0] , \U884/ackb , \U884/nack , \U884/acka , \U884/U1127/n5 , 
        \U884/U1127/n1 , \U884/U1127/n2 , \U884/U1127/n3 , \U884/U1127/n4 , 
        \c[3] , \c[2] , \c[1] , \c[0] , dsela, dsel, csel, \U884/U1118_0_/nr , 
        nca, \U884/U1118_0_/nd , \U884/U1118_0_/n2 , \U884/U1118_1_/nr , 
        \U884/U1118_1_/nd , \U884/U1118_1_/n2 , \U884/U1118_2_/nr , 
        \U884/U1118_2_/nd , \U884/U1118_2_/n2 , \U884/U1118_3_/nr , 
        \U884/U1118_3_/nd , \U884/U1118_3_/n2 , \U884/U1117_0_/nr , nda, 
        \U884/U1117_0_/nd , \U884/U1117_0_/n2 , \U884/U1117_1_/nr , 
        \U884/U1117_1_/nd , \U884/U1117_1_/n2 , \U884/U1117_2_/nr , 
        \U884/U1117_2_/nd , \U884/U1117_2_/n2 , \U884/U1117_3_/nr , 
        \U884/U1117_3_/nd , \U884/U1117_3_/n2 , \U888/s , \U888/r , 
        \U888/nback , \U888/naack , \U888/reset , \U887/s , \U887/r , 
        \U887/nback , \U887/naack , \U887/reset , \U885/s , \U885/r , 
        \U885/nback , \U885/naack , \U885/reset , \U877/x , \U877/reset , 
        \U877/y , \U877/U590/U25/U1/clr , net135, \cl[3] , \cl[1] , 
        \U877/U590/U25/U1/ob , n1, \U877/U589/U25/U1/clr , \cl[0] , 
        \U877/U589/U25/U1/ob , \U877/U588/U25/U1/clr , \cl[2] , 
        \U877/U588/U25/U1/ob , \U877/U591/U25/U1/clr , \U877/U591/U25/U1/ob , 
        \U876/x , \U876/reset , \U876/y , \U876/U590/U25/U1/clr , 
        \U876/U590/U25/U1/ob , \U876/U589/U25/U1/clr , \U876/U589/U25/U1/ob , 
        \U876/U588/U25/U1/clr , \U876/U588/U25/U1/ob , \U876/U591/U25/U1/clr , 
        \U876/U591/U25/U1/ob , \U2/x , \U2/reset , \U2/y , 
        \U2/U590/U25/U1/clr , \U2/U590/U25/U1/ob , \U2/U589/U25/U1/clr , 
        \U2/U589/U25/U1/ob , \U2/U588/U25/U1/clr , \U2/U588/U25/U1/ob , 
        \U2/U591/U25/U1/clr , \U2/U591/U25/U1/ob , \U1/x , \U1/reset , \U1/y , 
        \U1/U590/U25/U1/clr , \U1/U590/U25/U1/ob , \U1/U589/U25/U1/clr , 
        \U1/U589/U25/U1/ob , \U1/U588/U25/U1/clr , \U1/U588/U25/U1/ob , 
        \U1/U591/U25/U1/clr , \U1/U591/U25/U1/ob , \U881/nack[1] , 
        \U881/nack[0] ;
    buf_2 U897 ( .x(nbReset), .a(nReset) );
    and4_1 \U894/U12  ( .x(eop), .a(ncla), .b(csela), .c(asela), .d(i[4]) );
    inv_1 \U891/U1126/U3  ( .x(\U891/reset ), .a(nbReset) );
    inv_1 \U891/U1139/U3  ( .x(\U891/neopack ), .a(eop) );
    nand3_1 \U891/U1131/U9  ( .x(\U891/iay ), .a(\U891/neopack ), .b(
        \U891/naack[0] ), .c(\U891/naack[1] ) );
    nor3_1 \U891/U1128/U27  ( .x(\U891/U1128/nb ), .a(\U891/reset ), .b(\b[3] 
        ), .c(\b[2] ) );
    nor2_1 \U891/U1128/U26  ( .x(\U891/U1128/na ), .a(\b[1] ), .b(\b[0] ) );
    nand2_2 \U891/U1128/U29  ( .x(\U891/ackb ), .a(\U891/U1128/nb ), .b(
        \U891/U1128/na ) );
    nor2_1 \U891/U1133/U5  ( .x(\U891/naack[0] ), .a(\a[3] ), .b(\a[2] ) );
    nor2_1 \U891/U1108/U5  ( .x(\U891/nack ), .a(\U891/acka ), .b(\U891/ackb )
         );
    nor2_1 \U891/U1134/U5  ( .x(\U891/naack[1] ), .a(\a[1] ), .b(\a[0] ) );
    nor2_2 \U891/U914/U6  ( .x(nia), .a(\U891/iay ), .b(\U891/ackb ) );
    nand2_1 \U891/U1130/U5  ( .x(\U891/acka ), .a(\U891/naack[0] ), .b(
        \U891/naack[1] ) );
    ao222_4 \U891/U1121/U1/U1  ( .x(bsela), .a(\U891/nack ), .b(bsel), .c(
        \U891/nack ), .d(bsela), .e(bsel), .f(bsela) );
    ao222_4 \U891/U1120/U1/U1  ( .x(asela), .a(asel), .b(\U891/nack ), .c(asel
        ), .d(asela), .e(\U891/nack ), .f(asela) );
    nor3_1 \U891/U1118_0_/Unr  ( .x(\U891/U1118_0_/nr ), .a(i[0]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_0_/Und  ( .x(\U891/U1118_0_/nd ), .a(i[0]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_0_/U1  ( .x(\U891/U1118_0_/n2 ), .a(\U891/U1118_0_/n2 ), 
        .b(\U891/U1118_0_/nr ), .c(\U891/U1118_0_/nd ) );
    inv_2 \U891/U1118_0_/U3  ( .x(\a[0] ), .a(\U891/U1118_0_/n2 ) );
    nor3_1 \U891/U1118_1_/Unr  ( .x(\U891/U1118_1_/nr ), .a(i[1]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_1_/Und  ( .x(\U891/U1118_1_/nd ), .a(i[1]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_1_/U1  ( .x(\U891/U1118_1_/n2 ), .a(\U891/U1118_1_/n2 ), 
        .b(\U891/U1118_1_/nr ), .c(\U891/U1118_1_/nd ) );
    inv_2 \U891/U1118_1_/U3  ( .x(\a[1] ), .a(\U891/U1118_1_/n2 ) );
    nor3_1 \U891/U1118_2_/Unr  ( .x(\U891/U1118_2_/nr ), .a(i[2]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_2_/Und  ( .x(\U891/U1118_2_/nd ), .a(i[2]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_2_/U1  ( .x(\U891/U1118_2_/n2 ), .a(\U891/U1118_2_/n2 ), 
        .b(\U891/U1118_2_/nr ), .c(\U891/U1118_2_/nd ) );
    inv_2 \U891/U1118_2_/U3  ( .x(\a[2] ), .a(\U891/U1118_2_/n2 ) );
    nor3_1 \U891/U1118_3_/Unr  ( .x(\U891/U1118_3_/nr ), .a(i[3]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_3_/Und  ( .x(\U891/U1118_3_/nd ), .a(i[3]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_3_/U1  ( .x(\U891/U1118_3_/n2 ), .a(\U891/U1118_3_/n2 ), 
        .b(\U891/U1118_3_/nr ), .c(\U891/U1118_3_/nd ) );
    inv_2 \U891/U1118_3_/U3  ( .x(\a[3] ), .a(\U891/U1118_3_/n2 ) );
    nor3_1 \U891/U1117_0_/Unr  ( .x(\U891/U1117_0_/nr ), .a(i[0]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_0_/Und  ( .x(\U891/U1117_0_/nd ), .a(i[0]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_0_/U1  ( .x(\U891/U1117_0_/n2 ), .a(\U891/U1117_0_/n2 ), 
        .b(\U891/U1117_0_/nr ), .c(\U891/U1117_0_/nd ) );
    inv_2 \U891/U1117_0_/U3  ( .x(\b[0] ), .a(\U891/U1117_0_/n2 ) );
    nor3_1 \U891/U1117_1_/Unr  ( .x(\U891/U1117_1_/nr ), .a(i[1]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_1_/Und  ( .x(\U891/U1117_1_/nd ), .a(i[1]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_1_/U1  ( .x(\U891/U1117_1_/n2 ), .a(\U891/U1117_1_/n2 ), 
        .b(\U891/U1117_1_/nr ), .c(\U891/U1117_1_/nd ) );
    inv_2 \U891/U1117_1_/U3  ( .x(\b[1] ), .a(\U891/U1117_1_/n2 ) );
    nor3_1 \U891/U1117_2_/Unr  ( .x(\U891/U1117_2_/nr ), .a(i[2]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_2_/Und  ( .x(\U891/U1117_2_/nd ), .a(i[2]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_2_/U1  ( .x(\U891/U1117_2_/n2 ), .a(\U891/U1117_2_/n2 ), 
        .b(\U891/U1117_2_/nr ), .c(\U891/U1117_2_/nd ) );
    inv_2 \U891/U1117_2_/U3  ( .x(\b[2] ), .a(\U891/U1117_2_/n2 ) );
    nor3_1 \U891/U1117_3_/Unr  ( .x(\U891/U1117_3_/nr ), .a(i[3]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_3_/Und  ( .x(\U891/U1117_3_/nd ), .a(i[3]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_3_/U1  ( .x(\U891/U1117_3_/n2 ), .a(\U891/U1117_3_/n2 ), 
        .b(\U891/U1117_3_/nr ), .c(\U891/U1117_3_/nd ) );
    inv_2 \U891/U1117_3_/U3  ( .x(\b[3] ), .a(\U891/U1117_3_/n2 ) );
    inv_1 \U886/U1126/U3  ( .x(\U886/reset ), .a(nbReset) );
    nor3_1 \U886/U1128/U27  ( .x(\U886/U1128/nb ), .a(\U886/reset ), .b(\f[3] 
        ), .c(\f[2] ) );
    nor2_1 \U886/U1128/U26  ( .x(\U886/U1128/na ), .a(\f[1] ), .b(\f[0] ) );
    nand2_2 \U886/U1128/U29  ( .x(\U886/ackb ), .a(\U886/U1128/nb ), .b(
        \U886/U1128/na ) );
    nor2_1 \U886/U1108/U5  ( .x(\U886/nack ), .a(\U886/acka ), .b(\U886/ackb )
         );
    nor2_2 \U886/U914/U6  ( .x(nba), .a(\U886/acka ), .b(\U886/ackb ) );
    and4_1 \U886/U1127/U25  ( .x(\U886/U1127/n5 ), .a(\U886/U1127/n1 ), .b(
        \U886/U1127/n2 ), .c(\U886/U1127/n3 ), .d(\U886/U1127/n4 ) );
    inv_1 \U886/U1127/U1  ( .x(\U886/U1127/n1 ), .a(\e[3] ) );
    inv_1 \U886/U1127/U2  ( .x(\U886/U1127/n2 ), .a(\e[2] ) );
    inv_1 \U886/U1127/U3  ( .x(\U886/U1127/n3 ), .a(\e[1] ) );
    inv_1 \U886/U1127/U4  ( .x(\U886/U1127/n4 ), .a(\e[0] ) );
    inv_2 \U886/U1127/U5  ( .x(\U886/acka ), .a(\U886/U1127/n5 ) );
    ao222_2 \U886/U1121/U19/U1/U1  ( .x(fsela), .a(\U886/nack ), .b(fsel), .c(
        \U886/nack ), .d(fsela), .e(fsel), .f(fsela) );
    ao222_2 \U886/U1120/U19/U1/U1  ( .x(esela), .a(esel), .b(\U886/nack ), .c(
        esel), .d(esela), .e(\U886/nack ), .f(esela) );
    nor3_1 \U886/U1118_0_/Unr  ( .x(\U886/U1118_0_/nr ), .a(\b[0] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_0_/Und  ( .x(\U886/U1118_0_/nd ), .a(\b[0] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_0_/U1  ( .x(\U886/U1118_0_/n2 ), .a(\U886/U1118_0_/n2 ), 
        .b(\U886/U1118_0_/nr ), .c(\U886/U1118_0_/nd ) );
    inv_2 \U886/U1118_0_/U3  ( .x(\e[0] ), .a(\U886/U1118_0_/n2 ) );
    nor3_1 \U886/U1118_1_/Unr  ( .x(\U886/U1118_1_/nr ), .a(\b[1] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_1_/Und  ( .x(\U886/U1118_1_/nd ), .a(\b[1] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_1_/U1  ( .x(\U886/U1118_1_/n2 ), .a(\U886/U1118_1_/n2 ), 
        .b(\U886/U1118_1_/nr ), .c(\U886/U1118_1_/nd ) );
    inv_2 \U886/U1118_1_/U3  ( .x(\e[1] ), .a(\U886/U1118_1_/n2 ) );
    nor3_1 \U886/U1118_2_/Unr  ( .x(\U886/U1118_2_/nr ), .a(\b[2] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_2_/Und  ( .x(\U886/U1118_2_/nd ), .a(\b[2] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_2_/U1  ( .x(\U886/U1118_2_/n2 ), .a(\U886/U1118_2_/n2 ), 
        .b(\U886/U1118_2_/nr ), .c(\U886/U1118_2_/nd ) );
    inv_2 \U886/U1118_2_/U3  ( .x(\e[2] ), .a(\U886/U1118_2_/n2 ) );
    nor3_1 \U886/U1118_3_/Unr  ( .x(\U886/U1118_3_/nr ), .a(\b[3] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_3_/Und  ( .x(\U886/U1118_3_/nd ), .a(\b[3] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_3_/U1  ( .x(\U886/U1118_3_/n2 ), .a(\U886/U1118_3_/n2 ), 
        .b(\U886/U1118_3_/nr ), .c(\U886/U1118_3_/nd ) );
    inv_2 \U886/U1118_3_/U3  ( .x(\e[3] ), .a(\U886/U1118_3_/n2 ) );
    nor3_1 \U886/U1117_0_/Unr  ( .x(\U886/U1117_0_/nr ), .a(\b[0] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_0_/Und  ( .x(\U886/U1117_0_/nd ), .a(\b[0] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_0_/U1  ( .x(\U886/U1117_0_/n2 ), .a(\U886/U1117_0_/n2 ), 
        .b(\U886/U1117_0_/nr ), .c(\U886/U1117_0_/nd ) );
    inv_2 \U886/U1117_0_/U3  ( .x(\f[0] ), .a(\U886/U1117_0_/n2 ) );
    nor3_1 \U886/U1117_1_/Unr  ( .x(\U886/U1117_1_/nr ), .a(\b[1] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_1_/Und  ( .x(\U886/U1117_1_/nd ), .a(\b[1] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_1_/U1  ( .x(\U886/U1117_1_/n2 ), .a(\U886/U1117_1_/n2 ), 
        .b(\U886/U1117_1_/nr ), .c(\U886/U1117_1_/nd ) );
    inv_2 \U886/U1117_1_/U3  ( .x(\f[1] ), .a(\U886/U1117_1_/n2 ) );
    nor3_1 \U886/U1117_2_/Unr  ( .x(\U886/U1117_2_/nr ), .a(\b[2] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_2_/Und  ( .x(\U886/U1117_2_/nd ), .a(\b[2] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_2_/U1  ( .x(\U886/U1117_2_/n2 ), .a(\U886/U1117_2_/n2 ), 
        .b(\U886/U1117_2_/nr ), .c(\U886/U1117_2_/nd ) );
    inv_2 \U886/U1117_2_/U3  ( .x(\f[2] ), .a(\U886/U1117_2_/n2 ) );
    nor3_1 \U886/U1117_3_/Unr  ( .x(\U886/U1117_3_/nr ), .a(\b[3] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_3_/Und  ( .x(\U886/U1117_3_/nd ), .a(\b[3] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_3_/U1  ( .x(\U886/U1117_3_/n2 ), .a(\U886/U1117_3_/n2 ), 
        .b(\U886/U1117_3_/nr ), .c(\U886/U1117_3_/nd ) );
    inv_2 \U886/U1117_3_/U3  ( .x(\f[3] ), .a(\U886/U1117_3_/n2 ) );
    inv_1 \U884/U1126/U3  ( .x(\U884/reset ), .a(nbReset) );
    nor3_1 \U884/U1128/U27  ( .x(\U884/U1128/nb ), .a(\U884/reset ), .b(\d[3] 
        ), .c(\d[2] ) );
    nor2_1 \U884/U1128/U26  ( .x(\U884/U1128/na ), .a(\d[1] ), .b(\d[0] ) );
    nand2_2 \U884/U1128/U29  ( .x(\U884/ackb ), .a(\U884/U1128/nb ), .b(
        \U884/U1128/na ) );
    nor2_1 \U884/U1108/U5  ( .x(\U884/nack ), .a(\U884/acka ), .b(\U884/ackb )
         );
    nor2_2 \U884/U914/U6  ( .x(naa), .a(\U884/acka ), .b(\U884/ackb ) );
    and4_1 \U884/U1127/U25  ( .x(\U884/U1127/n5 ), .a(\U884/U1127/n1 ), .b(
        \U884/U1127/n2 ), .c(\U884/U1127/n3 ), .d(\U884/U1127/n4 ) );
    inv_1 \U884/U1127/U1  ( .x(\U884/U1127/n1 ), .a(\c[3] ) );
    inv_1 \U884/U1127/U2  ( .x(\U884/U1127/n2 ), .a(\c[2] ) );
    inv_1 \U884/U1127/U3  ( .x(\U884/U1127/n3 ), .a(\c[1] ) );
    inv_1 \U884/U1127/U4  ( .x(\U884/U1127/n4 ), .a(\c[0] ) );
    inv_2 \U884/U1127/U5  ( .x(\U884/acka ), .a(\U884/U1127/n5 ) );
    ao222_2 \U884/U1121/U19/U1/U1  ( .x(dsela), .a(\U884/nack ), .b(dsel), .c(
        \U884/nack ), .d(dsela), .e(dsel), .f(dsela) );
    ao222_2 \U884/U1120/U19/U1/U1  ( .x(csela), .a(csel), .b(\U884/nack ), .c(
        csel), .d(csela), .e(\U884/nack ), .f(csela) );
    nor3_1 \U884/U1118_0_/Unr  ( .x(\U884/U1118_0_/nr ), .a(\a[0] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_0_/Und  ( .x(\U884/U1118_0_/nd ), .a(\a[0] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_0_/U1  ( .x(\U884/U1118_0_/n2 ), .a(\U884/U1118_0_/n2 ), 
        .b(\U884/U1118_0_/nr ), .c(\U884/U1118_0_/nd ) );
    inv_2 \U884/U1118_0_/U3  ( .x(\c[0] ), .a(\U884/U1118_0_/n2 ) );
    nor3_1 \U884/U1118_1_/Unr  ( .x(\U884/U1118_1_/nr ), .a(\a[1] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_1_/Und  ( .x(\U884/U1118_1_/nd ), .a(\a[1] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_1_/U1  ( .x(\U884/U1118_1_/n2 ), .a(\U884/U1118_1_/n2 ), 
        .b(\U884/U1118_1_/nr ), .c(\U884/U1118_1_/nd ) );
    inv_2 \U884/U1118_1_/U3  ( .x(\c[1] ), .a(\U884/U1118_1_/n2 ) );
    nor3_1 \U884/U1118_2_/Unr  ( .x(\U884/U1118_2_/nr ), .a(\a[2] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_2_/Und  ( .x(\U884/U1118_2_/nd ), .a(\a[2] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_2_/U1  ( .x(\U884/U1118_2_/n2 ), .a(\U884/U1118_2_/n2 ), 
        .b(\U884/U1118_2_/nr ), .c(\U884/U1118_2_/nd ) );
    inv_2 \U884/U1118_2_/U3  ( .x(\c[2] ), .a(\U884/U1118_2_/n2 ) );
    nor3_1 \U884/U1118_3_/Unr  ( .x(\U884/U1118_3_/nr ), .a(\a[3] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_3_/Und  ( .x(\U884/U1118_3_/nd ), .a(\a[3] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_3_/U1  ( .x(\U884/U1118_3_/n2 ), .a(\U884/U1118_3_/n2 ), 
        .b(\U884/U1118_3_/nr ), .c(\U884/U1118_3_/nd ) );
    inv_2 \U884/U1118_3_/U3  ( .x(\c[3] ), .a(\U884/U1118_3_/n2 ) );
    nor3_1 \U884/U1117_0_/Unr  ( .x(\U884/U1117_0_/nr ), .a(\a[0] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_0_/Und  ( .x(\U884/U1117_0_/nd ), .a(\a[0] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_0_/U1  ( .x(\U884/U1117_0_/n2 ), .a(\U884/U1117_0_/n2 ), 
        .b(\U884/U1117_0_/nr ), .c(\U884/U1117_0_/nd ) );
    inv_2 \U884/U1117_0_/U3  ( .x(\d[0] ), .a(\U884/U1117_0_/n2 ) );
    nor3_1 \U884/U1117_1_/Unr  ( .x(\U884/U1117_1_/nr ), .a(\a[1] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_1_/Und  ( .x(\U884/U1117_1_/nd ), .a(\a[1] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_1_/U1  ( .x(\U884/U1117_1_/n2 ), .a(\U884/U1117_1_/n2 ), 
        .b(\U884/U1117_1_/nr ), .c(\U884/U1117_1_/nd ) );
    inv_2 \U884/U1117_1_/U3  ( .x(\d[1] ), .a(\U884/U1117_1_/n2 ) );
    nor3_1 \U884/U1117_2_/Unr  ( .x(\U884/U1117_2_/nr ), .a(\a[2] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_2_/Und  ( .x(\U884/U1117_2_/nd ), .a(\a[2] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_2_/U1  ( .x(\U884/U1117_2_/n2 ), .a(\U884/U1117_2_/n2 ), 
        .b(\U884/U1117_2_/nr ), .c(\U884/U1117_2_/nd ) );
    inv_2 \U884/U1117_2_/U3  ( .x(\d[2] ), .a(\U884/U1117_2_/n2 ) );
    nor3_1 \U884/U1117_3_/Unr  ( .x(\U884/U1117_3_/nr ), .a(\a[3] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_3_/Und  ( .x(\U884/U1117_3_/nd ), .a(\a[3] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_3_/U1  ( .x(\U884/U1117_3_/n2 ), .a(\U884/U1117_3_/n2 ), 
        .b(\U884/U1117_3_/nr ), .c(\U884/U1117_3_/nd ) );
    inv_2 \U884/U1117_3_/U3  ( .x(\d[3] ), .a(\U884/U1117_3_/n2 ) );
    nand2_1 \U888/U1128/U5  ( .x(\U888/s ), .a(\U888/r ), .b(\U888/nback ) );
    nand2_1 \U888/U1103/U5  ( .x(\U888/r ), .a(\U888/naack ), .b(\U888/s ) );
    inv_1 \U888/U1111/U3  ( .x(\U888/reset ), .a(nbReset) );
    inv_1 \U888/U1112/U3  ( .x(\U888/naack ), .a(esela) );
    nor2_1 \U888/U1127/U5  ( .x(\U888/nback ), .a(fsela), .b(\U888/reset ) );
    and2_2 \U888/U1129/U8  ( .x(esel), .a(\U888/nback ), .b(\U888/s ) );
    and2_2 \U888/U1124/U8  ( .x(fsel), .a(\U888/r ), .b(\U888/naack ) );
    nand2_1 \U887/U1128/U5  ( .x(\U887/s ), .a(\U887/r ), .b(\U887/nback ) );
    nand2_1 \U887/U1103/U5  ( .x(\U887/r ), .a(\U887/naack ), .b(\U887/s ) );
    inv_1 \U887/U1111/U3  ( .x(\U887/reset ), .a(nbReset) );
    inv_1 \U887/U1112/U3  ( .x(\U887/naack ), .a(csela) );
    nor2_1 \U887/U1127/U5  ( .x(\U887/nback ), .a(dsela), .b(\U887/reset ) );
    and2_2 \U887/U1129/U8  ( .x(csel), .a(\U887/nback ), .b(\U887/s ) );
    and2_2 \U887/U1124/U8  ( .x(dsel), .a(\U887/r ), .b(\U887/naack ) );
    nand2_1 \U885/U1128/U5  ( .x(\U885/s ), .a(\U885/r ), .b(\U885/nback ) );
    nand2_1 \U885/U1103/U5  ( .x(\U885/r ), .a(\U885/naack ), .b(\U885/s ) );
    inv_1 \U885/U1111/U3  ( .x(\U885/reset ), .a(nbReset) );
    inv_1 \U885/U1112/U3  ( .x(\U885/naack ), .a(asela) );
    nor2_1 \U885/U1127/U5  ( .x(\U885/nback ), .a(bsela), .b(\U885/reset ) );
    and2_2 \U885/U1129/U8  ( .x(asel), .a(\U885/nback ), .b(\U885/s ) );
    and2_2 \U885/U1124/U8  ( .x(bsel), .a(\U885/r ), .b(\U885/naack ) );
    nor3_1 \U877/U594/U7  ( .x(\U877/x ), .a(ol[7]), .b(\U877/reset ), .c(oh
        [7]) );
    nor3_1 \U877/U593/U7  ( .x(\U877/y ), .a(ol[6]), .b(\U877/reset ), .c(oh
        [6]) );
    inv_1 \U877/U604/U3  ( .x(\U877/reset ), .a(nbReset) );
    oa31_1 \U877/U590/U25/U1/Uclr  ( .x(\U877/U590/U25/U1/clr ), .a(net135), 
        .b(\cl[3] ), .c(\cl[1] ), .d(oh[6]) );
    oaoi211_1 \U877/U590/U25/U1/Uaoi  ( .x(\U877/U590/U25/U1/ob ), .a(\cl[3] ), 
        .b(\cl[1] ), .c(n1), .d(\U877/U590/U25/U1/clr ) );
    inv_2 \U877/U590/U25/U1/Ui  ( .x(oh[6]), .a(\U877/U590/U25/U1/ob ) );
    oa31_1 \U877/U589/U25/U1/Uclr  ( .x(\U877/U589/U25/U1/clr ), .a(net135), 
        .b(\cl[1] ), .c(\cl[0] ), .d(ol[7]) );
    oaoi211_1 \U877/U589/U25/U1/Uaoi  ( .x(\U877/U589/U25/U1/ob ), .a(\cl[1] ), 
        .b(\cl[0] ), .c(n1), .d(\U877/U589/U25/U1/clr ) );
    inv_2 \U877/U589/U25/U1/Ui  ( .x(ol[7]), .a(\U877/U589/U25/U1/ob ) );
    oa31_1 \U877/U588/U25/U1/Uclr  ( .x(\U877/U588/U25/U1/clr ), .a(net135), 
        .b(\cl[3] ), .c(\cl[2] ), .d(oh[7]) );
    oaoi211_1 \U877/U588/U25/U1/Uaoi  ( .x(\U877/U588/U25/U1/ob ), .a(\cl[3] ), 
        .b(\cl[2] ), .c(n1), .d(\U877/U588/U25/U1/clr ) );
    inv_2 \U877/U588/U25/U1/Ui  ( .x(oh[7]), .a(\U877/U588/U25/U1/ob ) );
    oa31_1 \U877/U591/U25/U1/Uclr  ( .x(\U877/U591/U25/U1/clr ), .a(net135), 
        .b(\cl[2] ), .c(\cl[0] ), .d(ol[6]) );
    oaoi211_1 \U877/U591/U25/U1/Uaoi  ( .x(\U877/U591/U25/U1/ob ), .a(\cl[2] ), 
        .b(\cl[0] ), .c(n1), .d(\U877/U591/U25/U1/clr ) );
    inv_2 \U877/U591/U25/U1/Ui  ( .x(ol[6]), .a(\U877/U591/U25/U1/ob ) );
    ao222_2 \U877/U592/U19/U1/U1  ( .x(ncla), .a(\U877/x ), .b(\U877/y ), .c(
        \U877/x ), .d(ncla), .e(\U877/y ), .f(ncla) );
    nor3_1 \U876/U594/U7  ( .x(\U876/x ), .a(ol[3]), .b(\U876/reset ), .c(oh
        [3]) );
    nor3_1 \U876/U593/U7  ( .x(\U876/y ), .a(ol[2]), .b(\U876/reset ), .c(oh
        [2]) );
    inv_1 \U876/U604/U3  ( .x(\U876/reset ), .a(nbReset) );
    oa31_1 \U876/U590/U25/U1/Uclr  ( .x(\U876/U590/U25/U1/clr ), .a(net135), 
        .b(\d[3] ), .c(\d[1] ), .d(oh[2]) );
    oaoi211_1 \U876/U590/U25/U1/Uaoi  ( .x(\U876/U590/U25/U1/ob ), .a(\d[3] ), 
        .b(\d[1] ), .c(n1), .d(\U876/U590/U25/U1/clr ) );
    inv_2 \U876/U590/U25/U1/Ui  ( .x(oh[2]), .a(\U876/U590/U25/U1/ob ) );
    oa31_1 \U876/U589/U25/U1/Uclr  ( .x(\U876/U589/U25/U1/clr ), .a(net135), 
        .b(\d[1] ), .c(\d[0] ), .d(ol[3]) );
    oaoi211_1 \U876/U589/U25/U1/Uaoi  ( .x(\U876/U589/U25/U1/ob ), .a(\d[1] ), 
        .b(\d[0] ), .c(n1), .d(\U876/U589/U25/U1/clr ) );
    inv_2 \U876/U589/U25/U1/Ui  ( .x(ol[3]), .a(\U876/U589/U25/U1/ob ) );
    oa31_1 \U876/U588/U25/U1/Uclr  ( .x(\U876/U588/U25/U1/clr ), .a(net135), 
        .b(\d[3] ), .c(\d[2] ), .d(oh[3]) );
    oaoi211_1 \U876/U588/U25/U1/Uaoi  ( .x(\U876/U588/U25/U1/ob ), .a(\d[3] ), 
        .b(\d[2] ), .c(n1), .d(\U876/U588/U25/U1/clr ) );
    inv_2 \U876/U588/U25/U1/Ui  ( .x(oh[3]), .a(\U876/U588/U25/U1/ob ) );
    oa31_1 \U876/U591/U25/U1/Uclr  ( .x(\U876/U591/U25/U1/clr ), .a(net135), 
        .b(\d[2] ), .c(\d[0] ), .d(ol[2]) );
    oaoi211_1 \U876/U591/U25/U1/Uaoi  ( .x(\U876/U591/U25/U1/ob ), .a(\d[2] ), 
        .b(\d[0] ), .c(n1), .d(\U876/U591/U25/U1/clr ) );
    inv_2 \U876/U591/U25/U1/Ui  ( .x(ol[2]), .a(\U876/U591/U25/U1/ob ) );
    ao222_2 \U876/U592/U19/U1/U1  ( .x(nda), .a(\U876/x ), .b(\U876/y ), .c(
        \U876/x ), .d(nda), .e(\U876/y ), .f(nda) );
    nor3_1 \U2/U594/U7  ( .x(\U2/x ), .a(ol[1]), .b(\U2/reset ), .c(oh[1]) );
    nor3_1 \U2/U593/U7  ( .x(\U2/y ), .a(ol[0]), .b(\U2/reset ), .c(oh[0]) );
    inv_1 \U2/U604/U3  ( .x(\U2/reset ), .a(nbReset) );
    oa31_1 \U2/U590/U25/U1/Uclr  ( .x(\U2/U590/U25/U1/clr ), .a(net135), .b(
        \f[3] ), .c(\f[1] ), .d(oh[0]) );
    oaoi211_1 \U2/U590/U25/U1/Uaoi  ( .x(\U2/U590/U25/U1/ob ), .a(\f[3] ), .b(
        \f[1] ), .c(n1), .d(\U2/U590/U25/U1/clr ) );
    inv_2 \U2/U590/U25/U1/Ui  ( .x(oh[0]), .a(\U2/U590/U25/U1/ob ) );
    oa31_1 \U2/U589/U25/U1/Uclr  ( .x(\U2/U589/U25/U1/clr ), .a(net135), .b(
        \f[1] ), .c(\f[0] ), .d(ol[1]) );
    oaoi211_1 \U2/U589/U25/U1/Uaoi  ( .x(\U2/U589/U25/U1/ob ), .a(\f[1] ), .b(
        \f[0] ), .c(n1), .d(\U2/U589/U25/U1/clr ) );
    inv_2 \U2/U589/U25/U1/Ui  ( .x(ol[1]), .a(\U2/U589/U25/U1/ob ) );
    oa31_1 \U2/U588/U25/U1/Uclr  ( .x(\U2/U588/U25/U1/clr ), .a(net135), .b(
        \f[3] ), .c(\f[2] ), .d(oh[1]) );
    oaoi211_1 \U2/U588/U25/U1/Uaoi  ( .x(\U2/U588/U25/U1/ob ), .a(\f[3] ), .b(
        \f[2] ), .c(n1), .d(\U2/U588/U25/U1/clr ) );
    inv_2 \U2/U588/U25/U1/Ui  ( .x(oh[1]), .a(\U2/U588/U25/U1/ob ) );
    oa31_1 \U2/U591/U25/U1/Uclr  ( .x(\U2/U591/U25/U1/clr ), .a(net135), .b(
        \f[2] ), .c(\f[0] ), .d(ol[0]) );
    oaoi211_1 \U2/U591/U25/U1/Uaoi  ( .x(\U2/U591/U25/U1/ob ), .a(\f[2] ), .b(
        \f[0] ), .c(n1), .d(\U2/U591/U25/U1/clr ) );
    inv_2 \U2/U591/U25/U1/Ui  ( .x(ol[0]), .a(\U2/U591/U25/U1/ob ) );
    ao222_2 \U2/U592/U19/U1/U1  ( .x(nfa), .a(\U2/x ), .b(\U2/y ), .c(\U2/x ), 
        .d(nfa), .e(\U2/y ), .f(nfa) );
    nor3_1 \U1/U594/U7  ( .x(\U1/x ), .a(ol[5]), .b(\U1/reset ), .c(oh[5]) );
    nor3_1 \U1/U593/U7  ( .x(\U1/y ), .a(ol[4]), .b(\U1/reset ), .c(oh[4]) );
    inv_1 \U1/U604/U3  ( .x(\U1/reset ), .a(nbReset) );
    oa31_1 \U1/U590/U25/U1/Uclr  ( .x(\U1/U590/U25/U1/clr ), .a(net135), .b(
        \e[3] ), .c(\e[1] ), .d(oh[4]) );
    oaoi211_1 \U1/U590/U25/U1/Uaoi  ( .x(\U1/U590/U25/U1/ob ), .a(\e[3] ), .b(
        \e[1] ), .c(n1), .d(\U1/U590/U25/U1/clr ) );
    inv_2 \U1/U590/U25/U1/Ui  ( .x(oh[4]), .a(\U1/U590/U25/U1/ob ) );
    oa31_1 \U1/U589/U25/U1/Uclr  ( .x(\U1/U589/U25/U1/clr ), .a(net135), .b(
        \e[1] ), .c(\e[0] ), .d(ol[5]) );
    oaoi211_1 \U1/U589/U25/U1/Uaoi  ( .x(\U1/U589/U25/U1/ob ), .a(\e[1] ), .b(
        \e[0] ), .c(n1), .d(\U1/U589/U25/U1/clr ) );
    inv_2 \U1/U589/U25/U1/Ui  ( .x(ol[5]), .a(\U1/U589/U25/U1/ob ) );
    oa31_1 \U1/U588/U25/U1/Uclr  ( .x(\U1/U588/U25/U1/clr ), .a(net135), .b(
        \e[3] ), .c(\e[2] ), .d(oh[5]) );
    oaoi211_1 \U1/U588/U25/U1/Uaoi  ( .x(\U1/U588/U25/U1/ob ), .a(\e[3] ), .b(
        \e[2] ), .c(n1), .d(\U1/U588/U25/U1/clr ) );
    inv_2 \U1/U588/U25/U1/Ui  ( .x(oh[5]), .a(\U1/U588/U25/U1/ob ) );
    oa31_1 \U1/U591/U25/U1/Uclr  ( .x(\U1/U591/U25/U1/clr ), .a(net135), .b(
        \e[2] ), .c(\e[0] ), .d(ol[4]) );
    oaoi211_1 \U1/U591/U25/U1/Uaoi  ( .x(\U1/U591/U25/U1/ob ), .a(\e[2] ), .b(
        \e[0] ), .c(n1), .d(\U1/U591/U25/U1/clr ) );
    inv_2 \U1/U591/U25/U1/Ui  ( .x(ol[4]), .a(\U1/U591/U25/U1/ob ) );
    ao222_2 \U1/U592/U19/U1/U1  ( .x(nea), .a(\U1/x ), .b(\U1/y ), .c(\U1/x ), 
        .d(nea), .e(\U1/y ), .f(nea) );
    and3_4 \U881/U20/U9  ( .x(nca), .a(\U881/nack[1] ), .b(\U881/nack[0] ), 
        .c(nbReset) );
    nor2_1 \U881/U18/U5  ( .x(\U881/nack[0] ), .a(\cl[3] ), .b(\cl[0] ) );
    nor2_1 \U881/U19/U5  ( .x(\U881/nack[1] ), .a(\cl[1] ), .b(\cl[2] ) );
    ao222_2 \U881/U15_0_/U19/U1/U1  ( .x(\cl[0] ), .a(\c[0] ), .b(ncla), .c(
        \c[0] ), .d(\cl[0] ), .e(ncla), .f(\cl[0] ) );
    ao222_2 \U881/U15_1_/U19/U1/U1  ( .x(\cl[1] ), .a(\c[1] ), .b(ncla), .c(
        \c[1] ), .d(\cl[1] ), .e(ncla), .f(\cl[1] ) );
    ao222_2 \U881/U15_2_/U19/U1/U1  ( .x(\cl[2] ), .a(\c[2] ), .b(ncla), .c(
        \c[2] ), .d(\cl[2] ), .e(ncla), .f(\cl[2] ) );
    ao222_2 \U881/U15_3_/U19/U1/U1  ( .x(\cl[3] ), .a(\c[3] ), .b(ncla), .c(
        \c[3] ), .d(\cl[3] ), .e(ncla), .f(\cl[3] ) );
    and2_5 U1 ( .x(n1), .a(nbReset), .b(noa) );
    and2_3 U2 ( .x(net135), .a(nbReset), .b(noa) );
endmodule


module chain_ic_ctrl_0 ( ack, candefer, eop, nstatack, pltxreq, routetxreq, 
    tok_ack, accept, candefer_ack, defer, eopack, lock, nReset, pltxack, 
    routetxack, tok_err, tok_ok );
input  [1:0] candefer_ack;
input  [1:0] lock;
input  accept, defer, eopack, nReset, pltxack, routetxack, tok_err, tok_ok;
output ack, candefer, eop, nstatack, pltxreq, routetxreq, tok_ack;
    wire net23, net25, net6, net19, net9, retry, net31, net24, net28, net27, 
        net7, net18, net13, net8, net11, net15, \U249/n5 , \U249/n1 , 
        \U249/n2 , \U249/n3 , \U249/n4 , txnodefer, net16, reset, net17, net29, 
        net12, txmaydefer, nlclear, net4, net22, net14, txlocked, net3, 
        \U286/U28/U1/clr , n1, \U286/U28/U1/set , \U285/U28/U1/clr , n2, 
        \U285/U28/U1/set , txunlocked, net2, txdone, net5, lockcleared, 
        \U262/U25/U1/clr , \U262/U25/U1/ob , \U284/U25/U1/clr , 
        \U284/U25/U1/ob , \U283/U25/U1/clr , net10, \U283/U25/U1/ob , net20, 
        \U289/Z , net21, \U287/Z , \U288/Z , \U149/nr , net30, \U149/nd , 
        \U149/n2 , \locked[0] , \locked[1] , lwrite, \U160/acb , net26, 
        \U160/U1/Z , \U136/nclear_latch , \U136/nwl , \U136/nulsense , 
        \U136/nlsense , \U136/nwh ;
    nand2_1 \U146/U5  ( .x(candefer), .a(net23), .b(net25) );
    or2_1 \U277/U12  ( .x(net6), .a(net19), .b(net9) );
    or2_1 \U264/U12  ( .x(retry), .a(net31), .b(net24) );
    or2_1 \U259/U12  ( .x(net28), .a(net27), .b(net7) );
    or2_1 \U140/U12  ( .x(net18), .a(net13), .b(net8) );
    or2_1 \U148/U12  ( .x(net11), .a(net15), .b(routetxack) );
    and4_1 \U249/U16  ( .x(\U249/n5 ), .a(\U249/n1 ), .b(\U249/n2 ), .c(
        \U249/n3 ), .d(\U249/n4 ) );
    inv_1 \U249/U1  ( .x(\U249/n1 ), .a(txnodefer) );
    inv_1 \U249/U2  ( .x(\U249/n2 ), .a(net16) );
    inv_1 \U249/U3  ( .x(\U249/n3 ), .a(net9) );
    inv_1 \U249/U4  ( .x(\U249/n4 ), .a(net19) );
    inv_1 \U249/U5  ( .x(ack), .a(\U249/n5 ) );
    nor3_2 \U40/U16  ( .x(nstatack), .a(net16), .b(reset), .c(retry) );
    nor3_2 \U275/U16  ( .x(net17), .a(net29), .b(reset), .c(tok_ack) );
    buf_3 \U290/U8  ( .x(net12), .a(txmaydefer) );
    nor2_1 \U154/U5  ( .x(nlclear), .a(net4), .b(net31) );
    or2_2 \U274/U12  ( .x(pltxreq), .a(net22), .b(net14) );
    or3_1 \U260/U12  ( .x(eop), .a(net31), .b(txlocked), .c(net4) );
    inv_1 \U147/U3  ( .x(net3), .a(net29) );
    inv_1 \U174/U3  ( .x(reset), .a(nReset) );
    aoai211_1 \U286/U28/U1/U1  ( .x(\U286/U28/U1/clr ), .a(net3), .b(n1), .c(
        net17), .d(net22) );
    nand3_1 \U286/U28/U1/U2  ( .x(\U286/U28/U1/set ), .a(net17), .b(net3), .c(
        n1) );
    nand2_2 \U286/U28/U1/U3  ( .x(net22), .a(\U286/U28/U1/clr ), .b(
        \U286/U28/U1/set ) );
    aoai211_1 \U285/U28/U1/U1  ( .x(\U285/U28/U1/clr ), .a(net3), .b(n2), .c(
        net17), .d(net14) );
    nand3_1 \U285/U28/U1/U2  ( .x(\U285/U28/U1/set ), .a(net17), .b(net3), .c(
        n2) );
    nand2_2 \U285/U28/U1/U3  ( .x(net14), .a(\U285/U28/U1/clr ), .b(
        \U285/U28/U1/set ) );
    ao222_1 \U254/U18/U1/U1  ( .x(net31), .a(defer), .b(txunlocked), .c(defer), 
        .d(net31), .e(txunlocked), .f(net31) );
    ao222_1 \U252/U18/U1/U1  ( .x(net19), .a(tok_err), .b(net12), .c(tok_err), 
        .d(net19), .e(net12), .f(net19) );
    ao222_1 \U276/U18/U1/U1  ( .x(net24), .a(txlocked), .b(defer), .c(txlocked
        ), .d(net24), .e(defer), .f(net24) );
    ao222_1 \U251/U18/U1/U1  ( .x(net9), .a(tok_ok), .b(net12), .c(tok_ok), 
        .d(net9), .e(net12), .f(net9) );
    ao222_1 \U235/U18/U1/U1  ( .x(tok_ack), .a(ack), .b(net2), .c(ack), .d(
        tok_ack), .e(net2), .f(tok_ack) );
    ao222_1 \U247/U18/U1/U1  ( .x(txnodefer), .a(txdone), .b(candefer_ack[0]), 
        .c(txdone), .d(txnodefer), .e(candefer_ack[0]), .f(txnodefer) );
    ao222_2 \U246/U19/U1/U1  ( .x(txlocked), .a(net14), .b(txdone), .c(net14), 
        .d(txlocked), .e(txdone), .f(txlocked) );
    ao222_2 \U245/U19/U1/U1  ( .x(txunlocked), .a(txdone), .b(net22), .c(
        txdone), .d(txunlocked), .e(net22), .f(txunlocked) );
    ao222_1 \U269/U18/U1/U1  ( .x(net2), .a(net28), .b(net18), .c(net28), .d(
        net2), .e(net18), .f(net2) );
    ao222_1 \U268/U18/U1/U1  ( .x(net5), .a(eopack), .b(lockcleared), .c(
        eopack), .d(net5), .e(lockcleared), .f(net5) );
    ao222_1 \U256/U18/U1/U1  ( .x(net4), .a(tok_err), .b(txunlocked), .c(
        tok_err), .d(net4), .e(txunlocked), .f(net4) );
    ao222_1 \U175/U18/U1/U1  ( .x(net29), .a(net2), .b(retry), .c(net2), .d(
        net29), .e(retry), .f(net29) );
    ao222_1 \U255/U18/U1/U1  ( .x(net8), .a(txlocked), .b(eopack), .c(txlocked
        ), .d(net8), .e(eopack), .f(net8) );
    ao222_2 \U248/U19/U1/U1  ( .x(txmaydefer), .a(candefer_ack[1]), .b(txdone), 
        .c(candefer_ack[1]), .d(txmaydefer), .e(txdone), .f(txmaydefer) );
    ao222_2 \U250/U19/U1/U1  ( .x(net16), .a(accept), .b(net12), .c(accept), 
        .d(net16), .e(net12), .f(net16) );
    oa31_1 \U262/U25/U1/Uclr  ( .x(\U262/U25/U1/clr ), .a(txunlocked), .b(net5
        ), .c(tok_ok), .d(net13) );
    oaoi211_1 \U262/U25/U1/Uaoi  ( .x(\U262/U25/U1/ob ), .a(net5), .b(tok_ok), 
        .c(txunlocked), .d(\U262/U25/U1/clr ) );
    inv_2 \U262/U25/U1/Ui  ( .x(net13), .a(\U262/U25/U1/ob ) );
    oa31_1 \U284/U25/U1/Uclr  ( .x(\U284/U25/U1/clr ), .a(txnodefer), .b(
        tok_ok), .c(tok_err), .d(net27) );
    oaoi211_1 \U284/U25/U1/Uaoi  ( .x(\U284/U25/U1/ob ), .a(tok_ok), .b(
        tok_err), .c(txnodefer), .d(\U284/U25/U1/clr ) );
    inv_2 \U284/U25/U1/Ui  ( .x(net27), .a(\U284/U25/U1/ob ) );
    oa31_1 \U283/U25/U1/Uclr  ( .x(\U283/U25/U1/clr ), .a(net10), .b(net6), 
        .c(retry), .d(net7) );
    oaoi211_1 \U283/U25/U1/Uaoi  ( .x(\U283/U25/U1/ob ), .a(net6), .b(retry), 
        .c(net10), .d(\U283/U25/U1/clr ) );
    inv_2 \U283/U25/U1/Ui  ( .x(net7), .a(\U283/U25/U1/ob ) );
    aoi21_1 \U289/U30/U1/U1  ( .x(net20), .a(\U289/Z ), .b(net16), .c(net12)
         );
    inv_1 \U289/U30/U1/U2  ( .x(\U289/Z ), .a(net20) );
    aoi21_1 \U287/U30/U1/U1  ( .x(net21), .a(\U287/Z ), .b(accept), .c(net12)
         );
    inv_1 \U287/U30/U1/U2  ( .x(\U287/Z ), .a(net21) );
    aoi222_1 \U288/U30/U1  ( .x(net10), .a(net20), .b(net21), .c(net20), .d(
        \U288/Z ), .e(net21), .f(\U288/Z ) );
    inv_1 \U288/U30/Uinv  ( .x(\U288/Z ), .a(net10) );
    nor3_1 \U149/Unr  ( .x(\U149/nr ), .a(pltxack), .b(net11), .c(net30) );
    nand3_1 \U149/Und  ( .x(\U149/nd ), .a(pltxack), .b(net11), .c(net30) );
    oa21_1 \U149/U1  ( .x(\U149/n2 ), .a(\U149/n2 ), .b(\U149/nr ), .c(
        \U149/nd ) );
    inv_2 \U149/U3  ( .x(txdone), .a(\U149/n2 ) );
    inv_1 \U133/U618/U3  ( .x(net23), .a(net15) );
    inv_1 \U133/U617/U3  ( .x(net25), .a(routetxreq) );
    ao23_1 \U133/U616/U21/U1/U1  ( .x(routetxreq), .a(pltxreq), .b(routetxreq), 
        .c(pltxreq), .d(\locked[0] ), .e(net23) );
    ao23_1 \U133/U615/U21/U1/U1  ( .x(net15), .a(pltxreq), .b(net15), .c(
        pltxreq), .d(\locked[1] ), .e(net25) );
    and2_1 \U160/U2/U8  ( .x(lwrite), .a(candefer), .b(\U160/acb ) );
    nor2_1 \U160/U3/U5  ( .x(net30), .a(\U160/acb ), .b(net26) );
    oai21_1 \U160/U1/U30/U1/U1  ( .x(\U160/acb ), .a(\U160/U1/Z ), .b(net26), 
        .c(candefer) );
    inv_1 \U160/U1/U30/U1/U2  ( .x(\U160/U1/Z ), .a(\U160/acb ) );
    nand3_2 \U136/U48/U16  ( .x(\locked[0] ), .a(\locked[1] ), .b(
        \U136/nclear_latch ), .c(\U136/nwl ) );
    nor2_0 \U136/U36/U5  ( .x(\U136/nulsense ), .a(\locked[1] ), .b(\U136/nwl 
        ) );
    nor2_0 \U136/U37/U5  ( .x(\U136/nlsense ), .a(\U136/nwh ), .b(\locked[0] )
         );
    and2_1 \U136/U76/U8  ( .x(\U136/nclear_latch ), .a(nReset), .b(nlclear) );
    nor2_1 \U136/U77/U5  ( .x(lockcleared), .a(nlclear), .b(\locked[1] ) );
    nand2_1 \U136/U14/U5  ( .x(\U136/nwl ), .a(lwrite), .b(n2) );
    nand2_1 \U136/U15/U5  ( .x(\U136/nwh ), .a(n1), .b(lwrite) );
    nand2_2 \U136/U47/U5  ( .x(\locked[1] ), .a(\U136/nwh ), .b(\locked[0] )
         );
    or2_4 \U136/U35/U12  ( .x(net26), .a(\U136/nlsense ), .b(\U136/nulsense )
         );
    buf_1 U1 ( .x(n1), .a(lock[1]) );
    buf_1 U2 ( .x(n2), .a(lock[0]) );
endmodule


module chain_selement_ga_33 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_34 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_35 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_36 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_40 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_37 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_41 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_38 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_39 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_32 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_dr8bit_completion_50 ( o, i );
input  [15:0] i;
output o;
    wire \nx[0] , \nx[1] , \nx[2] , \nx[3] , \ny[0] , \ny[1] , \ny[2] , 
        \ny[3] , y, x, \U6/Z , \U3/net3 , \U3/U20/Z , \U3/net2 , \U3/U21/Z , 
        \U3/U19/Z , \U5/net3 , \U5/U20/Z , \U5/net2 , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_51 ( o, i );
input  [15:0] i;
output o;
    wire \nx[0] , \nx[1] , \nx[2] , \nx[3] , \ny[0] , \ny[1] , \ny[2] , 
        \ny[3] , y, x, \U6/Z , \U3/net3 , \U3/U20/Z , \U3/net2 , \U3/U21/Z , 
        \U3/U19/Z , \U5/net3 , \U5/U20/Z , \U5/net2 , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_16 ( o, i );
input  [15:0] i;
output o;
    wire \nx[0] , \nx[1] , \nx[2] , \nx[3] , \ny[0] , \ny[1] , \ny[2] , 
        \ny[3] , y, x, \U6/Z , \U3/net3 , \U3/U20/Z , \U3/net2 , \U3/U21/Z , 
        \U3/U19/Z , \U5/net3 , \U5/U20/Z , \U5/net2 , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_19 ( o, i );
input  [15:0] i;
output o;
    wire \nx[0] , \nx[1] , \nx[2] , \nx[3] , \ny[0] , \ny[1] , \ny[2] , 
        \ny[3] , y, x, \U6/Z , \U3/net3 , \U3/U20/Z , \U3/net2 , \U3/U21/Z , 
        \U3/U19/Z , \U5/net3 , \U5/U20/Z , \U5/net2 , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_18 ( o, i );
input  [15:0] i;
output o;
    wire \nx[0] , \nx[1] , \nx[2] , \nx[3] , \ny[0] , \ny[1] , \ny[2] , 
        \ny[3] , y, x, \U6/Z , \U3/net3 , \U3/U20/Z , \U3/net2 , \U3/U21/Z , 
        \U3/U19/Z , \U5/net3 , \U5/U20/Z , \U5/net2 , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_17 ( o, i );
input  [15:0] i;
output o;
    wire \nx[0] , \nx[1] , \nx[2] , \nx[3] , \ny[0] , \ny[1] , \ny[2] , 
        \ny[3] , y, x, \U6/Z , \U3/net3 , \U3/U20/Z , \U3/net2 , \U3/U21/Z , 
        \U3/U19/Z , \U5/net3 , \U5/U20/Z , \U5/net2 , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr32bit_completion_2 ( o, i );
input  [63:0] i;
output o;
    wire \cd[3] , \cd[2] , \cd[1] , \cd[0] , ny, \U16/Z , nx, \U6/Z , \U15/Z ;
    chain_dr8bit_completion_16 U11 ( .o(\cd[3] ), .i({i[63], i[62], i[61], 
        i[60], i[59], i[58], i[57], i[56], i[31], i[30], i[29], i[28], i[27], 
        i[26], i[25], i[24]}) );
    chain_dr8bit_completion_19 U14 ( .o(\cd[2] ), .i({i[55], i[54], i[53], 
        i[52], i[51], i[50], i[49], i[48], i[23], i[22], i[21], i[20], i[19], 
        i[18], i[17], i[16]}) );
    chain_dr8bit_completion_18 U13 ( .o(\cd[1] ), .i({i[47], i[46], i[45], 
        i[44], i[43], i[42], i[41], i[40], i[15], i[14], i[13], i[12], i[11], 
        i[10], i[9], i[8]}) );
    chain_dr8bit_completion_17 U12 ( .o(\cd[0] ), .i({i[39], i[38], i[37], 
        i[36], i[35], i[34], i[33], i[32], i[7], i[6], i[5], i[4], i[3], i[2], 
        i[1], i[0]}) );
    aoi222_1 \U16/U30/U1  ( .x(ny), .a(\cd[0] ), .b(\cd[1] ), .c(\cd[0] ), .d(
        \U16/Z ), .e(\cd[1] ), .f(\U16/Z ) );
    inv_1 \U16/U30/Uinv  ( .x(\U16/Z ), .a(ny) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(ny), .b(nx), .c(ny), .d(\U6/Z ), .e(nx), 
        .f(\U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U15/U30/U1  ( .x(nx), .a(\cd[3] ), .b(\cd[2] ), .c(\cd[3] ), .d(
        \U15/Z ), .e(\cd[2] ), .f(\U15/Z ) );
    inv_1 \U15/U30/Uinv  ( .x(\U15/Z ), .a(nx) );
endmodule


module chain_dr8bit_completion_20 ( o, i );
input  [15:0] i;
output o;
    wire \nx[0] , \nx[1] , \nx[2] , \nx[3] , \ny[0] , \ny[1] , \ny[2] , 
        \ny[3] , y, x, \U6/Z , \U3/net3 , \U3/U20/Z , \U3/net2 , \U3/U21/Z , 
        \U3/U19/Z , \U5/net3 , \U5/U20/Z , \U5/net2 , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_23 ( o, i );
input  [15:0] i;
output o;
    wire \nx[0] , \nx[1] , \nx[2] , \nx[3] , \ny[0] , \ny[1] , \ny[2] , 
        \ny[3] , y, x, \U6/Z , \U3/net3 , \U3/U20/Z , \U3/net2 , \U3/U21/Z , 
        \U3/U19/Z , \U5/net3 , \U5/U20/Z , \U5/net2 , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_22 ( o, i );
input  [15:0] i;
output o;
    wire \nx[0] , \nx[1] , \nx[2] , \nx[3] , \ny[0] , \ny[1] , \ny[2] , 
        \ny[3] , y, x, \U6/Z , \U3/net3 , \U3/U20/Z , \U3/net2 , \U3/U21/Z , 
        \U3/U19/Z , \U5/net3 , \U5/U20/Z , \U5/net2 , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_21 ( o, i );
input  [15:0] i;
output o;
    wire \nx[0] , \nx[1] , \nx[2] , \nx[3] , \ny[0] , \ny[1] , \ny[2] , 
        \ny[3] , y, x, \U6/Z , \U3/net3 , \U3/U20/Z , \U3/net2 , \U3/U21/Z , 
        \U3/U19/Z , \U5/net3 , \U5/U20/Z , \U5/net2 , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr32bit_completion_3 ( o, i );
input  [63:0] i;
output o;
    wire \cd[3] , \cd[2] , \cd[1] , \cd[0] , ny, \U16/Z , nx, \U6/Z , \U15/Z ;
    chain_dr8bit_completion_20 U11 ( .o(\cd[3] ), .i({i[63], i[62], i[61], 
        i[60], i[59], i[58], i[57], i[56], i[31], i[30], i[29], i[28], i[27], 
        i[26], i[25], i[24]}) );
    chain_dr8bit_completion_23 U14 ( .o(\cd[2] ), .i({i[55], i[54], i[53], 
        i[52], i[51], i[50], i[49], i[48], i[23], i[22], i[21], i[20], i[19], 
        i[18], i[17], i[16]}) );
    chain_dr8bit_completion_22 U13 ( .o(\cd[1] ), .i({i[47], i[46], i[45], 
        i[44], i[43], i[42], i[41], i[40], i[15], i[14], i[13], i[12], i[11], 
        i[10], i[9], i[8]}) );
    chain_dr8bit_completion_21 U12 ( .o(\cd[0] ), .i({i[39], i[38], i[37], 
        i[36], i[35], i[34], i[33], i[32], i[7], i[6], i[5], i[4], i[3], i[2], 
        i[1], i[0]}) );
    aoi222_1 \U16/U30/U1  ( .x(ny), .a(\cd[0] ), .b(\cd[1] ), .c(\cd[0] ), .d(
        \U16/Z ), .e(\cd[1] ), .f(\U16/Z ) );
    inv_1 \U16/U30/Uinv  ( .x(\U16/Z ), .a(ny) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(ny), .b(nx), .c(ny), .d(\U6/Z ), .e(nx), 
        .f(\U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U15/U30/U1  ( .x(nx), .a(\cd[3] ), .b(\cd[2] ), .c(\cd[3] ), .d(
        \U15/Z ), .e(\cd[2] ), .f(\U15/Z ) );
    inv_1 \U15/U30/Uinv  ( .x(\U15/Z ), .a(nx) );
endmodule


module chain_icmux_0 ( ack, chainh, chainl, sendack, addr, col, itag, lock, 
    nReset, nia, pred, rnw, sendreq, seq, size, wd );
output [7:0] chainh;
output [7:0] chainl;
input  [63:0] addr;
input  [5:0] col;
input  [9:0] itag;
input  [1:0] lock;
input  [1:0] pred;
input  [1:0] rnw;
input  [1:0] seq;
input  [3:0] size;
input  [63:0] wd;
input  nReset, nia, sendreq;
output ack, sendack;
    wire net152, net146, net148, n1, net156, \bs[1] , net138, net160, \bs[2] , 
        net168, \bs[3] , net172, \bs[7] , net164, net132, \bs[4] , net289, 
        \bs[8] , net180, \bs[5] , net176, \bs[6] , \bs[0] , \hdr[4] , net185, 
        net187, net189, net191, net293, net131, \net246[15] , net265, 
        \net246[14] , \net246[13] , \net246[12] , \net246[11] , \net246[10] , 
        \net246[9] , \net246[8] , \net246[7] , \net246[6] , \net246[5] , 
        \net246[4] , \net246[3] , \net246[2] , \net246[1] , \net246[0] , 
        \net243[15] , net263, \net243[14] , \net243[13] , \net243[12] , 
        \net243[11] , \net243[10] , \net243[9] , \net243[8] , \net243[7] , 
        \net243[6] , \net243[5] , \net243[4] , \net243[3] , \net243[2] , 
        \net243[1] , \net243[0] , \net240[15] , net267, \net240[14] , 
        \net240[13] , \net240[12] , \net240[11] , \net240[10] , \net240[9] , 
        \net240[8] , \net240[7] , \net240[6] , \net240[5] , \net240[4] , 
        \net240[3] , \net240[2] , \net240[1] , \net240[0] , \net237[15] , 
        net269, \net237[14] , \net237[13] , \net237[12] , \net237[11] , 
        \net237[10] , \net237[9] , \net237[8] , \net237[7] , \net237[6] , 
        \net237[5] , \net237[2] , \net237[1] , \net237[0] , \net234[15] , 
        net259, \net234[14] , \net234[13] , \net234[12] , \net234[11] , 
        \net234[10] , \net234[9] , \net234[8] , \net234[7] , \net234[6] , 
        \net234[5] , \net234[4] , \net234[3] , \net234[2] , \net234[1] , 
        \net234[0] , \net231[15] , net253, \net231[14] , \net231[13] , 
        \net231[12] , \net231[11] , \net231[10] , \net231[9] , \net231[8] , 
        \net231[7] , \net231[6] , \net231[5] , \net231[4] , \net231[3] , 
        \net231[2] , \net231[1] , \net231[0] , \net228[15] , net255, 
        \net228[14] , \net228[13] , \net228[12] , \net228[11] , \net228[10] , 
        \net228[9] , \net228[8] , \net228[7] , \net228[6] , \net228[5] , 
        \net228[4] , \net228[3] , \net228[2] , \net228[1] , \net228[0] , 
        \net225[15] , net251, \net225[14] , \net225[13] , \net225[12] , 
        \net225[11] , \net225[10] , \net225[9] , \net225[8] , \net225[7] , 
        \net225[6] , \net225[5] , \net225[4] , \net225[3] , \net225[2] , 
        \net225[1] , \net225[0] , \net222[15] , net261, \net222[14] , 
        \net222[13] , \net222[12] , \net222[11] , \net222[10] , \net222[9] , 
        \net222[8] , \net222[7] , \net222[6] , \net222[5] , \net222[4] , 
        \net222[3] , \net222[2] , \net222[1] , \net222[0] , \net219[15] , 
        net249, \net219[14] , \net219[13] , \net219[12] , \net219[11] , 
        \net219[10] , \net219[9] , \net219[8] , \net219[7] , \net219[6] , 
        \net219[5] , \net219[4] , \net219[3] , \net219[2] , \net219[1] , 
        \net219[0] , \U40_0_/n3 , \U40_0_/n4 , \net217[15] , \U40_0_/n5 , 
        \U40_1_/n3 , \U40_1_/n4 , \net217[14] , \U40_1_/n5 , \U40_2_/n3 , 
        \U40_2_/n4 , \net217[13] , \U40_2_/n5 , \U40_3_/n3 , \U40_3_/n4 , 
        \net217[12] , \U40_3_/n5 , \U40_4_/n3 , \U40_4_/n4 , \net217[11] , 
        \U40_4_/n5 , \U40_5_/n3 , \U40_5_/n4 , \net217[10] , \U40_5_/n5 , 
        \U40_6_/n3 , \U40_6_/n4 , \net217[9] , \U40_6_/n5 , \U40_7_/n3 , 
        \U40_7_/n4 , \net217[8] , \U40_7_/n5 , \U40_8_/n3 , \U40_8_/n4 , 
        \net217[7] , \U40_8_/n5 , \U40_9_/n3 , \U40_9_/n4 , \net217[6] , 
        \U40_9_/n5 , \U40_10_/n3 , \U40_10_/n4 , \net217[5] , \U40_10_/n5 , 
        \U40_11_/n3 , \U40_11_/n4 , \net217[4] , \U40_11_/n5 , \U40_12_/n3 , 
        \U40_12_/n4 , \net217[3] , \U40_12_/n5 , \U40_13_/n3 , \U40_13_/n4 , 
        \net217[2] , \U40_13_/n5 , \U40_14_/n3 , \U40_14_/n4 , \net217[1] , 
        \U40_14_/n5 , \U40_15_/n3 , \U40_15_/n4 , \net217[0] , \U40_15_/n5 , 
        \U14_0_/n5 , \U14_0_/n1 , \U14_0_/n2 , \U14_0_/n3 , \U14_0_/n4 , 
        \net212[15] , \U14_1_/n5 , \U14_1_/n1 , \U14_1_/n2 , \U14_1_/n3 , 
        \U14_1_/n4 , \net212[14] , \U14_2_/n5 , \U14_2_/n1 , \U14_2_/n2 , 
        \U14_2_/n3 , \U14_2_/n4 , \net212[13] , \U14_3_/n5 , \U14_3_/n1 , 
        \U14_3_/n2 , \U14_3_/n3 , \U14_3_/n4 , \net212[12] , \U14_4_/n5 , 
        \U14_4_/n1 , \U14_4_/n2 , \U14_4_/n3 , \U14_4_/n4 , \net212[11] , 
        \U14_5_/n5 , \U14_5_/n1 , \U14_5_/n2 , \U14_5_/n3 , \U14_5_/n4 , 
        \net212[10] , \U14_6_/n5 , \U14_6_/n1 , \U14_6_/n2 , \U14_6_/n3 , 
        \U14_6_/n4 , \net212[9] , \U14_7_/n5 , \U14_7_/n1 , \U14_7_/n2 , 
        \U14_7_/n3 , \U14_7_/n4 , \net212[8] , \U14_8_/n5 , \U14_8_/n1 , 
        \U14_8_/n2 , \U14_8_/n3 , \U14_8_/n4 , \net212[7] , \U14_9_/n5 , 
        \U14_9_/n1 , \U14_9_/n2 , \U14_9_/n3 , \U14_9_/n4 , \net212[6] , 
        \U14_10_/n5 , \U14_10_/n1 , \U14_10_/n2 , \U14_10_/n3 , \U14_10_/n4 , 
        \net212[5] , \U14_11_/n1 , \U14_11_/n2 , \U14_11_/n4 , \net212[4] , 
        \U14_11_/n5 , \U14_12_/n1 , \U14_12_/n2 , \U14_12_/n4 , \net212[3] , 
        \U14_12_/n5 , \U14_13_/n5 , \U14_13_/n1 , \U14_13_/n2 , \U14_13_/n3 , 
        \U14_13_/n4 , \net212[2] , \U14_14_/n5 , \U14_14_/n1 , \U14_14_/n2 , 
        \U14_14_/n3 , \U14_14_/n4 , \net212[1] , \U14_15_/n5 , \U14_15_/n1 , 
        \U14_15_/n2 , \U14_15_/n3 , \U14_15_/n4 , \net212[0] , \U91_0_/n5 , 
        \U91_0_/n1 , \U91_0_/n2 , \U91_0_/n3 , \U91_0_/n4 , \net207[15] , 
        \U91_1_/n5 , \U91_1_/n1 , \U91_1_/n2 , \U91_1_/n3 , \U91_1_/n4 , 
        \net207[14] , \U91_2_/n5 , \U91_2_/n1 , \U91_2_/n2 , \U91_2_/n3 , 
        \U91_2_/n4 , \net207[13] , \U91_3_/n5 , \U91_3_/n1 , \U91_3_/n2 , 
        \U91_3_/n3 , \U91_3_/n4 , \net207[12] , \U91_4_/n5 , \U91_4_/n1 , 
        \U91_4_/n2 , \U91_4_/n3 , \U91_4_/n4 , \net207[11] , \U91_5_/n5 , 
        \U91_5_/n1 , \U91_5_/n2 , \U91_5_/n3 , \U91_5_/n4 , \net207[10] , 
        \U91_6_/n5 , \U91_6_/n1 , \U91_6_/n2 , \U91_6_/n3 , \U91_6_/n4 , 
        \net207[9] , \U91_7_/n5 , \U91_7_/n1 , \U91_7_/n2 , \U91_7_/n3 , 
        \U91_7_/n4 , \net207[8] , \U91_8_/n5 , \U91_8_/n1 , \U91_8_/n2 , 
        \U91_8_/n3 , \U91_8_/n4 , \net207[7] , \U91_9_/n5 , \U91_9_/n1 , 
        \U91_9_/n2 , \U91_9_/n3 , \U91_9_/n4 , \net207[6] , \U91_10_/n5 , 
        \U91_10_/n1 , \U91_10_/n2 , \U91_10_/n3 , \U91_10_/n4 , \net207[5] , 
        \U91_11_/n5 , \U91_11_/n1 , \U91_11_/n2 , \U91_11_/n3 , \U91_11_/n4 , 
        \net207[4] , \U91_12_/n5 , \U91_12_/n1 , \U91_12_/n2 , \U91_12_/n3 , 
        \U91_12_/n4 , \net207[3] , \U91_13_/n5 , \U91_13_/n1 , \U91_13_/n2 , 
        \U91_13_/n3 , \U91_13_/n4 , \net207[2] , \U91_14_/n5 , \U91_14_/n1 , 
        \U91_14_/n2 , \U91_14_/n3 , \U91_14_/n4 , \net207[1] , \U91_15_/n5 , 
        \U91_15_/n1 , \U91_15_/n2 , \U91_15_/n3 , \U91_15_/n4 , \net207[0] , 
        net198, net136, \U151/Z , \U148/U21/nr , \U148/U21/nd , \U148/U21/n2 ;
    chain_selement_ga_33 U163 ( .Aa(net152), .Br(net146), .Ar(net148), .Ba(n1)
         );
    chain_selement_ga_34 U164 ( .Aa(net156), .Br(\bs[1] ), .Ar(net152), .Ba(
        net138) );
    chain_selement_ga_35 U165 ( .Aa(net160), .Br(\bs[2] ), .Ar(net156), .Ba(n1
        ) );
    chain_selement_ga_36 U166 ( .Aa(net168), .Br(\bs[3] ), .Ar(net160), .Ba(
        net138) );
    chain_selement_ga_40 U170 ( .Aa(net172), .Br(\bs[7] ), .Ar(net164), .Ba(
        net138) );
    chain_selement_ga_37 U167 ( .Aa(net132), .Br(\bs[4] ), .Ar(net168), .Ba(
        net138) );
    chain_selement_ga_41 U171 ( .Aa(net289), .Br(\bs[8] ), .Ar(net172), .Ba(
        net138) );
    chain_selement_ga_38 U168 ( .Aa(net180), .Br(\bs[5] ), .Ar(net176), .Ba(
        net138) );
    chain_selement_ga_39 U169 ( .Aa(net164), .Br(\bs[6] ), .Ar(net180), .Ba(n1
        ) );
    chain_selement_ga_32 U161 ( .Aa(net148), .Br(\bs[0] ), .Ar(\hdr[4] ), .Ba(
        n1) );
    chain_dr8bit_completion_50 U119 ( .o(net185), .i({col[5], col[4], col[3], 
        itag[9], itag[8], itag[7], itag[6], itag[5], col[2], col[1], col[0], 
        itag[4], itag[3], itag[2], itag[1], itag[0]}) );
    chain_dr8bit_completion_51 U147 ( .o(net187), .i({size[3], size[2], rnw[1], 
        1'b0, 1'b0, lock[1], pred[1], seq[1], size[1], size[0], rnw[0], 
        \hdr[4] , \hdr[4] , lock[0], pred[0], seq[0]}) );
    chain_dr32bit_completion_2 U117 ( .o(net189), .i(wd) );
    chain_dr32bit_completion_3 U118 ( .o(net191), .i(addr) );
    or2_4 \U122/U12  ( .x(net293), .a(net189), .b(net131) );
    or2_4 \U53/U12  ( .x(sendack), .a(net131), .b(net289) );
    and2_1 \U32_0_/U8  ( .x(\net246[15] ), .a(itag[0]), .b(net265) );
    and2_1 \U32_1_/U8  ( .x(\net246[14] ), .a(itag[1]), .b(net265) );
    and2_1 \U32_2_/U8  ( .x(\net246[13] ), .a(itag[2]), .b(net265) );
    and2_1 \U32_3_/U8  ( .x(\net246[12] ), .a(itag[3]), .b(net265) );
    and2_1 \U32_4_/U8  ( .x(\net246[11] ), .a(itag[4]), .b(net265) );
    and2_1 \U32_5_/U8  ( .x(\net246[10] ), .a(col[0]), .b(net265) );
    and2_1 \U32_6_/U8  ( .x(\net246[9] ), .a(col[1]), .b(net265) );
    and2_1 \U32_7_/U8  ( .x(\net246[8] ), .a(col[2]), .b(net265) );
    and2_1 \U32_8_/U8  ( .x(\net246[7] ), .a(itag[5]), .b(net265) );
    and2_1 \U32_9_/U8  ( .x(\net246[6] ), .a(itag[6]), .b(net265) );
    and2_1 \U32_10_/U8  ( .x(\net246[5] ), .a(itag[7]), .b(net265) );
    and2_1 \U32_11_/U8  ( .x(\net246[4] ), .a(itag[8]), .b(net265) );
    and2_1 \U32_12_/U8  ( .x(\net246[3] ), .a(itag[9]), .b(net265) );
    and2_1 \U32_13_/U8  ( .x(\net246[2] ), .a(col[3]), .b(net265) );
    and2_1 \U32_14_/U8  ( .x(\net246[1] ), .a(col[4]), .b(net265) );
    and2_1 \U32_15_/U8  ( .x(\net246[0] ), .a(col[5]), .b(net265) );
    and2_1 \U76_0_/U8  ( .x(\net243[15] ), .a(wd[8]), .b(net263) );
    and2_1 \U76_1_/U8  ( .x(\net243[14] ), .a(wd[9]), .b(net263) );
    and2_1 \U76_2_/U8  ( .x(\net243[13] ), .a(wd[10]), .b(net263) );
    and2_1 \U76_3_/U8  ( .x(\net243[12] ), .a(wd[11]), .b(net263) );
    and2_1 \U76_4_/U8  ( .x(\net243[11] ), .a(wd[12]), .b(net263) );
    and2_1 \U76_5_/U8  ( .x(\net243[10] ), .a(wd[13]), .b(net263) );
    and2_1 \U76_6_/U8  ( .x(\net243[9] ), .a(wd[14]), .b(net263) );
    and2_1 \U76_7_/U8  ( .x(\net243[8] ), .a(wd[15]), .b(net263) );
    and2_1 \U76_8_/U8  ( .x(\net243[7] ), .a(wd[40]), .b(net263) );
    and2_1 \U76_9_/U8  ( .x(\net243[6] ), .a(wd[41]), .b(net263) );
    and2_1 \U76_10_/U8  ( .x(\net243[5] ), .a(wd[42]), .b(net263) );
    and2_1 \U76_11_/U8  ( .x(\net243[4] ), .a(wd[43]), .b(net263) );
    and2_1 \U76_12_/U8  ( .x(\net243[3] ), .a(wd[44]), .b(net263) );
    and2_1 \U76_13_/U8  ( .x(\net243[2] ), .a(wd[45]), .b(net263) );
    and2_1 \U76_14_/U8  ( .x(\net243[1] ), .a(wd[46]), .b(net263) );
    and2_1 \U76_15_/U8  ( .x(\net243[0] ), .a(wd[47]), .b(net263) );
    and2_1 \U80_0_/U8  ( .x(\net240[15] ), .a(wd[16]), .b(net267) );
    and2_1 \U80_1_/U8  ( .x(\net240[14] ), .a(wd[17]), .b(net267) );
    and2_1 \U80_2_/U8  ( .x(\net240[13] ), .a(wd[18]), .b(net267) );
    and2_1 \U80_3_/U8  ( .x(\net240[12] ), .a(wd[19]), .b(net267) );
    and2_1 \U80_4_/U8  ( .x(\net240[11] ), .a(wd[20]), .b(net267) );
    and2_1 \U80_5_/U8  ( .x(\net240[10] ), .a(wd[21]), .b(net267) );
    and2_1 \U80_6_/U8  ( .x(\net240[9] ), .a(wd[22]), .b(net267) );
    and2_1 \U80_7_/U8  ( .x(\net240[8] ), .a(wd[23]), .b(net267) );
    and2_1 \U80_8_/U8  ( .x(\net240[7] ), .a(wd[48]), .b(net267) );
    and2_1 \U80_9_/U8  ( .x(\net240[6] ), .a(wd[49]), .b(net267) );
    and2_1 \U80_10_/U8  ( .x(\net240[5] ), .a(wd[50]), .b(net267) );
    and2_1 \U80_11_/U8  ( .x(\net240[4] ), .a(wd[51]), .b(net267) );
    and2_1 \U80_12_/U8  ( .x(\net240[3] ), .a(wd[52]), .b(net267) );
    and2_1 \U80_13_/U8  ( .x(\net240[2] ), .a(wd[53]), .b(net267) );
    and2_1 \U80_14_/U8  ( .x(\net240[1] ), .a(wd[54]), .b(net267) );
    and2_1 \U80_15_/U8  ( .x(\net240[0] ), .a(wd[55]), .b(net267) );
    and2_1 \U128_0_/U8  ( .x(\net237[15] ), .a(seq[0]), .b(net269) );
    and2_1 \U128_1_/U8  ( .x(\net237[14] ), .a(pred[0]), .b(net269) );
    and2_1 \U128_2_/U8  ( .x(\net237[13] ), .a(lock[0]), .b(net269) );
    and2_1 \U128_3_/U8  ( .x(\net237[12] ), .a(\hdr[4] ), .b(net269) );
    and2_1 \U128_4_/U8  ( .x(\net237[11] ), .a(\hdr[4] ), .b(net269) );
    and2_1 \U128_5_/U8  ( .x(\net237[10] ), .a(rnw[0]), .b(net269) );
    and2_1 \U128_6_/U8  ( .x(\net237[9] ), .a(size[0]), .b(net269) );
    and2_1 \U128_7_/U8  ( .x(\net237[8] ), .a(size[1]), .b(net269) );
    and2_1 \U128_8_/U8  ( .x(\net237[7] ), .a(seq[1]), .b(net269) );
    and2_1 \U128_9_/U8  ( .x(\net237[6] ), .a(pred[1]), .b(net269) );
    and2_1 \U128_10_/U8  ( .x(\net237[5] ), .a(lock[1]), .b(net269) );
    and2_1 \U128_13_/U8  ( .x(\net237[2] ), .a(rnw[1]), .b(net269) );
    and2_1 \U128_14_/U8  ( .x(\net237[1] ), .a(size[2]), .b(net269) );
    and2_1 \U128_15_/U8  ( .x(\net237[0] ), .a(size[3]), .b(net269) );
    and2_1 \U37_0_/U8  ( .x(\net234[15] ), .a(addr[8]), .b(net259) );
    and2_1 \U37_1_/U8  ( .x(\net234[14] ), .a(addr[9]), .b(net259) );
    and2_1 \U37_2_/U8  ( .x(\net234[13] ), .a(addr[10]), .b(net259) );
    and2_1 \U37_3_/U8  ( .x(\net234[12] ), .a(addr[11]), .b(net259) );
    and2_1 \U37_4_/U8  ( .x(\net234[11] ), .a(addr[12]), .b(net259) );
    and2_1 \U37_5_/U8  ( .x(\net234[10] ), .a(addr[13]), .b(net259) );
    and2_1 \U37_6_/U8  ( .x(\net234[9] ), .a(addr[14]), .b(net259) );
    and2_1 \U37_7_/U8  ( .x(\net234[8] ), .a(addr[15]), .b(net259) );
    and2_1 \U37_8_/U8  ( .x(\net234[7] ), .a(addr[40]), .b(net259) );
    and2_1 \U37_9_/U8  ( .x(\net234[6] ), .a(addr[41]), .b(net259) );
    and2_1 \U37_10_/U8  ( .x(\net234[5] ), .a(addr[42]), .b(net259) );
    and2_1 \U37_11_/U8  ( .x(\net234[4] ), .a(addr[43]), .b(net259) );
    and2_1 \U37_12_/U8  ( .x(\net234[3] ), .a(addr[44]), .b(net259) );
    and2_1 \U37_13_/U8  ( .x(\net234[2] ), .a(addr[45]), .b(net259) );
    and2_1 \U37_14_/U8  ( .x(\net234[1] ), .a(addr[46]), .b(net259) );
    and2_1 \U37_15_/U8  ( .x(\net234[0] ), .a(addr[47]), .b(net259) );
    and2_1 \U33_0_/U8  ( .x(\net231[15] ), .a(addr[16]), .b(net253) );
    and2_1 \U33_1_/U8  ( .x(\net231[14] ), .a(addr[17]), .b(net253) );
    and2_1 \U33_2_/U8  ( .x(\net231[13] ), .a(addr[18]), .b(net253) );
    and2_1 \U33_3_/U8  ( .x(\net231[12] ), .a(addr[19]), .b(net253) );
    and2_1 \U33_4_/U8  ( .x(\net231[11] ), .a(addr[20]), .b(net253) );
    and2_1 \U33_5_/U8  ( .x(\net231[10] ), .a(addr[21]), .b(net253) );
    and2_1 \U33_6_/U8  ( .x(\net231[9] ), .a(addr[22]), .b(net253) );
    and2_1 \U33_7_/U8  ( .x(\net231[8] ), .a(addr[23]), .b(net253) );
    and2_1 \U33_8_/U8  ( .x(\net231[7] ), .a(addr[48]), .b(net253) );
    and2_1 \U33_9_/U8  ( .x(\net231[6] ), .a(addr[49]), .b(net253) );
    and2_1 \U33_10_/U8  ( .x(\net231[5] ), .a(addr[50]), .b(net253) );
    and2_1 \U33_11_/U8  ( .x(\net231[4] ), .a(addr[51]), .b(net253) );
    and2_1 \U33_12_/U8  ( .x(\net231[3] ), .a(addr[52]), .b(net253) );
    and2_1 \U33_13_/U8  ( .x(\net231[2] ), .a(addr[53]), .b(net253) );
    and2_1 \U33_14_/U8  ( .x(\net231[1] ), .a(addr[54]), .b(net253) );
    and2_1 \U33_15_/U8  ( .x(\net231[0] ), .a(addr[55]), .b(net253) );
    and2_1 \U81_0_/U8  ( .x(\net228[15] ), .a(wd[24]), .b(net255) );
    and2_1 \U81_1_/U8  ( .x(\net228[14] ), .a(wd[25]), .b(net255) );
    and2_1 \U81_2_/U8  ( .x(\net228[13] ), .a(wd[26]), .b(net255) );
    and2_1 \U81_3_/U8  ( .x(\net228[12] ), .a(wd[27]), .b(net255) );
    and2_1 \U81_4_/U8  ( .x(\net228[11] ), .a(wd[28]), .b(net255) );
    and2_1 \U81_5_/U8  ( .x(\net228[10] ), .a(wd[29]), .b(net255) );
    and2_1 \U81_6_/U8  ( .x(\net228[9] ), .a(wd[30]), .b(net255) );
    and2_1 \U81_7_/U8  ( .x(\net228[8] ), .a(wd[31]), .b(net255) );
    and2_1 \U81_8_/U8  ( .x(\net228[7] ), .a(wd[56]), .b(net255) );
    and2_1 \U81_9_/U8  ( .x(\net228[6] ), .a(wd[57]), .b(net255) );
    and2_1 \U81_10_/U8  ( .x(\net228[5] ), .a(wd[58]), .b(net255) );
    and2_1 \U81_11_/U8  ( .x(\net228[4] ), .a(wd[59]), .b(net255) );
    and2_1 \U81_12_/U8  ( .x(\net228[3] ), .a(wd[60]), .b(net255) );
    and2_1 \U81_13_/U8  ( .x(\net228[2] ), .a(wd[61]), .b(net255) );
    and2_1 \U81_14_/U8  ( .x(\net228[1] ), .a(wd[62]), .b(net255) );
    and2_1 \U81_15_/U8  ( .x(\net228[0] ), .a(wd[63]), .b(net255) );
    and2_1 \U34_0_/U8  ( .x(\net225[15] ), .a(addr[0]), .b(net251) );
    and2_1 \U34_1_/U8  ( .x(\net225[14] ), .a(addr[1]), .b(net251) );
    and2_1 \U34_2_/U8  ( .x(\net225[13] ), .a(addr[2]), .b(net251) );
    and2_1 \U34_3_/U8  ( .x(\net225[12] ), .a(addr[3]), .b(net251) );
    and2_1 \U34_4_/U8  ( .x(\net225[11] ), .a(addr[4]), .b(net251) );
    and2_1 \U34_5_/U8  ( .x(\net225[10] ), .a(addr[5]), .b(net251) );
    and2_1 \U34_6_/U8  ( .x(\net225[9] ), .a(addr[6]), .b(net251) );
    and2_1 \U34_7_/U8  ( .x(\net225[8] ), .a(addr[7]), .b(net251) );
    and2_1 \U34_8_/U8  ( .x(\net225[7] ), .a(addr[32]), .b(net251) );
    and2_1 \U34_9_/U8  ( .x(\net225[6] ), .a(addr[33]), .b(net251) );
    and2_1 \U34_10_/U8  ( .x(\net225[5] ), .a(addr[34]), .b(net251) );
    and2_1 \U34_11_/U8  ( .x(\net225[4] ), .a(addr[35]), .b(net251) );
    and2_1 \U34_12_/U8  ( .x(\net225[3] ), .a(addr[36]), .b(net251) );
    and2_1 \U34_13_/U8  ( .x(\net225[2] ), .a(addr[37]), .b(net251) );
    and2_1 \U34_14_/U8  ( .x(\net225[1] ), .a(addr[38]), .b(net251) );
    and2_1 \U34_15_/U8  ( .x(\net225[0] ), .a(addr[39]), .b(net251) );
    and2_1 \U30_0_/U8  ( .x(\net222[15] ), .a(addr[24]), .b(net261) );
    and2_1 \U30_1_/U8  ( .x(\net222[14] ), .a(addr[25]), .b(net261) );
    and2_1 \U30_2_/U8  ( .x(\net222[13] ), .a(addr[26]), .b(net261) );
    and2_1 \U30_3_/U8  ( .x(\net222[12] ), .a(addr[27]), .b(net261) );
    and2_1 \U30_4_/U8  ( .x(\net222[11] ), .a(addr[28]), .b(net261) );
    and2_1 \U30_5_/U8  ( .x(\net222[10] ), .a(addr[29]), .b(net261) );
    and2_1 \U30_6_/U8  ( .x(\net222[9] ), .a(addr[30]), .b(net261) );
    and2_1 \U30_7_/U8  ( .x(\net222[8] ), .a(addr[31]), .b(net261) );
    and2_1 \U30_8_/U8  ( .x(\net222[7] ), .a(addr[56]), .b(net261) );
    and2_1 \U30_9_/U8  ( .x(\net222[6] ), .a(addr[57]), .b(net261) );
    and2_1 \U30_10_/U8  ( .x(\net222[5] ), .a(addr[58]), .b(net261) );
    and2_1 \U30_11_/U8  ( .x(\net222[4] ), .a(addr[59]), .b(net261) );
    and2_1 \U30_12_/U8  ( .x(\net222[3] ), .a(addr[60]), .b(net261) );
    and2_1 \U30_13_/U8  ( .x(\net222[2] ), .a(addr[61]), .b(net261) );
    and2_1 \U30_14_/U8  ( .x(\net222[1] ), .a(addr[62]), .b(net261) );
    and2_1 \U30_15_/U8  ( .x(\net222[0] ), .a(addr[63]), .b(net261) );
    and2_1 \U82_0_/U8  ( .x(\net219[15] ), .a(wd[0]), .b(net249) );
    and2_1 \U82_1_/U8  ( .x(\net219[14] ), .a(wd[1]), .b(net249) );
    and2_1 \U82_2_/U8  ( .x(\net219[13] ), .a(wd[2]), .b(net249) );
    and2_1 \U82_3_/U8  ( .x(\net219[12] ), .a(wd[3]), .b(net249) );
    and2_1 \U82_4_/U8  ( .x(\net219[11] ), .a(wd[4]), .b(net249) );
    and2_1 \U82_5_/U8  ( .x(\net219[10] ), .a(wd[5]), .b(net249) );
    and2_1 \U82_6_/U8  ( .x(\net219[9] ), .a(wd[6]), .b(net249) );
    and2_1 \U82_7_/U8  ( .x(\net219[8] ), .a(wd[7]), .b(net249) );
    and2_1 \U82_8_/U8  ( .x(\net219[7] ), .a(wd[32]), .b(net249) );
    and2_1 \U82_9_/U8  ( .x(\net219[6] ), .a(wd[33]), .b(net249) );
    and2_1 \U82_10_/U8  ( .x(\net219[5] ), .a(wd[34]), .b(net249) );
    and2_1 \U82_11_/U8  ( .x(\net219[4] ), .a(wd[35]), .b(net249) );
    and2_1 \U82_12_/U8  ( .x(\net219[3] ), .a(wd[36]), .b(net249) );
    and2_1 \U82_13_/U8  ( .x(\net219[2] ), .a(wd[37]), .b(net249) );
    and2_1 \U82_14_/U8  ( .x(\net219[1] ), .a(wd[38]), .b(net249) );
    and2_1 \U82_15_/U8  ( .x(\net219[0] ), .a(wd[39]), .b(net249) );
    inv_1 \U40_0_/U3  ( .x(\U40_0_/n3 ), .a(\net225[15] ) );
    inv_1 \U40_0_/U4  ( .x(\U40_0_/n4 ), .a(\net234[15] ) );
    inv_1 \U40_0_/U5  ( .x(\net217[15] ), .a(\U40_0_/n5 ) );
    inv_1 \U40_1_/U3  ( .x(\U40_1_/n3 ), .a(\net225[14] ) );
    inv_1 \U40_1_/U4  ( .x(\U40_1_/n4 ), .a(\net234[14] ) );
    inv_1 \U40_1_/U5  ( .x(\net217[14] ), .a(\U40_1_/n5 ) );
    inv_1 \U40_2_/U3  ( .x(\U40_2_/n3 ), .a(\net225[13] ) );
    inv_1 \U40_2_/U4  ( .x(\U40_2_/n4 ), .a(\net234[13] ) );
    inv_1 \U40_2_/U5  ( .x(\net217[13] ), .a(\U40_2_/n5 ) );
    inv_1 \U40_3_/U3  ( .x(\U40_3_/n3 ), .a(\net225[12] ) );
    inv_1 \U40_3_/U4  ( .x(\U40_3_/n4 ), .a(\net234[12] ) );
    inv_1 \U40_3_/U5  ( .x(\net217[12] ), .a(\U40_3_/n5 ) );
    inv_1 \U40_4_/U3  ( .x(\U40_4_/n3 ), .a(\net225[11] ) );
    inv_1 \U40_4_/U4  ( .x(\U40_4_/n4 ), .a(\net234[11] ) );
    inv_1 \U40_4_/U5  ( .x(\net217[11] ), .a(\U40_4_/n5 ) );
    inv_1 \U40_5_/U3  ( .x(\U40_5_/n3 ), .a(\net225[10] ) );
    inv_1 \U40_5_/U4  ( .x(\U40_5_/n4 ), .a(\net234[10] ) );
    inv_1 \U40_5_/U5  ( .x(\net217[10] ), .a(\U40_5_/n5 ) );
    inv_1 \U40_6_/U3  ( .x(\U40_6_/n3 ), .a(\net225[9] ) );
    inv_1 \U40_6_/U4  ( .x(\U40_6_/n4 ), .a(\net234[9] ) );
    inv_1 \U40_6_/U5  ( .x(\net217[9] ), .a(\U40_6_/n5 ) );
    inv_1 \U40_7_/U3  ( .x(\U40_7_/n3 ), .a(\net225[8] ) );
    inv_1 \U40_7_/U4  ( .x(\U40_7_/n4 ), .a(\net234[8] ) );
    inv_1 \U40_7_/U5  ( .x(\net217[8] ), .a(\U40_7_/n5 ) );
    inv_1 \U40_8_/U3  ( .x(\U40_8_/n3 ), .a(\net225[7] ) );
    inv_1 \U40_8_/U4  ( .x(\U40_8_/n4 ), .a(\net234[7] ) );
    inv_1 \U40_8_/U5  ( .x(\net217[7] ), .a(\U40_8_/n5 ) );
    inv_1 \U40_9_/U3  ( .x(\U40_9_/n3 ), .a(\net225[6] ) );
    inv_1 \U40_9_/U4  ( .x(\U40_9_/n4 ), .a(\net234[6] ) );
    inv_1 \U40_9_/U5  ( .x(\net217[6] ), .a(\U40_9_/n5 ) );
    inv_1 \U40_10_/U3  ( .x(\U40_10_/n3 ), .a(\net225[5] ) );
    inv_1 \U40_10_/U4  ( .x(\U40_10_/n4 ), .a(\net234[5] ) );
    inv_1 \U40_10_/U5  ( .x(\net217[5] ), .a(\U40_10_/n5 ) );
    inv_1 \U40_11_/U3  ( .x(\U40_11_/n3 ), .a(\net225[4] ) );
    inv_1 \U40_11_/U4  ( .x(\U40_11_/n4 ), .a(\net234[4] ) );
    inv_1 \U40_11_/U5  ( .x(\net217[4] ), .a(\U40_11_/n5 ) );
    inv_1 \U40_12_/U3  ( .x(\U40_12_/n3 ), .a(\net225[3] ) );
    inv_1 \U40_12_/U4  ( .x(\U40_12_/n4 ), .a(\net234[3] ) );
    inv_1 \U40_12_/U5  ( .x(\net217[3] ), .a(\U40_12_/n5 ) );
    inv_1 \U40_13_/U3  ( .x(\U40_13_/n3 ), .a(\net225[2] ) );
    inv_1 \U40_13_/U4  ( .x(\U40_13_/n4 ), .a(\net234[2] ) );
    inv_1 \U40_13_/U5  ( .x(\net217[2] ), .a(\U40_13_/n5 ) );
    inv_1 \U40_14_/U3  ( .x(\U40_14_/n3 ), .a(\net225[1] ) );
    inv_1 \U40_14_/U4  ( .x(\U40_14_/n4 ), .a(\net234[1] ) );
    inv_1 \U40_14_/U5  ( .x(\net217[1] ), .a(\U40_14_/n5 ) );
    inv_1 \U40_15_/U3  ( .x(\U40_15_/n3 ), .a(\net225[0] ) );
    inv_1 \U40_15_/U4  ( .x(\U40_15_/n4 ), .a(\net234[0] ) );
    inv_1 \U40_15_/U5  ( .x(\net217[0] ), .a(\U40_15_/n5 ) );
    and4_1 \U14_0_/U16  ( .x(\U14_0_/n5 ), .a(\U14_0_/n1 ), .b(\U14_0_/n2 ), 
        .c(\U14_0_/n3 ), .d(\U14_0_/n4 ) );
    inv_1 \U14_0_/U1  ( .x(\U14_0_/n1 ), .a(\net231[15] ) );
    inv_1 \U14_0_/U2  ( .x(\U14_0_/n2 ), .a(\net222[15] ) );
    inv_1 \U14_0_/U3  ( .x(\U14_0_/n3 ), .a(\net237[15] ) );
    inv_1 \U14_0_/U4  ( .x(\U14_0_/n4 ), .a(\net246[15] ) );
    inv_1 \U14_0_/U5  ( .x(\net212[15] ), .a(\U14_0_/n5 ) );
    and4_1 \U14_1_/U16  ( .x(\U14_1_/n5 ), .a(\U14_1_/n1 ), .b(\U14_1_/n2 ), 
        .c(\U14_1_/n3 ), .d(\U14_1_/n4 ) );
    inv_1 \U14_1_/U1  ( .x(\U14_1_/n1 ), .a(\net231[14] ) );
    inv_1 \U14_1_/U2  ( .x(\U14_1_/n2 ), .a(\net222[14] ) );
    inv_1 \U14_1_/U3  ( .x(\U14_1_/n3 ), .a(\net237[14] ) );
    inv_1 \U14_1_/U4  ( .x(\U14_1_/n4 ), .a(\net246[14] ) );
    inv_1 \U14_1_/U5  ( .x(\net212[14] ), .a(\U14_1_/n5 ) );
    and4_1 \U14_2_/U16  ( .x(\U14_2_/n5 ), .a(\U14_2_/n1 ), .b(\U14_2_/n2 ), 
        .c(\U14_2_/n3 ), .d(\U14_2_/n4 ) );
    inv_1 \U14_2_/U1  ( .x(\U14_2_/n1 ), .a(\net231[13] ) );
    inv_1 \U14_2_/U2  ( .x(\U14_2_/n2 ), .a(\net222[13] ) );
    inv_1 \U14_2_/U3  ( .x(\U14_2_/n3 ), .a(\net237[13] ) );
    inv_1 \U14_2_/U4  ( .x(\U14_2_/n4 ), .a(\net246[13] ) );
    inv_1 \U14_2_/U5  ( .x(\net212[13] ), .a(\U14_2_/n5 ) );
    and4_1 \U14_3_/U16  ( .x(\U14_3_/n5 ), .a(\U14_3_/n1 ), .b(\U14_3_/n2 ), 
        .c(\U14_3_/n3 ), .d(\U14_3_/n4 ) );
    inv_1 \U14_3_/U1  ( .x(\U14_3_/n1 ), .a(\net231[12] ) );
    inv_1 \U14_3_/U2  ( .x(\U14_3_/n2 ), .a(\net222[12] ) );
    inv_1 \U14_3_/U3  ( .x(\U14_3_/n3 ), .a(\net237[12] ) );
    inv_1 \U14_3_/U4  ( .x(\U14_3_/n4 ), .a(\net246[12] ) );
    inv_1 \U14_3_/U5  ( .x(\net212[12] ), .a(\U14_3_/n5 ) );
    and4_1 \U14_4_/U16  ( .x(\U14_4_/n5 ), .a(\U14_4_/n1 ), .b(\U14_4_/n2 ), 
        .c(\U14_4_/n3 ), .d(\U14_4_/n4 ) );
    inv_1 \U14_4_/U1  ( .x(\U14_4_/n1 ), .a(\net231[11] ) );
    inv_1 \U14_4_/U2  ( .x(\U14_4_/n2 ), .a(\net222[11] ) );
    inv_1 \U14_4_/U3  ( .x(\U14_4_/n3 ), .a(\net237[11] ) );
    inv_1 \U14_4_/U4  ( .x(\U14_4_/n4 ), .a(\net246[11] ) );
    inv_1 \U14_4_/U5  ( .x(\net212[11] ), .a(\U14_4_/n5 ) );
    and4_1 \U14_5_/U16  ( .x(\U14_5_/n5 ), .a(\U14_5_/n1 ), .b(\U14_5_/n2 ), 
        .c(\U14_5_/n3 ), .d(\U14_5_/n4 ) );
    inv_1 \U14_5_/U1  ( .x(\U14_5_/n1 ), .a(\net231[10] ) );
    inv_1 \U14_5_/U2  ( .x(\U14_5_/n2 ), .a(\net222[10] ) );
    inv_1 \U14_5_/U3  ( .x(\U14_5_/n3 ), .a(\net237[10] ) );
    inv_1 \U14_5_/U4  ( .x(\U14_5_/n4 ), .a(\net246[10] ) );
    inv_1 \U14_5_/U5  ( .x(\net212[10] ), .a(\U14_5_/n5 ) );
    and4_1 \U14_6_/U16  ( .x(\U14_6_/n5 ), .a(\U14_6_/n1 ), .b(\U14_6_/n2 ), 
        .c(\U14_6_/n3 ), .d(\U14_6_/n4 ) );
    inv_1 \U14_6_/U1  ( .x(\U14_6_/n1 ), .a(\net231[9] ) );
    inv_1 \U14_6_/U2  ( .x(\U14_6_/n2 ), .a(\net222[9] ) );
    inv_1 \U14_6_/U3  ( .x(\U14_6_/n3 ), .a(\net237[9] ) );
    inv_1 \U14_6_/U4  ( .x(\U14_6_/n4 ), .a(\net246[9] ) );
    inv_1 \U14_6_/U5  ( .x(\net212[9] ), .a(\U14_6_/n5 ) );
    and4_1 \U14_7_/U16  ( .x(\U14_7_/n5 ), .a(\U14_7_/n1 ), .b(\U14_7_/n2 ), 
        .c(\U14_7_/n3 ), .d(\U14_7_/n4 ) );
    inv_1 \U14_7_/U1  ( .x(\U14_7_/n1 ), .a(\net231[8] ) );
    inv_1 \U14_7_/U2  ( .x(\U14_7_/n2 ), .a(\net222[8] ) );
    inv_1 \U14_7_/U3  ( .x(\U14_7_/n3 ), .a(\net237[8] ) );
    inv_1 \U14_7_/U4  ( .x(\U14_7_/n4 ), .a(\net246[8] ) );
    inv_1 \U14_7_/U5  ( .x(\net212[8] ), .a(\U14_7_/n5 ) );
    and4_1 \U14_8_/U16  ( .x(\U14_8_/n5 ), .a(\U14_8_/n1 ), .b(\U14_8_/n2 ), 
        .c(\U14_8_/n3 ), .d(\U14_8_/n4 ) );
    inv_1 \U14_8_/U1  ( .x(\U14_8_/n1 ), .a(\net231[7] ) );
    inv_1 \U14_8_/U2  ( .x(\U14_8_/n2 ), .a(\net222[7] ) );
    inv_1 \U14_8_/U3  ( .x(\U14_8_/n3 ), .a(\net237[7] ) );
    inv_1 \U14_8_/U4  ( .x(\U14_8_/n4 ), .a(\net246[7] ) );
    inv_1 \U14_8_/U5  ( .x(\net212[7] ), .a(\U14_8_/n5 ) );
    and4_1 \U14_9_/U16  ( .x(\U14_9_/n5 ), .a(\U14_9_/n1 ), .b(\U14_9_/n2 ), 
        .c(\U14_9_/n3 ), .d(\U14_9_/n4 ) );
    inv_1 \U14_9_/U1  ( .x(\U14_9_/n1 ), .a(\net231[6] ) );
    inv_1 \U14_9_/U2  ( .x(\U14_9_/n2 ), .a(\net222[6] ) );
    inv_1 \U14_9_/U3  ( .x(\U14_9_/n3 ), .a(\net237[6] ) );
    inv_1 \U14_9_/U4  ( .x(\U14_9_/n4 ), .a(\net246[6] ) );
    inv_1 \U14_9_/U5  ( .x(\net212[6] ), .a(\U14_9_/n5 ) );
    and4_1 \U14_10_/U16  ( .x(\U14_10_/n5 ), .a(\U14_10_/n1 ), .b(\U14_10_/n2 
        ), .c(\U14_10_/n3 ), .d(\U14_10_/n4 ) );
    inv_1 \U14_10_/U1  ( .x(\U14_10_/n1 ), .a(\net231[5] ) );
    inv_1 \U14_10_/U2  ( .x(\U14_10_/n2 ), .a(\net222[5] ) );
    inv_1 \U14_10_/U3  ( .x(\U14_10_/n3 ), .a(\net237[5] ) );
    inv_1 \U14_10_/U4  ( .x(\U14_10_/n4 ), .a(\net246[5] ) );
    inv_1 \U14_10_/U5  ( .x(\net212[5] ), .a(\U14_10_/n5 ) );
    inv_1 \U14_11_/U1  ( .x(\U14_11_/n1 ), .a(\net231[4] ) );
    inv_1 \U14_11_/U2  ( .x(\U14_11_/n2 ), .a(\net222[4] ) );
    inv_1 \U14_11_/U4  ( .x(\U14_11_/n4 ), .a(\net246[4] ) );
    inv_1 \U14_11_/U5  ( .x(\net212[4] ), .a(\U14_11_/n5 ) );
    inv_1 \U14_12_/U1  ( .x(\U14_12_/n1 ), .a(\net231[3] ) );
    inv_1 \U14_12_/U2  ( .x(\U14_12_/n2 ), .a(\net222[3] ) );
    inv_1 \U14_12_/U4  ( .x(\U14_12_/n4 ), .a(\net246[3] ) );
    inv_1 \U14_12_/U5  ( .x(\net212[3] ), .a(\U14_12_/n5 ) );
    and4_1 \U14_13_/U16  ( .x(\U14_13_/n5 ), .a(\U14_13_/n1 ), .b(\U14_13_/n2 
        ), .c(\U14_13_/n3 ), .d(\U14_13_/n4 ) );
    inv_1 \U14_13_/U1  ( .x(\U14_13_/n1 ), .a(\net231[2] ) );
    inv_1 \U14_13_/U2  ( .x(\U14_13_/n2 ), .a(\net222[2] ) );
    inv_1 \U14_13_/U3  ( .x(\U14_13_/n3 ), .a(\net237[2] ) );
    inv_1 \U14_13_/U4  ( .x(\U14_13_/n4 ), .a(\net246[2] ) );
    inv_1 \U14_13_/U5  ( .x(\net212[2] ), .a(\U14_13_/n5 ) );
    and4_1 \U14_14_/U16  ( .x(\U14_14_/n5 ), .a(\U14_14_/n1 ), .b(\U14_14_/n2 
        ), .c(\U14_14_/n3 ), .d(\U14_14_/n4 ) );
    inv_1 \U14_14_/U1  ( .x(\U14_14_/n1 ), .a(\net231[1] ) );
    inv_1 \U14_14_/U2  ( .x(\U14_14_/n2 ), .a(\net222[1] ) );
    inv_1 \U14_14_/U3  ( .x(\U14_14_/n3 ), .a(\net237[1] ) );
    inv_1 \U14_14_/U4  ( .x(\U14_14_/n4 ), .a(\net246[1] ) );
    inv_1 \U14_14_/U5  ( .x(\net212[1] ), .a(\U14_14_/n5 ) );
    and4_1 \U14_15_/U16  ( .x(\U14_15_/n5 ), .a(\U14_15_/n1 ), .b(\U14_15_/n2 
        ), .c(\U14_15_/n3 ), .d(\U14_15_/n4 ) );
    inv_1 \U14_15_/U1  ( .x(\U14_15_/n1 ), .a(\net231[0] ) );
    inv_1 \U14_15_/U2  ( .x(\U14_15_/n2 ), .a(\net222[0] ) );
    inv_1 \U14_15_/U3  ( .x(\U14_15_/n3 ), .a(\net237[0] ) );
    inv_1 \U14_15_/U4  ( .x(\U14_15_/n4 ), .a(\net246[0] ) );
    inv_1 \U14_15_/U5  ( .x(\net212[0] ), .a(\U14_15_/n5 ) );
    and4_1 \U91_0_/U16  ( .x(\U91_0_/n5 ), .a(\U91_0_/n1 ), .b(\U91_0_/n2 ), 
        .c(\U91_0_/n3 ), .d(\U91_0_/n4 ) );
    inv_1 \U91_0_/U1  ( .x(\U91_0_/n1 ), .a(\net219[15] ) );
    inv_1 \U91_0_/U2  ( .x(\U91_0_/n2 ), .a(\net243[15] ) );
    inv_1 \U91_0_/U3  ( .x(\U91_0_/n3 ), .a(\net240[15] ) );
    inv_1 \U91_0_/U4  ( .x(\U91_0_/n4 ), .a(\net228[15] ) );
    inv_1 \U91_0_/U5  ( .x(\net207[15] ), .a(\U91_0_/n5 ) );
    and4_1 \U91_1_/U16  ( .x(\U91_1_/n5 ), .a(\U91_1_/n1 ), .b(\U91_1_/n2 ), 
        .c(\U91_1_/n3 ), .d(\U91_1_/n4 ) );
    inv_1 \U91_1_/U1  ( .x(\U91_1_/n1 ), .a(\net219[14] ) );
    inv_1 \U91_1_/U2  ( .x(\U91_1_/n2 ), .a(\net243[14] ) );
    inv_1 \U91_1_/U3  ( .x(\U91_1_/n3 ), .a(\net240[14] ) );
    inv_1 \U91_1_/U4  ( .x(\U91_1_/n4 ), .a(\net228[14] ) );
    inv_1 \U91_1_/U5  ( .x(\net207[14] ), .a(\U91_1_/n5 ) );
    and4_1 \U91_2_/U16  ( .x(\U91_2_/n5 ), .a(\U91_2_/n1 ), .b(\U91_2_/n2 ), 
        .c(\U91_2_/n3 ), .d(\U91_2_/n4 ) );
    inv_1 \U91_2_/U1  ( .x(\U91_2_/n1 ), .a(\net219[13] ) );
    inv_1 \U91_2_/U2  ( .x(\U91_2_/n2 ), .a(\net243[13] ) );
    inv_1 \U91_2_/U3  ( .x(\U91_2_/n3 ), .a(\net240[13] ) );
    inv_1 \U91_2_/U4  ( .x(\U91_2_/n4 ), .a(\net228[13] ) );
    inv_1 \U91_2_/U5  ( .x(\net207[13] ), .a(\U91_2_/n5 ) );
    and4_1 \U91_3_/U16  ( .x(\U91_3_/n5 ), .a(\U91_3_/n1 ), .b(\U91_3_/n2 ), 
        .c(\U91_3_/n3 ), .d(\U91_3_/n4 ) );
    inv_1 \U91_3_/U1  ( .x(\U91_3_/n1 ), .a(\net219[12] ) );
    inv_1 \U91_3_/U2  ( .x(\U91_3_/n2 ), .a(\net243[12] ) );
    inv_1 \U91_3_/U3  ( .x(\U91_3_/n3 ), .a(\net240[12] ) );
    inv_1 \U91_3_/U4  ( .x(\U91_3_/n4 ), .a(\net228[12] ) );
    inv_1 \U91_3_/U5  ( .x(\net207[12] ), .a(\U91_3_/n5 ) );
    and4_1 \U91_4_/U16  ( .x(\U91_4_/n5 ), .a(\U91_4_/n1 ), .b(\U91_4_/n2 ), 
        .c(\U91_4_/n3 ), .d(\U91_4_/n4 ) );
    inv_1 \U91_4_/U1  ( .x(\U91_4_/n1 ), .a(\net219[11] ) );
    inv_1 \U91_4_/U2  ( .x(\U91_4_/n2 ), .a(\net243[11] ) );
    inv_1 \U91_4_/U3  ( .x(\U91_4_/n3 ), .a(\net240[11] ) );
    inv_1 \U91_4_/U4  ( .x(\U91_4_/n4 ), .a(\net228[11] ) );
    inv_1 \U91_4_/U5  ( .x(\net207[11] ), .a(\U91_4_/n5 ) );
    and4_1 \U91_5_/U16  ( .x(\U91_5_/n5 ), .a(\U91_5_/n1 ), .b(\U91_5_/n2 ), 
        .c(\U91_5_/n3 ), .d(\U91_5_/n4 ) );
    inv_1 \U91_5_/U1  ( .x(\U91_5_/n1 ), .a(\net219[10] ) );
    inv_1 \U91_5_/U2  ( .x(\U91_5_/n2 ), .a(\net243[10] ) );
    inv_1 \U91_5_/U3  ( .x(\U91_5_/n3 ), .a(\net240[10] ) );
    inv_1 \U91_5_/U4  ( .x(\U91_5_/n4 ), .a(\net228[10] ) );
    inv_1 \U91_5_/U5  ( .x(\net207[10] ), .a(\U91_5_/n5 ) );
    and4_1 \U91_6_/U16  ( .x(\U91_6_/n5 ), .a(\U91_6_/n1 ), .b(\U91_6_/n2 ), 
        .c(\U91_6_/n3 ), .d(\U91_6_/n4 ) );
    inv_1 \U91_6_/U1  ( .x(\U91_6_/n1 ), .a(\net219[9] ) );
    inv_1 \U91_6_/U2  ( .x(\U91_6_/n2 ), .a(\net243[9] ) );
    inv_1 \U91_6_/U3  ( .x(\U91_6_/n3 ), .a(\net240[9] ) );
    inv_1 \U91_6_/U4  ( .x(\U91_6_/n4 ), .a(\net228[9] ) );
    inv_1 \U91_6_/U5  ( .x(\net207[9] ), .a(\U91_6_/n5 ) );
    and4_1 \U91_7_/U16  ( .x(\U91_7_/n5 ), .a(\U91_7_/n1 ), .b(\U91_7_/n2 ), 
        .c(\U91_7_/n3 ), .d(\U91_7_/n4 ) );
    inv_1 \U91_7_/U1  ( .x(\U91_7_/n1 ), .a(\net219[8] ) );
    inv_1 \U91_7_/U2  ( .x(\U91_7_/n2 ), .a(\net243[8] ) );
    inv_1 \U91_7_/U3  ( .x(\U91_7_/n3 ), .a(\net240[8] ) );
    inv_1 \U91_7_/U4  ( .x(\U91_7_/n4 ), .a(\net228[8] ) );
    inv_1 \U91_7_/U5  ( .x(\net207[8] ), .a(\U91_7_/n5 ) );
    and4_1 \U91_8_/U16  ( .x(\U91_8_/n5 ), .a(\U91_8_/n1 ), .b(\U91_8_/n2 ), 
        .c(\U91_8_/n3 ), .d(\U91_8_/n4 ) );
    inv_1 \U91_8_/U1  ( .x(\U91_8_/n1 ), .a(\net219[7] ) );
    inv_1 \U91_8_/U2  ( .x(\U91_8_/n2 ), .a(\net243[7] ) );
    inv_1 \U91_8_/U3  ( .x(\U91_8_/n3 ), .a(\net240[7] ) );
    inv_1 \U91_8_/U4  ( .x(\U91_8_/n4 ), .a(\net228[7] ) );
    inv_1 \U91_8_/U5  ( .x(\net207[7] ), .a(\U91_8_/n5 ) );
    and4_1 \U91_9_/U16  ( .x(\U91_9_/n5 ), .a(\U91_9_/n1 ), .b(\U91_9_/n2 ), 
        .c(\U91_9_/n3 ), .d(\U91_9_/n4 ) );
    inv_1 \U91_9_/U1  ( .x(\U91_9_/n1 ), .a(\net219[6] ) );
    inv_1 \U91_9_/U2  ( .x(\U91_9_/n2 ), .a(\net243[6] ) );
    inv_1 \U91_9_/U3  ( .x(\U91_9_/n3 ), .a(\net240[6] ) );
    inv_1 \U91_9_/U4  ( .x(\U91_9_/n4 ), .a(\net228[6] ) );
    inv_1 \U91_9_/U5  ( .x(\net207[6] ), .a(\U91_9_/n5 ) );
    and4_1 \U91_10_/U16  ( .x(\U91_10_/n5 ), .a(\U91_10_/n1 ), .b(\U91_10_/n2 
        ), .c(\U91_10_/n3 ), .d(\U91_10_/n4 ) );
    inv_1 \U91_10_/U1  ( .x(\U91_10_/n1 ), .a(\net219[5] ) );
    inv_1 \U91_10_/U2  ( .x(\U91_10_/n2 ), .a(\net243[5] ) );
    inv_1 \U91_10_/U3  ( .x(\U91_10_/n3 ), .a(\net240[5] ) );
    inv_1 \U91_10_/U4  ( .x(\U91_10_/n4 ), .a(\net228[5] ) );
    inv_1 \U91_10_/U5  ( .x(\net207[5] ), .a(\U91_10_/n5 ) );
    and4_1 \U91_11_/U16  ( .x(\U91_11_/n5 ), .a(\U91_11_/n1 ), .b(\U91_11_/n2 
        ), .c(\U91_11_/n3 ), .d(\U91_11_/n4 ) );
    inv_1 \U91_11_/U1  ( .x(\U91_11_/n1 ), .a(\net219[4] ) );
    inv_1 \U91_11_/U2  ( .x(\U91_11_/n2 ), .a(\net243[4] ) );
    inv_1 \U91_11_/U3  ( .x(\U91_11_/n3 ), .a(\net240[4] ) );
    inv_1 \U91_11_/U4  ( .x(\U91_11_/n4 ), .a(\net228[4] ) );
    inv_1 \U91_11_/U5  ( .x(\net207[4] ), .a(\U91_11_/n5 ) );
    and4_1 \U91_12_/U16  ( .x(\U91_12_/n5 ), .a(\U91_12_/n1 ), .b(\U91_12_/n2 
        ), .c(\U91_12_/n3 ), .d(\U91_12_/n4 ) );
    inv_1 \U91_12_/U1  ( .x(\U91_12_/n1 ), .a(\net219[3] ) );
    inv_1 \U91_12_/U2  ( .x(\U91_12_/n2 ), .a(\net243[3] ) );
    inv_1 \U91_12_/U3  ( .x(\U91_12_/n3 ), .a(\net240[3] ) );
    inv_1 \U91_12_/U4  ( .x(\U91_12_/n4 ), .a(\net228[3] ) );
    inv_1 \U91_12_/U5  ( .x(\net207[3] ), .a(\U91_12_/n5 ) );
    and4_1 \U91_13_/U16  ( .x(\U91_13_/n5 ), .a(\U91_13_/n1 ), .b(\U91_13_/n2 
        ), .c(\U91_13_/n3 ), .d(\U91_13_/n4 ) );
    inv_1 \U91_13_/U1  ( .x(\U91_13_/n1 ), .a(\net219[2] ) );
    inv_1 \U91_13_/U2  ( .x(\U91_13_/n2 ), .a(\net243[2] ) );
    inv_1 \U91_13_/U3  ( .x(\U91_13_/n3 ), .a(\net240[2] ) );
    inv_1 \U91_13_/U4  ( .x(\U91_13_/n4 ), .a(\net228[2] ) );
    inv_1 \U91_13_/U5  ( .x(\net207[2] ), .a(\U91_13_/n5 ) );
    and4_1 \U91_14_/U16  ( .x(\U91_14_/n5 ), .a(\U91_14_/n1 ), .b(\U91_14_/n2 
        ), .c(\U91_14_/n3 ), .d(\U91_14_/n4 ) );
    inv_1 \U91_14_/U1  ( .x(\U91_14_/n1 ), .a(\net219[1] ) );
    inv_1 \U91_14_/U2  ( .x(\U91_14_/n2 ), .a(\net243[1] ) );
    inv_1 \U91_14_/U3  ( .x(\U91_14_/n3 ), .a(\net240[1] ) );
    inv_1 \U91_14_/U4  ( .x(\U91_14_/n4 ), .a(\net228[1] ) );
    inv_1 \U91_14_/U5  ( .x(\net207[1] ), .a(\U91_14_/n5 ) );
    and4_1 \U91_15_/U16  ( .x(\U91_15_/n5 ), .a(\U91_15_/n1 ), .b(\U91_15_/n2 
        ), .c(\U91_15_/n3 ), .d(\U91_15_/n4 ) );
    inv_1 \U91_15_/U1  ( .x(\U91_15_/n1 ), .a(\net219[0] ) );
    inv_1 \U91_15_/U2  ( .x(\U91_15_/n2 ), .a(\net243[0] ) );
    inv_1 \U91_15_/U3  ( .x(\U91_15_/n3 ), .a(\net240[0] ) );
    inv_1 \U91_15_/U4  ( .x(\U91_15_/n4 ), .a(\net228[0] ) );
    inv_1 \U91_15_/U5  ( .x(\net207[0] ), .a(\U91_15_/n5 ) );
    or3_2 \U93_0_/U12  ( .x(chainl[0]), .a(\net207[15] ), .b(\net217[15] ), 
        .c(\net212[15] ) );
    or3_2 \U93_1_/U12  ( .x(chainl[1]), .a(\net207[14] ), .b(\net217[14] ), 
        .c(\net212[14] ) );
    or3_2 \U93_2_/U12  ( .x(chainl[2]), .a(\net207[13] ), .b(\net217[13] ), 
        .c(\net212[13] ) );
    or3_2 \U93_3_/U12  ( .x(chainl[3]), .a(\net207[12] ), .b(\net217[12] ), 
        .c(\net212[12] ) );
    or3_2 \U93_4_/U12  ( .x(chainl[4]), .a(\net207[11] ), .b(\net217[11] ), 
        .c(\net212[11] ) );
    or3_2 \U93_5_/U12  ( .x(chainl[5]), .a(\net207[10] ), .b(\net217[10] ), 
        .c(\net212[10] ) );
    or3_2 \U93_6_/U12  ( .x(chainl[6]), .a(\net207[9] ), .b(\net217[9] ), .c(
        \net212[9] ) );
    or3_2 \U93_7_/U12  ( .x(chainl[7]), .a(\net207[8] ), .b(\net217[8] ), .c(
        \net212[8] ) );
    or3_2 \U93_8_/U12  ( .x(chainh[0]), .a(\net207[7] ), .b(\net217[7] ), .c(
        \net212[7] ) );
    or3_2 \U93_9_/U12  ( .x(chainh[1]), .a(\net207[6] ), .b(\net217[6] ), .c(
        \net212[6] ) );
    or3_2 \U93_10_/U12  ( .x(chainh[2]), .a(\net207[5] ), .b(\net217[5] ), .c(
        \net212[5] ) );
    or3_2 \U93_11_/U12  ( .x(chainh[3]), .a(\net207[4] ), .b(\net217[4] ), .c(
        \net212[4] ) );
    or3_2 \U93_12_/U12  ( .x(chainh[4]), .a(\net207[3] ), .b(\net217[3] ), .c(
        \net212[3] ) );
    or3_2 \U93_13_/U12  ( .x(chainh[5]), .a(\net207[2] ), .b(\net217[2] ), .c(
        \net212[2] ) );
    or3_2 \U93_14_/U12  ( .x(chainh[6]), .a(\net207[1] ), .b(\net217[1] ), .c(
        \net212[1] ) );
    or3_2 \U93_15_/U12  ( .x(chainh[7]), .a(\net207[0] ), .b(\net217[0] ), .c(
        \net212[0] ) );
    inv_1 \U152/U3  ( .x(net198), .a(sendreq) );
    ao23_1 \U158/U19/U21/U1/U1  ( .x(net131), .a(net132), .b(net131), .c(
        net132), .d(rnw[1]), .e(rnw[1]) );
    ao23_1 \U157/U19/U21/U1/U1  ( .x(net176), .a(net132), .b(net176), .c(
        net132), .d(rnw[0]), .e(rnw[0]) );
    ao222_1 \U123/U18/U1/U1  ( .x(net136), .a(net185), .b(net187), .c(net185), 
        .d(net136), .e(net187), .f(net136) );
    aoi21_1 \U151/U30/U1/U1  ( .x(\hdr[4] ), .a(\U151/Z ), .b(net138), .c(
        net198) );
    inv_1 \U151/U30/U1/U2  ( .x(\U151/Z ), .a(\hdr[4] ) );
    nor3_1 \U148/U21/Unr  ( .x(\U148/U21/nr ), .a(net191), .b(net136), .c(
        net293) );
    nand3_1 \U148/U21/Und  ( .x(\U148/U21/nd ), .a(net191), .b(net136), .c(
        net293) );
    oa21_1 \U148/U21/U1  ( .x(\U148/U21/n2 ), .a(\U148/U21/n2 ), .b(
        \U148/U21/nr ), .c(\U148/U21/nd ) );
    inv_1 \U148/U21/U3  ( .x(ack), .a(\U148/U21/n2 ) );
    buf_3 U1 ( .x(n1), .a(net138) );
    buf_3 U2 ( .x(net138), .a(nia) );
    buf_3 U3 ( .x(net269), .a(net146) );
    buf_3 U4 ( .x(net255), .a(\bs[5] ) );
    buf_3 U5 ( .x(net253), .a(\bs[2] ) );
    buf_3 U6 ( .x(net267), .a(\bs[6] ) );
    buf_3 U7 ( .x(net263), .a(\bs[7] ) );
    buf_3 U8 ( .x(net249), .a(\bs[8] ) );
    buf_3 U9 ( .x(net251), .a(\bs[4] ) );
    buf_3 U10 ( .x(net265), .a(\bs[0] ) );
    buf_3 U11 ( .x(net261), .a(\bs[1] ) );
    buf_3 U12 ( .x(net259), .a(\bs[3] ) );
    and2_1 U13 ( .x(\U40_2_/n5 ), .a(\U40_2_/n3 ), .b(\U40_2_/n4 ) );
    and2_1 U14 ( .x(\U40_1_/n5 ), .a(\U40_1_/n3 ), .b(\U40_1_/n4 ) );
    and2_1 U15 ( .x(\U40_9_/n5 ), .a(\U40_9_/n3 ), .b(\U40_9_/n4 ) );
    and2_1 U16 ( .x(\U40_8_/n5 ), .a(\U40_8_/n3 ), .b(\U40_8_/n4 ) );
    and2_1 U17 ( .x(\U40_13_/n5 ), .a(\U40_13_/n3 ), .b(\U40_13_/n4 ) );
    and2_1 U18 ( .x(\U40_0_/n5 ), .a(\U40_0_/n3 ), .b(\U40_0_/n4 ) );
    and2_1 U19 ( .x(\U40_5_/n5 ), .a(\U40_5_/n3 ), .b(\U40_5_/n4 ) );
    and2_1 U20 ( .x(\U40_4_/n5 ), .a(\U40_4_/n3 ), .b(\U40_4_/n4 ) );
    and3_1 U21 ( .x(\U14_12_/n5 ), .a(\U14_12_/n2 ), .b(\U14_12_/n4 ), .c(
        \U14_12_/n1 ) );
    and2_1 U22 ( .x(\U40_12_/n5 ), .a(\U40_12_/n3 ), .b(\U40_12_/n4 ) );
    and2_1 U23 ( .x(\U40_3_/n5 ), .a(\U40_3_/n3 ), .b(\U40_3_/n4 ) );
    and3_1 U24 ( .x(\U14_11_/n5 ), .a(\U14_11_/n2 ), .b(\U14_11_/n4 ), .c(
        \U14_11_/n1 ) );
    and2_1 U25 ( .x(\U40_11_/n5 ), .a(\U40_11_/n3 ), .b(\U40_11_/n4 ) );
    and2_1 U26 ( .x(\U40_10_/n5 ), .a(\U40_10_/n3 ), .b(\U40_10_/n4 ) );
    and2_1 U27 ( .x(\U40_15_/n5 ), .a(\U40_15_/n3 ), .b(\U40_15_/n4 ) );
    and2_1 U28 ( .x(\U40_7_/n5 ), .a(\U40_7_/n3 ), .b(\U40_7_/n4 ) );
    and2_1 U29 ( .x(\U40_6_/n5 ), .a(\U40_6_/n3 ), .b(\U40_6_/n4 ) );
    and2_1 U30 ( .x(\U40_14_/n5 ), .a(\U40_14_/n3 ), .b(\U40_14_/n4 ) );
endmodule


module chain_dr2fr_byte_0 ( eop_ack, ia, o, eop, ih, il, nReset, noa );
output [4:0] o;
input  [7:0] ih;
input  [7:0] il;
input  eop, nReset, noa;
output eop_ack, ia;
    wire eop_ack_wire, nbReset, eop_pass, nxa, naa, nlowack, \twobitack[0] , 
        \twobitack[1] , nhighack, \twobitack[2] , \twobitack[3] , \U1018/Z , 
        \U1270/net189 , \U1270/net192 , \U1270/net191 , net199, \U1270/net190 , 
        \U1270/U1141/Z , \U1268/net189 , \U1268/net192 , \U1268/net191 , 
        net194, \U1268/net190 , \U1268/U1141/Z , \U1224/nack[0] , \x[3] , 
        \x[2] , \U1224/nack[1] , \x[1] , \U1224/net4 , \x[0] , 
        \U1224/U1125/U28/U1/clr , asel, \U1224/U1125/U28/U1/set , 
        \U1224/U1122/U28/U1/clr , csel, nca, \U1224/U1122/U28/U1/set , 
        \U1224/U916_0_/U25/U1/clr , \a[0] , \c[0] , \U1224/U916_0_/U25/U1/ob , 
        \U1224/U916_1_/U25/U1/clr , \a[1] , \c[1] , \U1224/U916_1_/U25/U1/ob , 
        \U1224/U916_2_/U25/U1/clr , \a[2] , \c[2] , \U1224/U916_2_/U25/U1/ob , 
        \U1224/U916_3_/U25/U1/clr , \a[3] , \c[3] , \U1224/U916_3_/U25/U1/ob , 
        \U1209/nack[0] , \U1209/nack[1] , \U1209/net4 , 
        \U1209/U1125/U28/U1/clr , xsel, \U1209/U1125/U28/U1/set , 
        \U1209/U1122/U28/U1/clr , ysel, nyla, \U1209/U1122/U28/U1/set , 
        \U1209/U916_0_/U25/U1/clr , \yl[0] , \U1209/U916_0_/U25/U1/ob , 
        \U1209/U916_1_/U25/U1/clr , \yl[1] , \U1209/U916_1_/U25/U1/ob , 
        \U1209/U916_2_/U25/U1/clr , \yl[2] , \U1209/U916_2_/U25/U1/ob , 
        \U1209/U916_3_/U25/U1/clr , \yl[3] , \U1209/U916_3_/U25/U1/ob , 
        \U1213/nack[0] , \y[3] , \y[2] , \U1213/nack[1] , \y[1] , \U1213/net4 , 
        \y[0] , \U1213/U1125/U28/U1/clr , bsel, nba, \U1213/U1125/U28/U1/set , 
        \U1213/U1122/U28/U1/clr , dsel, nda, \U1213/U1122/U28/U1/set , 
        \U1213/U916_0_/U25/U1/clr , nya, \b[0] , \d[0] , 
        \U1213/U916_0_/U25/U1/ob , \U1213/U916_1_/U25/U1/clr , \b[1] , \d[1] , 
        \U1213/U916_1_/U25/U1/ob , \U1213/U916_2_/U25/U1/clr , \b[2] , \d[2] , 
        \U1213/U916_2_/U25/U1/ob , \U1213/U916_3_/U25/U1/clr , \b[3] , \d[3] , 
        \U1213/U916_3_/U25/U1/ob , \cdh[0] , \cdh[1] , \cdl[0] , \cdl[1] , 
        \cdh[2] , \cdh[3] , \cdl[2] , \cdl[3] , cg, \U1296/ng , net195, 
        \U1296/U1384/Z , \U1296/U1386/U25/U1/clr , \U1296/U1386/U25/U1/ob , dg, 
        \U1298/ng , net193, \U1298/U1384/Z , \U1298/U1386/U25/U1/clr , 
        \U1298/U1386/U25/U1/ob , bg, \U1306/ng , \U1306/U1384/Z , 
        \U1306/U1386/U25/U1/clr , \U1306/U1386/U25/U1/ob , ag, \U1295/ng , 
        \U1295/U1384/Z , \U1295/U1386/U25/U1/clr , \U1295/U1386/U25/U1/ob , 
        \U1297/s , \U1297/r , \U1297/nback , \U1297/naack , \U1297/reset , 
        \U1297/U1128/U28/U1/clr , \U1297/U1128/U28/U1/set , 
        \U1297/U1127/U28/U1/clr , \U1297/U1127/U28/U1/set , \U1300/s , 
        \U1300/r , \U1300/nback , \U1300/naack , \U1300/reset , 
        \U1300/U1128/U28/U1/clr , \U1300/U1128/U28/U1/set , 
        \U1300/U1127/U28/U1/clr , \U1300/U1127/U28/U1/set , 
        \U1289/U1150/U28/U1/clr , \U1289/bnreset , \U1289/U1150/U28/U1/set , 
        \U1289/U1152/U28/U1/clr , \U1289/U1152/U28/U1/set , 
        \U1289/U1149/U28/U1/clr , \U1289/U1149/U28/U1/set , 
        \U1289/U1151/U28/U1/clr , \U1289/U1151/U28/U1/set , 
        \U1289/U1148/net189 , \U1289/U1148/net192 , \U1289/U1148/net191 , 
        \U1289/U1148/net190 , \U1289/U1148/U1141/Z , \U1271/U1150/U28/U1/clr , 
        \U1271/bnreset , \U1271/U1150/U28/U1/set , \U1271/U1152/U28/U1/clr , 
        \U1271/U1152/U28/U1/set , \U1271/U1149/U28/U1/clr , 
        \U1271/U1149/U28/U1/set , \U1271/U1151/U28/U1/clr , 
        \U1271/U1151/U28/U1/set , \U1271/U1148/net189 , \U1271/U1148/net192 , 
        \U1271/U1148/net191 , \U1271/U1148/net190 , \U1271/U1148/U1141/Z , 
        \U1225/s , \U1225/r , \U1225/nback , \U1225/naack , \U1225/reset , 
        \U1308/nack[1] , \U1308/nack[0] ;
    assign eop_ack = eop_ack_wire;
    assign o[4] = eop_ack_wire;
    buf_2 U1231 ( .x(nbReset), .a(nReset) );
    and3_1 \U1194/U9  ( .x(eop_pass), .a(nxa), .b(naa), .c(eop) );
    ao222_1 \U1301/U18/U1/U1  ( .x(nlowack), .a(\twobitack[0] ), .b(
        \twobitack[1] ), .c(\twobitack[0] ), .d(nlowack), .e(\twobitack[1] ), 
        .f(nlowack) );
    ao222_1 \U1302/U18/U1/U1  ( .x(nhighack), .a(\twobitack[2] ), .b(
        \twobitack[3] ), .c(\twobitack[2] ), .d(nhighack), .e(\twobitack[3] ), 
        .f(nhighack) );
    aoi222_1 \U1018/U30/U1  ( .x(ia), .a(nhighack), .b(nlowack), .c(nhighack), 
        .d(\U1018/Z ), .e(nlowack), .f(\U1018/Z ) );
    inv_1 \U1018/U30/Uinv  ( .x(\U1018/Z ), .a(ia) );
    ao222_2 \U1038/U19/U1/U1  ( .x(eop_ack_wire), .a(eop_pass), .b(noa), .c(
        eop_pass), .d(eop_ack_wire), .e(noa), .f(eop_ack_wire) );
    inv_1 \U1270/U1147/U3  ( .x(\U1270/net189 ), .a(nbReset) );
    nor2_1 \U1270/U582/U5  ( .x(\U1270/net192 ), .a(il[4]), .b(ih[4]) );
    nor2_1 \U1270/U580/U5  ( .x(\U1270/net191 ), .a(il[5]), .b(ih[5]) );
    nor2_2 \U1270/U1146/U6  ( .x(net199), .a(\U1270/net190 ), .b(
        \U1270/net189 ) );
    aoi222_1 \U1270/U1141/U30/U1  ( .x(\U1270/net190 ), .a(\U1270/net191 ), 
        .b(\U1270/net192 ), .c(\U1270/net191 ), .d(\U1270/U1141/Z ), .e(
        \U1270/net192 ), .f(\U1270/U1141/Z ) );
    inv_1 \U1270/U1141/U30/Uinv  ( .x(\U1270/U1141/Z ), .a(\U1270/net190 ) );
    inv_1 \U1268/U1147/U3  ( .x(\U1268/net189 ), .a(nbReset) );
    nor2_1 \U1268/U582/U5  ( .x(\U1268/net192 ), .a(il[6]), .b(ih[6]) );
    nor2_1 \U1268/U580/U5  ( .x(\U1268/net191 ), .a(il[7]), .b(ih[7]) );
    nor2_2 \U1268/U1146/U6  ( .x(net194), .a(\U1268/net190 ), .b(
        \U1268/net189 ) );
    aoi222_1 \U1268/U1141/U30/U1  ( .x(\U1268/net190 ), .a(\U1268/net191 ), 
        .b(\U1268/net192 ), .c(\U1268/net191 ), .d(\U1268/U1141/Z ), .e(
        \U1268/net192 ), .f(\U1268/U1141/Z ) );
    inv_1 \U1268/U1141/U30/Uinv  ( .x(\U1268/U1141/Z ), .a(\U1268/net190 ) );
    nor2_1 \U1224/U1128/U5  ( .x(\U1224/nack[0] ), .a(\x[3] ), .b(\x[2] ) );
    nor3_1 \U1224/U1127/U7  ( .x(\U1224/nack[1] ), .a(\x[1] ), .b(\U1224/net4 
        ), .c(\x[0] ) );
    inv_1 \U1224/U907/U3  ( .x(\U1224/net4 ), .a(nbReset) );
    aoai211_1 \U1224/U1125/U28/U1/U1  ( .x(\U1224/U1125/U28/U1/clr ), .a(
        \U1224/nack[1] ), .b(\U1224/nack[0] ), .c(asel), .d(naa) );
    nand3_1 \U1224/U1125/U28/U1/U2  ( .x(\U1224/U1125/U28/U1/set ), .a(asel), 
        .b(\U1224/nack[1] ), .c(\U1224/nack[0] ) );
    nand2_2 \U1224/U1125/U28/U1/U3  ( .x(naa), .a(\U1224/U1125/U28/U1/clr ), 
        .b(\U1224/U1125/U28/U1/set ) );
    aoai211_1 \U1224/U1122/U28/U1/U1  ( .x(\U1224/U1122/U28/U1/clr ), .a(
        \U1224/nack[0] ), .b(\U1224/nack[1] ), .c(csel), .d(nca) );
    nand3_1 \U1224/U1122/U28/U1/U2  ( .x(\U1224/U1122/U28/U1/set ), .a(csel), 
        .b(\U1224/nack[0] ), .c(\U1224/nack[1] ) );
    nand2_2 \U1224/U1122/U28/U1/U3  ( .x(nca), .a(\U1224/U1122/U28/U1/clr ), 
        .b(\U1224/U1122/U28/U1/set ) );
    oa31_1 \U1224/U916_0_/U25/U1/Uclr  ( .x(\U1224/U916_0_/U25/U1/clr ), .a(
        nxa), .b(\a[0] ), .c(\c[0] ), .d(\x[0] ) );
    oaoi211_1 \U1224/U916_0_/U25/U1/Uaoi  ( .x(\U1224/U916_0_/U25/U1/ob ), .a(
        \a[0] ), .b(\c[0] ), .c(nxa), .d(\U1224/U916_0_/U25/U1/clr ) );
    inv_2 \U1224/U916_0_/U25/U1/Ui  ( .x(\x[0] ), .a(\U1224/U916_0_/U25/U1/ob 
        ) );
    oa31_1 \U1224/U916_1_/U25/U1/Uclr  ( .x(\U1224/U916_1_/U25/U1/clr ), .a(
        nxa), .b(\a[1] ), .c(\c[1] ), .d(\x[1] ) );
    oaoi211_1 \U1224/U916_1_/U25/U1/Uaoi  ( .x(\U1224/U916_1_/U25/U1/ob ), .a(
        \a[1] ), .b(\c[1] ), .c(nxa), .d(\U1224/U916_1_/U25/U1/clr ) );
    inv_2 \U1224/U916_1_/U25/U1/Ui  ( .x(\x[1] ), .a(\U1224/U916_1_/U25/U1/ob 
        ) );
    oa31_1 \U1224/U916_2_/U25/U1/Uclr  ( .x(\U1224/U916_2_/U25/U1/clr ), .a(
        nxa), .b(\a[2] ), .c(\c[2] ), .d(\x[2] ) );
    oaoi211_1 \U1224/U916_2_/U25/U1/Uaoi  ( .x(\U1224/U916_2_/U25/U1/ob ), .a(
        \a[2] ), .b(\c[2] ), .c(nxa), .d(\U1224/U916_2_/U25/U1/clr ) );
    inv_2 \U1224/U916_2_/U25/U1/Ui  ( .x(\x[2] ), .a(\U1224/U916_2_/U25/U1/ob 
        ) );
    oa31_1 \U1224/U916_3_/U25/U1/Uclr  ( .x(\U1224/U916_3_/U25/U1/clr ), .a(
        nxa), .b(\a[3] ), .c(\c[3] ), .d(\x[3] ) );
    oaoi211_1 \U1224/U916_3_/U25/U1/Uaoi  ( .x(\U1224/U916_3_/U25/U1/ob ), .a(
        \a[3] ), .b(\c[3] ), .c(nxa), .d(\U1224/U916_3_/U25/U1/clr ) );
    inv_2 \U1224/U916_3_/U25/U1/Ui  ( .x(\x[3] ), .a(\U1224/U916_3_/U25/U1/ob 
        ) );
    nor2_1 \U1209/U1128/U5  ( .x(\U1209/nack[0] ), .a(o[3]), .b(o[2]) );
    nor3_1 \U1209/U1127/U7  ( .x(\U1209/nack[1] ), .a(o[1]), .b(\U1209/net4 ), 
        .c(o[0]) );
    inv_1 \U1209/U907/U3  ( .x(\U1209/net4 ), .a(nbReset) );
    aoai211_1 \U1209/U1125/U28/U1/U1  ( .x(\U1209/U1125/U28/U1/clr ), .a(
        \U1209/nack[1] ), .b(\U1209/nack[0] ), .c(xsel), .d(nxa) );
    nand3_1 \U1209/U1125/U28/U1/U2  ( .x(\U1209/U1125/U28/U1/set ), .a(xsel), 
        .b(\U1209/nack[1] ), .c(\U1209/nack[0] ) );
    nand2_2 \U1209/U1125/U28/U1/U3  ( .x(nxa), .a(\U1209/U1125/U28/U1/clr ), 
        .b(\U1209/U1125/U28/U1/set ) );
    aoai211_1 \U1209/U1122/U28/U1/U1  ( .x(\U1209/U1122/U28/U1/clr ), .a(
        \U1209/nack[0] ), .b(\U1209/nack[1] ), .c(ysel), .d(nyla) );
    nand3_1 \U1209/U1122/U28/U1/U2  ( .x(\U1209/U1122/U28/U1/set ), .a(ysel), 
        .b(\U1209/nack[0] ), .c(\U1209/nack[1] ) );
    nand2_2 \U1209/U1122/U28/U1/U3  ( .x(nyla), .a(\U1209/U1122/U28/U1/clr ), 
        .b(\U1209/U1122/U28/U1/set ) );
    oa31_1 \U1209/U916_0_/U25/U1/Uclr  ( .x(\U1209/U916_0_/U25/U1/clr ), .a(
        noa), .b(\x[0] ), .c(\yl[0] ), .d(o[0]) );
    oaoi211_1 \U1209/U916_0_/U25/U1/Uaoi  ( .x(\U1209/U916_0_/U25/U1/ob ), .a(
        \x[0] ), .b(\yl[0] ), .c(noa), .d(\U1209/U916_0_/U25/U1/clr ) );
    inv_2 \U1209/U916_0_/U25/U1/Ui  ( .x(o[0]), .a(\U1209/U916_0_/U25/U1/ob )
         );
    oa31_1 \U1209/U916_1_/U25/U1/Uclr  ( .x(\U1209/U916_1_/U25/U1/clr ), .a(
        noa), .b(\x[1] ), .c(\yl[1] ), .d(o[1]) );
    oaoi211_1 \U1209/U916_1_/U25/U1/Uaoi  ( .x(\U1209/U916_1_/U25/U1/ob ), .a(
        \x[1] ), .b(\yl[1] ), .c(noa), .d(\U1209/U916_1_/U25/U1/clr ) );
    inv_2 \U1209/U916_1_/U25/U1/Ui  ( .x(o[1]), .a(\U1209/U916_1_/U25/U1/ob )
         );
    oa31_1 \U1209/U916_2_/U25/U1/Uclr  ( .x(\U1209/U916_2_/U25/U1/clr ), .a(
        noa), .b(\x[2] ), .c(\yl[2] ), .d(o[2]) );
    oaoi211_1 \U1209/U916_2_/U25/U1/Uaoi  ( .x(\U1209/U916_2_/U25/U1/ob ), .a(
        \x[2] ), .b(\yl[2] ), .c(noa), .d(\U1209/U916_2_/U25/U1/clr ) );
    inv_2 \U1209/U916_2_/U25/U1/Ui  ( .x(o[2]), .a(\U1209/U916_2_/U25/U1/ob )
         );
    oa31_1 \U1209/U916_3_/U25/U1/Uclr  ( .x(\U1209/U916_3_/U25/U1/clr ), .a(
        noa), .b(\x[3] ), .c(\yl[3] ), .d(o[3]) );
    oaoi211_1 \U1209/U916_3_/U25/U1/Uaoi  ( .x(\U1209/U916_3_/U25/U1/ob ), .a(
        \x[3] ), .b(\yl[3] ), .c(noa), .d(\U1209/U916_3_/U25/U1/clr ) );
    inv_2 \U1209/U916_3_/U25/U1/Ui  ( .x(o[3]), .a(\U1209/U916_3_/U25/U1/ob )
         );
    nor2_1 \U1213/U1128/U5  ( .x(\U1213/nack[0] ), .a(\y[3] ), .b(\y[2] ) );
    nor3_1 \U1213/U1127/U7  ( .x(\U1213/nack[1] ), .a(\y[1] ), .b(\U1213/net4 
        ), .c(\y[0] ) );
    inv_1 \U1213/U907/U3  ( .x(\U1213/net4 ), .a(nbReset) );
    aoai211_1 \U1213/U1125/U28/U1/U1  ( .x(\U1213/U1125/U28/U1/clr ), .a(
        \U1213/nack[1] ), .b(\U1213/nack[0] ), .c(bsel), .d(nba) );
    nand3_1 \U1213/U1125/U28/U1/U2  ( .x(\U1213/U1125/U28/U1/set ), .a(bsel), 
        .b(\U1213/nack[1] ), .c(\U1213/nack[0] ) );
    nand2_2 \U1213/U1125/U28/U1/U3  ( .x(nba), .a(\U1213/U1125/U28/U1/clr ), 
        .b(\U1213/U1125/U28/U1/set ) );
    aoai211_1 \U1213/U1122/U28/U1/U1  ( .x(\U1213/U1122/U28/U1/clr ), .a(
        \U1213/nack[0] ), .b(\U1213/nack[1] ), .c(dsel), .d(nda) );
    nand3_1 \U1213/U1122/U28/U1/U2  ( .x(\U1213/U1122/U28/U1/set ), .a(dsel), 
        .b(\U1213/nack[0] ), .c(\U1213/nack[1] ) );
    nand2_2 \U1213/U1122/U28/U1/U3  ( .x(nda), .a(\U1213/U1122/U28/U1/clr ), 
        .b(\U1213/U1122/U28/U1/set ) );
    oa31_1 \U1213/U916_0_/U25/U1/Uclr  ( .x(\U1213/U916_0_/U25/U1/clr ), .a(
        nya), .b(\b[0] ), .c(\d[0] ), .d(\y[0] ) );
    oaoi211_1 \U1213/U916_0_/U25/U1/Uaoi  ( .x(\U1213/U916_0_/U25/U1/ob ), .a(
        \b[0] ), .b(\d[0] ), .c(nya), .d(\U1213/U916_0_/U25/U1/clr ) );
    inv_2 \U1213/U916_0_/U25/U1/Ui  ( .x(\y[0] ), .a(\U1213/U916_0_/U25/U1/ob 
        ) );
    oa31_1 \U1213/U916_1_/U25/U1/Uclr  ( .x(\U1213/U916_1_/U25/U1/clr ), .a(
        nya), .b(\b[1] ), .c(\d[1] ), .d(\y[1] ) );
    oaoi211_1 \U1213/U916_1_/U25/U1/Uaoi  ( .x(\U1213/U916_1_/U25/U1/ob ), .a(
        \b[1] ), .b(\d[1] ), .c(nya), .d(\U1213/U916_1_/U25/U1/clr ) );
    inv_2 \U1213/U916_1_/U25/U1/Ui  ( .x(\y[1] ), .a(\U1213/U916_1_/U25/U1/ob 
        ) );
    oa31_1 \U1213/U916_2_/U25/U1/Uclr  ( .x(\U1213/U916_2_/U25/U1/clr ), .a(
        nya), .b(\b[2] ), .c(\d[2] ), .d(\y[2] ) );
    oaoi211_1 \U1213/U916_2_/U25/U1/Uaoi  ( .x(\U1213/U916_2_/U25/U1/ob ), .a(
        \b[2] ), .b(\d[2] ), .c(nya), .d(\U1213/U916_2_/U25/U1/clr ) );
    inv_2 \U1213/U916_2_/U25/U1/Ui  ( .x(\y[2] ), .a(\U1213/U916_2_/U25/U1/ob 
        ) );
    oa31_1 \U1213/U916_3_/U25/U1/Uclr  ( .x(\U1213/U916_3_/U25/U1/clr ), .a(
        nya), .b(\b[3] ), .c(\d[3] ), .d(\y[3] ) );
    oaoi211_1 \U1213/U916_3_/U25/U1/Uaoi  ( .x(\U1213/U916_3_/U25/U1/ob ), .a(
        \b[3] ), .b(\d[3] ), .c(nya), .d(\U1213/U916_3_/U25/U1/clr ) );
    inv_2 \U1213/U916_3_/U25/U1/Ui  ( .x(\y[3] ), .a(\U1213/U916_3_/U25/U1/ob 
        ) );
    and3_2 \U1210/U1138/U9  ( .x(\d[3] ), .a(\cdh[0] ), .b(nda), .c(\cdh[1] )
         );
    and3_2 \U1210/U1137/U9  ( .x(\d[2] ), .a(\cdl[0] ), .b(nda), .c(\cdh[1] )
         );
    and3_2 \U1210/U1139/U9  ( .x(\d[1] ), .a(\cdh[0] ), .b(nda), .c(\cdl[1] )
         );
    and3_2 \U1210/U1136/U9  ( .x(\d[0] ), .a(\cdl[0] ), .b(nda), .c(\cdl[1] )
         );
    and3_2 \U1162/U1138/U9  ( .x(\a[3] ), .a(ih[6]), .b(naa), .c(ih[7]) );
    and3_2 \U1162/U1137/U9  ( .x(\a[2] ), .a(il[6]), .b(naa), .c(ih[7]) );
    and3_2 \U1162/U1139/U9  ( .x(\a[1] ), .a(ih[6]), .b(naa), .c(il[7]) );
    and3_2 \U1162/U1136/U9  ( .x(\a[0] ), .a(il[6]), .b(naa), .c(il[7]) );
    and3_2 \U1211/U1138/U9  ( .x(\b[3] ), .a(ih[4]), .b(nba), .c(ih[5]) );
    and3_2 \U1211/U1137/U9  ( .x(\b[2] ), .a(il[4]), .b(nba), .c(ih[5]) );
    and3_2 \U1211/U1139/U9  ( .x(\b[1] ), .a(ih[4]), .b(nba), .c(il[5]) );
    and3_2 \U1211/U1136/U9  ( .x(\b[0] ), .a(il[4]), .b(nba), .c(il[5]) );
    and3_2 \U1163/U1138/U9  ( .x(\c[3] ), .a(\cdh[2] ), .b(nca), .c(\cdh[3] )
         );
    and3_2 \U1163/U1137/U9  ( .x(\c[2] ), .a(\cdl[2] ), .b(nca), .c(\cdh[3] )
         );
    and3_2 \U1163/U1139/U9  ( .x(\c[1] ), .a(\cdh[2] ), .b(nca), .c(\cdl[3] )
         );
    and3_2 \U1163/U1136/U9  ( .x(\c[0] ), .a(\cdl[2] ), .b(nca), .c(\cdl[3] )
         );
    and2_1 \U1296/U1385/U8  ( .x(cg), .a(nbReset), .b(\U1296/ng ) );
    aoi222_1 \U1296/U1384/U30/U1  ( .x(\U1296/ng ), .a(nca), .b(net195), .c(
        nca), .d(\U1296/U1384/Z ), .e(net195), .f(\U1296/U1384/Z ) );
    inv_1 \U1296/U1384/U30/Uinv  ( .x(\U1296/U1384/Z ), .a(\U1296/ng ) );
    oa31_1 \U1296/U1386/U25/U1/Uclr  ( .x(\U1296/U1386/U25/U1/clr ), .a(
        \twobitack[2] ), .b(cg), .c(nca), .d(net195) );
    oaoi211_1 \U1296/U1386/U25/U1/Uaoi  ( .x(\U1296/U1386/U25/U1/ob ), .a(cg), 
        .b(nca), .c(\twobitack[2] ), .d(\U1296/U1386/U25/U1/clr ) );
    inv_2 \U1296/U1386/U25/U1/Ui  ( .x(net195), .a(\U1296/U1386/U25/U1/ob ) );
    and2_1 \U1298/U1385/U8  ( .x(dg), .a(nbReset), .b(\U1298/ng ) );
    aoi222_1 \U1298/U1384/U30/U1  ( .x(\U1298/ng ), .a(nda), .b(net193), .c(
        nda), .d(\U1298/U1384/Z ), .e(net193), .f(\U1298/U1384/Z ) );
    inv_1 \U1298/U1384/U30/Uinv  ( .x(\U1298/U1384/Z ), .a(\U1298/ng ) );
    oa31_1 \U1298/U1386/U25/U1/Uclr  ( .x(\U1298/U1386/U25/U1/clr ), .a(
        \twobitack[0] ), .b(dg), .c(nda), .d(net193) );
    oaoi211_1 \U1298/U1386/U25/U1/Uaoi  ( .x(\U1298/U1386/U25/U1/ob ), .a(dg), 
        .b(nda), .c(\twobitack[0] ), .d(\U1298/U1386/U25/U1/clr ) );
    inv_2 \U1298/U1386/U25/U1/Ui  ( .x(net193), .a(\U1298/U1386/U25/U1/ob ) );
    and2_1 \U1306/U1385/U8  ( .x(bg), .a(nbReset), .b(\U1306/ng ) );
    aoi222_1 \U1306/U1384/U30/U1  ( .x(\U1306/ng ), .a(nba), .b(\twobitack[1] 
        ), .c(nba), .d(\U1306/U1384/Z ), .e(\twobitack[1] ), .f(
        \U1306/U1384/Z ) );
    inv_1 \U1306/U1384/U30/Uinv  ( .x(\U1306/U1384/Z ), .a(\U1306/ng ) );
    oa31_1 \U1306/U1386/U25/U1/Uclr  ( .x(\U1306/U1386/U25/U1/clr ), .a(net199
        ), .b(bg), .c(nba), .d(\twobitack[1] ) );
    oaoi211_1 \U1306/U1386/U25/U1/Uaoi  ( .x(\U1306/U1386/U25/U1/ob ), .a(bg), 
        .b(nba), .c(net199), .d(\U1306/U1386/U25/U1/clr ) );
    inv_2 \U1306/U1386/U25/U1/Ui  ( .x(\twobitack[1] ), .a(
        \U1306/U1386/U25/U1/ob ) );
    and2_1 \U1295/U1385/U8  ( .x(ag), .a(nbReset), .b(\U1295/ng ) );
    aoi222_1 \U1295/U1384/U30/U1  ( .x(\U1295/ng ), .a(naa), .b(\twobitack[3] 
        ), .c(naa), .d(\U1295/U1384/Z ), .e(\twobitack[3] ), .f(
        \U1295/U1384/Z ) );
    inv_1 \U1295/U1384/U30/Uinv  ( .x(\U1295/U1384/Z ), .a(\U1295/ng ) );
    oa31_1 \U1295/U1386/U25/U1/Uclr  ( .x(\U1295/U1386/U25/U1/clr ), .a(net194
        ), .b(ag), .c(naa), .d(\twobitack[3] ) );
    oaoi211_1 \U1295/U1386/U25/U1/Uaoi  ( .x(\U1295/U1386/U25/U1/ob ), .a(ag), 
        .b(naa), .c(net194), .d(\U1295/U1386/U25/U1/clr ) );
    inv_2 \U1295/U1386/U25/U1/Ui  ( .x(\twobitack[3] ), .a(
        \U1295/U1386/U25/U1/ob ) );
    nand2_1 \U1297/U1131/U5  ( .x(\U1297/s ), .a(\U1297/r ), .b(\U1297/nback )
         );
    nand2_1 \U1297/U1103/U5  ( .x(\U1297/r ), .a(\U1297/naack ), .b(\U1297/s )
         );
    inv_1 \U1297/U1111/U3  ( .x(\U1297/reset ), .a(nbReset) );
    inv_1 \U1297/U1112/U3  ( .x(\U1297/naack ), .a(naa) );
    nor2_1 \U1297/U1130/U5  ( .x(\U1297/nback ), .a(nca), .b(\U1297/reset ) );
    aoai211_1 \U1297/U1128/U28/U1/U1  ( .x(\U1297/U1128/U28/U1/clr ), .a(
        \U1297/r ), .b(\U1297/naack ), .c(cg), .d(csel) );
    nand3_1 \U1297/U1128/U28/U1/U2  ( .x(\U1297/U1128/U28/U1/set ), .a(cg), 
        .b(\U1297/r ), .c(\U1297/naack ) );
    nand2_2 \U1297/U1128/U28/U1/U3  ( .x(csel), .a(\U1297/U1128/U28/U1/clr ), 
        .b(\U1297/U1128/U28/U1/set ) );
    aoai211_1 \U1297/U1127/U28/U1/U1  ( .x(\U1297/U1127/U28/U1/clr ), .a(
        \U1297/s ), .b(\U1297/nback ), .c(ag), .d(asel) );
    nand3_1 \U1297/U1127/U28/U1/U2  ( .x(\U1297/U1127/U28/U1/set ), .a(ag), 
        .b(\U1297/s ), .c(\U1297/nback ) );
    nand2_2 \U1297/U1127/U28/U1/U3  ( .x(asel), .a(\U1297/U1127/U28/U1/clr ), 
        .b(\U1297/U1127/U28/U1/set ) );
    nand2_1 \U1300/U1131/U5  ( .x(\U1300/s ), .a(\U1300/r ), .b(\U1300/nback )
         );
    nand2_1 \U1300/U1103/U5  ( .x(\U1300/r ), .a(\U1300/naack ), .b(\U1300/s )
         );
    inv_1 \U1300/U1111/U3  ( .x(\U1300/reset ), .a(nbReset) );
    inv_1 \U1300/U1112/U3  ( .x(\U1300/naack ), .a(nba) );
    nor2_1 \U1300/U1130/U5  ( .x(\U1300/nback ), .a(nda), .b(\U1300/reset ) );
    aoai211_1 \U1300/U1128/U28/U1/U1  ( .x(\U1300/U1128/U28/U1/clr ), .a(
        \U1300/r ), .b(\U1300/naack ), .c(dg), .d(dsel) );
    nand3_1 \U1300/U1128/U28/U1/U2  ( .x(\U1300/U1128/U28/U1/set ), .a(dg), 
        .b(\U1300/r ), .c(\U1300/naack ) );
    nand2_2 \U1300/U1128/U28/U1/U3  ( .x(dsel), .a(\U1300/U1128/U28/U1/clr ), 
        .b(\U1300/U1128/U28/U1/set ) );
    aoai211_1 \U1300/U1127/U28/U1/U1  ( .x(\U1300/U1127/U28/U1/clr ), .a(
        \U1300/s ), .b(\U1300/nback ), .c(bg), .d(bsel) );
    nand3_1 \U1300/U1127/U28/U1/U2  ( .x(\U1300/U1127/U28/U1/set ), .a(bg), 
        .b(\U1300/s ), .c(\U1300/nback ) );
    nand2_2 \U1300/U1127/U28/U1/U3  ( .x(bsel), .a(\U1300/U1127/U28/U1/clr ), 
        .b(\U1300/U1127/U28/U1/set ) );
    aoai211_1 \U1289/U1150/U28/U1/U1  ( .x(\U1289/U1150/U28/U1/clr ), .a(il[2]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdl[2] ) );
    nand3_1 \U1289/U1150/U28/U1/U2  ( .x(\U1289/U1150/U28/U1/set ), .a(net195), 
        .b(il[2]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1150/U28/U1/U3  ( .x(\cdl[2] ), .a(
        \U1289/U1150/U28/U1/clr ), .b(\U1289/U1150/U28/U1/set ) );
    aoai211_1 \U1289/U1152/U28/U1/U1  ( .x(\U1289/U1152/U28/U1/clr ), .a(il[3]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdl[3] ) );
    nand3_1 \U1289/U1152/U28/U1/U2  ( .x(\U1289/U1152/U28/U1/set ), .a(net195), 
        .b(il[3]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1152/U28/U1/U3  ( .x(\cdl[3] ), .a(
        \U1289/U1152/U28/U1/clr ), .b(\U1289/U1152/U28/U1/set ) );
    aoai211_1 \U1289/U1149/U28/U1/U1  ( .x(\U1289/U1149/U28/U1/clr ), .a(ih[2]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdh[2] ) );
    nand3_1 \U1289/U1149/U28/U1/U2  ( .x(\U1289/U1149/U28/U1/set ), .a(net195), 
        .b(ih[2]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1149/U28/U1/U3  ( .x(\cdh[2] ), .a(
        \U1289/U1149/U28/U1/clr ), .b(\U1289/U1149/U28/U1/set ) );
    aoai211_1 \U1289/U1151/U28/U1/U1  ( .x(\U1289/U1151/U28/U1/clr ), .a(ih[3]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdh[3] ) );
    nand3_1 \U1289/U1151/U28/U1/U2  ( .x(\U1289/U1151/U28/U1/set ), .a(net195), 
        .b(ih[3]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1151/U28/U1/U3  ( .x(\cdh[3] ), .a(
        \U1289/U1151/U28/U1/clr ), .b(\U1289/U1151/U28/U1/set ) );
    inv_1 \U1289/U1148/U1147/U3  ( .x(\U1289/U1148/net189 ), .a(
        \U1289/bnreset ) );
    nor2_1 \U1289/U1148/U582/U5  ( .x(\U1289/U1148/net192 ), .a(\cdl[3] ), .b(
        \cdh[3] ) );
    nor2_1 \U1289/U1148/U580/U5  ( .x(\U1289/U1148/net191 ), .a(\cdl[2] ), .b(
        \cdh[2] ) );
    nor2_2 \U1289/U1148/U1146/U6  ( .x(\twobitack[2] ), .a(
        \U1289/U1148/net190 ), .b(\U1289/U1148/net189 ) );
    aoi222_1 \U1289/U1148/U1141/U30/U1  ( .x(\U1289/U1148/net190 ), .a(
        \U1289/U1148/net191 ), .b(\U1289/U1148/net192 ), .c(
        \U1289/U1148/net191 ), .d(\U1289/U1148/U1141/Z ), .e(
        \U1289/U1148/net192 ), .f(\U1289/U1148/U1141/Z ) );
    inv_1 \U1289/U1148/U1141/U30/Uinv  ( .x(\U1289/U1148/U1141/Z ), .a(
        \U1289/U1148/net190 ) );
    aoai211_1 \U1271/U1150/U28/U1/U1  ( .x(\U1271/U1150/U28/U1/clr ), .a(il[0]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdl[0] ) );
    nand3_1 \U1271/U1150/U28/U1/U2  ( .x(\U1271/U1150/U28/U1/set ), .a(net193), 
        .b(il[0]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1150/U28/U1/U3  ( .x(\cdl[0] ), .a(
        \U1271/U1150/U28/U1/clr ), .b(\U1271/U1150/U28/U1/set ) );
    aoai211_1 \U1271/U1152/U28/U1/U1  ( .x(\U1271/U1152/U28/U1/clr ), .a(il[1]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdl[1] ) );
    nand3_1 \U1271/U1152/U28/U1/U2  ( .x(\U1271/U1152/U28/U1/set ), .a(net193), 
        .b(il[1]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1152/U28/U1/U3  ( .x(\cdl[1] ), .a(
        \U1271/U1152/U28/U1/clr ), .b(\U1271/U1152/U28/U1/set ) );
    aoai211_1 \U1271/U1149/U28/U1/U1  ( .x(\U1271/U1149/U28/U1/clr ), .a(ih[0]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdh[0] ) );
    nand3_1 \U1271/U1149/U28/U1/U2  ( .x(\U1271/U1149/U28/U1/set ), .a(net193), 
        .b(ih[0]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1149/U28/U1/U3  ( .x(\cdh[0] ), .a(
        \U1271/U1149/U28/U1/clr ), .b(\U1271/U1149/U28/U1/set ) );
    aoai211_1 \U1271/U1151/U28/U1/U1  ( .x(\U1271/U1151/U28/U1/clr ), .a(ih[1]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdh[1] ) );
    nand3_1 \U1271/U1151/U28/U1/U2  ( .x(\U1271/U1151/U28/U1/set ), .a(net193), 
        .b(ih[1]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1151/U28/U1/U3  ( .x(\cdh[1] ), .a(
        \U1271/U1151/U28/U1/clr ), .b(\U1271/U1151/U28/U1/set ) );
    inv_1 \U1271/U1148/U1147/U3  ( .x(\U1271/U1148/net189 ), .a(
        \U1271/bnreset ) );
    nor2_1 \U1271/U1148/U582/U5  ( .x(\U1271/U1148/net192 ), .a(\cdl[1] ), .b(
        \cdh[1] ) );
    nor2_1 \U1271/U1148/U580/U5  ( .x(\U1271/U1148/net191 ), .a(\cdl[0] ), .b(
        \cdh[0] ) );
    nor2_2 \U1271/U1148/U1146/U6  ( .x(\twobitack[0] ), .a(
        \U1271/U1148/net190 ), .b(\U1271/U1148/net189 ) );
    aoi222_1 \U1271/U1148/U1141/U30/U1  ( .x(\U1271/U1148/net190 ), .a(
        \U1271/U1148/net191 ), .b(\U1271/U1148/net192 ), .c(
        \U1271/U1148/net191 ), .d(\U1271/U1148/U1141/Z ), .e(
        \U1271/U1148/net192 ), .f(\U1271/U1148/U1141/Z ) );
    inv_1 \U1271/U1148/U1141/U30/Uinv  ( .x(\U1271/U1148/U1141/Z ), .a(
        \U1271/U1148/net190 ) );
    nand2_1 \U1225/U1128/U5  ( .x(\U1225/s ), .a(\U1225/r ), .b(\U1225/nback )
         );
    nand2_1 \U1225/U1103/U5  ( .x(\U1225/r ), .a(\U1225/naack ), .b(\U1225/s )
         );
    inv_1 \U1225/U1111/U3  ( .x(\U1225/reset ), .a(nbReset) );
    inv_1 \U1225/U1112/U3  ( .x(\U1225/naack ), .a(nxa) );
    nor2_1 \U1225/U1127/U5  ( .x(\U1225/nback ), .a(nyla), .b(\U1225/reset )
         );
    and2_2 \U1225/U1129/U8  ( .x(xsel), .a(\U1225/nback ), .b(\U1225/s ) );
    and2_2 \U1225/U1124/U8  ( .x(ysel), .a(\U1225/r ), .b(\U1225/naack ) );
    and3_4 \U1308/U20/U9  ( .x(nya), .a(\U1308/nack[1] ), .b(\U1308/nack[0] ), 
        .c(nbReset) );
    nor2_1 \U1308/U18/U5  ( .x(\U1308/nack[0] ), .a(\yl[3] ), .b(\yl[0] ) );
    nor2_1 \U1308/U19/U5  ( .x(\U1308/nack[1] ), .a(\yl[1] ), .b(\yl[2] ) );
    ao222_2 \U1308/U15_0_/U19/U1/U1  ( .x(\yl[0] ), .a(\y[0] ), .b(nyla), .c(
        \y[0] ), .d(\yl[0] ), .e(nyla), .f(\yl[0] ) );
    ao222_2 \U1308/U15_1_/U19/U1/U1  ( .x(\yl[1] ), .a(\y[1] ), .b(nyla), .c(
        \y[1] ), .d(\yl[1] ), .e(nyla), .f(\yl[1] ) );
    ao222_2 \U1308/U15_2_/U19/U1/U1  ( .x(\yl[2] ), .a(\y[2] ), .b(nyla), .c(
        \y[2] ), .d(\yl[2] ), .e(nyla), .f(\yl[2] ) );
    ao222_2 \U1308/U15_3_/U19/U1/U1  ( .x(\yl[3] ), .a(\y[3] ), .b(nyla), .c(
        \y[3] ), .d(\yl[3] ), .e(nyla), .f(\yl[3] ) );
    buf_3 U1 ( .x(\U1271/bnreset ), .a(nbReset) );
    buf_3 U2 ( .x(\U1289/bnreset ), .a(nbReset) );
endmodule


module chain_mergepackets_0 ( naa, nba, o, a, b, nReset, noa );
output [4:0] o;
input  [4:0] a;
input  [4:0] b;
input  nReset, noa;
output naa, nba;
    wire as, seta, asel, bsel, setb, reset, \noack[1] , \noack[0] , 
        \U916_0_/U25/U1/clr , \U916_0_/U25/U1/ob , \U916_1_/U25/U1/clr , 
        \U916_1_/U25/U1/ob , \U916_2_/U25/U1/clr , \U916_2_/U25/U1/ob , 
        \U916_3_/U25/U1/clr , \U916_3_/U25/U1/ob ;
    and2_1 \U1155/U8  ( .x(as), .a(seta), .b(asel) );
    nand2_1 \U1145/U5  ( .x(asel), .a(bsel), .b(seta) );
    nand2_1 \U1103/U5  ( .x(bsel), .a(setb), .b(asel) );
    inv_1 \U1135/U3  ( .x(reset), .a(nReset) );
    inv_1 \U1134/U3  ( .x(setb), .a(a[4]) );
    and3_2 \U1154/U9  ( .x(naa), .a(\noack[1] ), .b(\noack[0] ), .c(as) );
    nor3_1 \U1127/U7  ( .x(\noack[0] ), .a(o[1]), .b(reset), .c(o[0]) );
    nor2_1 \U1132/U5  ( .x(\noack[1] ), .a(o[3]), .b(o[2]) );
    oa31_1 \U916_0_/U25/U1/Uclr  ( .x(\U916_0_/U25/U1/clr ), .a(noa), .b(a[0]), 
        .c(b[0]), .d(o[0]) );
    oaoi211_1 \U916_0_/U25/U1/Uaoi  ( .x(\U916_0_/U25/U1/ob ), .a(a[0]), .b(b
        [0]), .c(noa), .d(\U916_0_/U25/U1/clr ) );
    inv_2 \U916_0_/U25/U1/Ui  ( .x(o[0]), .a(\U916_0_/U25/U1/ob ) );
    oa31_1 \U916_1_/U25/U1/Uclr  ( .x(\U916_1_/U25/U1/clr ), .a(noa), .b(a[1]), 
        .c(b[1]), .d(o[1]) );
    oaoi211_1 \U916_1_/U25/U1/Uaoi  ( .x(\U916_1_/U25/U1/ob ), .a(a[1]), .b(b
        [1]), .c(noa), .d(\U916_1_/U25/U1/clr ) );
    inv_2 \U916_1_/U25/U1/Ui  ( .x(o[1]), .a(\U916_1_/U25/U1/ob ) );
    oa31_1 \U916_2_/U25/U1/Uclr  ( .x(\U916_2_/U25/U1/clr ), .a(noa), .b(a[2]), 
        .c(b[2]), .d(o[2]) );
    oaoi211_1 \U916_2_/U25/U1/Uaoi  ( .x(\U916_2_/U25/U1/ob ), .a(a[2]), .b(b
        [2]), .c(noa), .d(\U916_2_/U25/U1/clr ) );
    inv_2 \U916_2_/U25/U1/Ui  ( .x(o[2]), .a(\U916_2_/U25/U1/ob ) );
    oa31_1 \U916_3_/U25/U1/Uclr  ( .x(\U916_3_/U25/U1/clr ), .a(noa), .b(a[3]), 
        .c(b[3]), .d(o[3]) );
    oaoi211_1 \U916_3_/U25/U1/Uaoi  ( .x(\U916_3_/U25/U1/ob ), .a(a[3]), .b(b
        [3]), .c(noa), .d(\U916_3_/U25/U1/clr ) );
    inv_2 \U916_3_/U25/U1/Ui  ( .x(o[3]), .a(\U916_3_/U25/U1/ob ) );
    ao222_2 \U1148/U19/U1/U1  ( .x(o[4]), .a(noa), .b(b[4]), .c(noa), .d(o[4]), 
        .e(b[4]), .f(o[4]) );
    aoi21_1 \U1153/U11  ( .x(seta), .a(o[4]), .b(setb), .c(reset) );
    and3_3 U1 ( .x(nba), .a(bsel), .b(\noack[0] ), .c(\noack[1] ) );
endmodule


module initiator_iport ( cack, chaincommand, err, nchainresponseack, nrouteack, 
    rd, routetxreq, rrnw, a, chainresponse, col, crnw, itag, lock, nReset, 
    nchaincommandack, pred, rack, route, routetxack, seq, size, wd );
output [4:0] chaincommand;
output [1:0] err;
output [63:0] rd;
output [1:0] rrnw;
input  [63:0] a;
input  [4:0] chainresponse;
input  [5:0] col;
input  [1:0] crnw;
input  [9:0] itag;
input  [1:0] lock;
input  [1:0] pred;
input  [4:0] route;
input  [1:0] seq;
input  [3:0] size;
input  [63:0] wd;
input  nReset, nchaincommandack, rack, routetxack;
output cack, nchainresponseack, nrouteack, routetxreq;
    wire nircba, nResetb, responseack, rstatusack, \irbl[7] , \irbl[6] , 
        \irbl[5] , \irbl[4] , \irbl[3] , \irbl[2] , \irbl[1] , \irbl[0] , 
        \irbh[7] , \irbh[6] , \irbh[5] , \irbh[4] , \irbh[3] , \irbh[2] , 
        \irbh[1] , \irbh[0] , \rstatus[1] , \rstatus[0] , ictrlack, 
        \can_defer[0] , net116, ncstatusack, pltxreq, tok_ack, \cstatus[0] , 
        \cstatus[1] , net115, net128, pltxack, icmdack, nicba, \icbl[7] , 
        \icbl[6] , \icbl[5] , \icbl[4] , \icbl[3] , \icbl[2] , \icbl[1] , 
        \icbl[0] , \icbh[7] , \icbh[6] , \icbh[5] , \icbh[4] , \icbh[3] , 
        \icbh[2] , \icbh[1] , \icbh[0] , nipayloadack, \ipayload[4] , 
        \ipayload[3] , \ipayload[2] , \ipayload[1] , \ipayload[0] , net170, 
        reset, net165, \U1662/U28/U1/clr , \U1662/U28/U1/set ;
    chain_irdemuxNew_0 U1442 ( .err(err), .ncback(nircba), .rd(rd), .rnw(rrnw), 
        .status({\rstatus[1] , \rstatus[0] }), .cbh({\irbh[7] , \irbh[6] , 
        \irbh[5] , \irbh[4] , \irbh[3] , \irbh[2] , \irbh[1] , \irbh[0] }), 
        .cbl({\irbl[7] , \irbl[6] , \irbl[5] , \irbl[4] , \irbl[3] , \irbl[2] , 
        \irbl[1] , \irbl[0] }), .nReset(nResetb), .nack(responseack), 
        .statusack(rstatusack) );
    chain_fr2dr_byte_3 chain_decoder ( .nia(nchainresponseack), .oh({\irbh[7] , 
        \irbh[6] , \irbh[5] , \irbh[4] , \irbh[3] , \irbh[2] , \irbh[1] , 
        \irbh[0] }), .ol({\irbl[7] , \irbl[6] , \irbl[5] , \irbl[4] , 
        \irbl[3] , \irbl[2] , \irbl[1] , \irbl[0] }), .i(chainresponse), 
        .nReset(nResetb), .noa(nircba) );
    chain_ic_ctrl_0 cmd_ctrl ( .ack(ictrlack), .candefer(\can_defer[0] ), 
        .eop(net116), .nstatack(ncstatusack), .pltxreq(pltxreq), .routetxreq(
        routetxreq), .tok_ack(tok_ack), .accept(\cstatus[0] ), .candefer_ack({
        1'b0, \can_defer[0] }), .defer(\cstatus[1] ), .eopack(net115), .lock(
        lock), .nReset(net128), .pltxack(pltxack), .routetxack(routetxack), 
        .tok_err(err[1]), .tok_ok(err[0]) );
    chain_icmux_0 cmd_mux ( .ack(icmdack), .chainh({\icbh[7] , \icbh[6] , 
        \icbh[5] , \icbh[4] , \icbh[3] , \icbh[2] , \icbh[1] , \icbh[0] }), 
        .chainl({\icbl[7] , \icbl[6] , \icbl[5] , \icbl[4] , \icbl[3] , 
        \icbl[2] , \icbl[1] , \icbl[0] }), .sendack(pltxack), .addr(a), .col(
        col), .itag(itag), .lock(lock), .nReset(net128), .nia(nicba), .pred(
        pred), .rnw(crnw), .sendreq(pltxreq), .seq(seq), .size(size), .wd(wd)
         );
    chain_dr2fr_byte_0 U1604 ( .eop_ack(net115), .ia(nicba), .o({\ipayload[4] , 
        \ipayload[3] , \ipayload[2] , \ipayload[1] , \ipayload[0] }), .eop(
        net116), .ih({\icbh[7] , \icbh[6] , \icbh[5] , \icbh[4] , \icbh[3] , 
        \icbh[2] , \icbh[1] , \icbh[0] }), .il({\icbl[7] , \icbl[6] , 
        \icbl[5] , \icbl[4] , \icbl[3] , \icbl[2] , \icbl[1] , \icbl[0] }), 
        .nReset(net128), .noa(nipayloadack) );
    chain_mergepackets_0 U1605 ( .naa(nrouteack), .nba(nipayloadack), .o(
        chaincommand), .a(route), .b({\ipayload[4] , \ipayload[3] , 
        \ipayload[2] , \ipayload[1] , \ipayload[0] }), .nReset(net128), .noa(
        nchaincommandack) );
    and2_1 U1676 ( .x(cack), .a(net170), .b(nResetb) );
    inv_4 \U1643/U3  ( .x(net128), .a(reset) );
    or2_4 \U1660/U12  ( .x(net165), .a(\cstatus[0] ), .b(\cstatus[1] ) );
    or2_1 \U1661/U12  ( .x(rstatusack), .a(net165), .b(reset) );
    ao222_2 \status_pipe_0_/U19/U1/U1  ( .x(\cstatus[0] ), .a(\rstatus[0] ), 
        .b(ncstatusack), .c(\rstatus[0] ), .d(\cstatus[0] ), .e(ncstatusack), 
        .f(\cstatus[0] ) );
    ao222_2 \status_pipe_1_/U19/U1/U1  ( .x(\cstatus[1] ), .a(\rstatus[1] ), 
        .b(ncstatusack), .c(\rstatus[1] ), .d(\cstatus[1] ), .e(ncstatusack), 
        .f(\cstatus[1] ) );
    ao222_1 \U1609/U18/U1/U1  ( .x(net170), .a(ictrlack), .b(icmdack), .c(
        ictrlack), .d(net170), .e(icmdack), .f(net170) );
    aoai211_1 \U1662/U28/U1/U1  ( .x(\U1662/U28/U1/clr ), .a(rack), .b(nResetb
        ), .c(tok_ack), .d(responseack) );
    nand3_1 \U1662/U28/U1/U2  ( .x(\U1662/U28/U1/set ), .a(tok_ack), .b(rack), 
        .c(nResetb) );
    nand2_2 \U1662/U28/U1/U3  ( .x(responseack), .a(\U1662/U28/U1/clr ), .b(
        \U1662/U28/U1/set ) );
    inv_2 U1 ( .x(reset), .a(nResetb) );
    buf_3 U2 ( .x(nResetb), .a(nReset) );
endmodule


module master_if_iport ( nReset, mc_req, mc_we, mc_mult, mc_prd, mc_seq, mc_ts, 
    mc_sel, mc_adr, mc_dat, mc_ack, mr_req, mr_we, mr_err, mr_rty, mr_acc, 
    mr_ts, mr_sel, mr_dat, mr_ack, chaincommand, nchaincommandack, 
    chainresponse, nchainresponseack, e_bare, e_dm, e_im, e_wish, r_bare, r_dm, 
    r_im, r_wish, tag_id, force_bare );
input  [2:0] mc_ts;
input  [3:0] mc_sel;
input  [31:0] mc_adr;
input  [31:0] mc_dat;
output [2:0] mr_ts;
output [3:0] mr_sel;
output [31:0] mr_dat;
output [4:0] chaincommand;
input  [4:0] chainresponse;
input  [3:0] e_bare;
input  [3:0] e_dm;
input  [3:0] e_im;
input  [3:0] e_wish;
input  [3:0] r_bare;
input  [3:0] r_dm;
input  [3:0] r_im;
input  [3:0] r_wish;
input  [4:0] tag_id;
input  nReset, mc_req, mc_we, mc_mult, mc_prd, mc_seq, mr_ack, 
    nchaincommandack, force_bare;
output mc_ack, mr_req, mr_we, mr_err, mr_rty, mr_acc, nchainresponseack;
    wire reset, ci_ack, ri_ack, \ri_rnw[1] , \ri_rnw[0] , \ri_err[1] , 
        \ri_err[0] , \ri_rd[63] , \ri_rd[62] , \ri_rd[61] , \ri_rd[60] , 
        \ri_rd[59] , \ri_rd[58] , \ri_rd[57] , \ri_rd[56] , \ri_rd[55] , 
        \ri_rd[54] , \ri_rd[53] , \ri_rd[52] , \ri_rd[51] , \ri_rd[50] , 
        \ri_rd[49] , \ri_rd[48] , \ri_rd[47] , \ri_rd[46] , \ri_rd[45] , 
        \ri_rd[44] , \ri_rd[43] , \ri_rd[42] , \ri_rd[41] , \ri_rd[40] , 
        \ri_rd[39] , \ri_rd[38] , \ri_rd[37] , \ri_rd[36] , \ri_rd[35] , 
        \ri_rd[34] , \ri_rd[33] , \ri_rd[32] , \ri_rd[31] , \ri_rd[30] , 
        \ri_rd[29] , \ri_rd[28] , \ri_rd[27] , \ri_rd[26] , \ri_rd[25] , 
        \ri_rd[24] , \ri_rd[23] , \ri_rd[22] , \ri_rd[21] , \ri_rd[20] , 
        \ri_rd[19] , \ri_rd[18] , \ri_rd[17] , \ri_rd[16] , \ri_rd[15] , 
        \ri_rd[14] , \ri_rd[13] , \ri_rd[12] , \ri_rd[11] , \ri_rd[10] , 
        \ri_rd[9] , \ri_rd[8] , \ri_rd[7] , \ri_rd[6] , \ri_rd[5] , \ri_rd[4] , 
        \ri_rd[3] , \ri_rd[2] , \ri_rd[1] , \ri_rd[0] , \ci_col[5] , 
        \ci_col[4] , \ci_col[3] , \ci_col[2] , \ci_col[1] , \ci_col[0] , 
        \ci_rnw[1] , \ci_rnw[0] , \ci_a[63] , \ci_a[62] , \ci_a[61] , 
        \ci_a[60] , \ci_a[59] , \ci_a[58] , \ci_a[57] , \ci_a[56] , \ci_a[55] , 
        \ci_a[54] , \ci_a[53] , \ci_a[52] , \ci_a[51] , \ci_a[50] , \ci_a[49] , 
        \ci_a[48] , \ci_a[47] , \ci_a[46] , \ci_a[45] , \ci_a[44] , \ci_a[43] , 
        \ci_a[42] , \ci_a[41] , \ci_a[40] , \ci_a[39] , \ci_a[38] , \ci_a[37] , 
        \ci_a[36] , \ci_a[35] , \ci_a[34] , \ci_a[33] , \ci_a[32] , \ci_a[31] , 
        \ci_a[30] , \ci_a[29] , \ci_a[28] , \ci_a[27] , \ci_a[26] , \ci_a[25] , 
        \ci_a[24] , \ci_a[23] , \ci_a[22] , \ci_a[21] , \ci_a[20] , \ci_a[19] , 
        \ci_a[18] , \ci_a[17] , \ci_a[16] , \ci_a[15] , \ci_a[14] , \ci_a[13] , 
        \ci_a[12] , \ci_a[11] , \ci_a[10] , \ci_a[9] , \ci_a[8] , \ci_a[7] , 
        \ci_a[6] , \ci_a[5] , \ci_a[4] , \ci_a[3] , \ci_a[2] , \ci_a[1] , 
        \ci_a[0] , \ci_lock[1] , \ci_lock[0] , \ci_wd[63] , \ci_wd[62] , 
        \ci_wd[61] , \ci_wd[60] , \ci_wd[59] , \ci_wd[58] , \ci_wd[57] , 
        \ci_wd[56] , \ci_wd[55] , \ci_wd[54] , \ci_wd[53] , \ci_wd[52] , 
        \ci_wd[51] , \ci_wd[50] , \ci_wd[49] , \ci_wd[48] , \ci_wd[47] , 
        \ci_wd[46] , \ci_wd[45] , \ci_wd[44] , \ci_wd[43] , \ci_wd[42] , 
        \ci_wd[41] , \ci_wd[40] , \ci_wd[39] , \ci_wd[38] , \ci_wd[37] , 
        \ci_wd[36] , \ci_wd[35] , \ci_wd[34] , \ci_wd[33] , \ci_wd[32] , 
        \ci_wd[31] , \ci_wd[30] , \ci_wd[29] , \ci_wd[28] , \ci_wd[27] , 
        \ci_wd[26] , \ci_wd[25] , \ci_wd[24] , \ci_wd[23] , \ci_wd[22] , 
        \ci_wd[21] , \ci_wd[20] , \ci_wd[19] , \ci_wd[18] , \ci_wd[17] , 
        \ci_wd[16] , \ci_wd[15] , \ci_wd[14] , \ci_wd[13] , \ci_wd[12] , 
        \ci_wd[11] , \ci_wd[10] , \ci_wd[9] , \ci_wd[8] , \ci_wd[7] , 
        \ci_wd[6] , \ci_wd[5] , \ci_wd[4] , \ci_wd[3] , \ci_wd[2] , \ci_wd[1] , 
        \ci_wd[0] , \ci_itag[9] , \ci_itag[8] , \ci_itag[7] , \ci_itag[6] , 
        \ci_itag[5] , \ci_itag[4] , \ci_itag[3] , \ci_itag[2] , \ci_itag[1] , 
        \ci_itag[0] , \ci_size[3] , \ci_size[2] , \ci_size[1] , \ci_size[0] , 
        \ci_pred[1] , \ci_pred[0] , \ci_seq[1] , \ci_seq[0] , \i_rl[3] , 
        \i_rl[2] , \i_rl[1] , \i_rl[0] , \i_rh[3] , \i_rh[2] , \i_rh[1] , 
        SYNOPSYS_UNCONNECTED_2, \i_el[3] , \i_el[2] , \i_el[1] , \i_el[0] , 
        SYNOPSYS_UNCONNECTED_1, \i_eh[2] , \i_eh[1] , \i_eh[0] , routetx_ack, 
        nroute_ack, routetx_req, \route[4] , SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4, \route[1] , \route[0] ;
    assign mr_rty = 1'b0;
    assign mr_acc = 1'b0;
    assign mr_ts[2] = 1'b0;
    assign mr_ts[1] = 1'b0;
    assign mr_ts[0] = 1'b0;
    assign mr_sel[3] = 1'b0;
    assign mr_sel[2] = 1'b0;
    assign mr_sel[1] = 1'b0;
    assign mr_sel[0] = 1'b0;
    inv_2 U1 ( .x(reset), .a(nReset) );
    m2cp_iport master2chainif ( .req_in(mc_req), .ts_o(mc_ts), .sel_o(mc_sel), 
        .mult_o(mc_mult), .we_o(mc_we), .prd_o(mc_prd), .seq_o(mc_seq), 
        .adr_o(mc_adr), .dat_o(mc_dat), .ain(mc_ack), .ic_seq({\ci_seq[1] , 
        \ci_seq[0] }), .ic_pred({\ci_pred[1] , \ci_pred[0] }), .ic_size({
        \ci_size[3] , \ci_size[2] , \ci_size[1] , \ci_size[0] }), .ic_itag({
        \ci_itag[9] , \ci_itag[8] , \ci_itag[7] , \ci_itag[6] , \ci_itag[5] , 
        \ci_itag[4] , \ci_itag[3] , \ci_itag[2] , \ci_itag[1] , \ci_itag[0] }), 
        .ic_wd({\ci_wd[63] , \ci_wd[62] , \ci_wd[61] , \ci_wd[60] , 
        \ci_wd[59] , \ci_wd[58] , \ci_wd[57] , \ci_wd[56] , \ci_wd[55] , 
        \ci_wd[54] , \ci_wd[53] , \ci_wd[52] , \ci_wd[51] , \ci_wd[50] , 
        \ci_wd[49] , \ci_wd[48] , \ci_wd[47] , \ci_wd[46] , \ci_wd[45] , 
        \ci_wd[44] , \ci_wd[43] , \ci_wd[42] , \ci_wd[41] , \ci_wd[40] , 
        \ci_wd[39] , \ci_wd[38] , \ci_wd[37] , \ci_wd[36] , \ci_wd[35] , 
        \ci_wd[34] , \ci_wd[33] , \ci_wd[32] , \ci_wd[31] , \ci_wd[30] , 
        \ci_wd[29] , \ci_wd[28] , \ci_wd[27] , \ci_wd[26] , \ci_wd[25] , 
        \ci_wd[24] , \ci_wd[23] , \ci_wd[22] , \ci_wd[21] , \ci_wd[20] , 
        \ci_wd[19] , \ci_wd[18] , \ci_wd[17] , \ci_wd[16] , \ci_wd[15] , 
        \ci_wd[14] , \ci_wd[13] , \ci_wd[12] , \ci_wd[11] , \ci_wd[10] , 
        \ci_wd[9] , \ci_wd[8] , \ci_wd[7] , \ci_wd[6] , \ci_wd[5] , \ci_wd[4] , 
        \ci_wd[3] , \ci_wd[2] , \ci_wd[1] , \ci_wd[0] }), .ic_lock({
        \ci_lock[1] , \ci_lock[0] }), .ic_a({\ci_a[63] , \ci_a[62] , 
        \ci_a[61] , \ci_a[60] , \ci_a[59] , \ci_a[58] , \ci_a[57] , \ci_a[56] , 
        \ci_a[55] , \ci_a[54] , \ci_a[53] , \ci_a[52] , \ci_a[51] , \ci_a[50] , 
        \ci_a[49] , \ci_a[48] , \ci_a[47] , \ci_a[46] , \ci_a[45] , \ci_a[44] , 
        \ci_a[43] , \ci_a[42] , \ci_a[41] , \ci_a[40] , \ci_a[39] , \ci_a[38] , 
        \ci_a[37] , \ci_a[36] , \ci_a[35] , \ci_a[34] , \ci_a[33] , \ci_a[32] , 
        \ci_a[31] , \ci_a[30] , \ci_a[29] , \ci_a[28] , \ci_a[27] , \ci_a[26] , 
        \ci_a[25] , \ci_a[24] , \ci_a[23] , \ci_a[22] , \ci_a[21] , \ci_a[20] , 
        \ci_a[19] , \ci_a[18] , \ci_a[17] , \ci_a[16] , \ci_a[15] , \ci_a[14] , 
        \ci_a[13] , \ci_a[12] , \ci_a[11] , \ci_a[10] , \ci_a[9] , \ci_a[8] , 
        \ci_a[7] , \ci_a[6] , \ci_a[5] , \ci_a[4] , \ci_a[3] , \ci_a[2] , 
        \ci_a[1] , \ci_a[0] }), .ic_rnw({\ci_rnw[1] , \ci_rnw[0] }), .ic_col({
        \ci_col[5] , \ci_col[4] , \ci_col[3] , \ci_col[2] , \ci_col[1] , 
        \ci_col[0] }), .ic_ack(ci_ack), .req_out(mr_req), .we_i(mr_we), 
        .err_i(mr_err), .dat_i(mr_dat), .aout(mr_ack), .ir_rd({\ri_rd[63] , 
        \ri_rd[62] , \ri_rd[61] , \ri_rd[60] , \ri_rd[59] , \ri_rd[58] , 
        \ri_rd[57] , \ri_rd[56] , \ri_rd[55] , \ri_rd[54] , \ri_rd[53] , 
        \ri_rd[52] , \ri_rd[51] , \ri_rd[50] , \ri_rd[49] , \ri_rd[48] , 
        \ri_rd[47] , \ri_rd[46] , \ri_rd[45] , \ri_rd[44] , \ri_rd[43] , 
        \ri_rd[42] , \ri_rd[41] , \ri_rd[40] , \ri_rd[39] , \ri_rd[38] , 
        \ri_rd[37] , \ri_rd[36] , \ri_rd[35] , \ri_rd[34] , \ri_rd[33] , 
        \ri_rd[32] , \ri_rd[31] , \ri_rd[30] , \ri_rd[29] , \ri_rd[28] , 
        \ri_rd[27] , \ri_rd[26] , \ri_rd[25] , \ri_rd[24] , \ri_rd[23] , 
        \ri_rd[22] , \ri_rd[21] , \ri_rd[20] , \ri_rd[19] , \ri_rd[18] , 
        \ri_rd[17] , \ri_rd[16] , \ri_rd[15] , \ri_rd[14] , \ri_rd[13] , 
        \ri_rd[12] , \ri_rd[11] , \ri_rd[10] , \ri_rd[9] , \ri_rd[8] , 
        \ri_rd[7] , \ri_rd[6] , \ri_rd[5] , \ri_rd[4] , \ri_rd[3] , \ri_rd[2] , 
        \ri_rd[1] , \ri_rd[0] }), .ir_err({\ri_err[1] , \ri_err[0] }), 
        .ir_rnw({\ri_rnw[1] , \ri_rnw[0] }), .ir_ack(ri_ack), .tag_id(tag_id), 
        .reset(reset) );
    i_adec_iport dec ( .e_h({SYNOPSYS_UNCONNECTED_1, \i_eh[2] , \i_eh[1] , 
        \i_eh[0] }), .e_l({\i_el[3] , \i_el[2] , \i_el[1] , \i_el[0] }), .r_h(
        {\i_rh[3] , \i_rh[2] , \i_rh[1] , SYNOPSYS_UNCONNECTED_2}), .r_l({
        \i_rl[3] , \i_rl[2] , \i_rl[1] , \i_rl[0] }), .ah({\ci_a[63] , 
        \ci_a[62] , \ci_a[61] , \ci_a[60] , \ci_a[59] , \ci_a[58] , \ci_a[57] , 
        \ci_a[56] , \ci_a[55] , \ci_a[54] , \ci_a[53] , \ci_a[52] , \ci_a[51] , 
        \ci_a[50] , \ci_a[49] , \ci_a[48] , \ci_a[47] , \ci_a[46] , \ci_a[45] , 
        \ci_a[44] , \ci_a[43] , \ci_a[42] , \ci_a[41] , \ci_a[40] , \ci_a[39] , 
        \ci_a[38] , \ci_a[37] , \ci_a[36] , \ci_a[35] , \ci_a[34] , \ci_a[33] , 
        \ci_a[32] }), .al({\ci_a[31] , \ci_a[30] , \ci_a[29] , \ci_a[28] , 
        \ci_a[27] , \ci_a[26] , \ci_a[25] , \ci_a[24] , \ci_a[23] , \ci_a[22] , 
        \ci_a[21] , \ci_a[20] , \ci_a[19] , \ci_a[18] , \ci_a[17] , \ci_a[16] , 
        \ci_a[15] , \ci_a[14] , \ci_a[13] , \ci_a[12] , \ci_a[11] , \ci_a[10] , 
        \ci_a[9] , \ci_a[8] , \ci_a[7] , \ci_a[6] , \ci_a[5] , \ci_a[4] , 
        \ci_a[3] , \ci_a[2] , \ci_a[1] , \ci_a[0] }), .e_bare(e_bare), .e_dm(
        e_dm), .e_im(e_im), .e_wish(e_wish), .r_bare(r_bare), .r_dm(r_dm), 
        .r_im(r_im), .r_wish(r_wish), .force_bare(force_bare) );
    route_tx_iport rt ( .o({\route[4] , SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4, \route[1] , \route[0] }), .rtxack(routetx_ack), 
        .e_h({1'b0, \i_eh[2] , \i_eh[1] , \i_eh[0] }), .e_l({\i_el[3] , 
        \i_el[2] , \i_el[1] , \i_el[0] }), .noa(nroute_ack), .r_h({\i_rh[3] , 
        \i_rh[2] , \i_rh[1] , 1'b0}), .r_l({\i_rl[3] , \i_rl[2] , \i_rl[1] , 
        \i_rl[0] }), .rtxreq(routetx_req) );
    initiator_iport it ( .cack(ci_ack), .chaincommand(chaincommand), .err({
        \ri_err[1] , \ri_err[0] }), .nchainresponseack(nchainresponseack), 
        .nrouteack(nroute_ack), .rd({\ri_rd[63] , \ri_rd[62] , \ri_rd[61] , 
        \ri_rd[60] , \ri_rd[59] , \ri_rd[58] , \ri_rd[57] , \ri_rd[56] , 
        \ri_rd[55] , \ri_rd[54] , \ri_rd[53] , \ri_rd[52] , \ri_rd[51] , 
        \ri_rd[50] , \ri_rd[49] , \ri_rd[48] , \ri_rd[47] , \ri_rd[46] , 
        \ri_rd[45] , \ri_rd[44] , \ri_rd[43] , \ri_rd[42] , \ri_rd[41] , 
        \ri_rd[40] , \ri_rd[39] , \ri_rd[38] , \ri_rd[37] , \ri_rd[36] , 
        \ri_rd[35] , \ri_rd[34] , \ri_rd[33] , \ri_rd[32] , \ri_rd[31] , 
        \ri_rd[30] , \ri_rd[29] , \ri_rd[28] , \ri_rd[27] , \ri_rd[26] , 
        \ri_rd[25] , \ri_rd[24] , \ri_rd[23] , \ri_rd[22] , \ri_rd[21] , 
        \ri_rd[20] , \ri_rd[19] , \ri_rd[18] , \ri_rd[17] , \ri_rd[16] , 
        \ri_rd[15] , \ri_rd[14] , \ri_rd[13] , \ri_rd[12] , \ri_rd[11] , 
        \ri_rd[10] , \ri_rd[9] , \ri_rd[8] , \ri_rd[7] , \ri_rd[6] , 
        \ri_rd[5] , \ri_rd[4] , \ri_rd[3] , \ri_rd[2] , \ri_rd[1] , \ri_rd[0] 
        }), .routetxreq(routetx_req), .rrnw({\ri_rnw[1] , \ri_rnw[0] }), .a({
        \ci_a[63] , \ci_a[62] , \ci_a[61] , \ci_a[60] , \ci_a[59] , \ci_a[58] , 
        \ci_a[57] , \ci_a[56] , \ci_a[55] , \ci_a[54] , \ci_a[53] , \ci_a[52] , 
        \ci_a[51] , \ci_a[50] , \ci_a[49] , \ci_a[48] , \ci_a[47] , \ci_a[46] , 
        \ci_a[45] , \ci_a[44] , \ci_a[43] , \ci_a[42] , \ci_a[41] , \ci_a[40] , 
        \ci_a[39] , \ci_a[38] , \ci_a[37] , \ci_a[36] , \ci_a[35] , \ci_a[34] , 
        \ci_a[33] , \ci_a[32] , \ci_a[31] , \ci_a[30] , \ci_a[29] , \ci_a[28] , 
        \ci_a[27] , \ci_a[26] , \ci_a[25] , \ci_a[24] , \ci_a[23] , \ci_a[22] , 
        \ci_a[21] , \ci_a[20] , \ci_a[19] , \ci_a[18] , \ci_a[17] , \ci_a[16] , 
        \ci_a[15] , \ci_a[14] , \ci_a[13] , \ci_a[12] , \ci_a[11] , \ci_a[10] , 
        \ci_a[9] , \ci_a[8] , \ci_a[7] , \ci_a[6] , \ci_a[5] , \ci_a[4] , 
        \ci_a[3] , \ci_a[2] , \ci_a[1] , \ci_a[0] }), .chainresponse(
        chainresponse), .col({\ci_col[5] , \ci_col[4] , \ci_col[3] , 
        \ci_col[2] , \ci_col[1] , \ci_col[0] }), .crnw({\ci_rnw[1] , 
        \ci_rnw[0] }), .itag({\ci_itag[9] , \ci_itag[8] , \ci_itag[7] , 
        \ci_itag[6] , \ci_itag[5] , \ci_itag[4] , \ci_itag[3] , \ci_itag[2] , 
        \ci_itag[1] , \ci_itag[0] }), .lock({\ci_lock[1] , \ci_lock[0] }), 
        .nReset(nReset), .nchaincommandack(nchaincommandack), .pred({
        \ci_pred[1] , \ci_pred[0] }), .rack(ri_ack), .route({\route[4] , 1'b0, 
        1'b0, \route[1] , \route[0] }), .routetxack(routetx_ack), .seq({
        \ci_seq[1] , \ci_seq[0] }), .size({\ci_size[3] , \ci_size[2] , 
        \ci_size[1] , \ci_size[0] }), .wd({\ci_wd[63] , \ci_wd[62] , 
        \ci_wd[61] , \ci_wd[60] , \ci_wd[59] , \ci_wd[58] , \ci_wd[57] , 
        \ci_wd[56] , \ci_wd[55] , \ci_wd[54] , \ci_wd[53] , \ci_wd[52] , 
        \ci_wd[51] , \ci_wd[50] , \ci_wd[49] , \ci_wd[48] , \ci_wd[47] , 
        \ci_wd[46] , \ci_wd[45] , \ci_wd[44] , \ci_wd[43] , \ci_wd[42] , 
        \ci_wd[41] , \ci_wd[40] , \ci_wd[39] , \ci_wd[38] , \ci_wd[37] , 
        \ci_wd[36] , \ci_wd[35] , \ci_wd[34] , \ci_wd[33] , \ci_wd[32] , 
        \ci_wd[31] , \ci_wd[30] , \ci_wd[29] , \ci_wd[28] , \ci_wd[27] , 
        \ci_wd[26] , \ci_wd[25] , \ci_wd[24] , \ci_wd[23] , \ci_wd[22] , 
        \ci_wd[21] , \ci_wd[20] , \ci_wd[19] , \ci_wd[18] , \ci_wd[17] , 
        \ci_wd[16] , \ci_wd[15] , \ci_wd[14] , \ci_wd[13] , \ci_wd[12] , 
        \ci_wd[11] , \ci_wd[10] , \ci_wd[9] , \ci_wd[8] , \ci_wd[7] , 
        \ci_wd[6] , \ci_wd[5] , \ci_wd[4] , \ci_wd[3] , \ci_wd[2] , \ci_wd[1] , 
        \ci_wd[0] }) );
endmodule


module matched_delay_m2cp_com_dport ( x, a );
input  a;
output x;
    wire n2;
    buf_1 I1 ( .x(n2), .a(a) );
    buf_16 U1 ( .x(x), .a(n2) );
endmodule


module sr2dr_word_3 ( i, req, h, l );
input  [31:0] i;
output [31:0] h;
output [31:0] l;
input  req;
    wire \U31/ni , \U31/nh , \U31/nl , n9, n1, n2, \U30/ni , \U30/nh , 
        \U30/nl , n8, \U29/ni , \U29/nh , \U29/nl , \U28/ni , \U28/nh , 
        \U28/nl , \U27/ni , \U27/nh , \U27/nl , \U26/ni , \U26/nh , \U26/nl , 
        n7, n4, \U25/ni , \U25/nh , \U25/nl , \U24/ni , \U24/nh , \U24/nl , 
        \U23/ni , \U23/nh , \U23/nl , n3, \U22/ni , \U22/nh , \U22/nl , n6, 
        \U21/ni , \U21/nh , \U21/nl , \U20/ni , \U20/nh , \U20/nl , n5, 
        \U19/ni , \U19/nh , \U19/nl , \U18/ni , \U18/nh , \U18/nl , \U17/ni , 
        \U17/nh , \U17/nl , \U16/ni , \U16/nh , \U16/nl , \U15/ni , \U15/nh , 
        \U15/nl , \U14/ni , \U14/nh , \U14/nl , \U13/ni , \U13/nh , \U13/nl , 
        \U12/ni , \U12/nh , \U12/nl , \U11/ni , \U11/nh , \U11/nl , \U10/ni , 
        \U10/nh , \U10/nl , \U9/ni , \U9/nh , \U9/nl , \U8/ni , \U8/nh , 
        \U8/nl , \U7/ni , \U7/nh , \U7/nl , \U6/ni , \U6/nh , \U6/nl , \U5/ni , 
        \U5/nh , \U5/nl , \U4/ni , \U4/nh , \U4/nl , \U3/ni , \U3/nh , \U3/nl , 
        \U2/ni , \U2/nh , \U2/nl , \U1/ni , \U1/nh , \U1/nl , \U0/ni , \U0/nh , 
        \U0/nl , n12, n11, n10;
    inv_1 \U31/Uii  ( .x(\U31/ni ), .a(i[31]) );
    inv_1 \U31/Uih  ( .x(\U31/nh ), .a(h[31]) );
    inv_1 \U31/Uil  ( .x(\U31/nl ), .a(l[31]) );
    ao23_1 \U31/Ucl/U1/U1  ( .x(l[31]), .a(n9), .b(l[31]), .c(n1), .d(\U31/ni 
        ), .e(\U31/nh ) );
    ao23_1 \U31/Uch/U1/U1  ( .x(h[31]), .a(n9), .b(h[31]), .c(n2), .d(i[31]), 
        .e(\U31/nl ) );
    inv_1 \U30/Uii  ( .x(\U30/ni ), .a(i[30]) );
    inv_1 \U30/Uih  ( .x(\U30/nh ), .a(h[30]) );
    inv_1 \U30/Uil  ( .x(\U30/nl ), .a(l[30]) );
    ao23_1 \U30/Ucl/U1/U1  ( .x(l[30]), .a(n8), .b(l[30]), .c(n1), .d(\U30/ni 
        ), .e(\U30/nh ) );
    ao23_1 \U30/Uch/U1/U1  ( .x(h[30]), .a(n8), .b(h[30]), .c(n1), .d(i[30]), 
        .e(\U30/nl ) );
    inv_1 \U29/Uii  ( .x(\U29/ni ), .a(i[29]) );
    inv_1 \U29/Uih  ( .x(\U29/nh ), .a(h[29]) );
    inv_1 \U29/Uil  ( .x(\U29/nl ), .a(l[29]) );
    ao23_1 \U29/Ucl/U1/U1  ( .x(l[29]), .a(n8), .b(l[29]), .c(n1), .d(\U29/ni 
        ), .e(\U29/nh ) );
    ao23_1 \U29/Uch/U1/U1  ( .x(h[29]), .a(n8), .b(h[29]), .c(n2), .d(i[29]), 
        .e(\U29/nl ) );
    inv_1 \U28/Uii  ( .x(\U28/ni ), .a(i[28]) );
    inv_1 \U28/Uih  ( .x(\U28/nh ), .a(h[28]) );
    inv_1 \U28/Uil  ( .x(\U28/nl ), .a(l[28]) );
    ao23_1 \U28/Ucl/U1/U1  ( .x(l[28]), .a(n8), .b(l[28]), .c(n2), .d(\U28/ni 
        ), .e(\U28/nh ) );
    ao23_1 \U28/Uch/U1/U1  ( .x(h[28]), .a(n8), .b(h[28]), .c(n2), .d(i[28]), 
        .e(\U28/nl ) );
    inv_1 \U27/Uii  ( .x(\U27/ni ), .a(i[27]) );
    inv_1 \U27/Uih  ( .x(\U27/nh ), .a(h[27]) );
    inv_1 \U27/Uil  ( .x(\U27/nl ), .a(l[27]) );
    ao23_1 \U27/Ucl/U1/U1  ( .x(l[27]), .a(n8), .b(l[27]), .c(n2), .d(\U27/ni 
        ), .e(\U27/nh ) );
    ao23_1 \U27/Uch/U1/U1  ( .x(h[27]), .a(n8), .b(h[27]), .c(n2), .d(i[27]), 
        .e(\U27/nl ) );
    inv_1 \U26/Uii  ( .x(\U26/ni ), .a(i[26]) );
    inv_1 \U26/Uih  ( .x(\U26/nh ), .a(h[26]) );
    inv_1 \U26/Uil  ( .x(\U26/nl ), .a(l[26]) );
    ao23_1 \U26/Ucl/U1/U1  ( .x(l[26]), .a(n7), .b(l[26]), .c(n2), .d(\U26/ni 
        ), .e(\U26/nh ) );
    ao23_1 \U26/Uch/U1/U1  ( .x(h[26]), .a(n7), .b(h[26]), .c(n4), .d(i[26]), 
        .e(\U26/nl ) );
    inv_1 \U25/Uii  ( .x(\U25/ni ), .a(i[25]) );
    inv_1 \U25/Uih  ( .x(\U25/nh ), .a(h[25]) );
    inv_1 \U25/Uil  ( .x(\U25/nl ), .a(l[25]) );
    ao23_1 \U25/Ucl/U1/U1  ( .x(l[25]), .a(n7), .b(l[25]), .c(n4), .d(\U25/ni 
        ), .e(\U25/nh ) );
    ao23_1 \U25/Uch/U1/U1  ( .x(h[25]), .a(n7), .b(h[25]), .c(n4), .d(i[25]), 
        .e(\U25/nl ) );
    inv_1 \U24/Uii  ( .x(\U24/ni ), .a(i[24]) );
    inv_1 \U24/Uih  ( .x(\U24/nh ), .a(h[24]) );
    inv_1 \U24/Uil  ( .x(\U24/nl ), .a(l[24]) );
    ao23_1 \U24/Ucl/U1/U1  ( .x(l[24]), .a(n7), .b(l[24]), .c(n4), .d(\U24/ni 
        ), .e(\U24/nh ) );
    ao23_1 \U24/Uch/U1/U1  ( .x(h[24]), .a(n7), .b(h[24]), .c(n4), .d(i[24]), 
        .e(\U24/nl ) );
    inv_1 \U23/Uii  ( .x(\U23/ni ), .a(i[23]) );
    inv_1 \U23/Uih  ( .x(\U23/nh ), .a(h[23]) );
    inv_1 \U23/Uil  ( .x(\U23/nl ), .a(l[23]) );
    ao23_1 \U23/Ucl/U1/U1  ( .x(l[23]), .a(n7), .b(l[23]), .c(n3), .d(\U23/ni 
        ), .e(\U23/nh ) );
    ao23_1 \U23/Uch/U1/U1  ( .x(h[23]), .a(n7), .b(h[23]), .c(n3), .d(i[23]), 
        .e(\U23/nl ) );
    inv_1 \U22/Uii  ( .x(\U22/ni ), .a(i[22]) );
    inv_1 \U22/Uih  ( .x(\U22/nh ), .a(h[22]) );
    inv_1 \U22/Uil  ( .x(\U22/nl ), .a(l[22]) );
    ao23_1 \U22/Ucl/U1/U1  ( .x(l[22]), .a(n6), .b(l[22]), .c(n3), .d(\U22/ni 
        ), .e(\U22/nh ) );
    ao23_1 \U22/Uch/U1/U1  ( .x(h[22]), .a(n6), .b(h[22]), .c(n3), .d(i[22]), 
        .e(\U22/nl ) );
    inv_1 \U21/Uii  ( .x(\U21/ni ), .a(i[21]) );
    inv_1 \U21/Uih  ( .x(\U21/nh ), .a(h[21]) );
    inv_1 \U21/Uil  ( .x(\U21/nl ), .a(l[21]) );
    ao23_1 \U21/Ucl/U1/U1  ( .x(l[21]), .a(n6), .b(l[21]), .c(n3), .d(\U21/ni 
        ), .e(\U21/nh ) );
    ao23_1 \U21/Uch/U1/U1  ( .x(h[21]), .a(n6), .b(h[21]), .c(n3), .d(i[21]), 
        .e(\U21/nl ) );
    inv_1 \U20/Uii  ( .x(\U20/ni ), .a(i[20]) );
    inv_1 \U20/Uih  ( .x(\U20/nh ), .a(h[20]) );
    inv_1 \U20/Uil  ( .x(\U20/nl ), .a(l[20]) );
    ao23_1 \U20/Ucl/U1/U1  ( .x(l[20]), .a(n6), .b(l[20]), .c(n5), .d(\U20/ni 
        ), .e(\U20/nh ) );
    ao23_1 \U20/Uch/U1/U1  ( .x(h[20]), .a(n6), .b(h[20]), .c(n4), .d(i[20]), 
        .e(\U20/nl ) );
    inv_1 \U19/Uii  ( .x(\U19/ni ), .a(i[19]) );
    inv_1 \U19/Uih  ( .x(\U19/nh ), .a(h[19]) );
    inv_1 \U19/Uil  ( .x(\U19/nl ), .a(l[19]) );
    ao23_1 \U19/Ucl/U1/U1  ( .x(l[19]), .a(n6), .b(l[19]), .c(n4), .d(\U19/ni 
        ), .e(\U19/nh ) );
    ao23_1 \U19/Uch/U1/U1  ( .x(h[19]), .a(n6), .b(h[19]), .c(n4), .d(i[19]), 
        .e(\U19/nl ) );
    inv_1 \U18/Uii  ( .x(\U18/ni ), .a(i[18]) );
    inv_1 \U18/Uih  ( .x(\U18/nh ), .a(h[18]) );
    inv_1 \U18/Uil  ( .x(\U18/nl ), .a(l[18]) );
    ao23_1 \U18/Ucl/U1/U1  ( .x(l[18]), .a(n5), .b(l[18]), .c(n5), .d(\U18/ni 
        ), .e(\U18/nh ) );
    ao23_1 \U18/Uch/U1/U1  ( .x(h[18]), .a(n5), .b(h[18]), .c(n5), .d(i[18]), 
        .e(\U18/nl ) );
    inv_1 \U17/Uii  ( .x(\U17/ni ), .a(i[17]) );
    inv_1 \U17/Uih  ( .x(\U17/nh ), .a(h[17]) );
    inv_1 \U17/Uil  ( .x(\U17/nl ), .a(l[17]) );
    ao23_1 \U17/Ucl/U1/U1  ( .x(l[17]), .a(n6), .b(l[17]), .c(n5), .d(\U17/ni 
        ), .e(\U17/nh ) );
    ao23_1 \U17/Uch/U1/U1  ( .x(h[17]), .a(n7), .b(h[17]), .c(n4), .d(i[17]), 
        .e(\U17/nl ) );
    inv_1 \U16/Uii  ( .x(\U16/ni ), .a(i[16]) );
    inv_1 \U16/Uih  ( .x(\U16/nh ), .a(h[16]) );
    inv_1 \U16/Uil  ( .x(\U16/nl ), .a(l[16]) );
    ao23_1 \U16/Ucl/U1/U1  ( .x(l[16]), .a(n9), .b(l[16]), .c(n3), .d(\U16/ni 
        ), .e(\U16/nh ) );
    ao23_1 \U16/Uch/U1/U1  ( .x(h[16]), .a(n9), .b(h[16]), .c(n1), .d(i[16]), 
        .e(\U16/nl ) );
    inv_1 \U15/Uii  ( .x(\U15/ni ), .a(i[15]) );
    inv_1 \U15/Uih  ( .x(\U15/nh ), .a(h[15]) );
    inv_1 \U15/Uil  ( .x(\U15/nl ), .a(l[15]) );
    ao23_1 \U15/Ucl/U1/U1  ( .x(l[15]), .a(n8), .b(l[15]), .c(n1), .d(\U15/ni 
        ), .e(\U15/nh ) );
    ao23_1 \U15/Uch/U1/U1  ( .x(h[15]), .a(n7), .b(h[15]), .c(n1), .d(i[15]), 
        .e(\U15/nl ) );
    inv_1 \U14/Uii  ( .x(\U14/ni ), .a(i[14]) );
    inv_1 \U14/Uih  ( .x(\U14/nh ), .a(h[14]) );
    inv_1 \U14/Uil  ( .x(\U14/nl ), .a(l[14]) );
    ao23_1 \U14/Ucl/U1/U1  ( .x(l[14]), .a(n6), .b(l[14]), .c(n1), .d(\U14/ni 
        ), .e(\U14/nh ) );
    ao23_1 \U14/Uch/U1/U1  ( .x(h[14]), .a(n6), .b(h[14]), .c(n3), .d(i[14]), 
        .e(\U14/nl ) );
    inv_1 \U13/Uii  ( .x(\U13/ni ), .a(i[13]) );
    inv_1 \U13/Uih  ( .x(\U13/nh ), .a(h[13]) );
    inv_1 \U13/Uil  ( .x(\U13/nl ), .a(l[13]) );
    ao23_1 \U13/Ucl/U1/U1  ( .x(l[13]), .a(n6), .b(l[13]), .c(n4), .d(\U13/ni 
        ), .e(\U13/nh ) );
    ao23_1 \U13/Uch/U1/U1  ( .x(h[13]), .a(n6), .b(h[13]), .c(n4), .d(i[13]), 
        .e(\U13/nl ) );
    inv_1 \U12/Uii  ( .x(\U12/ni ), .a(i[12]) );
    inv_1 \U12/Uih  ( .x(\U12/nh ), .a(h[12]) );
    inv_1 \U12/Uil  ( .x(\U12/nl ), .a(l[12]) );
    ao23_1 \U12/Ucl/U1/U1  ( .x(l[12]), .a(n5), .b(l[12]), .c(n4), .d(\U12/ni 
        ), .e(\U12/nh ) );
    ao23_1 \U12/Uch/U1/U1  ( .x(h[12]), .a(n5), .b(h[12]), .c(n4), .d(i[12]), 
        .e(\U12/nl ) );
    inv_1 \U11/Uii  ( .x(\U11/ni ), .a(i[11]) );
    inv_1 \U11/Uih  ( .x(\U11/nh ), .a(h[11]) );
    inv_1 \U11/Uil  ( .x(\U11/nl ), .a(l[11]) );
    ao23_1 \U11/Ucl/U1/U1  ( .x(l[11]), .a(n5), .b(l[11]), .c(n4), .d(\U11/ni 
        ), .e(\U11/nh ) );
    ao23_1 \U11/Uch/U1/U1  ( .x(h[11]), .a(n5), .b(h[11]), .c(n4), .d(i[11]), 
        .e(\U11/nl ) );
    inv_1 \U10/Uii  ( .x(\U10/ni ), .a(i[10]) );
    inv_1 \U10/Uih  ( .x(\U10/nh ), .a(h[10]) );
    inv_1 \U10/Uil  ( .x(\U10/nl ), .a(l[10]) );
    ao23_1 \U10/Ucl/U1/U1  ( .x(l[10]), .a(n5), .b(l[10]), .c(n3), .d(\U10/ni 
        ), .e(\U10/nh ) );
    ao23_1 \U10/Uch/U1/U1  ( .x(h[10]), .a(n5), .b(h[10]), .c(n3), .d(i[10]), 
        .e(\U10/nl ) );
    inv_1 \U9/Uii  ( .x(\U9/ni ), .a(i[9]) );
    inv_1 \U9/Uih  ( .x(\U9/nh ), .a(h[9]) );
    inv_1 \U9/Uil  ( .x(\U9/nl ), .a(l[9]) );
    ao23_1 \U9/Ucl/U1/U1  ( .x(l[9]), .a(n5), .b(l[9]), .c(n3), .d(\U9/ni ), 
        .e(\U9/nh ) );
    ao23_1 \U9/Uch/U1/U1  ( .x(h[9]), .a(n5), .b(h[9]), .c(n3), .d(i[9]), .e(
        \U9/nl ) );
    inv_1 \U8/Uii  ( .x(\U8/ni ), .a(i[8]) );
    inv_1 \U8/Uih  ( .x(\U8/nh ), .a(h[8]) );
    inv_1 \U8/Uil  ( .x(\U8/nl ), .a(l[8]) );
    ao23_1 \U8/Ucl/U1/U1  ( .x(l[8]), .a(n5), .b(l[8]), .c(n3), .d(\U8/ni ), 
        .e(\U8/nh ) );
    ao23_1 \U8/Uch/U1/U1  ( .x(h[8]), .a(n5), .b(h[8]), .c(n3), .d(i[8]), .e(
        \U8/nl ) );
    inv_1 \U7/Uii  ( .x(\U7/ni ), .a(i[7]) );
    inv_1 \U7/Uih  ( .x(\U7/nh ), .a(h[7]) );
    inv_1 \U7/Uil  ( .x(\U7/nl ), .a(l[7]) );
    ao23_1 \U7/Ucl/U1/U1  ( .x(l[7]), .a(n7), .b(l[7]), .c(n3), .d(\U7/ni ), 
        .e(\U7/nh ) );
    ao23_1 \U7/Uch/U1/U1  ( .x(h[7]), .a(n7), .b(h[7]), .c(n2), .d(i[7]), .e(
        \U7/nl ) );
    inv_1 \U6/Uii  ( .x(\U6/ni ), .a(i[6]) );
    inv_1 \U6/Uih  ( .x(\U6/nh ), .a(h[6]) );
    inv_1 \U6/Uil  ( .x(\U6/nl ), .a(l[6]) );
    ao23_1 \U6/Ucl/U1/U1  ( .x(l[6]), .a(n7), .b(l[6]), .c(n2), .d(\U6/ni ), 
        .e(\U6/nh ) );
    ao23_1 \U6/Uch/U1/U1  ( .x(h[6]), .a(n7), .b(h[6]), .c(n2), .d(i[6]), .e(
        \U6/nl ) );
    inv_1 \U5/Uii  ( .x(\U5/ni ), .a(i[5]) );
    inv_1 \U5/Uih  ( .x(\U5/nh ), .a(h[5]) );
    inv_1 \U5/Uil  ( .x(\U5/nl ), .a(l[5]) );
    ao23_1 \U5/Ucl/U1/U1  ( .x(l[5]), .a(n7), .b(l[5]), .c(n2), .d(\U5/ni ), 
        .e(\U5/nh ) );
    ao23_1 \U5/Uch/U1/U1  ( .x(h[5]), .a(n7), .b(h[5]), .c(n2), .d(i[5]), .e(
        \U5/nl ) );
    inv_1 \U4/Uii  ( .x(\U4/ni ), .a(i[4]) );
    inv_1 \U4/Uih  ( .x(\U4/nh ), .a(h[4]) );
    inv_1 \U4/Uil  ( .x(\U4/nl ), .a(l[4]) );
    ao23_1 \U4/Ucl/U1/U1  ( .x(l[4]), .a(n6), .b(l[4]), .c(n2), .d(\U4/ni ), 
        .e(\U4/nh ) );
    ao23_1 \U4/Uch/U1/U1  ( .x(h[4]), .a(n6), .b(h[4]), .c(n2), .d(i[4]), .e(
        \U4/nl ) );
    inv_1 \U3/Uii  ( .x(\U3/ni ), .a(i[3]) );
    inv_1 \U3/Uih  ( .x(\U3/nh ), .a(h[3]) );
    inv_1 \U3/Uil  ( .x(\U3/nl ), .a(l[3]) );
    ao23_1 \U3/Ucl/U1/U1  ( .x(l[3]), .a(n6), .b(l[3]), .c(n2), .d(\U3/ni ), 
        .e(\U3/nh ) );
    ao23_1 \U3/Uch/U1/U1  ( .x(h[3]), .a(n8), .b(h[3]), .c(n1), .d(i[3]), .e(
        \U3/nl ) );
    inv_1 \U2/Uii  ( .x(\U2/ni ), .a(i[2]) );
    inv_1 \U2/Uih  ( .x(\U2/nh ), .a(h[2]) );
    inv_1 \U2/Uil  ( .x(\U2/nl ), .a(l[2]) );
    ao23_1 \U2/Ucl/U1/U1  ( .x(l[2]), .a(n8), .b(l[2]), .c(n1), .d(\U2/ni ), 
        .e(\U2/nh ) );
    ao23_1 \U2/Uch/U1/U1  ( .x(h[2]), .a(n8), .b(h[2]), .c(n1), .d(i[2]), .e(
        \U2/nl ) );
    inv_1 \U1/Uii  ( .x(\U1/ni ), .a(i[1]) );
    inv_1 \U1/Uih  ( .x(\U1/nh ), .a(h[1]) );
    inv_1 \U1/Uil  ( .x(\U1/nl ), .a(l[1]) );
    ao23_1 \U1/Ucl/U1/U1  ( .x(l[1]), .a(n8), .b(l[1]), .c(n1), .d(\U1/ni ), 
        .e(\U1/nh ) );
    ao23_1 \U1/Uch/U1/U1  ( .x(h[1]), .a(n8), .b(h[1]), .c(n1), .d(i[1]), .e(
        \U1/nl ) );
    inv_1 \U0/Uii  ( .x(\U0/ni ), .a(i[0]) );
    inv_1 \U0/Uih  ( .x(\U0/nh ), .a(h[0]) );
    inv_1 \U0/Uil  ( .x(\U0/nl ), .a(l[0]) );
    ao23_1 \U0/Ucl/U1/U1  ( .x(l[0]), .a(n8), .b(l[0]), .c(n1), .d(\U0/ni ), 
        .e(\U0/nh ) );
    ao23_1 \U0/Uch/U1/U1  ( .x(h[0]), .a(n8), .b(h[0]), .c(n1), .d(i[0]), .e(
        \U0/nl ) );
    buf_16 U1 ( .x(n1), .a(n12) );
    buf_16 U2 ( .x(n2), .a(n12) );
    buf_16 U3 ( .x(n3), .a(n12) );
    buf_16 U4 ( .x(n4), .a(n11) );
    buf_16 U5 ( .x(n5), .a(n11) );
    buf_16 U6 ( .x(n6), .a(n11) );
    buf_16 U7 ( .x(n7), .a(n10) );
    buf_16 U8 ( .x(n8), .a(n10) );
    buf_16 U9 ( .x(n9), .a(n10) );
    buf_16 U10 ( .x(n10), .a(req) );
    buf_16 U11 ( .x(n11), .a(req) );
    buf_16 U12 ( .x(n12), .a(req) );
endmodule


module sr2dr_word_2 ( i, req, h, l );
input  [31:0] i;
output [31:0] h;
output [31:0] l;
input  req;
    wire \U31/ni , \U31/nh , \U31/nl , n9, n1, n2, \U30/ni , \U30/nh , 
        \U30/nl , n8, \U29/ni , \U29/nh , \U29/nl , \U28/ni , \U28/nh , 
        \U28/nl , \U27/ni , \U27/nh , \U27/nl , \U26/ni , \U26/nh , \U26/nl , 
        n7, n4, \U25/ni , \U25/nh , \U25/nl , \U24/ni , \U24/nh , \U24/nl , 
        \U23/ni , \U23/nh , \U23/nl , n3, \U22/ni , \U22/nh , \U22/nl , n6, 
        \U21/ni , \U21/nh , \U21/nl , \U20/ni , \U20/nh , \U20/nl , n5, 
        \U19/ni , \U19/nh , \U19/nl , \U18/ni , \U18/nh , \U18/nl , \U17/ni , 
        \U17/nh , \U17/nl , \U16/ni , \U16/nh , \U16/nl , \U15/ni , \U15/nh , 
        \U15/nl , \U14/ni , \U14/nh , \U14/nl , \U13/ni , \U13/nh , \U13/nl , 
        \U12/ni , \U12/nh , \U12/nl , \U11/ni , \U11/nh , \U11/nl , \U10/ni , 
        \U10/nh , \U10/nl , \U9/ni , \U9/nh , \U9/nl , \U8/ni , \U8/nh , 
        \U8/nl , \U7/ni , \U7/nh , \U7/nl , \U6/ni , \U6/nh , \U6/nl , \U5/ni , 
        \U5/nh , \U5/nl , \U4/ni , \U4/nh , \U4/nl , \U3/ni , \U3/nh , \U3/nl , 
        \U2/ni , \U2/nh , \U2/nl , \U1/ni , \U1/nh , \U1/nl , \U0/ni , \U0/nh , 
        \U0/nl , n12, n11, n10;
    inv_1 \U31/Uii  ( .x(\U31/ni ), .a(i[31]) );
    inv_1 \U31/Uih  ( .x(\U31/nh ), .a(h[31]) );
    inv_1 \U31/Uil  ( .x(\U31/nl ), .a(l[31]) );
    ao23_1 \U31/Ucl/U1/U1  ( .x(l[31]), .a(n9), .b(l[31]), .c(n1), .d(\U31/ni 
        ), .e(\U31/nh ) );
    ao23_1 \U31/Uch/U1/U1  ( .x(h[31]), .a(n9), .b(h[31]), .c(n2), .d(i[31]), 
        .e(\U31/nl ) );
    inv_1 \U30/Uii  ( .x(\U30/ni ), .a(i[30]) );
    inv_1 \U30/Uih  ( .x(\U30/nh ), .a(h[30]) );
    inv_1 \U30/Uil  ( .x(\U30/nl ), .a(l[30]) );
    ao23_1 \U30/Ucl/U1/U1  ( .x(l[30]), .a(n8), .b(l[30]), .c(n1), .d(\U30/ni 
        ), .e(\U30/nh ) );
    ao23_1 \U30/Uch/U1/U1  ( .x(h[30]), .a(n8), .b(h[30]), .c(n1), .d(i[30]), 
        .e(\U30/nl ) );
    inv_1 \U29/Uii  ( .x(\U29/ni ), .a(i[29]) );
    inv_1 \U29/Uih  ( .x(\U29/nh ), .a(h[29]) );
    inv_1 \U29/Uil  ( .x(\U29/nl ), .a(l[29]) );
    ao23_1 \U29/Ucl/U1/U1  ( .x(l[29]), .a(n8), .b(l[29]), .c(n1), .d(\U29/ni 
        ), .e(\U29/nh ) );
    ao23_1 \U29/Uch/U1/U1  ( .x(h[29]), .a(n8), .b(h[29]), .c(n2), .d(i[29]), 
        .e(\U29/nl ) );
    inv_1 \U28/Uii  ( .x(\U28/ni ), .a(i[28]) );
    inv_1 \U28/Uih  ( .x(\U28/nh ), .a(h[28]) );
    inv_1 \U28/Uil  ( .x(\U28/nl ), .a(l[28]) );
    ao23_1 \U28/Ucl/U1/U1  ( .x(l[28]), .a(n8), .b(l[28]), .c(n2), .d(\U28/ni 
        ), .e(\U28/nh ) );
    ao23_1 \U28/Uch/U1/U1  ( .x(h[28]), .a(n8), .b(h[28]), .c(n2), .d(i[28]), 
        .e(\U28/nl ) );
    inv_1 \U27/Uii  ( .x(\U27/ni ), .a(i[27]) );
    inv_1 \U27/Uih  ( .x(\U27/nh ), .a(h[27]) );
    inv_1 \U27/Uil  ( .x(\U27/nl ), .a(l[27]) );
    ao23_1 \U27/Ucl/U1/U1  ( .x(l[27]), .a(n8), .b(l[27]), .c(n2), .d(\U27/ni 
        ), .e(\U27/nh ) );
    ao23_1 \U27/Uch/U1/U1  ( .x(h[27]), .a(n8), .b(h[27]), .c(n2), .d(i[27]), 
        .e(\U27/nl ) );
    inv_1 \U26/Uii  ( .x(\U26/ni ), .a(i[26]) );
    inv_1 \U26/Uih  ( .x(\U26/nh ), .a(h[26]) );
    inv_1 \U26/Uil  ( .x(\U26/nl ), .a(l[26]) );
    ao23_1 \U26/Ucl/U1/U1  ( .x(l[26]), .a(n7), .b(l[26]), .c(n2), .d(\U26/ni 
        ), .e(\U26/nh ) );
    ao23_1 \U26/Uch/U1/U1  ( .x(h[26]), .a(n7), .b(h[26]), .c(n4), .d(i[26]), 
        .e(\U26/nl ) );
    inv_1 \U25/Uii  ( .x(\U25/ni ), .a(i[25]) );
    inv_1 \U25/Uih  ( .x(\U25/nh ), .a(h[25]) );
    inv_1 \U25/Uil  ( .x(\U25/nl ), .a(l[25]) );
    ao23_1 \U25/Ucl/U1/U1  ( .x(l[25]), .a(n7), .b(l[25]), .c(n4), .d(\U25/ni 
        ), .e(\U25/nh ) );
    ao23_1 \U25/Uch/U1/U1  ( .x(h[25]), .a(n7), .b(h[25]), .c(n4), .d(i[25]), 
        .e(\U25/nl ) );
    inv_1 \U24/Uii  ( .x(\U24/ni ), .a(i[24]) );
    inv_1 \U24/Uih  ( .x(\U24/nh ), .a(h[24]) );
    inv_1 \U24/Uil  ( .x(\U24/nl ), .a(l[24]) );
    ao23_1 \U24/Ucl/U1/U1  ( .x(l[24]), .a(n7), .b(l[24]), .c(n4), .d(\U24/ni 
        ), .e(\U24/nh ) );
    ao23_1 \U24/Uch/U1/U1  ( .x(h[24]), .a(n7), .b(h[24]), .c(n4), .d(i[24]), 
        .e(\U24/nl ) );
    inv_1 \U23/Uii  ( .x(\U23/ni ), .a(i[23]) );
    inv_1 \U23/Uih  ( .x(\U23/nh ), .a(h[23]) );
    inv_1 \U23/Uil  ( .x(\U23/nl ), .a(l[23]) );
    ao23_1 \U23/Ucl/U1/U1  ( .x(l[23]), .a(n7), .b(l[23]), .c(n3), .d(\U23/ni 
        ), .e(\U23/nh ) );
    ao23_1 \U23/Uch/U1/U1  ( .x(h[23]), .a(n7), .b(h[23]), .c(n3), .d(i[23]), 
        .e(\U23/nl ) );
    inv_1 \U22/Uii  ( .x(\U22/ni ), .a(i[22]) );
    inv_1 \U22/Uih  ( .x(\U22/nh ), .a(h[22]) );
    inv_1 \U22/Uil  ( .x(\U22/nl ), .a(l[22]) );
    ao23_1 \U22/Ucl/U1/U1  ( .x(l[22]), .a(n6), .b(l[22]), .c(n3), .d(\U22/ni 
        ), .e(\U22/nh ) );
    ao23_1 \U22/Uch/U1/U1  ( .x(h[22]), .a(n6), .b(h[22]), .c(n3), .d(i[22]), 
        .e(\U22/nl ) );
    inv_1 \U21/Uii  ( .x(\U21/ni ), .a(i[21]) );
    inv_1 \U21/Uih  ( .x(\U21/nh ), .a(h[21]) );
    inv_1 \U21/Uil  ( .x(\U21/nl ), .a(l[21]) );
    ao23_1 \U21/Ucl/U1/U1  ( .x(l[21]), .a(n6), .b(l[21]), .c(n3), .d(\U21/ni 
        ), .e(\U21/nh ) );
    ao23_1 \U21/Uch/U1/U1  ( .x(h[21]), .a(n6), .b(h[21]), .c(n3), .d(i[21]), 
        .e(\U21/nl ) );
    inv_1 \U20/Uii  ( .x(\U20/ni ), .a(i[20]) );
    inv_1 \U20/Uih  ( .x(\U20/nh ), .a(h[20]) );
    inv_1 \U20/Uil  ( .x(\U20/nl ), .a(l[20]) );
    ao23_1 \U20/Ucl/U1/U1  ( .x(l[20]), .a(n6), .b(l[20]), .c(n5), .d(\U20/ni 
        ), .e(\U20/nh ) );
    ao23_1 \U20/Uch/U1/U1  ( .x(h[20]), .a(n6), .b(h[20]), .c(n4), .d(i[20]), 
        .e(\U20/nl ) );
    inv_1 \U19/Uii  ( .x(\U19/ni ), .a(i[19]) );
    inv_1 \U19/Uih  ( .x(\U19/nh ), .a(h[19]) );
    inv_1 \U19/Uil  ( .x(\U19/nl ), .a(l[19]) );
    ao23_1 \U19/Ucl/U1/U1  ( .x(l[19]), .a(n6), .b(l[19]), .c(n4), .d(\U19/ni 
        ), .e(\U19/nh ) );
    ao23_1 \U19/Uch/U1/U1  ( .x(h[19]), .a(n6), .b(h[19]), .c(n4), .d(i[19]), 
        .e(\U19/nl ) );
    inv_1 \U18/Uii  ( .x(\U18/ni ), .a(i[18]) );
    inv_1 \U18/Uih  ( .x(\U18/nh ), .a(h[18]) );
    inv_1 \U18/Uil  ( .x(\U18/nl ), .a(l[18]) );
    ao23_1 \U18/Ucl/U1/U1  ( .x(l[18]), .a(n5), .b(l[18]), .c(n5), .d(\U18/ni 
        ), .e(\U18/nh ) );
    ao23_1 \U18/Uch/U1/U1  ( .x(h[18]), .a(n5), .b(h[18]), .c(n5), .d(i[18]), 
        .e(\U18/nl ) );
    inv_1 \U17/Uii  ( .x(\U17/ni ), .a(i[17]) );
    inv_1 \U17/Uih  ( .x(\U17/nh ), .a(h[17]) );
    inv_1 \U17/Uil  ( .x(\U17/nl ), .a(l[17]) );
    ao23_1 \U17/Ucl/U1/U1  ( .x(l[17]), .a(n6), .b(l[17]), .c(n5), .d(\U17/ni 
        ), .e(\U17/nh ) );
    ao23_1 \U17/Uch/U1/U1  ( .x(h[17]), .a(n7), .b(h[17]), .c(n4), .d(i[17]), 
        .e(\U17/nl ) );
    inv_1 \U16/Uii  ( .x(\U16/ni ), .a(i[16]) );
    inv_1 \U16/Uih  ( .x(\U16/nh ), .a(h[16]) );
    inv_1 \U16/Uil  ( .x(\U16/nl ), .a(l[16]) );
    ao23_1 \U16/Ucl/U1/U1  ( .x(l[16]), .a(n9), .b(l[16]), .c(n3), .d(\U16/ni 
        ), .e(\U16/nh ) );
    ao23_1 \U16/Uch/U1/U1  ( .x(h[16]), .a(n9), .b(h[16]), .c(n1), .d(i[16]), 
        .e(\U16/nl ) );
    inv_1 \U15/Uii  ( .x(\U15/ni ), .a(i[15]) );
    inv_1 \U15/Uih  ( .x(\U15/nh ), .a(h[15]) );
    inv_1 \U15/Uil  ( .x(\U15/nl ), .a(l[15]) );
    ao23_1 \U15/Ucl/U1/U1  ( .x(l[15]), .a(n8), .b(l[15]), .c(n1), .d(\U15/ni 
        ), .e(\U15/nh ) );
    ao23_1 \U15/Uch/U1/U1  ( .x(h[15]), .a(n7), .b(h[15]), .c(n1), .d(i[15]), 
        .e(\U15/nl ) );
    inv_1 \U14/Uii  ( .x(\U14/ni ), .a(i[14]) );
    inv_1 \U14/Uih  ( .x(\U14/nh ), .a(h[14]) );
    inv_1 \U14/Uil  ( .x(\U14/nl ), .a(l[14]) );
    ao23_1 \U14/Ucl/U1/U1  ( .x(l[14]), .a(n6), .b(l[14]), .c(n1), .d(\U14/ni 
        ), .e(\U14/nh ) );
    ao23_1 \U14/Uch/U1/U1  ( .x(h[14]), .a(n6), .b(h[14]), .c(n3), .d(i[14]), 
        .e(\U14/nl ) );
    inv_1 \U13/Uii  ( .x(\U13/ni ), .a(i[13]) );
    inv_1 \U13/Uih  ( .x(\U13/nh ), .a(h[13]) );
    inv_1 \U13/Uil  ( .x(\U13/nl ), .a(l[13]) );
    ao23_1 \U13/Ucl/U1/U1  ( .x(l[13]), .a(n6), .b(l[13]), .c(n4), .d(\U13/ni 
        ), .e(\U13/nh ) );
    ao23_1 \U13/Uch/U1/U1  ( .x(h[13]), .a(n6), .b(h[13]), .c(n4), .d(i[13]), 
        .e(\U13/nl ) );
    inv_1 \U12/Uii  ( .x(\U12/ni ), .a(i[12]) );
    inv_1 \U12/Uih  ( .x(\U12/nh ), .a(h[12]) );
    inv_1 \U12/Uil  ( .x(\U12/nl ), .a(l[12]) );
    ao23_1 \U12/Ucl/U1/U1  ( .x(l[12]), .a(n5), .b(l[12]), .c(n4), .d(\U12/ni 
        ), .e(\U12/nh ) );
    ao23_1 \U12/Uch/U1/U1  ( .x(h[12]), .a(n5), .b(h[12]), .c(n4), .d(i[12]), 
        .e(\U12/nl ) );
    inv_1 \U11/Uii  ( .x(\U11/ni ), .a(i[11]) );
    inv_1 \U11/Uih  ( .x(\U11/nh ), .a(h[11]) );
    inv_1 \U11/Uil  ( .x(\U11/nl ), .a(l[11]) );
    ao23_1 \U11/Ucl/U1/U1  ( .x(l[11]), .a(n5), .b(l[11]), .c(n4), .d(\U11/ni 
        ), .e(\U11/nh ) );
    ao23_1 \U11/Uch/U1/U1  ( .x(h[11]), .a(n5), .b(h[11]), .c(n4), .d(i[11]), 
        .e(\U11/nl ) );
    inv_1 \U10/Uii  ( .x(\U10/ni ), .a(i[10]) );
    inv_1 \U10/Uih  ( .x(\U10/nh ), .a(h[10]) );
    inv_1 \U10/Uil  ( .x(\U10/nl ), .a(l[10]) );
    ao23_1 \U10/Ucl/U1/U1  ( .x(l[10]), .a(n5), .b(l[10]), .c(n3), .d(\U10/ni 
        ), .e(\U10/nh ) );
    ao23_1 \U10/Uch/U1/U1  ( .x(h[10]), .a(n5), .b(h[10]), .c(n3), .d(i[10]), 
        .e(\U10/nl ) );
    inv_1 \U9/Uii  ( .x(\U9/ni ), .a(i[9]) );
    inv_1 \U9/Uih  ( .x(\U9/nh ), .a(h[9]) );
    inv_1 \U9/Uil  ( .x(\U9/nl ), .a(l[9]) );
    ao23_1 \U9/Ucl/U1/U1  ( .x(l[9]), .a(n5), .b(l[9]), .c(n3), .d(\U9/ni ), 
        .e(\U9/nh ) );
    ao23_1 \U9/Uch/U1/U1  ( .x(h[9]), .a(n5), .b(h[9]), .c(n3), .d(i[9]), .e(
        \U9/nl ) );
    inv_1 \U8/Uii  ( .x(\U8/ni ), .a(i[8]) );
    inv_1 \U8/Uih  ( .x(\U8/nh ), .a(h[8]) );
    inv_1 \U8/Uil  ( .x(\U8/nl ), .a(l[8]) );
    ao23_1 \U8/Ucl/U1/U1  ( .x(l[8]), .a(n5), .b(l[8]), .c(n3), .d(\U8/ni ), 
        .e(\U8/nh ) );
    ao23_1 \U8/Uch/U1/U1  ( .x(h[8]), .a(n5), .b(h[8]), .c(n3), .d(i[8]), .e(
        \U8/nl ) );
    inv_1 \U7/Uii  ( .x(\U7/ni ), .a(i[7]) );
    inv_1 \U7/Uih  ( .x(\U7/nh ), .a(h[7]) );
    inv_1 \U7/Uil  ( .x(\U7/nl ), .a(l[7]) );
    ao23_1 \U7/Ucl/U1/U1  ( .x(l[7]), .a(n7), .b(l[7]), .c(n3), .d(\U7/ni ), 
        .e(\U7/nh ) );
    ao23_1 \U7/Uch/U1/U1  ( .x(h[7]), .a(n7), .b(h[7]), .c(n2), .d(i[7]), .e(
        \U7/nl ) );
    inv_1 \U6/Uii  ( .x(\U6/ni ), .a(i[6]) );
    inv_1 \U6/Uih  ( .x(\U6/nh ), .a(h[6]) );
    inv_1 \U6/Uil  ( .x(\U6/nl ), .a(l[6]) );
    ao23_1 \U6/Ucl/U1/U1  ( .x(l[6]), .a(n7), .b(l[6]), .c(n2), .d(\U6/ni ), 
        .e(\U6/nh ) );
    ao23_1 \U6/Uch/U1/U1  ( .x(h[6]), .a(n7), .b(h[6]), .c(n2), .d(i[6]), .e(
        \U6/nl ) );
    inv_1 \U5/Uii  ( .x(\U5/ni ), .a(i[5]) );
    inv_1 \U5/Uih  ( .x(\U5/nh ), .a(h[5]) );
    inv_1 \U5/Uil  ( .x(\U5/nl ), .a(l[5]) );
    ao23_1 \U5/Ucl/U1/U1  ( .x(l[5]), .a(n7), .b(l[5]), .c(n2), .d(\U5/ni ), 
        .e(\U5/nh ) );
    ao23_1 \U5/Uch/U1/U1  ( .x(h[5]), .a(n7), .b(h[5]), .c(n2), .d(i[5]), .e(
        \U5/nl ) );
    inv_1 \U4/Uii  ( .x(\U4/ni ), .a(i[4]) );
    inv_1 \U4/Uih  ( .x(\U4/nh ), .a(h[4]) );
    inv_1 \U4/Uil  ( .x(\U4/nl ), .a(l[4]) );
    ao23_1 \U4/Ucl/U1/U1  ( .x(l[4]), .a(n6), .b(l[4]), .c(n2), .d(\U4/ni ), 
        .e(\U4/nh ) );
    ao23_1 \U4/Uch/U1/U1  ( .x(h[4]), .a(n6), .b(h[4]), .c(n2), .d(i[4]), .e(
        \U4/nl ) );
    inv_1 \U3/Uii  ( .x(\U3/ni ), .a(i[3]) );
    inv_1 \U3/Uih  ( .x(\U3/nh ), .a(h[3]) );
    inv_1 \U3/Uil  ( .x(\U3/nl ), .a(l[3]) );
    ao23_1 \U3/Ucl/U1/U1  ( .x(l[3]), .a(n6), .b(l[3]), .c(n2), .d(\U3/ni ), 
        .e(\U3/nh ) );
    ao23_1 \U3/Uch/U1/U1  ( .x(h[3]), .a(n8), .b(h[3]), .c(n1), .d(i[3]), .e(
        \U3/nl ) );
    inv_1 \U2/Uii  ( .x(\U2/ni ), .a(i[2]) );
    inv_1 \U2/Uih  ( .x(\U2/nh ), .a(h[2]) );
    inv_1 \U2/Uil  ( .x(\U2/nl ), .a(l[2]) );
    ao23_1 \U2/Ucl/U1/U1  ( .x(l[2]), .a(n8), .b(l[2]), .c(n1), .d(\U2/ni ), 
        .e(\U2/nh ) );
    ao23_1 \U2/Uch/U1/U1  ( .x(h[2]), .a(n8), .b(h[2]), .c(n1), .d(i[2]), .e(
        \U2/nl ) );
    inv_1 \U1/Uii  ( .x(\U1/ni ), .a(i[1]) );
    inv_1 \U1/Uih  ( .x(\U1/nh ), .a(h[1]) );
    inv_1 \U1/Uil  ( .x(\U1/nl ), .a(l[1]) );
    ao23_1 \U1/Ucl/U1/U1  ( .x(l[1]), .a(n8), .b(l[1]), .c(n1), .d(\U1/ni ), 
        .e(\U1/nh ) );
    ao23_1 \U1/Uch/U1/U1  ( .x(h[1]), .a(n8), .b(h[1]), .c(n1), .d(i[1]), .e(
        \U1/nl ) );
    inv_1 \U0/Uii  ( .x(\U0/ni ), .a(i[0]) );
    inv_1 \U0/Uih  ( .x(\U0/nh ), .a(h[0]) );
    inv_1 \U0/Uil  ( .x(\U0/nl ), .a(l[0]) );
    ao23_1 \U0/Ucl/U1/U1  ( .x(l[0]), .a(n8), .b(l[0]), .c(n1), .d(\U0/ni ), 
        .e(\U0/nh ) );
    ao23_1 \U0/Uch/U1/U1  ( .x(h[0]), .a(n8), .b(h[0]), .c(n1), .d(i[0]), .e(
        \U0/nl ) );
    buf_16 U1 ( .x(n1), .a(n12) );
    buf_16 U2 ( .x(n2), .a(n12) );
    buf_16 U3 ( .x(n3), .a(n12) );
    buf_16 U4 ( .x(n4), .a(n11) );
    buf_16 U5 ( .x(n5), .a(n11) );
    buf_16 U6 ( .x(n6), .a(n11) );
    buf_16 U7 ( .x(n7), .a(n10) );
    buf_16 U8 ( .x(n8), .a(n10) );
    buf_16 U9 ( .x(n9), .a(n10) );
    buf_16 U10 ( .x(n10), .a(req) );
    buf_16 U11 ( .x(n11), .a(req) );
    buf_16 U12 ( .x(n12), .a(req) );
endmodule


module latch_ctrl_1 ( rin, ain, rout, aout, en, reset );
input  rin, aout, reset;
output ain, rout, en;
    wire nreset, na, n1, a, N6, N5, n_rout, n3, \c_rout/ob ;
    inv_1 U0 ( .x(nreset), .a(reset) );
    nor2_1 U1 ( .x(ain), .a(na), .b(n1) );
    inv_1 U2 ( .x(na), .a(a) );
    inv_1 U3 ( .x(N6), .a(N5) );
    inv_1 U4 ( .x(rout), .a(n_rout) );
    and2_1 C9 ( .x(n3), .a(na), .b(N6) );
    or2_1 C11 ( .x(N5), .a(rout), .b(aout) );
    oa21_1 \c_na/__tmp99/U1  ( .x(a), .a(n1), .b(a), .c(rin) );
    oai21_1 \c_rout/U1  ( .x(\c_rout/ob ), .a(aout), .b(n_rout), .c(na) );
    nand2_1 \c_rout/U2  ( .x(n_rout), .a(nreset), .b(\c_rout/ob ) );
    buf_1 U5 ( .x(en), .a(n3) );
    buf_1 U6 ( .x(n1), .a(n3) );
endmodule


module matched_delay_m2cp_resp_dport ( x, a );
input  a;
output x;
    assign x = a;
endmodule


module m2cp_dport ( req_in, ts_o, sel_o, mult_o, we_o, prd_o, seq_o, adr_o, 
    dat_o, ain, ic_seq, ic_pred, ic_size, ic_itag, ic_wd, ic_lock, ic_a, 
    ic_rnw, ic_col, ic_ack, req_out, ts_i, we_i, err_i, rty_i, acc_i, dat_i, 
    aout, ir_rd, ir_err, ir_rnw, ir_ack, tag_id, reset );
input  [2:0] ts_o;
input  [3:0] sel_o;
input  [31:0] adr_o;
input  [31:0] dat_o;
output [1:0] ic_seq;
output [1:0] ic_pred;
output [3:0] ic_size;
output [9:0] ic_itag;
output [63:0] ic_wd;
output [1:0] ic_lock;
output [63:0] ic_a;
output [1:0] ic_rnw;
output [5:0] ic_col;
output [2:0] ts_i;
output [31:0] dat_i;
input  [63:0] ir_rd;
input  [1:0] ir_err;
input  [1:0] ir_rnw;
input  [4:0] tag_id;
input  req_in, mult_o, we_o, prd_o, seq_o, ic_ack, aout, reset;
output ain, req_out, we_i, err_i, rty_i, acc_i, ir_ack;
    wire req_in_delayed, n8, \data[15] , \data[14] , \data[13] , \data[12] , 
        \data[11] , \data[10] , \data[9] , \data[8] , \data[7] , \data[6] , 
        \data[5] , \data[4] , \data[3] , \data[2] , \data[1] , \data[0] , 
        complete_delayed, en, _28_net_, n72, _26_net_, n77, _25_net_, n78, 
        _27_net_, _24_net_, n112, n124, n118, n206, n208, n210, n197, n199, 
        n202, n201, n203, n204, \size[1] , n83, n84, n89, n205, n64, n2, n90, 
        n97, n198, n3, n98, n87, n63, n4, n88, n85, n5, n86, n290, n289, n288, 
        n79, n277, n270, n273, n276, n266, n269, n283, n282, n281, n298, n70, 
        n68, n213, n223, n80, n291, n284, n287, n280, n99, n100, n95, n96, n93, 
        n94, n91, n92, n81, all_r, n69, n300, n294, n302, n296, n306, n292, 
        n304, low_ir_rd, n73, n74, n75, n76, complete, n82, n200, n207, n209, 
        n211, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, 
        n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, 
        n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, 
        n259, n260, n261, n262, n263, n265, n264, n268, n267, n272, n271, n275, 
        n274, n279, n278, n286, n285, n293, n295, n297, n299, n301, n303, n305, 
        n307, n222, n221, n220, n219, n218, n217, n216, n215, all_w, n65, n214, 
        high_ir_rd, \size[0] , n212, n308, n182, n179, n176, n173, n194, n191, 
        n188, n185, n158, n155, n152, n149, n170, n167, n164, n161, n134, n131, 
        n128, n125, n146, n143, n140, n137, n110, n107, n104, n101, n122, n119, 
        n116, n113, n183, n184, n180, n181, n177, n178, n174, n175, n195, n196, 
        n192, n193, n189, n190, n186, n187, n159, n160, n156, n157, n153, n154, 
        n150, n151, n171, n172, n168, n169, n165, n166, n162, n163, n135, n136, 
        n132, n133, n129, n130, n126, n127, n147, n148, n144, n145, n141, n142, 
        n138, n139, n111, n108, n109, n105, n106, n102, n103, n123, n120, n121, 
        n117, n114, n115, n7, n6, n1, comp_basic, \all_read/__tmp99/loop , 
        comp_rd, \Ucol2/ni , \Ucol2/nh , \Ucol2/nl , n11, \Ucol1/ni , 
        \Ucol1/nh , \Ucol1/nl , n9, \Ucol0/ni , \Ucol0/nh , \Ucol0/nl , n10, 
        \Utag4/ni , \Utag4/nh , \Utag4/nl , \Utag3/ni , \Utag3/nh , \Utag3/nl , 
        \Utag2/ni , \Utag2/nh , \Utag2/nl , \Utag1/ni , \Utag1/nh , \Utag1/nl , 
        \Utag0/ni , \Utag0/nh , \Utag0/nl , \Usze1/ni , \Usze1/nh , \Usze1/nl , 
        \Usze0/ni , \Usze0/nh , \Usze0/nl , \Urnw/ni , \Urnw/nh , \Urnw/nl , 
        \Ulock/ni , \Ulock/nh , \Ulock/nl , \Upred/ni , \Upred/nh , \Upred/nl , 
        \Useq/ni , \Useq/nh , \Useq/nl ;
    assign ain = ic_ack;
    assign ts_i[2] = 1'b0;
    assign ts_i[1] = 1'b0;
    assign ts_i[0] = 1'b0;
    assign rty_i = 1'b0;
    assign acc_i = 1'b0;
    matched_delay_m2cp_com_dport U130 ( .x(req_in_delayed), .a(req_in) );
    sr2dr_word_3 Uwd ( .i({dat_o[31], dat_o[30], dat_o[29], dat_o[28], 
        dat_o[27], dat_o[26], dat_o[25], dat_o[24], dat_o[23], dat_o[22], 
        dat_o[21], dat_o[20], dat_o[19], dat_o[18], dat_o[17], dat_o[16], 
        \data[15] , \data[14] , \data[13] , \data[12] , \data[11] , \data[10] , 
        \data[9] , \data[8] , \data[7] , \data[6] , \data[5] , \data[4] , 
        \data[3] , \data[2] , \data[1] , \data[0] }), .req(n8), .h(ic_wd
        [63:32]), .l(ic_wd[31:0]) );
    sr2dr_word_2 Ua ( .i(adr_o), .req(n8), .h(ic_a[63:32]), .l(ic_a[31:0]) );
    latch_ctrl_1 lc ( .rin(complete_delayed), .ain(ir_ack), .rout(req_out), 
        .aout(aout), .en(en), .reset(reset) );
    nand2i_1 U59 ( .x(_28_net_), .a(ir_err[1]), .b(n72) );
    nand2_1 U61 ( .x(_26_net_), .a(n72), .b(n77) );
    nand2i_1 U112 ( .x(_25_net_), .a(ir_err[1]), .b(n78) );
    and2_1 U274 ( .x(_27_net_), .a(ir_rnw[1]), .b(ir_err[0]) );
    inv_1 U275 ( .x(_24_net_), .a(we_o) );
    inv_1 U2 ( .x(n112), .a(ir_rd[4]) );
    inv_1 U3 ( .x(n124), .a(ir_rd[0]) );
    inv_1 U4 ( .x(n118), .a(ir_rd[2]) );
    inv_1 U5 ( .x(n206), .a(dat_o[28]) );
    inv_1 U6 ( .x(n208), .a(dat_o[27]) );
    inv_1 U7 ( .x(n210), .a(dat_o[26]) );
    inv_1 U8 ( .x(n197), .a(dat_o[25]) );
    inv_1 U9 ( .x(n199), .a(dat_o[24]) );
    inv_1 U10 ( .x(n202), .a(dat_o[15]) );
    inv_1 U11 ( .x(n201), .a(dat_o[31]) );
    inv_1 U12 ( .x(n203), .a(dat_o[30]) );
    inv_1 U13 ( .x(n204), .a(dat_o[29]) );
    nor2_1 U14 ( .x(\size[1] ), .a(n83), .b(n84) );
    inv_1 U15 ( .x(n72), .a(ir_rnw[0]) );
    oa21_1 U16 ( .x(n89), .a(n205), .b(n64), .c(n2) );
    inv_1 U24 ( .x(n2), .a(n90) );
    inv_1 U17 ( .x(n205), .a(dat_o[13]) );
    inv_1 U18 ( .x(n64), .a(sel_o[1]) );
    oa21_1 U19 ( .x(n97), .a(n198), .b(n64), .c(n3) );
    inv_1 U276 ( .x(n3), .a(n98) );
    inv_1 U20 ( .x(n198), .a(dat_o[9]) );
    oa21_1 U21 ( .x(n87), .a(n63), .b(n64), .c(n4) );
    inv_1 U277 ( .x(n4), .a(n88) );
    inv_1 U22 ( .x(n63), .a(dat_o[14]) );
    oa21_1 U23 ( .x(n85), .a(n202), .b(n64), .c(n5) );
    inv_1 U278 ( .x(n5), .a(n86) );
    nand2_1 U25 ( .x(n290), .a(n289), .b(n288) );
    nand2_1 U26 ( .x(n79), .a(n277), .b(n270) );
    nor2_1 U27 ( .x(n277), .a(n273), .b(n276) );
    nor2_1 U28 ( .x(n270), .a(n266), .b(n269) );
    nand2_1 U29 ( .x(n283), .a(n282), .b(n281) );
    nand2_1 U30 ( .x(n298), .a(dat_o[20]), .b(n70) );
    inv_1 U31 ( .x(n70), .a(n68) );
    nand2_1 U32 ( .x(n213), .a(n223), .b(sel_o[1]) );
    nand2_1 U33 ( .x(n80), .a(n291), .b(n284) );
    nor2_1 U34 ( .x(n291), .a(n287), .b(n290) );
    nor2_1 U35 ( .x(n284), .a(n280), .b(n283) );
    aoi21_1 U36 ( .x(n99), .a(dat_o[8]), .b(sel_o[1]), .c(n100) );
    aoi21_1 U37 ( .x(n95), .a(dat_o[10]), .b(sel_o[1]), .c(n96) );
    aoi21_1 U38 ( .x(n93), .a(dat_o[11]), .b(sel_o[1]), .c(n94) );
    aoi21_1 U39 ( .x(n91), .a(dat_o[12]), .b(sel_o[1]), .c(n92) );
    inv_1 U40 ( .x(n81), .a(all_r) );
    nand2_1 U42 ( .x(n84), .a(sel_o[0]), .b(sel_o[1]) );
    inv_1 U45 ( .x(n68), .a(sel_o[2]) );
    inv_1 U46 ( .x(n69), .a(n68) );
    nand2_1 U48 ( .x(n83), .a(n70), .b(sel_o[3]) );
    nand2_1 U51 ( .x(n300), .a(dat_o[19]), .b(n69) );
    nand2_1 U52 ( .x(n294), .a(dat_o[22]), .b(n69) );
    nand2_1 U53 ( .x(n302), .a(dat_o[18]), .b(n69) );
    nand2_1 U54 ( .x(n296), .a(dat_o[21]), .b(n69) );
    nand2_1 U55 ( .x(n306), .a(dat_o[16]), .b(n69) );
    nand2_1 U56 ( .x(n292), .a(dat_o[23]), .b(n69) );
    nand2_1 U57 ( .x(n304), .a(dat_o[17]), .b(n69) );
    nand4_1 U60 ( .x(low_ir_rd), .a(n73), .b(n74), .c(n75), .d(n76) );
    nand2_1 U62 ( .x(complete), .a(n81), .b(n82) );
    matched_delay_m2cp_resp_dport mdel ( .x(complete_delayed), .a(complete) );
    inv_1 U63 ( .x(n200), .a(dat_o[8]) );
    inv_1 U64 ( .x(n207), .a(dat_o[12]) );
    inv_1 U65 ( .x(n209), .a(dat_o[11]) );
    inv_1 U66 ( .x(n211), .a(dat_o[10]) );
    nand4_1 U67 ( .x(n224), .a(n225), .b(n226), .c(n227), .d(n228) );
    nand4_1 U68 ( .x(n229), .a(n230), .b(n231), .c(n232), .d(n233) );
    nor2_1 U69 ( .x(n76), .a(n224), .b(n229) );
    nand4_1 U70 ( .x(n234), .a(n235), .b(n236), .c(n237), .d(n238) );
    nand4_1 U71 ( .x(n239), .a(n240), .b(n241), .c(n242), .d(n243) );
    nor2_1 U72 ( .x(n75), .a(n234), .b(n239) );
    nand4_1 U73 ( .x(n244), .a(n245), .b(n246), .c(n247), .d(n248) );
    nand4_1 U74 ( .x(n249), .a(n250), .b(n251), .c(n252), .d(n253) );
    nor2_1 U75 ( .x(n74), .a(n244), .b(n249) );
    nand4_1 U76 ( .x(n254), .a(n255), .b(n256), .c(n257), .d(n258) );
    nand4_1 U77 ( .x(n259), .a(n260), .b(n261), .c(n262), .d(n263) );
    nor2_1 U78 ( .x(n73), .a(n254), .b(n259) );
    nand2_1 U79 ( .x(n266), .a(n265), .b(n264) );
    nand2_1 U80 ( .x(n269), .a(n268), .b(n267) );
    nand2_1 U81 ( .x(n273), .a(n272), .b(n271) );
    nand2_1 U82 ( .x(n276), .a(n275), .b(n274) );
    nand2_1 U83 ( .x(n280), .a(n279), .b(n278) );
    nand2_1 U84 ( .x(n287), .a(n286), .b(n285) );
    nand2_1 U85 ( .x(n86), .a(n292), .b(n293) );
    nand2_1 U86 ( .x(n88), .a(n294), .b(n295) );
    nand2_1 U87 ( .x(n90), .a(n296), .b(n297) );
    nand2_1 U88 ( .x(n92), .a(n298), .b(n299) );
    nand2_1 U89 ( .x(n94), .a(n300), .b(n301) );
    nand2_1 U90 ( .x(n96), .a(n302), .b(n303) );
    nand2_1 U91 ( .x(n98), .a(n304), .b(n305) );
    nand2_1 U92 ( .x(n100), .a(n306), .b(n307) );
    inv_1 U93 ( .x(n222), .a(dat_o[0]) );
    inv_1 U94 ( .x(n221), .a(dat_o[1]) );
    inv_1 U95 ( .x(n220), .a(dat_o[2]) );
    inv_1 U96 ( .x(n219), .a(dat_o[3]) );
    inv_1 U97 ( .x(n218), .a(dat_o[4]) );
    inv_1 U98 ( .x(n217), .a(dat_o[5]) );
    inv_1 U99 ( .x(n216), .a(dat_o[6]) );
    inv_1 U100 ( .x(n215), .a(dat_o[7]) );
    inv_1 U101 ( .x(n77), .a(ir_rnw[1]) );
    inv_1 U103 ( .x(n82), .a(all_w) );
    nand2_1 U104 ( .x(n293), .a(dat_o[31]), .b(sel_o[3]) );
    nand2_1 U109 ( .x(n303), .a(dat_o[26]), .b(sel_o[3]) );
    nand2_1 U110 ( .x(n305), .a(dat_o[25]), .b(sel_o[3]) );
    nand2_1 U111 ( .x(n307), .a(dat_o[24]), .b(sel_o[3]) );
    mux2i_1 U113 ( .x(\data[0] ), .d0(n99), .sl(n65), .d1(n222) );
    mux2i_1 U114 ( .x(\data[10] ), .d0(n211), .sl(n214), .d1(n210) );
    mux2i_1 U115 ( .x(\data[11] ), .d0(n209), .sl(n214), .d1(n208) );
    mux2i_1 U116 ( .x(\data[12] ), .d0(n207), .sl(n214), .d1(n206) );
    mux2i_1 U117 ( .x(\data[13] ), .d0(n205), .sl(n214), .d1(n204) );
    mux2i_1 U118 ( .x(\data[14] ), .d0(n63), .sl(n214), .d1(n203) );
    mux2i_1 U119 ( .x(\data[15] ), .d0(n202), .sl(n214), .d1(n201) );
    mux2i_1 U120 ( .x(\data[1] ), .d0(n97), .sl(n65), .d1(n221) );
    mux2i_1 U121 ( .x(\data[2] ), .d0(n95), .sl(n65), .d1(n220) );
    mux2i_1 U122 ( .x(\data[3] ), .d0(n93), .sl(n65), .d1(n219) );
    mux2i_1 U123 ( .x(\data[4] ), .d0(n91), .sl(n65), .d1(n218) );
    mux2i_1 U124 ( .x(\data[5] ), .d0(n89), .sl(n65), .d1(n217) );
    mux2i_1 U125 ( .x(\data[6] ), .d0(n87), .sl(n65), .d1(n216) );
    mux2i_1 U126 ( .x(\data[7] ), .d0(n85), .sl(n65), .d1(n215) );
    mux2i_1 U127 ( .x(\data[8] ), .d0(n200), .sl(n214), .d1(n199) );
    mux2i_1 U128 ( .x(\data[9] ), .d0(n198), .sl(n214), .d1(n197) );
    nor2_1 U129 ( .x(high_ir_rd), .a(n79), .b(n80) );
    mux2i_1 U131 ( .x(\size[0] ), .d0(n212), .sl(n65), .d1(n213) );
    nand2i_1 U132 ( .x(n308), .a(sel_o[1]), .b(n70) );
    inv_1 U133 ( .x(n255), .a(n182) );
    inv_1 U134 ( .x(n256), .a(n179) );
    inv_1 U135 ( .x(n257), .a(n176) );
    inv_1 U136 ( .x(n258), .a(n173) );
    inv_1 U137 ( .x(n260), .a(n194) );
    inv_1 U138 ( .x(n261), .a(n191) );
    inv_1 U139 ( .x(n262), .a(n188) );
    inv_1 U140 ( .x(n263), .a(n185) );
    inv_1 U141 ( .x(n245), .a(n158) );
    inv_1 U142 ( .x(n246), .a(n155) );
    inv_1 U143 ( .x(n247), .a(n152) );
    inv_1 U144 ( .x(n248), .a(n149) );
    inv_1 U145 ( .x(n250), .a(n170) );
    inv_1 U146 ( .x(n251), .a(n167) );
    inv_1 U147 ( .x(n252), .a(n164) );
    inv_1 U148 ( .x(n253), .a(n161) );
    inv_1 U149 ( .x(n235), .a(n134) );
    inv_1 U150 ( .x(n236), .a(n131) );
    inv_1 U151 ( .x(n237), .a(n128) );
    inv_1 U152 ( .x(n238), .a(n125) );
    inv_1 U153 ( .x(n240), .a(n146) );
    inv_1 U154 ( .x(n241), .a(n143) );
    inv_1 U155 ( .x(n242), .a(n140) );
    inv_1 U156 ( .x(n243), .a(n137) );
    inv_1 U157 ( .x(n225), .a(n110) );
    inv_1 U158 ( .x(n226), .a(n107) );
    inv_1 U159 ( .x(n227), .a(n104) );
    inv_1 U160 ( .x(n228), .a(n101) );
    inv_1 U161 ( .x(n230), .a(n122) );
    inv_1 U162 ( .x(n231), .a(n119) );
    inv_1 U163 ( .x(n232), .a(n116) );
    inv_1 U164 ( .x(n233), .a(n113) );
    nor2_1 U165 ( .x(n272), .a(n252), .b(n253) );
    nor2_1 U166 ( .x(n271), .a(n250), .b(n251) );
    nor2_1 U167 ( .x(n275), .a(n247), .b(n248) );
    nor2_1 U168 ( .x(n274), .a(n245), .b(n246) );
    nor2_1 U169 ( .x(n265), .a(n262), .b(n263) );
    nor2_1 U170 ( .x(n264), .a(n260), .b(n261) );
    nor2_1 U171 ( .x(n268), .a(n257), .b(n258) );
    nor2_1 U172 ( .x(n267), .a(n255), .b(n256) );
    nor2_1 U173 ( .x(n286), .a(n232), .b(n233) );
    nor2_1 U174 ( .x(n285), .a(n230), .b(n231) );
    nor2_1 U175 ( .x(n289), .a(n227), .b(n228) );
    nor2_1 U176 ( .x(n288), .a(n225), .b(n226) );
    nor2_1 U177 ( .x(n279), .a(n242), .b(n243) );
    nor2_1 U178 ( .x(n278), .a(n240), .b(n241) );
    nor2_1 U179 ( .x(n282), .a(n237), .b(n238) );
    nor2_1 U180 ( .x(n281), .a(n235), .b(n236) );
    nand2_1 U181 ( .x(n182), .a(n183), .b(n184) );
    nand2_1 U182 ( .x(n179), .a(n180), .b(n181) );
    nand2_1 U183 ( .x(n176), .a(n177), .b(n178) );
    nand2_1 U184 ( .x(n173), .a(n174), .b(n175) );
    nand2_1 U185 ( .x(n194), .a(n195), .b(n196) );
    nand2_1 U186 ( .x(n191), .a(n192), .b(n193) );
    nand2_1 U187 ( .x(n188), .a(n189), .b(n190) );
    nand2_1 U188 ( .x(n185), .a(n186), .b(n187) );
    nand2_1 U189 ( .x(n158), .a(n159), .b(n160) );
    nand2_1 U190 ( .x(n155), .a(n156), .b(n157) );
    nand2_1 U191 ( .x(n152), .a(n153), .b(n154) );
    nand2_1 U192 ( .x(n149), .a(n150), .b(n151) );
    nand2_1 U193 ( .x(n170), .a(n171), .b(n172) );
    nand2_1 U194 ( .x(n167), .a(n168), .b(n169) );
    nand2_1 U195 ( .x(n164), .a(n165), .b(n166) );
    nand2_1 U196 ( .x(n161), .a(n162), .b(n163) );
    nand2_1 U197 ( .x(n134), .a(n135), .b(n136) );
    nand2_1 U198 ( .x(n131), .a(n132), .b(n133) );
    nand2_1 U199 ( .x(n128), .a(n129), .b(n130) );
    nand2_1 U200 ( .x(n125), .a(n126), .b(n127) );
    nand2_1 U201 ( .x(n146), .a(n147), .b(n148) );
    nand2_1 U202 ( .x(n143), .a(n144), .b(n145) );
    nand2_1 U203 ( .x(n140), .a(n141), .b(n142) );
    nand2_1 U204 ( .x(n137), .a(n138), .b(n139) );
    nand2_1 U205 ( .x(n110), .a(n111), .b(n112) );
    nand2_1 U206 ( .x(n107), .a(n108), .b(n109) );
    nand2_1 U207 ( .x(n104), .a(n105), .b(n106) );
    nand2_1 U208 ( .x(n101), .a(n102), .b(n103) );
    nand2_1 U209 ( .x(n122), .a(n123), .b(n124) );
    nand2_1 U210 ( .x(n119), .a(n120), .b(n121) );
    nand2_1 U211 ( .x(n116), .a(n117), .b(n118) );
    nand2_1 U212 ( .x(n113), .a(n114), .b(n115) );
    inv_1 U213 ( .x(n183), .a(ir_rd[60]) );
    inv_1 U214 ( .x(n184), .a(ir_rd[28]) );
    inv_1 U215 ( .x(n180), .a(ir_rd[61]) );
    inv_1 U216 ( .x(n181), .a(ir_rd[29]) );
    inv_1 U217 ( .x(n177), .a(ir_rd[62]) );
    inv_1 U218 ( .x(n178), .a(ir_rd[30]) );
    inv_1 U219 ( .x(n174), .a(ir_rd[63]) );
    inv_1 U220 ( .x(n175), .a(ir_rd[31]) );
    inv_1 U221 ( .x(n195), .a(ir_rd[56]) );
    inv_1 U222 ( .x(n196), .a(ir_rd[24]) );
    inv_1 U223 ( .x(n192), .a(ir_rd[57]) );
    inv_1 U224 ( .x(n193), .a(ir_rd[25]) );
    inv_1 U225 ( .x(n189), .a(ir_rd[58]) );
    inv_1 U226 ( .x(n190), .a(ir_rd[26]) );
    inv_1 U227 ( .x(n186), .a(ir_rd[59]) );
    inv_1 U228 ( .x(n187), .a(ir_rd[27]) );
    inv_1 U229 ( .x(n159), .a(ir_rd[52]) );
    inv_1 U230 ( .x(n160), .a(ir_rd[20]) );
    inv_1 U231 ( .x(n156), .a(ir_rd[53]) );
    inv_1 U232 ( .x(n157), .a(ir_rd[21]) );
    inv_1 U233 ( .x(n153), .a(ir_rd[54]) );
    inv_1 U234 ( .x(n154), .a(ir_rd[22]) );
    inv_1 U235 ( .x(n150), .a(ir_rd[55]) );
    inv_1 U236 ( .x(n151), .a(ir_rd[23]) );
    inv_1 U237 ( .x(n171), .a(ir_rd[48]) );
    inv_1 U238 ( .x(n172), .a(ir_rd[16]) );
    inv_1 U239 ( .x(n168), .a(ir_rd[49]) );
    inv_1 U240 ( .x(n169), .a(ir_rd[17]) );
    inv_1 U241 ( .x(n165), .a(ir_rd[50]) );
    inv_1 U242 ( .x(n166), .a(ir_rd[18]) );
    inv_1 U243 ( .x(n162), .a(ir_rd[51]) );
    inv_1 U244 ( .x(n163), .a(ir_rd[19]) );
    inv_1 U245 ( .x(n135), .a(ir_rd[44]) );
    inv_1 U246 ( .x(n136), .a(ir_rd[12]) );
    inv_1 U247 ( .x(n132), .a(ir_rd[45]) );
    inv_1 U248 ( .x(n133), .a(ir_rd[13]) );
    inv_1 U249 ( .x(n129), .a(ir_rd[46]) );
    inv_1 U250 ( .x(n130), .a(ir_rd[14]) );
    inv_1 U251 ( .x(n126), .a(ir_rd[47]) );
    inv_1 U252 ( .x(n127), .a(ir_rd[15]) );
    inv_1 U253 ( .x(n147), .a(ir_rd[40]) );
    inv_1 U254 ( .x(n148), .a(ir_rd[8]) );
    inv_1 U255 ( .x(n144), .a(ir_rd[41]) );
    inv_1 U256 ( .x(n145), .a(ir_rd[9]) );
    inv_1 U257 ( .x(n141), .a(ir_rd[42]) );
    inv_1 U258 ( .x(n142), .a(ir_rd[10]) );
    inv_1 U259 ( .x(n138), .a(ir_rd[43]) );
    inv_1 U260 ( .x(n139), .a(ir_rd[11]) );
    inv_1 U261 ( .x(n111), .a(ir_rd[36]) );
    inv_1 U262 ( .x(n108), .a(ir_rd[37]) );
    inv_1 U263 ( .x(n109), .a(ir_rd[5]) );
    inv_1 U264 ( .x(n105), .a(ir_rd[38]) );
    inv_1 U265 ( .x(n106), .a(ir_rd[6]) );
    inv_1 U266 ( .x(n102), .a(ir_rd[39]) );
    inv_1 U267 ( .x(n103), .a(ir_rd[7]) );
    inv_1 U268 ( .x(n123), .a(ir_rd[32]) );
    inv_1 U269 ( .x(n120), .a(ir_rd[33]) );
    inv_1 U270 ( .x(n121), .a(ir_rd[1]) );
    inv_1 U271 ( .x(n117), .a(ir_rd[34]) );
    inv_1 U272 ( .x(n114), .a(ir_rd[35]) );
    inv_1 U273 ( .x(n115), .a(ir_rd[3]) );
    latn_1 \dat_i_reg[30]  ( .q(dat_i[30]), .d(ir_rd[62]), .g(n7) );
    latn_1 \dat_i_reg[28]  ( .q(dat_i[28]), .d(ir_rd[60]), .g(n7) );
    latn_1 \dat_i_reg[27]  ( .q(dat_i[27]), .d(ir_rd[59]), .g(n7) );
    latn_1 \dat_i_reg[26]  ( .q(dat_i[26]), .d(ir_rd[58]), .g(n7) );
    latn_1 \dat_i_reg[25]  ( .q(dat_i[25]), .d(ir_rd[57]), .g(n7) );
    latn_1 \dat_i_reg[24]  ( .q(dat_i[24]), .d(ir_rd[56]), .g(n7) );
    latn_1 \dat_i_reg[22]  ( .q(dat_i[22]), .d(ir_rd[54]), .g(n7) );
    latn_1 \dat_i_reg[20]  ( .q(dat_i[20]), .d(ir_rd[52]), .g(n7) );
    latn_1 \dat_i_reg[19]  ( .q(dat_i[19]), .d(ir_rd[51]), .g(n7) );
    latn_1 \dat_i_reg[18]  ( .q(dat_i[18]), .d(ir_rd[50]), .g(n7) );
    latn_1 \dat_i_reg[17]  ( .q(dat_i[17]), .d(ir_rd[49]), .g(n7) );
    latn_1 \dat_i_reg[16]  ( .q(dat_i[16]), .d(ir_rd[48]), .g(n6) );
    latn_1 \dat_i_reg[14]  ( .q(dat_i[14]), .d(ir_rd[46]), .g(n6) );
    latn_1 \dat_i_reg[12]  ( .q(dat_i[12]), .d(ir_rd[44]), .g(n6) );
    latn_1 \dat_i_reg[10]  ( .q(dat_i[10]), .d(ir_rd[42]), .g(n6) );
    latn_1 \dat_i_reg[8]  ( .q(dat_i[8]), .d(ir_rd[40]), .g(n6) );
    latn_1 \dat_i_reg[6]  ( .q(dat_i[6]), .d(ir_rd[38]), .g(n6) );
    latn_1 \dat_i_reg[4]  ( .q(dat_i[4]), .d(ir_rd[36]), .g(n6) );
    latn_1 \dat_i_reg[3]  ( .q(dat_i[3]), .d(ir_rd[35]), .g(n1) );
    latn_1 \dat_i_reg[2]  ( .q(dat_i[2]), .d(ir_rd[34]), .g(n1) );
    latn_1 \dat_i_reg[1]  ( .q(dat_i[1]), .d(ir_rd[33]), .g(n1) );
    latn_1 \dat_i_reg[0]  ( .q(dat_i[0]), .d(ir_rd[32]), .g(n1) );
    latn_1 we_i_reg ( .q(we_i), .d(ir_rnw[0]), .g(n1) );
    latn_1 err_i_reg ( .q(err_i), .d(ir_err[1]), .g(n1) );
    latn_1 \dat_i_reg[13]  ( .q(dat_i[13]), .d(ir_rd[45]), .g(n6) );
    latn_1 \dat_i_reg[5]  ( .q(dat_i[5]), .d(ir_rd[37]), .g(n1) );
    latn_1 \dat_i_reg[15]  ( .q(dat_i[15]), .d(ir_rd[47]), .g(n6) );
    latn_1 \dat_i_reg[7]  ( .q(dat_i[7]), .d(ir_rd[39]), .g(n1) );
    latn_1 \dat_i_reg[29]  ( .q(dat_i[29]), .d(ir_rd[61]), .g(n6) );
    latn_1 \dat_i_reg[21]  ( .q(dat_i[21]), .d(ir_rd[53]), .g(n1) );
    latn_1 \dat_i_reg[31]  ( .q(dat_i[31]), .d(ir_rd[63]), .g(n6) );
    latn_1 \dat_i_reg[23]  ( .q(dat_i[23]), .d(ir_rd[55]), .g(n1) );
    latn_1 \dat_i_reg[9]  ( .q(dat_i[9]), .d(ir_rd[41]), .g(n6) );
    latn_1 \dat_i_reg[11]  ( .q(dat_i[11]), .d(ir_rd[43]), .g(n1) );
    oa21_1 \all_write/__tmp99/U1  ( .x(all_w), .a(_28_net_), .b(all_w), .c(
        comp_basic) );
    ao31_1 \all_read/__tmp99/aoi  ( .x(\all_read/__tmp99/loop ), .a(comp_basic
        ), .b(comp_rd), .c(_27_net_), .d(all_r) );
    oa21_1 \all_read/__tmp99/outGate  ( .x(all_r), .a(comp_basic), .b(comp_rd), 
        .c(\all_read/__tmp99/loop ) );
    ao222_1 \rd/__tmp99/U1  ( .x(comp_rd), .a(high_ir_rd), .b(low_ir_rd), .c(
        high_ir_rd), .d(comp_rd), .e(low_ir_rd), .f(comp_rd) );
    ao222_1 \basic/__tmp99/U1  ( .x(comp_basic), .a(_25_net_), .b(_26_net_), 
        .c(_25_net_), .d(comp_basic), .e(_26_net_), .f(comp_basic) );
    inv_1 \Ucol2/Uii  ( .x(\Ucol2/ni ), .a(ts_o[2]) );
    inv_1 \Ucol2/Uih  ( .x(\Ucol2/nh ), .a(ic_col[5]) );
    inv_1 \Ucol2/Uil  ( .x(\Ucol2/nl ), .a(ic_col[2]) );
    ao23_1 \Ucol2/Ucl/U1/U1  ( .x(ic_col[2]), .a(n11), .b(ic_col[2]), .c(n8), 
        .d(\Ucol2/ni ), .e(\Ucol2/nh ) );
    ao23_1 \Ucol2/Uch/U1/U1  ( .x(ic_col[5]), .a(n11), .b(ic_col[5]), .c(n8), 
        .d(ts_o[2]), .e(\Ucol2/nl ) );
    inv_1 \Ucol1/Uii  ( .x(\Ucol1/ni ), .a(ts_o[1]) );
    inv_1 \Ucol1/Uih  ( .x(\Ucol1/nh ), .a(ic_col[4]) );
    inv_1 \Ucol1/Uil  ( .x(\Ucol1/nl ), .a(ic_col[1]) );
    ao23_1 \Ucol1/Ucl/U1/U1  ( .x(ic_col[1]), .a(n11), .b(ic_col[1]), .c(n8), 
        .d(\Ucol1/ni ), .e(\Ucol1/nh ) );
    ao23_1 \Ucol1/Uch/U1/U1  ( .x(ic_col[4]), .a(n11), .b(ic_col[4]), .c(n9), 
        .d(ts_o[1]), .e(\Ucol1/nl ) );
    inv_1 \Ucol0/Uii  ( .x(\Ucol0/ni ), .a(ts_o[0]) );
    inv_1 \Ucol0/Uih  ( .x(\Ucol0/nh ), .a(ic_col[3]) );
    inv_1 \Ucol0/Uil  ( .x(\Ucol0/nl ), .a(ic_col[0]) );
    ao23_1 \Ucol0/Ucl/U1/U1  ( .x(ic_col[0]), .a(n11), .b(ic_col[0]), .c(n10), 
        .d(\Ucol0/ni ), .e(\Ucol0/nh ) );
    ao23_1 \Ucol0/Uch/U1/U1  ( .x(ic_col[3]), .a(n11), .b(ic_col[3]), .c(n9), 
        .d(ts_o[0]), .e(\Ucol0/nl ) );
    inv_1 \Utag4/Uii  ( .x(\Utag4/ni ), .a(tag_id[4]) );
    inv_1 \Utag4/Uih  ( .x(\Utag4/nh ), .a(ic_itag[9]) );
    inv_1 \Utag4/Uil  ( .x(\Utag4/nl ), .a(ic_itag[4]) );
    ao23_1 \Utag4/Ucl/U1/U1  ( .x(ic_itag[4]), .a(n11), .b(ic_itag[4]), .c(n9), 
        .d(\Utag4/ni ), .e(\Utag4/nh ) );
    ao23_1 \Utag4/Uch/U1/U1  ( .x(ic_itag[9]), .a(n10), .b(ic_itag[9]), .c(n9), 
        .d(tag_id[4]), .e(\Utag4/nl ) );
    inv_1 \Utag3/Uii  ( .x(\Utag3/ni ), .a(tag_id[3]) );
    inv_1 \Utag3/Uih  ( .x(\Utag3/nh ), .a(ic_itag[8]) );
    inv_1 \Utag3/Uil  ( .x(\Utag3/nl ), .a(ic_itag[3]) );
    ao23_1 \Utag3/Ucl/U1/U1  ( .x(ic_itag[3]), .a(n10), .b(ic_itag[3]), .c(n9), 
        .d(\Utag3/ni ), .e(\Utag3/nh ) );
    ao23_1 \Utag3/Uch/U1/U1  ( .x(ic_itag[8]), .a(n10), .b(ic_itag[8]), .c(n9), 
        .d(tag_id[3]), .e(\Utag3/nl ) );
    inv_1 \Utag2/Uii  ( .x(\Utag2/ni ), .a(tag_id[2]) );
    inv_1 \Utag2/Uih  ( .x(\Utag2/nh ), .a(ic_itag[7]) );
    inv_1 \Utag2/Uil  ( .x(\Utag2/nl ), .a(ic_itag[2]) );
    ao23_1 \Utag2/Ucl/U1/U1  ( .x(ic_itag[2]), .a(n10), .b(ic_itag[2]), .c(n9), 
        .d(\Utag2/ni ), .e(\Utag2/nh ) );
    ao23_1 \Utag2/Uch/U1/U1  ( .x(ic_itag[7]), .a(n10), .b(ic_itag[7]), .c(n10
        ), .d(tag_id[2]), .e(\Utag2/nl ) );
    inv_1 \Utag1/Uii  ( .x(\Utag1/ni ), .a(tag_id[1]) );
    inv_1 \Utag1/Uih  ( .x(\Utag1/nh ), .a(ic_itag[6]) );
    inv_1 \Utag1/Uil  ( .x(\Utag1/nl ), .a(ic_itag[1]) );
    ao23_1 \Utag1/Ucl/U1/U1  ( .x(ic_itag[1]), .a(n11), .b(ic_itag[1]), .c(n9), 
        .d(\Utag1/ni ), .e(\Utag1/nh ) );
    ao23_1 \Utag1/Uch/U1/U1  ( .x(ic_itag[6]), .a(n11), .b(ic_itag[6]), .c(n9), 
        .d(tag_id[1]), .e(\Utag1/nl ) );
    inv_1 \Utag0/Uii  ( .x(\Utag0/ni ), .a(tag_id[0]) );
    inv_1 \Utag0/Uih  ( .x(\Utag0/nh ), .a(ic_itag[5]) );
    inv_1 \Utag0/Uil  ( .x(\Utag0/nl ), .a(ic_itag[0]) );
    ao23_1 \Utag0/Ucl/U1/U1  ( .x(ic_itag[0]), .a(n11), .b(ic_itag[0]), .c(n8), 
        .d(\Utag0/ni ), .e(\Utag0/nh ) );
    ao23_1 \Utag0/Uch/U1/U1  ( .x(ic_itag[5]), .a(n10), .b(ic_itag[5]), .c(n8), 
        .d(tag_id[0]), .e(\Utag0/nl ) );
    inv_1 \Usze1/Uii  ( .x(\Usze1/ni ), .a(\size[1] ) );
    inv_1 \Usze1/Uih  ( .x(\Usze1/nh ), .a(ic_size[3]) );
    inv_1 \Usze1/Uil  ( .x(\Usze1/nl ), .a(ic_size[1]) );
    ao23_1 \Usze1/Ucl/U1/U1  ( .x(ic_size[1]), .a(n10), .b(ic_size[1]), .c(n9), 
        .d(\Usze1/ni ), .e(\Usze1/nh ) );
    ao23_1 \Usze1/Uch/U1/U1  ( .x(ic_size[3]), .a(n10), .b(ic_size[3]), .c(n9), 
        .d(\size[1] ), .e(\Usze1/nl ) );
    inv_1 \Usze0/Uii  ( .x(\Usze0/ni ), .a(\size[0] ) );
    inv_1 \Usze0/Uih  ( .x(\Usze0/nh ), .a(ic_size[2]) );
    inv_1 \Usze0/Uil  ( .x(\Usze0/nl ), .a(ic_size[0]) );
    ao23_1 \Usze0/Ucl/U1/U1  ( .x(ic_size[0]), .a(n10), .b(ic_size[0]), .c(n9), 
        .d(\Usze0/ni ), .e(\Usze0/nh ) );
    ao23_1 \Usze0/Uch/U1/U1  ( .x(ic_size[2]), .a(n10), .b(ic_size[2]), .c(n9), 
        .d(\size[0] ), .e(\Usze0/nl ) );
    inv_1 \Urnw/Uii  ( .x(\Urnw/ni ), .a(_24_net_) );
    inv_1 \Urnw/Uih  ( .x(\Urnw/nh ), .a(ic_rnw[1]) );
    inv_1 \Urnw/Uil  ( .x(\Urnw/nl ), .a(ic_rnw[0]) );
    ao23_1 \Urnw/Ucl/U1/U1  ( .x(ic_rnw[0]), .a(n10), .b(ic_rnw[0]), .c(n9), 
        .d(\Urnw/ni ), .e(\Urnw/nh ) );
    ao23_1 \Urnw/Uch/U1/U1  ( .x(ic_rnw[1]), .a(n10), .b(ic_rnw[1]), .c(n9), 
        .d(_24_net_), .e(\Urnw/nl ) );
    inv_1 \Ulock/Uii  ( .x(\Ulock/ni ), .a(mult_o) );
    inv_1 \Ulock/Uih  ( .x(\Ulock/nh ), .a(ic_lock[1]) );
    inv_1 \Ulock/Uil  ( .x(\Ulock/nl ), .a(ic_lock[0]) );
    ao23_1 \Ulock/Ucl/U1/U1  ( .x(ic_lock[0]), .a(n11), .b(ic_lock[0]), .c(n9), 
        .d(\Ulock/ni ), .e(\Ulock/nh ) );
    ao23_1 \Ulock/Uch/U1/U1  ( .x(ic_lock[1]), .a(n11), .b(ic_lock[1]), .c(n8), 
        .d(mult_o), .e(\Ulock/nl ) );
    inv_1 \Upred/Uii  ( .x(\Upred/ni ), .a(prd_o) );
    inv_1 \Upred/Uih  ( .x(\Upred/nh ), .a(ic_pred[1]) );
    inv_1 \Upred/Uil  ( .x(\Upred/nl ), .a(ic_pred[0]) );
    ao23_1 \Upred/Ucl/U1/U1  ( .x(ic_pred[0]), .a(n11), .b(ic_pred[0]), .c(n8), 
        .d(\Upred/ni ), .e(\Upred/nh ) );
    ao23_1 \Upred/Uch/U1/U1  ( .x(ic_pred[1]), .a(n10), .b(ic_pred[1]), .c(n8), 
        .d(prd_o), .e(\Upred/nl ) );
    inv_1 \Useq/Uii  ( .x(\Useq/ni ), .a(seq_o) );
    inv_1 \Useq/Uih  ( .x(\Useq/nh ), .a(ic_seq[1]) );
    inv_1 \Useq/Uil  ( .x(\Useq/nl ), .a(ic_seq[0]) );
    ao23_1 \Useq/Ucl/U1/U1  ( .x(ic_seq[0]), .a(n10), .b(ic_seq[0]), .c(n8), 
        .d(\Useq/ni ), .e(\Useq/nh ) );
    ao23_1 \Useq/Uch/U1/U1  ( .x(ic_seq[1]), .a(n11), .b(ic_seq[1]), .c(n8), 
        .d(seq_o), .e(\Useq/nl ) );
    buf_3 U1 ( .x(n1), .a(en) );
    buf_3 U41 ( .x(n7), .a(en) );
    buf_3 U43 ( .x(n6), .a(en) );
    inv_2 U44 ( .x(n214), .a(n308) );
    buf_3 U47 ( .x(n65), .a(sel_o[0]) );
    nand3i_0 U49 ( .x(n212), .a(sel_o[1]), .b(sel_o[3]), .c(n70) );
    nor2_0 U50 ( .x(n223), .a(n70), .b(sel_o[3]) );
    nand2_0 U58 ( .x(n297), .a(dat_o[29]), .b(sel_o[3]) );
    nand2_0 U102 ( .x(n301), .a(dat_o[27]), .b(sel_o[3]) );
    nand2_0 U105 ( .x(n299), .a(dat_o[28]), .b(sel_o[3]) );
    nand2_0 U106 ( .x(n295), .a(dat_o[30]), .b(sel_o[3]) );
    inv_0 U107 ( .x(n78), .a(ir_err[0]) );
    buf_16 U108 ( .x(n8), .a(req_in_delayed) );
    buf_16 U279 ( .x(n9), .a(req_in_delayed) );
    buf_16 U280 ( .x(n10), .a(req_in_delayed) );
    buf_16 U281 ( .x(n11), .a(req_in_delayed) );
endmodule


module i_adec_dport ( e_h, e_l, r_h, r_l, ah, al, e_bare, e_dm, e_im, e_wish, 
    r_bare, r_dm, r_im, r_wish, force_bare );
output [3:0] e_h;
output [3:0] e_l;
output [3:0] r_h;
output [3:0] r_l;
input  [31:0] ah;
input  [31:0] al;
input  [3:0] e_bare;
input  [3:0] e_dm;
input  [3:0] e_im;
input  [3:0] e_wish;
input  [3:0] r_bare;
input  [3:0] r_dm;
input  [3:0] r_im;
input  [3:0] r_wish;
input  force_bare;
    wire e_h_2, e_h_0, e_l_3, e_l_2, e_l_0, wish_i, n6, bare_i, im_i, n7, dm_i, 
        \r_l[2] , \r_l[0] , n1, n2, n3, \r_l[3] , n12;
    assign e_h[3] = 1'b0;
    assign e_h[2] = e_h_2;
    assign e_h[0] = e_h_0;
    assign e_l[3] = e_l_3;
    assign e_l[2] = e_l_2;
    assign e_l[0] = e_l_0;
    assign r_h[3] = e_l_2;
    assign r_h[2] = e_h_0;
    assign r_h[0] = 1'b0;
    assign r_l[3] = e_h_2;
    assign r_l[2] = e_l_0;
    assign r_l[0] = e_l_3;
    ao222_1 \U1632/U18/U1/U1  ( .x(wish_i), .a(n6), .b(al[30]), .c(n6), .d(
        wish_i), .e(al[30]), .f(wish_i) );
    ao222_1 \U1633/U18/U1/U1  ( .x(bare_i), .a(n6), .b(ah[30]), .c(n6), .d(
        bare_i), .e(ah[30]), .f(bare_i) );
    ao222_1 \U1634/U18/U1/U1  ( .x(im_i), .a(al[11]), .b(n7), .c(al[11]), .d(
        im_i), .e(n7), .f(im_i) );
    ao222_1 \U1635/U18/U1/U1  ( .x(dm_i), .a(ah[11]), .b(n7), .c(ah[11]), .d(
        dm_i), .e(n7), .f(dm_i) );
    or3_1 U1 ( .x(\r_l[2] ), .a(wish_i), .b(bare_i), .c(force_bare) );
    or2_1 U2 ( .x(r_l[1]), .a(e_l_0), .b(im_i) );
    or2_1 U3 ( .x(\r_l[0] ), .a(dm_i), .b(r_l[1]) );
    nor2_0 U4 ( .x(n1), .a(bare_i), .b(force_bare) );
    aoi21_1 U6 ( .x(n2), .a(n3), .b(im_i), .c(r_h[1]) );
    inv_0 U8 ( .x(n3), .a(force_bare) );
    nor2i_0 U9 ( .x(\r_l[3] ), .a(wish_i), .b(force_bare) );
    nor2i_0 U10 ( .x(n12), .a(dm_i), .b(force_bare) );
    inv_0 U11 ( .x(e_h[1]), .a(n1) );
    buf_1 U15 ( .x(n6), .a(ah[31]) );
    buf_1 U16 ( .x(n7), .a(al[31]) );
    nand2_2 U17 ( .x(e_l_2), .a(n2), .b(n1) );
    buf_1 U18 ( .x(r_h[1]), .a(n12) );
    inv_2 U19 ( .x(e_h_0), .a(n2) );
    buf_3 U20 ( .x(e_l_3), .a(\r_l[0] ) );
    buf_3 U21 ( .x(e_l_0), .a(\r_l[2] ) );
    buf_3 U22 ( .x(e_h_2), .a(\r_l[3] ) );
    nand2i_2 U23 ( .x(e_l[1]), .a(e_h_2), .b(n2) );
endmodule


module chain_selement_ga_8 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_symbol_4 ( o, txack, txack_last, e, oa, r, txreq );
output [2:0] o;
input  [1:0] e;
input  [1:0] r;
input  oa, txreq;
output txack, txack_last;
    wire ack, net10, \c[0] , \c[1] ;
    chain_selement_ga_8 U1239 ( .Aa(ack), .Br(net10), .Ar(txreq), .Ba(oa) );
    and2_1 \U1229_0_/U8  ( .x(o[0]), .a(\c[0] ), .b(net10) );
    and2_1 \U1229_1_/U8  ( .x(o[1]), .a(\c[1] ), .b(net10) );
    and2_1 \U1229_2_/U8  ( .x(o[2]), .a(e[1]), .b(net10) );
    ao23_1 \U1251/U19/U21/U1/U1  ( .x(txack_last), .a(ack), .b(txack_last), 
        .c(ack), .d(e[1]), .e(e[1]) );
    ao23_1 \U1250/U19/U21/U1/U1  ( .x(txack), .a(ack), .b(txack), .c(ack), .d(
        e[0]), .e(e[0]) );
    ao222_1 \U1210/U18/U1/U1  ( .x(\c[0] ), .a(e[0]), .b(r[0]), .c(e[0]), .d(
        \c[0] ), .e(r[0]), .f(\c[0] ) );
    ao222_1 \U1209/U18/U1/U1  ( .x(\c[1] ), .a(e[0]), .b(r[1]), .c(e[0]), .d(
        \c[1] ), .e(r[1]), .f(\c[1] ) );
endmodule


module chain_selement_ga_9 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_symbol_5 ( o, txack, txack_last, e, oa, r, txreq );
output [2:0] o;
input  [1:0] e;
input  [1:0] r;
input  oa, txreq;
output txack, txack_last;
    wire ack, net10, \c[0] , \c[1] ;
    chain_selement_ga_9 U1239 ( .Aa(ack), .Br(net10), .Ar(txreq), .Ba(oa) );
    and2_1 \U1229_0_/U8  ( .x(o[0]), .a(\c[0] ), .b(net10) );
    and2_1 \U1229_1_/U8  ( .x(o[1]), .a(\c[1] ), .b(net10) );
    and2_1 \U1229_2_/U8  ( .x(o[2]), .a(e[1]), .b(net10) );
    ao23_1 \U1251/U19/U21/U1/U1  ( .x(txack_last), .a(ack), .b(txack_last), 
        .c(ack), .d(e[1]), .e(e[1]) );
    ao23_1 \U1250/U19/U21/U1/U1  ( .x(txack), .a(ack), .b(txack), .c(ack), .d(
        e[0]), .e(e[0]) );
    ao222_1 \U1210/U18/U1/U1  ( .x(\c[0] ), .a(e[0]), .b(r[0]), .c(e[0]), .d(
        \c[0] ), .e(r[0]), .f(\c[0] ) );
    ao222_1 \U1209/U18/U1/U1  ( .x(\c[1] ), .a(e[0]), .b(r[1]), .c(e[0]), .d(
        \c[1] ), .e(r[1]), .f(\c[1] ) );
endmodule


module chain_selement_ga_10 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_symbol_6 ( o, txack, txack_last, e, oa, r, txreq );
output [2:0] o;
input  [1:0] e;
input  [1:0] r;
input  oa, txreq;
output txack, txack_last;
    wire ack, net10, \c[0] , \c[1] ;
    chain_selement_ga_10 U1239 ( .Aa(ack), .Br(net10), .Ar(txreq), .Ba(oa) );
    and2_1 \U1229_0_/U8  ( .x(o[0]), .a(\c[0] ), .b(net10) );
    and2_1 \U1229_1_/U8  ( .x(o[1]), .a(\c[1] ), .b(net10) );
    and2_1 \U1229_2_/U8  ( .x(o[2]), .a(e[1]), .b(net10) );
    ao23_1 \U1251/U19/U21/U1/U1  ( .x(txack_last), .a(ack), .b(txack_last), 
        .c(ack), .d(e[1]), .e(e[1]) );
    ao23_1 \U1250/U19/U21/U1/U1  ( .x(txack), .a(ack), .b(txack), .c(ack), .d(
        e[0]), .e(e[0]) );
    ao222_1 \U1210/U18/U1/U1  ( .x(\c[0] ), .a(e[0]), .b(r[0]), .c(e[0]), .d(
        \c[0] ), .e(r[0]), .f(\c[0] ) );
    ao222_1 \U1209/U18/U1/U1  ( .x(\c[1] ), .a(e[0]), .b(r[1]), .c(e[0]), .d(
        \c[1] ), .e(r[1]), .f(\c[1] ) );
endmodule


module chain_selement_ga_11 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_symbol_7 ( o, txack, txack_last, e, oa, r, txreq );
output [2:0] o;
input  [1:0] e;
input  [1:0] r;
input  oa, txreq;
output txack, txack_last;
    wire ack, net10, \c[0] , \c[1] ;
    chain_selement_ga_11 U1239 ( .Aa(ack), .Br(net10), .Ar(txreq), .Ba(oa) );
    and2_1 \U1229_0_/U8  ( .x(o[0]), .a(\c[0] ), .b(net10) );
    and2_1 \U1229_1_/U8  ( .x(o[1]), .a(\c[1] ), .b(net10) );
    and2_1 \U1229_2_/U8  ( .x(o[2]), .a(e[1]), .b(net10) );
    ao23_1 \U1251/U19/U21/U1/U1  ( .x(txack_last), .a(ack), .b(txack_last), 
        .c(ack), .d(e[1]), .e(e[1]) );
    ao23_1 \U1250/U19/U21/U1/U1  ( .x(txack), .a(ack), .b(txack), .c(ack), .d(
        e[0]), .e(e[0]) );
    ao222_1 \U1210/U18/U1/U1  ( .x(\c[0] ), .a(e[0]), .b(r[0]), .c(e[0]), .d(
        \c[0] ), .e(r[0]), .f(\c[0] ) );
    ao222_1 \U1209/U18/U1/U1  ( .x(\c[1] ), .a(e[0]), .b(r[1]), .c(e[0]), .d(
        \c[1] ), .e(r[1]), .f(\c[1] ) );
endmodule


module chain_selement_ga_78 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_tx_dport ( o, rtxack, e_h, e_l, noa, r_h, r_l, rtxreq );
output [4:0] o;
input  [3:0] e_h;
input  [3:0] e_l;
input  [3:0] r_h;
input  [3:0] r_l;
input  noa, rtxreq;
output rtxack;
    wire net33, \last[4] , net60, \r3[2] , \r3[1] , \r3[0] , net40, \last[3] , 
        \r2[2] , \r2[1] , \r2[0] , net47, \last[2] , \r1[2] , \r1[1] , \r1[0] , 
        net50, \last[1] , \r0[2] , \r0[1] , \r0[0] , \last[0] , eopsym, 
        \I8/nb , \I8/na , \net55[1] , \net55[0] , \net52[1] , \net52[0] , 
        \I11/nc , \I11/nb , \I11/na , net16, net11, net9, net6, 
        \I7_0_/U25/U1/clr , \I7_0_/U25/U1/ob , \I7_1_/U25/U1/clr , 
        \I7_1_/U25/U1/ob ;
    assign o[3] = 1'b0;
    assign o[2] = 1'b0;
    route_symbol_4 I0 ( .o({\r3[2] , \r3[1] , \r3[0] }), .txack(net33), 
        .txack_last(\last[4] ), .e({e_h[3], e_l[3]}), .oa(net60), .r({r_h[3], 
        r_l[3]}), .txreq(rtxreq) );
    route_symbol_5 I1 ( .o({\r2[2] , \r2[1] , \r2[0] }), .txack(net40), 
        .txack_last(\last[3] ), .e({e_h[2], e_l[2]}), .oa(net60), .r({r_h[2], 
        r_l[2]}), .txreq(net33) );
    route_symbol_6 I2 ( .o({\r1[2] , \r1[1] , \r1[0] }), .txack(net47), 
        .txack_last(\last[2] ), .e({e_h[1], e_l[1]}), .oa(net60), .r({r_h[1], 
        r_l[1]}), .txreq(net40) );
    route_symbol_7 I3 ( .o({\r0[2] , \r0[1] , \r0[0] }), .txack(net50), 
        .txack_last(\last[1] ), .e({e_h[0], e_l[0]}), .oa(net60), .r({r_h[0], 
        r_l[0]}), .txreq(net47) );
    chain_selement_ga_78 I9 ( .Aa(\last[0] ), .Br(eopsym), .Ar(net50), .Ba(
        net60) );
    nor3_1 \I8/U27  ( .x(\I8/nb ), .a(o[4]), .b(1'b0), .c(1'b0) );
    nor2_1 \I8/U26  ( .x(\I8/na ), .a(o[1]), .b(o[0]) );
    nand2_2 \I8/U29  ( .x(net60), .a(\I8/nb ), .b(\I8/na ) );
    or2_1 \I13_0_/U12  ( .x(\net55[1] ), .a(\r1[0] ), .b(\r0[0] ) );
    or2_1 \I13_1_/U12  ( .x(\net55[0] ), .a(\r1[1] ), .b(\r0[1] ) );
    or2_1 \I14_0_/U12  ( .x(\net52[1] ), .a(\r3[0] ), .b(\r2[0] ) );
    or2_1 \I14_1_/U12  ( .x(\net52[0] ), .a(\r3[1] ), .b(\r2[1] ) );
    nand3_1 \I11/U31  ( .x(rtxack), .a(\I11/nc ), .b(\I11/nb ), .c(\I11/na )
         );
    inv_1 \I11/U33  ( .x(\I11/nc ), .a(\last[0] ) );
    nor2_1 \I11/U26  ( .x(\I11/na ), .a(\last[3] ), .b(\last[4] ) );
    nor2_1 \I11/U32  ( .x(\I11/nb ), .a(\last[1] ), .b(\last[2] ) );
    nor2_1 \I16/U5  ( .x(net16), .a(\r1[2] ), .b(\r0[2] ) );
    nor2_1 \I5/U5  ( .x(net11), .a(\r3[2] ), .b(\r2[2] ) );
    nand3_1 \I17/U9  ( .x(net9), .a(net6), .b(net11), .c(net16) );
    inv_1 \I18/U3  ( .x(net6), .a(eopsym) );
    oa31_1 \I7_0_/U25/U1/Uclr  ( .x(\I7_0_/U25/U1/clr ), .a(noa), .b(
        \net55[1] ), .c(\net52[1] ), .d(o[0]) );
    oaoi211_1 \I7_0_/U25/U1/Uaoi  ( .x(\I7_0_/U25/U1/ob ), .a(\net55[1] ), .b(
        \net52[1] ), .c(noa), .d(\I7_0_/U25/U1/clr ) );
    inv_2 \I7_0_/U25/U1/Ui  ( .x(o[0]), .a(\I7_0_/U25/U1/ob ) );
    oa31_1 \I7_1_/U25/U1/Uclr  ( .x(\I7_1_/U25/U1/clr ), .a(noa), .b(
        \net55[0] ), .c(\net52[0] ), .d(o[1]) );
    oaoi211_1 \I7_1_/U25/U1/Uaoi  ( .x(\I7_1_/U25/U1/ob ), .a(\net55[0] ), .b(
        \net52[0] ), .c(noa), .d(\I7_1_/U25/U1/clr ) );
    inv_2 \I7_1_/U25/U1/Ui  ( .x(o[1]), .a(\I7_1_/U25/U1/ob ) );
    ao222_1 \I15/U18/U1/U1  ( .x(o[4]), .a(noa), .b(net9), .c(noa), .d(o[4]), 
        .e(net9), .f(o[4]) );
endmodule


module chain_irdemuxNew_1 ( err, ncback, rd, rnw, status, cbh, cbl, nReset, 
    nack, statusack );
output [1:0] err;
output [63:0] rd;
output [1:0] rnw;
output [1:0] status;
input  [7:0] cbh;
input  [7:0] cbl;
input  nReset, nack, statusack;
output ncback;
    wire bpullcd, pullcd, net162, reset, pkt_normal, \opc_l[2] , \opc_l[1] , 
        net150, \opc_h[1] , pkt_done, write, net193, \ncd[0] , \ncd[1] , 
        \ncd[2] , \ncd[3] , \ncd[4] , \ncd[5] , \ncd[6] , \ncd[7] , 
        start_receiving, notify, net176, net86, net172, net173, net171, net169, 
        net170, net168, net166, net167, \U1664/x[3] , \U1664/U28/Z , 
        \U1664/x[0] , \U1664/U32/Z , \U1664/x[2] , \U1664/U29/Z , \U1664/y[0] , 
        \U1664/x[1] , \U1664/U33/Z , \U1664/y[1] , \U1664/U30/Z , 
        \U1664/U31/Z , \U1664/U37/Z , \U1697/U21/nr , net149, \U1697/U21/nd , 
        \U1697/U21/n2 , \U307/U21/nr , \U307/U21/nd , \U307/U21/n2 , 
        \U1698/nr , \U1698/nd , \U1698/n2 , read, n17, \opc_h[0] , n18, 
        \opc_l[0] , net0187, net0208, \I6/latch , \I6/nlocalcd , \I6/localcd , 
        \I6/ncd[0] , \I6/ncd[1] , \I6/ncd[2] , \I6/oh[2] , \I6/ncd[3] , 
        \I6/ol[3] , \I6/oh[3] , \I6/ncd[4] , \I6/ol[4] , \I6/oh[4] , 
        \I6/ncd[5] , \I6/ncd[6] , \I6/ol[6] , \I6/oh[6] , \I6/ncd[7] , 
        \I6/ol[7] , \I6/oh[7] , \I6/ctrlack_internal , \I6/acb , \I6/ba , 
        \I6/driveh , net139, \I6/drivel , n12, n13, \I6/U4/U28/U1/clr , 
        \I6/U4/U28/U1/set , \I6/U1/Z , n14, \I6/U1664/x[3] , \I6/U1664/U28/Z , 
        \I6/U1664/x[0] , \I6/U1664/U32/Z , \I6/U1664/x[2] , \I6/U1664/U29/Z , 
        \I6/U1664/y[0] , \I6/U1664/x[1] , \I6/U1664/U33/Z , \I6/U1664/y[1] , 
        \I6/U1664/U30/Z , \I6/U1664/U31/Z , \I6/U1664/U37/Z , \I6/U1669/nr , 
        \I6/U1669/nd , \I6/U1669/n2 , \U1667/latch , \U1667/nlocalcd , 
        \U1667/localcd , \U1667/ncd[0] , \U1667/ncd[1] , \U1667/ncd[2] , 
        \U1667/ncd[3] , \U1667/ncd[4] , \U1667/ncd[5] , \U1667/ncd[6] , 
        \U1667/ncd[7] , \U1667/ctrlack_internal , \U1667/acb , \U1667/ba , 
        \U1667/driveh , read_lhw, \U1667/drivel , n11, n10, 
        \U1667/U4/U28/U1/clr , \U1667/U4/U28/U1/set , \U1667/U1/Z , 
        \U1667/U1664/x[3] , \U1667/U1664/U28/Z , \U1667/U1664/x[0] , 
        \U1667/U1664/U32/Z , \U1667/U1664/x[2] , \U1667/U1664/U29/Z , 
        \U1667/U1664/y[0] , \U1667/U1664/x[1] , \U1667/U1664/U33/Z , 
        \U1667/U1664/y[1] , \U1667/U1664/U30/Z , \U1667/U1664/U31/Z , 
        \U1667/U1664/U37/Z , \U1667/U1669/nr , \U1667/U1669/nd , 
        \U1667/U1669/n2 , \U1650/latch , \U1650/nlocalcd , \U1650/localcd , 
        \U1650/ncd[0] , \U1650/ol[0] , \U1650/oh[0] , \U1650/ncd[1] , 
        \U1650/ol[1] , \U1650/oh[1] , \U1650/ncd[2] , \U1650/ol[2] , 
        \U1650/oh[2] , \U1650/ncd[3] , \U1650/ol[3] , \U1650/oh[3] , 
        \U1650/ncd[4] , \U1650/ol[4] , \U1650/oh[4] , \U1650/ncd[5] , 
        \col_l[0] , \col_h[0] , \U1650/ncd[6] , \col_l[1] , \col_h[1] , 
        \U1650/ncd[7] , \col_l[2] , \col_h[2] , \U1650/ctrlack_internal , 
        \U1650/acb , \U1650/ba , \U1650/driveh , \U1650/drivel , n7, n9, n8, 
        \U1650/U4/U28/U1/clr , \U1650/U4/U28/U1/set , \U1650/U1/Z , 
        \U1650/U1664/x[3] , \U1650/U1664/U28/Z , \U1650/U1664/x[0] , 
        \U1650/U1664/U32/Z , \U1650/U1664/x[2] , \U1650/U1664/U29/Z , 
        \U1650/U1664/y[0] , \U1650/U1664/x[1] , \U1650/U1664/U33/Z , 
        \U1650/U1664/y[1] , \U1650/U1664/U30/Z , \U1650/U1664/U31/Z , 
        \U1650/U1664/U37/Z , \U1650/U1669/nr , \U1650/U1669/nd , 
        \U1650/U1669/n2 , \U1666/latch , \U1666/nlocalcd , \U1666/localcd , 
        \U1666/ncd[0] , \U1666/ncd[1] , \U1666/ncd[2] , \U1666/ncd[3] , 
        \U1666/ncd[4] , \U1666/ncd[5] , \U1666/ncd[6] , \U1666/ncd[7] , 
        \U1666/ctrlack_internal , \U1666/acb , \U1666/ba , \U1666/driveh , 
        \U1666/drivel , n6, n5, \U1666/U4/U28/U1/clr , \U1666/U4/U28/U1/set , 
        \U1666/U1/Z , \U1666/U1664/x[3] , \U1666/U1664/U28/Z , 
        \U1666/U1664/x[0] , \U1666/U1664/U32/Z , \U1666/U1664/x[2] , 
        \U1666/U1664/U29/Z , \U1666/U1664/y[0] , \U1666/U1664/x[1] , 
        \U1666/U1664/U33/Z , \U1666/U1664/y[1] , \U1666/U1664/U30/Z , 
        \U1666/U1664/U31/Z , \U1666/U1664/U37/Z , \U1666/U1669/nr , 
        \U1666/U1669/nd , \U1666/U1669/n2 , net94, \I1/latch , \I1/nlocalcd , 
        \I1/localcd , \I1/ncd[0] , \I1/ncd[1] , \I1/ncd[2] , \I1/ncd[3] , 
        \I1/ncd[4] , \I1/ncd[5] , \I1/ncd[6] , \I1/ncd[7] , 
        \I1/ctrlack_internal , \I1/acb , \I1/ba , \I1/driveh , net103, 
        \I1/drivel , n4, n3, \I1/U4/U28/U1/clr , \I1/U4/U28/U1/set , \I1/U1/Z , 
        \I1/U1664/x[3] , \I1/U1664/U28/Z , \I1/U1664/x[0] , \I1/U1664/U32/Z , 
        \I1/U1664/x[2] , \I1/U1664/U29/Z , \I1/U1664/y[0] , \I1/U1664/x[1] , 
        \I1/U1664/U33/Z , \I1/U1664/y[1] , \I1/U1664/U30/Z , \I1/U1664/U31/Z , 
        \I1/U1664/U37/Z , \I1/U1669/nr , \I1/U1669/nd , \I1/U1669/n2 , 
        \I2/latch , \I2/nlocalcd , \I2/localcd , \I2/ncd[0] , \I2/ncd[1] , 
        \I2/ncd[2] , \I2/ncd[3] , \I2/ncd[4] , \I2/ncd[5] , \I2/ncd[6] , 
        \I2/ncd[7] , \I2/ctrlack_internal , \I2/acb , \I2/ba , \I2/driveh , 
        \I2/drivel , n2, n1, \I2/U4/U28/U1/clr , \I2/U4/U28/U1/set , \I2/U1/Z , 
        \I2/U1664/x[3] , \I2/U1664/U28/Z , \I2/U1664/x[0] , \I2/U1664/U32/Z , 
        \I2/U1664/x[2] , \I2/U1664/U29/Z , \I2/U1664/y[0] , \I2/U1664/x[1] , 
        \I2/U1664/U33/Z , \I2/U1664/y[1] , \I2/U1664/U30/Z , \I2/U1664/U31/Z , 
        \I2/U1664/U37/Z , \I2/U1669/nr , \I2/U1669/nd , \I2/U1669/n2 ;
    buf_1 U262 ( .x(bpullcd), .a(pullcd) );
    or2_4 \U1674/U12  ( .x(net162), .a(nack), .b(reset) );
    and2_4 \U1785/U8  ( .x(pkt_normal), .a(\opc_l[2] ), .b(\opc_l[1] ) );
    and2_4 \U1777/U8  ( .x(net150), .a(\opc_l[2] ), .b(\opc_h[1] ) );
    or3_1 \U1813/U12  ( .x(pkt_done), .a(write), .b(reset), .c(net193) );
    nor2_1 \U1651_0_/U5  ( .x(\ncd[0] ), .a(cbh[0]), .b(cbl[0]) );
    nor2_1 \U1651_1_/U5  ( .x(\ncd[1] ), .a(cbh[1]), .b(cbl[1]) );
    nor2_1 \U1651_2_/U5  ( .x(\ncd[2] ), .a(cbh[2]), .b(cbl[2]) );
    nor2_1 \U1651_3_/U5  ( .x(\ncd[3] ), .a(cbh[3]), .b(cbl[3]) );
    nor2_1 \U1651_4_/U5  ( .x(\ncd[4] ), .a(cbh[4]), .b(cbl[4]) );
    nor2_1 \U1651_5_/U5  ( .x(\ncd[5] ), .a(cbh[5]), .b(cbl[5]) );
    nor2_1 \U1651_6_/U5  ( .x(\ncd[6] ), .a(cbh[6]), .b(cbl[6]) );
    nor2_1 \U1651_7_/U5  ( .x(\ncd[7] ), .a(cbh[7]), .b(cbl[7]) );
    nor2_1 \U1812/U5  ( .x(start_receiving), .a(notify), .b(net176) );
    nor2_1 \I7/U5  ( .x(net86), .a(net172), .b(net173) );
    nor2_1 \I4/U5  ( .x(net171), .a(net169), .b(net170) );
    nor2_1 \I3/U5  ( .x(net168), .a(net166), .b(net167) );
    inv_2 \U1675/U3  ( .x(reset), .a(nReset) );
    nand3_2 \U193/U16  ( .x(ncback), .a(net86), .b(net171), .c(net168) );
    ao222_1 \U1811/U18/U1/U1  ( .x(net176), .a(net162), .b(pkt_done), .c(
        net162), .d(net176), .e(pkt_done), .f(net176) );
    aoi222_1 \U1664/U28/U30/U1  ( .x(\U1664/x[3] ), .a(\ncd[7] ), .b(\ncd[6] ), 
        .c(\ncd[7] ), .d(\U1664/U28/Z ), .e(\ncd[6] ), .f(\U1664/U28/Z ) );
    inv_1 \U1664/U28/U30/Uinv  ( .x(\U1664/U28/Z ), .a(\U1664/x[3] ) );
    aoi222_1 \U1664/U32/U30/U1  ( .x(\U1664/x[0] ), .a(\ncd[1] ), .b(\ncd[0] ), 
        .c(\ncd[1] ), .d(\U1664/U32/Z ), .e(\ncd[0] ), .f(\U1664/U32/Z ) );
    inv_1 \U1664/U32/U30/Uinv  ( .x(\U1664/U32/Z ), .a(\U1664/x[0] ) );
    aoi222_1 \U1664/U29/U30/U1  ( .x(\U1664/x[2] ), .a(\ncd[5] ), .b(\ncd[4] ), 
        .c(\ncd[5] ), .d(\U1664/U29/Z ), .e(\ncd[4] ), .f(\U1664/U29/Z ) );
    inv_1 \U1664/U29/U30/Uinv  ( .x(\U1664/U29/Z ), .a(\U1664/x[2] ) );
    aoi222_1 \U1664/U33/U30/U1  ( .x(\U1664/y[0] ), .a(\U1664/x[1] ), .b(
        \U1664/x[0] ), .c(\U1664/x[1] ), .d(\U1664/U33/Z ), .e(\U1664/x[0] ), 
        .f(\U1664/U33/Z ) );
    inv_1 \U1664/U33/U30/Uinv  ( .x(\U1664/U33/Z ), .a(\U1664/y[0] ) );
    aoi222_1 \U1664/U30/U30/U1  ( .x(\U1664/y[1] ), .a(\U1664/x[3] ), .b(
        \U1664/x[2] ), .c(\U1664/x[3] ), .d(\U1664/U30/Z ), .e(\U1664/x[2] ), 
        .f(\U1664/U30/Z ) );
    inv_1 \U1664/U30/U30/Uinv  ( .x(\U1664/U30/Z ), .a(\U1664/y[1] ) );
    aoi222_1 \U1664/U31/U30/U1  ( .x(\U1664/x[1] ), .a(\ncd[3] ), .b(\ncd[2] ), 
        .c(\ncd[3] ), .d(\U1664/U31/Z ), .e(\ncd[2] ), .f(\U1664/U31/Z ) );
    inv_1 \U1664/U31/U30/Uinv  ( .x(\U1664/U31/Z ), .a(\U1664/x[1] ) );
    aoi222_1 \U1664/U37/U30/U1  ( .x(pullcd), .a(\U1664/y[0] ), .b(
        \U1664/y[1] ), .c(\U1664/y[0] ), .d(\U1664/U37/Z ), .e(\U1664/y[1] ), 
        .f(\U1664/U37/Z ) );
    inv_1 \U1664/U37/U30/Uinv  ( .x(\U1664/U37/Z ), .a(pullcd) );
    nor3_1 \U1697/U21/Unr  ( .x(\U1697/U21/nr ), .a(rnw[0]), .b(pkt_normal), 
        .c(net149) );
    nand3_1 \U1697/U21/Und  ( .x(\U1697/U21/nd ), .a(rnw[0]), .b(pkt_normal), 
        .c(net149) );
    oa21_1 \U1697/U21/U1  ( .x(\U1697/U21/n2 ), .a(\U1697/U21/n2 ), .b(
        \U1697/U21/nr ), .c(\U1697/U21/nd ) );
    inv_1 \U1697/U21/U3  ( .x(write), .a(\U1697/U21/n2 ) );
    nor3_1 \U307/U21/Unr  ( .x(\U307/U21/nr ), .a(net149), .b(net150), .c(
        statusack) );
    nand3_1 \U307/U21/Und  ( .x(\U307/U21/nd ), .a(net149), .b(net150), .c(
        statusack) );
    oa21_1 \U307/U21/U1  ( .x(\U307/U21/n2 ), .a(\U307/U21/n2 ), .b(
        \U307/U21/nr ), .c(\U307/U21/nd ) );
    inv_1 \U307/U21/U3  ( .x(notify), .a(\U307/U21/n2 ) );
    nor3_1 \U1698/Unr  ( .x(\U1698/nr ), .a(rnw[1]), .b(pkt_normal), .c(net149
        ) );
    nand3_1 \U1698/Und  ( .x(\U1698/nd ), .a(rnw[1]), .b(pkt_normal), .c(
        net149) );
    oa21_1 \U1698/U1  ( .x(\U1698/n2 ), .a(\U1698/n2 ), .b(\U1698/nr ), .c(
        \U1698/nd ) );
    inv_2 \U1698/U3  ( .x(read), .a(\U1698/n2 ) );
    and2_1 \U1756/U1754/U8  ( .x(n17), .a(\opc_h[0] ), .b(pkt_normal) );
    and2_1 \U1756/U1755/U8  ( .x(n18), .a(\opc_l[0] ), .b(pkt_normal) );
    and2_1 \U1800/U1754/U8  ( .x(rnw[1]), .a(net0187), .b(pkt_normal) );
    and2_1 \U1800/U1755/U8  ( .x(rnw[0]), .a(net0208), .b(pkt_normal) );
    and2_1 \U1758/U1754/U8  ( .x(status[1]), .a(\opc_h[0] ), .b(net150) );
    and2_1 \U1758/U1755/U8  ( .x(status[0]), .a(\opc_l[0] ), .b(net150) );
    buf_2 \I6/U1653  ( .x(\I6/latch ), .a(net173) );
    nor2_1 \I6/U264/U5  ( .x(\I6/nlocalcd ), .a(reset), .b(\I6/localcd ) );
    nor2_1 \I6/U1659_0_/U5  ( .x(\I6/ncd[0] ), .a(\opc_l[0] ), .b(\opc_h[0] )
         );
    nor2_1 \I6/U1659_1_/U5  ( .x(\I6/ncd[1] ), .a(\opc_l[1] ), .b(\opc_h[1] )
         );
    nor2_1 \I6/U1659_2_/U5  ( .x(\I6/ncd[2] ), .a(\opc_l[2] ), .b(\I6/oh[2] )
         );
    nor2_1 \I6/U1659_3_/U5  ( .x(\I6/ncd[3] ), .a(\I6/ol[3] ), .b(\I6/oh[3] )
         );
    nor2_1 \I6/U1659_4_/U5  ( .x(\I6/ncd[4] ), .a(\I6/ol[4] ), .b(\I6/oh[4] )
         );
    nor2_1 \I6/U1659_5_/U5  ( .x(\I6/ncd[5] ), .a(net0208), .b(net0187) );
    nor2_1 \I6/U1659_6_/U5  ( .x(\I6/ncd[6] ), .a(\I6/ol[6] ), .b(\I6/oh[6] )
         );
    nor2_1 \I6/U1659_7_/U5  ( .x(\I6/ncd[7] ), .a(\I6/ol[7] ), .b(\I6/oh[7] )
         );
    nor2_1 \I6/U3/U5  ( .x(\I6/ctrlack_internal ), .a(\I6/acb ), .b(\I6/ba )
         );
    buf_2 \I6/U1665/U7  ( .x(\I6/driveh ), .a(net139) );
    buf_2 \I6/U1666/U7  ( .x(\I6/drivel ), .a(net139) );
    ao23_1 \I6/U1658_0_/U21/U1/U1  ( .x(\opc_l[0] ), .a(\I6/driveh ), .b(
        \opc_l[0] ), .c(\I6/driveh ), .d(cbl[0]), .e(n12) );
    ao23_1 \I6/U1658_1_/U21/U1/U1  ( .x(\opc_l[1] ), .a(\I6/driveh ), .b(
        \opc_l[1] ), .c(\I6/drivel ), .d(cbl[1]), .e(n12) );
    ao23_1 \I6/U1658_2_/U21/U1/U1  ( .x(\opc_l[2] ), .a(\I6/drivel ), .b(
        \opc_l[2] ), .c(n13), .d(cbl[2]), .e(n12) );
    ao23_1 \I6/U1658_3_/U21/U1/U1  ( .x(\I6/ol[3] ), .a(\I6/drivel ), .b(
        \I6/ol[3] ), .c(\I6/drivel ), .d(cbl[3]), .e(\I6/latch ) );
    ao23_1 \I6/U1658_4_/U21/U1/U1  ( .x(\I6/ol[4] ), .a(n13), .b(\I6/ol[4] ), 
        .c(n13), .d(cbl[4]), .e(\I6/latch ) );
    ao23_1 \I6/U1658_5_/U21/U1/U1  ( .x(net0208), .a(\I6/driveh ), .b(net0208), 
        .c(\I6/driveh ), .d(cbl[5]), .e(\I6/latch ) );
    ao23_1 \I6/U1658_6_/U21/U1/U1  ( .x(\I6/ol[6] ), .a(n13), .b(\I6/ol[6] ), 
        .c(n13), .d(cbl[6]), .e(\I6/latch ) );
    ao23_1 \I6/U1658_7_/U21/U1/U1  ( .x(\I6/ol[7] ), .a(n13), .b(\I6/ol[7] ), 
        .c(\I6/driveh ), .d(cbl[7]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_0_/U21/U1/U1  ( .x(\opc_h[0] ), .a(n13), .b(\opc_h[0] ), 
        .c(\I6/drivel ), .d(cbh[0]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_1_/U21/U1/U1  ( .x(\opc_h[1] ), .a(\I6/driveh ), .b(
        \opc_h[1] ), .c(n13), .d(cbh[1]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_2_/U21/U1/U1  ( .x(\I6/oh[2] ), .a(\I6/driveh ), .b(
        \I6/oh[2] ), .c(n13), .d(cbh[2]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_3_/U21/U1/U1  ( .x(\I6/oh[3] ), .a(\I6/drivel ), .b(
        \I6/oh[3] ), .c(\I6/drivel ), .d(cbh[3]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_4_/U21/U1/U1  ( .x(\I6/oh[4] ), .a(n13), .b(\I6/oh[4] ), 
        .c(\I6/driveh ), .d(cbh[4]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_5_/U21/U1/U1  ( .x(net0187), .a(\I6/driveh ), .b(net0187), 
        .c(\I6/driveh ), .d(cbh[5]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_6_/U21/U1/U1  ( .x(\I6/oh[6] ), .a(\I6/drivel ), .b(
        \I6/oh[6] ), .c(\I6/drivel ), .d(cbh[6]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_7_/U21/U1/U1  ( .x(\I6/oh[7] ), .a(\I6/drivel ), .b(
        \I6/oh[7] ), .c(n13), .d(cbh[7]), .e(\I6/latch ) );
    aoai211_1 \I6/U4/U28/U1/U1  ( .x(\I6/U4/U28/U1/clr ), .a(net139), .b(
        \I6/acb ), .c(\I6/nlocalcd ), .d(net173) );
    nand3_1 \I6/U4/U28/U1/U2  ( .x(\I6/U4/U28/U1/set ), .a(\I6/nlocalcd ), .b(
        net139), .c(\I6/acb ) );
    nand2_2 \I6/U4/U28/U1/U3  ( .x(net173), .a(\I6/U4/U28/U1/clr ), .b(
        \I6/U4/U28/U1/set ) );
    oai21_1 \I6/U1/U30/U1/U1  ( .x(\I6/acb ), .a(\I6/U1/Z ), .b(\I6/ba ), .c(
        net139) );
    inv_1 \I6/U1/U30/U1/U2  ( .x(\I6/U1/Z ), .a(\I6/acb ) );
    ao222_1 \I6/U5/U18/U1/U1  ( .x(\I6/ba ), .a(\I6/latch ), .b(n14), .c(
        \I6/latch ), .d(\I6/ba ), .e(n14), .f(\I6/ba ) );
    aoi222_1 \I6/U1664/U28/U30/U1  ( .x(\I6/U1664/x[3] ), .a(\I6/ncd[7] ), .b(
        \I6/ncd[6] ), .c(\I6/ncd[7] ), .d(\I6/U1664/U28/Z ), .e(\I6/ncd[6] ), 
        .f(\I6/U1664/U28/Z ) );
    inv_1 \I6/U1664/U28/U30/Uinv  ( .x(\I6/U1664/U28/Z ), .a(\I6/U1664/x[3] )
         );
    aoi222_1 \I6/U1664/U32/U30/U1  ( .x(\I6/U1664/x[0] ), .a(\I6/ncd[1] ), .b(
        \I6/ncd[0] ), .c(\I6/ncd[1] ), .d(\I6/U1664/U32/Z ), .e(\I6/ncd[0] ), 
        .f(\I6/U1664/U32/Z ) );
    inv_1 \I6/U1664/U32/U30/Uinv  ( .x(\I6/U1664/U32/Z ), .a(\I6/U1664/x[0] )
         );
    aoi222_1 \I6/U1664/U29/U30/U1  ( .x(\I6/U1664/x[2] ), .a(\I6/ncd[5] ), .b(
        \I6/ncd[4] ), .c(\I6/ncd[5] ), .d(\I6/U1664/U29/Z ), .e(\I6/ncd[4] ), 
        .f(\I6/U1664/U29/Z ) );
    inv_1 \I6/U1664/U29/U30/Uinv  ( .x(\I6/U1664/U29/Z ), .a(\I6/U1664/x[2] )
         );
    aoi222_1 \I6/U1664/U33/U30/U1  ( .x(\I6/U1664/y[0] ), .a(\I6/U1664/x[1] ), 
        .b(\I6/U1664/x[0] ), .c(\I6/U1664/x[1] ), .d(\I6/U1664/U33/Z ), .e(
        \I6/U1664/x[0] ), .f(\I6/U1664/U33/Z ) );
    inv_1 \I6/U1664/U33/U30/Uinv  ( .x(\I6/U1664/U33/Z ), .a(\I6/U1664/y[0] )
         );
    aoi222_1 \I6/U1664/U30/U30/U1  ( .x(\I6/U1664/y[1] ), .a(\I6/U1664/x[3] ), 
        .b(\I6/U1664/x[2] ), .c(\I6/U1664/x[3] ), .d(\I6/U1664/U30/Z ), .e(
        \I6/U1664/x[2] ), .f(\I6/U1664/U30/Z ) );
    inv_1 \I6/U1664/U30/U30/Uinv  ( .x(\I6/U1664/U30/Z ), .a(\I6/U1664/y[1] )
         );
    aoi222_1 \I6/U1664/U31/U30/U1  ( .x(\I6/U1664/x[1] ), .a(\I6/ncd[3] ), .b(
        \I6/ncd[2] ), .c(\I6/ncd[3] ), .d(\I6/U1664/U31/Z ), .e(\I6/ncd[2] ), 
        .f(\I6/U1664/U31/Z ) );
    inv_1 \I6/U1664/U31/U30/Uinv  ( .x(\I6/U1664/U31/Z ), .a(\I6/U1664/x[1] )
         );
    aoi222_1 \I6/U1664/U37/U30/U1  ( .x(\I6/localcd ), .a(\I6/U1664/y[0] ), 
        .b(\I6/U1664/y[1] ), .c(\I6/U1664/y[0] ), .d(\I6/U1664/U37/Z ), .e(
        \I6/U1664/y[1] ), .f(\I6/U1664/U37/Z ) );
    inv_1 \I6/U1664/U37/U30/Uinv  ( .x(\I6/U1664/U37/Z ), .a(\I6/localcd ) );
    nor3_1 \I6/U1669/Unr  ( .x(\I6/U1669/nr ), .a(\I6/ctrlack_internal ), .b(
        n13), .c(\I6/drivel ) );
    nand3_1 \I6/U1669/Und  ( .x(\I6/U1669/nd ), .a(\I6/ctrlack_internal ), .b(
        \I6/driveh ), .c(\I6/drivel ) );
    oa21_1 \I6/U1669/U1  ( .x(\I6/U1669/n2 ), .a(\I6/U1669/n2 ), .b(
        \I6/U1669/nr ), .c(\I6/U1669/nd ) );
    inv_2 \I6/U1669/U3  ( .x(net149), .a(\I6/U1669/n2 ) );
    buf_2 \U1667/U1653  ( .x(\U1667/latch ), .a(net167) );
    nor2_1 \U1667/U264/U5  ( .x(\U1667/nlocalcd ), .a(reset), .b(
        \U1667/localcd ) );
    nor2_1 \U1667/U1659_0_/U5  ( .x(\U1667/ncd[0] ), .a(rd[0]), .b(rd[32]) );
    nor2_1 \U1667/U1659_1_/U5  ( .x(\U1667/ncd[1] ), .a(rd[1]), .b(rd[33]) );
    nor2_1 \U1667/U1659_2_/U5  ( .x(\U1667/ncd[2] ), .a(rd[2]), .b(rd[34]) );
    nor2_1 \U1667/U1659_3_/U5  ( .x(\U1667/ncd[3] ), .a(rd[3]), .b(rd[35]) );
    nor2_1 \U1667/U1659_4_/U5  ( .x(\U1667/ncd[4] ), .a(rd[4]), .b(rd[36]) );
    nor2_1 \U1667/U1659_5_/U5  ( .x(\U1667/ncd[5] ), .a(rd[5]), .b(rd[37]) );
    nor2_1 \U1667/U1659_6_/U5  ( .x(\U1667/ncd[6] ), .a(rd[6]), .b(rd[38]) );
    nor2_1 \U1667/U1659_7_/U5  ( .x(\U1667/ncd[7] ), .a(rd[7]), .b(rd[39]) );
    nor2_1 \U1667/U3/U5  ( .x(\U1667/ctrlack_internal ), .a(\U1667/acb ), .b(
        \U1667/ba ) );
    buf_2 \U1667/U1665/U7  ( .x(\U1667/driveh ), .a(read_lhw) );
    buf_2 \U1667/U1666/U7  ( .x(\U1667/drivel ), .a(read_lhw) );
    ao23_1 \U1667/U1658_0_/U21/U1/U1  ( .x(rd[0]), .a(n11), .b(rd[0]), .c(
        \U1667/drivel ), .d(cbl[0]), .e(n10) );
    ao23_1 \U1667/U1658_1_/U21/U1/U1  ( .x(rd[1]), .a(n11), .b(rd[1]), .c(
        \U1667/driveh ), .d(cbl[1]), .e(n10) );
    ao23_1 \U1667/U1658_2_/U21/U1/U1  ( .x(rd[2]), .a(\U1667/driveh ), .b(rd
        [2]), .c(n11), .d(cbl[2]), .e(n10) );
    ao23_1 \U1667/U1658_3_/U21/U1/U1  ( .x(rd[3]), .a(n11), .b(rd[3]), .c(
        \U1667/driveh ), .d(cbl[3]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1658_4_/U21/U1/U1  ( .x(rd[4]), .a(\U1667/drivel ), .b(rd
        [4]), .c(n11), .d(cbl[4]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1658_5_/U21/U1/U1  ( .x(rd[5]), .a(\U1667/drivel ), .b(rd
        [5]), .c(n11), .d(cbl[5]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1658_6_/U21/U1/U1  ( .x(rd[6]), .a(\U1667/driveh ), .b(rd
        [6]), .c(\U1667/drivel ), .d(cbl[6]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1658_7_/U21/U1/U1  ( .x(rd[7]), .a(\U1667/driveh ), .b(rd
        [7]), .c(\U1667/driveh ), .d(cbl[7]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_0_/U21/U1/U1  ( .x(rd[32]), .a(\U1667/drivel ), .b(rd
        [32]), .c(n11), .d(cbh[0]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_1_/U21/U1/U1  ( .x(rd[33]), .a(\U1667/driveh ), .b(rd
        [33]), .c(\U1667/drivel ), .d(cbh[1]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_2_/U21/U1/U1  ( .x(rd[34]), .a(\U1667/drivel ), .b(rd
        [34]), .c(\U1667/drivel ), .d(cbh[2]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_3_/U21/U1/U1  ( .x(rd[35]), .a(\U1667/driveh ), .b(rd
        [35]), .c(\U1667/driveh ), .d(cbh[3]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_4_/U21/U1/U1  ( .x(rd[36]), .a(\U1667/drivel ), .b(rd
        [36]), .c(\U1667/driveh ), .d(cbh[4]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_5_/U21/U1/U1  ( .x(rd[37]), .a(\U1667/driveh ), .b(rd
        [37]), .c(n11), .d(cbh[5]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_6_/U21/U1/U1  ( .x(rd[38]), .a(n11), .b(rd[38]), .c(
        \U1667/drivel ), .d(cbh[6]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_7_/U21/U1/U1  ( .x(rd[39]), .a(n11), .b(rd[39]), .c(
        n11), .d(cbh[7]), .e(\U1667/latch ) );
    aoai211_1 \U1667/U4/U28/U1/U1  ( .x(\U1667/U4/U28/U1/clr ), .a(read_lhw), 
        .b(\U1667/acb ), .c(\U1667/nlocalcd ), .d(net167) );
    nand3_1 \U1667/U4/U28/U1/U2  ( .x(\U1667/U4/U28/U1/set ), .a(
        \U1667/nlocalcd ), .b(read_lhw), .c(\U1667/acb ) );
    nand2_2 \U1667/U4/U28/U1/U3  ( .x(net167), .a(\U1667/U4/U28/U1/clr ), .b(
        \U1667/U4/U28/U1/set ) );
    oai21_1 \U1667/U1/U30/U1/U1  ( .x(\U1667/acb ), .a(\U1667/U1/Z ), .b(
        \U1667/ba ), .c(read_lhw) );
    inv_1 \U1667/U1/U30/U1/U2  ( .x(\U1667/U1/Z ), .a(\U1667/acb ) );
    ao222_1 \U1667/U5/U18/U1/U1  ( .x(\U1667/ba ), .a(\U1667/latch ), .b(n14), 
        .c(\U1667/latch ), .d(\U1667/ba ), .e(n14), .f(\U1667/ba ) );
    aoi222_1 \U1667/U1664/U28/U30/U1  ( .x(\U1667/U1664/x[3] ), .a(
        \U1667/ncd[7] ), .b(\U1667/ncd[6] ), .c(\U1667/ncd[7] ), .d(
        \U1667/U1664/U28/Z ), .e(\U1667/ncd[6] ), .f(\U1667/U1664/U28/Z ) );
    inv_1 \U1667/U1664/U28/U30/Uinv  ( .x(\U1667/U1664/U28/Z ), .a(
        \U1667/U1664/x[3] ) );
    aoi222_1 \U1667/U1664/U32/U30/U1  ( .x(\U1667/U1664/x[0] ), .a(
        \U1667/ncd[1] ), .b(\U1667/ncd[0] ), .c(\U1667/ncd[1] ), .d(
        \U1667/U1664/U32/Z ), .e(\U1667/ncd[0] ), .f(\U1667/U1664/U32/Z ) );
    inv_1 \U1667/U1664/U32/U30/Uinv  ( .x(\U1667/U1664/U32/Z ), .a(
        \U1667/U1664/x[0] ) );
    aoi222_1 \U1667/U1664/U29/U30/U1  ( .x(\U1667/U1664/x[2] ), .a(
        \U1667/ncd[5] ), .b(\U1667/ncd[4] ), .c(\U1667/ncd[5] ), .d(
        \U1667/U1664/U29/Z ), .e(\U1667/ncd[4] ), .f(\U1667/U1664/U29/Z ) );
    inv_1 \U1667/U1664/U29/U30/Uinv  ( .x(\U1667/U1664/U29/Z ), .a(
        \U1667/U1664/x[2] ) );
    aoi222_1 \U1667/U1664/U33/U30/U1  ( .x(\U1667/U1664/y[0] ), .a(
        \U1667/U1664/x[1] ), .b(\U1667/U1664/x[0] ), .c(\U1667/U1664/x[1] ), 
        .d(\U1667/U1664/U33/Z ), .e(\U1667/U1664/x[0] ), .f(
        \U1667/U1664/U33/Z ) );
    inv_1 \U1667/U1664/U33/U30/Uinv  ( .x(\U1667/U1664/U33/Z ), .a(
        \U1667/U1664/y[0] ) );
    aoi222_1 \U1667/U1664/U30/U30/U1  ( .x(\U1667/U1664/y[1] ), .a(
        \U1667/U1664/x[3] ), .b(\U1667/U1664/x[2] ), .c(\U1667/U1664/x[3] ), 
        .d(\U1667/U1664/U30/Z ), .e(\U1667/U1664/x[2] ), .f(
        \U1667/U1664/U30/Z ) );
    inv_1 \U1667/U1664/U30/U30/Uinv  ( .x(\U1667/U1664/U30/Z ), .a(
        \U1667/U1664/y[1] ) );
    aoi222_1 \U1667/U1664/U31/U30/U1  ( .x(\U1667/U1664/x[1] ), .a(
        \U1667/ncd[3] ), .b(\U1667/ncd[2] ), .c(\U1667/ncd[3] ), .d(
        \U1667/U1664/U31/Z ), .e(\U1667/ncd[2] ), .f(\U1667/U1664/U31/Z ) );
    inv_1 \U1667/U1664/U31/U30/Uinv  ( .x(\U1667/U1664/U31/Z ), .a(
        \U1667/U1664/x[1] ) );
    aoi222_1 \U1667/U1664/U37/U30/U1  ( .x(\U1667/localcd ), .a(
        \U1667/U1664/y[0] ), .b(\U1667/U1664/y[1] ), .c(\U1667/U1664/y[0] ), 
        .d(\U1667/U1664/U37/Z ), .e(\U1667/U1664/y[1] ), .f(
        \U1667/U1664/U37/Z ) );
    inv_1 \U1667/U1664/U37/U30/Uinv  ( .x(\U1667/U1664/U37/Z ), .a(
        \U1667/localcd ) );
    nor3_1 \U1667/U1669/Unr  ( .x(\U1667/U1669/nr ), .a(
        \U1667/ctrlack_internal ), .b(n11), .c(\U1667/drivel ) );
    nand3_1 \U1667/U1669/Und  ( .x(\U1667/U1669/nd ), .a(
        \U1667/ctrlack_internal ), .b(\U1667/driveh ), .c(\U1667/drivel ) );
    oa21_1 \U1667/U1669/U1  ( .x(\U1667/U1669/n2 ), .a(\U1667/U1669/n2 ), .b(
        \U1667/U1669/nr ), .c(\U1667/U1669/nd ) );
    inv_2 \U1667/U1669/U3  ( .x(net193), .a(\U1667/U1669/n2 ) );
    buf_2 \U1650/U1653  ( .x(\U1650/latch ), .a(net172) );
    nor2_1 \U1650/U264/U5  ( .x(\U1650/nlocalcd ), .a(reset), .b(
        \U1650/localcd ) );
    nor2_1 \U1650/U1659_0_/U5  ( .x(\U1650/ncd[0] ), .a(\U1650/ol[0] ), .b(
        \U1650/oh[0] ) );
    nor2_1 \U1650/U1659_1_/U5  ( .x(\U1650/ncd[1] ), .a(\U1650/ol[1] ), .b(
        \U1650/oh[1] ) );
    nor2_1 \U1650/U1659_2_/U5  ( .x(\U1650/ncd[2] ), .a(\U1650/ol[2] ), .b(
        \U1650/oh[2] ) );
    nor2_1 \U1650/U1659_3_/U5  ( .x(\U1650/ncd[3] ), .a(\U1650/ol[3] ), .b(
        \U1650/oh[3] ) );
    nor2_1 \U1650/U1659_4_/U5  ( .x(\U1650/ncd[4] ), .a(\U1650/ol[4] ), .b(
        \U1650/oh[4] ) );
    nor2_1 \U1650/U1659_5_/U5  ( .x(\U1650/ncd[5] ), .a(\col_l[0] ), .b(
        \col_h[0] ) );
    nor2_1 \U1650/U1659_6_/U5  ( .x(\U1650/ncd[6] ), .a(\col_l[1] ), .b(
        \col_h[1] ) );
    nor2_1 \U1650/U1659_7_/U5  ( .x(\U1650/ncd[7] ), .a(\col_l[2] ), .b(
        \col_h[2] ) );
    nor2_1 \U1650/U3/U5  ( .x(\U1650/ctrlack_internal ), .a(\U1650/acb ), .b(
        \U1650/ba ) );
    buf_2 \U1650/U1665/U7  ( .x(\U1650/driveh ), .a(start_receiving) );
    buf_2 \U1650/U1666/U7  ( .x(\U1650/drivel ), .a(start_receiving) );
    ao23_1 \U1650/U1658_0_/U21/U1/U1  ( .x(\U1650/ol[0] ), .a(\U1650/drivel ), 
        .b(\U1650/ol[0] ), .c(\U1650/drivel ), .d(cbl[0]), .e(n7) );
    ao23_1 \U1650/U1658_1_/U21/U1/U1  ( .x(\U1650/ol[1] ), .a(\U1650/drivel ), 
        .b(\U1650/ol[1] ), .c(\U1650/drivel ), .d(cbl[1]), .e(n7) );
    ao23_1 \U1650/U1658_2_/U21/U1/U1  ( .x(\U1650/ol[2] ), .a(\U1650/drivel ), 
        .b(\U1650/ol[2] ), .c(\U1650/drivel ), .d(cbl[2]), .e(n7) );
    ao23_1 \U1650/U1658_3_/U21/U1/U1  ( .x(\U1650/ol[3] ), .a(n9), .b(
        \U1650/ol[3] ), .c(\U1650/drivel ), .d(cbl[3]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1658_4_/U21/U1/U1  ( .x(\U1650/ol[4] ), .a(\U1650/drivel ), 
        .b(\U1650/ol[4] ), .c(\U1650/drivel ), .d(cbl[4]), .e(\U1650/latch )
         );
    ao23_1 \U1650/U1658_5_/U21/U1/U1  ( .x(\col_l[0] ), .a(\U1650/drivel ), 
        .b(\col_l[0] ), .c(\U1650/drivel ), .d(cbl[5]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1658_6_/U21/U1/U1  ( .x(\col_l[1] ), .a(n9), .b(\col_l[1] ), 
        .c(\U1650/drivel ), .d(cbl[6]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1658_7_/U21/U1/U1  ( .x(\col_l[2] ), .a(n9), .b(\col_l[2] ), 
        .c(\U1650/drivel ), .d(cbl[7]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1651_0_/U21/U1/U1  ( .x(\U1650/oh[0] ), .a(\U1650/driveh ), 
        .b(\U1650/oh[0] ), .c(\U1650/driveh ), .d(cbh[0]), .e(\U1650/latch )
         );
    ao23_1 \U1650/U1651_1_/U21/U1/U1  ( .x(\U1650/oh[1] ), .a(\U1650/driveh ), 
        .b(\U1650/oh[1] ), .c(\U1650/driveh ), .d(cbh[1]), .e(\U1650/latch )
         );
    ao23_1 \U1650/U1651_2_/U21/U1/U1  ( .x(\U1650/oh[2] ), .a(\U1650/driveh ), 
        .b(\U1650/oh[2] ), .c(\U1650/driveh ), .d(cbh[2]), .e(\U1650/latch )
         );
    ao23_1 \U1650/U1651_3_/U21/U1/U1  ( .x(\U1650/oh[3] ), .a(n8), .b(
        \U1650/oh[3] ), .c(\U1650/driveh ), .d(cbh[3]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1651_4_/U21/U1/U1  ( .x(\U1650/oh[4] ), .a(n8), .b(
        \U1650/oh[4] ), .c(\U1650/driveh ), .d(cbh[4]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1651_5_/U21/U1/U1  ( .x(\col_h[0] ), .a(\U1650/driveh ), 
        .b(\col_h[0] ), .c(\U1650/driveh ), .d(cbh[5]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1651_6_/U21/U1/U1  ( .x(\col_h[1] ), .a(n8), .b(\col_h[1] ), 
        .c(\U1650/driveh ), .d(cbh[6]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1651_7_/U21/U1/U1  ( .x(\col_h[2] ), .a(\U1650/driveh ), 
        .b(\col_h[2] ), .c(\U1650/driveh ), .d(cbh[7]), .e(\U1650/latch ) );
    aoai211_1 \U1650/U4/U28/U1/U1  ( .x(\U1650/U4/U28/U1/clr ), .a(
        start_receiving), .b(\U1650/acb ), .c(\U1650/nlocalcd ), .d(net172) );
    nand3_1 \U1650/U4/U28/U1/U2  ( .x(\U1650/U4/U28/U1/set ), .a(
        \U1650/nlocalcd ), .b(start_receiving), .c(\U1650/acb ) );
    nand2_2 \U1650/U4/U28/U1/U3  ( .x(net172), .a(\U1650/U4/U28/U1/clr ), .b(
        \U1650/U4/U28/U1/set ) );
    oai21_1 \U1650/U1/U30/U1/U1  ( .x(\U1650/acb ), .a(\U1650/U1/Z ), .b(
        \U1650/ba ), .c(start_receiving) );
    inv_1 \U1650/U1/U30/U1/U2  ( .x(\U1650/U1/Z ), .a(\U1650/acb ) );
    ao222_1 \U1650/U5/U18/U1/U1  ( .x(\U1650/ba ), .a(\U1650/latch ), .b(n14), 
        .c(\U1650/latch ), .d(\U1650/ba ), .e(n14), .f(\U1650/ba ) );
    aoi222_1 \U1650/U1664/U28/U30/U1  ( .x(\U1650/U1664/x[3] ), .a(
        \U1650/ncd[7] ), .b(\U1650/ncd[6] ), .c(\U1650/ncd[7] ), .d(
        \U1650/U1664/U28/Z ), .e(\U1650/ncd[6] ), .f(\U1650/U1664/U28/Z ) );
    inv_1 \U1650/U1664/U28/U30/Uinv  ( .x(\U1650/U1664/U28/Z ), .a(
        \U1650/U1664/x[3] ) );
    aoi222_1 \U1650/U1664/U32/U30/U1  ( .x(\U1650/U1664/x[0] ), .a(
        \U1650/ncd[1] ), .b(\U1650/ncd[0] ), .c(\U1650/ncd[1] ), .d(
        \U1650/U1664/U32/Z ), .e(\U1650/ncd[0] ), .f(\U1650/U1664/U32/Z ) );
    inv_1 \U1650/U1664/U32/U30/Uinv  ( .x(\U1650/U1664/U32/Z ), .a(
        \U1650/U1664/x[0] ) );
    aoi222_1 \U1650/U1664/U29/U30/U1  ( .x(\U1650/U1664/x[2] ), .a(
        \U1650/ncd[5] ), .b(\U1650/ncd[4] ), .c(\U1650/ncd[5] ), .d(
        \U1650/U1664/U29/Z ), .e(\U1650/ncd[4] ), .f(\U1650/U1664/U29/Z ) );
    inv_1 \U1650/U1664/U29/U30/Uinv  ( .x(\U1650/U1664/U29/Z ), .a(
        \U1650/U1664/x[2] ) );
    aoi222_1 \U1650/U1664/U33/U30/U1  ( .x(\U1650/U1664/y[0] ), .a(
        \U1650/U1664/x[1] ), .b(\U1650/U1664/x[0] ), .c(\U1650/U1664/x[1] ), 
        .d(\U1650/U1664/U33/Z ), .e(\U1650/U1664/x[0] ), .f(
        \U1650/U1664/U33/Z ) );
    inv_1 \U1650/U1664/U33/U30/Uinv  ( .x(\U1650/U1664/U33/Z ), .a(
        \U1650/U1664/y[0] ) );
    aoi222_1 \U1650/U1664/U30/U30/U1  ( .x(\U1650/U1664/y[1] ), .a(
        \U1650/U1664/x[3] ), .b(\U1650/U1664/x[2] ), .c(\U1650/U1664/x[3] ), 
        .d(\U1650/U1664/U30/Z ), .e(\U1650/U1664/x[2] ), .f(
        \U1650/U1664/U30/Z ) );
    inv_1 \U1650/U1664/U30/U30/Uinv  ( .x(\U1650/U1664/U30/Z ), .a(
        \U1650/U1664/y[1] ) );
    aoi222_1 \U1650/U1664/U31/U30/U1  ( .x(\U1650/U1664/x[1] ), .a(
        \U1650/ncd[3] ), .b(\U1650/ncd[2] ), .c(\U1650/ncd[3] ), .d(
        \U1650/U1664/U31/Z ), .e(\U1650/ncd[2] ), .f(\U1650/U1664/U31/Z ) );
    inv_1 \U1650/U1664/U31/U30/Uinv  ( .x(\U1650/U1664/U31/Z ), .a(
        \U1650/U1664/x[1] ) );
    aoi222_1 \U1650/U1664/U37/U30/U1  ( .x(\U1650/localcd ), .a(
        \U1650/U1664/y[0] ), .b(\U1650/U1664/y[1] ), .c(\U1650/U1664/y[0] ), 
        .d(\U1650/U1664/U37/Z ), .e(\U1650/U1664/y[1] ), .f(
        \U1650/U1664/U37/Z ) );
    inv_1 \U1650/U1664/U37/U30/Uinv  ( .x(\U1650/U1664/U37/Z ), .a(
        \U1650/localcd ) );
    nor3_1 \U1650/U1669/Unr  ( .x(\U1650/U1669/nr ), .a(
        \U1650/ctrlack_internal ), .b(\U1650/drivel ), .c(\U1650/driveh ) );
    nand3_1 \U1650/U1669/Und  ( .x(\U1650/U1669/nd ), .a(
        \U1650/ctrlack_internal ), .b(\U1650/drivel ), .c(\U1650/driveh ) );
    oa21_1 \U1650/U1669/U1  ( .x(\U1650/U1669/n2 ), .a(\U1650/U1669/n2 ), .b(
        \U1650/U1669/nr ), .c(\U1650/U1669/nd ) );
    inv_2 \U1650/U1669/U3  ( .x(net139), .a(\U1650/U1669/n2 ) );
    buf_2 \U1666/U1653  ( .x(\U1666/latch ), .a(net169) );
    nor2_1 \U1666/U264/U5  ( .x(\U1666/nlocalcd ), .a(reset), .b(
        \U1666/localcd ) );
    nor2_1 \U1666/U1659_0_/U5  ( .x(\U1666/ncd[0] ), .a(rd[24]), .b(rd[56]) );
    nor2_1 \U1666/U1659_1_/U5  ( .x(\U1666/ncd[1] ), .a(rd[25]), .b(rd[57]) );
    nor2_1 \U1666/U1659_2_/U5  ( .x(\U1666/ncd[2] ), .a(rd[26]), .b(rd[58]) );
    nor2_1 \U1666/U1659_3_/U5  ( .x(\U1666/ncd[3] ), .a(rd[27]), .b(rd[59]) );
    nor2_1 \U1666/U1659_4_/U5  ( .x(\U1666/ncd[4] ), .a(rd[28]), .b(rd[60]) );
    nor2_1 \U1666/U1659_5_/U5  ( .x(\U1666/ncd[5] ), .a(rd[29]), .b(rd[61]) );
    nor2_1 \U1666/U1659_6_/U5  ( .x(\U1666/ncd[6] ), .a(rd[30]), .b(rd[62]) );
    nor2_1 \U1666/U1659_7_/U5  ( .x(\U1666/ncd[7] ), .a(rd[31]), .b(rd[63]) );
    nor2_1 \U1666/U3/U5  ( .x(\U1666/ctrlack_internal ), .a(\U1666/acb ), .b(
        \U1666/ba ) );
    buf_2 \U1666/U1665/U7  ( .x(\U1666/driveh ), .a(read) );
    buf_2 \U1666/U1666/U7  ( .x(\U1666/drivel ), .a(read) );
    ao23_1 \U1666/U1658_0_/U21/U1/U1  ( .x(rd[24]), .a(n6), .b(rd[24]), .c(
        \U1666/drivel ), .d(cbl[0]), .e(n5) );
    ao23_1 \U1666/U1658_1_/U21/U1/U1  ( .x(rd[25]), .a(n6), .b(rd[25]), .c(
        \U1666/driveh ), .d(cbl[1]), .e(n5) );
    ao23_1 \U1666/U1658_2_/U21/U1/U1  ( .x(rd[26]), .a(\U1666/driveh ), .b(rd
        [26]), .c(n6), .d(cbl[2]), .e(n5) );
    ao23_1 \U1666/U1658_3_/U21/U1/U1  ( .x(rd[27]), .a(n6), .b(rd[27]), .c(
        \U1666/driveh ), .d(cbl[3]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1658_4_/U21/U1/U1  ( .x(rd[28]), .a(\U1666/drivel ), .b(rd
        [28]), .c(n6), .d(cbl[4]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1658_5_/U21/U1/U1  ( .x(rd[29]), .a(\U1666/drivel ), .b(rd
        [29]), .c(n6), .d(cbl[5]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1658_6_/U21/U1/U1  ( .x(rd[30]), .a(\U1666/driveh ), .b(rd
        [30]), .c(\U1666/drivel ), .d(cbl[6]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1658_7_/U21/U1/U1  ( .x(rd[31]), .a(\U1666/driveh ), .b(rd
        [31]), .c(\U1666/driveh ), .d(cbl[7]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_0_/U21/U1/U1  ( .x(rd[56]), .a(\U1666/drivel ), .b(rd
        [56]), .c(n6), .d(cbh[0]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_1_/U21/U1/U1  ( .x(rd[57]), .a(\U1666/driveh ), .b(rd
        [57]), .c(\U1666/drivel ), .d(cbh[1]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_2_/U21/U1/U1  ( .x(rd[58]), .a(\U1666/drivel ), .b(rd
        [58]), .c(\U1666/drivel ), .d(cbh[2]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_3_/U21/U1/U1  ( .x(rd[59]), .a(\U1666/driveh ), .b(rd
        [59]), .c(\U1666/driveh ), .d(cbh[3]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_4_/U21/U1/U1  ( .x(rd[60]), .a(\U1666/drivel ), .b(rd
        [60]), .c(\U1666/driveh ), .d(cbh[4]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_5_/U21/U1/U1  ( .x(rd[61]), .a(\U1666/driveh ), .b(rd
        [61]), .c(n6), .d(cbh[5]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_6_/U21/U1/U1  ( .x(rd[62]), .a(n6), .b(rd[62]), .c(
        \U1666/drivel ), .d(cbh[6]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_7_/U21/U1/U1  ( .x(rd[63]), .a(n6), .b(rd[63]), .c(n6), 
        .d(cbh[7]), .e(\U1666/latch ) );
    aoai211_1 \U1666/U4/U28/U1/U1  ( .x(\U1666/U4/U28/U1/clr ), .a(read), .b(
        \U1666/acb ), .c(\U1666/nlocalcd ), .d(net169) );
    nand3_1 \U1666/U4/U28/U1/U2  ( .x(\U1666/U4/U28/U1/set ), .a(
        \U1666/nlocalcd ), .b(read), .c(\U1666/acb ) );
    nand2_2 \U1666/U4/U28/U1/U3  ( .x(net169), .a(\U1666/U4/U28/U1/clr ), .b(
        \U1666/U4/U28/U1/set ) );
    oai21_1 \U1666/U1/U30/U1/U1  ( .x(\U1666/acb ), .a(\U1666/U1/Z ), .b(
        \U1666/ba ), .c(read) );
    inv_1 \U1666/U1/U30/U1/U2  ( .x(\U1666/U1/Z ), .a(\U1666/acb ) );
    ao222_1 \U1666/U5/U18/U1/U1  ( .x(\U1666/ba ), .a(\U1666/latch ), .b(n14), 
        .c(\U1666/latch ), .d(\U1666/ba ), .e(n14), .f(\U1666/ba ) );
    aoi222_1 \U1666/U1664/U28/U30/U1  ( .x(\U1666/U1664/x[3] ), .a(
        \U1666/ncd[7] ), .b(\U1666/ncd[6] ), .c(\U1666/ncd[7] ), .d(
        \U1666/U1664/U28/Z ), .e(\U1666/ncd[6] ), .f(\U1666/U1664/U28/Z ) );
    inv_1 \U1666/U1664/U28/U30/Uinv  ( .x(\U1666/U1664/U28/Z ), .a(
        \U1666/U1664/x[3] ) );
    aoi222_1 \U1666/U1664/U32/U30/U1  ( .x(\U1666/U1664/x[0] ), .a(
        \U1666/ncd[1] ), .b(\U1666/ncd[0] ), .c(\U1666/ncd[1] ), .d(
        \U1666/U1664/U32/Z ), .e(\U1666/ncd[0] ), .f(\U1666/U1664/U32/Z ) );
    inv_1 \U1666/U1664/U32/U30/Uinv  ( .x(\U1666/U1664/U32/Z ), .a(
        \U1666/U1664/x[0] ) );
    aoi222_1 \U1666/U1664/U29/U30/U1  ( .x(\U1666/U1664/x[2] ), .a(
        \U1666/ncd[5] ), .b(\U1666/ncd[4] ), .c(\U1666/ncd[5] ), .d(
        \U1666/U1664/U29/Z ), .e(\U1666/ncd[4] ), .f(\U1666/U1664/U29/Z ) );
    inv_1 \U1666/U1664/U29/U30/Uinv  ( .x(\U1666/U1664/U29/Z ), .a(
        \U1666/U1664/x[2] ) );
    aoi222_1 \U1666/U1664/U33/U30/U1  ( .x(\U1666/U1664/y[0] ), .a(
        \U1666/U1664/x[1] ), .b(\U1666/U1664/x[0] ), .c(\U1666/U1664/x[1] ), 
        .d(\U1666/U1664/U33/Z ), .e(\U1666/U1664/x[0] ), .f(
        \U1666/U1664/U33/Z ) );
    inv_1 \U1666/U1664/U33/U30/Uinv  ( .x(\U1666/U1664/U33/Z ), .a(
        \U1666/U1664/y[0] ) );
    aoi222_1 \U1666/U1664/U30/U30/U1  ( .x(\U1666/U1664/y[1] ), .a(
        \U1666/U1664/x[3] ), .b(\U1666/U1664/x[2] ), .c(\U1666/U1664/x[3] ), 
        .d(\U1666/U1664/U30/Z ), .e(\U1666/U1664/x[2] ), .f(
        \U1666/U1664/U30/Z ) );
    inv_1 \U1666/U1664/U30/U30/Uinv  ( .x(\U1666/U1664/U30/Z ), .a(
        \U1666/U1664/y[1] ) );
    aoi222_1 \U1666/U1664/U31/U30/U1  ( .x(\U1666/U1664/x[1] ), .a(
        \U1666/ncd[3] ), .b(\U1666/ncd[2] ), .c(\U1666/ncd[3] ), .d(
        \U1666/U1664/U31/Z ), .e(\U1666/ncd[2] ), .f(\U1666/U1664/U31/Z ) );
    inv_1 \U1666/U1664/U31/U30/Uinv  ( .x(\U1666/U1664/U31/Z ), .a(
        \U1666/U1664/x[1] ) );
    aoi222_1 \U1666/U1664/U37/U30/U1  ( .x(\U1666/localcd ), .a(
        \U1666/U1664/y[0] ), .b(\U1666/U1664/y[1] ), .c(\U1666/U1664/y[0] ), 
        .d(\U1666/U1664/U37/Z ), .e(\U1666/U1664/y[1] ), .f(
        \U1666/U1664/U37/Z ) );
    inv_1 \U1666/U1664/U37/U30/Uinv  ( .x(\U1666/U1664/U37/Z ), .a(
        \U1666/localcd ) );
    nor3_1 \U1666/U1669/Unr  ( .x(\U1666/U1669/nr ), .a(
        \U1666/ctrlack_internal ), .b(n6), .c(\U1666/drivel ) );
    nand3_1 \U1666/U1669/Und  ( .x(\U1666/U1669/nd ), .a(
        \U1666/ctrlack_internal ), .b(\U1666/driveh ), .c(\U1666/drivel ) );
    oa21_1 \U1666/U1669/U1  ( .x(\U1666/U1669/n2 ), .a(\U1666/U1669/n2 ), .b(
        \U1666/U1669/nr ), .c(\U1666/U1669/nd ) );
    inv_2 \U1666/U1669/U3  ( .x(net94), .a(\U1666/U1669/n2 ) );
    buf_2 \I1/U1653  ( .x(\I1/latch ), .a(net166) );
    nor2_1 \I1/U264/U5  ( .x(\I1/nlocalcd ), .a(reset), .b(\I1/localcd ) );
    nor2_1 \I1/U1659_0_/U5  ( .x(\I1/ncd[0] ), .a(rd[8]), .b(rd[40]) );
    nor2_1 \I1/U1659_1_/U5  ( .x(\I1/ncd[1] ), .a(rd[9]), .b(rd[41]) );
    nor2_1 \I1/U1659_2_/U5  ( .x(\I1/ncd[2] ), .a(rd[10]), .b(rd[42]) );
    nor2_1 \I1/U1659_3_/U5  ( .x(\I1/ncd[3] ), .a(rd[11]), .b(rd[43]) );
    nor2_1 \I1/U1659_4_/U5  ( .x(\I1/ncd[4] ), .a(rd[12]), .b(rd[44]) );
    nor2_1 \I1/U1659_5_/U5  ( .x(\I1/ncd[5] ), .a(rd[13]), .b(rd[45]) );
    nor2_1 \I1/U1659_6_/U5  ( .x(\I1/ncd[6] ), .a(rd[14]), .b(rd[46]) );
    nor2_1 \I1/U1659_7_/U5  ( .x(\I1/ncd[7] ), .a(rd[15]), .b(rd[47]) );
    nor2_1 \I1/U3/U5  ( .x(\I1/ctrlack_internal ), .a(\I1/acb ), .b(\I1/ba )
         );
    buf_2 \I1/U1665/U7  ( .x(\I1/driveh ), .a(net103) );
    buf_2 \I1/U1666/U7  ( .x(\I1/drivel ), .a(net103) );
    ao23_1 \I1/U1658_0_/U21/U1/U1  ( .x(rd[8]), .a(n4), .b(rd[8]), .c(
        \I1/drivel ), .d(cbl[0]), .e(n3) );
    ao23_1 \I1/U1658_1_/U21/U1/U1  ( .x(rd[9]), .a(n4), .b(rd[9]), .c(
        \I1/driveh ), .d(cbl[1]), .e(n3) );
    ao23_1 \I1/U1658_2_/U21/U1/U1  ( .x(rd[10]), .a(\I1/driveh ), .b(rd[10]), 
        .c(n4), .d(cbl[2]), .e(n3) );
    ao23_1 \I1/U1658_3_/U21/U1/U1  ( .x(rd[11]), .a(n4), .b(rd[11]), .c(
        \I1/driveh ), .d(cbl[3]), .e(\I1/latch ) );
    ao23_1 \I1/U1658_4_/U21/U1/U1  ( .x(rd[12]), .a(\I1/drivel ), .b(rd[12]), 
        .c(n4), .d(cbl[4]), .e(\I1/latch ) );
    ao23_1 \I1/U1658_5_/U21/U1/U1  ( .x(rd[13]), .a(\I1/drivel ), .b(rd[13]), 
        .c(n4), .d(cbl[5]), .e(\I1/latch ) );
    ao23_1 \I1/U1658_6_/U21/U1/U1  ( .x(rd[14]), .a(\I1/driveh ), .b(rd[14]), 
        .c(\I1/drivel ), .d(cbl[6]), .e(\I1/latch ) );
    ao23_1 \I1/U1658_7_/U21/U1/U1  ( .x(rd[15]), .a(\I1/driveh ), .b(rd[15]), 
        .c(\I1/driveh ), .d(cbl[7]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_0_/U21/U1/U1  ( .x(rd[40]), .a(\I1/drivel ), .b(rd[40]), 
        .c(n4), .d(cbh[0]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_1_/U21/U1/U1  ( .x(rd[41]), .a(\I1/driveh ), .b(rd[41]), 
        .c(\I1/drivel ), .d(cbh[1]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_2_/U21/U1/U1  ( .x(rd[42]), .a(\I1/drivel ), .b(rd[42]), 
        .c(\I1/drivel ), .d(cbh[2]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_3_/U21/U1/U1  ( .x(rd[43]), .a(\I1/driveh ), .b(rd[43]), 
        .c(\I1/driveh ), .d(cbh[3]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_4_/U21/U1/U1  ( .x(rd[44]), .a(\I1/drivel ), .b(rd[44]), 
        .c(\I1/driveh ), .d(cbh[4]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_5_/U21/U1/U1  ( .x(rd[45]), .a(\I1/driveh ), .b(rd[45]), 
        .c(n4), .d(cbh[5]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_6_/U21/U1/U1  ( .x(rd[46]), .a(n4), .b(rd[46]), .c(
        \I1/drivel ), .d(cbh[6]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_7_/U21/U1/U1  ( .x(rd[47]), .a(n4), .b(rd[47]), .c(n4), 
        .d(cbh[7]), .e(\I1/latch ) );
    aoai211_1 \I1/U4/U28/U1/U1  ( .x(\I1/U4/U28/U1/clr ), .a(net103), .b(
        \I1/acb ), .c(\I1/nlocalcd ), .d(net166) );
    nand3_1 \I1/U4/U28/U1/U2  ( .x(\I1/U4/U28/U1/set ), .a(\I1/nlocalcd ), .b(
        net103), .c(\I1/acb ) );
    nand2_2 \I1/U4/U28/U1/U3  ( .x(net166), .a(\I1/U4/U28/U1/clr ), .b(
        \I1/U4/U28/U1/set ) );
    oai21_1 \I1/U1/U30/U1/U1  ( .x(\I1/acb ), .a(\I1/U1/Z ), .b(\I1/ba ), .c(
        net103) );
    inv_1 \I1/U1/U30/U1/U2  ( .x(\I1/U1/Z ), .a(\I1/acb ) );
    ao222_1 \I1/U5/U18/U1/U1  ( .x(\I1/ba ), .a(\I1/latch ), .b(n14), .c(
        \I1/latch ), .d(\I1/ba ), .e(n14), .f(\I1/ba ) );
    aoi222_1 \I1/U1664/U28/U30/U1  ( .x(\I1/U1664/x[3] ), .a(\I1/ncd[7] ), .b(
        \I1/ncd[6] ), .c(\I1/ncd[7] ), .d(\I1/U1664/U28/Z ), .e(\I1/ncd[6] ), 
        .f(\I1/U1664/U28/Z ) );
    inv_1 \I1/U1664/U28/U30/Uinv  ( .x(\I1/U1664/U28/Z ), .a(\I1/U1664/x[3] )
         );
    aoi222_1 \I1/U1664/U32/U30/U1  ( .x(\I1/U1664/x[0] ), .a(\I1/ncd[1] ), .b(
        \I1/ncd[0] ), .c(\I1/ncd[1] ), .d(\I1/U1664/U32/Z ), .e(\I1/ncd[0] ), 
        .f(\I1/U1664/U32/Z ) );
    inv_1 \I1/U1664/U32/U30/Uinv  ( .x(\I1/U1664/U32/Z ), .a(\I1/U1664/x[0] )
         );
    aoi222_1 \I1/U1664/U29/U30/U1  ( .x(\I1/U1664/x[2] ), .a(\I1/ncd[5] ), .b(
        \I1/ncd[4] ), .c(\I1/ncd[5] ), .d(\I1/U1664/U29/Z ), .e(\I1/ncd[4] ), 
        .f(\I1/U1664/U29/Z ) );
    inv_1 \I1/U1664/U29/U30/Uinv  ( .x(\I1/U1664/U29/Z ), .a(\I1/U1664/x[2] )
         );
    aoi222_1 \I1/U1664/U33/U30/U1  ( .x(\I1/U1664/y[0] ), .a(\I1/U1664/x[1] ), 
        .b(\I1/U1664/x[0] ), .c(\I1/U1664/x[1] ), .d(\I1/U1664/U33/Z ), .e(
        \I1/U1664/x[0] ), .f(\I1/U1664/U33/Z ) );
    inv_1 \I1/U1664/U33/U30/Uinv  ( .x(\I1/U1664/U33/Z ), .a(\I1/U1664/y[0] )
         );
    aoi222_1 \I1/U1664/U30/U30/U1  ( .x(\I1/U1664/y[1] ), .a(\I1/U1664/x[3] ), 
        .b(\I1/U1664/x[2] ), .c(\I1/U1664/x[3] ), .d(\I1/U1664/U30/Z ), .e(
        \I1/U1664/x[2] ), .f(\I1/U1664/U30/Z ) );
    inv_1 \I1/U1664/U30/U30/Uinv  ( .x(\I1/U1664/U30/Z ), .a(\I1/U1664/y[1] )
         );
    aoi222_1 \I1/U1664/U31/U30/U1  ( .x(\I1/U1664/x[1] ), .a(\I1/ncd[3] ), .b(
        \I1/ncd[2] ), .c(\I1/ncd[3] ), .d(\I1/U1664/U31/Z ), .e(\I1/ncd[2] ), 
        .f(\I1/U1664/U31/Z ) );
    inv_1 \I1/U1664/U31/U30/Uinv  ( .x(\I1/U1664/U31/Z ), .a(\I1/U1664/x[1] )
         );
    aoi222_1 \I1/U1664/U37/U30/U1  ( .x(\I1/localcd ), .a(\I1/U1664/y[0] ), 
        .b(\I1/U1664/y[1] ), .c(\I1/U1664/y[0] ), .d(\I1/U1664/U37/Z ), .e(
        \I1/U1664/y[1] ), .f(\I1/U1664/U37/Z ) );
    inv_1 \I1/U1664/U37/U30/Uinv  ( .x(\I1/U1664/U37/Z ), .a(\I1/localcd ) );
    nor3_1 \I1/U1669/Unr  ( .x(\I1/U1669/nr ), .a(\I1/ctrlack_internal ), .b(
        n4), .c(\I1/drivel ) );
    nand3_1 \I1/U1669/Und  ( .x(\I1/U1669/nd ), .a(\I1/ctrlack_internal ), .b(
        \I1/driveh ), .c(\I1/drivel ) );
    oa21_1 \I1/U1669/U1  ( .x(\I1/U1669/n2 ), .a(\I1/U1669/n2 ), .b(
        \I1/U1669/nr ), .c(\I1/U1669/nd ) );
    inv_2 \I1/U1669/U3  ( .x(read_lhw), .a(\I1/U1669/n2 ) );
    buf_2 \I2/U1653  ( .x(\I2/latch ), .a(net170) );
    nor2_1 \I2/U264/U5  ( .x(\I2/nlocalcd ), .a(reset), .b(\I2/localcd ) );
    nor2_1 \I2/U1659_0_/U5  ( .x(\I2/ncd[0] ), .a(rd[16]), .b(rd[48]) );
    nor2_1 \I2/U1659_1_/U5  ( .x(\I2/ncd[1] ), .a(rd[17]), .b(rd[49]) );
    nor2_1 \I2/U1659_2_/U5  ( .x(\I2/ncd[2] ), .a(rd[18]), .b(rd[50]) );
    nor2_1 \I2/U1659_3_/U5  ( .x(\I2/ncd[3] ), .a(rd[19]), .b(rd[51]) );
    nor2_1 \I2/U1659_4_/U5  ( .x(\I2/ncd[4] ), .a(rd[20]), .b(rd[52]) );
    nor2_1 \I2/U1659_5_/U5  ( .x(\I2/ncd[5] ), .a(rd[21]), .b(rd[53]) );
    nor2_1 \I2/U1659_6_/U5  ( .x(\I2/ncd[6] ), .a(rd[22]), .b(rd[54]) );
    nor2_1 \I2/U1659_7_/U5  ( .x(\I2/ncd[7] ), .a(rd[23]), .b(rd[55]) );
    nor2_1 \I2/U3/U5  ( .x(\I2/ctrlack_internal ), .a(\I2/acb ), .b(\I2/ba )
         );
    buf_2 \I2/U1665/U7  ( .x(\I2/driveh ), .a(net94) );
    buf_2 \I2/U1666/U7  ( .x(\I2/drivel ), .a(net94) );
    ao23_1 \I2/U1658_0_/U21/U1/U1  ( .x(rd[16]), .a(n2), .b(rd[16]), .c(
        \I2/drivel ), .d(cbl[0]), .e(n1) );
    ao23_1 \I2/U1658_1_/U21/U1/U1  ( .x(rd[17]), .a(n2), .b(rd[17]), .c(
        \I2/driveh ), .d(cbl[1]), .e(n1) );
    ao23_1 \I2/U1658_2_/U21/U1/U1  ( .x(rd[18]), .a(\I2/driveh ), .b(rd[18]), 
        .c(n2), .d(cbl[2]), .e(n1) );
    ao23_1 \I2/U1658_3_/U21/U1/U1  ( .x(rd[19]), .a(n2), .b(rd[19]), .c(
        \I2/driveh ), .d(cbl[3]), .e(\I2/latch ) );
    ao23_1 \I2/U1658_4_/U21/U1/U1  ( .x(rd[20]), .a(\I2/drivel ), .b(rd[20]), 
        .c(n2), .d(cbl[4]), .e(\I2/latch ) );
    ao23_1 \I2/U1658_5_/U21/U1/U1  ( .x(rd[21]), .a(\I2/drivel ), .b(rd[21]), 
        .c(n2), .d(cbl[5]), .e(\I2/latch ) );
    ao23_1 \I2/U1658_6_/U21/U1/U1  ( .x(rd[22]), .a(\I2/driveh ), .b(rd[22]), 
        .c(\I2/drivel ), .d(cbl[6]), .e(\I2/latch ) );
    ao23_1 \I2/U1658_7_/U21/U1/U1  ( .x(rd[23]), .a(\I2/driveh ), .b(rd[23]), 
        .c(\I2/driveh ), .d(cbl[7]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_0_/U21/U1/U1  ( .x(rd[48]), .a(\I2/drivel ), .b(rd[48]), 
        .c(n2), .d(cbh[0]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_1_/U21/U1/U1  ( .x(rd[49]), .a(\I2/driveh ), .b(rd[49]), 
        .c(\I2/drivel ), .d(cbh[1]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_2_/U21/U1/U1  ( .x(rd[50]), .a(\I2/drivel ), .b(rd[50]), 
        .c(\I2/drivel ), .d(cbh[2]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_3_/U21/U1/U1  ( .x(rd[51]), .a(\I2/driveh ), .b(rd[51]), 
        .c(\I2/driveh ), .d(cbh[3]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_4_/U21/U1/U1  ( .x(rd[52]), .a(\I2/drivel ), .b(rd[52]), 
        .c(\I2/driveh ), .d(cbh[4]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_5_/U21/U1/U1  ( .x(rd[53]), .a(\I2/driveh ), .b(rd[53]), 
        .c(n2), .d(cbh[5]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_6_/U21/U1/U1  ( .x(rd[54]), .a(n2), .b(rd[54]), .c(
        \I2/drivel ), .d(cbh[6]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_7_/U21/U1/U1  ( .x(rd[55]), .a(n2), .b(rd[55]), .c(n2), 
        .d(cbh[7]), .e(\I2/latch ) );
    aoai211_1 \I2/U4/U28/U1/U1  ( .x(\I2/U4/U28/U1/clr ), .a(net94), .b(
        \I2/acb ), .c(\I2/nlocalcd ), .d(net170) );
    nand3_1 \I2/U4/U28/U1/U2  ( .x(\I2/U4/U28/U1/set ), .a(\I2/nlocalcd ), .b(
        net94), .c(\I2/acb ) );
    nand2_2 \I2/U4/U28/U1/U3  ( .x(net170), .a(\I2/U4/U28/U1/clr ), .b(
        \I2/U4/U28/U1/set ) );
    oai21_1 \I2/U1/U30/U1/U1  ( .x(\I2/acb ), .a(\I2/U1/Z ), .b(\I2/ba ), .c(
        net94) );
    inv_1 \I2/U1/U30/U1/U2  ( .x(\I2/U1/Z ), .a(\I2/acb ) );
    ao222_1 \I2/U5/U18/U1/U1  ( .x(\I2/ba ), .a(\I2/latch ), .b(n14), .c(
        \I2/latch ), .d(\I2/ba ), .e(n14), .f(\I2/ba ) );
    aoi222_1 \I2/U1664/U28/U30/U1  ( .x(\I2/U1664/x[3] ), .a(\I2/ncd[7] ), .b(
        \I2/ncd[6] ), .c(\I2/ncd[7] ), .d(\I2/U1664/U28/Z ), .e(\I2/ncd[6] ), 
        .f(\I2/U1664/U28/Z ) );
    inv_1 \I2/U1664/U28/U30/Uinv  ( .x(\I2/U1664/U28/Z ), .a(\I2/U1664/x[3] )
         );
    aoi222_1 \I2/U1664/U32/U30/U1  ( .x(\I2/U1664/x[0] ), .a(\I2/ncd[1] ), .b(
        \I2/ncd[0] ), .c(\I2/ncd[1] ), .d(\I2/U1664/U32/Z ), .e(\I2/ncd[0] ), 
        .f(\I2/U1664/U32/Z ) );
    inv_1 \I2/U1664/U32/U30/Uinv  ( .x(\I2/U1664/U32/Z ), .a(\I2/U1664/x[0] )
         );
    aoi222_1 \I2/U1664/U29/U30/U1  ( .x(\I2/U1664/x[2] ), .a(\I2/ncd[5] ), .b(
        \I2/ncd[4] ), .c(\I2/ncd[5] ), .d(\I2/U1664/U29/Z ), .e(\I2/ncd[4] ), 
        .f(\I2/U1664/U29/Z ) );
    inv_1 \I2/U1664/U29/U30/Uinv  ( .x(\I2/U1664/U29/Z ), .a(\I2/U1664/x[2] )
         );
    aoi222_1 \I2/U1664/U33/U30/U1  ( .x(\I2/U1664/y[0] ), .a(\I2/U1664/x[1] ), 
        .b(\I2/U1664/x[0] ), .c(\I2/U1664/x[1] ), .d(\I2/U1664/U33/Z ), .e(
        \I2/U1664/x[0] ), .f(\I2/U1664/U33/Z ) );
    inv_1 \I2/U1664/U33/U30/Uinv  ( .x(\I2/U1664/U33/Z ), .a(\I2/U1664/y[0] )
         );
    aoi222_1 \I2/U1664/U30/U30/U1  ( .x(\I2/U1664/y[1] ), .a(\I2/U1664/x[3] ), 
        .b(\I2/U1664/x[2] ), .c(\I2/U1664/x[3] ), .d(\I2/U1664/U30/Z ), .e(
        \I2/U1664/x[2] ), .f(\I2/U1664/U30/Z ) );
    inv_1 \I2/U1664/U30/U30/Uinv  ( .x(\I2/U1664/U30/Z ), .a(\I2/U1664/y[1] )
         );
    aoi222_1 \I2/U1664/U31/U30/U1  ( .x(\I2/U1664/x[1] ), .a(\I2/ncd[3] ), .b(
        \I2/ncd[2] ), .c(\I2/ncd[3] ), .d(\I2/U1664/U31/Z ), .e(\I2/ncd[2] ), 
        .f(\I2/U1664/U31/Z ) );
    inv_1 \I2/U1664/U31/U30/Uinv  ( .x(\I2/U1664/U31/Z ), .a(\I2/U1664/x[1] )
         );
    aoi222_1 \I2/U1664/U37/U30/U1  ( .x(\I2/localcd ), .a(\I2/U1664/y[0] ), 
        .b(\I2/U1664/y[1] ), .c(\I2/U1664/y[0] ), .d(\I2/U1664/U37/Z ), .e(
        \I2/U1664/y[1] ), .f(\I2/U1664/U37/Z ) );
    inv_1 \I2/U1664/U37/U30/Uinv  ( .x(\I2/U1664/U37/Z ), .a(\I2/localcd ) );
    nor3_1 \I2/U1669/Unr  ( .x(\I2/U1669/nr ), .a(\I2/ctrlack_internal ), .b(
        n2), .c(\I2/drivel ) );
    nand3_1 \I2/U1669/Und  ( .x(\I2/U1669/nd ), .a(\I2/ctrlack_internal ), .b(
        \I2/driveh ), .c(\I2/drivel ) );
    oa21_1 \I2/U1669/U1  ( .x(\I2/U1669/n2 ), .a(\I2/U1669/n2 ), .b(
        \I2/U1669/nr ), .c(\I2/U1669/nd ) );
    inv_2 \I2/U1669/U3  ( .x(net103), .a(\I2/U1669/n2 ) );
    buf_1 U1 ( .x(n1), .a(\I2/latch ) );
    buf_2 U2 ( .x(n2), .a(net94) );
    buf_1 U3 ( .x(n3), .a(\I1/latch ) );
    buf_2 U4 ( .x(n4), .a(net103) );
    buf_1 U5 ( .x(n5), .a(\U1666/latch ) );
    buf_2 U6 ( .x(n6), .a(read) );
    buf_1 U7 ( .x(n7), .a(\U1650/latch ) );
    buf_1 U8 ( .x(n8), .a(\U1650/driveh ) );
    buf_1 U9 ( .x(n9), .a(\U1650/drivel ) );
    buf_1 U10 ( .x(n10), .a(\U1667/latch ) );
    buf_2 U11 ( .x(n11), .a(read_lhw) );
    buf_1 U12 ( .x(n12), .a(\I6/latch ) );
    buf_2 U13 ( .x(n13), .a(net139) );
    buf_3 U14 ( .x(n14), .a(bpullcd) );
    buf_3 U15 ( .x(err[1]), .a(n17) );
    buf_3 U16 ( .x(err[0]), .a(n18) );
endmodule


module chain_fr2dr_byte_4 ( nia, oh, ol, i, nReset, noa );
output [7:0] oh;
output [7:0] ol;
input  [4:0] i;
input  nReset, noa;
output nia;
    wire nbReset, eop, ncla, csela, asela, \U891/reset , \U891/neopack , 
        \U891/iay , \U891/naack[0] , \U891/naack[1] , \U891/U1128/nb , \b[3] , 
        \b[2] , \U891/U1128/na , \b[1] , \b[0] , \U891/ackb , \a[3] , \a[2] , 
        \U891/nack , \U891/acka , \a[1] , \a[0] , bsela, bsel, asel, 
        \U891/U1118_0_/nr , naa, \U891/U1118_0_/nd , \U891/U1118_0_/n2 , 
        \U891/U1118_1_/nr , \U891/U1118_1_/nd , \U891/U1118_1_/n2 , 
        \U891/U1118_2_/nr , \U891/U1118_2_/nd , \U891/U1118_2_/n2 , 
        \U891/U1118_3_/nr , \U891/U1118_3_/nd , \U891/U1118_3_/n2 , 
        \U891/U1117_0_/nr , nba, \U891/U1117_0_/nd , \U891/U1117_0_/n2 , 
        \U891/U1117_1_/nr , \U891/U1117_1_/nd , \U891/U1117_1_/n2 , 
        \U891/U1117_2_/nr , \U891/U1117_2_/nd , \U891/U1117_2_/n2 , 
        \U891/U1117_3_/nr , \U891/U1117_3_/nd , \U891/U1117_3_/n2 , 
        \U886/reset , \U886/U1128/nb , \f[3] , \f[2] , \U886/U1128/na , \f[1] , 
        \f[0] , \U886/ackb , \U886/nack , \U886/acka , \U886/U1127/n5 , 
        \U886/U1127/n1 , \U886/U1127/n2 , \U886/U1127/n3 , \U886/U1127/n4 , 
        \e[3] , \e[2] , \e[1] , \e[0] , fsela, fsel, esela, esel, 
        \U886/U1118_0_/nr , nea, \U886/U1118_0_/nd , \U886/U1118_0_/n2 , 
        \U886/U1118_1_/nr , \U886/U1118_1_/nd , \U886/U1118_1_/n2 , 
        \U886/U1118_2_/nr , \U886/U1118_2_/nd , \U886/U1118_2_/n2 , 
        \U886/U1118_3_/nr , \U886/U1118_3_/nd , \U886/U1118_3_/n2 , 
        \U886/U1117_0_/nr , nfa, \U886/U1117_0_/nd , \U886/U1117_0_/n2 , 
        \U886/U1117_1_/nr , \U886/U1117_1_/nd , \U886/U1117_1_/n2 , 
        \U886/U1117_2_/nr , \U886/U1117_2_/nd , \U886/U1117_2_/n2 , 
        \U886/U1117_3_/nr , \U886/U1117_3_/nd , \U886/U1117_3_/n2 , 
        \U884/reset , \U884/U1128/nb , \d[3] , \d[2] , \U884/U1128/na , \d[1] , 
        \d[0] , \U884/ackb , \U884/nack , \U884/acka , \U884/U1127/n5 , 
        \U884/U1127/n1 , \U884/U1127/n2 , \U884/U1127/n3 , \U884/U1127/n4 , 
        \c[3] , \c[2] , \c[1] , \c[0] , dsela, dsel, csel, \U884/U1118_0_/nr , 
        nca, \U884/U1118_0_/nd , \U884/U1118_0_/n2 , \U884/U1118_1_/nr , 
        \U884/U1118_1_/nd , \U884/U1118_1_/n2 , \U884/U1118_2_/nr , 
        \U884/U1118_2_/nd , \U884/U1118_2_/n2 , \U884/U1118_3_/nr , 
        \U884/U1118_3_/nd , \U884/U1118_3_/n2 , \U884/U1117_0_/nr , nda, 
        \U884/U1117_0_/nd , \U884/U1117_0_/n2 , \U884/U1117_1_/nr , 
        \U884/U1117_1_/nd , \U884/U1117_1_/n2 , \U884/U1117_2_/nr , 
        \U884/U1117_2_/nd , \U884/U1117_2_/n2 , \U884/U1117_3_/nr , 
        \U884/U1117_3_/nd , \U884/U1117_3_/n2 , \U888/s , \U888/r , 
        \U888/nback , \U888/naack , \U888/reset , \U887/s , \U887/r , 
        \U887/nback , \U887/naack , \U887/reset , \U885/s , \U885/r , 
        \U885/nback , \U885/naack , \U885/reset , \U877/x , \U877/reset , 
        \U877/y , \U877/U590/U25/U1/clr , net135, \cl[3] , \cl[1] , 
        \U877/U590/U25/U1/ob , n1, \U877/U589/U25/U1/clr , \cl[0] , 
        \U877/U589/U25/U1/ob , \U877/U588/U25/U1/clr , \cl[2] , 
        \U877/U588/U25/U1/ob , \U877/U591/U25/U1/clr , \U877/U591/U25/U1/ob , 
        \U876/x , \U876/reset , \U876/y , \U876/U590/U25/U1/clr , 
        \U876/U590/U25/U1/ob , \U876/U589/U25/U1/clr , \U876/U589/U25/U1/ob , 
        \U876/U588/U25/U1/clr , \U876/U588/U25/U1/ob , \U876/U591/U25/U1/clr , 
        \U876/U591/U25/U1/ob , \U2/x , \U2/reset , \U2/y , 
        \U2/U590/U25/U1/clr , \U2/U590/U25/U1/ob , \U2/U589/U25/U1/clr , 
        \U2/U589/U25/U1/ob , \U2/U588/U25/U1/clr , \U2/U588/U25/U1/ob , 
        \U2/U591/U25/U1/clr , \U2/U591/U25/U1/ob , \U1/x , \U1/reset , \U1/y , 
        \U1/U590/U25/U1/clr , \U1/U590/U25/U1/ob , \U1/U589/U25/U1/clr , 
        \U1/U589/U25/U1/ob , \U1/U588/U25/U1/clr , \U1/U588/U25/U1/ob , 
        \U1/U591/U25/U1/clr , \U1/U591/U25/U1/ob , \U881/nack[1] , 
        \U881/nack[0] ;
    buf_2 U897 ( .x(nbReset), .a(nReset) );
    and4_1 \U894/U12  ( .x(eop), .a(ncla), .b(csela), .c(asela), .d(i[4]) );
    inv_1 \U891/U1126/U3  ( .x(\U891/reset ), .a(nbReset) );
    inv_1 \U891/U1139/U3  ( .x(\U891/neopack ), .a(eop) );
    nand3_1 \U891/U1131/U9  ( .x(\U891/iay ), .a(\U891/neopack ), .b(
        \U891/naack[0] ), .c(\U891/naack[1] ) );
    nor3_1 \U891/U1128/U27  ( .x(\U891/U1128/nb ), .a(\U891/reset ), .b(\b[3] 
        ), .c(\b[2] ) );
    nor2_1 \U891/U1128/U26  ( .x(\U891/U1128/na ), .a(\b[1] ), .b(\b[0] ) );
    nand2_2 \U891/U1128/U29  ( .x(\U891/ackb ), .a(\U891/U1128/nb ), .b(
        \U891/U1128/na ) );
    nor2_1 \U891/U1133/U5  ( .x(\U891/naack[0] ), .a(\a[3] ), .b(\a[2] ) );
    nor2_1 \U891/U1108/U5  ( .x(\U891/nack ), .a(\U891/acka ), .b(\U891/ackb )
         );
    nor2_1 \U891/U1134/U5  ( .x(\U891/naack[1] ), .a(\a[1] ), .b(\a[0] ) );
    nor2_2 \U891/U914/U6  ( .x(nia), .a(\U891/iay ), .b(\U891/ackb ) );
    nand2_1 \U891/U1130/U5  ( .x(\U891/acka ), .a(\U891/naack[0] ), .b(
        \U891/naack[1] ) );
    ao222_4 \U891/U1121/U1/U1  ( .x(bsela), .a(\U891/nack ), .b(bsel), .c(
        \U891/nack ), .d(bsela), .e(bsel), .f(bsela) );
    ao222_4 \U891/U1120/U1/U1  ( .x(asela), .a(asel), .b(\U891/nack ), .c(asel
        ), .d(asela), .e(\U891/nack ), .f(asela) );
    nor3_1 \U891/U1118_0_/Unr  ( .x(\U891/U1118_0_/nr ), .a(i[0]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_0_/Und  ( .x(\U891/U1118_0_/nd ), .a(i[0]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_0_/U1  ( .x(\U891/U1118_0_/n2 ), .a(\U891/U1118_0_/n2 ), 
        .b(\U891/U1118_0_/nr ), .c(\U891/U1118_0_/nd ) );
    inv_2 \U891/U1118_0_/U3  ( .x(\a[0] ), .a(\U891/U1118_0_/n2 ) );
    nor3_1 \U891/U1118_1_/Unr  ( .x(\U891/U1118_1_/nr ), .a(i[1]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_1_/Und  ( .x(\U891/U1118_1_/nd ), .a(i[1]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_1_/U1  ( .x(\U891/U1118_1_/n2 ), .a(\U891/U1118_1_/n2 ), 
        .b(\U891/U1118_1_/nr ), .c(\U891/U1118_1_/nd ) );
    inv_2 \U891/U1118_1_/U3  ( .x(\a[1] ), .a(\U891/U1118_1_/n2 ) );
    nor3_1 \U891/U1118_2_/Unr  ( .x(\U891/U1118_2_/nr ), .a(i[2]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_2_/Und  ( .x(\U891/U1118_2_/nd ), .a(i[2]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_2_/U1  ( .x(\U891/U1118_2_/n2 ), .a(\U891/U1118_2_/n2 ), 
        .b(\U891/U1118_2_/nr ), .c(\U891/U1118_2_/nd ) );
    inv_2 \U891/U1118_2_/U3  ( .x(\a[2] ), .a(\U891/U1118_2_/n2 ) );
    nor3_1 \U891/U1118_3_/Unr  ( .x(\U891/U1118_3_/nr ), .a(i[3]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_3_/Und  ( .x(\U891/U1118_3_/nd ), .a(i[3]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_3_/U1  ( .x(\U891/U1118_3_/n2 ), .a(\U891/U1118_3_/n2 ), 
        .b(\U891/U1118_3_/nr ), .c(\U891/U1118_3_/nd ) );
    inv_2 \U891/U1118_3_/U3  ( .x(\a[3] ), .a(\U891/U1118_3_/n2 ) );
    nor3_1 \U891/U1117_0_/Unr  ( .x(\U891/U1117_0_/nr ), .a(i[0]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_0_/Und  ( .x(\U891/U1117_0_/nd ), .a(i[0]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_0_/U1  ( .x(\U891/U1117_0_/n2 ), .a(\U891/U1117_0_/n2 ), 
        .b(\U891/U1117_0_/nr ), .c(\U891/U1117_0_/nd ) );
    inv_2 \U891/U1117_0_/U3  ( .x(\b[0] ), .a(\U891/U1117_0_/n2 ) );
    nor3_1 \U891/U1117_1_/Unr  ( .x(\U891/U1117_1_/nr ), .a(i[1]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_1_/Und  ( .x(\U891/U1117_1_/nd ), .a(i[1]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_1_/U1  ( .x(\U891/U1117_1_/n2 ), .a(\U891/U1117_1_/n2 ), 
        .b(\U891/U1117_1_/nr ), .c(\U891/U1117_1_/nd ) );
    inv_2 \U891/U1117_1_/U3  ( .x(\b[1] ), .a(\U891/U1117_1_/n2 ) );
    nor3_1 \U891/U1117_2_/Unr  ( .x(\U891/U1117_2_/nr ), .a(i[2]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_2_/Und  ( .x(\U891/U1117_2_/nd ), .a(i[2]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_2_/U1  ( .x(\U891/U1117_2_/n2 ), .a(\U891/U1117_2_/n2 ), 
        .b(\U891/U1117_2_/nr ), .c(\U891/U1117_2_/nd ) );
    inv_2 \U891/U1117_2_/U3  ( .x(\b[2] ), .a(\U891/U1117_2_/n2 ) );
    nor3_1 \U891/U1117_3_/Unr  ( .x(\U891/U1117_3_/nr ), .a(i[3]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_3_/Und  ( .x(\U891/U1117_3_/nd ), .a(i[3]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_3_/U1  ( .x(\U891/U1117_3_/n2 ), .a(\U891/U1117_3_/n2 ), 
        .b(\U891/U1117_3_/nr ), .c(\U891/U1117_3_/nd ) );
    inv_2 \U891/U1117_3_/U3  ( .x(\b[3] ), .a(\U891/U1117_3_/n2 ) );
    inv_1 \U886/U1126/U3  ( .x(\U886/reset ), .a(nbReset) );
    nor3_1 \U886/U1128/U27  ( .x(\U886/U1128/nb ), .a(\U886/reset ), .b(\f[3] 
        ), .c(\f[2] ) );
    nor2_1 \U886/U1128/U26  ( .x(\U886/U1128/na ), .a(\f[1] ), .b(\f[0] ) );
    nand2_2 \U886/U1128/U29  ( .x(\U886/ackb ), .a(\U886/U1128/nb ), .b(
        \U886/U1128/na ) );
    nor2_1 \U886/U1108/U5  ( .x(\U886/nack ), .a(\U886/acka ), .b(\U886/ackb )
         );
    nor2_2 \U886/U914/U6  ( .x(nba), .a(\U886/acka ), .b(\U886/ackb ) );
    and4_1 \U886/U1127/U25  ( .x(\U886/U1127/n5 ), .a(\U886/U1127/n1 ), .b(
        \U886/U1127/n2 ), .c(\U886/U1127/n3 ), .d(\U886/U1127/n4 ) );
    inv_1 \U886/U1127/U1  ( .x(\U886/U1127/n1 ), .a(\e[3] ) );
    inv_1 \U886/U1127/U2  ( .x(\U886/U1127/n2 ), .a(\e[2] ) );
    inv_1 \U886/U1127/U3  ( .x(\U886/U1127/n3 ), .a(\e[1] ) );
    inv_1 \U886/U1127/U4  ( .x(\U886/U1127/n4 ), .a(\e[0] ) );
    inv_2 \U886/U1127/U5  ( .x(\U886/acka ), .a(\U886/U1127/n5 ) );
    ao222_2 \U886/U1121/U19/U1/U1  ( .x(fsela), .a(\U886/nack ), .b(fsel), .c(
        \U886/nack ), .d(fsela), .e(fsel), .f(fsela) );
    ao222_2 \U886/U1120/U19/U1/U1  ( .x(esela), .a(esel), .b(\U886/nack ), .c(
        esel), .d(esela), .e(\U886/nack ), .f(esela) );
    nor3_1 \U886/U1118_0_/Unr  ( .x(\U886/U1118_0_/nr ), .a(\b[0] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_0_/Und  ( .x(\U886/U1118_0_/nd ), .a(\b[0] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_0_/U1  ( .x(\U886/U1118_0_/n2 ), .a(\U886/U1118_0_/n2 ), 
        .b(\U886/U1118_0_/nr ), .c(\U886/U1118_0_/nd ) );
    inv_2 \U886/U1118_0_/U3  ( .x(\e[0] ), .a(\U886/U1118_0_/n2 ) );
    nor3_1 \U886/U1118_1_/Unr  ( .x(\U886/U1118_1_/nr ), .a(\b[1] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_1_/Und  ( .x(\U886/U1118_1_/nd ), .a(\b[1] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_1_/U1  ( .x(\U886/U1118_1_/n2 ), .a(\U886/U1118_1_/n2 ), 
        .b(\U886/U1118_1_/nr ), .c(\U886/U1118_1_/nd ) );
    inv_2 \U886/U1118_1_/U3  ( .x(\e[1] ), .a(\U886/U1118_1_/n2 ) );
    nor3_1 \U886/U1118_2_/Unr  ( .x(\U886/U1118_2_/nr ), .a(\b[2] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_2_/Und  ( .x(\U886/U1118_2_/nd ), .a(\b[2] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_2_/U1  ( .x(\U886/U1118_2_/n2 ), .a(\U886/U1118_2_/n2 ), 
        .b(\U886/U1118_2_/nr ), .c(\U886/U1118_2_/nd ) );
    inv_2 \U886/U1118_2_/U3  ( .x(\e[2] ), .a(\U886/U1118_2_/n2 ) );
    nor3_1 \U886/U1118_3_/Unr  ( .x(\U886/U1118_3_/nr ), .a(\b[3] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_3_/Und  ( .x(\U886/U1118_3_/nd ), .a(\b[3] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_3_/U1  ( .x(\U886/U1118_3_/n2 ), .a(\U886/U1118_3_/n2 ), 
        .b(\U886/U1118_3_/nr ), .c(\U886/U1118_3_/nd ) );
    inv_2 \U886/U1118_3_/U3  ( .x(\e[3] ), .a(\U886/U1118_3_/n2 ) );
    nor3_1 \U886/U1117_0_/Unr  ( .x(\U886/U1117_0_/nr ), .a(\b[0] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_0_/Und  ( .x(\U886/U1117_0_/nd ), .a(\b[0] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_0_/U1  ( .x(\U886/U1117_0_/n2 ), .a(\U886/U1117_0_/n2 ), 
        .b(\U886/U1117_0_/nr ), .c(\U886/U1117_0_/nd ) );
    inv_2 \U886/U1117_0_/U3  ( .x(\f[0] ), .a(\U886/U1117_0_/n2 ) );
    nor3_1 \U886/U1117_1_/Unr  ( .x(\U886/U1117_1_/nr ), .a(\b[1] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_1_/Und  ( .x(\U886/U1117_1_/nd ), .a(\b[1] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_1_/U1  ( .x(\U886/U1117_1_/n2 ), .a(\U886/U1117_1_/n2 ), 
        .b(\U886/U1117_1_/nr ), .c(\U886/U1117_1_/nd ) );
    inv_2 \U886/U1117_1_/U3  ( .x(\f[1] ), .a(\U886/U1117_1_/n2 ) );
    nor3_1 \U886/U1117_2_/Unr  ( .x(\U886/U1117_2_/nr ), .a(\b[2] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_2_/Und  ( .x(\U886/U1117_2_/nd ), .a(\b[2] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_2_/U1  ( .x(\U886/U1117_2_/n2 ), .a(\U886/U1117_2_/n2 ), 
        .b(\U886/U1117_2_/nr ), .c(\U886/U1117_2_/nd ) );
    inv_2 \U886/U1117_2_/U3  ( .x(\f[2] ), .a(\U886/U1117_2_/n2 ) );
    nor3_1 \U886/U1117_3_/Unr  ( .x(\U886/U1117_3_/nr ), .a(\b[3] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_3_/Und  ( .x(\U886/U1117_3_/nd ), .a(\b[3] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_3_/U1  ( .x(\U886/U1117_3_/n2 ), .a(\U886/U1117_3_/n2 ), 
        .b(\U886/U1117_3_/nr ), .c(\U886/U1117_3_/nd ) );
    inv_2 \U886/U1117_3_/U3  ( .x(\f[3] ), .a(\U886/U1117_3_/n2 ) );
    inv_1 \U884/U1126/U3  ( .x(\U884/reset ), .a(nbReset) );
    nor3_1 \U884/U1128/U27  ( .x(\U884/U1128/nb ), .a(\U884/reset ), .b(\d[3] 
        ), .c(\d[2] ) );
    nor2_1 \U884/U1128/U26  ( .x(\U884/U1128/na ), .a(\d[1] ), .b(\d[0] ) );
    nand2_2 \U884/U1128/U29  ( .x(\U884/ackb ), .a(\U884/U1128/nb ), .b(
        \U884/U1128/na ) );
    nor2_1 \U884/U1108/U5  ( .x(\U884/nack ), .a(\U884/acka ), .b(\U884/ackb )
         );
    nor2_2 \U884/U914/U6  ( .x(naa), .a(\U884/acka ), .b(\U884/ackb ) );
    and4_1 \U884/U1127/U25  ( .x(\U884/U1127/n5 ), .a(\U884/U1127/n1 ), .b(
        \U884/U1127/n2 ), .c(\U884/U1127/n3 ), .d(\U884/U1127/n4 ) );
    inv_1 \U884/U1127/U1  ( .x(\U884/U1127/n1 ), .a(\c[3] ) );
    inv_1 \U884/U1127/U2  ( .x(\U884/U1127/n2 ), .a(\c[2] ) );
    inv_1 \U884/U1127/U3  ( .x(\U884/U1127/n3 ), .a(\c[1] ) );
    inv_1 \U884/U1127/U4  ( .x(\U884/U1127/n4 ), .a(\c[0] ) );
    inv_2 \U884/U1127/U5  ( .x(\U884/acka ), .a(\U884/U1127/n5 ) );
    ao222_2 \U884/U1121/U19/U1/U1  ( .x(dsela), .a(\U884/nack ), .b(dsel), .c(
        \U884/nack ), .d(dsela), .e(dsel), .f(dsela) );
    ao222_2 \U884/U1120/U19/U1/U1  ( .x(csela), .a(csel), .b(\U884/nack ), .c(
        csel), .d(csela), .e(\U884/nack ), .f(csela) );
    nor3_1 \U884/U1118_0_/Unr  ( .x(\U884/U1118_0_/nr ), .a(\a[0] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_0_/Und  ( .x(\U884/U1118_0_/nd ), .a(\a[0] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_0_/U1  ( .x(\U884/U1118_0_/n2 ), .a(\U884/U1118_0_/n2 ), 
        .b(\U884/U1118_0_/nr ), .c(\U884/U1118_0_/nd ) );
    inv_2 \U884/U1118_0_/U3  ( .x(\c[0] ), .a(\U884/U1118_0_/n2 ) );
    nor3_1 \U884/U1118_1_/Unr  ( .x(\U884/U1118_1_/nr ), .a(\a[1] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_1_/Und  ( .x(\U884/U1118_1_/nd ), .a(\a[1] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_1_/U1  ( .x(\U884/U1118_1_/n2 ), .a(\U884/U1118_1_/n2 ), 
        .b(\U884/U1118_1_/nr ), .c(\U884/U1118_1_/nd ) );
    inv_2 \U884/U1118_1_/U3  ( .x(\c[1] ), .a(\U884/U1118_1_/n2 ) );
    nor3_1 \U884/U1118_2_/Unr  ( .x(\U884/U1118_2_/nr ), .a(\a[2] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_2_/Und  ( .x(\U884/U1118_2_/nd ), .a(\a[2] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_2_/U1  ( .x(\U884/U1118_2_/n2 ), .a(\U884/U1118_2_/n2 ), 
        .b(\U884/U1118_2_/nr ), .c(\U884/U1118_2_/nd ) );
    inv_2 \U884/U1118_2_/U3  ( .x(\c[2] ), .a(\U884/U1118_2_/n2 ) );
    nor3_1 \U884/U1118_3_/Unr  ( .x(\U884/U1118_3_/nr ), .a(\a[3] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_3_/Und  ( .x(\U884/U1118_3_/nd ), .a(\a[3] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_3_/U1  ( .x(\U884/U1118_3_/n2 ), .a(\U884/U1118_3_/n2 ), 
        .b(\U884/U1118_3_/nr ), .c(\U884/U1118_3_/nd ) );
    inv_2 \U884/U1118_3_/U3  ( .x(\c[3] ), .a(\U884/U1118_3_/n2 ) );
    nor3_1 \U884/U1117_0_/Unr  ( .x(\U884/U1117_0_/nr ), .a(\a[0] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_0_/Und  ( .x(\U884/U1117_0_/nd ), .a(\a[0] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_0_/U1  ( .x(\U884/U1117_0_/n2 ), .a(\U884/U1117_0_/n2 ), 
        .b(\U884/U1117_0_/nr ), .c(\U884/U1117_0_/nd ) );
    inv_2 \U884/U1117_0_/U3  ( .x(\d[0] ), .a(\U884/U1117_0_/n2 ) );
    nor3_1 \U884/U1117_1_/Unr  ( .x(\U884/U1117_1_/nr ), .a(\a[1] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_1_/Und  ( .x(\U884/U1117_1_/nd ), .a(\a[1] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_1_/U1  ( .x(\U884/U1117_1_/n2 ), .a(\U884/U1117_1_/n2 ), 
        .b(\U884/U1117_1_/nr ), .c(\U884/U1117_1_/nd ) );
    inv_2 \U884/U1117_1_/U3  ( .x(\d[1] ), .a(\U884/U1117_1_/n2 ) );
    nor3_1 \U884/U1117_2_/Unr  ( .x(\U884/U1117_2_/nr ), .a(\a[2] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_2_/Und  ( .x(\U884/U1117_2_/nd ), .a(\a[2] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_2_/U1  ( .x(\U884/U1117_2_/n2 ), .a(\U884/U1117_2_/n2 ), 
        .b(\U884/U1117_2_/nr ), .c(\U884/U1117_2_/nd ) );
    inv_2 \U884/U1117_2_/U3  ( .x(\d[2] ), .a(\U884/U1117_2_/n2 ) );
    nor3_1 \U884/U1117_3_/Unr  ( .x(\U884/U1117_3_/nr ), .a(\a[3] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_3_/Und  ( .x(\U884/U1117_3_/nd ), .a(\a[3] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_3_/U1  ( .x(\U884/U1117_3_/n2 ), .a(\U884/U1117_3_/n2 ), 
        .b(\U884/U1117_3_/nr ), .c(\U884/U1117_3_/nd ) );
    inv_2 \U884/U1117_3_/U3  ( .x(\d[3] ), .a(\U884/U1117_3_/n2 ) );
    nand2_1 \U888/U1128/U5  ( .x(\U888/s ), .a(\U888/r ), .b(\U888/nback ) );
    nand2_1 \U888/U1103/U5  ( .x(\U888/r ), .a(\U888/naack ), .b(\U888/s ) );
    inv_1 \U888/U1111/U3  ( .x(\U888/reset ), .a(nbReset) );
    inv_1 \U888/U1112/U3  ( .x(\U888/naack ), .a(esela) );
    nor2_1 \U888/U1127/U5  ( .x(\U888/nback ), .a(fsela), .b(\U888/reset ) );
    and2_2 \U888/U1129/U8  ( .x(esel), .a(\U888/nback ), .b(\U888/s ) );
    and2_2 \U888/U1124/U8  ( .x(fsel), .a(\U888/r ), .b(\U888/naack ) );
    nand2_1 \U887/U1128/U5  ( .x(\U887/s ), .a(\U887/r ), .b(\U887/nback ) );
    nand2_1 \U887/U1103/U5  ( .x(\U887/r ), .a(\U887/naack ), .b(\U887/s ) );
    inv_1 \U887/U1111/U3  ( .x(\U887/reset ), .a(nbReset) );
    inv_1 \U887/U1112/U3  ( .x(\U887/naack ), .a(csela) );
    nor2_1 \U887/U1127/U5  ( .x(\U887/nback ), .a(dsela), .b(\U887/reset ) );
    and2_2 \U887/U1129/U8  ( .x(csel), .a(\U887/nback ), .b(\U887/s ) );
    and2_2 \U887/U1124/U8  ( .x(dsel), .a(\U887/r ), .b(\U887/naack ) );
    nand2_1 \U885/U1128/U5  ( .x(\U885/s ), .a(\U885/r ), .b(\U885/nback ) );
    nand2_1 \U885/U1103/U5  ( .x(\U885/r ), .a(\U885/naack ), .b(\U885/s ) );
    inv_1 \U885/U1111/U3  ( .x(\U885/reset ), .a(nbReset) );
    inv_1 \U885/U1112/U3  ( .x(\U885/naack ), .a(asela) );
    nor2_1 \U885/U1127/U5  ( .x(\U885/nback ), .a(bsela), .b(\U885/reset ) );
    and2_2 \U885/U1129/U8  ( .x(asel), .a(\U885/nback ), .b(\U885/s ) );
    and2_2 \U885/U1124/U8  ( .x(bsel), .a(\U885/r ), .b(\U885/naack ) );
    nor3_1 \U877/U594/U7  ( .x(\U877/x ), .a(ol[7]), .b(\U877/reset ), .c(oh
        [7]) );
    nor3_1 \U877/U593/U7  ( .x(\U877/y ), .a(ol[6]), .b(\U877/reset ), .c(oh
        [6]) );
    inv_1 \U877/U604/U3  ( .x(\U877/reset ), .a(nbReset) );
    oa31_1 \U877/U590/U25/U1/Uclr  ( .x(\U877/U590/U25/U1/clr ), .a(net135), 
        .b(\cl[3] ), .c(\cl[1] ), .d(oh[6]) );
    oaoi211_1 \U877/U590/U25/U1/Uaoi  ( .x(\U877/U590/U25/U1/ob ), .a(\cl[3] ), 
        .b(\cl[1] ), .c(n1), .d(\U877/U590/U25/U1/clr ) );
    inv_2 \U877/U590/U25/U1/Ui  ( .x(oh[6]), .a(\U877/U590/U25/U1/ob ) );
    oa31_1 \U877/U589/U25/U1/Uclr  ( .x(\U877/U589/U25/U1/clr ), .a(net135), 
        .b(\cl[1] ), .c(\cl[0] ), .d(ol[7]) );
    oaoi211_1 \U877/U589/U25/U1/Uaoi  ( .x(\U877/U589/U25/U1/ob ), .a(\cl[1] ), 
        .b(\cl[0] ), .c(n1), .d(\U877/U589/U25/U1/clr ) );
    inv_2 \U877/U589/U25/U1/Ui  ( .x(ol[7]), .a(\U877/U589/U25/U1/ob ) );
    oa31_1 \U877/U588/U25/U1/Uclr  ( .x(\U877/U588/U25/U1/clr ), .a(net135), 
        .b(\cl[3] ), .c(\cl[2] ), .d(oh[7]) );
    oaoi211_1 \U877/U588/U25/U1/Uaoi  ( .x(\U877/U588/U25/U1/ob ), .a(\cl[3] ), 
        .b(\cl[2] ), .c(n1), .d(\U877/U588/U25/U1/clr ) );
    inv_2 \U877/U588/U25/U1/Ui  ( .x(oh[7]), .a(\U877/U588/U25/U1/ob ) );
    oa31_1 \U877/U591/U25/U1/Uclr  ( .x(\U877/U591/U25/U1/clr ), .a(net135), 
        .b(\cl[2] ), .c(\cl[0] ), .d(ol[6]) );
    oaoi211_1 \U877/U591/U25/U1/Uaoi  ( .x(\U877/U591/U25/U1/ob ), .a(\cl[2] ), 
        .b(\cl[0] ), .c(n1), .d(\U877/U591/U25/U1/clr ) );
    inv_2 \U877/U591/U25/U1/Ui  ( .x(ol[6]), .a(\U877/U591/U25/U1/ob ) );
    ao222_2 \U877/U592/U19/U1/U1  ( .x(ncla), .a(\U877/x ), .b(\U877/y ), .c(
        \U877/x ), .d(ncla), .e(\U877/y ), .f(ncla) );
    nor3_1 \U876/U594/U7  ( .x(\U876/x ), .a(ol[3]), .b(\U876/reset ), .c(oh
        [3]) );
    nor3_1 \U876/U593/U7  ( .x(\U876/y ), .a(ol[2]), .b(\U876/reset ), .c(oh
        [2]) );
    inv_1 \U876/U604/U3  ( .x(\U876/reset ), .a(nbReset) );
    oa31_1 \U876/U590/U25/U1/Uclr  ( .x(\U876/U590/U25/U1/clr ), .a(net135), 
        .b(\d[3] ), .c(\d[1] ), .d(oh[2]) );
    oaoi211_1 \U876/U590/U25/U1/Uaoi  ( .x(\U876/U590/U25/U1/ob ), .a(\d[3] ), 
        .b(\d[1] ), .c(n1), .d(\U876/U590/U25/U1/clr ) );
    inv_2 \U876/U590/U25/U1/Ui  ( .x(oh[2]), .a(\U876/U590/U25/U1/ob ) );
    oa31_1 \U876/U589/U25/U1/Uclr  ( .x(\U876/U589/U25/U1/clr ), .a(net135), 
        .b(\d[1] ), .c(\d[0] ), .d(ol[3]) );
    oaoi211_1 \U876/U589/U25/U1/Uaoi  ( .x(\U876/U589/U25/U1/ob ), .a(\d[1] ), 
        .b(\d[0] ), .c(n1), .d(\U876/U589/U25/U1/clr ) );
    inv_2 \U876/U589/U25/U1/Ui  ( .x(ol[3]), .a(\U876/U589/U25/U1/ob ) );
    oa31_1 \U876/U588/U25/U1/Uclr  ( .x(\U876/U588/U25/U1/clr ), .a(net135), 
        .b(\d[3] ), .c(\d[2] ), .d(oh[3]) );
    oaoi211_1 \U876/U588/U25/U1/Uaoi  ( .x(\U876/U588/U25/U1/ob ), .a(\d[3] ), 
        .b(\d[2] ), .c(n1), .d(\U876/U588/U25/U1/clr ) );
    inv_2 \U876/U588/U25/U1/Ui  ( .x(oh[3]), .a(\U876/U588/U25/U1/ob ) );
    oa31_1 \U876/U591/U25/U1/Uclr  ( .x(\U876/U591/U25/U1/clr ), .a(net135), 
        .b(\d[2] ), .c(\d[0] ), .d(ol[2]) );
    oaoi211_1 \U876/U591/U25/U1/Uaoi  ( .x(\U876/U591/U25/U1/ob ), .a(\d[2] ), 
        .b(\d[0] ), .c(n1), .d(\U876/U591/U25/U1/clr ) );
    inv_2 \U876/U591/U25/U1/Ui  ( .x(ol[2]), .a(\U876/U591/U25/U1/ob ) );
    ao222_2 \U876/U592/U19/U1/U1  ( .x(nda), .a(\U876/x ), .b(\U876/y ), .c(
        \U876/x ), .d(nda), .e(\U876/y ), .f(nda) );
    nor3_1 \U2/U594/U7  ( .x(\U2/x ), .a(ol[1]), .b(\U2/reset ), .c(oh[1]) );
    nor3_1 \U2/U593/U7  ( .x(\U2/y ), .a(ol[0]), .b(\U2/reset ), .c(oh[0]) );
    inv_1 \U2/U604/U3  ( .x(\U2/reset ), .a(nbReset) );
    oa31_1 \U2/U590/U25/U1/Uclr  ( .x(\U2/U590/U25/U1/clr ), .a(net135), .b(
        \f[3] ), .c(\f[1] ), .d(oh[0]) );
    oaoi211_1 \U2/U590/U25/U1/Uaoi  ( .x(\U2/U590/U25/U1/ob ), .a(\f[3] ), .b(
        \f[1] ), .c(n1), .d(\U2/U590/U25/U1/clr ) );
    inv_2 \U2/U590/U25/U1/Ui  ( .x(oh[0]), .a(\U2/U590/U25/U1/ob ) );
    oa31_1 \U2/U589/U25/U1/Uclr  ( .x(\U2/U589/U25/U1/clr ), .a(net135), .b(
        \f[1] ), .c(\f[0] ), .d(ol[1]) );
    oaoi211_1 \U2/U589/U25/U1/Uaoi  ( .x(\U2/U589/U25/U1/ob ), .a(\f[1] ), .b(
        \f[0] ), .c(n1), .d(\U2/U589/U25/U1/clr ) );
    inv_2 \U2/U589/U25/U1/Ui  ( .x(ol[1]), .a(\U2/U589/U25/U1/ob ) );
    oa31_1 \U2/U588/U25/U1/Uclr  ( .x(\U2/U588/U25/U1/clr ), .a(net135), .b(
        \f[3] ), .c(\f[2] ), .d(oh[1]) );
    oaoi211_1 \U2/U588/U25/U1/Uaoi  ( .x(\U2/U588/U25/U1/ob ), .a(\f[3] ), .b(
        \f[2] ), .c(n1), .d(\U2/U588/U25/U1/clr ) );
    inv_2 \U2/U588/U25/U1/Ui  ( .x(oh[1]), .a(\U2/U588/U25/U1/ob ) );
    oa31_1 \U2/U591/U25/U1/Uclr  ( .x(\U2/U591/U25/U1/clr ), .a(net135), .b(
        \f[2] ), .c(\f[0] ), .d(ol[0]) );
    oaoi211_1 \U2/U591/U25/U1/Uaoi  ( .x(\U2/U591/U25/U1/ob ), .a(\f[2] ), .b(
        \f[0] ), .c(n1), .d(\U2/U591/U25/U1/clr ) );
    inv_2 \U2/U591/U25/U1/Ui  ( .x(ol[0]), .a(\U2/U591/U25/U1/ob ) );
    ao222_2 \U2/U592/U19/U1/U1  ( .x(nfa), .a(\U2/x ), .b(\U2/y ), .c(\U2/x ), 
        .d(nfa), .e(\U2/y ), .f(nfa) );
    nor3_1 \U1/U594/U7  ( .x(\U1/x ), .a(ol[5]), .b(\U1/reset ), .c(oh[5]) );
    nor3_1 \U1/U593/U7  ( .x(\U1/y ), .a(ol[4]), .b(\U1/reset ), .c(oh[4]) );
    inv_1 \U1/U604/U3  ( .x(\U1/reset ), .a(nbReset) );
    oa31_1 \U1/U590/U25/U1/Uclr  ( .x(\U1/U590/U25/U1/clr ), .a(net135), .b(
        \e[3] ), .c(\e[1] ), .d(oh[4]) );
    oaoi211_1 \U1/U590/U25/U1/Uaoi  ( .x(\U1/U590/U25/U1/ob ), .a(\e[3] ), .b(
        \e[1] ), .c(n1), .d(\U1/U590/U25/U1/clr ) );
    inv_2 \U1/U590/U25/U1/Ui  ( .x(oh[4]), .a(\U1/U590/U25/U1/ob ) );
    oa31_1 \U1/U589/U25/U1/Uclr  ( .x(\U1/U589/U25/U1/clr ), .a(net135), .b(
        \e[1] ), .c(\e[0] ), .d(ol[5]) );
    oaoi211_1 \U1/U589/U25/U1/Uaoi  ( .x(\U1/U589/U25/U1/ob ), .a(\e[1] ), .b(
        \e[0] ), .c(n1), .d(\U1/U589/U25/U1/clr ) );
    inv_2 \U1/U589/U25/U1/Ui  ( .x(ol[5]), .a(\U1/U589/U25/U1/ob ) );
    oa31_1 \U1/U588/U25/U1/Uclr  ( .x(\U1/U588/U25/U1/clr ), .a(net135), .b(
        \e[3] ), .c(\e[2] ), .d(oh[5]) );
    oaoi211_1 \U1/U588/U25/U1/Uaoi  ( .x(\U1/U588/U25/U1/ob ), .a(\e[3] ), .b(
        \e[2] ), .c(n1), .d(\U1/U588/U25/U1/clr ) );
    inv_2 \U1/U588/U25/U1/Ui  ( .x(oh[5]), .a(\U1/U588/U25/U1/ob ) );
    oa31_1 \U1/U591/U25/U1/Uclr  ( .x(\U1/U591/U25/U1/clr ), .a(net135), .b(
        \e[2] ), .c(\e[0] ), .d(ol[4]) );
    oaoi211_1 \U1/U591/U25/U1/Uaoi  ( .x(\U1/U591/U25/U1/ob ), .a(\e[2] ), .b(
        \e[0] ), .c(n1), .d(\U1/U591/U25/U1/clr ) );
    inv_2 \U1/U591/U25/U1/Ui  ( .x(ol[4]), .a(\U1/U591/U25/U1/ob ) );
    ao222_2 \U1/U592/U19/U1/U1  ( .x(nea), .a(\U1/x ), .b(\U1/y ), .c(\U1/x ), 
        .d(nea), .e(\U1/y ), .f(nea) );
    and3_4 \U881/U20/U9  ( .x(nca), .a(\U881/nack[1] ), .b(\U881/nack[0] ), 
        .c(nbReset) );
    nor2_1 \U881/U18/U5  ( .x(\U881/nack[0] ), .a(\cl[3] ), .b(\cl[0] ) );
    nor2_1 \U881/U19/U5  ( .x(\U881/nack[1] ), .a(\cl[1] ), .b(\cl[2] ) );
    ao222_2 \U881/U15_0_/U19/U1/U1  ( .x(\cl[0] ), .a(\c[0] ), .b(ncla), .c(
        \c[0] ), .d(\cl[0] ), .e(ncla), .f(\cl[0] ) );
    ao222_2 \U881/U15_1_/U19/U1/U1  ( .x(\cl[1] ), .a(\c[1] ), .b(ncla), .c(
        \c[1] ), .d(\cl[1] ), .e(ncla), .f(\cl[1] ) );
    ao222_2 \U881/U15_2_/U19/U1/U1  ( .x(\cl[2] ), .a(\c[2] ), .b(ncla), .c(
        \c[2] ), .d(\cl[2] ), .e(ncla), .f(\cl[2] ) );
    ao222_2 \U881/U15_3_/U19/U1/U1  ( .x(\cl[3] ), .a(\c[3] ), .b(ncla), .c(
        \c[3] ), .d(\cl[3] ), .e(ncla), .f(\cl[3] ) );
    and2_5 U1 ( .x(n1), .a(nbReset), .b(noa) );
    and2_3 U2 ( .x(net135), .a(nbReset), .b(noa) );
endmodule


module chain_ic_ctrl_1 ( ack, candefer, eop, nstatack, pltxreq, routetxreq, 
    tok_ack, accept, candefer_ack, defer, eopack, lock, nReset, pltxack, 
    routetxack, tok_err, tok_ok );
input  [1:0] candefer_ack;
input  [1:0] lock;
input  accept, defer, eopack, nReset, pltxack, routetxack, tok_err, tok_ok;
output ack, candefer, eop, nstatack, pltxreq, routetxreq, tok_ack;
    wire net23, net25, net6, net19, net9, retry, net31, net24, net28, net27, 
        net7, net18, net13, net8, net11, net15, \U249/n5 , \U249/n1 , 
        \U249/n2 , \U249/n3 , \U249/n4 , txnodefer, net16, reset, net17, net29, 
        net12, txmaydefer, nlclear, net4, net22, net14, txlocked, net3, 
        \U286/U28/U1/clr , n1, \U286/U28/U1/set , \U285/U28/U1/clr , n2, 
        \U285/U28/U1/set , txunlocked, net2, txdone, net5, lockcleared, 
        \U262/U25/U1/clr , \U262/U25/U1/ob , \U284/U25/U1/clr , 
        \U284/U25/U1/ob , \U283/U25/U1/clr , net10, \U283/U25/U1/ob , net20, 
        \U289/Z , net21, \U287/Z , \U288/Z , \U149/nr , net30, \U149/nd , 
        \U149/n2 , \locked[0] , \locked[1] , lwrite, \U160/acb , net26, 
        \U160/U1/Z , \U136/nclear_latch , \U136/nwl , \U136/nulsense , 
        \U136/nlsense , \U136/nwh ;
    nand2_1 \U146/U5  ( .x(candefer), .a(net23), .b(net25) );
    or2_1 \U277/U12  ( .x(net6), .a(net19), .b(net9) );
    or2_1 \U264/U12  ( .x(retry), .a(net31), .b(net24) );
    or2_1 \U259/U12  ( .x(net28), .a(net27), .b(net7) );
    or2_1 \U140/U12  ( .x(net18), .a(net13), .b(net8) );
    or2_1 \U148/U12  ( .x(net11), .a(net15), .b(routetxack) );
    and4_1 \U249/U16  ( .x(\U249/n5 ), .a(\U249/n1 ), .b(\U249/n2 ), .c(
        \U249/n3 ), .d(\U249/n4 ) );
    inv_1 \U249/U1  ( .x(\U249/n1 ), .a(txnodefer) );
    inv_1 \U249/U2  ( .x(\U249/n2 ), .a(net16) );
    inv_1 \U249/U3  ( .x(\U249/n3 ), .a(net9) );
    inv_1 \U249/U4  ( .x(\U249/n4 ), .a(net19) );
    inv_1 \U249/U5  ( .x(ack), .a(\U249/n5 ) );
    nor3_2 \U40/U16  ( .x(nstatack), .a(net16), .b(reset), .c(retry) );
    nor3_2 \U275/U16  ( .x(net17), .a(net29), .b(reset), .c(tok_ack) );
    buf_3 \U290/U8  ( .x(net12), .a(txmaydefer) );
    nor2_1 \U154/U5  ( .x(nlclear), .a(net4), .b(net31) );
    or2_2 \U274/U12  ( .x(pltxreq), .a(net22), .b(net14) );
    or3_1 \U260/U12  ( .x(eop), .a(net31), .b(txlocked), .c(net4) );
    inv_1 \U147/U3  ( .x(net3), .a(net29) );
    inv_1 \U174/U3  ( .x(reset), .a(nReset) );
    aoai211_1 \U286/U28/U1/U1  ( .x(\U286/U28/U1/clr ), .a(net3), .b(n1), .c(
        net17), .d(net22) );
    nand3_1 \U286/U28/U1/U2  ( .x(\U286/U28/U1/set ), .a(net17), .b(net3), .c(
        n1) );
    nand2_2 \U286/U28/U1/U3  ( .x(net22), .a(\U286/U28/U1/clr ), .b(
        \U286/U28/U1/set ) );
    aoai211_1 \U285/U28/U1/U1  ( .x(\U285/U28/U1/clr ), .a(net3), .b(n2), .c(
        net17), .d(net14) );
    nand3_1 \U285/U28/U1/U2  ( .x(\U285/U28/U1/set ), .a(net17), .b(net3), .c(
        n2) );
    nand2_2 \U285/U28/U1/U3  ( .x(net14), .a(\U285/U28/U1/clr ), .b(
        \U285/U28/U1/set ) );
    ao222_1 \U254/U18/U1/U1  ( .x(net31), .a(defer), .b(txunlocked), .c(defer), 
        .d(net31), .e(txunlocked), .f(net31) );
    ao222_1 \U252/U18/U1/U1  ( .x(net19), .a(tok_err), .b(net12), .c(tok_err), 
        .d(net19), .e(net12), .f(net19) );
    ao222_1 \U276/U18/U1/U1  ( .x(net24), .a(txlocked), .b(defer), .c(txlocked
        ), .d(net24), .e(defer), .f(net24) );
    ao222_1 \U251/U18/U1/U1  ( .x(net9), .a(tok_ok), .b(net12), .c(tok_ok), 
        .d(net9), .e(net12), .f(net9) );
    ao222_1 \U235/U18/U1/U1  ( .x(tok_ack), .a(ack), .b(net2), .c(ack), .d(
        tok_ack), .e(net2), .f(tok_ack) );
    ao222_1 \U247/U18/U1/U1  ( .x(txnodefer), .a(txdone), .b(candefer_ack[0]), 
        .c(txdone), .d(txnodefer), .e(candefer_ack[0]), .f(txnodefer) );
    ao222_2 \U246/U19/U1/U1  ( .x(txlocked), .a(net14), .b(txdone), .c(net14), 
        .d(txlocked), .e(txdone), .f(txlocked) );
    ao222_2 \U245/U19/U1/U1  ( .x(txunlocked), .a(txdone), .b(net22), .c(
        txdone), .d(txunlocked), .e(net22), .f(txunlocked) );
    ao222_1 \U269/U18/U1/U1  ( .x(net2), .a(net28), .b(net18), .c(net28), .d(
        net2), .e(net18), .f(net2) );
    ao222_1 \U268/U18/U1/U1  ( .x(net5), .a(eopack), .b(lockcleared), .c(
        eopack), .d(net5), .e(lockcleared), .f(net5) );
    ao222_1 \U256/U18/U1/U1  ( .x(net4), .a(tok_err), .b(txunlocked), .c(
        tok_err), .d(net4), .e(txunlocked), .f(net4) );
    ao222_1 \U175/U18/U1/U1  ( .x(net29), .a(net2), .b(retry), .c(net2), .d(
        net29), .e(retry), .f(net29) );
    ao222_1 \U255/U18/U1/U1  ( .x(net8), .a(txlocked), .b(eopack), .c(txlocked
        ), .d(net8), .e(eopack), .f(net8) );
    ao222_2 \U248/U19/U1/U1  ( .x(txmaydefer), .a(candefer_ack[1]), .b(txdone), 
        .c(candefer_ack[1]), .d(txmaydefer), .e(txdone), .f(txmaydefer) );
    ao222_2 \U250/U19/U1/U1  ( .x(net16), .a(accept), .b(net12), .c(accept), 
        .d(net16), .e(net12), .f(net16) );
    oa31_1 \U262/U25/U1/Uclr  ( .x(\U262/U25/U1/clr ), .a(txunlocked), .b(net5
        ), .c(tok_ok), .d(net13) );
    oaoi211_1 \U262/U25/U1/Uaoi  ( .x(\U262/U25/U1/ob ), .a(net5), .b(tok_ok), 
        .c(txunlocked), .d(\U262/U25/U1/clr ) );
    inv_2 \U262/U25/U1/Ui  ( .x(net13), .a(\U262/U25/U1/ob ) );
    oa31_1 \U284/U25/U1/Uclr  ( .x(\U284/U25/U1/clr ), .a(txnodefer), .b(
        tok_ok), .c(tok_err), .d(net27) );
    oaoi211_1 \U284/U25/U1/Uaoi  ( .x(\U284/U25/U1/ob ), .a(tok_ok), .b(
        tok_err), .c(txnodefer), .d(\U284/U25/U1/clr ) );
    inv_2 \U284/U25/U1/Ui  ( .x(net27), .a(\U284/U25/U1/ob ) );
    oa31_1 \U283/U25/U1/Uclr  ( .x(\U283/U25/U1/clr ), .a(net10), .b(net6), 
        .c(retry), .d(net7) );
    oaoi211_1 \U283/U25/U1/Uaoi  ( .x(\U283/U25/U1/ob ), .a(net6), .b(retry), 
        .c(net10), .d(\U283/U25/U1/clr ) );
    inv_2 \U283/U25/U1/Ui  ( .x(net7), .a(\U283/U25/U1/ob ) );
    aoi21_1 \U289/U30/U1/U1  ( .x(net20), .a(\U289/Z ), .b(net16), .c(net12)
         );
    inv_1 \U289/U30/U1/U2  ( .x(\U289/Z ), .a(net20) );
    aoi21_1 \U287/U30/U1/U1  ( .x(net21), .a(\U287/Z ), .b(accept), .c(net12)
         );
    inv_1 \U287/U30/U1/U2  ( .x(\U287/Z ), .a(net21) );
    aoi222_1 \U288/U30/U1  ( .x(net10), .a(net20), .b(net21), .c(net20), .d(
        \U288/Z ), .e(net21), .f(\U288/Z ) );
    inv_1 \U288/U30/Uinv  ( .x(\U288/Z ), .a(net10) );
    nor3_1 \U149/Unr  ( .x(\U149/nr ), .a(pltxack), .b(net11), .c(net30) );
    nand3_1 \U149/Und  ( .x(\U149/nd ), .a(pltxack), .b(net11), .c(net30) );
    oa21_1 \U149/U1  ( .x(\U149/n2 ), .a(\U149/n2 ), .b(\U149/nr ), .c(
        \U149/nd ) );
    inv_2 \U149/U3  ( .x(txdone), .a(\U149/n2 ) );
    inv_1 \U133/U618/U3  ( .x(net23), .a(net15) );
    inv_1 \U133/U617/U3  ( .x(net25), .a(routetxreq) );
    ao23_1 \U133/U616/U21/U1/U1  ( .x(routetxreq), .a(pltxreq), .b(routetxreq), 
        .c(pltxreq), .d(\locked[0] ), .e(net23) );
    ao23_1 \U133/U615/U21/U1/U1  ( .x(net15), .a(pltxreq), .b(net15), .c(
        pltxreq), .d(\locked[1] ), .e(net25) );
    and2_1 \U160/U2/U8  ( .x(lwrite), .a(candefer), .b(\U160/acb ) );
    nor2_1 \U160/U3/U5  ( .x(net30), .a(\U160/acb ), .b(net26) );
    oai21_1 \U160/U1/U30/U1/U1  ( .x(\U160/acb ), .a(\U160/U1/Z ), .b(net26), 
        .c(candefer) );
    inv_1 \U160/U1/U30/U1/U2  ( .x(\U160/U1/Z ), .a(\U160/acb ) );
    nand3_2 \U136/U48/U16  ( .x(\locked[0] ), .a(\locked[1] ), .b(
        \U136/nclear_latch ), .c(\U136/nwl ) );
    nor2_0 \U136/U36/U5  ( .x(\U136/nulsense ), .a(\locked[1] ), .b(\U136/nwl 
        ) );
    nor2_0 \U136/U37/U5  ( .x(\U136/nlsense ), .a(\U136/nwh ), .b(\locked[0] )
         );
    and2_1 \U136/U76/U8  ( .x(\U136/nclear_latch ), .a(nReset), .b(nlclear) );
    nor2_1 \U136/U77/U5  ( .x(lockcleared), .a(nlclear), .b(\locked[1] ) );
    nand2_1 \U136/U14/U5  ( .x(\U136/nwl ), .a(lwrite), .b(n2) );
    nand2_1 \U136/U15/U5  ( .x(\U136/nwh ), .a(n1), .b(lwrite) );
    nand2_2 \U136/U47/U5  ( .x(\locked[1] ), .a(\U136/nwh ), .b(\locked[0] )
         );
    or2_4 \U136/U35/U12  ( .x(net26), .a(\U136/nlsense ), .b(\U136/nulsense )
         );
    buf_1 U1 ( .x(n1), .a(lock[1]) );
    buf_1 U2 ( .x(n2), .a(lock[0]) );
endmodule


module chain_selement_ga_43 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_44 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_45 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_46 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_50 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_47 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_51 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_48 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_49 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_42 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_dr8bit_completion_52 ( o, i );
input  [15:0] i;
output o;
    wire \nx[0] , \nx[1] , \nx[2] , \nx[3] , \ny[0] , \ny[1] , \ny[2] , 
        \ny[3] , y, x, \U6/Z , \U3/net3 , \U3/U20/Z , \U3/net2 , \U3/U21/Z , 
        \U3/U19/Z , \U5/net3 , \U5/U20/Z , \U5/net2 , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_53 ( o, i );
input  [15:0] i;
output o;
    wire \nx[0] , \nx[1] , \nx[2] , \nx[3] , \ny[0] , \ny[1] , \ny[2] , 
        \ny[3] , y, x, \U6/Z , \U3/net3 , \U3/U20/Z , \U3/net2 , \U3/U21/Z , 
        \U3/U19/Z , \U5/net3 , \U5/U20/Z , \U5/net2 , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_24 ( o, i );
input  [15:0] i;
output o;
    wire \nx[0] , \nx[1] , \nx[2] , \nx[3] , \ny[0] , \ny[1] , \ny[2] , 
        \ny[3] , y, x, \U6/Z , \U3/net3 , \U3/U20/Z , \U3/net2 , \U3/U21/Z , 
        \U3/U19/Z , \U5/net3 , \U5/U20/Z , \U5/net2 , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_27 ( o, i );
input  [15:0] i;
output o;
    wire \nx[0] , \nx[1] , \nx[2] , \nx[3] , \ny[0] , \ny[1] , \ny[2] , 
        \ny[3] , y, x, \U6/Z , \U3/net3 , \U3/U20/Z , \U3/net2 , \U3/U21/Z , 
        \U3/U19/Z , \U5/net3 , \U5/U20/Z , \U5/net2 , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_26 ( o, i );
input  [15:0] i;
output o;
    wire \nx[0] , \nx[1] , \nx[2] , \nx[3] , \ny[0] , \ny[1] , \ny[2] , 
        \ny[3] , y, x, \U6/Z , \U3/net3 , \U3/U20/Z , \U3/net2 , \U3/U21/Z , 
        \U3/U19/Z , \U5/net3 , \U5/U20/Z , \U5/net2 , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_25 ( o, i );
input  [15:0] i;
output o;
    wire \nx[0] , \nx[1] , \nx[2] , \nx[3] , \ny[0] , \ny[1] , \ny[2] , 
        \ny[3] , y, x, \U6/Z , \U3/net3 , \U3/U20/Z , \U3/net2 , \U3/U21/Z , 
        \U3/U19/Z , \U5/net3 , \U5/U20/Z , \U5/net2 , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr32bit_completion_4 ( o, i );
input  [63:0] i;
output o;
    wire \cd[3] , \cd[2] , \cd[1] , \cd[0] , ny, \U16/Z , nx, \U6/Z , \U15/Z ;
    chain_dr8bit_completion_24 U11 ( .o(\cd[3] ), .i({i[63], i[62], i[61], 
        i[60], i[59], i[58], i[57], i[56], i[31], i[30], i[29], i[28], i[27], 
        i[26], i[25], i[24]}) );
    chain_dr8bit_completion_27 U14 ( .o(\cd[2] ), .i({i[55], i[54], i[53], 
        i[52], i[51], i[50], i[49], i[48], i[23], i[22], i[21], i[20], i[19], 
        i[18], i[17], i[16]}) );
    chain_dr8bit_completion_26 U13 ( .o(\cd[1] ), .i({i[47], i[46], i[45], 
        i[44], i[43], i[42], i[41], i[40], i[15], i[14], i[13], i[12], i[11], 
        i[10], i[9], i[8]}) );
    chain_dr8bit_completion_25 U12 ( .o(\cd[0] ), .i({i[39], i[38], i[37], 
        i[36], i[35], i[34], i[33], i[32], i[7], i[6], i[5], i[4], i[3], i[2], 
        i[1], i[0]}) );
    aoi222_1 \U16/U30/U1  ( .x(ny), .a(\cd[0] ), .b(\cd[1] ), .c(\cd[0] ), .d(
        \U16/Z ), .e(\cd[1] ), .f(\U16/Z ) );
    inv_1 \U16/U30/Uinv  ( .x(\U16/Z ), .a(ny) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(ny), .b(nx), .c(ny), .d(\U6/Z ), .e(nx), 
        .f(\U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U15/U30/U1  ( .x(nx), .a(\cd[3] ), .b(\cd[2] ), .c(\cd[3] ), .d(
        \U15/Z ), .e(\cd[2] ), .f(\U15/Z ) );
    inv_1 \U15/U30/Uinv  ( .x(\U15/Z ), .a(nx) );
endmodule


module chain_dr8bit_completion_28 ( o, i );
input  [15:0] i;
output o;
    wire \nx[0] , \nx[1] , \nx[2] , \nx[3] , \ny[0] , \ny[1] , \ny[2] , 
        \ny[3] , y, x, \U6/Z , \U3/net3 , \U3/U20/Z , \U3/net2 , \U3/U21/Z , 
        \U3/U19/Z , \U5/net3 , \U5/U20/Z , \U5/net2 , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_31 ( o, i );
input  [15:0] i;
output o;
    wire \nx[0] , \nx[1] , \nx[2] , \nx[3] , \ny[0] , \ny[1] , \ny[2] , 
        \ny[3] , y, x, \U6/Z , \U3/net3 , \U3/U20/Z , \U3/net2 , \U3/U21/Z , 
        \U3/U19/Z , \U5/net3 , \U5/U20/Z , \U5/net2 , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_30 ( o, i );
input  [15:0] i;
output o;
    wire \nx[0] , \nx[1] , \nx[2] , \nx[3] , \ny[0] , \ny[1] , \ny[2] , 
        \ny[3] , y, x, \U6/Z , \U3/net3 , \U3/U20/Z , \U3/net2 , \U3/U21/Z , 
        \U3/U19/Z , \U5/net3 , \U5/U20/Z , \U5/net2 , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_29 ( o, i );
input  [15:0] i;
output o;
    wire \nx[0] , \nx[1] , \nx[2] , \nx[3] , \ny[0] , \ny[1] , \ny[2] , 
        \ny[3] , y, x, \U6/Z , \U3/net3 , \U3/U20/Z , \U3/net2 , \U3/U21/Z , 
        \U3/U19/Z , \U5/net3 , \U5/U20/Z , \U5/net2 , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr32bit_completion_5 ( o, i );
input  [63:0] i;
output o;
    wire \cd[3] , \cd[2] , \cd[1] , \cd[0] , ny, \U16/Z , nx, \U6/Z , \U15/Z ;
    chain_dr8bit_completion_28 U11 ( .o(\cd[3] ), .i({i[63], i[62], i[61], 
        i[60], i[59], i[58], i[57], i[56], i[31], i[30], i[29], i[28], i[27], 
        i[26], i[25], i[24]}) );
    chain_dr8bit_completion_31 U14 ( .o(\cd[2] ), .i({i[55], i[54], i[53], 
        i[52], i[51], i[50], i[49], i[48], i[23], i[22], i[21], i[20], i[19], 
        i[18], i[17], i[16]}) );
    chain_dr8bit_completion_30 U13 ( .o(\cd[1] ), .i({i[47], i[46], i[45], 
        i[44], i[43], i[42], i[41], i[40], i[15], i[14], i[13], i[12], i[11], 
        i[10], i[9], i[8]}) );
    chain_dr8bit_completion_29 U12 ( .o(\cd[0] ), .i({i[39], i[38], i[37], 
        i[36], i[35], i[34], i[33], i[32], i[7], i[6], i[5], i[4], i[3], i[2], 
        i[1], i[0]}) );
    aoi222_1 \U16/U30/U1  ( .x(ny), .a(\cd[0] ), .b(\cd[1] ), .c(\cd[0] ), .d(
        \U16/Z ), .e(\cd[1] ), .f(\U16/Z ) );
    inv_1 \U16/U30/Uinv  ( .x(\U16/Z ), .a(ny) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(ny), .b(nx), .c(ny), .d(\U6/Z ), .e(nx), 
        .f(\U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U15/U30/U1  ( .x(nx), .a(\cd[3] ), .b(\cd[2] ), .c(\cd[3] ), .d(
        \U15/Z ), .e(\cd[2] ), .f(\U15/Z ) );
    inv_1 \U15/U30/Uinv  ( .x(\U15/Z ), .a(nx) );
endmodule


module chain_icmux_1 ( ack, chainh, chainl, sendack, addr, col, itag, lock, 
    nReset, nia, pred, rnw, sendreq, seq, size, wd );
output [7:0] chainh;
output [7:0] chainl;
input  [63:0] addr;
input  [5:0] col;
input  [9:0] itag;
input  [1:0] lock;
input  [1:0] pred;
input  [1:0] rnw;
input  [1:0] seq;
input  [3:0] size;
input  [63:0] wd;
input  nReset, nia, sendreq;
output ack, sendack;
    wire net152, net146, net148, n1, net156, \bs[1] , net138, net160, \bs[2] , 
        net168, \bs[3] , net172, \bs[7] , net164, net132, \bs[4] , net289, 
        \bs[8] , net180, \bs[5] , net176, \bs[6] , \bs[0] , \hdr[4] , net185, 
        net187, net189, net191, net293, net131, \net246[15] , net265, 
        \net246[14] , \net246[13] , \net246[12] , \net246[11] , \net246[10] , 
        \net246[9] , \net246[8] , \net246[7] , \net246[6] , \net246[5] , 
        \net246[4] , \net246[3] , \net246[2] , \net246[1] , \net246[0] , 
        \net243[15] , net263, \net243[14] , \net243[13] , \net243[12] , 
        \net243[11] , \net243[10] , \net243[9] , \net243[8] , \net243[7] , 
        \net243[6] , \net243[5] , \net243[4] , \net243[3] , \net243[2] , 
        \net243[1] , \net243[0] , \net240[15] , net267, \net240[14] , 
        \net240[13] , \net240[12] , \net240[11] , \net240[10] , \net240[9] , 
        \net240[8] , \net240[7] , \net240[6] , \net240[5] , \net240[4] , 
        \net240[3] , \net240[2] , \net240[1] , \net240[0] , \net237[15] , 
        net269, \net237[14] , \net237[13] , \net237[12] , \net237[11] , 
        \net237[10] , \net237[9] , \net237[8] , \net237[7] , \net237[6] , 
        \net237[5] , \net237[2] , \net237[1] , \net237[0] , \net234[15] , 
        net259, \net234[14] , \net234[13] , \net234[12] , \net234[11] , 
        \net234[10] , \net234[9] , \net234[8] , \net234[7] , \net234[6] , 
        \net234[5] , \net234[4] , \net234[3] , \net234[2] , \net234[1] , 
        \net234[0] , \net231[15] , net253, \net231[14] , \net231[13] , 
        \net231[12] , \net231[11] , \net231[10] , \net231[9] , \net231[8] , 
        \net231[7] , \net231[6] , \net231[5] , \net231[4] , \net231[3] , 
        \net231[2] , \net231[1] , \net231[0] , \net228[15] , net255, 
        \net228[14] , \net228[13] , \net228[12] , \net228[11] , \net228[10] , 
        \net228[9] , \net228[8] , \net228[7] , \net228[6] , \net228[5] , 
        \net228[4] , \net228[3] , \net228[2] , \net228[1] , \net228[0] , 
        \net225[15] , net251, \net225[14] , \net225[13] , \net225[12] , 
        \net225[11] , \net225[10] , \net225[9] , \net225[8] , \net225[7] , 
        \net225[6] , \net225[5] , \net225[4] , \net225[3] , \net225[2] , 
        \net225[1] , \net225[0] , \net222[15] , net261, \net222[14] , 
        \net222[13] , \net222[12] , \net222[11] , \net222[10] , \net222[9] , 
        \net222[8] , \net222[7] , \net222[6] , \net222[5] , \net222[4] , 
        \net222[3] , \net222[2] , \net222[1] , \net222[0] , \net219[15] , 
        net249, \net219[14] , \net219[13] , \net219[12] , \net219[11] , 
        \net219[10] , \net219[9] , \net219[8] , \net219[7] , \net219[6] , 
        \net219[5] , \net219[4] , \net219[3] , \net219[2] , \net219[1] , 
        \net219[0] , \U40_0_/n3 , \U40_0_/n4 , \net217[15] , \U40_0_/n5 , 
        \U40_1_/n3 , \U40_1_/n4 , \net217[14] , \U40_1_/n5 , \U40_2_/n3 , 
        \U40_2_/n4 , \net217[13] , \U40_2_/n5 , \U40_3_/n3 , \U40_3_/n4 , 
        \net217[12] , \U40_3_/n5 , \U40_4_/n3 , \U40_4_/n4 , \net217[11] , 
        \U40_4_/n5 , \U40_5_/n3 , \U40_5_/n4 , \net217[10] , \U40_5_/n5 , 
        \U40_6_/n3 , \U40_6_/n4 , \net217[9] , \U40_6_/n5 , \U40_7_/n3 , 
        \U40_7_/n4 , \net217[8] , \U40_7_/n5 , \U40_8_/n3 , \U40_8_/n4 , 
        \net217[7] , \U40_8_/n5 , \U40_9_/n3 , \U40_9_/n4 , \net217[6] , 
        \U40_9_/n5 , \U40_10_/n3 , \U40_10_/n4 , \net217[5] , \U40_10_/n5 , 
        \U40_11_/n3 , \U40_11_/n4 , \net217[4] , \U40_11_/n5 , \U40_12_/n3 , 
        \U40_12_/n4 , \net217[3] , \U40_12_/n5 , \U40_13_/n3 , \U40_13_/n4 , 
        \net217[2] , \U40_13_/n5 , \U40_14_/n3 , \U40_14_/n4 , \net217[1] , 
        \U40_14_/n5 , \U40_15_/n3 , \U40_15_/n4 , \net217[0] , \U40_15_/n5 , 
        \U14_0_/n5 , \U14_0_/n1 , \U14_0_/n2 , \U14_0_/n3 , \U14_0_/n4 , 
        \net212[15] , \U14_1_/n5 , \U14_1_/n1 , \U14_1_/n2 , \U14_1_/n3 , 
        \U14_1_/n4 , \net212[14] , \U14_2_/n5 , \U14_2_/n1 , \U14_2_/n2 , 
        \U14_2_/n3 , \U14_2_/n4 , \net212[13] , \U14_3_/n5 , \U14_3_/n1 , 
        \U14_3_/n2 , \U14_3_/n3 , \U14_3_/n4 , \net212[12] , \U14_4_/n5 , 
        \U14_4_/n1 , \U14_4_/n2 , \U14_4_/n3 , \U14_4_/n4 , \net212[11] , 
        \U14_5_/n5 , \U14_5_/n1 , \U14_5_/n2 , \U14_5_/n3 , \U14_5_/n4 , 
        \net212[10] , \U14_6_/n5 , \U14_6_/n1 , \U14_6_/n2 , \U14_6_/n3 , 
        \U14_6_/n4 , \net212[9] , \U14_7_/n5 , \U14_7_/n1 , \U14_7_/n2 , 
        \U14_7_/n3 , \U14_7_/n4 , \net212[8] , \U14_8_/n5 , \U14_8_/n1 , 
        \U14_8_/n2 , \U14_8_/n3 , \U14_8_/n4 , \net212[7] , \U14_9_/n5 , 
        \U14_9_/n1 , \U14_9_/n2 , \U14_9_/n3 , \U14_9_/n4 , \net212[6] , 
        \U14_10_/n5 , \U14_10_/n1 , \U14_10_/n2 , \U14_10_/n3 , \U14_10_/n4 , 
        \net212[5] , \U14_11_/n1 , \U14_11_/n2 , \U14_11_/n4 , \net212[4] , 
        \U14_11_/n5 , \U14_12_/n1 , \U14_12_/n2 , \U14_12_/n4 , \net212[3] , 
        \U14_12_/n5 , \U14_13_/n5 , \U14_13_/n1 , \U14_13_/n2 , \U14_13_/n3 , 
        \U14_13_/n4 , \net212[2] , \U14_14_/n5 , \U14_14_/n1 , \U14_14_/n2 , 
        \U14_14_/n3 , \U14_14_/n4 , \net212[1] , \U14_15_/n5 , \U14_15_/n1 , 
        \U14_15_/n2 , \U14_15_/n3 , \U14_15_/n4 , \net212[0] , \U91_0_/n5 , 
        \U91_0_/n1 , \U91_0_/n2 , \U91_0_/n3 , \U91_0_/n4 , \net207[15] , 
        \U91_1_/n5 , \U91_1_/n1 , \U91_1_/n2 , \U91_1_/n3 , \U91_1_/n4 , 
        \net207[14] , \U91_2_/n5 , \U91_2_/n1 , \U91_2_/n2 , \U91_2_/n3 , 
        \U91_2_/n4 , \net207[13] , \U91_3_/n5 , \U91_3_/n1 , \U91_3_/n2 , 
        \U91_3_/n3 , \U91_3_/n4 , \net207[12] , \U91_4_/n5 , \U91_4_/n1 , 
        \U91_4_/n2 , \U91_4_/n3 , \U91_4_/n4 , \net207[11] , \U91_5_/n5 , 
        \U91_5_/n1 , \U91_5_/n2 , \U91_5_/n3 , \U91_5_/n4 , \net207[10] , 
        \U91_6_/n5 , \U91_6_/n1 , \U91_6_/n2 , \U91_6_/n3 , \U91_6_/n4 , 
        \net207[9] , \U91_7_/n5 , \U91_7_/n1 , \U91_7_/n2 , \U91_7_/n3 , 
        \U91_7_/n4 , \net207[8] , \U91_8_/n5 , \U91_8_/n1 , \U91_8_/n2 , 
        \U91_8_/n3 , \U91_8_/n4 , \net207[7] , \U91_9_/n5 , \U91_9_/n1 , 
        \U91_9_/n2 , \U91_9_/n3 , \U91_9_/n4 , \net207[6] , \U91_10_/n5 , 
        \U91_10_/n1 , \U91_10_/n2 , \U91_10_/n3 , \U91_10_/n4 , \net207[5] , 
        \U91_11_/n5 , \U91_11_/n1 , \U91_11_/n2 , \U91_11_/n3 , \U91_11_/n4 , 
        \net207[4] , \U91_12_/n5 , \U91_12_/n1 , \U91_12_/n2 , \U91_12_/n3 , 
        \U91_12_/n4 , \net207[3] , \U91_13_/n5 , \U91_13_/n1 , \U91_13_/n2 , 
        \U91_13_/n3 , \U91_13_/n4 , \net207[2] , \U91_14_/n5 , \U91_14_/n1 , 
        \U91_14_/n2 , \U91_14_/n3 , \U91_14_/n4 , \net207[1] , \U91_15_/n5 , 
        \U91_15_/n1 , \U91_15_/n2 , \U91_15_/n3 , \U91_15_/n4 , \net207[0] , 
        net198, net136, \U151/Z , \U148/U21/nr , \U148/U21/nd , \U148/U21/n2 ;
    chain_selement_ga_43 U163 ( .Aa(net152), .Br(net146), .Ar(net148), .Ba(n1)
         );
    chain_selement_ga_44 U164 ( .Aa(net156), .Br(\bs[1] ), .Ar(net152), .Ba(
        net138) );
    chain_selement_ga_45 U165 ( .Aa(net160), .Br(\bs[2] ), .Ar(net156), .Ba(n1
        ) );
    chain_selement_ga_46 U166 ( .Aa(net168), .Br(\bs[3] ), .Ar(net160), .Ba(
        net138) );
    chain_selement_ga_50 U170 ( .Aa(net172), .Br(\bs[7] ), .Ar(net164), .Ba(
        net138) );
    chain_selement_ga_47 U167 ( .Aa(net132), .Br(\bs[4] ), .Ar(net168), .Ba(
        net138) );
    chain_selement_ga_51 U171 ( .Aa(net289), .Br(\bs[8] ), .Ar(net172), .Ba(
        net138) );
    chain_selement_ga_48 U168 ( .Aa(net180), .Br(\bs[5] ), .Ar(net176), .Ba(
        net138) );
    chain_selement_ga_49 U169 ( .Aa(net164), .Br(\bs[6] ), .Ar(net180), .Ba(n1
        ) );
    chain_selement_ga_42 U161 ( .Aa(net148), .Br(\bs[0] ), .Ar(\hdr[4] ), .Ba(
        n1) );
    chain_dr8bit_completion_52 U119 ( .o(net185), .i({col[5], col[4], col[3], 
        itag[9], itag[8], itag[7], itag[6], itag[5], col[2], col[1], col[0], 
        itag[4], itag[3], itag[2], itag[1], itag[0]}) );
    chain_dr8bit_completion_53 U147 ( .o(net187), .i({size[3], size[2], rnw[1], 
        1'b0, 1'b0, lock[1], pred[1], seq[1], size[1], size[0], rnw[0], 
        \hdr[4] , \hdr[4] , lock[0], pred[0], seq[0]}) );
    chain_dr32bit_completion_4 U117 ( .o(net189), .i(wd) );
    chain_dr32bit_completion_5 U118 ( .o(net191), .i(addr) );
    or2_4 \U122/U12  ( .x(net293), .a(net189), .b(net131) );
    or2_4 \U53/U12  ( .x(sendack), .a(net131), .b(net289) );
    and2_1 \U32_0_/U8  ( .x(\net246[15] ), .a(itag[0]), .b(net265) );
    and2_1 \U32_1_/U8  ( .x(\net246[14] ), .a(itag[1]), .b(net265) );
    and2_1 \U32_2_/U8  ( .x(\net246[13] ), .a(itag[2]), .b(net265) );
    and2_1 \U32_3_/U8  ( .x(\net246[12] ), .a(itag[3]), .b(net265) );
    and2_1 \U32_4_/U8  ( .x(\net246[11] ), .a(itag[4]), .b(net265) );
    and2_1 \U32_5_/U8  ( .x(\net246[10] ), .a(col[0]), .b(net265) );
    and2_1 \U32_6_/U8  ( .x(\net246[9] ), .a(col[1]), .b(net265) );
    and2_1 \U32_7_/U8  ( .x(\net246[8] ), .a(col[2]), .b(net265) );
    and2_1 \U32_8_/U8  ( .x(\net246[7] ), .a(itag[5]), .b(net265) );
    and2_1 \U32_9_/U8  ( .x(\net246[6] ), .a(itag[6]), .b(net265) );
    and2_1 \U32_10_/U8  ( .x(\net246[5] ), .a(itag[7]), .b(net265) );
    and2_1 \U32_11_/U8  ( .x(\net246[4] ), .a(itag[8]), .b(net265) );
    and2_1 \U32_12_/U8  ( .x(\net246[3] ), .a(itag[9]), .b(net265) );
    and2_1 \U32_13_/U8  ( .x(\net246[2] ), .a(col[3]), .b(net265) );
    and2_1 \U32_14_/U8  ( .x(\net246[1] ), .a(col[4]), .b(net265) );
    and2_1 \U32_15_/U8  ( .x(\net246[0] ), .a(col[5]), .b(net265) );
    and2_1 \U76_0_/U8  ( .x(\net243[15] ), .a(wd[8]), .b(net263) );
    and2_1 \U76_1_/U8  ( .x(\net243[14] ), .a(wd[9]), .b(net263) );
    and2_1 \U76_2_/U8  ( .x(\net243[13] ), .a(wd[10]), .b(net263) );
    and2_1 \U76_3_/U8  ( .x(\net243[12] ), .a(wd[11]), .b(net263) );
    and2_1 \U76_4_/U8  ( .x(\net243[11] ), .a(wd[12]), .b(net263) );
    and2_1 \U76_5_/U8  ( .x(\net243[10] ), .a(wd[13]), .b(net263) );
    and2_1 \U76_6_/U8  ( .x(\net243[9] ), .a(wd[14]), .b(net263) );
    and2_1 \U76_7_/U8  ( .x(\net243[8] ), .a(wd[15]), .b(net263) );
    and2_1 \U76_8_/U8  ( .x(\net243[7] ), .a(wd[40]), .b(net263) );
    and2_1 \U76_9_/U8  ( .x(\net243[6] ), .a(wd[41]), .b(net263) );
    and2_1 \U76_10_/U8  ( .x(\net243[5] ), .a(wd[42]), .b(net263) );
    and2_1 \U76_11_/U8  ( .x(\net243[4] ), .a(wd[43]), .b(net263) );
    and2_1 \U76_12_/U8  ( .x(\net243[3] ), .a(wd[44]), .b(net263) );
    and2_1 \U76_13_/U8  ( .x(\net243[2] ), .a(wd[45]), .b(net263) );
    and2_1 \U76_14_/U8  ( .x(\net243[1] ), .a(wd[46]), .b(net263) );
    and2_1 \U76_15_/U8  ( .x(\net243[0] ), .a(wd[47]), .b(net263) );
    and2_1 \U80_0_/U8  ( .x(\net240[15] ), .a(wd[16]), .b(net267) );
    and2_1 \U80_1_/U8  ( .x(\net240[14] ), .a(wd[17]), .b(net267) );
    and2_1 \U80_2_/U8  ( .x(\net240[13] ), .a(wd[18]), .b(net267) );
    and2_1 \U80_3_/U8  ( .x(\net240[12] ), .a(wd[19]), .b(net267) );
    and2_1 \U80_4_/U8  ( .x(\net240[11] ), .a(wd[20]), .b(net267) );
    and2_1 \U80_5_/U8  ( .x(\net240[10] ), .a(wd[21]), .b(net267) );
    and2_1 \U80_6_/U8  ( .x(\net240[9] ), .a(wd[22]), .b(net267) );
    and2_1 \U80_7_/U8  ( .x(\net240[8] ), .a(wd[23]), .b(net267) );
    and2_1 \U80_8_/U8  ( .x(\net240[7] ), .a(wd[48]), .b(net267) );
    and2_1 \U80_9_/U8  ( .x(\net240[6] ), .a(wd[49]), .b(net267) );
    and2_1 \U80_10_/U8  ( .x(\net240[5] ), .a(wd[50]), .b(net267) );
    and2_1 \U80_11_/U8  ( .x(\net240[4] ), .a(wd[51]), .b(net267) );
    and2_1 \U80_12_/U8  ( .x(\net240[3] ), .a(wd[52]), .b(net267) );
    and2_1 \U80_13_/U8  ( .x(\net240[2] ), .a(wd[53]), .b(net267) );
    and2_1 \U80_14_/U8  ( .x(\net240[1] ), .a(wd[54]), .b(net267) );
    and2_1 \U80_15_/U8  ( .x(\net240[0] ), .a(wd[55]), .b(net267) );
    and2_1 \U128_0_/U8  ( .x(\net237[15] ), .a(seq[0]), .b(net269) );
    and2_1 \U128_1_/U8  ( .x(\net237[14] ), .a(pred[0]), .b(net269) );
    and2_1 \U128_2_/U8  ( .x(\net237[13] ), .a(lock[0]), .b(net269) );
    and2_1 \U128_3_/U8  ( .x(\net237[12] ), .a(\hdr[4] ), .b(net269) );
    and2_1 \U128_4_/U8  ( .x(\net237[11] ), .a(\hdr[4] ), .b(net269) );
    and2_1 \U128_5_/U8  ( .x(\net237[10] ), .a(rnw[0]), .b(net269) );
    and2_1 \U128_6_/U8  ( .x(\net237[9] ), .a(size[0]), .b(net269) );
    and2_1 \U128_7_/U8  ( .x(\net237[8] ), .a(size[1]), .b(net269) );
    and2_1 \U128_8_/U8  ( .x(\net237[7] ), .a(seq[1]), .b(net269) );
    and2_1 \U128_9_/U8  ( .x(\net237[6] ), .a(pred[1]), .b(net269) );
    and2_1 \U128_10_/U8  ( .x(\net237[5] ), .a(lock[1]), .b(net269) );
    and2_1 \U128_13_/U8  ( .x(\net237[2] ), .a(rnw[1]), .b(net269) );
    and2_1 \U128_14_/U8  ( .x(\net237[1] ), .a(size[2]), .b(net269) );
    and2_1 \U128_15_/U8  ( .x(\net237[0] ), .a(size[3]), .b(net269) );
    and2_1 \U37_0_/U8  ( .x(\net234[15] ), .a(addr[8]), .b(net259) );
    and2_1 \U37_1_/U8  ( .x(\net234[14] ), .a(addr[9]), .b(net259) );
    and2_1 \U37_2_/U8  ( .x(\net234[13] ), .a(addr[10]), .b(net259) );
    and2_1 \U37_3_/U8  ( .x(\net234[12] ), .a(addr[11]), .b(net259) );
    and2_1 \U37_4_/U8  ( .x(\net234[11] ), .a(addr[12]), .b(net259) );
    and2_1 \U37_5_/U8  ( .x(\net234[10] ), .a(addr[13]), .b(net259) );
    and2_1 \U37_6_/U8  ( .x(\net234[9] ), .a(addr[14]), .b(net259) );
    and2_1 \U37_7_/U8  ( .x(\net234[8] ), .a(addr[15]), .b(net259) );
    and2_1 \U37_8_/U8  ( .x(\net234[7] ), .a(addr[40]), .b(net259) );
    and2_1 \U37_9_/U8  ( .x(\net234[6] ), .a(addr[41]), .b(net259) );
    and2_1 \U37_10_/U8  ( .x(\net234[5] ), .a(addr[42]), .b(net259) );
    and2_1 \U37_11_/U8  ( .x(\net234[4] ), .a(addr[43]), .b(net259) );
    and2_1 \U37_12_/U8  ( .x(\net234[3] ), .a(addr[44]), .b(net259) );
    and2_1 \U37_13_/U8  ( .x(\net234[2] ), .a(addr[45]), .b(net259) );
    and2_1 \U37_14_/U8  ( .x(\net234[1] ), .a(addr[46]), .b(net259) );
    and2_1 \U37_15_/U8  ( .x(\net234[0] ), .a(addr[47]), .b(net259) );
    and2_1 \U33_0_/U8  ( .x(\net231[15] ), .a(addr[16]), .b(net253) );
    and2_1 \U33_1_/U8  ( .x(\net231[14] ), .a(addr[17]), .b(net253) );
    and2_1 \U33_2_/U8  ( .x(\net231[13] ), .a(addr[18]), .b(net253) );
    and2_1 \U33_3_/U8  ( .x(\net231[12] ), .a(addr[19]), .b(net253) );
    and2_1 \U33_4_/U8  ( .x(\net231[11] ), .a(addr[20]), .b(net253) );
    and2_1 \U33_5_/U8  ( .x(\net231[10] ), .a(addr[21]), .b(net253) );
    and2_1 \U33_6_/U8  ( .x(\net231[9] ), .a(addr[22]), .b(net253) );
    and2_1 \U33_7_/U8  ( .x(\net231[8] ), .a(addr[23]), .b(net253) );
    and2_1 \U33_8_/U8  ( .x(\net231[7] ), .a(addr[48]), .b(net253) );
    and2_1 \U33_9_/U8  ( .x(\net231[6] ), .a(addr[49]), .b(net253) );
    and2_1 \U33_10_/U8  ( .x(\net231[5] ), .a(addr[50]), .b(net253) );
    and2_1 \U33_11_/U8  ( .x(\net231[4] ), .a(addr[51]), .b(net253) );
    and2_1 \U33_12_/U8  ( .x(\net231[3] ), .a(addr[52]), .b(net253) );
    and2_1 \U33_13_/U8  ( .x(\net231[2] ), .a(addr[53]), .b(net253) );
    and2_1 \U33_14_/U8  ( .x(\net231[1] ), .a(addr[54]), .b(net253) );
    and2_1 \U33_15_/U8  ( .x(\net231[0] ), .a(addr[55]), .b(net253) );
    and2_1 \U81_0_/U8  ( .x(\net228[15] ), .a(wd[24]), .b(net255) );
    and2_1 \U81_1_/U8  ( .x(\net228[14] ), .a(wd[25]), .b(net255) );
    and2_1 \U81_2_/U8  ( .x(\net228[13] ), .a(wd[26]), .b(net255) );
    and2_1 \U81_3_/U8  ( .x(\net228[12] ), .a(wd[27]), .b(net255) );
    and2_1 \U81_4_/U8  ( .x(\net228[11] ), .a(wd[28]), .b(net255) );
    and2_1 \U81_5_/U8  ( .x(\net228[10] ), .a(wd[29]), .b(net255) );
    and2_1 \U81_6_/U8  ( .x(\net228[9] ), .a(wd[30]), .b(net255) );
    and2_1 \U81_7_/U8  ( .x(\net228[8] ), .a(wd[31]), .b(net255) );
    and2_1 \U81_8_/U8  ( .x(\net228[7] ), .a(wd[56]), .b(net255) );
    and2_1 \U81_9_/U8  ( .x(\net228[6] ), .a(wd[57]), .b(net255) );
    and2_1 \U81_10_/U8  ( .x(\net228[5] ), .a(wd[58]), .b(net255) );
    and2_1 \U81_11_/U8  ( .x(\net228[4] ), .a(wd[59]), .b(net255) );
    and2_1 \U81_12_/U8  ( .x(\net228[3] ), .a(wd[60]), .b(net255) );
    and2_1 \U81_13_/U8  ( .x(\net228[2] ), .a(wd[61]), .b(net255) );
    and2_1 \U81_14_/U8  ( .x(\net228[1] ), .a(wd[62]), .b(net255) );
    and2_1 \U81_15_/U8  ( .x(\net228[0] ), .a(wd[63]), .b(net255) );
    and2_1 \U34_0_/U8  ( .x(\net225[15] ), .a(addr[0]), .b(net251) );
    and2_1 \U34_1_/U8  ( .x(\net225[14] ), .a(addr[1]), .b(net251) );
    and2_1 \U34_2_/U8  ( .x(\net225[13] ), .a(addr[2]), .b(net251) );
    and2_1 \U34_3_/U8  ( .x(\net225[12] ), .a(addr[3]), .b(net251) );
    and2_1 \U34_4_/U8  ( .x(\net225[11] ), .a(addr[4]), .b(net251) );
    and2_1 \U34_5_/U8  ( .x(\net225[10] ), .a(addr[5]), .b(net251) );
    and2_1 \U34_6_/U8  ( .x(\net225[9] ), .a(addr[6]), .b(net251) );
    and2_1 \U34_7_/U8  ( .x(\net225[8] ), .a(addr[7]), .b(net251) );
    and2_1 \U34_8_/U8  ( .x(\net225[7] ), .a(addr[32]), .b(net251) );
    and2_1 \U34_9_/U8  ( .x(\net225[6] ), .a(addr[33]), .b(net251) );
    and2_1 \U34_10_/U8  ( .x(\net225[5] ), .a(addr[34]), .b(net251) );
    and2_1 \U34_11_/U8  ( .x(\net225[4] ), .a(addr[35]), .b(net251) );
    and2_1 \U34_12_/U8  ( .x(\net225[3] ), .a(addr[36]), .b(net251) );
    and2_1 \U34_13_/U8  ( .x(\net225[2] ), .a(addr[37]), .b(net251) );
    and2_1 \U34_14_/U8  ( .x(\net225[1] ), .a(addr[38]), .b(net251) );
    and2_1 \U34_15_/U8  ( .x(\net225[0] ), .a(addr[39]), .b(net251) );
    and2_1 \U30_0_/U8  ( .x(\net222[15] ), .a(addr[24]), .b(net261) );
    and2_1 \U30_1_/U8  ( .x(\net222[14] ), .a(addr[25]), .b(net261) );
    and2_1 \U30_2_/U8  ( .x(\net222[13] ), .a(addr[26]), .b(net261) );
    and2_1 \U30_3_/U8  ( .x(\net222[12] ), .a(addr[27]), .b(net261) );
    and2_1 \U30_4_/U8  ( .x(\net222[11] ), .a(addr[28]), .b(net261) );
    and2_1 \U30_5_/U8  ( .x(\net222[10] ), .a(addr[29]), .b(net261) );
    and2_1 \U30_6_/U8  ( .x(\net222[9] ), .a(addr[30]), .b(net261) );
    and2_1 \U30_7_/U8  ( .x(\net222[8] ), .a(addr[31]), .b(net261) );
    and2_1 \U30_8_/U8  ( .x(\net222[7] ), .a(addr[56]), .b(net261) );
    and2_1 \U30_9_/U8  ( .x(\net222[6] ), .a(addr[57]), .b(net261) );
    and2_1 \U30_10_/U8  ( .x(\net222[5] ), .a(addr[58]), .b(net261) );
    and2_1 \U30_11_/U8  ( .x(\net222[4] ), .a(addr[59]), .b(net261) );
    and2_1 \U30_12_/U8  ( .x(\net222[3] ), .a(addr[60]), .b(net261) );
    and2_1 \U30_13_/U8  ( .x(\net222[2] ), .a(addr[61]), .b(net261) );
    and2_1 \U30_14_/U8  ( .x(\net222[1] ), .a(addr[62]), .b(net261) );
    and2_1 \U30_15_/U8  ( .x(\net222[0] ), .a(addr[63]), .b(net261) );
    and2_1 \U82_0_/U8  ( .x(\net219[15] ), .a(wd[0]), .b(net249) );
    and2_1 \U82_1_/U8  ( .x(\net219[14] ), .a(wd[1]), .b(net249) );
    and2_1 \U82_2_/U8  ( .x(\net219[13] ), .a(wd[2]), .b(net249) );
    and2_1 \U82_3_/U8  ( .x(\net219[12] ), .a(wd[3]), .b(net249) );
    and2_1 \U82_4_/U8  ( .x(\net219[11] ), .a(wd[4]), .b(net249) );
    and2_1 \U82_5_/U8  ( .x(\net219[10] ), .a(wd[5]), .b(net249) );
    and2_1 \U82_6_/U8  ( .x(\net219[9] ), .a(wd[6]), .b(net249) );
    and2_1 \U82_7_/U8  ( .x(\net219[8] ), .a(wd[7]), .b(net249) );
    and2_1 \U82_8_/U8  ( .x(\net219[7] ), .a(wd[32]), .b(net249) );
    and2_1 \U82_9_/U8  ( .x(\net219[6] ), .a(wd[33]), .b(net249) );
    and2_1 \U82_10_/U8  ( .x(\net219[5] ), .a(wd[34]), .b(net249) );
    and2_1 \U82_11_/U8  ( .x(\net219[4] ), .a(wd[35]), .b(net249) );
    and2_1 \U82_12_/U8  ( .x(\net219[3] ), .a(wd[36]), .b(net249) );
    and2_1 \U82_13_/U8  ( .x(\net219[2] ), .a(wd[37]), .b(net249) );
    and2_1 \U82_14_/U8  ( .x(\net219[1] ), .a(wd[38]), .b(net249) );
    and2_1 \U82_15_/U8  ( .x(\net219[0] ), .a(wd[39]), .b(net249) );
    inv_1 \U40_0_/U3  ( .x(\U40_0_/n3 ), .a(\net225[15] ) );
    inv_1 \U40_0_/U4  ( .x(\U40_0_/n4 ), .a(\net234[15] ) );
    inv_1 \U40_0_/U5  ( .x(\net217[15] ), .a(\U40_0_/n5 ) );
    inv_1 \U40_1_/U3  ( .x(\U40_1_/n3 ), .a(\net225[14] ) );
    inv_1 \U40_1_/U4  ( .x(\U40_1_/n4 ), .a(\net234[14] ) );
    inv_1 \U40_1_/U5  ( .x(\net217[14] ), .a(\U40_1_/n5 ) );
    inv_1 \U40_2_/U3  ( .x(\U40_2_/n3 ), .a(\net225[13] ) );
    inv_1 \U40_2_/U4  ( .x(\U40_2_/n4 ), .a(\net234[13] ) );
    inv_1 \U40_2_/U5  ( .x(\net217[13] ), .a(\U40_2_/n5 ) );
    inv_1 \U40_3_/U3  ( .x(\U40_3_/n3 ), .a(\net225[12] ) );
    inv_1 \U40_3_/U4  ( .x(\U40_3_/n4 ), .a(\net234[12] ) );
    inv_1 \U40_3_/U5  ( .x(\net217[12] ), .a(\U40_3_/n5 ) );
    inv_1 \U40_4_/U3  ( .x(\U40_4_/n3 ), .a(\net225[11] ) );
    inv_1 \U40_4_/U4  ( .x(\U40_4_/n4 ), .a(\net234[11] ) );
    inv_1 \U40_4_/U5  ( .x(\net217[11] ), .a(\U40_4_/n5 ) );
    inv_1 \U40_5_/U3  ( .x(\U40_5_/n3 ), .a(\net225[10] ) );
    inv_1 \U40_5_/U4  ( .x(\U40_5_/n4 ), .a(\net234[10] ) );
    inv_1 \U40_5_/U5  ( .x(\net217[10] ), .a(\U40_5_/n5 ) );
    inv_1 \U40_6_/U3  ( .x(\U40_6_/n3 ), .a(\net225[9] ) );
    inv_1 \U40_6_/U4  ( .x(\U40_6_/n4 ), .a(\net234[9] ) );
    inv_1 \U40_6_/U5  ( .x(\net217[9] ), .a(\U40_6_/n5 ) );
    inv_1 \U40_7_/U3  ( .x(\U40_7_/n3 ), .a(\net225[8] ) );
    inv_1 \U40_7_/U4  ( .x(\U40_7_/n4 ), .a(\net234[8] ) );
    inv_1 \U40_7_/U5  ( .x(\net217[8] ), .a(\U40_7_/n5 ) );
    inv_1 \U40_8_/U3  ( .x(\U40_8_/n3 ), .a(\net225[7] ) );
    inv_1 \U40_8_/U4  ( .x(\U40_8_/n4 ), .a(\net234[7] ) );
    inv_1 \U40_8_/U5  ( .x(\net217[7] ), .a(\U40_8_/n5 ) );
    inv_1 \U40_9_/U3  ( .x(\U40_9_/n3 ), .a(\net225[6] ) );
    inv_1 \U40_9_/U4  ( .x(\U40_9_/n4 ), .a(\net234[6] ) );
    inv_1 \U40_9_/U5  ( .x(\net217[6] ), .a(\U40_9_/n5 ) );
    inv_1 \U40_10_/U3  ( .x(\U40_10_/n3 ), .a(\net225[5] ) );
    inv_1 \U40_10_/U4  ( .x(\U40_10_/n4 ), .a(\net234[5] ) );
    inv_1 \U40_10_/U5  ( .x(\net217[5] ), .a(\U40_10_/n5 ) );
    inv_1 \U40_11_/U3  ( .x(\U40_11_/n3 ), .a(\net225[4] ) );
    inv_1 \U40_11_/U4  ( .x(\U40_11_/n4 ), .a(\net234[4] ) );
    inv_1 \U40_11_/U5  ( .x(\net217[4] ), .a(\U40_11_/n5 ) );
    inv_1 \U40_12_/U3  ( .x(\U40_12_/n3 ), .a(\net225[3] ) );
    inv_1 \U40_12_/U4  ( .x(\U40_12_/n4 ), .a(\net234[3] ) );
    inv_1 \U40_12_/U5  ( .x(\net217[3] ), .a(\U40_12_/n5 ) );
    inv_1 \U40_13_/U3  ( .x(\U40_13_/n3 ), .a(\net225[2] ) );
    inv_1 \U40_13_/U4  ( .x(\U40_13_/n4 ), .a(\net234[2] ) );
    inv_1 \U40_13_/U5  ( .x(\net217[2] ), .a(\U40_13_/n5 ) );
    inv_1 \U40_14_/U3  ( .x(\U40_14_/n3 ), .a(\net225[1] ) );
    inv_1 \U40_14_/U4  ( .x(\U40_14_/n4 ), .a(\net234[1] ) );
    inv_1 \U40_14_/U5  ( .x(\net217[1] ), .a(\U40_14_/n5 ) );
    inv_1 \U40_15_/U3  ( .x(\U40_15_/n3 ), .a(\net225[0] ) );
    inv_1 \U40_15_/U4  ( .x(\U40_15_/n4 ), .a(\net234[0] ) );
    inv_1 \U40_15_/U5  ( .x(\net217[0] ), .a(\U40_15_/n5 ) );
    and4_1 \U14_0_/U16  ( .x(\U14_0_/n5 ), .a(\U14_0_/n1 ), .b(\U14_0_/n2 ), 
        .c(\U14_0_/n3 ), .d(\U14_0_/n4 ) );
    inv_1 \U14_0_/U1  ( .x(\U14_0_/n1 ), .a(\net231[15] ) );
    inv_1 \U14_0_/U2  ( .x(\U14_0_/n2 ), .a(\net222[15] ) );
    inv_1 \U14_0_/U3  ( .x(\U14_0_/n3 ), .a(\net237[15] ) );
    inv_1 \U14_0_/U4  ( .x(\U14_0_/n4 ), .a(\net246[15] ) );
    inv_1 \U14_0_/U5  ( .x(\net212[15] ), .a(\U14_0_/n5 ) );
    and4_1 \U14_1_/U16  ( .x(\U14_1_/n5 ), .a(\U14_1_/n1 ), .b(\U14_1_/n2 ), 
        .c(\U14_1_/n3 ), .d(\U14_1_/n4 ) );
    inv_1 \U14_1_/U1  ( .x(\U14_1_/n1 ), .a(\net231[14] ) );
    inv_1 \U14_1_/U2  ( .x(\U14_1_/n2 ), .a(\net222[14] ) );
    inv_1 \U14_1_/U3  ( .x(\U14_1_/n3 ), .a(\net237[14] ) );
    inv_1 \U14_1_/U4  ( .x(\U14_1_/n4 ), .a(\net246[14] ) );
    inv_1 \U14_1_/U5  ( .x(\net212[14] ), .a(\U14_1_/n5 ) );
    and4_1 \U14_2_/U16  ( .x(\U14_2_/n5 ), .a(\U14_2_/n1 ), .b(\U14_2_/n2 ), 
        .c(\U14_2_/n3 ), .d(\U14_2_/n4 ) );
    inv_1 \U14_2_/U1  ( .x(\U14_2_/n1 ), .a(\net231[13] ) );
    inv_1 \U14_2_/U2  ( .x(\U14_2_/n2 ), .a(\net222[13] ) );
    inv_1 \U14_2_/U3  ( .x(\U14_2_/n3 ), .a(\net237[13] ) );
    inv_1 \U14_2_/U4  ( .x(\U14_2_/n4 ), .a(\net246[13] ) );
    inv_1 \U14_2_/U5  ( .x(\net212[13] ), .a(\U14_2_/n5 ) );
    and4_1 \U14_3_/U16  ( .x(\U14_3_/n5 ), .a(\U14_3_/n1 ), .b(\U14_3_/n2 ), 
        .c(\U14_3_/n3 ), .d(\U14_3_/n4 ) );
    inv_1 \U14_3_/U1  ( .x(\U14_3_/n1 ), .a(\net231[12] ) );
    inv_1 \U14_3_/U2  ( .x(\U14_3_/n2 ), .a(\net222[12] ) );
    inv_1 \U14_3_/U3  ( .x(\U14_3_/n3 ), .a(\net237[12] ) );
    inv_1 \U14_3_/U4  ( .x(\U14_3_/n4 ), .a(\net246[12] ) );
    inv_1 \U14_3_/U5  ( .x(\net212[12] ), .a(\U14_3_/n5 ) );
    and4_1 \U14_4_/U16  ( .x(\U14_4_/n5 ), .a(\U14_4_/n1 ), .b(\U14_4_/n2 ), 
        .c(\U14_4_/n3 ), .d(\U14_4_/n4 ) );
    inv_1 \U14_4_/U1  ( .x(\U14_4_/n1 ), .a(\net231[11] ) );
    inv_1 \U14_4_/U2  ( .x(\U14_4_/n2 ), .a(\net222[11] ) );
    inv_1 \U14_4_/U3  ( .x(\U14_4_/n3 ), .a(\net237[11] ) );
    inv_1 \U14_4_/U4  ( .x(\U14_4_/n4 ), .a(\net246[11] ) );
    inv_1 \U14_4_/U5  ( .x(\net212[11] ), .a(\U14_4_/n5 ) );
    and4_1 \U14_5_/U16  ( .x(\U14_5_/n5 ), .a(\U14_5_/n1 ), .b(\U14_5_/n2 ), 
        .c(\U14_5_/n3 ), .d(\U14_5_/n4 ) );
    inv_1 \U14_5_/U1  ( .x(\U14_5_/n1 ), .a(\net231[10] ) );
    inv_1 \U14_5_/U2  ( .x(\U14_5_/n2 ), .a(\net222[10] ) );
    inv_1 \U14_5_/U3  ( .x(\U14_5_/n3 ), .a(\net237[10] ) );
    inv_1 \U14_5_/U4  ( .x(\U14_5_/n4 ), .a(\net246[10] ) );
    inv_1 \U14_5_/U5  ( .x(\net212[10] ), .a(\U14_5_/n5 ) );
    and4_1 \U14_6_/U16  ( .x(\U14_6_/n5 ), .a(\U14_6_/n1 ), .b(\U14_6_/n2 ), 
        .c(\U14_6_/n3 ), .d(\U14_6_/n4 ) );
    inv_1 \U14_6_/U1  ( .x(\U14_6_/n1 ), .a(\net231[9] ) );
    inv_1 \U14_6_/U2  ( .x(\U14_6_/n2 ), .a(\net222[9] ) );
    inv_1 \U14_6_/U3  ( .x(\U14_6_/n3 ), .a(\net237[9] ) );
    inv_1 \U14_6_/U4  ( .x(\U14_6_/n4 ), .a(\net246[9] ) );
    inv_1 \U14_6_/U5  ( .x(\net212[9] ), .a(\U14_6_/n5 ) );
    and4_1 \U14_7_/U16  ( .x(\U14_7_/n5 ), .a(\U14_7_/n1 ), .b(\U14_7_/n2 ), 
        .c(\U14_7_/n3 ), .d(\U14_7_/n4 ) );
    inv_1 \U14_7_/U1  ( .x(\U14_7_/n1 ), .a(\net231[8] ) );
    inv_1 \U14_7_/U2  ( .x(\U14_7_/n2 ), .a(\net222[8] ) );
    inv_1 \U14_7_/U3  ( .x(\U14_7_/n3 ), .a(\net237[8] ) );
    inv_1 \U14_7_/U4  ( .x(\U14_7_/n4 ), .a(\net246[8] ) );
    inv_1 \U14_7_/U5  ( .x(\net212[8] ), .a(\U14_7_/n5 ) );
    and4_1 \U14_8_/U16  ( .x(\U14_8_/n5 ), .a(\U14_8_/n1 ), .b(\U14_8_/n2 ), 
        .c(\U14_8_/n3 ), .d(\U14_8_/n4 ) );
    inv_1 \U14_8_/U1  ( .x(\U14_8_/n1 ), .a(\net231[7] ) );
    inv_1 \U14_8_/U2  ( .x(\U14_8_/n2 ), .a(\net222[7] ) );
    inv_1 \U14_8_/U3  ( .x(\U14_8_/n3 ), .a(\net237[7] ) );
    inv_1 \U14_8_/U4  ( .x(\U14_8_/n4 ), .a(\net246[7] ) );
    inv_1 \U14_8_/U5  ( .x(\net212[7] ), .a(\U14_8_/n5 ) );
    and4_1 \U14_9_/U16  ( .x(\U14_9_/n5 ), .a(\U14_9_/n1 ), .b(\U14_9_/n2 ), 
        .c(\U14_9_/n3 ), .d(\U14_9_/n4 ) );
    inv_1 \U14_9_/U1  ( .x(\U14_9_/n1 ), .a(\net231[6] ) );
    inv_1 \U14_9_/U2  ( .x(\U14_9_/n2 ), .a(\net222[6] ) );
    inv_1 \U14_9_/U3  ( .x(\U14_9_/n3 ), .a(\net237[6] ) );
    inv_1 \U14_9_/U4  ( .x(\U14_9_/n4 ), .a(\net246[6] ) );
    inv_1 \U14_9_/U5  ( .x(\net212[6] ), .a(\U14_9_/n5 ) );
    and4_1 \U14_10_/U16  ( .x(\U14_10_/n5 ), .a(\U14_10_/n1 ), .b(\U14_10_/n2 
        ), .c(\U14_10_/n3 ), .d(\U14_10_/n4 ) );
    inv_1 \U14_10_/U1  ( .x(\U14_10_/n1 ), .a(\net231[5] ) );
    inv_1 \U14_10_/U2  ( .x(\U14_10_/n2 ), .a(\net222[5] ) );
    inv_1 \U14_10_/U3  ( .x(\U14_10_/n3 ), .a(\net237[5] ) );
    inv_1 \U14_10_/U4  ( .x(\U14_10_/n4 ), .a(\net246[5] ) );
    inv_1 \U14_10_/U5  ( .x(\net212[5] ), .a(\U14_10_/n5 ) );
    inv_1 \U14_11_/U1  ( .x(\U14_11_/n1 ), .a(\net231[4] ) );
    inv_1 \U14_11_/U2  ( .x(\U14_11_/n2 ), .a(\net222[4] ) );
    inv_1 \U14_11_/U4  ( .x(\U14_11_/n4 ), .a(\net246[4] ) );
    inv_1 \U14_11_/U5  ( .x(\net212[4] ), .a(\U14_11_/n5 ) );
    inv_1 \U14_12_/U1  ( .x(\U14_12_/n1 ), .a(\net231[3] ) );
    inv_1 \U14_12_/U2  ( .x(\U14_12_/n2 ), .a(\net222[3] ) );
    inv_1 \U14_12_/U4  ( .x(\U14_12_/n4 ), .a(\net246[3] ) );
    inv_1 \U14_12_/U5  ( .x(\net212[3] ), .a(\U14_12_/n5 ) );
    and4_1 \U14_13_/U16  ( .x(\U14_13_/n5 ), .a(\U14_13_/n1 ), .b(\U14_13_/n2 
        ), .c(\U14_13_/n3 ), .d(\U14_13_/n4 ) );
    inv_1 \U14_13_/U1  ( .x(\U14_13_/n1 ), .a(\net231[2] ) );
    inv_1 \U14_13_/U2  ( .x(\U14_13_/n2 ), .a(\net222[2] ) );
    inv_1 \U14_13_/U3  ( .x(\U14_13_/n3 ), .a(\net237[2] ) );
    inv_1 \U14_13_/U4  ( .x(\U14_13_/n4 ), .a(\net246[2] ) );
    inv_1 \U14_13_/U5  ( .x(\net212[2] ), .a(\U14_13_/n5 ) );
    and4_1 \U14_14_/U16  ( .x(\U14_14_/n5 ), .a(\U14_14_/n1 ), .b(\U14_14_/n2 
        ), .c(\U14_14_/n3 ), .d(\U14_14_/n4 ) );
    inv_1 \U14_14_/U1  ( .x(\U14_14_/n1 ), .a(\net231[1] ) );
    inv_1 \U14_14_/U2  ( .x(\U14_14_/n2 ), .a(\net222[1] ) );
    inv_1 \U14_14_/U3  ( .x(\U14_14_/n3 ), .a(\net237[1] ) );
    inv_1 \U14_14_/U4  ( .x(\U14_14_/n4 ), .a(\net246[1] ) );
    inv_1 \U14_14_/U5  ( .x(\net212[1] ), .a(\U14_14_/n5 ) );
    and4_1 \U14_15_/U16  ( .x(\U14_15_/n5 ), .a(\U14_15_/n1 ), .b(\U14_15_/n2 
        ), .c(\U14_15_/n3 ), .d(\U14_15_/n4 ) );
    inv_1 \U14_15_/U1  ( .x(\U14_15_/n1 ), .a(\net231[0] ) );
    inv_1 \U14_15_/U2  ( .x(\U14_15_/n2 ), .a(\net222[0] ) );
    inv_1 \U14_15_/U3  ( .x(\U14_15_/n3 ), .a(\net237[0] ) );
    inv_1 \U14_15_/U4  ( .x(\U14_15_/n4 ), .a(\net246[0] ) );
    inv_1 \U14_15_/U5  ( .x(\net212[0] ), .a(\U14_15_/n5 ) );
    and4_1 \U91_0_/U16  ( .x(\U91_0_/n5 ), .a(\U91_0_/n1 ), .b(\U91_0_/n2 ), 
        .c(\U91_0_/n3 ), .d(\U91_0_/n4 ) );
    inv_1 \U91_0_/U1  ( .x(\U91_0_/n1 ), .a(\net219[15] ) );
    inv_1 \U91_0_/U2  ( .x(\U91_0_/n2 ), .a(\net243[15] ) );
    inv_1 \U91_0_/U3  ( .x(\U91_0_/n3 ), .a(\net240[15] ) );
    inv_1 \U91_0_/U4  ( .x(\U91_0_/n4 ), .a(\net228[15] ) );
    inv_1 \U91_0_/U5  ( .x(\net207[15] ), .a(\U91_0_/n5 ) );
    and4_1 \U91_1_/U16  ( .x(\U91_1_/n5 ), .a(\U91_1_/n1 ), .b(\U91_1_/n2 ), 
        .c(\U91_1_/n3 ), .d(\U91_1_/n4 ) );
    inv_1 \U91_1_/U1  ( .x(\U91_1_/n1 ), .a(\net219[14] ) );
    inv_1 \U91_1_/U2  ( .x(\U91_1_/n2 ), .a(\net243[14] ) );
    inv_1 \U91_1_/U3  ( .x(\U91_1_/n3 ), .a(\net240[14] ) );
    inv_1 \U91_1_/U4  ( .x(\U91_1_/n4 ), .a(\net228[14] ) );
    inv_1 \U91_1_/U5  ( .x(\net207[14] ), .a(\U91_1_/n5 ) );
    and4_1 \U91_2_/U16  ( .x(\U91_2_/n5 ), .a(\U91_2_/n1 ), .b(\U91_2_/n2 ), 
        .c(\U91_2_/n3 ), .d(\U91_2_/n4 ) );
    inv_1 \U91_2_/U1  ( .x(\U91_2_/n1 ), .a(\net219[13] ) );
    inv_1 \U91_2_/U2  ( .x(\U91_2_/n2 ), .a(\net243[13] ) );
    inv_1 \U91_2_/U3  ( .x(\U91_2_/n3 ), .a(\net240[13] ) );
    inv_1 \U91_2_/U4  ( .x(\U91_2_/n4 ), .a(\net228[13] ) );
    inv_1 \U91_2_/U5  ( .x(\net207[13] ), .a(\U91_2_/n5 ) );
    and4_1 \U91_3_/U16  ( .x(\U91_3_/n5 ), .a(\U91_3_/n1 ), .b(\U91_3_/n2 ), 
        .c(\U91_3_/n3 ), .d(\U91_3_/n4 ) );
    inv_1 \U91_3_/U1  ( .x(\U91_3_/n1 ), .a(\net219[12] ) );
    inv_1 \U91_3_/U2  ( .x(\U91_3_/n2 ), .a(\net243[12] ) );
    inv_1 \U91_3_/U3  ( .x(\U91_3_/n3 ), .a(\net240[12] ) );
    inv_1 \U91_3_/U4  ( .x(\U91_3_/n4 ), .a(\net228[12] ) );
    inv_1 \U91_3_/U5  ( .x(\net207[12] ), .a(\U91_3_/n5 ) );
    and4_1 \U91_4_/U16  ( .x(\U91_4_/n5 ), .a(\U91_4_/n1 ), .b(\U91_4_/n2 ), 
        .c(\U91_4_/n3 ), .d(\U91_4_/n4 ) );
    inv_1 \U91_4_/U1  ( .x(\U91_4_/n1 ), .a(\net219[11] ) );
    inv_1 \U91_4_/U2  ( .x(\U91_4_/n2 ), .a(\net243[11] ) );
    inv_1 \U91_4_/U3  ( .x(\U91_4_/n3 ), .a(\net240[11] ) );
    inv_1 \U91_4_/U4  ( .x(\U91_4_/n4 ), .a(\net228[11] ) );
    inv_1 \U91_4_/U5  ( .x(\net207[11] ), .a(\U91_4_/n5 ) );
    and4_1 \U91_5_/U16  ( .x(\U91_5_/n5 ), .a(\U91_5_/n1 ), .b(\U91_5_/n2 ), 
        .c(\U91_5_/n3 ), .d(\U91_5_/n4 ) );
    inv_1 \U91_5_/U1  ( .x(\U91_5_/n1 ), .a(\net219[10] ) );
    inv_1 \U91_5_/U2  ( .x(\U91_5_/n2 ), .a(\net243[10] ) );
    inv_1 \U91_5_/U3  ( .x(\U91_5_/n3 ), .a(\net240[10] ) );
    inv_1 \U91_5_/U4  ( .x(\U91_5_/n4 ), .a(\net228[10] ) );
    inv_1 \U91_5_/U5  ( .x(\net207[10] ), .a(\U91_5_/n5 ) );
    and4_1 \U91_6_/U16  ( .x(\U91_6_/n5 ), .a(\U91_6_/n1 ), .b(\U91_6_/n2 ), 
        .c(\U91_6_/n3 ), .d(\U91_6_/n4 ) );
    inv_1 \U91_6_/U1  ( .x(\U91_6_/n1 ), .a(\net219[9] ) );
    inv_1 \U91_6_/U2  ( .x(\U91_6_/n2 ), .a(\net243[9] ) );
    inv_1 \U91_6_/U3  ( .x(\U91_6_/n3 ), .a(\net240[9] ) );
    inv_1 \U91_6_/U4  ( .x(\U91_6_/n4 ), .a(\net228[9] ) );
    inv_1 \U91_6_/U5  ( .x(\net207[9] ), .a(\U91_6_/n5 ) );
    and4_1 \U91_7_/U16  ( .x(\U91_7_/n5 ), .a(\U91_7_/n1 ), .b(\U91_7_/n2 ), 
        .c(\U91_7_/n3 ), .d(\U91_7_/n4 ) );
    inv_1 \U91_7_/U1  ( .x(\U91_7_/n1 ), .a(\net219[8] ) );
    inv_1 \U91_7_/U2  ( .x(\U91_7_/n2 ), .a(\net243[8] ) );
    inv_1 \U91_7_/U3  ( .x(\U91_7_/n3 ), .a(\net240[8] ) );
    inv_1 \U91_7_/U4  ( .x(\U91_7_/n4 ), .a(\net228[8] ) );
    inv_1 \U91_7_/U5  ( .x(\net207[8] ), .a(\U91_7_/n5 ) );
    and4_1 \U91_8_/U16  ( .x(\U91_8_/n5 ), .a(\U91_8_/n1 ), .b(\U91_8_/n2 ), 
        .c(\U91_8_/n3 ), .d(\U91_8_/n4 ) );
    inv_1 \U91_8_/U1  ( .x(\U91_8_/n1 ), .a(\net219[7] ) );
    inv_1 \U91_8_/U2  ( .x(\U91_8_/n2 ), .a(\net243[7] ) );
    inv_1 \U91_8_/U3  ( .x(\U91_8_/n3 ), .a(\net240[7] ) );
    inv_1 \U91_8_/U4  ( .x(\U91_8_/n4 ), .a(\net228[7] ) );
    inv_1 \U91_8_/U5  ( .x(\net207[7] ), .a(\U91_8_/n5 ) );
    and4_1 \U91_9_/U16  ( .x(\U91_9_/n5 ), .a(\U91_9_/n1 ), .b(\U91_9_/n2 ), 
        .c(\U91_9_/n3 ), .d(\U91_9_/n4 ) );
    inv_1 \U91_9_/U1  ( .x(\U91_9_/n1 ), .a(\net219[6] ) );
    inv_1 \U91_9_/U2  ( .x(\U91_9_/n2 ), .a(\net243[6] ) );
    inv_1 \U91_9_/U3  ( .x(\U91_9_/n3 ), .a(\net240[6] ) );
    inv_1 \U91_9_/U4  ( .x(\U91_9_/n4 ), .a(\net228[6] ) );
    inv_1 \U91_9_/U5  ( .x(\net207[6] ), .a(\U91_9_/n5 ) );
    and4_1 \U91_10_/U16  ( .x(\U91_10_/n5 ), .a(\U91_10_/n1 ), .b(\U91_10_/n2 
        ), .c(\U91_10_/n3 ), .d(\U91_10_/n4 ) );
    inv_1 \U91_10_/U1  ( .x(\U91_10_/n1 ), .a(\net219[5] ) );
    inv_1 \U91_10_/U2  ( .x(\U91_10_/n2 ), .a(\net243[5] ) );
    inv_1 \U91_10_/U3  ( .x(\U91_10_/n3 ), .a(\net240[5] ) );
    inv_1 \U91_10_/U4  ( .x(\U91_10_/n4 ), .a(\net228[5] ) );
    inv_1 \U91_10_/U5  ( .x(\net207[5] ), .a(\U91_10_/n5 ) );
    and4_1 \U91_11_/U16  ( .x(\U91_11_/n5 ), .a(\U91_11_/n1 ), .b(\U91_11_/n2 
        ), .c(\U91_11_/n3 ), .d(\U91_11_/n4 ) );
    inv_1 \U91_11_/U1  ( .x(\U91_11_/n1 ), .a(\net219[4] ) );
    inv_1 \U91_11_/U2  ( .x(\U91_11_/n2 ), .a(\net243[4] ) );
    inv_1 \U91_11_/U3  ( .x(\U91_11_/n3 ), .a(\net240[4] ) );
    inv_1 \U91_11_/U4  ( .x(\U91_11_/n4 ), .a(\net228[4] ) );
    inv_1 \U91_11_/U5  ( .x(\net207[4] ), .a(\U91_11_/n5 ) );
    and4_1 \U91_12_/U16  ( .x(\U91_12_/n5 ), .a(\U91_12_/n1 ), .b(\U91_12_/n2 
        ), .c(\U91_12_/n3 ), .d(\U91_12_/n4 ) );
    inv_1 \U91_12_/U1  ( .x(\U91_12_/n1 ), .a(\net219[3] ) );
    inv_1 \U91_12_/U2  ( .x(\U91_12_/n2 ), .a(\net243[3] ) );
    inv_1 \U91_12_/U3  ( .x(\U91_12_/n3 ), .a(\net240[3] ) );
    inv_1 \U91_12_/U4  ( .x(\U91_12_/n4 ), .a(\net228[3] ) );
    inv_1 \U91_12_/U5  ( .x(\net207[3] ), .a(\U91_12_/n5 ) );
    and4_1 \U91_13_/U16  ( .x(\U91_13_/n5 ), .a(\U91_13_/n1 ), .b(\U91_13_/n2 
        ), .c(\U91_13_/n3 ), .d(\U91_13_/n4 ) );
    inv_1 \U91_13_/U1  ( .x(\U91_13_/n1 ), .a(\net219[2] ) );
    inv_1 \U91_13_/U2  ( .x(\U91_13_/n2 ), .a(\net243[2] ) );
    inv_1 \U91_13_/U3  ( .x(\U91_13_/n3 ), .a(\net240[2] ) );
    inv_1 \U91_13_/U4  ( .x(\U91_13_/n4 ), .a(\net228[2] ) );
    inv_1 \U91_13_/U5  ( .x(\net207[2] ), .a(\U91_13_/n5 ) );
    and4_1 \U91_14_/U16  ( .x(\U91_14_/n5 ), .a(\U91_14_/n1 ), .b(\U91_14_/n2 
        ), .c(\U91_14_/n3 ), .d(\U91_14_/n4 ) );
    inv_1 \U91_14_/U1  ( .x(\U91_14_/n1 ), .a(\net219[1] ) );
    inv_1 \U91_14_/U2  ( .x(\U91_14_/n2 ), .a(\net243[1] ) );
    inv_1 \U91_14_/U3  ( .x(\U91_14_/n3 ), .a(\net240[1] ) );
    inv_1 \U91_14_/U4  ( .x(\U91_14_/n4 ), .a(\net228[1] ) );
    inv_1 \U91_14_/U5  ( .x(\net207[1] ), .a(\U91_14_/n5 ) );
    and4_1 \U91_15_/U16  ( .x(\U91_15_/n5 ), .a(\U91_15_/n1 ), .b(\U91_15_/n2 
        ), .c(\U91_15_/n3 ), .d(\U91_15_/n4 ) );
    inv_1 \U91_15_/U1  ( .x(\U91_15_/n1 ), .a(\net219[0] ) );
    inv_1 \U91_15_/U2  ( .x(\U91_15_/n2 ), .a(\net243[0] ) );
    inv_1 \U91_15_/U3  ( .x(\U91_15_/n3 ), .a(\net240[0] ) );
    inv_1 \U91_15_/U4  ( .x(\U91_15_/n4 ), .a(\net228[0] ) );
    inv_1 \U91_15_/U5  ( .x(\net207[0] ), .a(\U91_15_/n5 ) );
    or3_2 \U93_0_/U12  ( .x(chainl[0]), .a(\net207[15] ), .b(\net217[15] ), 
        .c(\net212[15] ) );
    or3_2 \U93_1_/U12  ( .x(chainl[1]), .a(\net207[14] ), .b(\net217[14] ), 
        .c(\net212[14] ) );
    or3_2 \U93_2_/U12  ( .x(chainl[2]), .a(\net207[13] ), .b(\net217[13] ), 
        .c(\net212[13] ) );
    or3_2 \U93_3_/U12  ( .x(chainl[3]), .a(\net207[12] ), .b(\net217[12] ), 
        .c(\net212[12] ) );
    or3_2 \U93_4_/U12  ( .x(chainl[4]), .a(\net207[11] ), .b(\net217[11] ), 
        .c(\net212[11] ) );
    or3_2 \U93_5_/U12  ( .x(chainl[5]), .a(\net207[10] ), .b(\net217[10] ), 
        .c(\net212[10] ) );
    or3_2 \U93_6_/U12  ( .x(chainl[6]), .a(\net207[9] ), .b(\net217[9] ), .c(
        \net212[9] ) );
    or3_2 \U93_7_/U12  ( .x(chainl[7]), .a(\net207[8] ), .b(\net217[8] ), .c(
        \net212[8] ) );
    or3_2 \U93_8_/U12  ( .x(chainh[0]), .a(\net207[7] ), .b(\net217[7] ), .c(
        \net212[7] ) );
    or3_2 \U93_9_/U12  ( .x(chainh[1]), .a(\net207[6] ), .b(\net217[6] ), .c(
        \net212[6] ) );
    or3_2 \U93_10_/U12  ( .x(chainh[2]), .a(\net207[5] ), .b(\net217[5] ), .c(
        \net212[5] ) );
    or3_2 \U93_11_/U12  ( .x(chainh[3]), .a(\net207[4] ), .b(\net217[4] ), .c(
        \net212[4] ) );
    or3_2 \U93_12_/U12  ( .x(chainh[4]), .a(\net207[3] ), .b(\net217[3] ), .c(
        \net212[3] ) );
    or3_2 \U93_13_/U12  ( .x(chainh[5]), .a(\net207[2] ), .b(\net217[2] ), .c(
        \net212[2] ) );
    or3_2 \U93_14_/U12  ( .x(chainh[6]), .a(\net207[1] ), .b(\net217[1] ), .c(
        \net212[1] ) );
    or3_2 \U93_15_/U12  ( .x(chainh[7]), .a(\net207[0] ), .b(\net217[0] ), .c(
        \net212[0] ) );
    inv_1 \U152/U3  ( .x(net198), .a(sendreq) );
    ao23_1 \U158/U19/U21/U1/U1  ( .x(net131), .a(net132), .b(net131), .c(
        net132), .d(rnw[1]), .e(rnw[1]) );
    ao23_1 \U157/U19/U21/U1/U1  ( .x(net176), .a(net132), .b(net176), .c(
        net132), .d(rnw[0]), .e(rnw[0]) );
    ao222_1 \U123/U18/U1/U1  ( .x(net136), .a(net185), .b(net187), .c(net185), 
        .d(net136), .e(net187), .f(net136) );
    aoi21_1 \U151/U30/U1/U1  ( .x(\hdr[4] ), .a(\U151/Z ), .b(net138), .c(
        net198) );
    inv_1 \U151/U30/U1/U2  ( .x(\U151/Z ), .a(\hdr[4] ) );
    nor3_1 \U148/U21/Unr  ( .x(\U148/U21/nr ), .a(net191), .b(net136), .c(
        net293) );
    nand3_1 \U148/U21/Und  ( .x(\U148/U21/nd ), .a(net191), .b(net136), .c(
        net293) );
    oa21_1 \U148/U21/U1  ( .x(\U148/U21/n2 ), .a(\U148/U21/n2 ), .b(
        \U148/U21/nr ), .c(\U148/U21/nd ) );
    inv_1 \U148/U21/U3  ( .x(ack), .a(\U148/U21/n2 ) );
    buf_3 U1 ( .x(n1), .a(net138) );
    buf_3 U2 ( .x(net138), .a(nia) );
    buf_3 U3 ( .x(net269), .a(net146) );
    buf_3 U4 ( .x(net255), .a(\bs[5] ) );
    buf_3 U5 ( .x(net267), .a(\bs[6] ) );
    buf_3 U6 ( .x(net263), .a(\bs[7] ) );
    buf_3 U7 ( .x(net249), .a(\bs[8] ) );
    buf_3 U8 ( .x(net253), .a(\bs[2] ) );
    buf_3 U9 ( .x(net251), .a(\bs[4] ) );
    buf_3 U10 ( .x(net259), .a(\bs[3] ) );
    buf_3 U11 ( .x(net261), .a(\bs[1] ) );
    buf_3 U12 ( .x(net265), .a(\bs[0] ) );
    and2_1 U13 ( .x(\U40_2_/n5 ), .a(\U40_2_/n3 ), .b(\U40_2_/n4 ) );
    and2_1 U14 ( .x(\U40_1_/n5 ), .a(\U40_1_/n3 ), .b(\U40_1_/n4 ) );
    and2_1 U15 ( .x(\U40_9_/n5 ), .a(\U40_9_/n3 ), .b(\U40_9_/n4 ) );
    and2_1 U16 ( .x(\U40_8_/n5 ), .a(\U40_8_/n3 ), .b(\U40_8_/n4 ) );
    and2_1 U17 ( .x(\U40_13_/n5 ), .a(\U40_13_/n3 ), .b(\U40_13_/n4 ) );
    and2_1 U18 ( .x(\U40_0_/n5 ), .a(\U40_0_/n3 ), .b(\U40_0_/n4 ) );
    and2_1 U19 ( .x(\U40_5_/n5 ), .a(\U40_5_/n3 ), .b(\U40_5_/n4 ) );
    and2_1 U20 ( .x(\U40_4_/n5 ), .a(\U40_4_/n3 ), .b(\U40_4_/n4 ) );
    and3_1 U21 ( .x(\U14_12_/n5 ), .a(\U14_12_/n2 ), .b(\U14_12_/n4 ), .c(
        \U14_12_/n1 ) );
    and2_1 U22 ( .x(\U40_12_/n5 ), .a(\U40_12_/n3 ), .b(\U40_12_/n4 ) );
    and2_1 U23 ( .x(\U40_3_/n5 ), .a(\U40_3_/n3 ), .b(\U40_3_/n4 ) );
    and3_1 U24 ( .x(\U14_11_/n5 ), .a(\U14_11_/n2 ), .b(\U14_11_/n4 ), .c(
        \U14_11_/n1 ) );
    and2_1 U25 ( .x(\U40_11_/n5 ), .a(\U40_11_/n3 ), .b(\U40_11_/n4 ) );
    and2_1 U26 ( .x(\U40_10_/n5 ), .a(\U40_10_/n3 ), .b(\U40_10_/n4 ) );
    and2_1 U27 ( .x(\U40_15_/n5 ), .a(\U40_15_/n3 ), .b(\U40_15_/n4 ) );
    and2_1 U28 ( .x(\U40_7_/n5 ), .a(\U40_7_/n3 ), .b(\U40_7_/n4 ) );
    and2_1 U29 ( .x(\U40_6_/n5 ), .a(\U40_6_/n3 ), .b(\U40_6_/n4 ) );
    and2_1 U30 ( .x(\U40_14_/n5 ), .a(\U40_14_/n3 ), .b(\U40_14_/n4 ) );
endmodule


module chain_dr2fr_byte_1 ( eop_ack, ia, o, eop, ih, il, nReset, noa );
output [4:0] o;
input  [7:0] ih;
input  [7:0] il;
input  eop, nReset, noa;
output eop_ack, ia;
    wire eop_ack_wire, nbReset, eop_pass, nxa, naa, nlowack, \twobitack[0] , 
        \twobitack[1] , nhighack, \twobitack[2] , \twobitack[3] , \U1018/Z , 
        \U1270/net189 , \U1270/net192 , \U1270/net191 , net199, \U1270/net190 , 
        \U1270/U1141/Z , \U1268/net189 , \U1268/net192 , \U1268/net191 , 
        net194, \U1268/net190 , \U1268/U1141/Z , \U1224/nack[0] , \x[3] , 
        \x[2] , \U1224/nack[1] , \x[1] , \U1224/net4 , \x[0] , 
        \U1224/U1125/U28/U1/clr , asel, \U1224/U1125/U28/U1/set , 
        \U1224/U1122/U28/U1/clr , csel, nca, \U1224/U1122/U28/U1/set , 
        \U1224/U916_0_/U25/U1/clr , \a[0] , \c[0] , \U1224/U916_0_/U25/U1/ob , 
        \U1224/U916_1_/U25/U1/clr , \a[1] , \c[1] , \U1224/U916_1_/U25/U1/ob , 
        \U1224/U916_2_/U25/U1/clr , \a[2] , \c[2] , \U1224/U916_2_/U25/U1/ob , 
        \U1224/U916_3_/U25/U1/clr , \a[3] , \c[3] , \U1224/U916_3_/U25/U1/ob , 
        \U1209/nack[0] , \U1209/nack[1] , \U1209/net4 , 
        \U1209/U1125/U28/U1/clr , xsel, \U1209/U1125/U28/U1/set , 
        \U1209/U1122/U28/U1/clr , ysel, nyla, \U1209/U1122/U28/U1/set , 
        \U1209/U916_0_/U25/U1/clr , \yl[0] , \U1209/U916_0_/U25/U1/ob , 
        \U1209/U916_1_/U25/U1/clr , \yl[1] , \U1209/U916_1_/U25/U1/ob , 
        \U1209/U916_2_/U25/U1/clr , \yl[2] , \U1209/U916_2_/U25/U1/ob , 
        \U1209/U916_3_/U25/U1/clr , \yl[3] , \U1209/U916_3_/U25/U1/ob , 
        \U1213/nack[0] , \y[3] , \y[2] , \U1213/nack[1] , \y[1] , \U1213/net4 , 
        \y[0] , \U1213/U1125/U28/U1/clr , bsel, nba, \U1213/U1125/U28/U1/set , 
        \U1213/U1122/U28/U1/clr , dsel, nda, \U1213/U1122/U28/U1/set , 
        \U1213/U916_0_/U25/U1/clr , nya, \b[0] , \d[0] , 
        \U1213/U916_0_/U25/U1/ob , \U1213/U916_1_/U25/U1/clr , \b[1] , \d[1] , 
        \U1213/U916_1_/U25/U1/ob , \U1213/U916_2_/U25/U1/clr , \b[2] , \d[2] , 
        \U1213/U916_2_/U25/U1/ob , \U1213/U916_3_/U25/U1/clr , \b[3] , \d[3] , 
        \U1213/U916_3_/U25/U1/ob , \cdh[0] , \cdh[1] , \cdl[0] , \cdl[1] , 
        \cdh[2] , \cdh[3] , \cdl[2] , \cdl[3] , cg, \U1296/ng , net195, 
        \U1296/U1384/Z , \U1296/U1386/U25/U1/clr , \U1296/U1386/U25/U1/ob , dg, 
        \U1298/ng , net193, \U1298/U1384/Z , \U1298/U1386/U25/U1/clr , 
        \U1298/U1386/U25/U1/ob , bg, \U1306/ng , \U1306/U1384/Z , 
        \U1306/U1386/U25/U1/clr , \U1306/U1386/U25/U1/ob , ag, \U1295/ng , 
        \U1295/U1384/Z , \U1295/U1386/U25/U1/clr , \U1295/U1386/U25/U1/ob , 
        \U1297/s , \U1297/r , \U1297/nback , \U1297/naack , \U1297/reset , 
        \U1297/U1128/U28/U1/clr , \U1297/U1128/U28/U1/set , 
        \U1297/U1127/U28/U1/clr , \U1297/U1127/U28/U1/set , \U1300/s , 
        \U1300/r , \U1300/nback , \U1300/naack , \U1300/reset , 
        \U1300/U1128/U28/U1/clr , \U1300/U1128/U28/U1/set , 
        \U1300/U1127/U28/U1/clr , \U1300/U1127/U28/U1/set , 
        \U1289/U1150/U28/U1/clr , \U1289/bnreset , \U1289/U1150/U28/U1/set , 
        \U1289/U1152/U28/U1/clr , \U1289/U1152/U28/U1/set , 
        \U1289/U1149/U28/U1/clr , \U1289/U1149/U28/U1/set , 
        \U1289/U1151/U28/U1/clr , \U1289/U1151/U28/U1/set , 
        \U1289/U1148/net189 , \U1289/U1148/net192 , \U1289/U1148/net191 , 
        \U1289/U1148/net190 , \U1289/U1148/U1141/Z , \U1271/U1150/U28/U1/clr , 
        \U1271/bnreset , \U1271/U1150/U28/U1/set , \U1271/U1152/U28/U1/clr , 
        \U1271/U1152/U28/U1/set , \U1271/U1149/U28/U1/clr , 
        \U1271/U1149/U28/U1/set , \U1271/U1151/U28/U1/clr , 
        \U1271/U1151/U28/U1/set , \U1271/U1148/net189 , \U1271/U1148/net192 , 
        \U1271/U1148/net191 , \U1271/U1148/net190 , \U1271/U1148/U1141/Z , 
        \U1225/s , \U1225/r , \U1225/nback , \U1225/naack , \U1225/reset , 
        \U1308/nack[1] , \U1308/nack[0] ;
    assign eop_ack = eop_ack_wire;
    assign o[4] = eop_ack_wire;
    buf_2 U1231 ( .x(nbReset), .a(nReset) );
    and3_1 \U1194/U9  ( .x(eop_pass), .a(nxa), .b(naa), .c(eop) );
    ao222_1 \U1301/U18/U1/U1  ( .x(nlowack), .a(\twobitack[0] ), .b(
        \twobitack[1] ), .c(\twobitack[0] ), .d(nlowack), .e(\twobitack[1] ), 
        .f(nlowack) );
    ao222_1 \U1302/U18/U1/U1  ( .x(nhighack), .a(\twobitack[2] ), .b(
        \twobitack[3] ), .c(\twobitack[2] ), .d(nhighack), .e(\twobitack[3] ), 
        .f(nhighack) );
    aoi222_1 \U1018/U30/U1  ( .x(ia), .a(nhighack), .b(nlowack), .c(nhighack), 
        .d(\U1018/Z ), .e(nlowack), .f(\U1018/Z ) );
    inv_1 \U1018/U30/Uinv  ( .x(\U1018/Z ), .a(ia) );
    ao222_2 \U1038/U19/U1/U1  ( .x(eop_ack_wire), .a(eop_pass), .b(noa), .c(
        eop_pass), .d(eop_ack_wire), .e(noa), .f(eop_ack_wire) );
    inv_1 \U1270/U1147/U3  ( .x(\U1270/net189 ), .a(nbReset) );
    nor2_1 \U1270/U582/U5  ( .x(\U1270/net192 ), .a(il[4]), .b(ih[4]) );
    nor2_1 \U1270/U580/U5  ( .x(\U1270/net191 ), .a(il[5]), .b(ih[5]) );
    nor2_2 \U1270/U1146/U6  ( .x(net199), .a(\U1270/net190 ), .b(
        \U1270/net189 ) );
    aoi222_1 \U1270/U1141/U30/U1  ( .x(\U1270/net190 ), .a(\U1270/net191 ), 
        .b(\U1270/net192 ), .c(\U1270/net191 ), .d(\U1270/U1141/Z ), .e(
        \U1270/net192 ), .f(\U1270/U1141/Z ) );
    inv_1 \U1270/U1141/U30/Uinv  ( .x(\U1270/U1141/Z ), .a(\U1270/net190 ) );
    inv_1 \U1268/U1147/U3  ( .x(\U1268/net189 ), .a(nbReset) );
    nor2_1 \U1268/U582/U5  ( .x(\U1268/net192 ), .a(il[6]), .b(ih[6]) );
    nor2_1 \U1268/U580/U5  ( .x(\U1268/net191 ), .a(il[7]), .b(ih[7]) );
    nor2_2 \U1268/U1146/U6  ( .x(net194), .a(\U1268/net190 ), .b(
        \U1268/net189 ) );
    aoi222_1 \U1268/U1141/U30/U1  ( .x(\U1268/net190 ), .a(\U1268/net191 ), 
        .b(\U1268/net192 ), .c(\U1268/net191 ), .d(\U1268/U1141/Z ), .e(
        \U1268/net192 ), .f(\U1268/U1141/Z ) );
    inv_1 \U1268/U1141/U30/Uinv  ( .x(\U1268/U1141/Z ), .a(\U1268/net190 ) );
    nor2_1 \U1224/U1128/U5  ( .x(\U1224/nack[0] ), .a(\x[3] ), .b(\x[2] ) );
    nor3_1 \U1224/U1127/U7  ( .x(\U1224/nack[1] ), .a(\x[1] ), .b(\U1224/net4 
        ), .c(\x[0] ) );
    inv_1 \U1224/U907/U3  ( .x(\U1224/net4 ), .a(nbReset) );
    aoai211_1 \U1224/U1125/U28/U1/U1  ( .x(\U1224/U1125/U28/U1/clr ), .a(
        \U1224/nack[1] ), .b(\U1224/nack[0] ), .c(asel), .d(naa) );
    nand3_1 \U1224/U1125/U28/U1/U2  ( .x(\U1224/U1125/U28/U1/set ), .a(asel), 
        .b(\U1224/nack[1] ), .c(\U1224/nack[0] ) );
    nand2_2 \U1224/U1125/U28/U1/U3  ( .x(naa), .a(\U1224/U1125/U28/U1/clr ), 
        .b(\U1224/U1125/U28/U1/set ) );
    aoai211_1 \U1224/U1122/U28/U1/U1  ( .x(\U1224/U1122/U28/U1/clr ), .a(
        \U1224/nack[0] ), .b(\U1224/nack[1] ), .c(csel), .d(nca) );
    nand3_1 \U1224/U1122/U28/U1/U2  ( .x(\U1224/U1122/U28/U1/set ), .a(csel), 
        .b(\U1224/nack[0] ), .c(\U1224/nack[1] ) );
    nand2_2 \U1224/U1122/U28/U1/U3  ( .x(nca), .a(\U1224/U1122/U28/U1/clr ), 
        .b(\U1224/U1122/U28/U1/set ) );
    oa31_1 \U1224/U916_0_/U25/U1/Uclr  ( .x(\U1224/U916_0_/U25/U1/clr ), .a(
        nxa), .b(\a[0] ), .c(\c[0] ), .d(\x[0] ) );
    oaoi211_1 \U1224/U916_0_/U25/U1/Uaoi  ( .x(\U1224/U916_0_/U25/U1/ob ), .a(
        \a[0] ), .b(\c[0] ), .c(nxa), .d(\U1224/U916_0_/U25/U1/clr ) );
    inv_2 \U1224/U916_0_/U25/U1/Ui  ( .x(\x[0] ), .a(\U1224/U916_0_/U25/U1/ob 
        ) );
    oa31_1 \U1224/U916_1_/U25/U1/Uclr  ( .x(\U1224/U916_1_/U25/U1/clr ), .a(
        nxa), .b(\a[1] ), .c(\c[1] ), .d(\x[1] ) );
    oaoi211_1 \U1224/U916_1_/U25/U1/Uaoi  ( .x(\U1224/U916_1_/U25/U1/ob ), .a(
        \a[1] ), .b(\c[1] ), .c(nxa), .d(\U1224/U916_1_/U25/U1/clr ) );
    inv_2 \U1224/U916_1_/U25/U1/Ui  ( .x(\x[1] ), .a(\U1224/U916_1_/U25/U1/ob 
        ) );
    oa31_1 \U1224/U916_2_/U25/U1/Uclr  ( .x(\U1224/U916_2_/U25/U1/clr ), .a(
        nxa), .b(\a[2] ), .c(\c[2] ), .d(\x[2] ) );
    oaoi211_1 \U1224/U916_2_/U25/U1/Uaoi  ( .x(\U1224/U916_2_/U25/U1/ob ), .a(
        \a[2] ), .b(\c[2] ), .c(nxa), .d(\U1224/U916_2_/U25/U1/clr ) );
    inv_2 \U1224/U916_2_/U25/U1/Ui  ( .x(\x[2] ), .a(\U1224/U916_2_/U25/U1/ob 
        ) );
    oa31_1 \U1224/U916_3_/U25/U1/Uclr  ( .x(\U1224/U916_3_/U25/U1/clr ), .a(
        nxa), .b(\a[3] ), .c(\c[3] ), .d(\x[3] ) );
    oaoi211_1 \U1224/U916_3_/U25/U1/Uaoi  ( .x(\U1224/U916_3_/U25/U1/ob ), .a(
        \a[3] ), .b(\c[3] ), .c(nxa), .d(\U1224/U916_3_/U25/U1/clr ) );
    inv_2 \U1224/U916_3_/U25/U1/Ui  ( .x(\x[3] ), .a(\U1224/U916_3_/U25/U1/ob 
        ) );
    nor2_1 \U1209/U1128/U5  ( .x(\U1209/nack[0] ), .a(o[3]), .b(o[2]) );
    nor3_1 \U1209/U1127/U7  ( .x(\U1209/nack[1] ), .a(o[1]), .b(\U1209/net4 ), 
        .c(o[0]) );
    inv_1 \U1209/U907/U3  ( .x(\U1209/net4 ), .a(nbReset) );
    aoai211_1 \U1209/U1125/U28/U1/U1  ( .x(\U1209/U1125/U28/U1/clr ), .a(
        \U1209/nack[1] ), .b(\U1209/nack[0] ), .c(xsel), .d(nxa) );
    nand3_1 \U1209/U1125/U28/U1/U2  ( .x(\U1209/U1125/U28/U1/set ), .a(xsel), 
        .b(\U1209/nack[1] ), .c(\U1209/nack[0] ) );
    nand2_2 \U1209/U1125/U28/U1/U3  ( .x(nxa), .a(\U1209/U1125/U28/U1/clr ), 
        .b(\U1209/U1125/U28/U1/set ) );
    aoai211_1 \U1209/U1122/U28/U1/U1  ( .x(\U1209/U1122/U28/U1/clr ), .a(
        \U1209/nack[0] ), .b(\U1209/nack[1] ), .c(ysel), .d(nyla) );
    nand3_1 \U1209/U1122/U28/U1/U2  ( .x(\U1209/U1122/U28/U1/set ), .a(ysel), 
        .b(\U1209/nack[0] ), .c(\U1209/nack[1] ) );
    nand2_2 \U1209/U1122/U28/U1/U3  ( .x(nyla), .a(\U1209/U1122/U28/U1/clr ), 
        .b(\U1209/U1122/U28/U1/set ) );
    oa31_1 \U1209/U916_0_/U25/U1/Uclr  ( .x(\U1209/U916_0_/U25/U1/clr ), .a(
        noa), .b(\x[0] ), .c(\yl[0] ), .d(o[0]) );
    oaoi211_1 \U1209/U916_0_/U25/U1/Uaoi  ( .x(\U1209/U916_0_/U25/U1/ob ), .a(
        \x[0] ), .b(\yl[0] ), .c(noa), .d(\U1209/U916_0_/U25/U1/clr ) );
    inv_2 \U1209/U916_0_/U25/U1/Ui  ( .x(o[0]), .a(\U1209/U916_0_/U25/U1/ob )
         );
    oa31_1 \U1209/U916_1_/U25/U1/Uclr  ( .x(\U1209/U916_1_/U25/U1/clr ), .a(
        noa), .b(\x[1] ), .c(\yl[1] ), .d(o[1]) );
    oaoi211_1 \U1209/U916_1_/U25/U1/Uaoi  ( .x(\U1209/U916_1_/U25/U1/ob ), .a(
        \x[1] ), .b(\yl[1] ), .c(noa), .d(\U1209/U916_1_/U25/U1/clr ) );
    inv_2 \U1209/U916_1_/U25/U1/Ui  ( .x(o[1]), .a(\U1209/U916_1_/U25/U1/ob )
         );
    oa31_1 \U1209/U916_2_/U25/U1/Uclr  ( .x(\U1209/U916_2_/U25/U1/clr ), .a(
        noa), .b(\x[2] ), .c(\yl[2] ), .d(o[2]) );
    oaoi211_1 \U1209/U916_2_/U25/U1/Uaoi  ( .x(\U1209/U916_2_/U25/U1/ob ), .a(
        \x[2] ), .b(\yl[2] ), .c(noa), .d(\U1209/U916_2_/U25/U1/clr ) );
    inv_2 \U1209/U916_2_/U25/U1/Ui  ( .x(o[2]), .a(\U1209/U916_2_/U25/U1/ob )
         );
    oa31_1 \U1209/U916_3_/U25/U1/Uclr  ( .x(\U1209/U916_3_/U25/U1/clr ), .a(
        noa), .b(\x[3] ), .c(\yl[3] ), .d(o[3]) );
    oaoi211_1 \U1209/U916_3_/U25/U1/Uaoi  ( .x(\U1209/U916_3_/U25/U1/ob ), .a(
        \x[3] ), .b(\yl[3] ), .c(noa), .d(\U1209/U916_3_/U25/U1/clr ) );
    inv_2 \U1209/U916_3_/U25/U1/Ui  ( .x(o[3]), .a(\U1209/U916_3_/U25/U1/ob )
         );
    nor2_1 \U1213/U1128/U5  ( .x(\U1213/nack[0] ), .a(\y[3] ), .b(\y[2] ) );
    nor3_1 \U1213/U1127/U7  ( .x(\U1213/nack[1] ), .a(\y[1] ), .b(\U1213/net4 
        ), .c(\y[0] ) );
    inv_1 \U1213/U907/U3  ( .x(\U1213/net4 ), .a(nbReset) );
    aoai211_1 \U1213/U1125/U28/U1/U1  ( .x(\U1213/U1125/U28/U1/clr ), .a(
        \U1213/nack[1] ), .b(\U1213/nack[0] ), .c(bsel), .d(nba) );
    nand3_1 \U1213/U1125/U28/U1/U2  ( .x(\U1213/U1125/U28/U1/set ), .a(bsel), 
        .b(\U1213/nack[1] ), .c(\U1213/nack[0] ) );
    nand2_2 \U1213/U1125/U28/U1/U3  ( .x(nba), .a(\U1213/U1125/U28/U1/clr ), 
        .b(\U1213/U1125/U28/U1/set ) );
    aoai211_1 \U1213/U1122/U28/U1/U1  ( .x(\U1213/U1122/U28/U1/clr ), .a(
        \U1213/nack[0] ), .b(\U1213/nack[1] ), .c(dsel), .d(nda) );
    nand3_1 \U1213/U1122/U28/U1/U2  ( .x(\U1213/U1122/U28/U1/set ), .a(dsel), 
        .b(\U1213/nack[0] ), .c(\U1213/nack[1] ) );
    nand2_2 \U1213/U1122/U28/U1/U3  ( .x(nda), .a(\U1213/U1122/U28/U1/clr ), 
        .b(\U1213/U1122/U28/U1/set ) );
    oa31_1 \U1213/U916_0_/U25/U1/Uclr  ( .x(\U1213/U916_0_/U25/U1/clr ), .a(
        nya), .b(\b[0] ), .c(\d[0] ), .d(\y[0] ) );
    oaoi211_1 \U1213/U916_0_/U25/U1/Uaoi  ( .x(\U1213/U916_0_/U25/U1/ob ), .a(
        \b[0] ), .b(\d[0] ), .c(nya), .d(\U1213/U916_0_/U25/U1/clr ) );
    inv_2 \U1213/U916_0_/U25/U1/Ui  ( .x(\y[0] ), .a(\U1213/U916_0_/U25/U1/ob 
        ) );
    oa31_1 \U1213/U916_1_/U25/U1/Uclr  ( .x(\U1213/U916_1_/U25/U1/clr ), .a(
        nya), .b(\b[1] ), .c(\d[1] ), .d(\y[1] ) );
    oaoi211_1 \U1213/U916_1_/U25/U1/Uaoi  ( .x(\U1213/U916_1_/U25/U1/ob ), .a(
        \b[1] ), .b(\d[1] ), .c(nya), .d(\U1213/U916_1_/U25/U1/clr ) );
    inv_2 \U1213/U916_1_/U25/U1/Ui  ( .x(\y[1] ), .a(\U1213/U916_1_/U25/U1/ob 
        ) );
    oa31_1 \U1213/U916_2_/U25/U1/Uclr  ( .x(\U1213/U916_2_/U25/U1/clr ), .a(
        nya), .b(\b[2] ), .c(\d[2] ), .d(\y[2] ) );
    oaoi211_1 \U1213/U916_2_/U25/U1/Uaoi  ( .x(\U1213/U916_2_/U25/U1/ob ), .a(
        \b[2] ), .b(\d[2] ), .c(nya), .d(\U1213/U916_2_/U25/U1/clr ) );
    inv_2 \U1213/U916_2_/U25/U1/Ui  ( .x(\y[2] ), .a(\U1213/U916_2_/U25/U1/ob 
        ) );
    oa31_1 \U1213/U916_3_/U25/U1/Uclr  ( .x(\U1213/U916_3_/U25/U1/clr ), .a(
        nya), .b(\b[3] ), .c(\d[3] ), .d(\y[3] ) );
    oaoi211_1 \U1213/U916_3_/U25/U1/Uaoi  ( .x(\U1213/U916_3_/U25/U1/ob ), .a(
        \b[3] ), .b(\d[3] ), .c(nya), .d(\U1213/U916_3_/U25/U1/clr ) );
    inv_2 \U1213/U916_3_/U25/U1/Ui  ( .x(\y[3] ), .a(\U1213/U916_3_/U25/U1/ob 
        ) );
    and3_2 \U1210/U1138/U9  ( .x(\d[3] ), .a(\cdh[0] ), .b(nda), .c(\cdh[1] )
         );
    and3_2 \U1210/U1137/U9  ( .x(\d[2] ), .a(\cdl[0] ), .b(nda), .c(\cdh[1] )
         );
    and3_2 \U1210/U1139/U9  ( .x(\d[1] ), .a(\cdh[0] ), .b(nda), .c(\cdl[1] )
         );
    and3_2 \U1210/U1136/U9  ( .x(\d[0] ), .a(\cdl[0] ), .b(nda), .c(\cdl[1] )
         );
    and3_2 \U1162/U1138/U9  ( .x(\a[3] ), .a(ih[6]), .b(naa), .c(ih[7]) );
    and3_2 \U1162/U1137/U9  ( .x(\a[2] ), .a(il[6]), .b(naa), .c(ih[7]) );
    and3_2 \U1162/U1139/U9  ( .x(\a[1] ), .a(ih[6]), .b(naa), .c(il[7]) );
    and3_2 \U1162/U1136/U9  ( .x(\a[0] ), .a(il[6]), .b(naa), .c(il[7]) );
    and3_2 \U1211/U1138/U9  ( .x(\b[3] ), .a(ih[4]), .b(nba), .c(ih[5]) );
    and3_2 \U1211/U1137/U9  ( .x(\b[2] ), .a(il[4]), .b(nba), .c(ih[5]) );
    and3_2 \U1211/U1139/U9  ( .x(\b[1] ), .a(ih[4]), .b(nba), .c(il[5]) );
    and3_2 \U1211/U1136/U9  ( .x(\b[0] ), .a(il[4]), .b(nba), .c(il[5]) );
    and3_2 \U1163/U1138/U9  ( .x(\c[3] ), .a(\cdh[2] ), .b(nca), .c(\cdh[3] )
         );
    and3_2 \U1163/U1137/U9  ( .x(\c[2] ), .a(\cdl[2] ), .b(nca), .c(\cdh[3] )
         );
    and3_2 \U1163/U1139/U9  ( .x(\c[1] ), .a(\cdh[2] ), .b(nca), .c(\cdl[3] )
         );
    and3_2 \U1163/U1136/U9  ( .x(\c[0] ), .a(\cdl[2] ), .b(nca), .c(\cdl[3] )
         );
    and2_1 \U1296/U1385/U8  ( .x(cg), .a(nbReset), .b(\U1296/ng ) );
    aoi222_1 \U1296/U1384/U30/U1  ( .x(\U1296/ng ), .a(nca), .b(net195), .c(
        nca), .d(\U1296/U1384/Z ), .e(net195), .f(\U1296/U1384/Z ) );
    inv_1 \U1296/U1384/U30/Uinv  ( .x(\U1296/U1384/Z ), .a(\U1296/ng ) );
    oa31_1 \U1296/U1386/U25/U1/Uclr  ( .x(\U1296/U1386/U25/U1/clr ), .a(
        \twobitack[2] ), .b(cg), .c(nca), .d(net195) );
    oaoi211_1 \U1296/U1386/U25/U1/Uaoi  ( .x(\U1296/U1386/U25/U1/ob ), .a(cg), 
        .b(nca), .c(\twobitack[2] ), .d(\U1296/U1386/U25/U1/clr ) );
    inv_2 \U1296/U1386/U25/U1/Ui  ( .x(net195), .a(\U1296/U1386/U25/U1/ob ) );
    and2_1 \U1298/U1385/U8  ( .x(dg), .a(nbReset), .b(\U1298/ng ) );
    aoi222_1 \U1298/U1384/U30/U1  ( .x(\U1298/ng ), .a(nda), .b(net193), .c(
        nda), .d(\U1298/U1384/Z ), .e(net193), .f(\U1298/U1384/Z ) );
    inv_1 \U1298/U1384/U30/Uinv  ( .x(\U1298/U1384/Z ), .a(\U1298/ng ) );
    oa31_1 \U1298/U1386/U25/U1/Uclr  ( .x(\U1298/U1386/U25/U1/clr ), .a(
        \twobitack[0] ), .b(dg), .c(nda), .d(net193) );
    oaoi211_1 \U1298/U1386/U25/U1/Uaoi  ( .x(\U1298/U1386/U25/U1/ob ), .a(dg), 
        .b(nda), .c(\twobitack[0] ), .d(\U1298/U1386/U25/U1/clr ) );
    inv_2 \U1298/U1386/U25/U1/Ui  ( .x(net193), .a(\U1298/U1386/U25/U1/ob ) );
    and2_1 \U1306/U1385/U8  ( .x(bg), .a(nbReset), .b(\U1306/ng ) );
    aoi222_1 \U1306/U1384/U30/U1  ( .x(\U1306/ng ), .a(nba), .b(\twobitack[1] 
        ), .c(nba), .d(\U1306/U1384/Z ), .e(\twobitack[1] ), .f(
        \U1306/U1384/Z ) );
    inv_1 \U1306/U1384/U30/Uinv  ( .x(\U1306/U1384/Z ), .a(\U1306/ng ) );
    oa31_1 \U1306/U1386/U25/U1/Uclr  ( .x(\U1306/U1386/U25/U1/clr ), .a(net199
        ), .b(bg), .c(nba), .d(\twobitack[1] ) );
    oaoi211_1 \U1306/U1386/U25/U1/Uaoi  ( .x(\U1306/U1386/U25/U1/ob ), .a(bg), 
        .b(nba), .c(net199), .d(\U1306/U1386/U25/U1/clr ) );
    inv_2 \U1306/U1386/U25/U1/Ui  ( .x(\twobitack[1] ), .a(
        \U1306/U1386/U25/U1/ob ) );
    and2_1 \U1295/U1385/U8  ( .x(ag), .a(nbReset), .b(\U1295/ng ) );
    aoi222_1 \U1295/U1384/U30/U1  ( .x(\U1295/ng ), .a(naa), .b(\twobitack[3] 
        ), .c(naa), .d(\U1295/U1384/Z ), .e(\twobitack[3] ), .f(
        \U1295/U1384/Z ) );
    inv_1 \U1295/U1384/U30/Uinv  ( .x(\U1295/U1384/Z ), .a(\U1295/ng ) );
    oa31_1 \U1295/U1386/U25/U1/Uclr  ( .x(\U1295/U1386/U25/U1/clr ), .a(net194
        ), .b(ag), .c(naa), .d(\twobitack[3] ) );
    oaoi211_1 \U1295/U1386/U25/U1/Uaoi  ( .x(\U1295/U1386/U25/U1/ob ), .a(ag), 
        .b(naa), .c(net194), .d(\U1295/U1386/U25/U1/clr ) );
    inv_2 \U1295/U1386/U25/U1/Ui  ( .x(\twobitack[3] ), .a(
        \U1295/U1386/U25/U1/ob ) );
    nand2_1 \U1297/U1131/U5  ( .x(\U1297/s ), .a(\U1297/r ), .b(\U1297/nback )
         );
    nand2_1 \U1297/U1103/U5  ( .x(\U1297/r ), .a(\U1297/naack ), .b(\U1297/s )
         );
    inv_1 \U1297/U1111/U3  ( .x(\U1297/reset ), .a(nbReset) );
    inv_1 \U1297/U1112/U3  ( .x(\U1297/naack ), .a(naa) );
    nor2_1 \U1297/U1130/U5  ( .x(\U1297/nback ), .a(nca), .b(\U1297/reset ) );
    aoai211_1 \U1297/U1128/U28/U1/U1  ( .x(\U1297/U1128/U28/U1/clr ), .a(
        \U1297/r ), .b(\U1297/naack ), .c(cg), .d(csel) );
    nand3_1 \U1297/U1128/U28/U1/U2  ( .x(\U1297/U1128/U28/U1/set ), .a(cg), 
        .b(\U1297/r ), .c(\U1297/naack ) );
    nand2_2 \U1297/U1128/U28/U1/U3  ( .x(csel), .a(\U1297/U1128/U28/U1/clr ), 
        .b(\U1297/U1128/U28/U1/set ) );
    aoai211_1 \U1297/U1127/U28/U1/U1  ( .x(\U1297/U1127/U28/U1/clr ), .a(
        \U1297/s ), .b(\U1297/nback ), .c(ag), .d(asel) );
    nand3_1 \U1297/U1127/U28/U1/U2  ( .x(\U1297/U1127/U28/U1/set ), .a(ag), 
        .b(\U1297/s ), .c(\U1297/nback ) );
    nand2_2 \U1297/U1127/U28/U1/U3  ( .x(asel), .a(\U1297/U1127/U28/U1/clr ), 
        .b(\U1297/U1127/U28/U1/set ) );
    nand2_1 \U1300/U1131/U5  ( .x(\U1300/s ), .a(\U1300/r ), .b(\U1300/nback )
         );
    nand2_1 \U1300/U1103/U5  ( .x(\U1300/r ), .a(\U1300/naack ), .b(\U1300/s )
         );
    inv_1 \U1300/U1111/U3  ( .x(\U1300/reset ), .a(nbReset) );
    inv_1 \U1300/U1112/U3  ( .x(\U1300/naack ), .a(nba) );
    nor2_1 \U1300/U1130/U5  ( .x(\U1300/nback ), .a(nda), .b(\U1300/reset ) );
    aoai211_1 \U1300/U1128/U28/U1/U1  ( .x(\U1300/U1128/U28/U1/clr ), .a(
        \U1300/r ), .b(\U1300/naack ), .c(dg), .d(dsel) );
    nand3_1 \U1300/U1128/U28/U1/U2  ( .x(\U1300/U1128/U28/U1/set ), .a(dg), 
        .b(\U1300/r ), .c(\U1300/naack ) );
    nand2_2 \U1300/U1128/U28/U1/U3  ( .x(dsel), .a(\U1300/U1128/U28/U1/clr ), 
        .b(\U1300/U1128/U28/U1/set ) );
    aoai211_1 \U1300/U1127/U28/U1/U1  ( .x(\U1300/U1127/U28/U1/clr ), .a(
        \U1300/s ), .b(\U1300/nback ), .c(bg), .d(bsel) );
    nand3_1 \U1300/U1127/U28/U1/U2  ( .x(\U1300/U1127/U28/U1/set ), .a(bg), 
        .b(\U1300/s ), .c(\U1300/nback ) );
    nand2_2 \U1300/U1127/U28/U1/U3  ( .x(bsel), .a(\U1300/U1127/U28/U1/clr ), 
        .b(\U1300/U1127/U28/U1/set ) );
    aoai211_1 \U1289/U1150/U28/U1/U1  ( .x(\U1289/U1150/U28/U1/clr ), .a(il[2]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdl[2] ) );
    nand3_1 \U1289/U1150/U28/U1/U2  ( .x(\U1289/U1150/U28/U1/set ), .a(net195), 
        .b(il[2]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1150/U28/U1/U3  ( .x(\cdl[2] ), .a(
        \U1289/U1150/U28/U1/clr ), .b(\U1289/U1150/U28/U1/set ) );
    aoai211_1 \U1289/U1152/U28/U1/U1  ( .x(\U1289/U1152/U28/U1/clr ), .a(il[3]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdl[3] ) );
    nand3_1 \U1289/U1152/U28/U1/U2  ( .x(\U1289/U1152/U28/U1/set ), .a(net195), 
        .b(il[3]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1152/U28/U1/U3  ( .x(\cdl[3] ), .a(
        \U1289/U1152/U28/U1/clr ), .b(\U1289/U1152/U28/U1/set ) );
    aoai211_1 \U1289/U1149/U28/U1/U1  ( .x(\U1289/U1149/U28/U1/clr ), .a(ih[2]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdh[2] ) );
    nand3_1 \U1289/U1149/U28/U1/U2  ( .x(\U1289/U1149/U28/U1/set ), .a(net195), 
        .b(ih[2]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1149/U28/U1/U3  ( .x(\cdh[2] ), .a(
        \U1289/U1149/U28/U1/clr ), .b(\U1289/U1149/U28/U1/set ) );
    aoai211_1 \U1289/U1151/U28/U1/U1  ( .x(\U1289/U1151/U28/U1/clr ), .a(ih[3]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdh[3] ) );
    nand3_1 \U1289/U1151/U28/U1/U2  ( .x(\U1289/U1151/U28/U1/set ), .a(net195), 
        .b(ih[3]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1151/U28/U1/U3  ( .x(\cdh[3] ), .a(
        \U1289/U1151/U28/U1/clr ), .b(\U1289/U1151/U28/U1/set ) );
    inv_1 \U1289/U1148/U1147/U3  ( .x(\U1289/U1148/net189 ), .a(
        \U1289/bnreset ) );
    nor2_1 \U1289/U1148/U582/U5  ( .x(\U1289/U1148/net192 ), .a(\cdl[3] ), .b(
        \cdh[3] ) );
    nor2_1 \U1289/U1148/U580/U5  ( .x(\U1289/U1148/net191 ), .a(\cdl[2] ), .b(
        \cdh[2] ) );
    nor2_2 \U1289/U1148/U1146/U6  ( .x(\twobitack[2] ), .a(
        \U1289/U1148/net190 ), .b(\U1289/U1148/net189 ) );
    aoi222_1 \U1289/U1148/U1141/U30/U1  ( .x(\U1289/U1148/net190 ), .a(
        \U1289/U1148/net191 ), .b(\U1289/U1148/net192 ), .c(
        \U1289/U1148/net191 ), .d(\U1289/U1148/U1141/Z ), .e(
        \U1289/U1148/net192 ), .f(\U1289/U1148/U1141/Z ) );
    inv_1 \U1289/U1148/U1141/U30/Uinv  ( .x(\U1289/U1148/U1141/Z ), .a(
        \U1289/U1148/net190 ) );
    aoai211_1 \U1271/U1150/U28/U1/U1  ( .x(\U1271/U1150/U28/U1/clr ), .a(il[0]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdl[0] ) );
    nand3_1 \U1271/U1150/U28/U1/U2  ( .x(\U1271/U1150/U28/U1/set ), .a(net193), 
        .b(il[0]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1150/U28/U1/U3  ( .x(\cdl[0] ), .a(
        \U1271/U1150/U28/U1/clr ), .b(\U1271/U1150/U28/U1/set ) );
    aoai211_1 \U1271/U1152/U28/U1/U1  ( .x(\U1271/U1152/U28/U1/clr ), .a(il[1]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdl[1] ) );
    nand3_1 \U1271/U1152/U28/U1/U2  ( .x(\U1271/U1152/U28/U1/set ), .a(net193), 
        .b(il[1]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1152/U28/U1/U3  ( .x(\cdl[1] ), .a(
        \U1271/U1152/U28/U1/clr ), .b(\U1271/U1152/U28/U1/set ) );
    aoai211_1 \U1271/U1149/U28/U1/U1  ( .x(\U1271/U1149/U28/U1/clr ), .a(ih[0]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdh[0] ) );
    nand3_1 \U1271/U1149/U28/U1/U2  ( .x(\U1271/U1149/U28/U1/set ), .a(net193), 
        .b(ih[0]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1149/U28/U1/U3  ( .x(\cdh[0] ), .a(
        \U1271/U1149/U28/U1/clr ), .b(\U1271/U1149/U28/U1/set ) );
    aoai211_1 \U1271/U1151/U28/U1/U1  ( .x(\U1271/U1151/U28/U1/clr ), .a(ih[1]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdh[1] ) );
    nand3_1 \U1271/U1151/U28/U1/U2  ( .x(\U1271/U1151/U28/U1/set ), .a(net193), 
        .b(ih[1]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1151/U28/U1/U3  ( .x(\cdh[1] ), .a(
        \U1271/U1151/U28/U1/clr ), .b(\U1271/U1151/U28/U1/set ) );
    inv_1 \U1271/U1148/U1147/U3  ( .x(\U1271/U1148/net189 ), .a(
        \U1271/bnreset ) );
    nor2_1 \U1271/U1148/U582/U5  ( .x(\U1271/U1148/net192 ), .a(\cdl[1] ), .b(
        \cdh[1] ) );
    nor2_1 \U1271/U1148/U580/U5  ( .x(\U1271/U1148/net191 ), .a(\cdl[0] ), .b(
        \cdh[0] ) );
    nor2_2 \U1271/U1148/U1146/U6  ( .x(\twobitack[0] ), .a(
        \U1271/U1148/net190 ), .b(\U1271/U1148/net189 ) );
    aoi222_1 \U1271/U1148/U1141/U30/U1  ( .x(\U1271/U1148/net190 ), .a(
        \U1271/U1148/net191 ), .b(\U1271/U1148/net192 ), .c(
        \U1271/U1148/net191 ), .d(\U1271/U1148/U1141/Z ), .e(
        \U1271/U1148/net192 ), .f(\U1271/U1148/U1141/Z ) );
    inv_1 \U1271/U1148/U1141/U30/Uinv  ( .x(\U1271/U1148/U1141/Z ), .a(
        \U1271/U1148/net190 ) );
    nand2_1 \U1225/U1128/U5  ( .x(\U1225/s ), .a(\U1225/r ), .b(\U1225/nback )
         );
    nand2_1 \U1225/U1103/U5  ( .x(\U1225/r ), .a(\U1225/naack ), .b(\U1225/s )
         );
    inv_1 \U1225/U1111/U3  ( .x(\U1225/reset ), .a(nbReset) );
    inv_1 \U1225/U1112/U3  ( .x(\U1225/naack ), .a(nxa) );
    nor2_1 \U1225/U1127/U5  ( .x(\U1225/nback ), .a(nyla), .b(\U1225/reset )
         );
    and2_2 \U1225/U1129/U8  ( .x(xsel), .a(\U1225/nback ), .b(\U1225/s ) );
    and2_2 \U1225/U1124/U8  ( .x(ysel), .a(\U1225/r ), .b(\U1225/naack ) );
    and3_4 \U1308/U20/U9  ( .x(nya), .a(\U1308/nack[1] ), .b(\U1308/nack[0] ), 
        .c(nbReset) );
    nor2_1 \U1308/U18/U5  ( .x(\U1308/nack[0] ), .a(\yl[3] ), .b(\yl[0] ) );
    nor2_1 \U1308/U19/U5  ( .x(\U1308/nack[1] ), .a(\yl[1] ), .b(\yl[2] ) );
    ao222_2 \U1308/U15_0_/U19/U1/U1  ( .x(\yl[0] ), .a(\y[0] ), .b(nyla), .c(
        \y[0] ), .d(\yl[0] ), .e(nyla), .f(\yl[0] ) );
    ao222_2 \U1308/U15_1_/U19/U1/U1  ( .x(\yl[1] ), .a(\y[1] ), .b(nyla), .c(
        \y[1] ), .d(\yl[1] ), .e(nyla), .f(\yl[1] ) );
    ao222_2 \U1308/U15_2_/U19/U1/U1  ( .x(\yl[2] ), .a(\y[2] ), .b(nyla), .c(
        \y[2] ), .d(\yl[2] ), .e(nyla), .f(\yl[2] ) );
    ao222_2 \U1308/U15_3_/U19/U1/U1  ( .x(\yl[3] ), .a(\y[3] ), .b(nyla), .c(
        \y[3] ), .d(\yl[3] ), .e(nyla), .f(\yl[3] ) );
    buf_3 U1 ( .x(\U1271/bnreset ), .a(nbReset) );
    buf_3 U2 ( .x(\U1289/bnreset ), .a(nbReset) );
endmodule


module chain_mergepackets_1 ( naa, nba, o, a, b, nReset, noa );
output [4:0] o;
input  [4:0] a;
input  [4:0] b;
input  nReset, noa;
output naa, nba;
    wire as, seta, asel, bsel, setb, reset, \noack[1] , \noack[0] , 
        \U916_0_/U25/U1/clr , \U916_0_/U25/U1/ob , \U916_1_/U25/U1/clr , 
        \U916_1_/U25/U1/ob , \U916_2_/U25/U1/clr , \U916_2_/U25/U1/ob , 
        \U916_3_/U25/U1/clr , \U916_3_/U25/U1/ob ;
    and2_1 \U1155/U8  ( .x(as), .a(seta), .b(asel) );
    nand2_1 \U1145/U5  ( .x(asel), .a(bsel), .b(seta) );
    nand2_1 \U1103/U5  ( .x(bsel), .a(setb), .b(asel) );
    inv_1 \U1135/U3  ( .x(reset), .a(nReset) );
    inv_1 \U1134/U3  ( .x(setb), .a(a[4]) );
    and3_2 \U1154/U9  ( .x(naa), .a(\noack[1] ), .b(\noack[0] ), .c(as) );
    nor3_1 \U1127/U7  ( .x(\noack[0] ), .a(o[1]), .b(reset), .c(o[0]) );
    nor2_1 \U1132/U5  ( .x(\noack[1] ), .a(o[3]), .b(o[2]) );
    oa31_1 \U916_0_/U25/U1/Uclr  ( .x(\U916_0_/U25/U1/clr ), .a(noa), .b(a[0]), 
        .c(b[0]), .d(o[0]) );
    oaoi211_1 \U916_0_/U25/U1/Uaoi  ( .x(\U916_0_/U25/U1/ob ), .a(a[0]), .b(b
        [0]), .c(noa), .d(\U916_0_/U25/U1/clr ) );
    inv_2 \U916_0_/U25/U1/Ui  ( .x(o[0]), .a(\U916_0_/U25/U1/ob ) );
    oa31_1 \U916_1_/U25/U1/Uclr  ( .x(\U916_1_/U25/U1/clr ), .a(noa), .b(a[1]), 
        .c(b[1]), .d(o[1]) );
    oaoi211_1 \U916_1_/U25/U1/Uaoi  ( .x(\U916_1_/U25/U1/ob ), .a(a[1]), .b(b
        [1]), .c(noa), .d(\U916_1_/U25/U1/clr ) );
    inv_2 \U916_1_/U25/U1/Ui  ( .x(o[1]), .a(\U916_1_/U25/U1/ob ) );
    oa31_1 \U916_2_/U25/U1/Uclr  ( .x(\U916_2_/U25/U1/clr ), .a(noa), .b(a[2]), 
        .c(b[2]), .d(o[2]) );
    oaoi211_1 \U916_2_/U25/U1/Uaoi  ( .x(\U916_2_/U25/U1/ob ), .a(a[2]), .b(b
        [2]), .c(noa), .d(\U916_2_/U25/U1/clr ) );
    inv_2 \U916_2_/U25/U1/Ui  ( .x(o[2]), .a(\U916_2_/U25/U1/ob ) );
    oa31_1 \U916_3_/U25/U1/Uclr  ( .x(\U916_3_/U25/U1/clr ), .a(noa), .b(a[3]), 
        .c(b[3]), .d(o[3]) );
    oaoi211_1 \U916_3_/U25/U1/Uaoi  ( .x(\U916_3_/U25/U1/ob ), .a(a[3]), .b(b
        [3]), .c(noa), .d(\U916_3_/U25/U1/clr ) );
    inv_2 \U916_3_/U25/U1/Ui  ( .x(o[3]), .a(\U916_3_/U25/U1/ob ) );
    ao222_2 \U1148/U19/U1/U1  ( .x(o[4]), .a(noa), .b(b[4]), .c(noa), .d(o[4]), 
        .e(b[4]), .f(o[4]) );
    aoi21_1 \U1153/U11  ( .x(seta), .a(o[4]), .b(setb), .c(reset) );
    and3_3 U1 ( .x(nba), .a(bsel), .b(\noack[0] ), .c(\noack[1] ) );
endmodule


module initiator_dport ( cack, chaincommand, err, nchainresponseack, nrouteack, 
    rd, routetxreq, rrnw, a, chainresponse, col, crnw, itag, lock, nReset, 
    nchaincommandack, pred, rack, route, routetxack, seq, size, wd );
output [4:0] chaincommand;
output [1:0] err;
output [63:0] rd;
output [1:0] rrnw;
input  [63:0] a;
input  [4:0] chainresponse;
input  [5:0] col;
input  [1:0] crnw;
input  [9:0] itag;
input  [1:0] lock;
input  [1:0] pred;
input  [4:0] route;
input  [1:0] seq;
input  [3:0] size;
input  [63:0] wd;
input  nReset, nchaincommandack, rack, routetxack;
output cack, nchainresponseack, nrouteack, routetxreq;
    wire nircba, nResetb, responseack, rstatusack, \irbl[7] , \irbl[6] , 
        \irbl[5] , \irbl[4] , \irbl[3] , \irbl[2] , \irbl[1] , \irbl[0] , 
        \irbh[7] , \irbh[6] , \irbh[5] , \irbh[4] , \irbh[3] , \irbh[2] , 
        \irbh[1] , \irbh[0] , \rstatus[1] , \rstatus[0] , ictrlack, 
        \can_defer[0] , net116, ncstatusack, pltxreq, tok_ack, \cstatus[0] , 
        \cstatus[1] , net115, net128, pltxack, icmdack, nicba, \icbl[7] , 
        \icbl[6] , \icbl[5] , \icbl[4] , \icbl[3] , \icbl[2] , \icbl[1] , 
        \icbl[0] , \icbh[7] , \icbh[6] , \icbh[5] , \icbh[4] , \icbh[3] , 
        \icbh[2] , \icbh[1] , \icbh[0] , nipayloadack, \ipayload[4] , 
        \ipayload[3] , \ipayload[2] , \ipayload[1] , \ipayload[0] , net170, 
        reset, net165, \U1662/U28/U1/clr , \U1662/U28/U1/set ;
    chain_irdemuxNew_1 U1442 ( .err(err), .ncback(nircba), .rd(rd), .rnw(rrnw), 
        .status({\rstatus[1] , \rstatus[0] }), .cbh({\irbh[7] , \irbh[6] , 
        \irbh[5] , \irbh[4] , \irbh[3] , \irbh[2] , \irbh[1] , \irbh[0] }), 
        .cbl({\irbl[7] , \irbl[6] , \irbl[5] , \irbl[4] , \irbl[3] , \irbl[2] , 
        \irbl[1] , \irbl[0] }), .nReset(nResetb), .nack(responseack), 
        .statusack(rstatusack) );
    chain_fr2dr_byte_4 chain_decoder ( .nia(nchainresponseack), .oh({\irbh[7] , 
        \irbh[6] , \irbh[5] , \irbh[4] , \irbh[3] , \irbh[2] , \irbh[1] , 
        \irbh[0] }), .ol({\irbl[7] , \irbl[6] , \irbl[5] , \irbl[4] , 
        \irbl[3] , \irbl[2] , \irbl[1] , \irbl[0] }), .i(chainresponse), 
        .nReset(nResetb), .noa(nircba) );
    chain_ic_ctrl_1 cmd_ctrl ( .ack(ictrlack), .candefer(\can_defer[0] ), 
        .eop(net116), .nstatack(ncstatusack), .pltxreq(pltxreq), .routetxreq(
        routetxreq), .tok_ack(tok_ack), .accept(\cstatus[0] ), .candefer_ack({
        1'b0, \can_defer[0] }), .defer(\cstatus[1] ), .eopack(net115), .lock(
        lock), .nReset(net128), .pltxack(pltxack), .routetxack(routetxack), 
        .tok_err(err[1]), .tok_ok(err[0]) );
    chain_icmux_1 cmd_mux ( .ack(icmdack), .chainh({\icbh[7] , \icbh[6] , 
        \icbh[5] , \icbh[4] , \icbh[3] , \icbh[2] , \icbh[1] , \icbh[0] }), 
        .chainl({\icbl[7] , \icbl[6] , \icbl[5] , \icbl[4] , \icbl[3] , 
        \icbl[2] , \icbl[1] , \icbl[0] }), .sendack(pltxack), .addr(a), .col(
        col), .itag(itag), .lock(lock), .nReset(net128), .nia(nicba), .pred(
        pred), .rnw(crnw), .sendreq(pltxreq), .seq(seq), .size(size), .wd(wd)
         );
    chain_dr2fr_byte_1 U1604 ( .eop_ack(net115), .ia(nicba), .o({\ipayload[4] , 
        \ipayload[3] , \ipayload[2] , \ipayload[1] , \ipayload[0] }), .eop(
        net116), .ih({\icbh[7] , \icbh[6] , \icbh[5] , \icbh[4] , \icbh[3] , 
        \icbh[2] , \icbh[1] , \icbh[0] }), .il({\icbl[7] , \icbl[6] , 
        \icbl[5] , \icbl[4] , \icbl[3] , \icbl[2] , \icbl[1] , \icbl[0] }), 
        .nReset(net128), .noa(nipayloadack) );
    chain_mergepackets_1 U1605 ( .naa(nrouteack), .nba(nipayloadack), .o(
        chaincommand), .a(route), .b({\ipayload[4] , \ipayload[3] , 
        \ipayload[2] , \ipayload[1] , \ipayload[0] }), .nReset(net128), .noa(
        nchaincommandack) );
    and2_1 U1676 ( .x(cack), .a(net170), .b(nResetb) );
    inv_4 \U1643/U3  ( .x(net128), .a(reset) );
    or2_4 \U1660/U12  ( .x(net165), .a(\cstatus[0] ), .b(\cstatus[1] ) );
    or2_1 \U1661/U12  ( .x(rstatusack), .a(net165), .b(reset) );
    ao222_2 \status_pipe_0_/U19/U1/U1  ( .x(\cstatus[0] ), .a(\rstatus[0] ), 
        .b(ncstatusack), .c(\rstatus[0] ), .d(\cstatus[0] ), .e(ncstatusack), 
        .f(\cstatus[0] ) );
    ao222_2 \status_pipe_1_/U19/U1/U1  ( .x(\cstatus[1] ), .a(\rstatus[1] ), 
        .b(ncstatusack), .c(\rstatus[1] ), .d(\cstatus[1] ), .e(ncstatusack), 
        .f(\cstatus[1] ) );
    ao222_1 \U1609/U18/U1/U1  ( .x(net170), .a(ictrlack), .b(icmdack), .c(
        ictrlack), .d(net170), .e(icmdack), .f(net170) );
    aoai211_1 \U1662/U28/U1/U1  ( .x(\U1662/U28/U1/clr ), .a(rack), .b(nResetb
        ), .c(tok_ack), .d(responseack) );
    nand3_1 \U1662/U28/U1/U2  ( .x(\U1662/U28/U1/set ), .a(tok_ack), .b(rack), 
        .c(nResetb) );
    nand2_2 \U1662/U28/U1/U3  ( .x(responseack), .a(\U1662/U28/U1/clr ), .b(
        \U1662/U28/U1/set ) );
    inv_2 U1 ( .x(reset), .a(nResetb) );
    buf_3 U2 ( .x(nResetb), .a(nReset) );
endmodule


module master_if_dport ( nReset, mc_req, mc_we, mc_mult, mc_prd, mc_seq, mc_ts, 
    mc_sel, mc_adr, mc_dat, mc_ack, mr_req, mr_we, mr_err, mr_rty, mr_acc, 
    mr_ts, mr_sel, mr_dat, mr_ack, chaincommand, nchaincommandack, 
    chainresponse, nchainresponseack, e_bare, e_dm, e_im, e_wish, r_bare, r_dm, 
    r_im, r_wish, tag_id, force_bare );
input  [2:0] mc_ts;
input  [3:0] mc_sel;
input  [31:0] mc_adr;
input  [31:0] mc_dat;
output [2:0] mr_ts;
output [3:0] mr_sel;
output [31:0] mr_dat;
output [4:0] chaincommand;
input  [4:0] chainresponse;
input  [3:0] e_bare;
input  [3:0] e_dm;
input  [3:0] e_im;
input  [3:0] e_wish;
input  [3:0] r_bare;
input  [3:0] r_dm;
input  [3:0] r_im;
input  [3:0] r_wish;
input  [4:0] tag_id;
input  nReset, mc_req, mc_we, mc_mult, mc_prd, mc_seq, mr_ack, 
    nchaincommandack, force_bare;
output mc_ack, mr_req, mr_we, mr_err, mr_rty, mr_acc, nchainresponseack;
    wire reset, ci_ack, ri_ack, \ri_rnw[1] , \ri_rnw[0] , \ri_err[1] , 
        \ri_err[0] , \ri_rd[63] , \ri_rd[62] , \ri_rd[61] , \ri_rd[60] , 
        \ri_rd[59] , \ri_rd[58] , \ri_rd[57] , \ri_rd[56] , \ri_rd[55] , 
        \ri_rd[54] , \ri_rd[53] , \ri_rd[52] , \ri_rd[51] , \ri_rd[50] , 
        \ri_rd[49] , \ri_rd[48] , \ri_rd[47] , \ri_rd[46] , \ri_rd[45] , 
        \ri_rd[44] , \ri_rd[43] , \ri_rd[42] , \ri_rd[41] , \ri_rd[40] , 
        \ri_rd[39] , \ri_rd[38] , \ri_rd[37] , \ri_rd[36] , \ri_rd[35] , 
        \ri_rd[34] , \ri_rd[33] , \ri_rd[32] , \ri_rd[31] , \ri_rd[30] , 
        \ri_rd[29] , \ri_rd[28] , \ri_rd[27] , \ri_rd[26] , \ri_rd[25] , 
        \ri_rd[24] , \ri_rd[23] , \ri_rd[22] , \ri_rd[21] , \ri_rd[20] , 
        \ri_rd[19] , \ri_rd[18] , \ri_rd[17] , \ri_rd[16] , \ri_rd[15] , 
        \ri_rd[14] , \ri_rd[13] , \ri_rd[12] , \ri_rd[11] , \ri_rd[10] , 
        \ri_rd[9] , \ri_rd[8] , \ri_rd[7] , \ri_rd[6] , \ri_rd[5] , \ri_rd[4] , 
        \ri_rd[3] , \ri_rd[2] , \ri_rd[1] , \ri_rd[0] , \ci_col[5] , 
        \ci_col[4] , \ci_col[3] , \ci_col[2] , \ci_col[1] , \ci_col[0] , 
        \ci_rnw[1] , \ci_rnw[0] , \ci_a[63] , \ci_a[62] , \ci_a[61] , 
        \ci_a[60] , \ci_a[59] , \ci_a[58] , \ci_a[57] , \ci_a[56] , \ci_a[55] , 
        \ci_a[54] , \ci_a[53] , \ci_a[52] , \ci_a[51] , \ci_a[50] , \ci_a[49] , 
        \ci_a[48] , \ci_a[47] , \ci_a[46] , \ci_a[45] , \ci_a[44] , \ci_a[43] , 
        \ci_a[42] , \ci_a[41] , \ci_a[40] , \ci_a[39] , \ci_a[38] , \ci_a[37] , 
        \ci_a[36] , \ci_a[35] , \ci_a[34] , \ci_a[33] , \ci_a[32] , \ci_a[31] , 
        \ci_a[30] , \ci_a[29] , \ci_a[28] , \ci_a[27] , \ci_a[26] , \ci_a[25] , 
        \ci_a[24] , \ci_a[23] , \ci_a[22] , \ci_a[21] , \ci_a[20] , \ci_a[19] , 
        \ci_a[18] , \ci_a[17] , \ci_a[16] , \ci_a[15] , \ci_a[14] , \ci_a[13] , 
        \ci_a[12] , \ci_a[11] , \ci_a[10] , \ci_a[9] , \ci_a[8] , \ci_a[7] , 
        \ci_a[6] , \ci_a[5] , \ci_a[4] , \ci_a[3] , \ci_a[2] , \ci_a[1] , 
        \ci_a[0] , \ci_lock[1] , \ci_lock[0] , \ci_wd[63] , \ci_wd[62] , 
        \ci_wd[61] , \ci_wd[60] , \ci_wd[59] , \ci_wd[58] , \ci_wd[57] , 
        \ci_wd[56] , \ci_wd[55] , \ci_wd[54] , \ci_wd[53] , \ci_wd[52] , 
        \ci_wd[51] , \ci_wd[50] , \ci_wd[49] , \ci_wd[48] , \ci_wd[47] , 
        \ci_wd[46] , \ci_wd[45] , \ci_wd[44] , \ci_wd[43] , \ci_wd[42] , 
        \ci_wd[41] , \ci_wd[40] , \ci_wd[39] , \ci_wd[38] , \ci_wd[37] , 
        \ci_wd[36] , \ci_wd[35] , \ci_wd[34] , \ci_wd[33] , \ci_wd[32] , 
        \ci_wd[31] , \ci_wd[30] , \ci_wd[29] , \ci_wd[28] , \ci_wd[27] , 
        \ci_wd[26] , \ci_wd[25] , \ci_wd[24] , \ci_wd[23] , \ci_wd[22] , 
        \ci_wd[21] , \ci_wd[20] , \ci_wd[19] , \ci_wd[18] , \ci_wd[17] , 
        \ci_wd[16] , \ci_wd[15] , \ci_wd[14] , \ci_wd[13] , \ci_wd[12] , 
        \ci_wd[11] , \ci_wd[10] , \ci_wd[9] , \ci_wd[8] , \ci_wd[7] , 
        \ci_wd[6] , \ci_wd[5] , \ci_wd[4] , \ci_wd[3] , \ci_wd[2] , \ci_wd[1] , 
        \ci_wd[0] , \ci_itag[9] , \ci_itag[8] , \ci_itag[7] , \ci_itag[6] , 
        \ci_itag[5] , \ci_itag[4] , \ci_itag[3] , \ci_itag[2] , \ci_itag[1] , 
        \ci_itag[0] , \ci_size[3] , \ci_size[2] , \ci_size[1] , \ci_size[0] , 
        \ci_pred[1] , \ci_pred[0] , \ci_seq[1] , \ci_seq[0] , \i_rl[3] , 
        \i_rl[2] , \i_rl[1] , \i_rl[0] , \i_rh[3] , \i_rh[2] , \i_rh[1] , 
        SYNOPSYS_UNCONNECTED_2, \i_el[3] , \i_el[2] , \i_el[1] , \i_el[0] , 
        SYNOPSYS_UNCONNECTED_1, \i_eh[2] , \i_eh[1] , \i_eh[0] , routetx_ack, 
        nroute_ack, routetx_req, \route[4] , SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4, \route[1] , \route[0] ;
    assign mr_rty = 1'b0;
    assign mr_acc = 1'b0;
    assign mr_ts[2] = 1'b0;
    assign mr_ts[1] = 1'b0;
    assign mr_ts[0] = 1'b0;
    assign mr_sel[3] = 1'b0;
    assign mr_sel[2] = 1'b0;
    assign mr_sel[1] = 1'b0;
    assign mr_sel[0] = 1'b0;
    inv_2 U1 ( .x(reset), .a(nReset) );
    m2cp_dport master2chainif ( .req_in(mc_req), .ts_o(mc_ts), .sel_o(mc_sel), 
        .mult_o(mc_mult), .we_o(mc_we), .prd_o(mc_prd), .seq_o(mc_seq), 
        .adr_o(mc_adr), .dat_o(mc_dat), .ain(mc_ack), .ic_seq({\ci_seq[1] , 
        \ci_seq[0] }), .ic_pred({\ci_pred[1] , \ci_pred[0] }), .ic_size({
        \ci_size[3] , \ci_size[2] , \ci_size[1] , \ci_size[0] }), .ic_itag({
        \ci_itag[9] , \ci_itag[8] , \ci_itag[7] , \ci_itag[6] , \ci_itag[5] , 
        \ci_itag[4] , \ci_itag[3] , \ci_itag[2] , \ci_itag[1] , \ci_itag[0] }), 
        .ic_wd({\ci_wd[63] , \ci_wd[62] , \ci_wd[61] , \ci_wd[60] , 
        \ci_wd[59] , \ci_wd[58] , \ci_wd[57] , \ci_wd[56] , \ci_wd[55] , 
        \ci_wd[54] , \ci_wd[53] , \ci_wd[52] , \ci_wd[51] , \ci_wd[50] , 
        \ci_wd[49] , \ci_wd[48] , \ci_wd[47] , \ci_wd[46] , \ci_wd[45] , 
        \ci_wd[44] , \ci_wd[43] , \ci_wd[42] , \ci_wd[41] , \ci_wd[40] , 
        \ci_wd[39] , \ci_wd[38] , \ci_wd[37] , \ci_wd[36] , \ci_wd[35] , 
        \ci_wd[34] , \ci_wd[33] , \ci_wd[32] , \ci_wd[31] , \ci_wd[30] , 
        \ci_wd[29] , \ci_wd[28] , \ci_wd[27] , \ci_wd[26] , \ci_wd[25] , 
        \ci_wd[24] , \ci_wd[23] , \ci_wd[22] , \ci_wd[21] , \ci_wd[20] , 
        \ci_wd[19] , \ci_wd[18] , \ci_wd[17] , \ci_wd[16] , \ci_wd[15] , 
        \ci_wd[14] , \ci_wd[13] , \ci_wd[12] , \ci_wd[11] , \ci_wd[10] , 
        \ci_wd[9] , \ci_wd[8] , \ci_wd[7] , \ci_wd[6] , \ci_wd[5] , \ci_wd[4] , 
        \ci_wd[3] , \ci_wd[2] , \ci_wd[1] , \ci_wd[0] }), .ic_lock({
        \ci_lock[1] , \ci_lock[0] }), .ic_a({\ci_a[63] , \ci_a[62] , 
        \ci_a[61] , \ci_a[60] , \ci_a[59] , \ci_a[58] , \ci_a[57] , \ci_a[56] , 
        \ci_a[55] , \ci_a[54] , \ci_a[53] , \ci_a[52] , \ci_a[51] , \ci_a[50] , 
        \ci_a[49] , \ci_a[48] , \ci_a[47] , \ci_a[46] , \ci_a[45] , \ci_a[44] , 
        \ci_a[43] , \ci_a[42] , \ci_a[41] , \ci_a[40] , \ci_a[39] , \ci_a[38] , 
        \ci_a[37] , \ci_a[36] , \ci_a[35] , \ci_a[34] , \ci_a[33] , \ci_a[32] , 
        \ci_a[31] , \ci_a[30] , \ci_a[29] , \ci_a[28] , \ci_a[27] , \ci_a[26] , 
        \ci_a[25] , \ci_a[24] , \ci_a[23] , \ci_a[22] , \ci_a[21] , \ci_a[20] , 
        \ci_a[19] , \ci_a[18] , \ci_a[17] , \ci_a[16] , \ci_a[15] , \ci_a[14] , 
        \ci_a[13] , \ci_a[12] , \ci_a[11] , \ci_a[10] , \ci_a[9] , \ci_a[8] , 
        \ci_a[7] , \ci_a[6] , \ci_a[5] , \ci_a[4] , \ci_a[3] , \ci_a[2] , 
        \ci_a[1] , \ci_a[0] }), .ic_rnw({\ci_rnw[1] , \ci_rnw[0] }), .ic_col({
        \ci_col[5] , \ci_col[4] , \ci_col[3] , \ci_col[2] , \ci_col[1] , 
        \ci_col[0] }), .ic_ack(ci_ack), .req_out(mr_req), .we_i(mr_we), 
        .err_i(mr_err), .dat_i(mr_dat), .aout(mr_ack), .ir_rd({\ri_rd[63] , 
        \ri_rd[62] , \ri_rd[61] , \ri_rd[60] , \ri_rd[59] , \ri_rd[58] , 
        \ri_rd[57] , \ri_rd[56] , \ri_rd[55] , \ri_rd[54] , \ri_rd[53] , 
        \ri_rd[52] , \ri_rd[51] , \ri_rd[50] , \ri_rd[49] , \ri_rd[48] , 
        \ri_rd[47] , \ri_rd[46] , \ri_rd[45] , \ri_rd[44] , \ri_rd[43] , 
        \ri_rd[42] , \ri_rd[41] , \ri_rd[40] , \ri_rd[39] , \ri_rd[38] , 
        \ri_rd[37] , \ri_rd[36] , \ri_rd[35] , \ri_rd[34] , \ri_rd[33] , 
        \ri_rd[32] , \ri_rd[31] , \ri_rd[30] , \ri_rd[29] , \ri_rd[28] , 
        \ri_rd[27] , \ri_rd[26] , \ri_rd[25] , \ri_rd[24] , \ri_rd[23] , 
        \ri_rd[22] , \ri_rd[21] , \ri_rd[20] , \ri_rd[19] , \ri_rd[18] , 
        \ri_rd[17] , \ri_rd[16] , \ri_rd[15] , \ri_rd[14] , \ri_rd[13] , 
        \ri_rd[12] , \ri_rd[11] , \ri_rd[10] , \ri_rd[9] , \ri_rd[8] , 
        \ri_rd[7] , \ri_rd[6] , \ri_rd[5] , \ri_rd[4] , \ri_rd[3] , \ri_rd[2] , 
        \ri_rd[1] , \ri_rd[0] }), .ir_err({\ri_err[1] , \ri_err[0] }), 
        .ir_rnw({\ri_rnw[1] , \ri_rnw[0] }), .ir_ack(ri_ack), .tag_id(tag_id), 
        .reset(reset) );
    i_adec_dport dec ( .e_h({SYNOPSYS_UNCONNECTED_1, \i_eh[2] , \i_eh[1] , 
        \i_eh[0] }), .e_l({\i_el[3] , \i_el[2] , \i_el[1] , \i_el[0] }), .r_h(
        {\i_rh[3] , \i_rh[2] , \i_rh[1] , SYNOPSYS_UNCONNECTED_2}), .r_l({
        \i_rl[3] , \i_rl[2] , \i_rl[1] , \i_rl[0] }), .ah({\ci_a[63] , 
        \ci_a[62] , \ci_a[61] , \ci_a[60] , \ci_a[59] , \ci_a[58] , \ci_a[57] , 
        \ci_a[56] , \ci_a[55] , \ci_a[54] , \ci_a[53] , \ci_a[52] , \ci_a[51] , 
        \ci_a[50] , \ci_a[49] , \ci_a[48] , \ci_a[47] , \ci_a[46] , \ci_a[45] , 
        \ci_a[44] , \ci_a[43] , \ci_a[42] , \ci_a[41] , \ci_a[40] , \ci_a[39] , 
        \ci_a[38] , \ci_a[37] , \ci_a[36] , \ci_a[35] , \ci_a[34] , \ci_a[33] , 
        \ci_a[32] }), .al({\ci_a[31] , \ci_a[30] , \ci_a[29] , \ci_a[28] , 
        \ci_a[27] , \ci_a[26] , \ci_a[25] , \ci_a[24] , \ci_a[23] , \ci_a[22] , 
        \ci_a[21] , \ci_a[20] , \ci_a[19] , \ci_a[18] , \ci_a[17] , \ci_a[16] , 
        \ci_a[15] , \ci_a[14] , \ci_a[13] , \ci_a[12] , \ci_a[11] , \ci_a[10] , 
        \ci_a[9] , \ci_a[8] , \ci_a[7] , \ci_a[6] , \ci_a[5] , \ci_a[4] , 
        \ci_a[3] , \ci_a[2] , \ci_a[1] , \ci_a[0] }), .e_bare(e_bare), .e_dm(
        e_dm), .e_im(e_im), .e_wish(e_wish), .r_bare(r_bare), .r_dm(r_dm), 
        .r_im(r_im), .r_wish(r_wish), .force_bare(force_bare) );
    route_tx_dport rt ( .o({\route[4] , SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4, \route[1] , \route[0] }), .rtxack(routetx_ack), 
        .e_h({1'b0, \i_eh[2] , \i_eh[1] , \i_eh[0] }), .e_l({\i_el[3] , 
        \i_el[2] , \i_el[1] , \i_el[0] }), .noa(nroute_ack), .r_h({\i_rh[3] , 
        \i_rh[2] , \i_rh[1] , 1'b0}), .r_l({\i_rl[3] , \i_rl[2] , \i_rl[1] , 
        \i_rl[0] }), .rtxreq(routetx_req) );
    initiator_dport it ( .cack(ci_ack), .chaincommand(chaincommand), .err({
        \ri_err[1] , \ri_err[0] }), .nchainresponseack(nchainresponseack), 
        .nrouteack(nroute_ack), .rd({\ri_rd[63] , \ri_rd[62] , \ri_rd[61] , 
        \ri_rd[60] , \ri_rd[59] , \ri_rd[58] , \ri_rd[57] , \ri_rd[56] , 
        \ri_rd[55] , \ri_rd[54] , \ri_rd[53] , \ri_rd[52] , \ri_rd[51] , 
        \ri_rd[50] , \ri_rd[49] , \ri_rd[48] , \ri_rd[47] , \ri_rd[46] , 
        \ri_rd[45] , \ri_rd[44] , \ri_rd[43] , \ri_rd[42] , \ri_rd[41] , 
        \ri_rd[40] , \ri_rd[39] , \ri_rd[38] , \ri_rd[37] , \ri_rd[36] , 
        \ri_rd[35] , \ri_rd[34] , \ri_rd[33] , \ri_rd[32] , \ri_rd[31] , 
        \ri_rd[30] , \ri_rd[29] , \ri_rd[28] , \ri_rd[27] , \ri_rd[26] , 
        \ri_rd[25] , \ri_rd[24] , \ri_rd[23] , \ri_rd[22] , \ri_rd[21] , 
        \ri_rd[20] , \ri_rd[19] , \ri_rd[18] , \ri_rd[17] , \ri_rd[16] , 
        \ri_rd[15] , \ri_rd[14] , \ri_rd[13] , \ri_rd[12] , \ri_rd[11] , 
        \ri_rd[10] , \ri_rd[9] , \ri_rd[8] , \ri_rd[7] , \ri_rd[6] , 
        \ri_rd[5] , \ri_rd[4] , \ri_rd[3] , \ri_rd[2] , \ri_rd[1] , \ri_rd[0] 
        }), .routetxreq(routetx_req), .rrnw({\ri_rnw[1] , \ri_rnw[0] }), .a({
        \ci_a[63] , \ci_a[62] , \ci_a[61] , \ci_a[60] , \ci_a[59] , \ci_a[58] , 
        \ci_a[57] , \ci_a[56] , \ci_a[55] , \ci_a[54] , \ci_a[53] , \ci_a[52] , 
        \ci_a[51] , \ci_a[50] , \ci_a[49] , \ci_a[48] , \ci_a[47] , \ci_a[46] , 
        \ci_a[45] , \ci_a[44] , \ci_a[43] , \ci_a[42] , \ci_a[41] , \ci_a[40] , 
        \ci_a[39] , \ci_a[38] , \ci_a[37] , \ci_a[36] , \ci_a[35] , \ci_a[34] , 
        \ci_a[33] , \ci_a[32] , \ci_a[31] , \ci_a[30] , \ci_a[29] , \ci_a[28] , 
        \ci_a[27] , \ci_a[26] , \ci_a[25] , \ci_a[24] , \ci_a[23] , \ci_a[22] , 
        \ci_a[21] , \ci_a[20] , \ci_a[19] , \ci_a[18] , \ci_a[17] , \ci_a[16] , 
        \ci_a[15] , \ci_a[14] , \ci_a[13] , \ci_a[12] , \ci_a[11] , \ci_a[10] , 
        \ci_a[9] , \ci_a[8] , \ci_a[7] , \ci_a[6] , \ci_a[5] , \ci_a[4] , 
        \ci_a[3] , \ci_a[2] , \ci_a[1] , \ci_a[0] }), .chainresponse(
        chainresponse), .col({\ci_col[5] , \ci_col[4] , \ci_col[3] , 
        \ci_col[2] , \ci_col[1] , \ci_col[0] }), .crnw({\ci_rnw[1] , 
        \ci_rnw[0] }), .itag({\ci_itag[9] , \ci_itag[8] , \ci_itag[7] , 
        \ci_itag[6] , \ci_itag[5] , \ci_itag[4] , \ci_itag[3] , \ci_itag[2] , 
        \ci_itag[1] , \ci_itag[0] }), .lock({\ci_lock[1] , \ci_lock[0] }), 
        .nReset(nReset), .nchaincommandack(nchaincommandack), .pred({
        \ci_pred[1] , \ci_pred[0] }), .rack(ri_ack), .route({\route[4] , 1'b0, 
        1'b0, \route[1] , \route[0] }), .routetxack(routetx_ack), .seq({
        \ci_seq[1] , \ci_seq[0] }), .size({\ci_size[3] , \ci_size[2] , 
        \ci_size[1] , \ci_size[0] }), .wd({\ci_wd[63] , \ci_wd[62] , 
        \ci_wd[61] , \ci_wd[60] , \ci_wd[59] , \ci_wd[58] , \ci_wd[57] , 
        \ci_wd[56] , \ci_wd[55] , \ci_wd[54] , \ci_wd[53] , \ci_wd[52] , 
        \ci_wd[51] , \ci_wd[50] , \ci_wd[49] , \ci_wd[48] , \ci_wd[47] , 
        \ci_wd[46] , \ci_wd[45] , \ci_wd[44] , \ci_wd[43] , \ci_wd[42] , 
        \ci_wd[41] , \ci_wd[40] , \ci_wd[39] , \ci_wd[38] , \ci_wd[37] , 
        \ci_wd[36] , \ci_wd[35] , \ci_wd[34] , \ci_wd[33] , \ci_wd[32] , 
        \ci_wd[31] , \ci_wd[30] , \ci_wd[29] , \ci_wd[28] , \ci_wd[27] , 
        \ci_wd[26] , \ci_wd[25] , \ci_wd[24] , \ci_wd[23] , \ci_wd[22] , 
        \ci_wd[21] , \ci_wd[20] , \ci_wd[19] , \ci_wd[18] , \ci_wd[17] , 
        \ci_wd[16] , \ci_wd[15] , \ci_wd[14] , \ci_wd[13] , \ci_wd[12] , 
        \ci_wd[11] , \ci_wd[10] , \ci_wd[9] , \ci_wd[8] , \ci_wd[7] , 
        \ci_wd[6] , \ci_wd[5] , \ci_wd[4] , \ci_wd[3] , \ci_wd[2] , \ci_wd[1] , 
        \ci_wd[0] }) );
endmodule


module matched_delay_m2cp_com_tic ( x, a );
input  a;
output x;
    wire n2;
    buf_1 I1 ( .x(n2), .a(a) );
    buf_16 U1 ( .x(x), .a(n2) );
endmodule


module sr2dr_word_5 ( i, req, h, l );
input  [31:0] i;
output [31:0] h;
output [31:0] l;
input  req;
    wire \U31/ni , \U31/nh , \U31/nl , n9, n1, n2, \U30/ni , \U30/nh , 
        \U30/nl , n8, \U29/ni , \U29/nh , \U29/nl , \U28/ni , \U28/nh , 
        \U28/nl , \U27/ni , \U27/nh , \U27/nl , \U26/ni , \U26/nh , \U26/nl , 
        n7, n4, \U25/ni , \U25/nh , \U25/nl , \U24/ni , \U24/nh , \U24/nl , 
        \U23/ni , \U23/nh , \U23/nl , n3, \U22/ni , \U22/nh , \U22/nl , n6, 
        \U21/ni , \U21/nh , \U21/nl , \U20/ni , \U20/nh , \U20/nl , n5, 
        \U19/ni , \U19/nh , \U19/nl , \U18/ni , \U18/nh , \U18/nl , \U17/ni , 
        \U17/nh , \U17/nl , \U16/ni , \U16/nh , \U16/nl , \U15/ni , \U15/nh , 
        \U15/nl , \U14/ni , \U14/nh , \U14/nl , \U13/ni , \U13/nh , \U13/nl , 
        \U12/ni , \U12/nh , \U12/nl , \U11/ni , \U11/nh , \U11/nl , \U10/ni , 
        \U10/nh , \U10/nl , \U9/ni , \U9/nh , \U9/nl , \U8/ni , \U8/nh , 
        \U8/nl , \U7/ni , \U7/nh , \U7/nl , \U6/ni , \U6/nh , \U6/nl , \U5/ni , 
        \U5/nh , \U5/nl , \U4/ni , \U4/nh , \U4/nl , \U3/ni , \U3/nh , \U3/nl , 
        \U2/ni , \U2/nh , \U2/nl , \U1/ni , \U1/nh , \U1/nl , \U0/ni , \U0/nh , 
        \U0/nl , n12, n11, n10;
    inv_1 \U31/Uii  ( .x(\U31/ni ), .a(i[31]) );
    inv_1 \U31/Uih  ( .x(\U31/nh ), .a(h[31]) );
    inv_1 \U31/Uil  ( .x(\U31/nl ), .a(l[31]) );
    ao23_1 \U31/Ucl/U1/U1  ( .x(l[31]), .a(n9), .b(l[31]), .c(n1), .d(\U31/ni 
        ), .e(\U31/nh ) );
    ao23_1 \U31/Uch/U1/U1  ( .x(h[31]), .a(n9), .b(h[31]), .c(n2), .d(i[31]), 
        .e(\U31/nl ) );
    inv_1 \U30/Uii  ( .x(\U30/ni ), .a(i[30]) );
    inv_1 \U30/Uih  ( .x(\U30/nh ), .a(h[30]) );
    inv_1 \U30/Uil  ( .x(\U30/nl ), .a(l[30]) );
    ao23_1 \U30/Ucl/U1/U1  ( .x(l[30]), .a(n8), .b(l[30]), .c(n1), .d(\U30/ni 
        ), .e(\U30/nh ) );
    ao23_1 \U30/Uch/U1/U1  ( .x(h[30]), .a(n8), .b(h[30]), .c(n1), .d(i[30]), 
        .e(\U30/nl ) );
    inv_1 \U29/Uii  ( .x(\U29/ni ), .a(i[29]) );
    inv_1 \U29/Uih  ( .x(\U29/nh ), .a(h[29]) );
    inv_1 \U29/Uil  ( .x(\U29/nl ), .a(l[29]) );
    ao23_1 \U29/Ucl/U1/U1  ( .x(l[29]), .a(n8), .b(l[29]), .c(n1), .d(\U29/ni 
        ), .e(\U29/nh ) );
    ao23_1 \U29/Uch/U1/U1  ( .x(h[29]), .a(n8), .b(h[29]), .c(n2), .d(i[29]), 
        .e(\U29/nl ) );
    inv_1 \U28/Uii  ( .x(\U28/ni ), .a(i[28]) );
    inv_1 \U28/Uih  ( .x(\U28/nh ), .a(h[28]) );
    inv_1 \U28/Uil  ( .x(\U28/nl ), .a(l[28]) );
    ao23_1 \U28/Ucl/U1/U1  ( .x(l[28]), .a(n8), .b(l[28]), .c(n2), .d(\U28/ni 
        ), .e(\U28/nh ) );
    ao23_1 \U28/Uch/U1/U1  ( .x(h[28]), .a(n8), .b(h[28]), .c(n2), .d(i[28]), 
        .e(\U28/nl ) );
    inv_1 \U27/Uii  ( .x(\U27/ni ), .a(i[27]) );
    inv_1 \U27/Uih  ( .x(\U27/nh ), .a(h[27]) );
    inv_1 \U27/Uil  ( .x(\U27/nl ), .a(l[27]) );
    ao23_1 \U27/Ucl/U1/U1  ( .x(l[27]), .a(n8), .b(l[27]), .c(n2), .d(\U27/ni 
        ), .e(\U27/nh ) );
    ao23_1 \U27/Uch/U1/U1  ( .x(h[27]), .a(n8), .b(h[27]), .c(n2), .d(i[27]), 
        .e(\U27/nl ) );
    inv_1 \U26/Uii  ( .x(\U26/ni ), .a(i[26]) );
    inv_1 \U26/Uih  ( .x(\U26/nh ), .a(h[26]) );
    inv_1 \U26/Uil  ( .x(\U26/nl ), .a(l[26]) );
    ao23_1 \U26/Ucl/U1/U1  ( .x(l[26]), .a(n7), .b(l[26]), .c(n2), .d(\U26/ni 
        ), .e(\U26/nh ) );
    ao23_1 \U26/Uch/U1/U1  ( .x(h[26]), .a(n7), .b(h[26]), .c(n4), .d(i[26]), 
        .e(\U26/nl ) );
    inv_1 \U25/Uii  ( .x(\U25/ni ), .a(i[25]) );
    inv_1 \U25/Uih  ( .x(\U25/nh ), .a(h[25]) );
    inv_1 \U25/Uil  ( .x(\U25/nl ), .a(l[25]) );
    ao23_1 \U25/Ucl/U1/U1  ( .x(l[25]), .a(n7), .b(l[25]), .c(n4), .d(\U25/ni 
        ), .e(\U25/nh ) );
    ao23_1 \U25/Uch/U1/U1  ( .x(h[25]), .a(n7), .b(h[25]), .c(n4), .d(i[25]), 
        .e(\U25/nl ) );
    inv_1 \U24/Uii  ( .x(\U24/ni ), .a(i[24]) );
    inv_1 \U24/Uih  ( .x(\U24/nh ), .a(h[24]) );
    inv_1 \U24/Uil  ( .x(\U24/nl ), .a(l[24]) );
    ao23_1 \U24/Ucl/U1/U1  ( .x(l[24]), .a(n7), .b(l[24]), .c(n4), .d(\U24/ni 
        ), .e(\U24/nh ) );
    ao23_1 \U24/Uch/U1/U1  ( .x(h[24]), .a(n7), .b(h[24]), .c(n4), .d(i[24]), 
        .e(\U24/nl ) );
    inv_1 \U23/Uii  ( .x(\U23/ni ), .a(i[23]) );
    inv_1 \U23/Uih  ( .x(\U23/nh ), .a(h[23]) );
    inv_1 \U23/Uil  ( .x(\U23/nl ), .a(l[23]) );
    ao23_1 \U23/Ucl/U1/U1  ( .x(l[23]), .a(n7), .b(l[23]), .c(n3), .d(\U23/ni 
        ), .e(\U23/nh ) );
    ao23_1 \U23/Uch/U1/U1  ( .x(h[23]), .a(n7), .b(h[23]), .c(n3), .d(i[23]), 
        .e(\U23/nl ) );
    inv_1 \U22/Uii  ( .x(\U22/ni ), .a(i[22]) );
    inv_1 \U22/Uih  ( .x(\U22/nh ), .a(h[22]) );
    inv_1 \U22/Uil  ( .x(\U22/nl ), .a(l[22]) );
    ao23_1 \U22/Ucl/U1/U1  ( .x(l[22]), .a(n6), .b(l[22]), .c(n3), .d(\U22/ni 
        ), .e(\U22/nh ) );
    ao23_1 \U22/Uch/U1/U1  ( .x(h[22]), .a(n6), .b(h[22]), .c(n3), .d(i[22]), 
        .e(\U22/nl ) );
    inv_1 \U21/Uii  ( .x(\U21/ni ), .a(i[21]) );
    inv_1 \U21/Uih  ( .x(\U21/nh ), .a(h[21]) );
    inv_1 \U21/Uil  ( .x(\U21/nl ), .a(l[21]) );
    ao23_1 \U21/Ucl/U1/U1  ( .x(l[21]), .a(n6), .b(l[21]), .c(n3), .d(\U21/ni 
        ), .e(\U21/nh ) );
    ao23_1 \U21/Uch/U1/U1  ( .x(h[21]), .a(n6), .b(h[21]), .c(n3), .d(i[21]), 
        .e(\U21/nl ) );
    inv_1 \U20/Uii  ( .x(\U20/ni ), .a(i[20]) );
    inv_1 \U20/Uih  ( .x(\U20/nh ), .a(h[20]) );
    inv_1 \U20/Uil  ( .x(\U20/nl ), .a(l[20]) );
    ao23_1 \U20/Ucl/U1/U1  ( .x(l[20]), .a(n6), .b(l[20]), .c(n5), .d(\U20/ni 
        ), .e(\U20/nh ) );
    ao23_1 \U20/Uch/U1/U1  ( .x(h[20]), .a(n6), .b(h[20]), .c(n4), .d(i[20]), 
        .e(\U20/nl ) );
    inv_1 \U19/Uii  ( .x(\U19/ni ), .a(i[19]) );
    inv_1 \U19/Uih  ( .x(\U19/nh ), .a(h[19]) );
    inv_1 \U19/Uil  ( .x(\U19/nl ), .a(l[19]) );
    ao23_1 \U19/Ucl/U1/U1  ( .x(l[19]), .a(n6), .b(l[19]), .c(n4), .d(\U19/ni 
        ), .e(\U19/nh ) );
    ao23_1 \U19/Uch/U1/U1  ( .x(h[19]), .a(n6), .b(h[19]), .c(n4), .d(i[19]), 
        .e(\U19/nl ) );
    inv_1 \U18/Uii  ( .x(\U18/ni ), .a(i[18]) );
    inv_1 \U18/Uih  ( .x(\U18/nh ), .a(h[18]) );
    inv_1 \U18/Uil  ( .x(\U18/nl ), .a(l[18]) );
    ao23_1 \U18/Ucl/U1/U1  ( .x(l[18]), .a(n5), .b(l[18]), .c(n5), .d(\U18/ni 
        ), .e(\U18/nh ) );
    ao23_1 \U18/Uch/U1/U1  ( .x(h[18]), .a(n5), .b(h[18]), .c(n5), .d(i[18]), 
        .e(\U18/nl ) );
    inv_1 \U17/Uii  ( .x(\U17/ni ), .a(i[17]) );
    inv_1 \U17/Uih  ( .x(\U17/nh ), .a(h[17]) );
    inv_1 \U17/Uil  ( .x(\U17/nl ), .a(l[17]) );
    ao23_1 \U17/Ucl/U1/U1  ( .x(l[17]), .a(n6), .b(l[17]), .c(n5), .d(\U17/ni 
        ), .e(\U17/nh ) );
    ao23_1 \U17/Uch/U1/U1  ( .x(h[17]), .a(n7), .b(h[17]), .c(n4), .d(i[17]), 
        .e(\U17/nl ) );
    inv_1 \U16/Uii  ( .x(\U16/ni ), .a(i[16]) );
    inv_1 \U16/Uih  ( .x(\U16/nh ), .a(h[16]) );
    inv_1 \U16/Uil  ( .x(\U16/nl ), .a(l[16]) );
    ao23_1 \U16/Ucl/U1/U1  ( .x(l[16]), .a(n9), .b(l[16]), .c(n3), .d(\U16/ni 
        ), .e(\U16/nh ) );
    ao23_1 \U16/Uch/U1/U1  ( .x(h[16]), .a(n9), .b(h[16]), .c(n1), .d(i[16]), 
        .e(\U16/nl ) );
    inv_1 \U15/Uii  ( .x(\U15/ni ), .a(i[15]) );
    inv_1 \U15/Uih  ( .x(\U15/nh ), .a(h[15]) );
    inv_1 \U15/Uil  ( .x(\U15/nl ), .a(l[15]) );
    ao23_1 \U15/Ucl/U1/U1  ( .x(l[15]), .a(n8), .b(l[15]), .c(n1), .d(\U15/ni 
        ), .e(\U15/nh ) );
    ao23_1 \U15/Uch/U1/U1  ( .x(h[15]), .a(n7), .b(h[15]), .c(n1), .d(i[15]), 
        .e(\U15/nl ) );
    inv_1 \U14/Uii  ( .x(\U14/ni ), .a(i[14]) );
    inv_1 \U14/Uih  ( .x(\U14/nh ), .a(h[14]) );
    inv_1 \U14/Uil  ( .x(\U14/nl ), .a(l[14]) );
    ao23_1 \U14/Ucl/U1/U1  ( .x(l[14]), .a(n6), .b(l[14]), .c(n1), .d(\U14/ni 
        ), .e(\U14/nh ) );
    ao23_1 \U14/Uch/U1/U1  ( .x(h[14]), .a(n6), .b(h[14]), .c(n3), .d(i[14]), 
        .e(\U14/nl ) );
    inv_1 \U13/Uii  ( .x(\U13/ni ), .a(i[13]) );
    inv_1 \U13/Uih  ( .x(\U13/nh ), .a(h[13]) );
    inv_1 \U13/Uil  ( .x(\U13/nl ), .a(l[13]) );
    ao23_1 \U13/Ucl/U1/U1  ( .x(l[13]), .a(n6), .b(l[13]), .c(n4), .d(\U13/ni 
        ), .e(\U13/nh ) );
    ao23_1 \U13/Uch/U1/U1  ( .x(h[13]), .a(n6), .b(h[13]), .c(n4), .d(i[13]), 
        .e(\U13/nl ) );
    inv_1 \U12/Uii  ( .x(\U12/ni ), .a(i[12]) );
    inv_1 \U12/Uih  ( .x(\U12/nh ), .a(h[12]) );
    inv_1 \U12/Uil  ( .x(\U12/nl ), .a(l[12]) );
    ao23_1 \U12/Ucl/U1/U1  ( .x(l[12]), .a(n5), .b(l[12]), .c(n4), .d(\U12/ni 
        ), .e(\U12/nh ) );
    ao23_1 \U12/Uch/U1/U1  ( .x(h[12]), .a(n5), .b(h[12]), .c(n4), .d(i[12]), 
        .e(\U12/nl ) );
    inv_1 \U11/Uii  ( .x(\U11/ni ), .a(i[11]) );
    inv_1 \U11/Uih  ( .x(\U11/nh ), .a(h[11]) );
    inv_1 \U11/Uil  ( .x(\U11/nl ), .a(l[11]) );
    ao23_1 \U11/Ucl/U1/U1  ( .x(l[11]), .a(n5), .b(l[11]), .c(n4), .d(\U11/ni 
        ), .e(\U11/nh ) );
    ao23_1 \U11/Uch/U1/U1  ( .x(h[11]), .a(n5), .b(h[11]), .c(n4), .d(i[11]), 
        .e(\U11/nl ) );
    inv_1 \U10/Uii  ( .x(\U10/ni ), .a(i[10]) );
    inv_1 \U10/Uih  ( .x(\U10/nh ), .a(h[10]) );
    inv_1 \U10/Uil  ( .x(\U10/nl ), .a(l[10]) );
    ao23_1 \U10/Ucl/U1/U1  ( .x(l[10]), .a(n5), .b(l[10]), .c(n3), .d(\U10/ni 
        ), .e(\U10/nh ) );
    ao23_1 \U10/Uch/U1/U1  ( .x(h[10]), .a(n5), .b(h[10]), .c(n3), .d(i[10]), 
        .e(\U10/nl ) );
    inv_1 \U9/Uii  ( .x(\U9/ni ), .a(i[9]) );
    inv_1 \U9/Uih  ( .x(\U9/nh ), .a(h[9]) );
    inv_1 \U9/Uil  ( .x(\U9/nl ), .a(l[9]) );
    ao23_1 \U9/Ucl/U1/U1  ( .x(l[9]), .a(n5), .b(l[9]), .c(n3), .d(\U9/ni ), 
        .e(\U9/nh ) );
    ao23_1 \U9/Uch/U1/U1  ( .x(h[9]), .a(n5), .b(h[9]), .c(n3), .d(i[9]), .e(
        \U9/nl ) );
    inv_1 \U8/Uii  ( .x(\U8/ni ), .a(i[8]) );
    inv_1 \U8/Uih  ( .x(\U8/nh ), .a(h[8]) );
    inv_1 \U8/Uil  ( .x(\U8/nl ), .a(l[8]) );
    ao23_1 \U8/Ucl/U1/U1  ( .x(l[8]), .a(n5), .b(l[8]), .c(n3), .d(\U8/ni ), 
        .e(\U8/nh ) );
    ao23_1 \U8/Uch/U1/U1  ( .x(h[8]), .a(n5), .b(h[8]), .c(n3), .d(i[8]), .e(
        \U8/nl ) );
    inv_1 \U7/Uii  ( .x(\U7/ni ), .a(i[7]) );
    inv_1 \U7/Uih  ( .x(\U7/nh ), .a(h[7]) );
    inv_1 \U7/Uil  ( .x(\U7/nl ), .a(l[7]) );
    ao23_1 \U7/Ucl/U1/U1  ( .x(l[7]), .a(n7), .b(l[7]), .c(n3), .d(\U7/ni ), 
        .e(\U7/nh ) );
    ao23_1 \U7/Uch/U1/U1  ( .x(h[7]), .a(n7), .b(h[7]), .c(n2), .d(i[7]), .e(
        \U7/nl ) );
    inv_1 \U6/Uii  ( .x(\U6/ni ), .a(i[6]) );
    inv_1 \U6/Uih  ( .x(\U6/nh ), .a(h[6]) );
    inv_1 \U6/Uil  ( .x(\U6/nl ), .a(l[6]) );
    ao23_1 \U6/Ucl/U1/U1  ( .x(l[6]), .a(n7), .b(l[6]), .c(n2), .d(\U6/ni ), 
        .e(\U6/nh ) );
    ao23_1 \U6/Uch/U1/U1  ( .x(h[6]), .a(n7), .b(h[6]), .c(n2), .d(i[6]), .e(
        \U6/nl ) );
    inv_1 \U5/Uii  ( .x(\U5/ni ), .a(i[5]) );
    inv_1 \U5/Uih  ( .x(\U5/nh ), .a(h[5]) );
    inv_1 \U5/Uil  ( .x(\U5/nl ), .a(l[5]) );
    ao23_1 \U5/Ucl/U1/U1  ( .x(l[5]), .a(n7), .b(l[5]), .c(n2), .d(\U5/ni ), 
        .e(\U5/nh ) );
    ao23_1 \U5/Uch/U1/U1  ( .x(h[5]), .a(n7), .b(h[5]), .c(n2), .d(i[5]), .e(
        \U5/nl ) );
    inv_1 \U4/Uii  ( .x(\U4/ni ), .a(i[4]) );
    inv_1 \U4/Uih  ( .x(\U4/nh ), .a(h[4]) );
    inv_1 \U4/Uil  ( .x(\U4/nl ), .a(l[4]) );
    ao23_1 \U4/Ucl/U1/U1  ( .x(l[4]), .a(n6), .b(l[4]), .c(n2), .d(\U4/ni ), 
        .e(\U4/nh ) );
    ao23_1 \U4/Uch/U1/U1  ( .x(h[4]), .a(n6), .b(h[4]), .c(n2), .d(i[4]), .e(
        \U4/nl ) );
    inv_1 \U3/Uii  ( .x(\U3/ni ), .a(i[3]) );
    inv_1 \U3/Uih  ( .x(\U3/nh ), .a(h[3]) );
    inv_1 \U3/Uil  ( .x(\U3/nl ), .a(l[3]) );
    ao23_1 \U3/Ucl/U1/U1  ( .x(l[3]), .a(n6), .b(l[3]), .c(n2), .d(\U3/ni ), 
        .e(\U3/nh ) );
    ao23_1 \U3/Uch/U1/U1  ( .x(h[3]), .a(n8), .b(h[3]), .c(n1), .d(i[3]), .e(
        \U3/nl ) );
    inv_1 \U2/Uii  ( .x(\U2/ni ), .a(i[2]) );
    inv_1 \U2/Uih  ( .x(\U2/nh ), .a(h[2]) );
    inv_1 \U2/Uil  ( .x(\U2/nl ), .a(l[2]) );
    ao23_1 \U2/Ucl/U1/U1  ( .x(l[2]), .a(n8), .b(l[2]), .c(n1), .d(\U2/ni ), 
        .e(\U2/nh ) );
    ao23_1 \U2/Uch/U1/U1  ( .x(h[2]), .a(n8), .b(h[2]), .c(n1), .d(i[2]), .e(
        \U2/nl ) );
    inv_1 \U1/Uii  ( .x(\U1/ni ), .a(i[1]) );
    inv_1 \U1/Uih  ( .x(\U1/nh ), .a(h[1]) );
    inv_1 \U1/Uil  ( .x(\U1/nl ), .a(l[1]) );
    ao23_1 \U1/Ucl/U1/U1  ( .x(l[1]), .a(n8), .b(l[1]), .c(n1), .d(\U1/ni ), 
        .e(\U1/nh ) );
    ao23_1 \U1/Uch/U1/U1  ( .x(h[1]), .a(n8), .b(h[1]), .c(n1), .d(i[1]), .e(
        \U1/nl ) );
    inv_1 \U0/Uii  ( .x(\U0/ni ), .a(i[0]) );
    inv_1 \U0/Uih  ( .x(\U0/nh ), .a(h[0]) );
    inv_1 \U0/Uil  ( .x(\U0/nl ), .a(l[0]) );
    ao23_1 \U0/Ucl/U1/U1  ( .x(l[0]), .a(n8), .b(l[0]), .c(n1), .d(\U0/ni ), 
        .e(\U0/nh ) );
    ao23_1 \U0/Uch/U1/U1  ( .x(h[0]), .a(n8), .b(h[0]), .c(n1), .d(i[0]), .e(
        \U0/nl ) );
    buf_16 U1 ( .x(n1), .a(n12) );
    buf_16 U2 ( .x(n2), .a(n12) );
    buf_16 U3 ( .x(n3), .a(n12) );
    buf_16 U4 ( .x(n4), .a(n11) );
    buf_16 U5 ( .x(n5), .a(n11) );
    buf_16 U6 ( .x(n6), .a(n11) );
    buf_16 U7 ( .x(n7), .a(n10) );
    buf_16 U8 ( .x(n8), .a(n10) );
    buf_16 U9 ( .x(n9), .a(n10) );
    buf_16 U10 ( .x(n10), .a(req) );
    buf_16 U11 ( .x(n11), .a(req) );
    buf_16 U12 ( .x(n12), .a(req) );
endmodule


module sr2dr_word_4 ( i, req, h, l );
input  [31:0] i;
output [31:0] h;
output [31:0] l;
input  req;
    wire \U31/ni , \U31/nh , \U31/nl , n9, n1, n2, \U30/ni , \U30/nh , 
        \U30/nl , n8, \U29/ni , \U29/nh , \U29/nl , \U28/ni , \U28/nh , 
        \U28/nl , \U27/ni , \U27/nh , \U27/nl , \U26/ni , \U26/nh , \U26/nl , 
        n7, n4, \U25/ni , \U25/nh , \U25/nl , \U24/ni , \U24/nh , \U24/nl , 
        \U23/ni , \U23/nh , \U23/nl , n3, \U22/ni , \U22/nh , \U22/nl , n6, 
        \U21/ni , \U21/nh , \U21/nl , \U20/ni , \U20/nh , \U20/nl , n5, 
        \U19/ni , \U19/nh , \U19/nl , \U18/ni , \U18/nh , \U18/nl , \U17/ni , 
        \U17/nh , \U17/nl , \U16/ni , \U16/nh , \U16/nl , \U15/ni , \U15/nh , 
        \U15/nl , \U14/ni , \U14/nh , \U14/nl , \U13/ni , \U13/nh , \U13/nl , 
        \U12/ni , \U12/nh , \U12/nl , \U11/ni , \U11/nh , \U11/nl , \U10/ni , 
        \U10/nh , \U10/nl , \U9/ni , \U9/nh , \U9/nl , \U8/ni , \U8/nh , 
        \U8/nl , \U7/ni , \U7/nh , \U7/nl , \U6/ni , \U6/nh , \U6/nl , \U5/ni , 
        \U5/nh , \U5/nl , \U4/ni , \U4/nh , \U4/nl , \U3/ni , \U3/nh , \U3/nl , 
        \U2/ni , \U2/nh , \U2/nl , \U1/ni , \U1/nh , \U1/nl , \U0/ni , \U0/nh , 
        \U0/nl , n12, n11, n10;
    inv_1 \U31/Uii  ( .x(\U31/ni ), .a(i[31]) );
    inv_1 \U31/Uih  ( .x(\U31/nh ), .a(h[31]) );
    inv_1 \U31/Uil  ( .x(\U31/nl ), .a(l[31]) );
    ao23_1 \U31/Ucl/U1/U1  ( .x(l[31]), .a(n9), .b(l[31]), .c(n1), .d(\U31/ni 
        ), .e(\U31/nh ) );
    ao23_1 \U31/Uch/U1/U1  ( .x(h[31]), .a(n9), .b(h[31]), .c(n2), .d(i[31]), 
        .e(\U31/nl ) );
    inv_1 \U30/Uii  ( .x(\U30/ni ), .a(i[30]) );
    inv_1 \U30/Uih  ( .x(\U30/nh ), .a(h[30]) );
    inv_1 \U30/Uil  ( .x(\U30/nl ), .a(l[30]) );
    ao23_1 \U30/Ucl/U1/U1  ( .x(l[30]), .a(n8), .b(l[30]), .c(n1), .d(\U30/ni 
        ), .e(\U30/nh ) );
    ao23_1 \U30/Uch/U1/U1  ( .x(h[30]), .a(n8), .b(h[30]), .c(n1), .d(i[30]), 
        .e(\U30/nl ) );
    inv_1 \U29/Uii  ( .x(\U29/ni ), .a(i[29]) );
    inv_1 \U29/Uih  ( .x(\U29/nh ), .a(h[29]) );
    inv_1 \U29/Uil  ( .x(\U29/nl ), .a(l[29]) );
    ao23_1 \U29/Ucl/U1/U1  ( .x(l[29]), .a(n8), .b(l[29]), .c(n1), .d(\U29/ni 
        ), .e(\U29/nh ) );
    ao23_1 \U29/Uch/U1/U1  ( .x(h[29]), .a(n8), .b(h[29]), .c(n2), .d(i[29]), 
        .e(\U29/nl ) );
    inv_1 \U28/Uii  ( .x(\U28/ni ), .a(i[28]) );
    inv_1 \U28/Uih  ( .x(\U28/nh ), .a(h[28]) );
    inv_1 \U28/Uil  ( .x(\U28/nl ), .a(l[28]) );
    ao23_1 \U28/Ucl/U1/U1  ( .x(l[28]), .a(n8), .b(l[28]), .c(n2), .d(\U28/ni 
        ), .e(\U28/nh ) );
    ao23_1 \U28/Uch/U1/U1  ( .x(h[28]), .a(n8), .b(h[28]), .c(n2), .d(i[28]), 
        .e(\U28/nl ) );
    inv_1 \U27/Uii  ( .x(\U27/ni ), .a(i[27]) );
    inv_1 \U27/Uih  ( .x(\U27/nh ), .a(h[27]) );
    inv_1 \U27/Uil  ( .x(\U27/nl ), .a(l[27]) );
    ao23_1 \U27/Ucl/U1/U1  ( .x(l[27]), .a(n8), .b(l[27]), .c(n2), .d(\U27/ni 
        ), .e(\U27/nh ) );
    ao23_1 \U27/Uch/U1/U1  ( .x(h[27]), .a(n8), .b(h[27]), .c(n2), .d(i[27]), 
        .e(\U27/nl ) );
    inv_1 \U26/Uii  ( .x(\U26/ni ), .a(i[26]) );
    inv_1 \U26/Uih  ( .x(\U26/nh ), .a(h[26]) );
    inv_1 \U26/Uil  ( .x(\U26/nl ), .a(l[26]) );
    ao23_1 \U26/Ucl/U1/U1  ( .x(l[26]), .a(n7), .b(l[26]), .c(n2), .d(\U26/ni 
        ), .e(\U26/nh ) );
    ao23_1 \U26/Uch/U1/U1  ( .x(h[26]), .a(n7), .b(h[26]), .c(n4), .d(i[26]), 
        .e(\U26/nl ) );
    inv_1 \U25/Uii  ( .x(\U25/ni ), .a(i[25]) );
    inv_1 \U25/Uih  ( .x(\U25/nh ), .a(h[25]) );
    inv_1 \U25/Uil  ( .x(\U25/nl ), .a(l[25]) );
    ao23_1 \U25/Ucl/U1/U1  ( .x(l[25]), .a(n7), .b(l[25]), .c(n4), .d(\U25/ni 
        ), .e(\U25/nh ) );
    ao23_1 \U25/Uch/U1/U1  ( .x(h[25]), .a(n7), .b(h[25]), .c(n4), .d(i[25]), 
        .e(\U25/nl ) );
    inv_1 \U24/Uii  ( .x(\U24/ni ), .a(i[24]) );
    inv_1 \U24/Uih  ( .x(\U24/nh ), .a(h[24]) );
    inv_1 \U24/Uil  ( .x(\U24/nl ), .a(l[24]) );
    ao23_1 \U24/Ucl/U1/U1  ( .x(l[24]), .a(n7), .b(l[24]), .c(n4), .d(\U24/ni 
        ), .e(\U24/nh ) );
    ao23_1 \U24/Uch/U1/U1  ( .x(h[24]), .a(n7), .b(h[24]), .c(n4), .d(i[24]), 
        .e(\U24/nl ) );
    inv_1 \U23/Uii  ( .x(\U23/ni ), .a(i[23]) );
    inv_1 \U23/Uih  ( .x(\U23/nh ), .a(h[23]) );
    inv_1 \U23/Uil  ( .x(\U23/nl ), .a(l[23]) );
    ao23_1 \U23/Ucl/U1/U1  ( .x(l[23]), .a(n7), .b(l[23]), .c(n3), .d(\U23/ni 
        ), .e(\U23/nh ) );
    ao23_1 \U23/Uch/U1/U1  ( .x(h[23]), .a(n7), .b(h[23]), .c(n3), .d(i[23]), 
        .e(\U23/nl ) );
    inv_1 \U22/Uii  ( .x(\U22/ni ), .a(i[22]) );
    inv_1 \U22/Uih  ( .x(\U22/nh ), .a(h[22]) );
    inv_1 \U22/Uil  ( .x(\U22/nl ), .a(l[22]) );
    ao23_1 \U22/Ucl/U1/U1  ( .x(l[22]), .a(n6), .b(l[22]), .c(n3), .d(\U22/ni 
        ), .e(\U22/nh ) );
    ao23_1 \U22/Uch/U1/U1  ( .x(h[22]), .a(n6), .b(h[22]), .c(n3), .d(i[22]), 
        .e(\U22/nl ) );
    inv_1 \U21/Uii  ( .x(\U21/ni ), .a(i[21]) );
    inv_1 \U21/Uih  ( .x(\U21/nh ), .a(h[21]) );
    inv_1 \U21/Uil  ( .x(\U21/nl ), .a(l[21]) );
    ao23_1 \U21/Ucl/U1/U1  ( .x(l[21]), .a(n6), .b(l[21]), .c(n3), .d(\U21/ni 
        ), .e(\U21/nh ) );
    ao23_1 \U21/Uch/U1/U1  ( .x(h[21]), .a(n6), .b(h[21]), .c(n3), .d(i[21]), 
        .e(\U21/nl ) );
    inv_1 \U20/Uii  ( .x(\U20/ni ), .a(i[20]) );
    inv_1 \U20/Uih  ( .x(\U20/nh ), .a(h[20]) );
    inv_1 \U20/Uil  ( .x(\U20/nl ), .a(l[20]) );
    ao23_1 \U20/Ucl/U1/U1  ( .x(l[20]), .a(n6), .b(l[20]), .c(n5), .d(\U20/ni 
        ), .e(\U20/nh ) );
    ao23_1 \U20/Uch/U1/U1  ( .x(h[20]), .a(n6), .b(h[20]), .c(n4), .d(i[20]), 
        .e(\U20/nl ) );
    inv_1 \U19/Uii  ( .x(\U19/ni ), .a(i[19]) );
    inv_1 \U19/Uih  ( .x(\U19/nh ), .a(h[19]) );
    inv_1 \U19/Uil  ( .x(\U19/nl ), .a(l[19]) );
    ao23_1 \U19/Ucl/U1/U1  ( .x(l[19]), .a(n6), .b(l[19]), .c(n4), .d(\U19/ni 
        ), .e(\U19/nh ) );
    ao23_1 \U19/Uch/U1/U1  ( .x(h[19]), .a(n6), .b(h[19]), .c(n4), .d(i[19]), 
        .e(\U19/nl ) );
    inv_1 \U18/Uii  ( .x(\U18/ni ), .a(i[18]) );
    inv_1 \U18/Uih  ( .x(\U18/nh ), .a(h[18]) );
    inv_1 \U18/Uil  ( .x(\U18/nl ), .a(l[18]) );
    ao23_1 \U18/Ucl/U1/U1  ( .x(l[18]), .a(n5), .b(l[18]), .c(n5), .d(\U18/ni 
        ), .e(\U18/nh ) );
    ao23_1 \U18/Uch/U1/U1  ( .x(h[18]), .a(n5), .b(h[18]), .c(n5), .d(i[18]), 
        .e(\U18/nl ) );
    inv_1 \U17/Uii  ( .x(\U17/ni ), .a(i[17]) );
    inv_1 \U17/Uih  ( .x(\U17/nh ), .a(h[17]) );
    inv_1 \U17/Uil  ( .x(\U17/nl ), .a(l[17]) );
    ao23_1 \U17/Ucl/U1/U1  ( .x(l[17]), .a(n6), .b(l[17]), .c(n5), .d(\U17/ni 
        ), .e(\U17/nh ) );
    ao23_1 \U17/Uch/U1/U1  ( .x(h[17]), .a(n7), .b(h[17]), .c(n4), .d(i[17]), 
        .e(\U17/nl ) );
    inv_1 \U16/Uii  ( .x(\U16/ni ), .a(i[16]) );
    inv_1 \U16/Uih  ( .x(\U16/nh ), .a(h[16]) );
    inv_1 \U16/Uil  ( .x(\U16/nl ), .a(l[16]) );
    ao23_1 \U16/Ucl/U1/U1  ( .x(l[16]), .a(n9), .b(l[16]), .c(n3), .d(\U16/ni 
        ), .e(\U16/nh ) );
    ao23_1 \U16/Uch/U1/U1  ( .x(h[16]), .a(n9), .b(h[16]), .c(n1), .d(i[16]), 
        .e(\U16/nl ) );
    inv_1 \U15/Uii  ( .x(\U15/ni ), .a(i[15]) );
    inv_1 \U15/Uih  ( .x(\U15/nh ), .a(h[15]) );
    inv_1 \U15/Uil  ( .x(\U15/nl ), .a(l[15]) );
    ao23_1 \U15/Ucl/U1/U1  ( .x(l[15]), .a(n8), .b(l[15]), .c(n1), .d(\U15/ni 
        ), .e(\U15/nh ) );
    ao23_1 \U15/Uch/U1/U1  ( .x(h[15]), .a(n7), .b(h[15]), .c(n1), .d(i[15]), 
        .e(\U15/nl ) );
    inv_1 \U14/Uii  ( .x(\U14/ni ), .a(i[14]) );
    inv_1 \U14/Uih  ( .x(\U14/nh ), .a(h[14]) );
    inv_1 \U14/Uil  ( .x(\U14/nl ), .a(l[14]) );
    ao23_1 \U14/Ucl/U1/U1  ( .x(l[14]), .a(n6), .b(l[14]), .c(n1), .d(\U14/ni 
        ), .e(\U14/nh ) );
    ao23_1 \U14/Uch/U1/U1  ( .x(h[14]), .a(n6), .b(h[14]), .c(n3), .d(i[14]), 
        .e(\U14/nl ) );
    inv_1 \U13/Uii  ( .x(\U13/ni ), .a(i[13]) );
    inv_1 \U13/Uih  ( .x(\U13/nh ), .a(h[13]) );
    inv_1 \U13/Uil  ( .x(\U13/nl ), .a(l[13]) );
    ao23_1 \U13/Ucl/U1/U1  ( .x(l[13]), .a(n6), .b(l[13]), .c(n4), .d(\U13/ni 
        ), .e(\U13/nh ) );
    ao23_1 \U13/Uch/U1/U1  ( .x(h[13]), .a(n6), .b(h[13]), .c(n4), .d(i[13]), 
        .e(\U13/nl ) );
    inv_1 \U12/Uii  ( .x(\U12/ni ), .a(i[12]) );
    inv_1 \U12/Uih  ( .x(\U12/nh ), .a(h[12]) );
    inv_1 \U12/Uil  ( .x(\U12/nl ), .a(l[12]) );
    ao23_1 \U12/Ucl/U1/U1  ( .x(l[12]), .a(n5), .b(l[12]), .c(n4), .d(\U12/ni 
        ), .e(\U12/nh ) );
    ao23_1 \U12/Uch/U1/U1  ( .x(h[12]), .a(n5), .b(h[12]), .c(n4), .d(i[12]), 
        .e(\U12/nl ) );
    inv_1 \U11/Uii  ( .x(\U11/ni ), .a(i[11]) );
    inv_1 \U11/Uih  ( .x(\U11/nh ), .a(h[11]) );
    inv_1 \U11/Uil  ( .x(\U11/nl ), .a(l[11]) );
    ao23_1 \U11/Ucl/U1/U1  ( .x(l[11]), .a(n5), .b(l[11]), .c(n4), .d(\U11/ni 
        ), .e(\U11/nh ) );
    ao23_1 \U11/Uch/U1/U1  ( .x(h[11]), .a(n5), .b(h[11]), .c(n4), .d(i[11]), 
        .e(\U11/nl ) );
    inv_1 \U10/Uii  ( .x(\U10/ni ), .a(i[10]) );
    inv_1 \U10/Uih  ( .x(\U10/nh ), .a(h[10]) );
    inv_1 \U10/Uil  ( .x(\U10/nl ), .a(l[10]) );
    ao23_1 \U10/Ucl/U1/U1  ( .x(l[10]), .a(n5), .b(l[10]), .c(n3), .d(\U10/ni 
        ), .e(\U10/nh ) );
    ao23_1 \U10/Uch/U1/U1  ( .x(h[10]), .a(n5), .b(h[10]), .c(n3), .d(i[10]), 
        .e(\U10/nl ) );
    inv_1 \U9/Uii  ( .x(\U9/ni ), .a(i[9]) );
    inv_1 \U9/Uih  ( .x(\U9/nh ), .a(h[9]) );
    inv_1 \U9/Uil  ( .x(\U9/nl ), .a(l[9]) );
    ao23_1 \U9/Ucl/U1/U1  ( .x(l[9]), .a(n5), .b(l[9]), .c(n3), .d(\U9/ni ), 
        .e(\U9/nh ) );
    ao23_1 \U9/Uch/U1/U1  ( .x(h[9]), .a(n5), .b(h[9]), .c(n3), .d(i[9]), .e(
        \U9/nl ) );
    inv_1 \U8/Uii  ( .x(\U8/ni ), .a(i[8]) );
    inv_1 \U8/Uih  ( .x(\U8/nh ), .a(h[8]) );
    inv_1 \U8/Uil  ( .x(\U8/nl ), .a(l[8]) );
    ao23_1 \U8/Ucl/U1/U1  ( .x(l[8]), .a(n5), .b(l[8]), .c(n3), .d(\U8/ni ), 
        .e(\U8/nh ) );
    ao23_1 \U8/Uch/U1/U1  ( .x(h[8]), .a(n5), .b(h[8]), .c(n3), .d(i[8]), .e(
        \U8/nl ) );
    inv_1 \U7/Uii  ( .x(\U7/ni ), .a(i[7]) );
    inv_1 \U7/Uih  ( .x(\U7/nh ), .a(h[7]) );
    inv_1 \U7/Uil  ( .x(\U7/nl ), .a(l[7]) );
    ao23_1 \U7/Ucl/U1/U1  ( .x(l[7]), .a(n7), .b(l[7]), .c(n3), .d(\U7/ni ), 
        .e(\U7/nh ) );
    ao23_1 \U7/Uch/U1/U1  ( .x(h[7]), .a(n7), .b(h[7]), .c(n2), .d(i[7]), .e(
        \U7/nl ) );
    inv_1 \U6/Uii  ( .x(\U6/ni ), .a(i[6]) );
    inv_1 \U6/Uih  ( .x(\U6/nh ), .a(h[6]) );
    inv_1 \U6/Uil  ( .x(\U6/nl ), .a(l[6]) );
    ao23_1 \U6/Ucl/U1/U1  ( .x(l[6]), .a(n7), .b(l[6]), .c(n2), .d(\U6/ni ), 
        .e(\U6/nh ) );
    ao23_1 \U6/Uch/U1/U1  ( .x(h[6]), .a(n7), .b(h[6]), .c(n2), .d(i[6]), .e(
        \U6/nl ) );
    inv_1 \U5/Uii  ( .x(\U5/ni ), .a(i[5]) );
    inv_1 \U5/Uih  ( .x(\U5/nh ), .a(h[5]) );
    inv_1 \U5/Uil  ( .x(\U5/nl ), .a(l[5]) );
    ao23_1 \U5/Ucl/U1/U1  ( .x(l[5]), .a(n7), .b(l[5]), .c(n2), .d(\U5/ni ), 
        .e(\U5/nh ) );
    ao23_1 \U5/Uch/U1/U1  ( .x(h[5]), .a(n7), .b(h[5]), .c(n2), .d(i[5]), .e(
        \U5/nl ) );
    inv_1 \U4/Uii  ( .x(\U4/ni ), .a(i[4]) );
    inv_1 \U4/Uih  ( .x(\U4/nh ), .a(h[4]) );
    inv_1 \U4/Uil  ( .x(\U4/nl ), .a(l[4]) );
    ao23_1 \U4/Ucl/U1/U1  ( .x(l[4]), .a(n6), .b(l[4]), .c(n2), .d(\U4/ni ), 
        .e(\U4/nh ) );
    ao23_1 \U4/Uch/U1/U1  ( .x(h[4]), .a(n6), .b(h[4]), .c(n2), .d(i[4]), .e(
        \U4/nl ) );
    inv_1 \U3/Uii  ( .x(\U3/ni ), .a(i[3]) );
    inv_1 \U3/Uih  ( .x(\U3/nh ), .a(h[3]) );
    inv_1 \U3/Uil  ( .x(\U3/nl ), .a(l[3]) );
    ao23_1 \U3/Ucl/U1/U1  ( .x(l[3]), .a(n6), .b(l[3]), .c(n2), .d(\U3/ni ), 
        .e(\U3/nh ) );
    ao23_1 \U3/Uch/U1/U1  ( .x(h[3]), .a(n8), .b(h[3]), .c(n1), .d(i[3]), .e(
        \U3/nl ) );
    inv_1 \U2/Uii  ( .x(\U2/ni ), .a(i[2]) );
    inv_1 \U2/Uih  ( .x(\U2/nh ), .a(h[2]) );
    inv_1 \U2/Uil  ( .x(\U2/nl ), .a(l[2]) );
    ao23_1 \U2/Ucl/U1/U1  ( .x(l[2]), .a(n8), .b(l[2]), .c(n1), .d(\U2/ni ), 
        .e(\U2/nh ) );
    ao23_1 \U2/Uch/U1/U1  ( .x(h[2]), .a(n8), .b(h[2]), .c(n1), .d(i[2]), .e(
        \U2/nl ) );
    inv_1 \U1/Uii  ( .x(\U1/ni ), .a(i[1]) );
    inv_1 \U1/Uih  ( .x(\U1/nh ), .a(h[1]) );
    inv_1 \U1/Uil  ( .x(\U1/nl ), .a(l[1]) );
    ao23_1 \U1/Ucl/U1/U1  ( .x(l[1]), .a(n8), .b(l[1]), .c(n1), .d(\U1/ni ), 
        .e(\U1/nh ) );
    ao23_1 \U1/Uch/U1/U1  ( .x(h[1]), .a(n8), .b(h[1]), .c(n1), .d(i[1]), .e(
        \U1/nl ) );
    inv_1 \U0/Uii  ( .x(\U0/ni ), .a(i[0]) );
    inv_1 \U0/Uih  ( .x(\U0/nh ), .a(h[0]) );
    inv_1 \U0/Uil  ( .x(\U0/nl ), .a(l[0]) );
    ao23_1 \U0/Ucl/U1/U1  ( .x(l[0]), .a(n8), .b(l[0]), .c(n1), .d(\U0/ni ), 
        .e(\U0/nh ) );
    ao23_1 \U0/Uch/U1/U1  ( .x(h[0]), .a(n8), .b(h[0]), .c(n1), .d(i[0]), .e(
        \U0/nl ) );
    buf_16 U1 ( .x(n1), .a(n12) );
    buf_16 U2 ( .x(n2), .a(n12) );
    buf_16 U3 ( .x(n3), .a(n12) );
    buf_16 U4 ( .x(n4), .a(n11) );
    buf_16 U5 ( .x(n5), .a(n11) );
    buf_16 U6 ( .x(n6), .a(n11) );
    buf_16 U7 ( .x(n7), .a(n10) );
    buf_16 U8 ( .x(n8), .a(n10) );
    buf_16 U9 ( .x(n9), .a(n10) );
    buf_16 U10 ( .x(n10), .a(req) );
    buf_16 U11 ( .x(n11), .a(req) );
    buf_16 U12 ( .x(n12), .a(req) );
endmodule


module latch_ctrl_2 ( rin, ain, rout, aout, en, reset );
input  rin, aout, reset;
output ain, rout, en;
    wire nreset, na, n1, a, N6, N5, n3, \c_rout/ob , n_rout;
    inv_1 U0 ( .x(nreset), .a(reset) );
    nor2_1 U1 ( .x(ain), .a(na), .b(n1) );
    inv_1 U2 ( .x(na), .a(a) );
    inv_1 U3 ( .x(N6), .a(N5) );
    and2_1 C9 ( .x(n3), .a(na), .b(N6) );
    or2_1 C11 ( .x(N5), .a(rout), .b(aout) );
    oa21_1 \c_na/__tmp99/U1  ( .x(a), .a(n1), .b(a), .c(rin) );
    oai21_1 \c_rout/U1  ( .x(\c_rout/ob ), .a(aout), .b(n_rout), .c(na) );
    nand2_1 \c_rout/U2  ( .x(n_rout), .a(nreset), .b(\c_rout/ob ) );
    buf_1 U4 ( .x(en), .a(n3) );
    inv_2 U5 ( .x(rout), .a(n_rout) );
    buf_1 U6 ( .x(n1), .a(n3) );
endmodule


module matched_delay_m2cp_resp_tic ( x, a );
input  a;
output x;
    assign x = a;
endmodule


module m2cp_tic ( req_in, ts_o, sel_o, mult_o, we_o, prd_o, seq_o, adr_o, 
    dat_o, ain, ic_seq, ic_pred, ic_size, ic_itag, ic_wd, ic_lock, ic_a, 
    ic_rnw, ic_col, ic_ack, req_out, ts_i, we_i, err_i, rty_i, acc_i, dat_i, 
    aout, ir_rd, ir_err, ir_rnw, ir_ack, tag_id, reset );
input  [2:0] ts_o;
input  [3:0] sel_o;
input  [31:0] adr_o;
input  [31:0] dat_o;
output [1:0] ic_seq;
output [1:0] ic_pred;
output [3:0] ic_size;
output [9:0] ic_itag;
output [63:0] ic_wd;
output [1:0] ic_lock;
output [63:0] ic_a;
output [1:0] ic_rnw;
output [5:0] ic_col;
output [2:0] ts_i;
output [31:0] dat_i;
input  [63:0] ir_rd;
input  [1:0] ir_err;
input  [1:0] ir_rnw;
input  [4:0] tag_id;
input  req_in, mult_o, we_o, prd_o, seq_o, ic_ack, aout, reset;
output ain, req_out, we_i, err_i, rty_i, acc_i, ir_ack;
    wire req_in_delayed, n8, \data[15] , \data[14] , \data[13] , \data[12] , 
        \data[11] , \data[10] , \data[9] , \data[8] , \data[7] , \data[6] , 
        \data[5] , \data[4] , \data[3] , \data[2] , \data[1] , \data[0] , 
        complete_delayed, en, _26_net_, n72, n77, _27_net_, _24_net_, n112, 
        n124, n118, n206, n208, n210, n197, n199, n202, n201, n203, n204, 
        \size[1] , n83, n84, n89, n205, n64, n2, n90, n97, n198, n3, n98, n87, 
        n63, n4, n88, n85, n5, n86, n290, n289, n288, n79, n277, n270, n273, 
        n276, n266, n269, n283, n282, n281, n298, n70, n68, n213, n223, n71, 
        n80, n291, n284, n287, n280, n99, n100, n95, n96, n93, n94, n91, n92, 
        n81, all_r, n65, n66, n67, n69, n212, n300, n294, n302, n296, n306, 
        n292, n304, low_ir_rd, n73, n74, n75, n76, complete, n82, n200, n207, 
        n209, n211, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, 
        n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, 
        n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, 
        n258, n259, n260, n261, n262, n263, n265, n264, n268, n267, n272, n271, 
        n275, n274, n279, n278, n286, n285, n293, n295, n297, n299, n301, n303, 
        n305, n307, n222, n221, n220, n219, n218, n217, n216, n215, all_w, 
        n214, high_ir_rd, \size[0] , n308, n182, n179, n176, n173, n194, n191, 
        n188, n185, n158, n155, n152, n149, n170, n167, n164, n161, n134, n131, 
        n128, n125, n146, n143, n140, n137, n110, n107, n104, n101, n122, n119, 
        n116, n113, n183, n184, n180, n181, n177, n178, n174, n175, n195, n196, 
        n192, n193, n189, n190, n186, n187, n159, n160, n156, n157, n153, n154, 
        n150, n151, n171, n172, n168, n169, n165, n166, n162, n163, n135, n136, 
        n132, n133, n129, n130, n126, n127, n147, n148, n144, n145, n141, n142, 
        n138, n139, n111, n108, n109, n105, n106, n102, n103, n123, n120, n121, 
        n117, n114, n115, n7, n6, n1, _28_net_, comp_basic, 
        \all_read/__tmp99/loop , comp_rd, _25_net_, \Ucol2/ni , \Ucol2/nh , 
        \Ucol2/nl , n11, \Ucol1/ni , \Ucol1/nh , \Ucol1/nl , n9, \Ucol0/ni , 
        \Ucol0/nh , \Ucol0/nl , n10, \Utag4/ni , \Utag4/nh , \Utag4/nl , 
        \Utag3/ni , \Utag3/nh , \Utag3/nl , \Utag2/ni , \Utag2/nh , \Utag2/nl , 
        \Utag1/ni , \Utag1/nh , \Utag1/nl , \Utag0/ni , \Utag0/nh , \Utag0/nl , 
        \Usze1/ni , \Usze1/nh , \Usze1/nl , \Usze0/ni , \Usze0/nh , \Usze0/nl , 
        \Urnw/ni , \Urnw/nh , \Urnw/nl , \Ulock/ni , \Ulock/nh , \Ulock/nl , 
        \Upred/ni , \Upred/nh , \Upred/nl , \Useq/ni , \Useq/nh , \Useq/nl , 
        n78;
    assign ain = ic_ack;
    assign ts_i[2] = 1'b0;
    assign ts_i[1] = 1'b0;
    assign ts_i[0] = 1'b0;
    assign rty_i = 1'b0;
    assign acc_i = 1'b0;
    matched_delay_m2cp_com_tic U130 ( .x(req_in_delayed), .a(req_in) );
    sr2dr_word_5 Uwd ( .i({dat_o[31], dat_o[30], dat_o[29], dat_o[28], 
        dat_o[27], dat_o[26], dat_o[25], dat_o[24], dat_o[23], dat_o[22], 
        dat_o[21], dat_o[20], dat_o[19], dat_o[18], dat_o[17], dat_o[16], 
        \data[15] , \data[14] , \data[13] , \data[12] , \data[11] , \data[10] , 
        \data[9] , \data[8] , \data[7] , \data[6] , \data[5] , \data[4] , 
        \data[3] , \data[2] , \data[1] , \data[0] }), .req(n8), .h(ic_wd
        [63:32]), .l(ic_wd[31:0]) );
    sr2dr_word_4 Ua ( .i(adr_o), .req(n8), .h(ic_a[63:32]), .l(ic_a[31:0]) );
    latch_ctrl_2 lc ( .rin(complete_delayed), .ain(ir_ack), .rout(req_out), 
        .aout(aout), .en(en), .reset(reset) );
    nand2_1 U61 ( .x(_26_net_), .a(n72), .b(n77) );
    and2_1 U274 ( .x(_27_net_), .a(ir_rnw[1]), .b(ir_err[0]) );
    inv_1 U275 ( .x(_24_net_), .a(we_o) );
    inv_1 U2 ( .x(n112), .a(ir_rd[4]) );
    inv_1 U3 ( .x(n124), .a(ir_rd[0]) );
    inv_1 U4 ( .x(n118), .a(ir_rd[2]) );
    inv_1 U5 ( .x(n206), .a(dat_o[28]) );
    inv_1 U6 ( .x(n208), .a(dat_o[27]) );
    inv_1 U7 ( .x(n210), .a(dat_o[26]) );
    inv_1 U8 ( .x(n197), .a(dat_o[25]) );
    inv_1 U9 ( .x(n199), .a(dat_o[24]) );
    inv_1 U10 ( .x(n202), .a(dat_o[15]) );
    inv_1 U11 ( .x(n201), .a(dat_o[31]) );
    inv_1 U12 ( .x(n203), .a(dat_o[30]) );
    inv_1 U13 ( .x(n204), .a(dat_o[29]) );
    nor2_1 U14 ( .x(\size[1] ), .a(n83), .b(n84) );
    inv_1 U15 ( .x(n72), .a(ir_rnw[0]) );
    oa21_1 U16 ( .x(n89), .a(n205), .b(n64), .c(n2) );
    inv_1 U24 ( .x(n2), .a(n90) );
    inv_1 U17 ( .x(n205), .a(dat_o[13]) );
    inv_1 U18 ( .x(n64), .a(sel_o[1]) );
    oa21_1 U19 ( .x(n97), .a(n198), .b(n64), .c(n3) );
    inv_1 U276 ( .x(n3), .a(n98) );
    inv_1 U20 ( .x(n198), .a(dat_o[9]) );
    oa21_1 U21 ( .x(n87), .a(n63), .b(n64), .c(n4) );
    inv_1 U277 ( .x(n4), .a(n88) );
    inv_1 U22 ( .x(n63), .a(dat_o[14]) );
    oa21_1 U23 ( .x(n85), .a(n202), .b(n64), .c(n5) );
    inv_1 U278 ( .x(n5), .a(n86) );
    nand2_1 U25 ( .x(n290), .a(n289), .b(n288) );
    nand2_1 U26 ( .x(n79), .a(n277), .b(n270) );
    nor2_1 U27 ( .x(n277), .a(n273), .b(n276) );
    nor2_1 U28 ( .x(n270), .a(n266), .b(n269) );
    nand2_1 U29 ( .x(n283), .a(n282), .b(n281) );
    nand2_1 U30 ( .x(n298), .a(dat_o[20]), .b(n70) );
    inv_1 U31 ( .x(n70), .a(n68) );
    nand2_1 U32 ( .x(n213), .a(n223), .b(n71) );
    nand2_1 U33 ( .x(n80), .a(n291), .b(n284) );
    nor2_1 U34 ( .x(n291), .a(n287), .b(n290) );
    nor2_1 U35 ( .x(n284), .a(n280), .b(n283) );
    aoi21_1 U36 ( .x(n99), .a(dat_o[8]), .b(n71), .c(n100) );
    aoi21_1 U37 ( .x(n95), .a(dat_o[10]), .b(n71), .c(n96) );
    aoi21_1 U38 ( .x(n93), .a(dat_o[11]), .b(n71), .c(n94) );
    aoi21_1 U39 ( .x(n91), .a(dat_o[12]), .b(n71), .c(n92) );
    inv_1 U40 ( .x(n81), .a(all_r) );
    buf_1 U41 ( .x(n65), .a(sel_o[0]) );
    nand2_1 U42 ( .x(n84), .a(sel_o[0]), .b(n71) );
    inv_1 U43 ( .x(n66), .a(sel_o[3]) );
    inv_1 U44 ( .x(n67), .a(n66) );
    inv_1 U45 ( .x(n68), .a(sel_o[2]) );
    inv_1 U46 ( .x(n69), .a(n68) );
    nand2_1 U48 ( .x(n83), .a(n70), .b(n67) );
    nand3i_1 U49 ( .x(n212), .a(sel_o[1]), .b(n67), .c(n70) );
    nor2_1 U50 ( .x(n223), .a(n70), .b(n67) );
    nand2_1 U51 ( .x(n300), .a(dat_o[19]), .b(n69) );
    nand2_1 U52 ( .x(n294), .a(dat_o[22]), .b(n69) );
    nand2_1 U53 ( .x(n302), .a(dat_o[18]), .b(n69) );
    nand2_1 U54 ( .x(n296), .a(dat_o[21]), .b(n69) );
    nand2_1 U55 ( .x(n306), .a(dat_o[16]), .b(n69) );
    nand2_1 U56 ( .x(n292), .a(dat_o[23]), .b(n69) );
    nand2_1 U57 ( .x(n304), .a(dat_o[17]), .b(n69) );
    buf_1 U58 ( .x(n71), .a(sel_o[1]) );
    nand4_1 U60 ( .x(low_ir_rd), .a(n73), .b(n74), .c(n75), .d(n76) );
    nand2_1 U62 ( .x(complete), .a(n81), .b(n82) );
    matched_delay_m2cp_resp_tic mdel ( .x(complete_delayed), .a(complete) );
    inv_1 U63 ( .x(n200), .a(dat_o[8]) );
    inv_1 U64 ( .x(n207), .a(dat_o[12]) );
    inv_1 U65 ( .x(n209), .a(dat_o[11]) );
    inv_1 U66 ( .x(n211), .a(dat_o[10]) );
    nand4_1 U67 ( .x(n224), .a(n225), .b(n226), .c(n227), .d(n228) );
    nand4_1 U68 ( .x(n229), .a(n230), .b(n231), .c(n232), .d(n233) );
    nor2_1 U69 ( .x(n76), .a(n224), .b(n229) );
    nand4_1 U70 ( .x(n234), .a(n235), .b(n236), .c(n237), .d(n238) );
    nand4_1 U71 ( .x(n239), .a(n240), .b(n241), .c(n242), .d(n243) );
    nor2_1 U72 ( .x(n75), .a(n234), .b(n239) );
    nand4_1 U73 ( .x(n244), .a(n245), .b(n246), .c(n247), .d(n248) );
    nand4_1 U74 ( .x(n249), .a(n250), .b(n251), .c(n252), .d(n253) );
    nor2_1 U75 ( .x(n74), .a(n244), .b(n249) );
    nand4_1 U76 ( .x(n254), .a(n255), .b(n256), .c(n257), .d(n258) );
    nand4_1 U77 ( .x(n259), .a(n260), .b(n261), .c(n262), .d(n263) );
    nor2_1 U78 ( .x(n73), .a(n254), .b(n259) );
    nand2_1 U79 ( .x(n266), .a(n265), .b(n264) );
    nand2_1 U80 ( .x(n269), .a(n268), .b(n267) );
    nand2_1 U81 ( .x(n273), .a(n272), .b(n271) );
    nand2_1 U82 ( .x(n276), .a(n275), .b(n274) );
    nand2_1 U83 ( .x(n280), .a(n279), .b(n278) );
    nand2_1 U84 ( .x(n287), .a(n286), .b(n285) );
    nand2_1 U85 ( .x(n86), .a(n292), .b(n293) );
    nand2_1 U86 ( .x(n88), .a(n294), .b(n295) );
    nand2_1 U87 ( .x(n90), .a(n296), .b(n297) );
    nand2_1 U88 ( .x(n92), .a(n298), .b(n299) );
    nand2_1 U89 ( .x(n94), .a(n300), .b(n301) );
    nand2_1 U90 ( .x(n96), .a(n302), .b(n303) );
    nand2_1 U91 ( .x(n98), .a(n304), .b(n305) );
    nand2_1 U92 ( .x(n100), .a(n306), .b(n307) );
    inv_1 U93 ( .x(n222), .a(dat_o[0]) );
    inv_1 U94 ( .x(n221), .a(dat_o[1]) );
    inv_1 U95 ( .x(n220), .a(dat_o[2]) );
    inv_1 U96 ( .x(n219), .a(dat_o[3]) );
    inv_1 U97 ( .x(n218), .a(dat_o[4]) );
    inv_1 U98 ( .x(n217), .a(dat_o[5]) );
    inv_1 U99 ( .x(n216), .a(dat_o[6]) );
    inv_1 U100 ( .x(n215), .a(dat_o[7]) );
    inv_1 U101 ( .x(n77), .a(ir_rnw[1]) );
    inv_1 U103 ( .x(n82), .a(all_w) );
    nand2_1 U104 ( .x(n293), .a(dat_o[31]), .b(n67) );
    nand2_1 U105 ( .x(n295), .a(dat_o[30]), .b(n67) );
    nand2_1 U106 ( .x(n297), .a(dat_o[29]), .b(n67) );
    nand2_1 U107 ( .x(n299), .a(dat_o[28]), .b(n67) );
    nand2_1 U108 ( .x(n301), .a(dat_o[27]), .b(n67) );
    nand2_1 U109 ( .x(n303), .a(dat_o[26]), .b(n67) );
    nand2_1 U110 ( .x(n305), .a(dat_o[25]), .b(n67) );
    nand2_1 U111 ( .x(n307), .a(dat_o[24]), .b(n67) );
    mux2i_1 U113 ( .x(\data[0] ), .d0(n99), .sl(n65), .d1(n222) );
    mux2i_1 U114 ( .x(\data[10] ), .d0(n211), .sl(n214), .d1(n210) );
    mux2i_1 U115 ( .x(\data[11] ), .d0(n209), .sl(n214), .d1(n208) );
    mux2i_1 U116 ( .x(\data[12] ), .d0(n207), .sl(n214), .d1(n206) );
    mux2i_1 U117 ( .x(\data[13] ), .d0(n205), .sl(n214), .d1(n204) );
    mux2i_1 U118 ( .x(\data[14] ), .d0(n63), .sl(n214), .d1(n203) );
    mux2i_1 U119 ( .x(\data[15] ), .d0(n202), .sl(n214), .d1(n201) );
    mux2i_1 U120 ( .x(\data[1] ), .d0(n97), .sl(n65), .d1(n221) );
    mux2i_1 U121 ( .x(\data[2] ), .d0(n95), .sl(n65), .d1(n220) );
    mux2i_1 U122 ( .x(\data[3] ), .d0(n93), .sl(n65), .d1(n219) );
    mux2i_1 U123 ( .x(\data[4] ), .d0(n91), .sl(n65), .d1(n218) );
    mux2i_1 U124 ( .x(\data[5] ), .d0(n89), .sl(n65), .d1(n217) );
    mux2i_1 U125 ( .x(\data[6] ), .d0(n87), .sl(n65), .d1(n216) );
    mux2i_1 U126 ( .x(\data[7] ), .d0(n85), .sl(n65), .d1(n215) );
    mux2i_1 U127 ( .x(\data[8] ), .d0(n200), .sl(n214), .d1(n199) );
    mux2i_1 U128 ( .x(\data[9] ), .d0(n198), .sl(n214), .d1(n197) );
    nor2_1 U129 ( .x(high_ir_rd), .a(n79), .b(n80) );
    mux2i_1 U131 ( .x(\size[0] ), .d0(n212), .sl(n65), .d1(n213) );
    nand2i_1 U132 ( .x(n308), .a(sel_o[1]), .b(n70) );
    inv_1 U133 ( .x(n255), .a(n182) );
    inv_1 U134 ( .x(n256), .a(n179) );
    inv_1 U135 ( .x(n257), .a(n176) );
    inv_1 U136 ( .x(n258), .a(n173) );
    inv_1 U137 ( .x(n260), .a(n194) );
    inv_1 U138 ( .x(n261), .a(n191) );
    inv_1 U139 ( .x(n262), .a(n188) );
    inv_1 U140 ( .x(n263), .a(n185) );
    inv_1 U141 ( .x(n245), .a(n158) );
    inv_1 U142 ( .x(n246), .a(n155) );
    inv_1 U143 ( .x(n247), .a(n152) );
    inv_1 U144 ( .x(n248), .a(n149) );
    inv_1 U145 ( .x(n250), .a(n170) );
    inv_1 U146 ( .x(n251), .a(n167) );
    inv_1 U147 ( .x(n252), .a(n164) );
    inv_1 U148 ( .x(n253), .a(n161) );
    inv_1 U149 ( .x(n235), .a(n134) );
    inv_1 U150 ( .x(n236), .a(n131) );
    inv_1 U151 ( .x(n237), .a(n128) );
    inv_1 U152 ( .x(n238), .a(n125) );
    inv_1 U153 ( .x(n240), .a(n146) );
    inv_1 U154 ( .x(n241), .a(n143) );
    inv_1 U155 ( .x(n242), .a(n140) );
    inv_1 U156 ( .x(n243), .a(n137) );
    inv_1 U157 ( .x(n225), .a(n110) );
    inv_1 U158 ( .x(n226), .a(n107) );
    inv_1 U159 ( .x(n227), .a(n104) );
    inv_1 U160 ( .x(n228), .a(n101) );
    inv_1 U161 ( .x(n230), .a(n122) );
    inv_1 U162 ( .x(n231), .a(n119) );
    inv_1 U163 ( .x(n232), .a(n116) );
    inv_1 U164 ( .x(n233), .a(n113) );
    nor2_1 U165 ( .x(n272), .a(n252), .b(n253) );
    nor2_1 U166 ( .x(n271), .a(n250), .b(n251) );
    nor2_1 U167 ( .x(n275), .a(n247), .b(n248) );
    nor2_1 U168 ( .x(n274), .a(n245), .b(n246) );
    nor2_1 U169 ( .x(n265), .a(n262), .b(n263) );
    nor2_1 U170 ( .x(n264), .a(n260), .b(n261) );
    nor2_1 U171 ( .x(n268), .a(n257), .b(n258) );
    nor2_1 U172 ( .x(n267), .a(n255), .b(n256) );
    nor2_1 U173 ( .x(n286), .a(n232), .b(n233) );
    nor2_1 U174 ( .x(n285), .a(n230), .b(n231) );
    nor2_1 U175 ( .x(n289), .a(n227), .b(n228) );
    nor2_1 U176 ( .x(n288), .a(n225), .b(n226) );
    nor2_1 U177 ( .x(n279), .a(n242), .b(n243) );
    nor2_1 U178 ( .x(n278), .a(n240), .b(n241) );
    nor2_1 U179 ( .x(n282), .a(n237), .b(n238) );
    nor2_1 U180 ( .x(n281), .a(n235), .b(n236) );
    nand2_1 U181 ( .x(n182), .a(n183), .b(n184) );
    nand2_1 U182 ( .x(n179), .a(n180), .b(n181) );
    nand2_1 U183 ( .x(n176), .a(n177), .b(n178) );
    nand2_1 U184 ( .x(n173), .a(n174), .b(n175) );
    nand2_1 U185 ( .x(n194), .a(n195), .b(n196) );
    nand2_1 U186 ( .x(n191), .a(n192), .b(n193) );
    nand2_1 U187 ( .x(n188), .a(n189), .b(n190) );
    nand2_1 U188 ( .x(n185), .a(n186), .b(n187) );
    nand2_1 U189 ( .x(n158), .a(n159), .b(n160) );
    nand2_1 U190 ( .x(n155), .a(n156), .b(n157) );
    nand2_1 U191 ( .x(n152), .a(n153), .b(n154) );
    nand2_1 U192 ( .x(n149), .a(n150), .b(n151) );
    nand2_1 U193 ( .x(n170), .a(n171), .b(n172) );
    nand2_1 U194 ( .x(n167), .a(n168), .b(n169) );
    nand2_1 U195 ( .x(n164), .a(n165), .b(n166) );
    nand2_1 U196 ( .x(n161), .a(n162), .b(n163) );
    nand2_1 U197 ( .x(n134), .a(n135), .b(n136) );
    nand2_1 U198 ( .x(n131), .a(n132), .b(n133) );
    nand2_1 U199 ( .x(n128), .a(n129), .b(n130) );
    nand2_1 U200 ( .x(n125), .a(n126), .b(n127) );
    nand2_1 U201 ( .x(n146), .a(n147), .b(n148) );
    nand2_1 U202 ( .x(n143), .a(n144), .b(n145) );
    nand2_1 U203 ( .x(n140), .a(n141), .b(n142) );
    nand2_1 U204 ( .x(n137), .a(n138), .b(n139) );
    nand2_1 U205 ( .x(n110), .a(n111), .b(n112) );
    nand2_1 U206 ( .x(n107), .a(n108), .b(n109) );
    nand2_1 U207 ( .x(n104), .a(n105), .b(n106) );
    nand2_1 U208 ( .x(n101), .a(n102), .b(n103) );
    nand2_1 U209 ( .x(n122), .a(n123), .b(n124) );
    nand2_1 U210 ( .x(n119), .a(n120), .b(n121) );
    nand2_1 U211 ( .x(n116), .a(n117), .b(n118) );
    nand2_1 U212 ( .x(n113), .a(n114), .b(n115) );
    inv_1 U213 ( .x(n183), .a(ir_rd[60]) );
    inv_1 U214 ( .x(n184), .a(ir_rd[28]) );
    inv_1 U215 ( .x(n180), .a(ir_rd[61]) );
    inv_1 U216 ( .x(n181), .a(ir_rd[29]) );
    inv_1 U217 ( .x(n177), .a(ir_rd[62]) );
    inv_1 U218 ( .x(n178), .a(ir_rd[30]) );
    inv_1 U219 ( .x(n174), .a(ir_rd[63]) );
    inv_1 U220 ( .x(n175), .a(ir_rd[31]) );
    inv_1 U221 ( .x(n195), .a(ir_rd[56]) );
    inv_1 U222 ( .x(n196), .a(ir_rd[24]) );
    inv_1 U223 ( .x(n192), .a(ir_rd[57]) );
    inv_1 U224 ( .x(n193), .a(ir_rd[25]) );
    inv_1 U225 ( .x(n189), .a(ir_rd[58]) );
    inv_1 U226 ( .x(n190), .a(ir_rd[26]) );
    inv_1 U227 ( .x(n186), .a(ir_rd[59]) );
    inv_1 U228 ( .x(n187), .a(ir_rd[27]) );
    inv_1 U229 ( .x(n159), .a(ir_rd[52]) );
    inv_1 U230 ( .x(n160), .a(ir_rd[20]) );
    inv_1 U231 ( .x(n156), .a(ir_rd[53]) );
    inv_1 U232 ( .x(n157), .a(ir_rd[21]) );
    inv_1 U233 ( .x(n153), .a(ir_rd[54]) );
    inv_1 U234 ( .x(n154), .a(ir_rd[22]) );
    inv_1 U235 ( .x(n150), .a(ir_rd[55]) );
    inv_1 U236 ( .x(n151), .a(ir_rd[23]) );
    inv_1 U237 ( .x(n171), .a(ir_rd[48]) );
    inv_1 U238 ( .x(n172), .a(ir_rd[16]) );
    inv_1 U239 ( .x(n168), .a(ir_rd[49]) );
    inv_1 U240 ( .x(n169), .a(ir_rd[17]) );
    inv_1 U241 ( .x(n165), .a(ir_rd[50]) );
    inv_1 U242 ( .x(n166), .a(ir_rd[18]) );
    inv_1 U243 ( .x(n162), .a(ir_rd[51]) );
    inv_1 U244 ( .x(n163), .a(ir_rd[19]) );
    inv_1 U245 ( .x(n135), .a(ir_rd[44]) );
    inv_1 U246 ( .x(n136), .a(ir_rd[12]) );
    inv_1 U247 ( .x(n132), .a(ir_rd[45]) );
    inv_1 U248 ( .x(n133), .a(ir_rd[13]) );
    inv_1 U249 ( .x(n129), .a(ir_rd[46]) );
    inv_1 U250 ( .x(n130), .a(ir_rd[14]) );
    inv_1 U251 ( .x(n126), .a(ir_rd[47]) );
    inv_1 U252 ( .x(n127), .a(ir_rd[15]) );
    inv_1 U253 ( .x(n147), .a(ir_rd[40]) );
    inv_1 U254 ( .x(n148), .a(ir_rd[8]) );
    inv_1 U255 ( .x(n144), .a(ir_rd[41]) );
    inv_1 U256 ( .x(n145), .a(ir_rd[9]) );
    inv_1 U257 ( .x(n141), .a(ir_rd[42]) );
    inv_1 U258 ( .x(n142), .a(ir_rd[10]) );
    inv_1 U259 ( .x(n138), .a(ir_rd[43]) );
    inv_1 U260 ( .x(n139), .a(ir_rd[11]) );
    inv_1 U261 ( .x(n111), .a(ir_rd[36]) );
    inv_1 U262 ( .x(n108), .a(ir_rd[37]) );
    inv_1 U263 ( .x(n109), .a(ir_rd[5]) );
    inv_1 U264 ( .x(n105), .a(ir_rd[38]) );
    inv_1 U265 ( .x(n106), .a(ir_rd[6]) );
    inv_1 U266 ( .x(n102), .a(ir_rd[39]) );
    inv_1 U267 ( .x(n103), .a(ir_rd[7]) );
    inv_1 U268 ( .x(n123), .a(ir_rd[32]) );
    inv_1 U269 ( .x(n120), .a(ir_rd[33]) );
    inv_1 U270 ( .x(n121), .a(ir_rd[1]) );
    inv_1 U271 ( .x(n117), .a(ir_rd[34]) );
    inv_1 U272 ( .x(n114), .a(ir_rd[35]) );
    inv_1 U273 ( .x(n115), .a(ir_rd[3]) );
    latn_1 \dat_i_reg[30]  ( .q(dat_i[30]), .d(ir_rd[62]), .g(n7) );
    latn_1 \dat_i_reg[28]  ( .q(dat_i[28]), .d(ir_rd[60]), .g(n7) );
    latn_1 \dat_i_reg[27]  ( .q(dat_i[27]), .d(ir_rd[59]), .g(n7) );
    latn_1 \dat_i_reg[26]  ( .q(dat_i[26]), .d(ir_rd[58]), .g(n7) );
    latn_1 \dat_i_reg[25]  ( .q(dat_i[25]), .d(ir_rd[57]), .g(n7) );
    latn_1 \dat_i_reg[24]  ( .q(dat_i[24]), .d(ir_rd[56]), .g(n7) );
    latn_1 \dat_i_reg[22]  ( .q(dat_i[22]), .d(ir_rd[54]), .g(n7) );
    latn_1 \dat_i_reg[20]  ( .q(dat_i[20]), .d(ir_rd[52]), .g(n7) );
    latn_1 \dat_i_reg[19]  ( .q(dat_i[19]), .d(ir_rd[51]), .g(n7) );
    latn_1 \dat_i_reg[18]  ( .q(dat_i[18]), .d(ir_rd[50]), .g(n7) );
    latn_1 \dat_i_reg[17]  ( .q(dat_i[17]), .d(ir_rd[49]), .g(n7) );
    latn_1 \dat_i_reg[16]  ( .q(dat_i[16]), .d(ir_rd[48]), .g(n6) );
    latn_1 \dat_i_reg[14]  ( .q(dat_i[14]), .d(ir_rd[46]), .g(n6) );
    latn_1 \dat_i_reg[12]  ( .q(dat_i[12]), .d(ir_rd[44]), .g(n6) );
    latn_1 \dat_i_reg[10]  ( .q(dat_i[10]), .d(ir_rd[42]), .g(n6) );
    latn_1 \dat_i_reg[8]  ( .q(dat_i[8]), .d(ir_rd[40]), .g(n6) );
    latn_1 \dat_i_reg[6]  ( .q(dat_i[6]), .d(ir_rd[38]), .g(n6) );
    latn_1 \dat_i_reg[4]  ( .q(dat_i[4]), .d(ir_rd[36]), .g(n6) );
    latn_1 \dat_i_reg[3]  ( .q(dat_i[3]), .d(ir_rd[35]), .g(n1) );
    latn_1 \dat_i_reg[2]  ( .q(dat_i[2]), .d(ir_rd[34]), .g(n1) );
    latn_1 \dat_i_reg[1]  ( .q(dat_i[1]), .d(ir_rd[33]), .g(n1) );
    latn_1 \dat_i_reg[0]  ( .q(dat_i[0]), .d(ir_rd[32]), .g(n1) );
    latn_1 we_i_reg ( .q(we_i), .d(ir_rnw[0]), .g(n1) );
    latn_1 err_i_reg ( .q(err_i), .d(ir_err[1]), .g(n1) );
    latn_1 \dat_i_reg[13]  ( .q(dat_i[13]), .d(ir_rd[45]), .g(n6) );
    latn_1 \dat_i_reg[5]  ( .q(dat_i[5]), .d(ir_rd[37]), .g(n1) );
    latn_1 \dat_i_reg[15]  ( .q(dat_i[15]), .d(ir_rd[47]), .g(n6) );
    latn_1 \dat_i_reg[7]  ( .q(dat_i[7]), .d(ir_rd[39]), .g(n1) );
    latn_1 \dat_i_reg[29]  ( .q(dat_i[29]), .d(ir_rd[61]), .g(n6) );
    latn_1 \dat_i_reg[21]  ( .q(dat_i[21]), .d(ir_rd[53]), .g(n1) );
    latn_1 \dat_i_reg[31]  ( .q(dat_i[31]), .d(ir_rd[63]), .g(n6) );
    latn_1 \dat_i_reg[23]  ( .q(dat_i[23]), .d(ir_rd[55]), .g(n1) );
    latn_1 \dat_i_reg[9]  ( .q(dat_i[9]), .d(ir_rd[41]), .g(n6) );
    latn_1 \dat_i_reg[11]  ( .q(dat_i[11]), .d(ir_rd[43]), .g(n1) );
    oa21_1 \all_write/__tmp99/U1  ( .x(all_w), .a(_28_net_), .b(all_w), .c(
        comp_basic) );
    ao31_1 \all_read/__tmp99/aoi  ( .x(\all_read/__tmp99/loop ), .a(comp_basic
        ), .b(comp_rd), .c(_27_net_), .d(all_r) );
    oa21_1 \all_read/__tmp99/outGate  ( .x(all_r), .a(comp_basic), .b(comp_rd), 
        .c(\all_read/__tmp99/loop ) );
    ao222_1 \rd/__tmp99/U1  ( .x(comp_rd), .a(high_ir_rd), .b(low_ir_rd), .c(
        high_ir_rd), .d(comp_rd), .e(low_ir_rd), .f(comp_rd) );
    ao222_1 \basic/__tmp99/U1  ( .x(comp_basic), .a(_25_net_), .b(_26_net_), 
        .c(_25_net_), .d(comp_basic), .e(_26_net_), .f(comp_basic) );
    inv_1 \Ucol2/Uii  ( .x(\Ucol2/ni ), .a(ts_o[2]) );
    inv_1 \Ucol2/Uih  ( .x(\Ucol2/nh ), .a(ic_col[5]) );
    inv_1 \Ucol2/Uil  ( .x(\Ucol2/nl ), .a(ic_col[2]) );
    ao23_1 \Ucol2/Ucl/U1/U1  ( .x(ic_col[2]), .a(n11), .b(ic_col[2]), .c(n8), 
        .d(\Ucol2/ni ), .e(\Ucol2/nh ) );
    ao23_1 \Ucol2/Uch/U1/U1  ( .x(ic_col[5]), .a(n11), .b(ic_col[5]), .c(n8), 
        .d(ts_o[2]), .e(\Ucol2/nl ) );
    inv_1 \Ucol1/Uii  ( .x(\Ucol1/ni ), .a(ts_o[1]) );
    inv_1 \Ucol1/Uih  ( .x(\Ucol1/nh ), .a(ic_col[4]) );
    inv_1 \Ucol1/Uil  ( .x(\Ucol1/nl ), .a(ic_col[1]) );
    ao23_1 \Ucol1/Ucl/U1/U1  ( .x(ic_col[1]), .a(n11), .b(ic_col[1]), .c(n8), 
        .d(\Ucol1/ni ), .e(\Ucol1/nh ) );
    ao23_1 \Ucol1/Uch/U1/U1  ( .x(ic_col[4]), .a(n11), .b(ic_col[4]), .c(n9), 
        .d(ts_o[1]), .e(\Ucol1/nl ) );
    inv_1 \Ucol0/Uii  ( .x(\Ucol0/ni ), .a(ts_o[0]) );
    inv_1 \Ucol0/Uih  ( .x(\Ucol0/nh ), .a(ic_col[3]) );
    inv_1 \Ucol0/Uil  ( .x(\Ucol0/nl ), .a(ic_col[0]) );
    ao23_1 \Ucol0/Ucl/U1/U1  ( .x(ic_col[0]), .a(n11), .b(ic_col[0]), .c(n10), 
        .d(\Ucol0/ni ), .e(\Ucol0/nh ) );
    ao23_1 \Ucol0/Uch/U1/U1  ( .x(ic_col[3]), .a(n11), .b(ic_col[3]), .c(n9), 
        .d(ts_o[0]), .e(\Ucol0/nl ) );
    inv_1 \Utag4/Uii  ( .x(\Utag4/ni ), .a(tag_id[4]) );
    inv_1 \Utag4/Uih  ( .x(\Utag4/nh ), .a(ic_itag[9]) );
    inv_1 \Utag4/Uil  ( .x(\Utag4/nl ), .a(ic_itag[4]) );
    ao23_1 \Utag4/Ucl/U1/U1  ( .x(ic_itag[4]), .a(n11), .b(ic_itag[4]), .c(n9), 
        .d(\Utag4/ni ), .e(\Utag4/nh ) );
    ao23_1 \Utag4/Uch/U1/U1  ( .x(ic_itag[9]), .a(n10), .b(ic_itag[9]), .c(n9), 
        .d(tag_id[4]), .e(\Utag4/nl ) );
    inv_1 \Utag3/Uii  ( .x(\Utag3/ni ), .a(tag_id[3]) );
    inv_1 \Utag3/Uih  ( .x(\Utag3/nh ), .a(ic_itag[8]) );
    inv_1 \Utag3/Uil  ( .x(\Utag3/nl ), .a(ic_itag[3]) );
    ao23_1 \Utag3/Ucl/U1/U1  ( .x(ic_itag[3]), .a(n10), .b(ic_itag[3]), .c(n9), 
        .d(\Utag3/ni ), .e(\Utag3/nh ) );
    ao23_1 \Utag3/Uch/U1/U1  ( .x(ic_itag[8]), .a(n10), .b(ic_itag[8]), .c(n9), 
        .d(tag_id[3]), .e(\Utag3/nl ) );
    inv_1 \Utag2/Uii  ( .x(\Utag2/ni ), .a(tag_id[2]) );
    inv_1 \Utag2/Uih  ( .x(\Utag2/nh ), .a(ic_itag[7]) );
    inv_1 \Utag2/Uil  ( .x(\Utag2/nl ), .a(ic_itag[2]) );
    ao23_1 \Utag2/Ucl/U1/U1  ( .x(ic_itag[2]), .a(n10), .b(ic_itag[2]), .c(n9), 
        .d(\Utag2/ni ), .e(\Utag2/nh ) );
    ao23_1 \Utag2/Uch/U1/U1  ( .x(ic_itag[7]), .a(n10), .b(ic_itag[7]), .c(n10
        ), .d(tag_id[2]), .e(\Utag2/nl ) );
    inv_1 \Utag1/Uii  ( .x(\Utag1/ni ), .a(tag_id[1]) );
    inv_1 \Utag1/Uih  ( .x(\Utag1/nh ), .a(ic_itag[6]) );
    inv_1 \Utag1/Uil  ( .x(\Utag1/nl ), .a(ic_itag[1]) );
    ao23_1 \Utag1/Ucl/U1/U1  ( .x(ic_itag[1]), .a(n11), .b(ic_itag[1]), .c(n9), 
        .d(\Utag1/ni ), .e(\Utag1/nh ) );
    ao23_1 \Utag1/Uch/U1/U1  ( .x(ic_itag[6]), .a(n11), .b(ic_itag[6]), .c(n9), 
        .d(tag_id[1]), .e(\Utag1/nl ) );
    inv_1 \Utag0/Uii  ( .x(\Utag0/ni ), .a(tag_id[0]) );
    inv_1 \Utag0/Uih  ( .x(\Utag0/nh ), .a(ic_itag[5]) );
    inv_1 \Utag0/Uil  ( .x(\Utag0/nl ), .a(ic_itag[0]) );
    ao23_1 \Utag0/Ucl/U1/U1  ( .x(ic_itag[0]), .a(n11), .b(ic_itag[0]), .c(n8), 
        .d(\Utag0/ni ), .e(\Utag0/nh ) );
    ao23_1 \Utag0/Uch/U1/U1  ( .x(ic_itag[5]), .a(n10), .b(ic_itag[5]), .c(n8), 
        .d(tag_id[0]), .e(\Utag0/nl ) );
    inv_1 \Usze1/Uii  ( .x(\Usze1/ni ), .a(\size[1] ) );
    inv_1 \Usze1/Uih  ( .x(\Usze1/nh ), .a(ic_size[3]) );
    inv_1 \Usze1/Uil  ( .x(\Usze1/nl ), .a(ic_size[1]) );
    ao23_1 \Usze1/Ucl/U1/U1  ( .x(ic_size[1]), .a(n10), .b(ic_size[1]), .c(n9), 
        .d(\Usze1/ni ), .e(\Usze1/nh ) );
    ao23_1 \Usze1/Uch/U1/U1  ( .x(ic_size[3]), .a(n10), .b(ic_size[3]), .c(n9), 
        .d(\size[1] ), .e(\Usze1/nl ) );
    inv_1 \Usze0/Uii  ( .x(\Usze0/ni ), .a(\size[0] ) );
    inv_1 \Usze0/Uih  ( .x(\Usze0/nh ), .a(ic_size[2]) );
    inv_1 \Usze0/Uil  ( .x(\Usze0/nl ), .a(ic_size[0]) );
    ao23_1 \Usze0/Ucl/U1/U1  ( .x(ic_size[0]), .a(n10), .b(ic_size[0]), .c(n9), 
        .d(\Usze0/ni ), .e(\Usze0/nh ) );
    ao23_1 \Usze0/Uch/U1/U1  ( .x(ic_size[2]), .a(n10), .b(ic_size[2]), .c(n9), 
        .d(\size[0] ), .e(\Usze0/nl ) );
    inv_1 \Urnw/Uii  ( .x(\Urnw/ni ), .a(_24_net_) );
    inv_1 \Urnw/Uih  ( .x(\Urnw/nh ), .a(ic_rnw[1]) );
    inv_1 \Urnw/Uil  ( .x(\Urnw/nl ), .a(ic_rnw[0]) );
    ao23_1 \Urnw/Ucl/U1/U1  ( .x(ic_rnw[0]), .a(n10), .b(ic_rnw[0]), .c(n9), 
        .d(\Urnw/ni ), .e(\Urnw/nh ) );
    ao23_1 \Urnw/Uch/U1/U1  ( .x(ic_rnw[1]), .a(n10), .b(ic_rnw[1]), .c(n9), 
        .d(_24_net_), .e(\Urnw/nl ) );
    inv_1 \Ulock/Uii  ( .x(\Ulock/ni ), .a(mult_o) );
    inv_1 \Ulock/Uih  ( .x(\Ulock/nh ), .a(ic_lock[1]) );
    inv_1 \Ulock/Uil  ( .x(\Ulock/nl ), .a(ic_lock[0]) );
    ao23_1 \Ulock/Ucl/U1/U1  ( .x(ic_lock[0]), .a(n11), .b(ic_lock[0]), .c(n9), 
        .d(\Ulock/ni ), .e(\Ulock/nh ) );
    ao23_1 \Ulock/Uch/U1/U1  ( .x(ic_lock[1]), .a(n11), .b(ic_lock[1]), .c(n8), 
        .d(mult_o), .e(\Ulock/nl ) );
    inv_1 \Upred/Uii  ( .x(\Upred/ni ), .a(prd_o) );
    inv_1 \Upred/Uih  ( .x(\Upred/nh ), .a(ic_pred[1]) );
    inv_1 \Upred/Uil  ( .x(\Upred/nl ), .a(ic_pred[0]) );
    ao23_1 \Upred/Ucl/U1/U1  ( .x(ic_pred[0]), .a(n11), .b(ic_pred[0]), .c(n8), 
        .d(\Upred/ni ), .e(\Upred/nh ) );
    ao23_1 \Upred/Uch/U1/U1  ( .x(ic_pred[1]), .a(n10), .b(ic_pred[1]), .c(n8), 
        .d(prd_o), .e(\Upred/nl ) );
    inv_1 \Useq/Uii  ( .x(\Useq/ni ), .a(seq_o) );
    inv_1 \Useq/Uih  ( .x(\Useq/nh ), .a(ic_seq[1]) );
    inv_1 \Useq/Uil  ( .x(\Useq/nl ), .a(ic_seq[0]) );
    ao23_1 \Useq/Ucl/U1/U1  ( .x(ic_seq[0]), .a(n10), .b(ic_seq[0]), .c(n8), 
        .d(\Useq/ni ), .e(\Useq/nh ) );
    ao23_1 \Useq/Uch/U1/U1  ( .x(ic_seq[1]), .a(n11), .b(ic_seq[1]), .c(n8), 
        .d(seq_o), .e(\Useq/nl ) );
    buf_3 U1 ( .x(n1), .a(en) );
    buf_3 U47 ( .x(n7), .a(en) );
    buf_3 U59 ( .x(n6), .a(en) );
    inv_2 U102 ( .x(n214), .a(n308) );
    inv_0 U112 ( .x(n78), .a(ir_err[0]) );
    nand2i_0 U279 ( .x(_28_net_), .a(ir_err[1]), .b(n72) );
    nand2i_0 U280 ( .x(_25_net_), .a(ir_err[1]), .b(n78) );
    buf_16 U281 ( .x(n8), .a(req_in_delayed) );
    buf_16 U282 ( .x(n9), .a(req_in_delayed) );
    buf_16 U283 ( .x(n10), .a(req_in_delayed) );
    buf_16 U284 ( .x(n11), .a(req_in_delayed) );
endmodule


module i_adec_tic ( e_h, e_l, r_h, r_l, ah, al, e_bare, e_dm, e_im, e_wish, 
    r_bare, r_dm, r_im, r_wish, force_bare );
output [3:0] e_h;
output [3:0] e_l;
output [3:0] r_h;
output [3:0] r_l;
input  [31:0] ah;
input  [31:0] al;
input  [3:0] e_bare;
input  [3:0] e_dm;
input  [3:0] e_im;
input  [3:0] e_wish;
input  [3:0] r_bare;
input  [3:0] r_dm;
input  [3:0] r_im;
input  [3:0] r_wish;
input  force_bare;
    wire e_h_0, e_l_3, e_l_2, e_l_0, wish_i, n6, bare_i, im_i, n7, dm_i, 
        \r_l[2] , \r_l[0] , n1, n2, n3, n15, n14, n12;
    assign e_h[3] = 1'b0;
    assign e_h[0] = e_h_0;
    assign e_l[3] = e_l_3;
    assign e_l[2] = e_l_2;
    assign e_l[0] = e_l_0;
    assign r_h[3] = e_l_2;
    assign r_h[2] = e_h_0;
    assign r_h[0] = 1'b0;
    assign r_l[2] = e_l_0;
    assign r_l[0] = e_l_3;
    ao222_1 \U1632/U18/U1/U1  ( .x(wish_i), .a(n6), .b(al[30]), .c(n6), .d(
        wish_i), .e(al[30]), .f(wish_i) );
    ao222_1 \U1633/U18/U1/U1  ( .x(bare_i), .a(n6), .b(ah[30]), .c(n6), .d(
        bare_i), .e(ah[30]), .f(bare_i) );
    ao222_1 \U1634/U18/U1/U1  ( .x(im_i), .a(al[11]), .b(n7), .c(al[11]), .d(
        im_i), .e(n7), .f(im_i) );
    ao222_1 \U1635/U18/U1/U1  ( .x(dm_i), .a(ah[11]), .b(n7), .c(ah[11]), .d(
        dm_i), .e(n7), .f(dm_i) );
    or3_1 U1 ( .x(\r_l[2] ), .a(wish_i), .b(bare_i), .c(force_bare) );
    or2_1 U2 ( .x(r_l[1]), .a(e_l_0), .b(im_i) );
    or2_1 U3 ( .x(\r_l[0] ), .a(dm_i), .b(r_l[1]) );
    nor2_0 U4 ( .x(n1), .a(bare_i), .b(force_bare) );
    aoi21_1 U6 ( .x(n2), .a(n3), .b(im_i), .c(r_h[1]) );
    inv_0 U8 ( .x(n3), .a(force_bare) );
    nor2i_0 U9 ( .x(n15), .a(wish_i), .b(force_bare) );
    nor2i_0 U10 ( .x(n14), .a(dm_i), .b(force_bare) );
    inv_0 U11 ( .x(e_h[1]), .a(n1) );
    buf_1 U15 ( .x(n6), .a(ah[31]) );
    buf_1 U16 ( .x(n7), .a(al[31]) );
    nand2_2 U17 ( .x(e_l_2), .a(n2), .b(n1) );
    buf_1 U18 ( .x(r_h[1]), .a(n14) );
    inv_2 U19 ( .x(e_h_0), .a(n2) );
    buf_3 U20 ( .x(e_l_3), .a(\r_l[0] ) );
    buf_3 U21 ( .x(e_l_0), .a(\r_l[2] ) );
    nand2i_2 U22 ( .x(e_l[1]), .a(n12), .b(n2) );
    buf_1 U23 ( .x(e_h[2]), .a(n15) );
    buf_1 U24 ( .x(r_l[3]), .a(n15) );
    buf_1 U25 ( .x(n12), .a(n15) );
endmodule


module chain_selement_ga_12 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_symbol_8 ( o, txack, txack_last, e, oa, r, txreq );
output [2:0] o;
input  [1:0] e;
input  [1:0] r;
input  oa, txreq;
output txack, txack_last;
    wire ack, net10, \c[0] , \c[1] ;
    chain_selement_ga_12 U1239 ( .Aa(ack), .Br(net10), .Ar(txreq), .Ba(oa) );
    and2_1 \U1229_0_/U8  ( .x(o[0]), .a(\c[0] ), .b(net10) );
    and2_1 \U1229_1_/U8  ( .x(o[1]), .a(\c[1] ), .b(net10) );
    and2_1 \U1229_2_/U8  ( .x(o[2]), .a(e[1]), .b(net10) );
    ao23_1 \U1251/U19/U21/U1/U1  ( .x(txack_last), .a(ack), .b(txack_last), 
        .c(ack), .d(e[1]), .e(e[1]) );
    ao23_1 \U1250/U19/U21/U1/U1  ( .x(txack), .a(ack), .b(txack), .c(ack), .d(
        e[0]), .e(e[0]) );
    ao222_1 \U1210/U18/U1/U1  ( .x(\c[0] ), .a(e[0]), .b(r[0]), .c(e[0]), .d(
        \c[0] ), .e(r[0]), .f(\c[0] ) );
    ao222_1 \U1209/U18/U1/U1  ( .x(\c[1] ), .a(e[0]), .b(r[1]), .c(e[0]), .d(
        \c[1] ), .e(r[1]), .f(\c[1] ) );
endmodule


module chain_selement_ga_13 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_symbol_9 ( o, txack, txack_last, e, oa, r, txreq );
output [2:0] o;
input  [1:0] e;
input  [1:0] r;
input  oa, txreq;
output txack, txack_last;
    wire ack, net10, \c[0] , \c[1] ;
    chain_selement_ga_13 U1239 ( .Aa(ack), .Br(net10), .Ar(txreq), .Ba(oa) );
    and2_1 \U1229_0_/U8  ( .x(o[0]), .a(\c[0] ), .b(net10) );
    and2_1 \U1229_1_/U8  ( .x(o[1]), .a(\c[1] ), .b(net10) );
    and2_1 \U1229_2_/U8  ( .x(o[2]), .a(e[1]), .b(net10) );
    ao23_1 \U1251/U19/U21/U1/U1  ( .x(txack_last), .a(ack), .b(txack_last), 
        .c(ack), .d(e[1]), .e(e[1]) );
    ao23_1 \U1250/U19/U21/U1/U1  ( .x(txack), .a(ack), .b(txack), .c(ack), .d(
        e[0]), .e(e[0]) );
    ao222_1 \U1210/U18/U1/U1  ( .x(\c[0] ), .a(e[0]), .b(r[0]), .c(e[0]), .d(
        \c[0] ), .e(r[0]), .f(\c[0] ) );
    ao222_1 \U1209/U18/U1/U1  ( .x(\c[1] ), .a(e[0]), .b(r[1]), .c(e[0]), .d(
        \c[1] ), .e(r[1]), .f(\c[1] ) );
endmodule


module chain_selement_ga_14 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_symbol_10 ( o, txack, txack_last, e, oa, r, txreq );
output [2:0] o;
input  [1:0] e;
input  [1:0] r;
input  oa, txreq;
output txack, txack_last;
    wire ack, net10, \c[0] , \c[1] ;
    chain_selement_ga_14 U1239 ( .Aa(ack), .Br(net10), .Ar(txreq), .Ba(oa) );
    and2_1 \U1229_0_/U8  ( .x(o[0]), .a(\c[0] ), .b(net10) );
    and2_1 \U1229_1_/U8  ( .x(o[1]), .a(\c[1] ), .b(net10) );
    and2_1 \U1229_2_/U8  ( .x(o[2]), .a(e[1]), .b(net10) );
    ao23_1 \U1251/U19/U21/U1/U1  ( .x(txack_last), .a(ack), .b(txack_last), 
        .c(ack), .d(e[1]), .e(e[1]) );
    ao23_1 \U1250/U19/U21/U1/U1  ( .x(txack), .a(ack), .b(txack), .c(ack), .d(
        e[0]), .e(e[0]) );
    ao222_1 \U1210/U18/U1/U1  ( .x(\c[0] ), .a(e[0]), .b(r[0]), .c(e[0]), .d(
        \c[0] ), .e(r[0]), .f(\c[0] ) );
    ao222_1 \U1209/U18/U1/U1  ( .x(\c[1] ), .a(e[0]), .b(r[1]), .c(e[0]), .d(
        \c[1] ), .e(r[1]), .f(\c[1] ) );
endmodule


module chain_selement_ga_15 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_symbol_11 ( o, txack, txack_last, e, oa, r, txreq );
output [2:0] o;
input  [1:0] e;
input  [1:0] r;
input  oa, txreq;
output txack, txack_last;
    wire ack, net10, \c[0] , \c[1] ;
    chain_selement_ga_15 U1239 ( .Aa(ack), .Br(net10), .Ar(txreq), .Ba(oa) );
    and2_1 \U1229_0_/U8  ( .x(o[0]), .a(\c[0] ), .b(net10) );
    and2_1 \U1229_1_/U8  ( .x(o[1]), .a(\c[1] ), .b(net10) );
    and2_1 \U1229_2_/U8  ( .x(o[2]), .a(e[1]), .b(net10) );
    ao23_1 \U1251/U19/U21/U1/U1  ( .x(txack_last), .a(ack), .b(txack_last), 
        .c(ack), .d(e[1]), .e(e[1]) );
    ao23_1 \U1250/U19/U21/U1/U1  ( .x(txack), .a(ack), .b(txack), .c(ack), .d(
        e[0]), .e(e[0]) );
    ao222_1 \U1210/U18/U1/U1  ( .x(\c[0] ), .a(e[0]), .b(r[0]), .c(e[0]), .d(
        \c[0] ), .e(r[0]), .f(\c[0] ) );
    ao222_1 \U1209/U18/U1/U1  ( .x(\c[1] ), .a(e[0]), .b(r[1]), .c(e[0]), .d(
        \c[1] ), .e(r[1]), .f(\c[1] ) );
endmodule


module chain_selement_ga_79 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_tx_tic ( o, rtxack, e_h, e_l, noa, r_h, r_l, rtxreq );
output [4:0] o;
input  [3:0] e_h;
input  [3:0] e_l;
input  [3:0] r_h;
input  [3:0] r_l;
input  noa, rtxreq;
output rtxack;
    wire net33, \last[4] , net60, \r3[2] , \r3[1] , \r3[0] , net40, \last[3] , 
        \r2[2] , \r2[1] , \r2[0] , net47, \last[2] , \r1[2] , \r1[1] , \r1[0] , 
        net50, \last[1] , \r0[2] , \r0[1] , \r0[0] , \last[0] , eopsym, 
        \I8/nb , \I8/na , \net55[1] , \net55[0] , \net52[1] , \net52[0] , 
        \I11/nc , \I11/nb , \I11/na , net16, net11, net9, net6, 
        \I7_0_/U25/U1/clr , \I7_0_/U25/U1/ob , \I7_1_/U25/U1/clr , 
        \I7_1_/U25/U1/ob ;
    assign o[3] = 1'b0;
    assign o[2] = 1'b0;
    route_symbol_8 I0 ( .o({\r3[2] , \r3[1] , \r3[0] }), .txack(net33), 
        .txack_last(\last[4] ), .e({e_h[3], e_l[3]}), .oa(net60), .r({r_h[3], 
        r_l[3]}), .txreq(rtxreq) );
    route_symbol_9 I1 ( .o({\r2[2] , \r2[1] , \r2[0] }), .txack(net40), 
        .txack_last(\last[3] ), .e({e_h[2], e_l[2]}), .oa(net60), .r({r_h[2], 
        r_l[2]}), .txreq(net33) );
    route_symbol_10 I2 ( .o({\r1[2] , \r1[1] , \r1[0] }), .txack(net47), 
        .txack_last(\last[2] ), .e({e_h[1], e_l[1]}), .oa(net60), .r({r_h[1], 
        r_l[1]}), .txreq(net40) );
    route_symbol_11 I3 ( .o({\r0[2] , \r0[1] , \r0[0] }), .txack(net50), 
        .txack_last(\last[1] ), .e({e_h[0], e_l[0]}), .oa(net60), .r({r_h[0], 
        r_l[0]}), .txreq(net47) );
    chain_selement_ga_79 I9 ( .Aa(\last[0] ), .Br(eopsym), .Ar(net50), .Ba(
        net60) );
    nor3_1 \I8/U27  ( .x(\I8/nb ), .a(o[4]), .b(1'b0), .c(1'b0) );
    nor2_1 \I8/U26  ( .x(\I8/na ), .a(o[1]), .b(o[0]) );
    nand2_2 \I8/U29  ( .x(net60), .a(\I8/nb ), .b(\I8/na ) );
    or2_1 \I13_0_/U12  ( .x(\net55[1] ), .a(\r1[0] ), .b(\r0[0] ) );
    or2_1 \I13_1_/U12  ( .x(\net55[0] ), .a(\r1[1] ), .b(\r0[1] ) );
    or2_1 \I14_0_/U12  ( .x(\net52[1] ), .a(\r3[0] ), .b(\r2[0] ) );
    or2_1 \I14_1_/U12  ( .x(\net52[0] ), .a(\r3[1] ), .b(\r2[1] ) );
    nand3_1 \I11/U31  ( .x(rtxack), .a(\I11/nc ), .b(\I11/nb ), .c(\I11/na )
         );
    inv_1 \I11/U33  ( .x(\I11/nc ), .a(\last[0] ) );
    nor2_1 \I11/U26  ( .x(\I11/na ), .a(\last[3] ), .b(\last[4] ) );
    nor2_1 \I11/U32  ( .x(\I11/nb ), .a(\last[1] ), .b(\last[2] ) );
    nor2_1 \I16/U5  ( .x(net16), .a(\r1[2] ), .b(\r0[2] ) );
    nor2_1 \I5/U5  ( .x(net11), .a(\r3[2] ), .b(\r2[2] ) );
    nand3_1 \I17/U9  ( .x(net9), .a(net6), .b(net11), .c(net16) );
    inv_1 \I18/U3  ( .x(net6), .a(eopsym) );
    oa31_1 \I7_0_/U25/U1/Uclr  ( .x(\I7_0_/U25/U1/clr ), .a(noa), .b(
        \net55[1] ), .c(\net52[1] ), .d(o[0]) );
    oaoi211_1 \I7_0_/U25/U1/Uaoi  ( .x(\I7_0_/U25/U1/ob ), .a(\net55[1] ), .b(
        \net52[1] ), .c(noa), .d(\I7_0_/U25/U1/clr ) );
    inv_2 \I7_0_/U25/U1/Ui  ( .x(o[0]), .a(\I7_0_/U25/U1/ob ) );
    oa31_1 \I7_1_/U25/U1/Uclr  ( .x(\I7_1_/U25/U1/clr ), .a(noa), .b(
        \net55[0] ), .c(\net52[0] ), .d(o[1]) );
    oaoi211_1 \I7_1_/U25/U1/Uaoi  ( .x(\I7_1_/U25/U1/ob ), .a(\net55[0] ), .b(
        \net52[0] ), .c(noa), .d(\I7_1_/U25/U1/clr ) );
    inv_2 \I7_1_/U25/U1/Ui  ( .x(o[1]), .a(\I7_1_/U25/U1/ob ) );
    ao222_1 \I15/U18/U1/U1  ( .x(o[4]), .a(noa), .b(net9), .c(noa), .d(o[4]), 
        .e(net9), .f(o[4]) );
endmodule


module chain_irdemuxNew_2 ( err, ncback, rd, rnw, status, cbh, cbl, nReset, 
    nack, statusack );
output [1:0] err;
output [63:0] rd;
output [1:0] rnw;
output [1:0] status;
input  [7:0] cbh;
input  [7:0] cbl;
input  nReset, nack, statusack;
output ncback;
    wire bpullcd, pullcd, net162, reset, pkt_normal, \opc_l[2] , \opc_l[1] , 
        net150, \opc_h[1] , pkt_done, write, net193, \ncd[0] , \ncd[1] , 
        \ncd[2] , \ncd[3] , \ncd[4] , \ncd[5] , \ncd[6] , \ncd[7] , 
        start_receiving, notify, net176, net86, net172, net173, net171, net169, 
        net170, net168, net166, net167, \U1664/x[3] , \U1664/U28/Z , 
        \U1664/x[0] , \U1664/U32/Z , \U1664/x[2] , \U1664/U29/Z , \U1664/y[0] , 
        \U1664/x[1] , \U1664/U33/Z , \U1664/y[1] , \U1664/U30/Z , 
        \U1664/U31/Z , \U1664/U37/Z , \U1697/U21/nr , net149, \U1697/U21/nd , 
        \U1697/U21/n2 , \U307/U21/nr , \U307/U21/nd , \U307/U21/n2 , 
        \U1698/nr , \U1698/nd , \U1698/n2 , read, n17, \opc_h[0] , n18, 
        \opc_l[0] , net0187, net0208, \I6/latch , \I6/nlocalcd , \I6/localcd , 
        \I6/ncd[0] , \I6/ncd[1] , \I6/ncd[2] , \I6/oh[2] , \I6/ncd[3] , 
        \I6/ol[3] , \I6/oh[3] , \I6/ncd[4] , \I6/ol[4] , \I6/oh[4] , 
        \I6/ncd[5] , \I6/ncd[6] , \I6/ol[6] , \I6/oh[6] , \I6/ncd[7] , 
        \I6/ol[7] , \I6/oh[7] , \I6/ctrlack_internal , \I6/acb , \I6/ba , 
        \I6/driveh , net139, \I6/drivel , n12, n13, \I6/U4/U28/U1/clr , 
        \I6/U4/U28/U1/set , \I6/U1/Z , n14, \I6/U1664/x[3] , \I6/U1664/U28/Z , 
        \I6/U1664/x[0] , \I6/U1664/U32/Z , \I6/U1664/x[2] , \I6/U1664/U29/Z , 
        \I6/U1664/y[0] , \I6/U1664/x[1] , \I6/U1664/U33/Z , \I6/U1664/y[1] , 
        \I6/U1664/U30/Z , \I6/U1664/U31/Z , \I6/U1664/U37/Z , \I6/U1669/nr , 
        \I6/U1669/nd , \I6/U1669/n2 , \U1667/latch , \U1667/nlocalcd , 
        \U1667/localcd , \U1667/ncd[0] , \U1667/ncd[1] , \U1667/ncd[2] , 
        \U1667/ncd[3] , \U1667/ncd[4] , \U1667/ncd[5] , \U1667/ncd[6] , 
        \U1667/ncd[7] , \U1667/ctrlack_internal , \U1667/acb , \U1667/ba , 
        \U1667/driveh , read_lhw, \U1667/drivel , n11, n10, 
        \U1667/U4/U28/U1/clr , \U1667/U4/U28/U1/set , \U1667/U1/Z , 
        \U1667/U1664/x[3] , \U1667/U1664/U28/Z , \U1667/U1664/x[0] , 
        \U1667/U1664/U32/Z , \U1667/U1664/x[2] , \U1667/U1664/U29/Z , 
        \U1667/U1664/y[0] , \U1667/U1664/x[1] , \U1667/U1664/U33/Z , 
        \U1667/U1664/y[1] , \U1667/U1664/U30/Z , \U1667/U1664/U31/Z , 
        \U1667/U1664/U37/Z , \U1667/U1669/nr , \U1667/U1669/nd , 
        \U1667/U1669/n2 , \U1650/latch , \U1650/nlocalcd , \U1650/localcd , 
        \U1650/ncd[0] , \U1650/ol[0] , \U1650/oh[0] , \U1650/ncd[1] , 
        \U1650/ol[1] , \U1650/oh[1] , \U1650/ncd[2] , \U1650/ol[2] , 
        \U1650/oh[2] , \U1650/ncd[3] , \U1650/ol[3] , \U1650/oh[3] , 
        \U1650/ncd[4] , \U1650/ol[4] , \U1650/oh[4] , \U1650/ncd[5] , 
        \col_l[0] , \col_h[0] , \U1650/ncd[6] , \col_l[1] , \col_h[1] , 
        \U1650/ncd[7] , \col_l[2] , \col_h[2] , \U1650/ctrlack_internal , 
        \U1650/acb , \U1650/ba , \U1650/driveh , \U1650/drivel , n7, n9, n8, 
        \U1650/U4/U28/U1/clr , \U1650/U4/U28/U1/set , \U1650/U1/Z , 
        \U1650/U1664/x[3] , \U1650/U1664/U28/Z , \U1650/U1664/x[0] , 
        \U1650/U1664/U32/Z , \U1650/U1664/x[2] , \U1650/U1664/U29/Z , 
        \U1650/U1664/y[0] , \U1650/U1664/x[1] , \U1650/U1664/U33/Z , 
        \U1650/U1664/y[1] , \U1650/U1664/U30/Z , \U1650/U1664/U31/Z , 
        \U1650/U1664/U37/Z , \U1650/U1669/nr , \U1650/U1669/nd , 
        \U1650/U1669/n2 , \U1666/latch , \U1666/nlocalcd , \U1666/localcd , 
        \U1666/ncd[0] , \U1666/ncd[1] , \U1666/ncd[2] , \U1666/ncd[3] , 
        \U1666/ncd[4] , \U1666/ncd[5] , \U1666/ncd[6] , \U1666/ncd[7] , 
        \U1666/ctrlack_internal , \U1666/acb , \U1666/ba , \U1666/driveh , 
        \U1666/drivel , n6, n5, \U1666/U4/U28/U1/clr , \U1666/U4/U28/U1/set , 
        \U1666/U1/Z , \U1666/U1664/x[3] , \U1666/U1664/U28/Z , 
        \U1666/U1664/x[0] , \U1666/U1664/U32/Z , \U1666/U1664/x[2] , 
        \U1666/U1664/U29/Z , \U1666/U1664/y[0] , \U1666/U1664/x[1] , 
        \U1666/U1664/U33/Z , \U1666/U1664/y[1] , \U1666/U1664/U30/Z , 
        \U1666/U1664/U31/Z , \U1666/U1664/U37/Z , \U1666/U1669/nr , 
        \U1666/U1669/nd , \U1666/U1669/n2 , net94, \I1/latch , \I1/nlocalcd , 
        \I1/localcd , \I1/ncd[0] , \I1/ncd[1] , \I1/ncd[2] , \I1/ncd[3] , 
        \I1/ncd[4] , \I1/ncd[5] , \I1/ncd[6] , \I1/ncd[7] , 
        \I1/ctrlack_internal , \I1/acb , \I1/ba , \I1/driveh , net103, 
        \I1/drivel , n4, n3, \I1/U4/U28/U1/clr , \I1/U4/U28/U1/set , \I1/U1/Z , 
        \I1/U1664/x[3] , \I1/U1664/U28/Z , \I1/U1664/x[0] , \I1/U1664/U32/Z , 
        \I1/U1664/x[2] , \I1/U1664/U29/Z , \I1/U1664/y[0] , \I1/U1664/x[1] , 
        \I1/U1664/U33/Z , \I1/U1664/y[1] , \I1/U1664/U30/Z , \I1/U1664/U31/Z , 
        \I1/U1664/U37/Z , \I1/U1669/nr , \I1/U1669/nd , \I1/U1669/n2 , 
        \I2/latch , \I2/nlocalcd , \I2/localcd , \I2/ncd[0] , \I2/ncd[1] , 
        \I2/ncd[2] , \I2/ncd[3] , \I2/ncd[4] , \I2/ncd[5] , \I2/ncd[6] , 
        \I2/ncd[7] , \I2/ctrlack_internal , \I2/acb , \I2/ba , \I2/driveh , 
        \I2/drivel , n2, n1, \I2/U4/U28/U1/clr , \I2/U4/U28/U1/set , \I2/U1/Z , 
        \I2/U1664/x[3] , \I2/U1664/U28/Z , \I2/U1664/x[0] , \I2/U1664/U32/Z , 
        \I2/U1664/x[2] , \I2/U1664/U29/Z , \I2/U1664/y[0] , \I2/U1664/x[1] , 
        \I2/U1664/U33/Z , \I2/U1664/y[1] , \I2/U1664/U30/Z , \I2/U1664/U31/Z , 
        \I2/U1664/U37/Z , \I2/U1669/nr , \I2/U1669/nd , \I2/U1669/n2 ;
    buf_1 U262 ( .x(bpullcd), .a(pullcd) );
    or2_4 \U1674/U12  ( .x(net162), .a(nack), .b(reset) );
    and2_4 \U1785/U8  ( .x(pkt_normal), .a(\opc_l[2] ), .b(\opc_l[1] ) );
    and2_4 \U1777/U8  ( .x(net150), .a(\opc_l[2] ), .b(\opc_h[1] ) );
    or3_1 \U1813/U12  ( .x(pkt_done), .a(write), .b(reset), .c(net193) );
    nor2_1 \U1651_0_/U5  ( .x(\ncd[0] ), .a(cbh[0]), .b(cbl[0]) );
    nor2_1 \U1651_1_/U5  ( .x(\ncd[1] ), .a(cbh[1]), .b(cbl[1]) );
    nor2_1 \U1651_2_/U5  ( .x(\ncd[2] ), .a(cbh[2]), .b(cbl[2]) );
    nor2_1 \U1651_3_/U5  ( .x(\ncd[3] ), .a(cbh[3]), .b(cbl[3]) );
    nor2_1 \U1651_4_/U5  ( .x(\ncd[4] ), .a(cbh[4]), .b(cbl[4]) );
    nor2_1 \U1651_5_/U5  ( .x(\ncd[5] ), .a(cbh[5]), .b(cbl[5]) );
    nor2_1 \U1651_6_/U5  ( .x(\ncd[6] ), .a(cbh[6]), .b(cbl[6]) );
    nor2_1 \U1651_7_/U5  ( .x(\ncd[7] ), .a(cbh[7]), .b(cbl[7]) );
    nor2_1 \U1812/U5  ( .x(start_receiving), .a(notify), .b(net176) );
    nor2_1 \I7/U5  ( .x(net86), .a(net172), .b(net173) );
    nor2_1 \I4/U5  ( .x(net171), .a(net169), .b(net170) );
    nor2_1 \I3/U5  ( .x(net168), .a(net166), .b(net167) );
    inv_2 \U1675/U3  ( .x(reset), .a(nReset) );
    nand3_2 \U193/U16  ( .x(ncback), .a(net86), .b(net171), .c(net168) );
    ao222_1 \U1811/U18/U1/U1  ( .x(net176), .a(net162), .b(pkt_done), .c(
        net162), .d(net176), .e(pkt_done), .f(net176) );
    aoi222_1 \U1664/U28/U30/U1  ( .x(\U1664/x[3] ), .a(\ncd[7] ), .b(\ncd[6] ), 
        .c(\ncd[7] ), .d(\U1664/U28/Z ), .e(\ncd[6] ), .f(\U1664/U28/Z ) );
    inv_1 \U1664/U28/U30/Uinv  ( .x(\U1664/U28/Z ), .a(\U1664/x[3] ) );
    aoi222_1 \U1664/U32/U30/U1  ( .x(\U1664/x[0] ), .a(\ncd[1] ), .b(\ncd[0] ), 
        .c(\ncd[1] ), .d(\U1664/U32/Z ), .e(\ncd[0] ), .f(\U1664/U32/Z ) );
    inv_1 \U1664/U32/U30/Uinv  ( .x(\U1664/U32/Z ), .a(\U1664/x[0] ) );
    aoi222_1 \U1664/U29/U30/U1  ( .x(\U1664/x[2] ), .a(\ncd[5] ), .b(\ncd[4] ), 
        .c(\ncd[5] ), .d(\U1664/U29/Z ), .e(\ncd[4] ), .f(\U1664/U29/Z ) );
    inv_1 \U1664/U29/U30/Uinv  ( .x(\U1664/U29/Z ), .a(\U1664/x[2] ) );
    aoi222_1 \U1664/U33/U30/U1  ( .x(\U1664/y[0] ), .a(\U1664/x[1] ), .b(
        \U1664/x[0] ), .c(\U1664/x[1] ), .d(\U1664/U33/Z ), .e(\U1664/x[0] ), 
        .f(\U1664/U33/Z ) );
    inv_1 \U1664/U33/U30/Uinv  ( .x(\U1664/U33/Z ), .a(\U1664/y[0] ) );
    aoi222_1 \U1664/U30/U30/U1  ( .x(\U1664/y[1] ), .a(\U1664/x[3] ), .b(
        \U1664/x[2] ), .c(\U1664/x[3] ), .d(\U1664/U30/Z ), .e(\U1664/x[2] ), 
        .f(\U1664/U30/Z ) );
    inv_1 \U1664/U30/U30/Uinv  ( .x(\U1664/U30/Z ), .a(\U1664/y[1] ) );
    aoi222_1 \U1664/U31/U30/U1  ( .x(\U1664/x[1] ), .a(\ncd[3] ), .b(\ncd[2] ), 
        .c(\ncd[3] ), .d(\U1664/U31/Z ), .e(\ncd[2] ), .f(\U1664/U31/Z ) );
    inv_1 \U1664/U31/U30/Uinv  ( .x(\U1664/U31/Z ), .a(\U1664/x[1] ) );
    aoi222_1 \U1664/U37/U30/U1  ( .x(pullcd), .a(\U1664/y[0] ), .b(
        \U1664/y[1] ), .c(\U1664/y[0] ), .d(\U1664/U37/Z ), .e(\U1664/y[1] ), 
        .f(\U1664/U37/Z ) );
    inv_1 \U1664/U37/U30/Uinv  ( .x(\U1664/U37/Z ), .a(pullcd) );
    nor3_1 \U1697/U21/Unr  ( .x(\U1697/U21/nr ), .a(rnw[0]), .b(pkt_normal), 
        .c(net149) );
    nand3_1 \U1697/U21/Und  ( .x(\U1697/U21/nd ), .a(rnw[0]), .b(pkt_normal), 
        .c(net149) );
    oa21_1 \U1697/U21/U1  ( .x(\U1697/U21/n2 ), .a(\U1697/U21/n2 ), .b(
        \U1697/U21/nr ), .c(\U1697/U21/nd ) );
    inv_1 \U1697/U21/U3  ( .x(write), .a(\U1697/U21/n2 ) );
    nor3_1 \U307/U21/Unr  ( .x(\U307/U21/nr ), .a(net149), .b(net150), .c(
        statusack) );
    nand3_1 \U307/U21/Und  ( .x(\U307/U21/nd ), .a(net149), .b(net150), .c(
        statusack) );
    oa21_1 \U307/U21/U1  ( .x(\U307/U21/n2 ), .a(\U307/U21/n2 ), .b(
        \U307/U21/nr ), .c(\U307/U21/nd ) );
    inv_1 \U307/U21/U3  ( .x(notify), .a(\U307/U21/n2 ) );
    nor3_1 \U1698/Unr  ( .x(\U1698/nr ), .a(rnw[1]), .b(pkt_normal), .c(net149
        ) );
    nand3_1 \U1698/Und  ( .x(\U1698/nd ), .a(rnw[1]), .b(pkt_normal), .c(
        net149) );
    oa21_1 \U1698/U1  ( .x(\U1698/n2 ), .a(\U1698/n2 ), .b(\U1698/nr ), .c(
        \U1698/nd ) );
    inv_2 \U1698/U3  ( .x(read), .a(\U1698/n2 ) );
    and2_1 \U1756/U1754/U8  ( .x(n17), .a(\opc_h[0] ), .b(pkt_normal) );
    and2_1 \U1756/U1755/U8  ( .x(n18), .a(\opc_l[0] ), .b(pkt_normal) );
    and2_1 \U1800/U1754/U8  ( .x(rnw[1]), .a(net0187), .b(pkt_normal) );
    and2_1 \U1800/U1755/U8  ( .x(rnw[0]), .a(net0208), .b(pkt_normal) );
    and2_1 \U1758/U1754/U8  ( .x(status[1]), .a(\opc_h[0] ), .b(net150) );
    and2_1 \U1758/U1755/U8  ( .x(status[0]), .a(\opc_l[0] ), .b(net150) );
    buf_2 \I6/U1653  ( .x(\I6/latch ), .a(net173) );
    nor2_1 \I6/U264/U5  ( .x(\I6/nlocalcd ), .a(reset), .b(\I6/localcd ) );
    nor2_1 \I6/U1659_0_/U5  ( .x(\I6/ncd[0] ), .a(\opc_l[0] ), .b(\opc_h[0] )
         );
    nor2_1 \I6/U1659_1_/U5  ( .x(\I6/ncd[1] ), .a(\opc_l[1] ), .b(\opc_h[1] )
         );
    nor2_1 \I6/U1659_2_/U5  ( .x(\I6/ncd[2] ), .a(\opc_l[2] ), .b(\I6/oh[2] )
         );
    nor2_1 \I6/U1659_3_/U5  ( .x(\I6/ncd[3] ), .a(\I6/ol[3] ), .b(\I6/oh[3] )
         );
    nor2_1 \I6/U1659_4_/U5  ( .x(\I6/ncd[4] ), .a(\I6/ol[4] ), .b(\I6/oh[4] )
         );
    nor2_1 \I6/U1659_5_/U5  ( .x(\I6/ncd[5] ), .a(net0208), .b(net0187) );
    nor2_1 \I6/U1659_6_/U5  ( .x(\I6/ncd[6] ), .a(\I6/ol[6] ), .b(\I6/oh[6] )
         );
    nor2_1 \I6/U1659_7_/U5  ( .x(\I6/ncd[7] ), .a(\I6/ol[7] ), .b(\I6/oh[7] )
         );
    nor2_1 \I6/U3/U5  ( .x(\I6/ctrlack_internal ), .a(\I6/acb ), .b(\I6/ba )
         );
    buf_2 \I6/U1665/U7  ( .x(\I6/driveh ), .a(net139) );
    buf_2 \I6/U1666/U7  ( .x(\I6/drivel ), .a(net139) );
    ao23_1 \I6/U1658_0_/U21/U1/U1  ( .x(\opc_l[0] ), .a(\I6/driveh ), .b(
        \opc_l[0] ), .c(\I6/driveh ), .d(cbl[0]), .e(n12) );
    ao23_1 \I6/U1658_1_/U21/U1/U1  ( .x(\opc_l[1] ), .a(\I6/driveh ), .b(
        \opc_l[1] ), .c(\I6/drivel ), .d(cbl[1]), .e(n12) );
    ao23_1 \I6/U1658_2_/U21/U1/U1  ( .x(\opc_l[2] ), .a(\I6/drivel ), .b(
        \opc_l[2] ), .c(n13), .d(cbl[2]), .e(n12) );
    ao23_1 \I6/U1658_3_/U21/U1/U1  ( .x(\I6/ol[3] ), .a(\I6/drivel ), .b(
        \I6/ol[3] ), .c(\I6/drivel ), .d(cbl[3]), .e(\I6/latch ) );
    ao23_1 \I6/U1658_4_/U21/U1/U1  ( .x(\I6/ol[4] ), .a(n13), .b(\I6/ol[4] ), 
        .c(n13), .d(cbl[4]), .e(\I6/latch ) );
    ao23_1 \I6/U1658_5_/U21/U1/U1  ( .x(net0208), .a(\I6/driveh ), .b(net0208), 
        .c(\I6/driveh ), .d(cbl[5]), .e(\I6/latch ) );
    ao23_1 \I6/U1658_6_/U21/U1/U1  ( .x(\I6/ol[6] ), .a(n13), .b(\I6/ol[6] ), 
        .c(n13), .d(cbl[6]), .e(\I6/latch ) );
    ao23_1 \I6/U1658_7_/U21/U1/U1  ( .x(\I6/ol[7] ), .a(n13), .b(\I6/ol[7] ), 
        .c(\I6/driveh ), .d(cbl[7]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_0_/U21/U1/U1  ( .x(\opc_h[0] ), .a(n13), .b(\opc_h[0] ), 
        .c(\I6/drivel ), .d(cbh[0]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_1_/U21/U1/U1  ( .x(\opc_h[1] ), .a(\I6/driveh ), .b(
        \opc_h[1] ), .c(n13), .d(cbh[1]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_2_/U21/U1/U1  ( .x(\I6/oh[2] ), .a(\I6/driveh ), .b(
        \I6/oh[2] ), .c(n13), .d(cbh[2]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_3_/U21/U1/U1  ( .x(\I6/oh[3] ), .a(\I6/drivel ), .b(
        \I6/oh[3] ), .c(\I6/drivel ), .d(cbh[3]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_4_/U21/U1/U1  ( .x(\I6/oh[4] ), .a(n13), .b(\I6/oh[4] ), 
        .c(\I6/driveh ), .d(cbh[4]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_5_/U21/U1/U1  ( .x(net0187), .a(\I6/driveh ), .b(net0187), 
        .c(\I6/driveh ), .d(cbh[5]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_6_/U21/U1/U1  ( .x(\I6/oh[6] ), .a(\I6/drivel ), .b(
        \I6/oh[6] ), .c(\I6/drivel ), .d(cbh[6]), .e(\I6/latch ) );
    ao23_1 \I6/U1651_7_/U21/U1/U1  ( .x(\I6/oh[7] ), .a(\I6/drivel ), .b(
        \I6/oh[7] ), .c(n13), .d(cbh[7]), .e(\I6/latch ) );
    aoai211_1 \I6/U4/U28/U1/U1  ( .x(\I6/U4/U28/U1/clr ), .a(net139), .b(
        \I6/acb ), .c(\I6/nlocalcd ), .d(net173) );
    nand3_1 \I6/U4/U28/U1/U2  ( .x(\I6/U4/U28/U1/set ), .a(\I6/nlocalcd ), .b(
        net139), .c(\I6/acb ) );
    nand2_2 \I6/U4/U28/U1/U3  ( .x(net173), .a(\I6/U4/U28/U1/clr ), .b(
        \I6/U4/U28/U1/set ) );
    oai21_1 \I6/U1/U30/U1/U1  ( .x(\I6/acb ), .a(\I6/U1/Z ), .b(\I6/ba ), .c(
        net139) );
    inv_1 \I6/U1/U30/U1/U2  ( .x(\I6/U1/Z ), .a(\I6/acb ) );
    ao222_1 \I6/U5/U18/U1/U1  ( .x(\I6/ba ), .a(\I6/latch ), .b(n14), .c(
        \I6/latch ), .d(\I6/ba ), .e(n14), .f(\I6/ba ) );
    aoi222_1 \I6/U1664/U28/U30/U1  ( .x(\I6/U1664/x[3] ), .a(\I6/ncd[7] ), .b(
        \I6/ncd[6] ), .c(\I6/ncd[7] ), .d(\I6/U1664/U28/Z ), .e(\I6/ncd[6] ), 
        .f(\I6/U1664/U28/Z ) );
    inv_1 \I6/U1664/U28/U30/Uinv  ( .x(\I6/U1664/U28/Z ), .a(\I6/U1664/x[3] )
         );
    aoi222_1 \I6/U1664/U32/U30/U1  ( .x(\I6/U1664/x[0] ), .a(\I6/ncd[1] ), .b(
        \I6/ncd[0] ), .c(\I6/ncd[1] ), .d(\I6/U1664/U32/Z ), .e(\I6/ncd[0] ), 
        .f(\I6/U1664/U32/Z ) );
    inv_1 \I6/U1664/U32/U30/Uinv  ( .x(\I6/U1664/U32/Z ), .a(\I6/U1664/x[0] )
         );
    aoi222_1 \I6/U1664/U29/U30/U1  ( .x(\I6/U1664/x[2] ), .a(\I6/ncd[5] ), .b(
        \I6/ncd[4] ), .c(\I6/ncd[5] ), .d(\I6/U1664/U29/Z ), .e(\I6/ncd[4] ), 
        .f(\I6/U1664/U29/Z ) );
    inv_1 \I6/U1664/U29/U30/Uinv  ( .x(\I6/U1664/U29/Z ), .a(\I6/U1664/x[2] )
         );
    aoi222_1 \I6/U1664/U33/U30/U1  ( .x(\I6/U1664/y[0] ), .a(\I6/U1664/x[1] ), 
        .b(\I6/U1664/x[0] ), .c(\I6/U1664/x[1] ), .d(\I6/U1664/U33/Z ), .e(
        \I6/U1664/x[0] ), .f(\I6/U1664/U33/Z ) );
    inv_1 \I6/U1664/U33/U30/Uinv  ( .x(\I6/U1664/U33/Z ), .a(\I6/U1664/y[0] )
         );
    aoi222_1 \I6/U1664/U30/U30/U1  ( .x(\I6/U1664/y[1] ), .a(\I6/U1664/x[3] ), 
        .b(\I6/U1664/x[2] ), .c(\I6/U1664/x[3] ), .d(\I6/U1664/U30/Z ), .e(
        \I6/U1664/x[2] ), .f(\I6/U1664/U30/Z ) );
    inv_1 \I6/U1664/U30/U30/Uinv  ( .x(\I6/U1664/U30/Z ), .a(\I6/U1664/y[1] )
         );
    aoi222_1 \I6/U1664/U31/U30/U1  ( .x(\I6/U1664/x[1] ), .a(\I6/ncd[3] ), .b(
        \I6/ncd[2] ), .c(\I6/ncd[3] ), .d(\I6/U1664/U31/Z ), .e(\I6/ncd[2] ), 
        .f(\I6/U1664/U31/Z ) );
    inv_1 \I6/U1664/U31/U30/Uinv  ( .x(\I6/U1664/U31/Z ), .a(\I6/U1664/x[1] )
         );
    aoi222_1 \I6/U1664/U37/U30/U1  ( .x(\I6/localcd ), .a(\I6/U1664/y[0] ), 
        .b(\I6/U1664/y[1] ), .c(\I6/U1664/y[0] ), .d(\I6/U1664/U37/Z ), .e(
        \I6/U1664/y[1] ), .f(\I6/U1664/U37/Z ) );
    inv_1 \I6/U1664/U37/U30/Uinv  ( .x(\I6/U1664/U37/Z ), .a(\I6/localcd ) );
    nor3_1 \I6/U1669/Unr  ( .x(\I6/U1669/nr ), .a(\I6/ctrlack_internal ), .b(
        n13), .c(\I6/drivel ) );
    nand3_1 \I6/U1669/Und  ( .x(\I6/U1669/nd ), .a(\I6/ctrlack_internal ), .b(
        \I6/driveh ), .c(\I6/drivel ) );
    oa21_1 \I6/U1669/U1  ( .x(\I6/U1669/n2 ), .a(\I6/U1669/n2 ), .b(
        \I6/U1669/nr ), .c(\I6/U1669/nd ) );
    inv_2 \I6/U1669/U3  ( .x(net149), .a(\I6/U1669/n2 ) );
    buf_2 \U1667/U1653  ( .x(\U1667/latch ), .a(net167) );
    nor2_1 \U1667/U264/U5  ( .x(\U1667/nlocalcd ), .a(reset), .b(
        \U1667/localcd ) );
    nor2_1 \U1667/U1659_0_/U5  ( .x(\U1667/ncd[0] ), .a(rd[0]), .b(rd[32]) );
    nor2_1 \U1667/U1659_1_/U5  ( .x(\U1667/ncd[1] ), .a(rd[1]), .b(rd[33]) );
    nor2_1 \U1667/U1659_2_/U5  ( .x(\U1667/ncd[2] ), .a(rd[2]), .b(rd[34]) );
    nor2_1 \U1667/U1659_3_/U5  ( .x(\U1667/ncd[3] ), .a(rd[3]), .b(rd[35]) );
    nor2_1 \U1667/U1659_4_/U5  ( .x(\U1667/ncd[4] ), .a(rd[4]), .b(rd[36]) );
    nor2_1 \U1667/U1659_5_/U5  ( .x(\U1667/ncd[5] ), .a(rd[5]), .b(rd[37]) );
    nor2_1 \U1667/U1659_6_/U5  ( .x(\U1667/ncd[6] ), .a(rd[6]), .b(rd[38]) );
    nor2_1 \U1667/U1659_7_/U5  ( .x(\U1667/ncd[7] ), .a(rd[7]), .b(rd[39]) );
    nor2_1 \U1667/U3/U5  ( .x(\U1667/ctrlack_internal ), .a(\U1667/acb ), .b(
        \U1667/ba ) );
    buf_2 \U1667/U1665/U7  ( .x(\U1667/driveh ), .a(read_lhw) );
    buf_2 \U1667/U1666/U7  ( .x(\U1667/drivel ), .a(read_lhw) );
    ao23_1 \U1667/U1658_0_/U21/U1/U1  ( .x(rd[0]), .a(n11), .b(rd[0]), .c(
        \U1667/drivel ), .d(cbl[0]), .e(n10) );
    ao23_1 \U1667/U1658_1_/U21/U1/U1  ( .x(rd[1]), .a(n11), .b(rd[1]), .c(
        \U1667/driveh ), .d(cbl[1]), .e(n10) );
    ao23_1 \U1667/U1658_2_/U21/U1/U1  ( .x(rd[2]), .a(\U1667/driveh ), .b(rd
        [2]), .c(n11), .d(cbl[2]), .e(n10) );
    ao23_1 \U1667/U1658_3_/U21/U1/U1  ( .x(rd[3]), .a(n11), .b(rd[3]), .c(
        \U1667/driveh ), .d(cbl[3]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1658_4_/U21/U1/U1  ( .x(rd[4]), .a(\U1667/drivel ), .b(rd
        [4]), .c(n11), .d(cbl[4]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1658_5_/U21/U1/U1  ( .x(rd[5]), .a(\U1667/drivel ), .b(rd
        [5]), .c(n11), .d(cbl[5]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1658_6_/U21/U1/U1  ( .x(rd[6]), .a(\U1667/driveh ), .b(rd
        [6]), .c(\U1667/drivel ), .d(cbl[6]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1658_7_/U21/U1/U1  ( .x(rd[7]), .a(\U1667/driveh ), .b(rd
        [7]), .c(\U1667/driveh ), .d(cbl[7]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_0_/U21/U1/U1  ( .x(rd[32]), .a(\U1667/drivel ), .b(rd
        [32]), .c(n11), .d(cbh[0]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_1_/U21/U1/U1  ( .x(rd[33]), .a(\U1667/driveh ), .b(rd
        [33]), .c(\U1667/drivel ), .d(cbh[1]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_2_/U21/U1/U1  ( .x(rd[34]), .a(\U1667/drivel ), .b(rd
        [34]), .c(\U1667/drivel ), .d(cbh[2]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_3_/U21/U1/U1  ( .x(rd[35]), .a(\U1667/driveh ), .b(rd
        [35]), .c(\U1667/driveh ), .d(cbh[3]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_4_/U21/U1/U1  ( .x(rd[36]), .a(\U1667/drivel ), .b(rd
        [36]), .c(\U1667/driveh ), .d(cbh[4]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_5_/U21/U1/U1  ( .x(rd[37]), .a(\U1667/driveh ), .b(rd
        [37]), .c(n11), .d(cbh[5]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_6_/U21/U1/U1  ( .x(rd[38]), .a(n11), .b(rd[38]), .c(
        \U1667/drivel ), .d(cbh[6]), .e(\U1667/latch ) );
    ao23_1 \U1667/U1651_7_/U21/U1/U1  ( .x(rd[39]), .a(n11), .b(rd[39]), .c(
        n11), .d(cbh[7]), .e(\U1667/latch ) );
    aoai211_1 \U1667/U4/U28/U1/U1  ( .x(\U1667/U4/U28/U1/clr ), .a(read_lhw), 
        .b(\U1667/acb ), .c(\U1667/nlocalcd ), .d(net167) );
    nand3_1 \U1667/U4/U28/U1/U2  ( .x(\U1667/U4/U28/U1/set ), .a(
        \U1667/nlocalcd ), .b(read_lhw), .c(\U1667/acb ) );
    nand2_2 \U1667/U4/U28/U1/U3  ( .x(net167), .a(\U1667/U4/U28/U1/clr ), .b(
        \U1667/U4/U28/U1/set ) );
    oai21_1 \U1667/U1/U30/U1/U1  ( .x(\U1667/acb ), .a(\U1667/U1/Z ), .b(
        \U1667/ba ), .c(read_lhw) );
    inv_1 \U1667/U1/U30/U1/U2  ( .x(\U1667/U1/Z ), .a(\U1667/acb ) );
    ao222_1 \U1667/U5/U18/U1/U1  ( .x(\U1667/ba ), .a(\U1667/latch ), .b(n14), 
        .c(\U1667/latch ), .d(\U1667/ba ), .e(n14), .f(\U1667/ba ) );
    aoi222_1 \U1667/U1664/U28/U30/U1  ( .x(\U1667/U1664/x[3] ), .a(
        \U1667/ncd[7] ), .b(\U1667/ncd[6] ), .c(\U1667/ncd[7] ), .d(
        \U1667/U1664/U28/Z ), .e(\U1667/ncd[6] ), .f(\U1667/U1664/U28/Z ) );
    inv_1 \U1667/U1664/U28/U30/Uinv  ( .x(\U1667/U1664/U28/Z ), .a(
        \U1667/U1664/x[3] ) );
    aoi222_1 \U1667/U1664/U32/U30/U1  ( .x(\U1667/U1664/x[0] ), .a(
        \U1667/ncd[1] ), .b(\U1667/ncd[0] ), .c(\U1667/ncd[1] ), .d(
        \U1667/U1664/U32/Z ), .e(\U1667/ncd[0] ), .f(\U1667/U1664/U32/Z ) );
    inv_1 \U1667/U1664/U32/U30/Uinv  ( .x(\U1667/U1664/U32/Z ), .a(
        \U1667/U1664/x[0] ) );
    aoi222_1 \U1667/U1664/U29/U30/U1  ( .x(\U1667/U1664/x[2] ), .a(
        \U1667/ncd[5] ), .b(\U1667/ncd[4] ), .c(\U1667/ncd[5] ), .d(
        \U1667/U1664/U29/Z ), .e(\U1667/ncd[4] ), .f(\U1667/U1664/U29/Z ) );
    inv_1 \U1667/U1664/U29/U30/Uinv  ( .x(\U1667/U1664/U29/Z ), .a(
        \U1667/U1664/x[2] ) );
    aoi222_1 \U1667/U1664/U33/U30/U1  ( .x(\U1667/U1664/y[0] ), .a(
        \U1667/U1664/x[1] ), .b(\U1667/U1664/x[0] ), .c(\U1667/U1664/x[1] ), 
        .d(\U1667/U1664/U33/Z ), .e(\U1667/U1664/x[0] ), .f(
        \U1667/U1664/U33/Z ) );
    inv_1 \U1667/U1664/U33/U30/Uinv  ( .x(\U1667/U1664/U33/Z ), .a(
        \U1667/U1664/y[0] ) );
    aoi222_1 \U1667/U1664/U30/U30/U1  ( .x(\U1667/U1664/y[1] ), .a(
        \U1667/U1664/x[3] ), .b(\U1667/U1664/x[2] ), .c(\U1667/U1664/x[3] ), 
        .d(\U1667/U1664/U30/Z ), .e(\U1667/U1664/x[2] ), .f(
        \U1667/U1664/U30/Z ) );
    inv_1 \U1667/U1664/U30/U30/Uinv  ( .x(\U1667/U1664/U30/Z ), .a(
        \U1667/U1664/y[1] ) );
    aoi222_1 \U1667/U1664/U31/U30/U1  ( .x(\U1667/U1664/x[1] ), .a(
        \U1667/ncd[3] ), .b(\U1667/ncd[2] ), .c(\U1667/ncd[3] ), .d(
        \U1667/U1664/U31/Z ), .e(\U1667/ncd[2] ), .f(\U1667/U1664/U31/Z ) );
    inv_1 \U1667/U1664/U31/U30/Uinv  ( .x(\U1667/U1664/U31/Z ), .a(
        \U1667/U1664/x[1] ) );
    aoi222_1 \U1667/U1664/U37/U30/U1  ( .x(\U1667/localcd ), .a(
        \U1667/U1664/y[0] ), .b(\U1667/U1664/y[1] ), .c(\U1667/U1664/y[0] ), 
        .d(\U1667/U1664/U37/Z ), .e(\U1667/U1664/y[1] ), .f(
        \U1667/U1664/U37/Z ) );
    inv_1 \U1667/U1664/U37/U30/Uinv  ( .x(\U1667/U1664/U37/Z ), .a(
        \U1667/localcd ) );
    nor3_1 \U1667/U1669/Unr  ( .x(\U1667/U1669/nr ), .a(
        \U1667/ctrlack_internal ), .b(n11), .c(\U1667/drivel ) );
    nand3_1 \U1667/U1669/Und  ( .x(\U1667/U1669/nd ), .a(
        \U1667/ctrlack_internal ), .b(\U1667/driveh ), .c(\U1667/drivel ) );
    oa21_1 \U1667/U1669/U1  ( .x(\U1667/U1669/n2 ), .a(\U1667/U1669/n2 ), .b(
        \U1667/U1669/nr ), .c(\U1667/U1669/nd ) );
    inv_2 \U1667/U1669/U3  ( .x(net193), .a(\U1667/U1669/n2 ) );
    buf_2 \U1650/U1653  ( .x(\U1650/latch ), .a(net172) );
    nor2_1 \U1650/U264/U5  ( .x(\U1650/nlocalcd ), .a(reset), .b(
        \U1650/localcd ) );
    nor2_1 \U1650/U1659_0_/U5  ( .x(\U1650/ncd[0] ), .a(\U1650/ol[0] ), .b(
        \U1650/oh[0] ) );
    nor2_1 \U1650/U1659_1_/U5  ( .x(\U1650/ncd[1] ), .a(\U1650/ol[1] ), .b(
        \U1650/oh[1] ) );
    nor2_1 \U1650/U1659_2_/U5  ( .x(\U1650/ncd[2] ), .a(\U1650/ol[2] ), .b(
        \U1650/oh[2] ) );
    nor2_1 \U1650/U1659_3_/U5  ( .x(\U1650/ncd[3] ), .a(\U1650/ol[3] ), .b(
        \U1650/oh[3] ) );
    nor2_1 \U1650/U1659_4_/U5  ( .x(\U1650/ncd[4] ), .a(\U1650/ol[4] ), .b(
        \U1650/oh[4] ) );
    nor2_1 \U1650/U1659_5_/U5  ( .x(\U1650/ncd[5] ), .a(\col_l[0] ), .b(
        \col_h[0] ) );
    nor2_1 \U1650/U1659_6_/U5  ( .x(\U1650/ncd[6] ), .a(\col_l[1] ), .b(
        \col_h[1] ) );
    nor2_1 \U1650/U1659_7_/U5  ( .x(\U1650/ncd[7] ), .a(\col_l[2] ), .b(
        \col_h[2] ) );
    nor2_1 \U1650/U3/U5  ( .x(\U1650/ctrlack_internal ), .a(\U1650/acb ), .b(
        \U1650/ba ) );
    buf_2 \U1650/U1665/U7  ( .x(\U1650/driveh ), .a(start_receiving) );
    buf_2 \U1650/U1666/U7  ( .x(\U1650/drivel ), .a(start_receiving) );
    ao23_1 \U1650/U1658_0_/U21/U1/U1  ( .x(\U1650/ol[0] ), .a(\U1650/drivel ), 
        .b(\U1650/ol[0] ), .c(\U1650/drivel ), .d(cbl[0]), .e(n7) );
    ao23_1 \U1650/U1658_1_/U21/U1/U1  ( .x(\U1650/ol[1] ), .a(\U1650/drivel ), 
        .b(\U1650/ol[1] ), .c(\U1650/drivel ), .d(cbl[1]), .e(n7) );
    ao23_1 \U1650/U1658_2_/U21/U1/U1  ( .x(\U1650/ol[2] ), .a(\U1650/drivel ), 
        .b(\U1650/ol[2] ), .c(\U1650/drivel ), .d(cbl[2]), .e(n7) );
    ao23_1 \U1650/U1658_3_/U21/U1/U1  ( .x(\U1650/ol[3] ), .a(n9), .b(
        \U1650/ol[3] ), .c(\U1650/drivel ), .d(cbl[3]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1658_4_/U21/U1/U1  ( .x(\U1650/ol[4] ), .a(\U1650/drivel ), 
        .b(\U1650/ol[4] ), .c(\U1650/drivel ), .d(cbl[4]), .e(\U1650/latch )
         );
    ao23_1 \U1650/U1658_5_/U21/U1/U1  ( .x(\col_l[0] ), .a(\U1650/drivel ), 
        .b(\col_l[0] ), .c(\U1650/drivel ), .d(cbl[5]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1658_6_/U21/U1/U1  ( .x(\col_l[1] ), .a(n9), .b(\col_l[1] ), 
        .c(\U1650/drivel ), .d(cbl[6]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1658_7_/U21/U1/U1  ( .x(\col_l[2] ), .a(n9), .b(\col_l[2] ), 
        .c(\U1650/drivel ), .d(cbl[7]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1651_0_/U21/U1/U1  ( .x(\U1650/oh[0] ), .a(\U1650/driveh ), 
        .b(\U1650/oh[0] ), .c(\U1650/driveh ), .d(cbh[0]), .e(\U1650/latch )
         );
    ao23_1 \U1650/U1651_1_/U21/U1/U1  ( .x(\U1650/oh[1] ), .a(\U1650/driveh ), 
        .b(\U1650/oh[1] ), .c(\U1650/driveh ), .d(cbh[1]), .e(\U1650/latch )
         );
    ao23_1 \U1650/U1651_2_/U21/U1/U1  ( .x(\U1650/oh[2] ), .a(\U1650/driveh ), 
        .b(\U1650/oh[2] ), .c(\U1650/driveh ), .d(cbh[2]), .e(\U1650/latch )
         );
    ao23_1 \U1650/U1651_3_/U21/U1/U1  ( .x(\U1650/oh[3] ), .a(n8), .b(
        \U1650/oh[3] ), .c(\U1650/driveh ), .d(cbh[3]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1651_4_/U21/U1/U1  ( .x(\U1650/oh[4] ), .a(n8), .b(
        \U1650/oh[4] ), .c(\U1650/driveh ), .d(cbh[4]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1651_5_/U21/U1/U1  ( .x(\col_h[0] ), .a(\U1650/driveh ), 
        .b(\col_h[0] ), .c(\U1650/driveh ), .d(cbh[5]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1651_6_/U21/U1/U1  ( .x(\col_h[1] ), .a(n8), .b(\col_h[1] ), 
        .c(\U1650/driveh ), .d(cbh[6]), .e(\U1650/latch ) );
    ao23_1 \U1650/U1651_7_/U21/U1/U1  ( .x(\col_h[2] ), .a(\U1650/driveh ), 
        .b(\col_h[2] ), .c(\U1650/driveh ), .d(cbh[7]), .e(\U1650/latch ) );
    aoai211_1 \U1650/U4/U28/U1/U1  ( .x(\U1650/U4/U28/U1/clr ), .a(
        start_receiving), .b(\U1650/acb ), .c(\U1650/nlocalcd ), .d(net172) );
    nand3_1 \U1650/U4/U28/U1/U2  ( .x(\U1650/U4/U28/U1/set ), .a(
        \U1650/nlocalcd ), .b(start_receiving), .c(\U1650/acb ) );
    nand2_2 \U1650/U4/U28/U1/U3  ( .x(net172), .a(\U1650/U4/U28/U1/clr ), .b(
        \U1650/U4/U28/U1/set ) );
    oai21_1 \U1650/U1/U30/U1/U1  ( .x(\U1650/acb ), .a(\U1650/U1/Z ), .b(
        \U1650/ba ), .c(start_receiving) );
    inv_1 \U1650/U1/U30/U1/U2  ( .x(\U1650/U1/Z ), .a(\U1650/acb ) );
    ao222_1 \U1650/U5/U18/U1/U1  ( .x(\U1650/ba ), .a(\U1650/latch ), .b(n14), 
        .c(\U1650/latch ), .d(\U1650/ba ), .e(n14), .f(\U1650/ba ) );
    aoi222_1 \U1650/U1664/U28/U30/U1  ( .x(\U1650/U1664/x[3] ), .a(
        \U1650/ncd[7] ), .b(\U1650/ncd[6] ), .c(\U1650/ncd[7] ), .d(
        \U1650/U1664/U28/Z ), .e(\U1650/ncd[6] ), .f(\U1650/U1664/U28/Z ) );
    inv_1 \U1650/U1664/U28/U30/Uinv  ( .x(\U1650/U1664/U28/Z ), .a(
        \U1650/U1664/x[3] ) );
    aoi222_1 \U1650/U1664/U32/U30/U1  ( .x(\U1650/U1664/x[0] ), .a(
        \U1650/ncd[1] ), .b(\U1650/ncd[0] ), .c(\U1650/ncd[1] ), .d(
        \U1650/U1664/U32/Z ), .e(\U1650/ncd[0] ), .f(\U1650/U1664/U32/Z ) );
    inv_1 \U1650/U1664/U32/U30/Uinv  ( .x(\U1650/U1664/U32/Z ), .a(
        \U1650/U1664/x[0] ) );
    aoi222_1 \U1650/U1664/U29/U30/U1  ( .x(\U1650/U1664/x[2] ), .a(
        \U1650/ncd[5] ), .b(\U1650/ncd[4] ), .c(\U1650/ncd[5] ), .d(
        \U1650/U1664/U29/Z ), .e(\U1650/ncd[4] ), .f(\U1650/U1664/U29/Z ) );
    inv_1 \U1650/U1664/U29/U30/Uinv  ( .x(\U1650/U1664/U29/Z ), .a(
        \U1650/U1664/x[2] ) );
    aoi222_1 \U1650/U1664/U33/U30/U1  ( .x(\U1650/U1664/y[0] ), .a(
        \U1650/U1664/x[1] ), .b(\U1650/U1664/x[0] ), .c(\U1650/U1664/x[1] ), 
        .d(\U1650/U1664/U33/Z ), .e(\U1650/U1664/x[0] ), .f(
        \U1650/U1664/U33/Z ) );
    inv_1 \U1650/U1664/U33/U30/Uinv  ( .x(\U1650/U1664/U33/Z ), .a(
        \U1650/U1664/y[0] ) );
    aoi222_1 \U1650/U1664/U30/U30/U1  ( .x(\U1650/U1664/y[1] ), .a(
        \U1650/U1664/x[3] ), .b(\U1650/U1664/x[2] ), .c(\U1650/U1664/x[3] ), 
        .d(\U1650/U1664/U30/Z ), .e(\U1650/U1664/x[2] ), .f(
        \U1650/U1664/U30/Z ) );
    inv_1 \U1650/U1664/U30/U30/Uinv  ( .x(\U1650/U1664/U30/Z ), .a(
        \U1650/U1664/y[1] ) );
    aoi222_1 \U1650/U1664/U31/U30/U1  ( .x(\U1650/U1664/x[1] ), .a(
        \U1650/ncd[3] ), .b(\U1650/ncd[2] ), .c(\U1650/ncd[3] ), .d(
        \U1650/U1664/U31/Z ), .e(\U1650/ncd[2] ), .f(\U1650/U1664/U31/Z ) );
    inv_1 \U1650/U1664/U31/U30/Uinv  ( .x(\U1650/U1664/U31/Z ), .a(
        \U1650/U1664/x[1] ) );
    aoi222_1 \U1650/U1664/U37/U30/U1  ( .x(\U1650/localcd ), .a(
        \U1650/U1664/y[0] ), .b(\U1650/U1664/y[1] ), .c(\U1650/U1664/y[0] ), 
        .d(\U1650/U1664/U37/Z ), .e(\U1650/U1664/y[1] ), .f(
        \U1650/U1664/U37/Z ) );
    inv_1 \U1650/U1664/U37/U30/Uinv  ( .x(\U1650/U1664/U37/Z ), .a(
        \U1650/localcd ) );
    nor3_1 \U1650/U1669/Unr  ( .x(\U1650/U1669/nr ), .a(
        \U1650/ctrlack_internal ), .b(\U1650/drivel ), .c(\U1650/driveh ) );
    nand3_1 \U1650/U1669/Und  ( .x(\U1650/U1669/nd ), .a(
        \U1650/ctrlack_internal ), .b(\U1650/drivel ), .c(\U1650/driveh ) );
    oa21_1 \U1650/U1669/U1  ( .x(\U1650/U1669/n2 ), .a(\U1650/U1669/n2 ), .b(
        \U1650/U1669/nr ), .c(\U1650/U1669/nd ) );
    inv_2 \U1650/U1669/U3  ( .x(net139), .a(\U1650/U1669/n2 ) );
    buf_2 \U1666/U1653  ( .x(\U1666/latch ), .a(net169) );
    nor2_1 \U1666/U264/U5  ( .x(\U1666/nlocalcd ), .a(reset), .b(
        \U1666/localcd ) );
    nor2_1 \U1666/U1659_0_/U5  ( .x(\U1666/ncd[0] ), .a(rd[24]), .b(rd[56]) );
    nor2_1 \U1666/U1659_1_/U5  ( .x(\U1666/ncd[1] ), .a(rd[25]), .b(rd[57]) );
    nor2_1 \U1666/U1659_2_/U5  ( .x(\U1666/ncd[2] ), .a(rd[26]), .b(rd[58]) );
    nor2_1 \U1666/U1659_3_/U5  ( .x(\U1666/ncd[3] ), .a(rd[27]), .b(rd[59]) );
    nor2_1 \U1666/U1659_4_/U5  ( .x(\U1666/ncd[4] ), .a(rd[28]), .b(rd[60]) );
    nor2_1 \U1666/U1659_5_/U5  ( .x(\U1666/ncd[5] ), .a(rd[29]), .b(rd[61]) );
    nor2_1 \U1666/U1659_6_/U5  ( .x(\U1666/ncd[6] ), .a(rd[30]), .b(rd[62]) );
    nor2_1 \U1666/U1659_7_/U5  ( .x(\U1666/ncd[7] ), .a(rd[31]), .b(rd[63]) );
    nor2_1 \U1666/U3/U5  ( .x(\U1666/ctrlack_internal ), .a(\U1666/acb ), .b(
        \U1666/ba ) );
    buf_2 \U1666/U1665/U7  ( .x(\U1666/driveh ), .a(read) );
    buf_2 \U1666/U1666/U7  ( .x(\U1666/drivel ), .a(read) );
    ao23_1 \U1666/U1658_0_/U21/U1/U1  ( .x(rd[24]), .a(n6), .b(rd[24]), .c(
        \U1666/drivel ), .d(cbl[0]), .e(n5) );
    ao23_1 \U1666/U1658_1_/U21/U1/U1  ( .x(rd[25]), .a(n6), .b(rd[25]), .c(
        \U1666/driveh ), .d(cbl[1]), .e(n5) );
    ao23_1 \U1666/U1658_2_/U21/U1/U1  ( .x(rd[26]), .a(\U1666/driveh ), .b(rd
        [26]), .c(n6), .d(cbl[2]), .e(n5) );
    ao23_1 \U1666/U1658_3_/U21/U1/U1  ( .x(rd[27]), .a(n6), .b(rd[27]), .c(
        \U1666/driveh ), .d(cbl[3]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1658_4_/U21/U1/U1  ( .x(rd[28]), .a(\U1666/drivel ), .b(rd
        [28]), .c(n6), .d(cbl[4]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1658_5_/U21/U1/U1  ( .x(rd[29]), .a(\U1666/drivel ), .b(rd
        [29]), .c(n6), .d(cbl[5]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1658_6_/U21/U1/U1  ( .x(rd[30]), .a(\U1666/driveh ), .b(rd
        [30]), .c(\U1666/drivel ), .d(cbl[6]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1658_7_/U21/U1/U1  ( .x(rd[31]), .a(\U1666/driveh ), .b(rd
        [31]), .c(\U1666/driveh ), .d(cbl[7]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_0_/U21/U1/U1  ( .x(rd[56]), .a(\U1666/drivel ), .b(rd
        [56]), .c(n6), .d(cbh[0]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_1_/U21/U1/U1  ( .x(rd[57]), .a(\U1666/driveh ), .b(rd
        [57]), .c(\U1666/drivel ), .d(cbh[1]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_2_/U21/U1/U1  ( .x(rd[58]), .a(\U1666/drivel ), .b(rd
        [58]), .c(\U1666/drivel ), .d(cbh[2]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_3_/U21/U1/U1  ( .x(rd[59]), .a(\U1666/driveh ), .b(rd
        [59]), .c(\U1666/driveh ), .d(cbh[3]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_4_/U21/U1/U1  ( .x(rd[60]), .a(\U1666/drivel ), .b(rd
        [60]), .c(\U1666/driveh ), .d(cbh[4]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_5_/U21/U1/U1  ( .x(rd[61]), .a(\U1666/driveh ), .b(rd
        [61]), .c(n6), .d(cbh[5]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_6_/U21/U1/U1  ( .x(rd[62]), .a(n6), .b(rd[62]), .c(
        \U1666/drivel ), .d(cbh[6]), .e(\U1666/latch ) );
    ao23_1 \U1666/U1651_7_/U21/U1/U1  ( .x(rd[63]), .a(n6), .b(rd[63]), .c(n6), 
        .d(cbh[7]), .e(\U1666/latch ) );
    aoai211_1 \U1666/U4/U28/U1/U1  ( .x(\U1666/U4/U28/U1/clr ), .a(read), .b(
        \U1666/acb ), .c(\U1666/nlocalcd ), .d(net169) );
    nand3_1 \U1666/U4/U28/U1/U2  ( .x(\U1666/U4/U28/U1/set ), .a(
        \U1666/nlocalcd ), .b(read), .c(\U1666/acb ) );
    nand2_2 \U1666/U4/U28/U1/U3  ( .x(net169), .a(\U1666/U4/U28/U1/clr ), .b(
        \U1666/U4/U28/U1/set ) );
    oai21_1 \U1666/U1/U30/U1/U1  ( .x(\U1666/acb ), .a(\U1666/U1/Z ), .b(
        \U1666/ba ), .c(read) );
    inv_1 \U1666/U1/U30/U1/U2  ( .x(\U1666/U1/Z ), .a(\U1666/acb ) );
    ao222_1 \U1666/U5/U18/U1/U1  ( .x(\U1666/ba ), .a(\U1666/latch ), .b(n14), 
        .c(\U1666/latch ), .d(\U1666/ba ), .e(n14), .f(\U1666/ba ) );
    aoi222_1 \U1666/U1664/U28/U30/U1  ( .x(\U1666/U1664/x[3] ), .a(
        \U1666/ncd[7] ), .b(\U1666/ncd[6] ), .c(\U1666/ncd[7] ), .d(
        \U1666/U1664/U28/Z ), .e(\U1666/ncd[6] ), .f(\U1666/U1664/U28/Z ) );
    inv_1 \U1666/U1664/U28/U30/Uinv  ( .x(\U1666/U1664/U28/Z ), .a(
        \U1666/U1664/x[3] ) );
    aoi222_1 \U1666/U1664/U32/U30/U1  ( .x(\U1666/U1664/x[0] ), .a(
        \U1666/ncd[1] ), .b(\U1666/ncd[0] ), .c(\U1666/ncd[1] ), .d(
        \U1666/U1664/U32/Z ), .e(\U1666/ncd[0] ), .f(\U1666/U1664/U32/Z ) );
    inv_1 \U1666/U1664/U32/U30/Uinv  ( .x(\U1666/U1664/U32/Z ), .a(
        \U1666/U1664/x[0] ) );
    aoi222_1 \U1666/U1664/U29/U30/U1  ( .x(\U1666/U1664/x[2] ), .a(
        \U1666/ncd[5] ), .b(\U1666/ncd[4] ), .c(\U1666/ncd[5] ), .d(
        \U1666/U1664/U29/Z ), .e(\U1666/ncd[4] ), .f(\U1666/U1664/U29/Z ) );
    inv_1 \U1666/U1664/U29/U30/Uinv  ( .x(\U1666/U1664/U29/Z ), .a(
        \U1666/U1664/x[2] ) );
    aoi222_1 \U1666/U1664/U33/U30/U1  ( .x(\U1666/U1664/y[0] ), .a(
        \U1666/U1664/x[1] ), .b(\U1666/U1664/x[0] ), .c(\U1666/U1664/x[1] ), 
        .d(\U1666/U1664/U33/Z ), .e(\U1666/U1664/x[0] ), .f(
        \U1666/U1664/U33/Z ) );
    inv_1 \U1666/U1664/U33/U30/Uinv  ( .x(\U1666/U1664/U33/Z ), .a(
        \U1666/U1664/y[0] ) );
    aoi222_1 \U1666/U1664/U30/U30/U1  ( .x(\U1666/U1664/y[1] ), .a(
        \U1666/U1664/x[3] ), .b(\U1666/U1664/x[2] ), .c(\U1666/U1664/x[3] ), 
        .d(\U1666/U1664/U30/Z ), .e(\U1666/U1664/x[2] ), .f(
        \U1666/U1664/U30/Z ) );
    inv_1 \U1666/U1664/U30/U30/Uinv  ( .x(\U1666/U1664/U30/Z ), .a(
        \U1666/U1664/y[1] ) );
    aoi222_1 \U1666/U1664/U31/U30/U1  ( .x(\U1666/U1664/x[1] ), .a(
        \U1666/ncd[3] ), .b(\U1666/ncd[2] ), .c(\U1666/ncd[3] ), .d(
        \U1666/U1664/U31/Z ), .e(\U1666/ncd[2] ), .f(\U1666/U1664/U31/Z ) );
    inv_1 \U1666/U1664/U31/U30/Uinv  ( .x(\U1666/U1664/U31/Z ), .a(
        \U1666/U1664/x[1] ) );
    aoi222_1 \U1666/U1664/U37/U30/U1  ( .x(\U1666/localcd ), .a(
        \U1666/U1664/y[0] ), .b(\U1666/U1664/y[1] ), .c(\U1666/U1664/y[0] ), 
        .d(\U1666/U1664/U37/Z ), .e(\U1666/U1664/y[1] ), .f(
        \U1666/U1664/U37/Z ) );
    inv_1 \U1666/U1664/U37/U30/Uinv  ( .x(\U1666/U1664/U37/Z ), .a(
        \U1666/localcd ) );
    nor3_1 \U1666/U1669/Unr  ( .x(\U1666/U1669/nr ), .a(
        \U1666/ctrlack_internal ), .b(n6), .c(\U1666/drivel ) );
    nand3_1 \U1666/U1669/Und  ( .x(\U1666/U1669/nd ), .a(
        \U1666/ctrlack_internal ), .b(\U1666/driveh ), .c(\U1666/drivel ) );
    oa21_1 \U1666/U1669/U1  ( .x(\U1666/U1669/n2 ), .a(\U1666/U1669/n2 ), .b(
        \U1666/U1669/nr ), .c(\U1666/U1669/nd ) );
    inv_2 \U1666/U1669/U3  ( .x(net94), .a(\U1666/U1669/n2 ) );
    buf_2 \I1/U1653  ( .x(\I1/latch ), .a(net166) );
    nor2_1 \I1/U264/U5  ( .x(\I1/nlocalcd ), .a(reset), .b(\I1/localcd ) );
    nor2_1 \I1/U1659_0_/U5  ( .x(\I1/ncd[0] ), .a(rd[8]), .b(rd[40]) );
    nor2_1 \I1/U1659_1_/U5  ( .x(\I1/ncd[1] ), .a(rd[9]), .b(rd[41]) );
    nor2_1 \I1/U1659_2_/U5  ( .x(\I1/ncd[2] ), .a(rd[10]), .b(rd[42]) );
    nor2_1 \I1/U1659_3_/U5  ( .x(\I1/ncd[3] ), .a(rd[11]), .b(rd[43]) );
    nor2_1 \I1/U1659_4_/U5  ( .x(\I1/ncd[4] ), .a(rd[12]), .b(rd[44]) );
    nor2_1 \I1/U1659_5_/U5  ( .x(\I1/ncd[5] ), .a(rd[13]), .b(rd[45]) );
    nor2_1 \I1/U1659_6_/U5  ( .x(\I1/ncd[6] ), .a(rd[14]), .b(rd[46]) );
    nor2_1 \I1/U1659_7_/U5  ( .x(\I1/ncd[7] ), .a(rd[15]), .b(rd[47]) );
    nor2_1 \I1/U3/U5  ( .x(\I1/ctrlack_internal ), .a(\I1/acb ), .b(\I1/ba )
         );
    buf_2 \I1/U1665/U7  ( .x(\I1/driveh ), .a(net103) );
    buf_2 \I1/U1666/U7  ( .x(\I1/drivel ), .a(net103) );
    ao23_1 \I1/U1658_0_/U21/U1/U1  ( .x(rd[8]), .a(n4), .b(rd[8]), .c(
        \I1/drivel ), .d(cbl[0]), .e(n3) );
    ao23_1 \I1/U1658_1_/U21/U1/U1  ( .x(rd[9]), .a(n4), .b(rd[9]), .c(
        \I1/driveh ), .d(cbl[1]), .e(n3) );
    ao23_1 \I1/U1658_2_/U21/U1/U1  ( .x(rd[10]), .a(\I1/driveh ), .b(rd[10]), 
        .c(n4), .d(cbl[2]), .e(n3) );
    ao23_1 \I1/U1658_3_/U21/U1/U1  ( .x(rd[11]), .a(n4), .b(rd[11]), .c(
        \I1/driveh ), .d(cbl[3]), .e(\I1/latch ) );
    ao23_1 \I1/U1658_4_/U21/U1/U1  ( .x(rd[12]), .a(\I1/drivel ), .b(rd[12]), 
        .c(n4), .d(cbl[4]), .e(\I1/latch ) );
    ao23_1 \I1/U1658_5_/U21/U1/U1  ( .x(rd[13]), .a(\I1/drivel ), .b(rd[13]), 
        .c(n4), .d(cbl[5]), .e(\I1/latch ) );
    ao23_1 \I1/U1658_6_/U21/U1/U1  ( .x(rd[14]), .a(\I1/driveh ), .b(rd[14]), 
        .c(\I1/drivel ), .d(cbl[6]), .e(\I1/latch ) );
    ao23_1 \I1/U1658_7_/U21/U1/U1  ( .x(rd[15]), .a(\I1/driveh ), .b(rd[15]), 
        .c(\I1/driveh ), .d(cbl[7]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_0_/U21/U1/U1  ( .x(rd[40]), .a(\I1/drivel ), .b(rd[40]), 
        .c(n4), .d(cbh[0]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_1_/U21/U1/U1  ( .x(rd[41]), .a(\I1/driveh ), .b(rd[41]), 
        .c(\I1/drivel ), .d(cbh[1]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_2_/U21/U1/U1  ( .x(rd[42]), .a(\I1/drivel ), .b(rd[42]), 
        .c(\I1/drivel ), .d(cbh[2]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_3_/U21/U1/U1  ( .x(rd[43]), .a(\I1/driveh ), .b(rd[43]), 
        .c(\I1/driveh ), .d(cbh[3]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_4_/U21/U1/U1  ( .x(rd[44]), .a(\I1/drivel ), .b(rd[44]), 
        .c(\I1/driveh ), .d(cbh[4]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_5_/U21/U1/U1  ( .x(rd[45]), .a(\I1/driveh ), .b(rd[45]), 
        .c(n4), .d(cbh[5]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_6_/U21/U1/U1  ( .x(rd[46]), .a(n4), .b(rd[46]), .c(
        \I1/drivel ), .d(cbh[6]), .e(\I1/latch ) );
    ao23_1 \I1/U1651_7_/U21/U1/U1  ( .x(rd[47]), .a(n4), .b(rd[47]), .c(n4), 
        .d(cbh[7]), .e(\I1/latch ) );
    aoai211_1 \I1/U4/U28/U1/U1  ( .x(\I1/U4/U28/U1/clr ), .a(net103), .b(
        \I1/acb ), .c(\I1/nlocalcd ), .d(net166) );
    nand3_1 \I1/U4/U28/U1/U2  ( .x(\I1/U4/U28/U1/set ), .a(\I1/nlocalcd ), .b(
        net103), .c(\I1/acb ) );
    nand2_2 \I1/U4/U28/U1/U3  ( .x(net166), .a(\I1/U4/U28/U1/clr ), .b(
        \I1/U4/U28/U1/set ) );
    oai21_1 \I1/U1/U30/U1/U1  ( .x(\I1/acb ), .a(\I1/U1/Z ), .b(\I1/ba ), .c(
        net103) );
    inv_1 \I1/U1/U30/U1/U2  ( .x(\I1/U1/Z ), .a(\I1/acb ) );
    ao222_1 \I1/U5/U18/U1/U1  ( .x(\I1/ba ), .a(\I1/latch ), .b(n14), .c(
        \I1/latch ), .d(\I1/ba ), .e(n14), .f(\I1/ba ) );
    aoi222_1 \I1/U1664/U28/U30/U1  ( .x(\I1/U1664/x[3] ), .a(\I1/ncd[7] ), .b(
        \I1/ncd[6] ), .c(\I1/ncd[7] ), .d(\I1/U1664/U28/Z ), .e(\I1/ncd[6] ), 
        .f(\I1/U1664/U28/Z ) );
    inv_1 \I1/U1664/U28/U30/Uinv  ( .x(\I1/U1664/U28/Z ), .a(\I1/U1664/x[3] )
         );
    aoi222_1 \I1/U1664/U32/U30/U1  ( .x(\I1/U1664/x[0] ), .a(\I1/ncd[1] ), .b(
        \I1/ncd[0] ), .c(\I1/ncd[1] ), .d(\I1/U1664/U32/Z ), .e(\I1/ncd[0] ), 
        .f(\I1/U1664/U32/Z ) );
    inv_1 \I1/U1664/U32/U30/Uinv  ( .x(\I1/U1664/U32/Z ), .a(\I1/U1664/x[0] )
         );
    aoi222_1 \I1/U1664/U29/U30/U1  ( .x(\I1/U1664/x[2] ), .a(\I1/ncd[5] ), .b(
        \I1/ncd[4] ), .c(\I1/ncd[5] ), .d(\I1/U1664/U29/Z ), .e(\I1/ncd[4] ), 
        .f(\I1/U1664/U29/Z ) );
    inv_1 \I1/U1664/U29/U30/Uinv  ( .x(\I1/U1664/U29/Z ), .a(\I1/U1664/x[2] )
         );
    aoi222_1 \I1/U1664/U33/U30/U1  ( .x(\I1/U1664/y[0] ), .a(\I1/U1664/x[1] ), 
        .b(\I1/U1664/x[0] ), .c(\I1/U1664/x[1] ), .d(\I1/U1664/U33/Z ), .e(
        \I1/U1664/x[0] ), .f(\I1/U1664/U33/Z ) );
    inv_1 \I1/U1664/U33/U30/Uinv  ( .x(\I1/U1664/U33/Z ), .a(\I1/U1664/y[0] )
         );
    aoi222_1 \I1/U1664/U30/U30/U1  ( .x(\I1/U1664/y[1] ), .a(\I1/U1664/x[3] ), 
        .b(\I1/U1664/x[2] ), .c(\I1/U1664/x[3] ), .d(\I1/U1664/U30/Z ), .e(
        \I1/U1664/x[2] ), .f(\I1/U1664/U30/Z ) );
    inv_1 \I1/U1664/U30/U30/Uinv  ( .x(\I1/U1664/U30/Z ), .a(\I1/U1664/y[1] )
         );
    aoi222_1 \I1/U1664/U31/U30/U1  ( .x(\I1/U1664/x[1] ), .a(\I1/ncd[3] ), .b(
        \I1/ncd[2] ), .c(\I1/ncd[3] ), .d(\I1/U1664/U31/Z ), .e(\I1/ncd[2] ), 
        .f(\I1/U1664/U31/Z ) );
    inv_1 \I1/U1664/U31/U30/Uinv  ( .x(\I1/U1664/U31/Z ), .a(\I1/U1664/x[1] )
         );
    aoi222_1 \I1/U1664/U37/U30/U1  ( .x(\I1/localcd ), .a(\I1/U1664/y[0] ), 
        .b(\I1/U1664/y[1] ), .c(\I1/U1664/y[0] ), .d(\I1/U1664/U37/Z ), .e(
        \I1/U1664/y[1] ), .f(\I1/U1664/U37/Z ) );
    inv_1 \I1/U1664/U37/U30/Uinv  ( .x(\I1/U1664/U37/Z ), .a(\I1/localcd ) );
    nor3_1 \I1/U1669/Unr  ( .x(\I1/U1669/nr ), .a(\I1/ctrlack_internal ), .b(
        n4), .c(\I1/drivel ) );
    nand3_1 \I1/U1669/Und  ( .x(\I1/U1669/nd ), .a(\I1/ctrlack_internal ), .b(
        \I1/driveh ), .c(\I1/drivel ) );
    oa21_1 \I1/U1669/U1  ( .x(\I1/U1669/n2 ), .a(\I1/U1669/n2 ), .b(
        \I1/U1669/nr ), .c(\I1/U1669/nd ) );
    inv_2 \I1/U1669/U3  ( .x(read_lhw), .a(\I1/U1669/n2 ) );
    buf_2 \I2/U1653  ( .x(\I2/latch ), .a(net170) );
    nor2_1 \I2/U264/U5  ( .x(\I2/nlocalcd ), .a(reset), .b(\I2/localcd ) );
    nor2_1 \I2/U1659_0_/U5  ( .x(\I2/ncd[0] ), .a(rd[16]), .b(rd[48]) );
    nor2_1 \I2/U1659_1_/U5  ( .x(\I2/ncd[1] ), .a(rd[17]), .b(rd[49]) );
    nor2_1 \I2/U1659_2_/U5  ( .x(\I2/ncd[2] ), .a(rd[18]), .b(rd[50]) );
    nor2_1 \I2/U1659_3_/U5  ( .x(\I2/ncd[3] ), .a(rd[19]), .b(rd[51]) );
    nor2_1 \I2/U1659_4_/U5  ( .x(\I2/ncd[4] ), .a(rd[20]), .b(rd[52]) );
    nor2_1 \I2/U1659_5_/U5  ( .x(\I2/ncd[5] ), .a(rd[21]), .b(rd[53]) );
    nor2_1 \I2/U1659_6_/U5  ( .x(\I2/ncd[6] ), .a(rd[22]), .b(rd[54]) );
    nor2_1 \I2/U1659_7_/U5  ( .x(\I2/ncd[7] ), .a(rd[23]), .b(rd[55]) );
    nor2_1 \I2/U3/U5  ( .x(\I2/ctrlack_internal ), .a(\I2/acb ), .b(\I2/ba )
         );
    buf_2 \I2/U1665/U7  ( .x(\I2/driveh ), .a(net94) );
    buf_2 \I2/U1666/U7  ( .x(\I2/drivel ), .a(net94) );
    ao23_1 \I2/U1658_0_/U21/U1/U1  ( .x(rd[16]), .a(n2), .b(rd[16]), .c(
        \I2/drivel ), .d(cbl[0]), .e(n1) );
    ao23_1 \I2/U1658_1_/U21/U1/U1  ( .x(rd[17]), .a(n2), .b(rd[17]), .c(
        \I2/driveh ), .d(cbl[1]), .e(n1) );
    ao23_1 \I2/U1658_2_/U21/U1/U1  ( .x(rd[18]), .a(\I2/driveh ), .b(rd[18]), 
        .c(n2), .d(cbl[2]), .e(n1) );
    ao23_1 \I2/U1658_3_/U21/U1/U1  ( .x(rd[19]), .a(n2), .b(rd[19]), .c(
        \I2/driveh ), .d(cbl[3]), .e(\I2/latch ) );
    ao23_1 \I2/U1658_4_/U21/U1/U1  ( .x(rd[20]), .a(\I2/drivel ), .b(rd[20]), 
        .c(n2), .d(cbl[4]), .e(\I2/latch ) );
    ao23_1 \I2/U1658_5_/U21/U1/U1  ( .x(rd[21]), .a(\I2/drivel ), .b(rd[21]), 
        .c(n2), .d(cbl[5]), .e(\I2/latch ) );
    ao23_1 \I2/U1658_6_/U21/U1/U1  ( .x(rd[22]), .a(\I2/driveh ), .b(rd[22]), 
        .c(\I2/drivel ), .d(cbl[6]), .e(\I2/latch ) );
    ao23_1 \I2/U1658_7_/U21/U1/U1  ( .x(rd[23]), .a(\I2/driveh ), .b(rd[23]), 
        .c(\I2/driveh ), .d(cbl[7]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_0_/U21/U1/U1  ( .x(rd[48]), .a(\I2/drivel ), .b(rd[48]), 
        .c(n2), .d(cbh[0]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_1_/U21/U1/U1  ( .x(rd[49]), .a(\I2/driveh ), .b(rd[49]), 
        .c(\I2/drivel ), .d(cbh[1]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_2_/U21/U1/U1  ( .x(rd[50]), .a(\I2/drivel ), .b(rd[50]), 
        .c(\I2/drivel ), .d(cbh[2]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_3_/U21/U1/U1  ( .x(rd[51]), .a(\I2/driveh ), .b(rd[51]), 
        .c(\I2/driveh ), .d(cbh[3]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_4_/U21/U1/U1  ( .x(rd[52]), .a(\I2/drivel ), .b(rd[52]), 
        .c(\I2/driveh ), .d(cbh[4]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_5_/U21/U1/U1  ( .x(rd[53]), .a(\I2/driveh ), .b(rd[53]), 
        .c(n2), .d(cbh[5]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_6_/U21/U1/U1  ( .x(rd[54]), .a(n2), .b(rd[54]), .c(
        \I2/drivel ), .d(cbh[6]), .e(\I2/latch ) );
    ao23_1 \I2/U1651_7_/U21/U1/U1  ( .x(rd[55]), .a(n2), .b(rd[55]), .c(n2), 
        .d(cbh[7]), .e(\I2/latch ) );
    aoai211_1 \I2/U4/U28/U1/U1  ( .x(\I2/U4/U28/U1/clr ), .a(net94), .b(
        \I2/acb ), .c(\I2/nlocalcd ), .d(net170) );
    nand3_1 \I2/U4/U28/U1/U2  ( .x(\I2/U4/U28/U1/set ), .a(\I2/nlocalcd ), .b(
        net94), .c(\I2/acb ) );
    nand2_2 \I2/U4/U28/U1/U3  ( .x(net170), .a(\I2/U4/U28/U1/clr ), .b(
        \I2/U4/U28/U1/set ) );
    oai21_1 \I2/U1/U30/U1/U1  ( .x(\I2/acb ), .a(\I2/U1/Z ), .b(\I2/ba ), .c(
        net94) );
    inv_1 \I2/U1/U30/U1/U2  ( .x(\I2/U1/Z ), .a(\I2/acb ) );
    ao222_1 \I2/U5/U18/U1/U1  ( .x(\I2/ba ), .a(\I2/latch ), .b(n14), .c(
        \I2/latch ), .d(\I2/ba ), .e(n14), .f(\I2/ba ) );
    aoi222_1 \I2/U1664/U28/U30/U1  ( .x(\I2/U1664/x[3] ), .a(\I2/ncd[7] ), .b(
        \I2/ncd[6] ), .c(\I2/ncd[7] ), .d(\I2/U1664/U28/Z ), .e(\I2/ncd[6] ), 
        .f(\I2/U1664/U28/Z ) );
    inv_1 \I2/U1664/U28/U30/Uinv  ( .x(\I2/U1664/U28/Z ), .a(\I2/U1664/x[3] )
         );
    aoi222_1 \I2/U1664/U32/U30/U1  ( .x(\I2/U1664/x[0] ), .a(\I2/ncd[1] ), .b(
        \I2/ncd[0] ), .c(\I2/ncd[1] ), .d(\I2/U1664/U32/Z ), .e(\I2/ncd[0] ), 
        .f(\I2/U1664/U32/Z ) );
    inv_1 \I2/U1664/U32/U30/Uinv  ( .x(\I2/U1664/U32/Z ), .a(\I2/U1664/x[0] )
         );
    aoi222_1 \I2/U1664/U29/U30/U1  ( .x(\I2/U1664/x[2] ), .a(\I2/ncd[5] ), .b(
        \I2/ncd[4] ), .c(\I2/ncd[5] ), .d(\I2/U1664/U29/Z ), .e(\I2/ncd[4] ), 
        .f(\I2/U1664/U29/Z ) );
    inv_1 \I2/U1664/U29/U30/Uinv  ( .x(\I2/U1664/U29/Z ), .a(\I2/U1664/x[2] )
         );
    aoi222_1 \I2/U1664/U33/U30/U1  ( .x(\I2/U1664/y[0] ), .a(\I2/U1664/x[1] ), 
        .b(\I2/U1664/x[0] ), .c(\I2/U1664/x[1] ), .d(\I2/U1664/U33/Z ), .e(
        \I2/U1664/x[0] ), .f(\I2/U1664/U33/Z ) );
    inv_1 \I2/U1664/U33/U30/Uinv  ( .x(\I2/U1664/U33/Z ), .a(\I2/U1664/y[0] )
         );
    aoi222_1 \I2/U1664/U30/U30/U1  ( .x(\I2/U1664/y[1] ), .a(\I2/U1664/x[3] ), 
        .b(\I2/U1664/x[2] ), .c(\I2/U1664/x[3] ), .d(\I2/U1664/U30/Z ), .e(
        \I2/U1664/x[2] ), .f(\I2/U1664/U30/Z ) );
    inv_1 \I2/U1664/U30/U30/Uinv  ( .x(\I2/U1664/U30/Z ), .a(\I2/U1664/y[1] )
         );
    aoi222_1 \I2/U1664/U31/U30/U1  ( .x(\I2/U1664/x[1] ), .a(\I2/ncd[3] ), .b(
        \I2/ncd[2] ), .c(\I2/ncd[3] ), .d(\I2/U1664/U31/Z ), .e(\I2/ncd[2] ), 
        .f(\I2/U1664/U31/Z ) );
    inv_1 \I2/U1664/U31/U30/Uinv  ( .x(\I2/U1664/U31/Z ), .a(\I2/U1664/x[1] )
         );
    aoi222_1 \I2/U1664/U37/U30/U1  ( .x(\I2/localcd ), .a(\I2/U1664/y[0] ), 
        .b(\I2/U1664/y[1] ), .c(\I2/U1664/y[0] ), .d(\I2/U1664/U37/Z ), .e(
        \I2/U1664/y[1] ), .f(\I2/U1664/U37/Z ) );
    inv_1 \I2/U1664/U37/U30/Uinv  ( .x(\I2/U1664/U37/Z ), .a(\I2/localcd ) );
    nor3_1 \I2/U1669/Unr  ( .x(\I2/U1669/nr ), .a(\I2/ctrlack_internal ), .b(
        n2), .c(\I2/drivel ) );
    nand3_1 \I2/U1669/Und  ( .x(\I2/U1669/nd ), .a(\I2/ctrlack_internal ), .b(
        \I2/driveh ), .c(\I2/drivel ) );
    oa21_1 \I2/U1669/U1  ( .x(\I2/U1669/n2 ), .a(\I2/U1669/n2 ), .b(
        \I2/U1669/nr ), .c(\I2/U1669/nd ) );
    inv_2 \I2/U1669/U3  ( .x(net103), .a(\I2/U1669/n2 ) );
    buf_1 U1 ( .x(n1), .a(\I2/latch ) );
    buf_2 U2 ( .x(n2), .a(net94) );
    buf_1 U3 ( .x(n3), .a(\I1/latch ) );
    buf_2 U4 ( .x(n4), .a(net103) );
    buf_1 U5 ( .x(n5), .a(\U1666/latch ) );
    buf_2 U6 ( .x(n6), .a(read) );
    buf_1 U7 ( .x(n7), .a(\U1650/latch ) );
    buf_1 U8 ( .x(n8), .a(\U1650/driveh ) );
    buf_1 U9 ( .x(n9), .a(\U1650/drivel ) );
    buf_1 U10 ( .x(n10), .a(\U1667/latch ) );
    buf_2 U11 ( .x(n11), .a(read_lhw) );
    buf_1 U12 ( .x(n12), .a(\I6/latch ) );
    buf_2 U13 ( .x(n13), .a(net139) );
    buf_3 U14 ( .x(n14), .a(bpullcd) );
    buf_3 U15 ( .x(err[0]), .a(n18) );
    buf_3 U16 ( .x(err[1]), .a(n17) );
endmodule


module chain_fr2dr_byte_5 ( nia, oh, ol, i, nReset, noa );
output [7:0] oh;
output [7:0] ol;
input  [4:0] i;
input  nReset, noa;
output nia;
    wire nbReset, eop, ncla, csela, asela, \U891/reset , \U891/neopack , 
        \U891/iay , \U891/naack[0] , \U891/naack[1] , \U891/U1128/nb , \b[3] , 
        \b[2] , \U891/U1128/na , \b[1] , \b[0] , \U891/ackb , \a[3] , \a[2] , 
        \U891/nack , \U891/acka , \a[1] , \a[0] , bsela, bsel, asel, 
        \U891/U1118_0_/nr , naa, \U891/U1118_0_/nd , \U891/U1118_0_/n2 , 
        \U891/U1118_1_/nr , \U891/U1118_1_/nd , \U891/U1118_1_/n2 , 
        \U891/U1118_2_/nr , \U891/U1118_2_/nd , \U891/U1118_2_/n2 , 
        \U891/U1118_3_/nr , \U891/U1118_3_/nd , \U891/U1118_3_/n2 , 
        \U891/U1117_0_/nr , nba, \U891/U1117_0_/nd , \U891/U1117_0_/n2 , 
        \U891/U1117_1_/nr , \U891/U1117_1_/nd , \U891/U1117_1_/n2 , 
        \U891/U1117_2_/nr , \U891/U1117_2_/nd , \U891/U1117_2_/n2 , 
        \U891/U1117_3_/nr , \U891/U1117_3_/nd , \U891/U1117_3_/n2 , 
        \U886/reset , \U886/U1128/nb , \f[3] , \f[2] , \U886/U1128/na , \f[1] , 
        \f[0] , \U886/ackb , \U886/nack , \U886/acka , \U886/U1127/n5 , 
        \U886/U1127/n1 , \U886/U1127/n2 , \U886/U1127/n3 , \U886/U1127/n4 , 
        \e[3] , \e[2] , \e[1] , \e[0] , fsela, fsel, esela, esel, 
        \U886/U1118_0_/nr , nea, \U886/U1118_0_/nd , \U886/U1118_0_/n2 , 
        \U886/U1118_1_/nr , \U886/U1118_1_/nd , \U886/U1118_1_/n2 , 
        \U886/U1118_2_/nr , \U886/U1118_2_/nd , \U886/U1118_2_/n2 , 
        \U886/U1118_3_/nr , \U886/U1118_3_/nd , \U886/U1118_3_/n2 , 
        \U886/U1117_0_/nr , nfa, \U886/U1117_0_/nd , \U886/U1117_0_/n2 , 
        \U886/U1117_1_/nr , \U886/U1117_1_/nd , \U886/U1117_1_/n2 , 
        \U886/U1117_2_/nr , \U886/U1117_2_/nd , \U886/U1117_2_/n2 , 
        \U886/U1117_3_/nr , \U886/U1117_3_/nd , \U886/U1117_3_/n2 , 
        \U884/reset , \U884/U1128/nb , \d[3] , \d[2] , \U884/U1128/na , \d[1] , 
        \d[0] , \U884/ackb , \U884/nack , \U884/acka , \U884/U1127/n5 , 
        \U884/U1127/n1 , \U884/U1127/n2 , \U884/U1127/n3 , \U884/U1127/n4 , 
        \c[3] , \c[2] , \c[1] , \c[0] , dsela, dsel, csel, \U884/U1118_0_/nr , 
        nca, \U884/U1118_0_/nd , \U884/U1118_0_/n2 , \U884/U1118_1_/nr , 
        \U884/U1118_1_/nd , \U884/U1118_1_/n2 , \U884/U1118_2_/nr , 
        \U884/U1118_2_/nd , \U884/U1118_2_/n2 , \U884/U1118_3_/nr , 
        \U884/U1118_3_/nd , \U884/U1118_3_/n2 , \U884/U1117_0_/nr , nda, 
        \U884/U1117_0_/nd , \U884/U1117_0_/n2 , \U884/U1117_1_/nr , 
        \U884/U1117_1_/nd , \U884/U1117_1_/n2 , \U884/U1117_2_/nr , 
        \U884/U1117_2_/nd , \U884/U1117_2_/n2 , \U884/U1117_3_/nr , 
        \U884/U1117_3_/nd , \U884/U1117_3_/n2 , \U888/s , \U888/r , 
        \U888/nback , \U888/naack , \U888/reset , \U887/s , \U887/r , 
        \U887/nback , \U887/naack , \U887/reset , \U885/s , \U885/r , 
        \U885/nback , \U885/naack , \U885/reset , \U877/x , \U877/reset , 
        \U877/y , \U877/U590/U25/U1/clr , net135, \cl[3] , \cl[1] , 
        \U877/U590/U25/U1/ob , n1, \U877/U589/U25/U1/clr , \cl[0] , 
        \U877/U589/U25/U1/ob , \U877/U588/U25/U1/clr , \cl[2] , 
        \U877/U588/U25/U1/ob , \U877/U591/U25/U1/clr , \U877/U591/U25/U1/ob , 
        \U876/x , \U876/reset , \U876/y , \U876/U590/U25/U1/clr , 
        \U876/U590/U25/U1/ob , \U876/U589/U25/U1/clr , \U876/U589/U25/U1/ob , 
        \U876/U588/U25/U1/clr , \U876/U588/U25/U1/ob , \U876/U591/U25/U1/clr , 
        \U876/U591/U25/U1/ob , \U2/x , \U2/reset , \U2/y , 
        \U2/U590/U25/U1/clr , \U2/U590/U25/U1/ob , \U2/U589/U25/U1/clr , 
        \U2/U589/U25/U1/ob , \U2/U588/U25/U1/clr , \U2/U588/U25/U1/ob , 
        \U2/U591/U25/U1/clr , \U2/U591/U25/U1/ob , \U1/x , \U1/reset , \U1/y , 
        \U1/U590/U25/U1/clr , \U1/U590/U25/U1/ob , \U1/U589/U25/U1/clr , 
        \U1/U589/U25/U1/ob , \U1/U588/U25/U1/clr , \U1/U588/U25/U1/ob , 
        \U1/U591/U25/U1/clr , \U1/U591/U25/U1/ob , \U881/nack[1] , 
        \U881/nack[0] ;
    buf_2 U897 ( .x(nbReset), .a(nReset) );
    and4_1 \U894/U12  ( .x(eop), .a(ncla), .b(csela), .c(asela), .d(i[4]) );
    inv_1 \U891/U1126/U3  ( .x(\U891/reset ), .a(nbReset) );
    inv_1 \U891/U1139/U3  ( .x(\U891/neopack ), .a(eop) );
    nand3_1 \U891/U1131/U9  ( .x(\U891/iay ), .a(\U891/neopack ), .b(
        \U891/naack[0] ), .c(\U891/naack[1] ) );
    nor3_1 \U891/U1128/U27  ( .x(\U891/U1128/nb ), .a(\U891/reset ), .b(\b[3] 
        ), .c(\b[2] ) );
    nor2_1 \U891/U1128/U26  ( .x(\U891/U1128/na ), .a(\b[1] ), .b(\b[0] ) );
    nand2_2 \U891/U1128/U29  ( .x(\U891/ackb ), .a(\U891/U1128/nb ), .b(
        \U891/U1128/na ) );
    nor2_1 \U891/U1133/U5  ( .x(\U891/naack[0] ), .a(\a[3] ), .b(\a[2] ) );
    nor2_1 \U891/U1108/U5  ( .x(\U891/nack ), .a(\U891/acka ), .b(\U891/ackb )
         );
    nor2_1 \U891/U1134/U5  ( .x(\U891/naack[1] ), .a(\a[1] ), .b(\a[0] ) );
    nor2_2 \U891/U914/U6  ( .x(nia), .a(\U891/iay ), .b(\U891/ackb ) );
    nand2_1 \U891/U1130/U5  ( .x(\U891/acka ), .a(\U891/naack[0] ), .b(
        \U891/naack[1] ) );
    ao222_4 \U891/U1121/U1/U1  ( .x(bsela), .a(\U891/nack ), .b(bsel), .c(
        \U891/nack ), .d(bsela), .e(bsel), .f(bsela) );
    ao222_4 \U891/U1120/U1/U1  ( .x(asela), .a(asel), .b(\U891/nack ), .c(asel
        ), .d(asela), .e(\U891/nack ), .f(asela) );
    nor3_1 \U891/U1118_0_/Unr  ( .x(\U891/U1118_0_/nr ), .a(i[0]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_0_/Und  ( .x(\U891/U1118_0_/nd ), .a(i[0]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_0_/U1  ( .x(\U891/U1118_0_/n2 ), .a(\U891/U1118_0_/n2 ), 
        .b(\U891/U1118_0_/nr ), .c(\U891/U1118_0_/nd ) );
    inv_2 \U891/U1118_0_/U3  ( .x(\a[0] ), .a(\U891/U1118_0_/n2 ) );
    nor3_1 \U891/U1118_1_/Unr  ( .x(\U891/U1118_1_/nr ), .a(i[1]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_1_/Und  ( .x(\U891/U1118_1_/nd ), .a(i[1]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_1_/U1  ( .x(\U891/U1118_1_/n2 ), .a(\U891/U1118_1_/n2 ), 
        .b(\U891/U1118_1_/nr ), .c(\U891/U1118_1_/nd ) );
    inv_2 \U891/U1118_1_/U3  ( .x(\a[1] ), .a(\U891/U1118_1_/n2 ) );
    nor3_1 \U891/U1118_2_/Unr  ( .x(\U891/U1118_2_/nr ), .a(i[2]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_2_/Und  ( .x(\U891/U1118_2_/nd ), .a(i[2]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_2_/U1  ( .x(\U891/U1118_2_/n2 ), .a(\U891/U1118_2_/n2 ), 
        .b(\U891/U1118_2_/nr ), .c(\U891/U1118_2_/nd ) );
    inv_2 \U891/U1118_2_/U3  ( .x(\a[2] ), .a(\U891/U1118_2_/n2 ) );
    nor3_1 \U891/U1118_3_/Unr  ( .x(\U891/U1118_3_/nr ), .a(i[3]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_3_/Und  ( .x(\U891/U1118_3_/nd ), .a(i[3]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_3_/U1  ( .x(\U891/U1118_3_/n2 ), .a(\U891/U1118_3_/n2 ), 
        .b(\U891/U1118_3_/nr ), .c(\U891/U1118_3_/nd ) );
    inv_2 \U891/U1118_3_/U3  ( .x(\a[3] ), .a(\U891/U1118_3_/n2 ) );
    nor3_1 \U891/U1117_0_/Unr  ( .x(\U891/U1117_0_/nr ), .a(i[0]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_0_/Und  ( .x(\U891/U1117_0_/nd ), .a(i[0]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_0_/U1  ( .x(\U891/U1117_0_/n2 ), .a(\U891/U1117_0_/n2 ), 
        .b(\U891/U1117_0_/nr ), .c(\U891/U1117_0_/nd ) );
    inv_2 \U891/U1117_0_/U3  ( .x(\b[0] ), .a(\U891/U1117_0_/n2 ) );
    nor3_1 \U891/U1117_1_/Unr  ( .x(\U891/U1117_1_/nr ), .a(i[1]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_1_/Und  ( .x(\U891/U1117_1_/nd ), .a(i[1]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_1_/U1  ( .x(\U891/U1117_1_/n2 ), .a(\U891/U1117_1_/n2 ), 
        .b(\U891/U1117_1_/nr ), .c(\U891/U1117_1_/nd ) );
    inv_2 \U891/U1117_1_/U3  ( .x(\b[1] ), .a(\U891/U1117_1_/n2 ) );
    nor3_1 \U891/U1117_2_/Unr  ( .x(\U891/U1117_2_/nr ), .a(i[2]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_2_/Und  ( .x(\U891/U1117_2_/nd ), .a(i[2]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_2_/U1  ( .x(\U891/U1117_2_/n2 ), .a(\U891/U1117_2_/n2 ), 
        .b(\U891/U1117_2_/nr ), .c(\U891/U1117_2_/nd ) );
    inv_2 \U891/U1117_2_/U3  ( .x(\b[2] ), .a(\U891/U1117_2_/n2 ) );
    nor3_1 \U891/U1117_3_/Unr  ( .x(\U891/U1117_3_/nr ), .a(i[3]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_3_/Und  ( .x(\U891/U1117_3_/nd ), .a(i[3]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_3_/U1  ( .x(\U891/U1117_3_/n2 ), .a(\U891/U1117_3_/n2 ), 
        .b(\U891/U1117_3_/nr ), .c(\U891/U1117_3_/nd ) );
    inv_2 \U891/U1117_3_/U3  ( .x(\b[3] ), .a(\U891/U1117_3_/n2 ) );
    inv_1 \U886/U1126/U3  ( .x(\U886/reset ), .a(nbReset) );
    nor3_1 \U886/U1128/U27  ( .x(\U886/U1128/nb ), .a(\U886/reset ), .b(\f[3] 
        ), .c(\f[2] ) );
    nor2_1 \U886/U1128/U26  ( .x(\U886/U1128/na ), .a(\f[1] ), .b(\f[0] ) );
    nand2_2 \U886/U1128/U29  ( .x(\U886/ackb ), .a(\U886/U1128/nb ), .b(
        \U886/U1128/na ) );
    nor2_1 \U886/U1108/U5  ( .x(\U886/nack ), .a(\U886/acka ), .b(\U886/ackb )
         );
    nor2_2 \U886/U914/U6  ( .x(nba), .a(\U886/acka ), .b(\U886/ackb ) );
    and4_1 \U886/U1127/U25  ( .x(\U886/U1127/n5 ), .a(\U886/U1127/n1 ), .b(
        \U886/U1127/n2 ), .c(\U886/U1127/n3 ), .d(\U886/U1127/n4 ) );
    inv_1 \U886/U1127/U1  ( .x(\U886/U1127/n1 ), .a(\e[3] ) );
    inv_1 \U886/U1127/U2  ( .x(\U886/U1127/n2 ), .a(\e[2] ) );
    inv_1 \U886/U1127/U3  ( .x(\U886/U1127/n3 ), .a(\e[1] ) );
    inv_1 \U886/U1127/U4  ( .x(\U886/U1127/n4 ), .a(\e[0] ) );
    inv_2 \U886/U1127/U5  ( .x(\U886/acka ), .a(\U886/U1127/n5 ) );
    ao222_2 \U886/U1121/U19/U1/U1  ( .x(fsela), .a(\U886/nack ), .b(fsel), .c(
        \U886/nack ), .d(fsela), .e(fsel), .f(fsela) );
    ao222_2 \U886/U1120/U19/U1/U1  ( .x(esela), .a(esel), .b(\U886/nack ), .c(
        esel), .d(esela), .e(\U886/nack ), .f(esela) );
    nor3_1 \U886/U1118_0_/Unr  ( .x(\U886/U1118_0_/nr ), .a(\b[0] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_0_/Und  ( .x(\U886/U1118_0_/nd ), .a(\b[0] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_0_/U1  ( .x(\U886/U1118_0_/n2 ), .a(\U886/U1118_0_/n2 ), 
        .b(\U886/U1118_0_/nr ), .c(\U886/U1118_0_/nd ) );
    inv_2 \U886/U1118_0_/U3  ( .x(\e[0] ), .a(\U886/U1118_0_/n2 ) );
    nor3_1 \U886/U1118_1_/Unr  ( .x(\U886/U1118_1_/nr ), .a(\b[1] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_1_/Und  ( .x(\U886/U1118_1_/nd ), .a(\b[1] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_1_/U1  ( .x(\U886/U1118_1_/n2 ), .a(\U886/U1118_1_/n2 ), 
        .b(\U886/U1118_1_/nr ), .c(\U886/U1118_1_/nd ) );
    inv_2 \U886/U1118_1_/U3  ( .x(\e[1] ), .a(\U886/U1118_1_/n2 ) );
    nor3_1 \U886/U1118_2_/Unr  ( .x(\U886/U1118_2_/nr ), .a(\b[2] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_2_/Und  ( .x(\U886/U1118_2_/nd ), .a(\b[2] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_2_/U1  ( .x(\U886/U1118_2_/n2 ), .a(\U886/U1118_2_/n2 ), 
        .b(\U886/U1118_2_/nr ), .c(\U886/U1118_2_/nd ) );
    inv_2 \U886/U1118_2_/U3  ( .x(\e[2] ), .a(\U886/U1118_2_/n2 ) );
    nor3_1 \U886/U1118_3_/Unr  ( .x(\U886/U1118_3_/nr ), .a(\b[3] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_3_/Und  ( .x(\U886/U1118_3_/nd ), .a(\b[3] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_3_/U1  ( .x(\U886/U1118_3_/n2 ), .a(\U886/U1118_3_/n2 ), 
        .b(\U886/U1118_3_/nr ), .c(\U886/U1118_3_/nd ) );
    inv_2 \U886/U1118_3_/U3  ( .x(\e[3] ), .a(\U886/U1118_3_/n2 ) );
    nor3_1 \U886/U1117_0_/Unr  ( .x(\U886/U1117_0_/nr ), .a(\b[0] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_0_/Und  ( .x(\U886/U1117_0_/nd ), .a(\b[0] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_0_/U1  ( .x(\U886/U1117_0_/n2 ), .a(\U886/U1117_0_/n2 ), 
        .b(\U886/U1117_0_/nr ), .c(\U886/U1117_0_/nd ) );
    inv_2 \U886/U1117_0_/U3  ( .x(\f[0] ), .a(\U886/U1117_0_/n2 ) );
    nor3_1 \U886/U1117_1_/Unr  ( .x(\U886/U1117_1_/nr ), .a(\b[1] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_1_/Und  ( .x(\U886/U1117_1_/nd ), .a(\b[1] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_1_/U1  ( .x(\U886/U1117_1_/n2 ), .a(\U886/U1117_1_/n2 ), 
        .b(\U886/U1117_1_/nr ), .c(\U886/U1117_1_/nd ) );
    inv_2 \U886/U1117_1_/U3  ( .x(\f[1] ), .a(\U886/U1117_1_/n2 ) );
    nor3_1 \U886/U1117_2_/Unr  ( .x(\U886/U1117_2_/nr ), .a(\b[2] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_2_/Und  ( .x(\U886/U1117_2_/nd ), .a(\b[2] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_2_/U1  ( .x(\U886/U1117_2_/n2 ), .a(\U886/U1117_2_/n2 ), 
        .b(\U886/U1117_2_/nr ), .c(\U886/U1117_2_/nd ) );
    inv_2 \U886/U1117_2_/U3  ( .x(\f[2] ), .a(\U886/U1117_2_/n2 ) );
    nor3_1 \U886/U1117_3_/Unr  ( .x(\U886/U1117_3_/nr ), .a(\b[3] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_3_/Und  ( .x(\U886/U1117_3_/nd ), .a(\b[3] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_3_/U1  ( .x(\U886/U1117_3_/n2 ), .a(\U886/U1117_3_/n2 ), 
        .b(\U886/U1117_3_/nr ), .c(\U886/U1117_3_/nd ) );
    inv_2 \U886/U1117_3_/U3  ( .x(\f[3] ), .a(\U886/U1117_3_/n2 ) );
    inv_1 \U884/U1126/U3  ( .x(\U884/reset ), .a(nbReset) );
    nor3_1 \U884/U1128/U27  ( .x(\U884/U1128/nb ), .a(\U884/reset ), .b(\d[3] 
        ), .c(\d[2] ) );
    nor2_1 \U884/U1128/U26  ( .x(\U884/U1128/na ), .a(\d[1] ), .b(\d[0] ) );
    nand2_2 \U884/U1128/U29  ( .x(\U884/ackb ), .a(\U884/U1128/nb ), .b(
        \U884/U1128/na ) );
    nor2_1 \U884/U1108/U5  ( .x(\U884/nack ), .a(\U884/acka ), .b(\U884/ackb )
         );
    nor2_2 \U884/U914/U6  ( .x(naa), .a(\U884/acka ), .b(\U884/ackb ) );
    and4_1 \U884/U1127/U25  ( .x(\U884/U1127/n5 ), .a(\U884/U1127/n1 ), .b(
        \U884/U1127/n2 ), .c(\U884/U1127/n3 ), .d(\U884/U1127/n4 ) );
    inv_1 \U884/U1127/U1  ( .x(\U884/U1127/n1 ), .a(\c[3] ) );
    inv_1 \U884/U1127/U2  ( .x(\U884/U1127/n2 ), .a(\c[2] ) );
    inv_1 \U884/U1127/U3  ( .x(\U884/U1127/n3 ), .a(\c[1] ) );
    inv_1 \U884/U1127/U4  ( .x(\U884/U1127/n4 ), .a(\c[0] ) );
    inv_2 \U884/U1127/U5  ( .x(\U884/acka ), .a(\U884/U1127/n5 ) );
    ao222_2 \U884/U1121/U19/U1/U1  ( .x(dsela), .a(\U884/nack ), .b(dsel), .c(
        \U884/nack ), .d(dsela), .e(dsel), .f(dsela) );
    ao222_2 \U884/U1120/U19/U1/U1  ( .x(csela), .a(csel), .b(\U884/nack ), .c(
        csel), .d(csela), .e(\U884/nack ), .f(csela) );
    nor3_1 \U884/U1118_0_/Unr  ( .x(\U884/U1118_0_/nr ), .a(\a[0] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_0_/Und  ( .x(\U884/U1118_0_/nd ), .a(\a[0] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_0_/U1  ( .x(\U884/U1118_0_/n2 ), .a(\U884/U1118_0_/n2 ), 
        .b(\U884/U1118_0_/nr ), .c(\U884/U1118_0_/nd ) );
    inv_2 \U884/U1118_0_/U3  ( .x(\c[0] ), .a(\U884/U1118_0_/n2 ) );
    nor3_1 \U884/U1118_1_/Unr  ( .x(\U884/U1118_1_/nr ), .a(\a[1] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_1_/Und  ( .x(\U884/U1118_1_/nd ), .a(\a[1] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_1_/U1  ( .x(\U884/U1118_1_/n2 ), .a(\U884/U1118_1_/n2 ), 
        .b(\U884/U1118_1_/nr ), .c(\U884/U1118_1_/nd ) );
    inv_2 \U884/U1118_1_/U3  ( .x(\c[1] ), .a(\U884/U1118_1_/n2 ) );
    nor3_1 \U884/U1118_2_/Unr  ( .x(\U884/U1118_2_/nr ), .a(\a[2] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_2_/Und  ( .x(\U884/U1118_2_/nd ), .a(\a[2] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_2_/U1  ( .x(\U884/U1118_2_/n2 ), .a(\U884/U1118_2_/n2 ), 
        .b(\U884/U1118_2_/nr ), .c(\U884/U1118_2_/nd ) );
    inv_2 \U884/U1118_2_/U3  ( .x(\c[2] ), .a(\U884/U1118_2_/n2 ) );
    nor3_1 \U884/U1118_3_/Unr  ( .x(\U884/U1118_3_/nr ), .a(\a[3] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_3_/Und  ( .x(\U884/U1118_3_/nd ), .a(\a[3] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_3_/U1  ( .x(\U884/U1118_3_/n2 ), .a(\U884/U1118_3_/n2 ), 
        .b(\U884/U1118_3_/nr ), .c(\U884/U1118_3_/nd ) );
    inv_2 \U884/U1118_3_/U3  ( .x(\c[3] ), .a(\U884/U1118_3_/n2 ) );
    nor3_1 \U884/U1117_0_/Unr  ( .x(\U884/U1117_0_/nr ), .a(\a[0] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_0_/Und  ( .x(\U884/U1117_0_/nd ), .a(\a[0] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_0_/U1  ( .x(\U884/U1117_0_/n2 ), .a(\U884/U1117_0_/n2 ), 
        .b(\U884/U1117_0_/nr ), .c(\U884/U1117_0_/nd ) );
    inv_2 \U884/U1117_0_/U3  ( .x(\d[0] ), .a(\U884/U1117_0_/n2 ) );
    nor3_1 \U884/U1117_1_/Unr  ( .x(\U884/U1117_1_/nr ), .a(\a[1] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_1_/Und  ( .x(\U884/U1117_1_/nd ), .a(\a[1] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_1_/U1  ( .x(\U884/U1117_1_/n2 ), .a(\U884/U1117_1_/n2 ), 
        .b(\U884/U1117_1_/nr ), .c(\U884/U1117_1_/nd ) );
    inv_2 \U884/U1117_1_/U3  ( .x(\d[1] ), .a(\U884/U1117_1_/n2 ) );
    nor3_1 \U884/U1117_2_/Unr  ( .x(\U884/U1117_2_/nr ), .a(\a[2] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_2_/Und  ( .x(\U884/U1117_2_/nd ), .a(\a[2] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_2_/U1  ( .x(\U884/U1117_2_/n2 ), .a(\U884/U1117_2_/n2 ), 
        .b(\U884/U1117_2_/nr ), .c(\U884/U1117_2_/nd ) );
    inv_2 \U884/U1117_2_/U3  ( .x(\d[2] ), .a(\U884/U1117_2_/n2 ) );
    nor3_1 \U884/U1117_3_/Unr  ( .x(\U884/U1117_3_/nr ), .a(\a[3] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_3_/Und  ( .x(\U884/U1117_3_/nd ), .a(\a[3] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_3_/U1  ( .x(\U884/U1117_3_/n2 ), .a(\U884/U1117_3_/n2 ), 
        .b(\U884/U1117_3_/nr ), .c(\U884/U1117_3_/nd ) );
    inv_2 \U884/U1117_3_/U3  ( .x(\d[3] ), .a(\U884/U1117_3_/n2 ) );
    nand2_1 \U888/U1128/U5  ( .x(\U888/s ), .a(\U888/r ), .b(\U888/nback ) );
    nand2_1 \U888/U1103/U5  ( .x(\U888/r ), .a(\U888/naack ), .b(\U888/s ) );
    inv_1 \U888/U1111/U3  ( .x(\U888/reset ), .a(nbReset) );
    inv_1 \U888/U1112/U3  ( .x(\U888/naack ), .a(esela) );
    nor2_1 \U888/U1127/U5  ( .x(\U888/nback ), .a(fsela), .b(\U888/reset ) );
    and2_2 \U888/U1129/U8  ( .x(esel), .a(\U888/nback ), .b(\U888/s ) );
    and2_2 \U888/U1124/U8  ( .x(fsel), .a(\U888/r ), .b(\U888/naack ) );
    nand2_1 \U887/U1128/U5  ( .x(\U887/s ), .a(\U887/r ), .b(\U887/nback ) );
    nand2_1 \U887/U1103/U5  ( .x(\U887/r ), .a(\U887/naack ), .b(\U887/s ) );
    inv_1 \U887/U1111/U3  ( .x(\U887/reset ), .a(nbReset) );
    inv_1 \U887/U1112/U3  ( .x(\U887/naack ), .a(csela) );
    nor2_1 \U887/U1127/U5  ( .x(\U887/nback ), .a(dsela), .b(\U887/reset ) );
    and2_2 \U887/U1129/U8  ( .x(csel), .a(\U887/nback ), .b(\U887/s ) );
    and2_2 \U887/U1124/U8  ( .x(dsel), .a(\U887/r ), .b(\U887/naack ) );
    nand2_1 \U885/U1128/U5  ( .x(\U885/s ), .a(\U885/r ), .b(\U885/nback ) );
    nand2_1 \U885/U1103/U5  ( .x(\U885/r ), .a(\U885/naack ), .b(\U885/s ) );
    inv_1 \U885/U1111/U3  ( .x(\U885/reset ), .a(nbReset) );
    inv_1 \U885/U1112/U3  ( .x(\U885/naack ), .a(asela) );
    nor2_1 \U885/U1127/U5  ( .x(\U885/nback ), .a(bsela), .b(\U885/reset ) );
    and2_2 \U885/U1129/U8  ( .x(asel), .a(\U885/nback ), .b(\U885/s ) );
    and2_2 \U885/U1124/U8  ( .x(bsel), .a(\U885/r ), .b(\U885/naack ) );
    nor3_1 \U877/U594/U7  ( .x(\U877/x ), .a(ol[7]), .b(\U877/reset ), .c(oh
        [7]) );
    nor3_1 \U877/U593/U7  ( .x(\U877/y ), .a(ol[6]), .b(\U877/reset ), .c(oh
        [6]) );
    inv_1 \U877/U604/U3  ( .x(\U877/reset ), .a(nbReset) );
    oa31_1 \U877/U590/U25/U1/Uclr  ( .x(\U877/U590/U25/U1/clr ), .a(net135), 
        .b(\cl[3] ), .c(\cl[1] ), .d(oh[6]) );
    oaoi211_1 \U877/U590/U25/U1/Uaoi  ( .x(\U877/U590/U25/U1/ob ), .a(\cl[3] ), 
        .b(\cl[1] ), .c(n1), .d(\U877/U590/U25/U1/clr ) );
    inv_2 \U877/U590/U25/U1/Ui  ( .x(oh[6]), .a(\U877/U590/U25/U1/ob ) );
    oa31_1 \U877/U589/U25/U1/Uclr  ( .x(\U877/U589/U25/U1/clr ), .a(net135), 
        .b(\cl[1] ), .c(\cl[0] ), .d(ol[7]) );
    oaoi211_1 \U877/U589/U25/U1/Uaoi  ( .x(\U877/U589/U25/U1/ob ), .a(\cl[1] ), 
        .b(\cl[0] ), .c(n1), .d(\U877/U589/U25/U1/clr ) );
    inv_2 \U877/U589/U25/U1/Ui  ( .x(ol[7]), .a(\U877/U589/U25/U1/ob ) );
    oa31_1 \U877/U588/U25/U1/Uclr  ( .x(\U877/U588/U25/U1/clr ), .a(net135), 
        .b(\cl[3] ), .c(\cl[2] ), .d(oh[7]) );
    oaoi211_1 \U877/U588/U25/U1/Uaoi  ( .x(\U877/U588/U25/U1/ob ), .a(\cl[3] ), 
        .b(\cl[2] ), .c(n1), .d(\U877/U588/U25/U1/clr ) );
    inv_2 \U877/U588/U25/U1/Ui  ( .x(oh[7]), .a(\U877/U588/U25/U1/ob ) );
    oa31_1 \U877/U591/U25/U1/Uclr  ( .x(\U877/U591/U25/U1/clr ), .a(net135), 
        .b(\cl[2] ), .c(\cl[0] ), .d(ol[6]) );
    oaoi211_1 \U877/U591/U25/U1/Uaoi  ( .x(\U877/U591/U25/U1/ob ), .a(\cl[2] ), 
        .b(\cl[0] ), .c(n1), .d(\U877/U591/U25/U1/clr ) );
    inv_2 \U877/U591/U25/U1/Ui  ( .x(ol[6]), .a(\U877/U591/U25/U1/ob ) );
    ao222_2 \U877/U592/U19/U1/U1  ( .x(ncla), .a(\U877/x ), .b(\U877/y ), .c(
        \U877/x ), .d(ncla), .e(\U877/y ), .f(ncla) );
    nor3_1 \U876/U594/U7  ( .x(\U876/x ), .a(ol[3]), .b(\U876/reset ), .c(oh
        [3]) );
    nor3_1 \U876/U593/U7  ( .x(\U876/y ), .a(ol[2]), .b(\U876/reset ), .c(oh
        [2]) );
    inv_1 \U876/U604/U3  ( .x(\U876/reset ), .a(nbReset) );
    oa31_1 \U876/U590/U25/U1/Uclr  ( .x(\U876/U590/U25/U1/clr ), .a(net135), 
        .b(\d[3] ), .c(\d[1] ), .d(oh[2]) );
    oaoi211_1 \U876/U590/U25/U1/Uaoi  ( .x(\U876/U590/U25/U1/ob ), .a(\d[3] ), 
        .b(\d[1] ), .c(n1), .d(\U876/U590/U25/U1/clr ) );
    inv_2 \U876/U590/U25/U1/Ui  ( .x(oh[2]), .a(\U876/U590/U25/U1/ob ) );
    oa31_1 \U876/U589/U25/U1/Uclr  ( .x(\U876/U589/U25/U1/clr ), .a(net135), 
        .b(\d[1] ), .c(\d[0] ), .d(ol[3]) );
    oaoi211_1 \U876/U589/U25/U1/Uaoi  ( .x(\U876/U589/U25/U1/ob ), .a(\d[1] ), 
        .b(\d[0] ), .c(n1), .d(\U876/U589/U25/U1/clr ) );
    inv_2 \U876/U589/U25/U1/Ui  ( .x(ol[3]), .a(\U876/U589/U25/U1/ob ) );
    oa31_1 \U876/U588/U25/U1/Uclr  ( .x(\U876/U588/U25/U1/clr ), .a(net135), 
        .b(\d[3] ), .c(\d[2] ), .d(oh[3]) );
    oaoi211_1 \U876/U588/U25/U1/Uaoi  ( .x(\U876/U588/U25/U1/ob ), .a(\d[3] ), 
        .b(\d[2] ), .c(n1), .d(\U876/U588/U25/U1/clr ) );
    inv_2 \U876/U588/U25/U1/Ui  ( .x(oh[3]), .a(\U876/U588/U25/U1/ob ) );
    oa31_1 \U876/U591/U25/U1/Uclr  ( .x(\U876/U591/U25/U1/clr ), .a(net135), 
        .b(\d[2] ), .c(\d[0] ), .d(ol[2]) );
    oaoi211_1 \U876/U591/U25/U1/Uaoi  ( .x(\U876/U591/U25/U1/ob ), .a(\d[2] ), 
        .b(\d[0] ), .c(n1), .d(\U876/U591/U25/U1/clr ) );
    inv_2 \U876/U591/U25/U1/Ui  ( .x(ol[2]), .a(\U876/U591/U25/U1/ob ) );
    ao222_2 \U876/U592/U19/U1/U1  ( .x(nda), .a(\U876/x ), .b(\U876/y ), .c(
        \U876/x ), .d(nda), .e(\U876/y ), .f(nda) );
    nor3_1 \U2/U594/U7  ( .x(\U2/x ), .a(ol[1]), .b(\U2/reset ), .c(oh[1]) );
    nor3_1 \U2/U593/U7  ( .x(\U2/y ), .a(ol[0]), .b(\U2/reset ), .c(oh[0]) );
    inv_1 \U2/U604/U3  ( .x(\U2/reset ), .a(nbReset) );
    oa31_1 \U2/U590/U25/U1/Uclr  ( .x(\U2/U590/U25/U1/clr ), .a(net135), .b(
        \f[3] ), .c(\f[1] ), .d(oh[0]) );
    oaoi211_1 \U2/U590/U25/U1/Uaoi  ( .x(\U2/U590/U25/U1/ob ), .a(\f[3] ), .b(
        \f[1] ), .c(n1), .d(\U2/U590/U25/U1/clr ) );
    inv_2 \U2/U590/U25/U1/Ui  ( .x(oh[0]), .a(\U2/U590/U25/U1/ob ) );
    oa31_1 \U2/U589/U25/U1/Uclr  ( .x(\U2/U589/U25/U1/clr ), .a(net135), .b(
        \f[1] ), .c(\f[0] ), .d(ol[1]) );
    oaoi211_1 \U2/U589/U25/U1/Uaoi  ( .x(\U2/U589/U25/U1/ob ), .a(\f[1] ), .b(
        \f[0] ), .c(n1), .d(\U2/U589/U25/U1/clr ) );
    inv_2 \U2/U589/U25/U1/Ui  ( .x(ol[1]), .a(\U2/U589/U25/U1/ob ) );
    oa31_1 \U2/U588/U25/U1/Uclr  ( .x(\U2/U588/U25/U1/clr ), .a(net135), .b(
        \f[3] ), .c(\f[2] ), .d(oh[1]) );
    oaoi211_1 \U2/U588/U25/U1/Uaoi  ( .x(\U2/U588/U25/U1/ob ), .a(\f[3] ), .b(
        \f[2] ), .c(n1), .d(\U2/U588/U25/U1/clr ) );
    inv_2 \U2/U588/U25/U1/Ui  ( .x(oh[1]), .a(\U2/U588/U25/U1/ob ) );
    oa31_1 \U2/U591/U25/U1/Uclr  ( .x(\U2/U591/U25/U1/clr ), .a(net135), .b(
        \f[2] ), .c(\f[0] ), .d(ol[0]) );
    oaoi211_1 \U2/U591/U25/U1/Uaoi  ( .x(\U2/U591/U25/U1/ob ), .a(\f[2] ), .b(
        \f[0] ), .c(n1), .d(\U2/U591/U25/U1/clr ) );
    inv_2 \U2/U591/U25/U1/Ui  ( .x(ol[0]), .a(\U2/U591/U25/U1/ob ) );
    ao222_2 \U2/U592/U19/U1/U1  ( .x(nfa), .a(\U2/x ), .b(\U2/y ), .c(\U2/x ), 
        .d(nfa), .e(\U2/y ), .f(nfa) );
    nor3_1 \U1/U594/U7  ( .x(\U1/x ), .a(ol[5]), .b(\U1/reset ), .c(oh[5]) );
    nor3_1 \U1/U593/U7  ( .x(\U1/y ), .a(ol[4]), .b(\U1/reset ), .c(oh[4]) );
    inv_1 \U1/U604/U3  ( .x(\U1/reset ), .a(nbReset) );
    oa31_1 \U1/U590/U25/U1/Uclr  ( .x(\U1/U590/U25/U1/clr ), .a(net135), .b(
        \e[3] ), .c(\e[1] ), .d(oh[4]) );
    oaoi211_1 \U1/U590/U25/U1/Uaoi  ( .x(\U1/U590/U25/U1/ob ), .a(\e[3] ), .b(
        \e[1] ), .c(n1), .d(\U1/U590/U25/U1/clr ) );
    inv_2 \U1/U590/U25/U1/Ui  ( .x(oh[4]), .a(\U1/U590/U25/U1/ob ) );
    oa31_1 \U1/U589/U25/U1/Uclr  ( .x(\U1/U589/U25/U1/clr ), .a(net135), .b(
        \e[1] ), .c(\e[0] ), .d(ol[5]) );
    oaoi211_1 \U1/U589/U25/U1/Uaoi  ( .x(\U1/U589/U25/U1/ob ), .a(\e[1] ), .b(
        \e[0] ), .c(n1), .d(\U1/U589/U25/U1/clr ) );
    inv_2 \U1/U589/U25/U1/Ui  ( .x(ol[5]), .a(\U1/U589/U25/U1/ob ) );
    oa31_1 \U1/U588/U25/U1/Uclr  ( .x(\U1/U588/U25/U1/clr ), .a(net135), .b(
        \e[3] ), .c(\e[2] ), .d(oh[5]) );
    oaoi211_1 \U1/U588/U25/U1/Uaoi  ( .x(\U1/U588/U25/U1/ob ), .a(\e[3] ), .b(
        \e[2] ), .c(n1), .d(\U1/U588/U25/U1/clr ) );
    inv_2 \U1/U588/U25/U1/Ui  ( .x(oh[5]), .a(\U1/U588/U25/U1/ob ) );
    oa31_1 \U1/U591/U25/U1/Uclr  ( .x(\U1/U591/U25/U1/clr ), .a(net135), .b(
        \e[2] ), .c(\e[0] ), .d(ol[4]) );
    oaoi211_1 \U1/U591/U25/U1/Uaoi  ( .x(\U1/U591/U25/U1/ob ), .a(\e[2] ), .b(
        \e[0] ), .c(n1), .d(\U1/U591/U25/U1/clr ) );
    inv_2 \U1/U591/U25/U1/Ui  ( .x(ol[4]), .a(\U1/U591/U25/U1/ob ) );
    ao222_2 \U1/U592/U19/U1/U1  ( .x(nea), .a(\U1/x ), .b(\U1/y ), .c(\U1/x ), 
        .d(nea), .e(\U1/y ), .f(nea) );
    and3_4 \U881/U20/U9  ( .x(nca), .a(\U881/nack[1] ), .b(\U881/nack[0] ), 
        .c(nbReset) );
    nor2_1 \U881/U18/U5  ( .x(\U881/nack[0] ), .a(\cl[3] ), .b(\cl[0] ) );
    nor2_1 \U881/U19/U5  ( .x(\U881/nack[1] ), .a(\cl[1] ), .b(\cl[2] ) );
    ao222_2 \U881/U15_0_/U19/U1/U1  ( .x(\cl[0] ), .a(\c[0] ), .b(ncla), .c(
        \c[0] ), .d(\cl[0] ), .e(ncla), .f(\cl[0] ) );
    ao222_2 \U881/U15_1_/U19/U1/U1  ( .x(\cl[1] ), .a(\c[1] ), .b(ncla), .c(
        \c[1] ), .d(\cl[1] ), .e(ncla), .f(\cl[1] ) );
    ao222_2 \U881/U15_2_/U19/U1/U1  ( .x(\cl[2] ), .a(\c[2] ), .b(ncla), .c(
        \c[2] ), .d(\cl[2] ), .e(ncla), .f(\cl[2] ) );
    ao222_2 \U881/U15_3_/U19/U1/U1  ( .x(\cl[3] ), .a(\c[3] ), .b(ncla), .c(
        \c[3] ), .d(\cl[3] ), .e(ncla), .f(\cl[3] ) );
    and2_5 U1 ( .x(n1), .a(nbReset), .b(noa) );
    and2_3 U2 ( .x(net135), .a(nbReset), .b(noa) );
endmodule


module chain_ic_ctrl_2 ( ack, candefer, eop, nstatack, pltxreq, routetxreq, 
    tok_ack, accept, candefer_ack, defer, eopack, lock, nReset, pltxack, 
    routetxack, tok_err, tok_ok );
input  [1:0] candefer_ack;
input  [1:0] lock;
input  accept, defer, eopack, nReset, pltxack, routetxack, tok_err, tok_ok;
output ack, candefer, eop, nstatack, pltxreq, routetxreq, tok_ack;
    wire net23, net25, net6, net19, net9, retry, net31, net24, net28, net27, 
        net7, net18, net13, net8, net11, net15, \U249/n5 , \U249/n1 , 
        \U249/n2 , \U249/n3 , \U249/n4 , txnodefer, net16, reset, net17, net29, 
        net12, txmaydefer, nlclear, net4, net22, net14, txlocked, net3, 
        \U286/U28/U1/clr , n1, \U286/U28/U1/set , \U285/U28/U1/clr , n2, 
        \U285/U28/U1/set , txunlocked, net2, txdone, net5, lockcleared, 
        \U262/U25/U1/clr , \U262/U25/U1/ob , \U284/U25/U1/clr , 
        \U284/U25/U1/ob , \U283/U25/U1/clr , net10, \U283/U25/U1/ob , net20, 
        \U289/Z , net21, \U287/Z , \U288/Z , \U149/nr , net30, \U149/nd , 
        \U149/n2 , \locked[0] , \locked[1] , lwrite, \U160/acb , net26, 
        \U160/U1/Z , \U136/nclear_latch , \U136/nwl , \U136/nulsense , 
        \U136/nlsense , \U136/nwh ;
    nand2_1 \U146/U5  ( .x(candefer), .a(net23), .b(net25) );
    or2_1 \U277/U12  ( .x(net6), .a(net19), .b(net9) );
    or2_1 \U264/U12  ( .x(retry), .a(net31), .b(net24) );
    or2_1 \U259/U12  ( .x(net28), .a(net27), .b(net7) );
    or2_1 \U140/U12  ( .x(net18), .a(net13), .b(net8) );
    or2_1 \U148/U12  ( .x(net11), .a(net15), .b(routetxack) );
    and4_1 \U249/U16  ( .x(\U249/n5 ), .a(\U249/n1 ), .b(\U249/n2 ), .c(
        \U249/n3 ), .d(\U249/n4 ) );
    inv_1 \U249/U1  ( .x(\U249/n1 ), .a(txnodefer) );
    inv_1 \U249/U2  ( .x(\U249/n2 ), .a(net16) );
    inv_1 \U249/U3  ( .x(\U249/n3 ), .a(net9) );
    inv_1 \U249/U4  ( .x(\U249/n4 ), .a(net19) );
    inv_1 \U249/U5  ( .x(ack), .a(\U249/n5 ) );
    nor3_2 \U40/U16  ( .x(nstatack), .a(net16), .b(reset), .c(retry) );
    nor3_2 \U275/U16  ( .x(net17), .a(net29), .b(reset), .c(tok_ack) );
    buf_3 \U290/U8  ( .x(net12), .a(txmaydefer) );
    nor2_1 \U154/U5  ( .x(nlclear), .a(net4), .b(net31) );
    or2_2 \U274/U12  ( .x(pltxreq), .a(net22), .b(net14) );
    or3_1 \U260/U12  ( .x(eop), .a(net31), .b(txlocked), .c(net4) );
    inv_1 \U147/U3  ( .x(net3), .a(net29) );
    inv_1 \U174/U3  ( .x(reset), .a(nReset) );
    aoai211_1 \U286/U28/U1/U1  ( .x(\U286/U28/U1/clr ), .a(net3), .b(n1), .c(
        net17), .d(net22) );
    nand3_1 \U286/U28/U1/U2  ( .x(\U286/U28/U1/set ), .a(net17), .b(net3), .c(
        n1) );
    nand2_2 \U286/U28/U1/U3  ( .x(net22), .a(\U286/U28/U1/clr ), .b(
        \U286/U28/U1/set ) );
    aoai211_1 \U285/U28/U1/U1  ( .x(\U285/U28/U1/clr ), .a(net3), .b(n2), .c(
        net17), .d(net14) );
    nand3_1 \U285/U28/U1/U2  ( .x(\U285/U28/U1/set ), .a(net17), .b(net3), .c(
        n2) );
    nand2_2 \U285/U28/U1/U3  ( .x(net14), .a(\U285/U28/U1/clr ), .b(
        \U285/U28/U1/set ) );
    ao222_1 \U254/U18/U1/U1  ( .x(net31), .a(defer), .b(txunlocked), .c(defer), 
        .d(net31), .e(txunlocked), .f(net31) );
    ao222_1 \U252/U18/U1/U1  ( .x(net19), .a(tok_err), .b(net12), .c(tok_err), 
        .d(net19), .e(net12), .f(net19) );
    ao222_1 \U276/U18/U1/U1  ( .x(net24), .a(txlocked), .b(defer), .c(txlocked
        ), .d(net24), .e(defer), .f(net24) );
    ao222_1 \U251/U18/U1/U1  ( .x(net9), .a(tok_ok), .b(net12), .c(tok_ok), 
        .d(net9), .e(net12), .f(net9) );
    ao222_1 \U235/U18/U1/U1  ( .x(tok_ack), .a(ack), .b(net2), .c(ack), .d(
        tok_ack), .e(net2), .f(tok_ack) );
    ao222_1 \U247/U18/U1/U1  ( .x(txnodefer), .a(txdone), .b(candefer_ack[0]), 
        .c(txdone), .d(txnodefer), .e(candefer_ack[0]), .f(txnodefer) );
    ao222_2 \U246/U19/U1/U1  ( .x(txlocked), .a(net14), .b(txdone), .c(net14), 
        .d(txlocked), .e(txdone), .f(txlocked) );
    ao222_2 \U245/U19/U1/U1  ( .x(txunlocked), .a(txdone), .b(net22), .c(
        txdone), .d(txunlocked), .e(net22), .f(txunlocked) );
    ao222_1 \U269/U18/U1/U1  ( .x(net2), .a(net28), .b(net18), .c(net28), .d(
        net2), .e(net18), .f(net2) );
    ao222_1 \U268/U18/U1/U1  ( .x(net5), .a(eopack), .b(lockcleared), .c(
        eopack), .d(net5), .e(lockcleared), .f(net5) );
    ao222_1 \U256/U18/U1/U1  ( .x(net4), .a(tok_err), .b(txunlocked), .c(
        tok_err), .d(net4), .e(txunlocked), .f(net4) );
    ao222_1 \U175/U18/U1/U1  ( .x(net29), .a(net2), .b(retry), .c(net2), .d(
        net29), .e(retry), .f(net29) );
    ao222_1 \U255/U18/U1/U1  ( .x(net8), .a(txlocked), .b(eopack), .c(txlocked
        ), .d(net8), .e(eopack), .f(net8) );
    ao222_2 \U248/U19/U1/U1  ( .x(txmaydefer), .a(candefer_ack[1]), .b(txdone), 
        .c(candefer_ack[1]), .d(txmaydefer), .e(txdone), .f(txmaydefer) );
    ao222_2 \U250/U19/U1/U1  ( .x(net16), .a(accept), .b(net12), .c(accept), 
        .d(net16), .e(net12), .f(net16) );
    oa31_1 \U262/U25/U1/Uclr  ( .x(\U262/U25/U1/clr ), .a(txunlocked), .b(net5
        ), .c(tok_ok), .d(net13) );
    oaoi211_1 \U262/U25/U1/Uaoi  ( .x(\U262/U25/U1/ob ), .a(net5), .b(tok_ok), 
        .c(txunlocked), .d(\U262/U25/U1/clr ) );
    inv_2 \U262/U25/U1/Ui  ( .x(net13), .a(\U262/U25/U1/ob ) );
    oa31_1 \U284/U25/U1/Uclr  ( .x(\U284/U25/U1/clr ), .a(txnodefer), .b(
        tok_ok), .c(tok_err), .d(net27) );
    oaoi211_1 \U284/U25/U1/Uaoi  ( .x(\U284/U25/U1/ob ), .a(tok_ok), .b(
        tok_err), .c(txnodefer), .d(\U284/U25/U1/clr ) );
    inv_2 \U284/U25/U1/Ui  ( .x(net27), .a(\U284/U25/U1/ob ) );
    oa31_1 \U283/U25/U1/Uclr  ( .x(\U283/U25/U1/clr ), .a(net10), .b(net6), 
        .c(retry), .d(net7) );
    oaoi211_1 \U283/U25/U1/Uaoi  ( .x(\U283/U25/U1/ob ), .a(net6), .b(retry), 
        .c(net10), .d(\U283/U25/U1/clr ) );
    inv_2 \U283/U25/U1/Ui  ( .x(net7), .a(\U283/U25/U1/ob ) );
    aoi21_1 \U289/U30/U1/U1  ( .x(net20), .a(\U289/Z ), .b(net16), .c(net12)
         );
    inv_1 \U289/U30/U1/U2  ( .x(\U289/Z ), .a(net20) );
    aoi21_1 \U287/U30/U1/U1  ( .x(net21), .a(\U287/Z ), .b(accept), .c(net12)
         );
    inv_1 \U287/U30/U1/U2  ( .x(\U287/Z ), .a(net21) );
    aoi222_1 \U288/U30/U1  ( .x(net10), .a(net20), .b(net21), .c(net20), .d(
        \U288/Z ), .e(net21), .f(\U288/Z ) );
    inv_1 \U288/U30/Uinv  ( .x(\U288/Z ), .a(net10) );
    nor3_1 \U149/Unr  ( .x(\U149/nr ), .a(pltxack), .b(net11), .c(net30) );
    nand3_1 \U149/Und  ( .x(\U149/nd ), .a(pltxack), .b(net11), .c(net30) );
    oa21_1 \U149/U1  ( .x(\U149/n2 ), .a(\U149/n2 ), .b(\U149/nr ), .c(
        \U149/nd ) );
    inv_2 \U149/U3  ( .x(txdone), .a(\U149/n2 ) );
    inv_1 \U133/U618/U3  ( .x(net23), .a(net15) );
    inv_1 \U133/U617/U3  ( .x(net25), .a(routetxreq) );
    ao23_1 \U133/U616/U21/U1/U1  ( .x(routetxreq), .a(pltxreq), .b(routetxreq), 
        .c(pltxreq), .d(\locked[0] ), .e(net23) );
    ao23_1 \U133/U615/U21/U1/U1  ( .x(net15), .a(pltxreq), .b(net15), .c(
        pltxreq), .d(\locked[1] ), .e(net25) );
    and2_1 \U160/U2/U8  ( .x(lwrite), .a(candefer), .b(\U160/acb ) );
    nor2_1 \U160/U3/U5  ( .x(net30), .a(\U160/acb ), .b(net26) );
    oai21_1 \U160/U1/U30/U1/U1  ( .x(\U160/acb ), .a(\U160/U1/Z ), .b(net26), 
        .c(candefer) );
    inv_1 \U160/U1/U30/U1/U2  ( .x(\U160/U1/Z ), .a(\U160/acb ) );
    nand3_2 \U136/U48/U16  ( .x(\locked[0] ), .a(\locked[1] ), .b(
        \U136/nclear_latch ), .c(\U136/nwl ) );
    nor2_0 \U136/U36/U5  ( .x(\U136/nulsense ), .a(\locked[1] ), .b(\U136/nwl 
        ) );
    nor2_0 \U136/U37/U5  ( .x(\U136/nlsense ), .a(\U136/nwh ), .b(\locked[0] )
         );
    and2_1 \U136/U76/U8  ( .x(\U136/nclear_latch ), .a(nReset), .b(nlclear) );
    nor2_1 \U136/U77/U5  ( .x(lockcleared), .a(nlclear), .b(\locked[1] ) );
    nand2_1 \U136/U14/U5  ( .x(\U136/nwl ), .a(lwrite), .b(n2) );
    nand2_1 \U136/U15/U5  ( .x(\U136/nwh ), .a(n1), .b(lwrite) );
    nand2_2 \U136/U47/U5  ( .x(\locked[1] ), .a(\U136/nwh ), .b(\locked[0] )
         );
    or2_4 \U136/U35/U12  ( .x(net26), .a(\U136/nlsense ), .b(\U136/nulsense )
         );
    buf_1 U1 ( .x(n1), .a(lock[1]) );
    buf_1 U2 ( .x(n2), .a(lock[0]) );
endmodule


module chain_selement_ga_53 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_54 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_55 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_56 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_60 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_57 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_61 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_58 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_59 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_52 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_dr8bit_completion_54 ( o, i );
input  [15:0] i;
output o;
    wire \nx[0] , \nx[1] , \nx[2] , \nx[3] , \ny[0] , \ny[1] , \ny[2] , 
        \ny[3] , y, x, \U6/Z , \U3/net3 , \U3/U20/Z , \U3/net2 , \U3/U21/Z , 
        \U3/U19/Z , \U5/net3 , \U5/U20/Z , \U5/net2 , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_55 ( o, i );
input  [15:0] i;
output o;
    wire \nx[0] , \nx[1] , \nx[2] , \nx[3] , \ny[0] , \ny[1] , \ny[2] , 
        \ny[3] , y, x, \U6/Z , \U3/net3 , \U3/U20/Z , \U3/net2 , \U3/U21/Z , 
        \U3/U19/Z , \U5/net3 , \U5/U20/Z , \U5/net2 , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_32 ( o, i );
input  [15:0] i;
output o;
    wire \nx[0] , \nx[1] , \nx[2] , \nx[3] , \ny[0] , \ny[1] , \ny[2] , 
        \ny[3] , y, x, \U6/Z , \U3/net3 , \U3/U20/Z , \U3/net2 , \U3/U21/Z , 
        \U3/U19/Z , \U5/net3 , \U5/U20/Z , \U5/net2 , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_35 ( o, i );
input  [15:0] i;
output o;
    wire \nx[0] , \nx[1] , \nx[2] , \nx[3] , \ny[0] , \ny[1] , \ny[2] , 
        \ny[3] , y, x, \U6/Z , \U3/net3 , \U3/U20/Z , \U3/net2 , \U3/U21/Z , 
        \U3/U19/Z , \U5/net3 , \U5/U20/Z , \U5/net2 , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_34 ( o, i );
input  [15:0] i;
output o;
    wire \nx[0] , \nx[1] , \nx[2] , \nx[3] , \ny[0] , \ny[1] , \ny[2] , 
        \ny[3] , y, x, \U6/Z , \U3/net3 , \U3/U20/Z , \U3/net2 , \U3/U21/Z , 
        \U3/U19/Z , \U5/net3 , \U5/U20/Z , \U5/net2 , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_33 ( o, i );
input  [15:0] i;
output o;
    wire \nx[0] , \nx[1] , \nx[2] , \nx[3] , \ny[0] , \ny[1] , \ny[2] , 
        \ny[3] , y, x, \U6/Z , \U3/net3 , \U3/U20/Z , \U3/net2 , \U3/U21/Z , 
        \U3/U19/Z , \U5/net3 , \U5/U20/Z , \U5/net2 , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr32bit_completion_6 ( o, i );
input  [63:0] i;
output o;
    wire \cd[3] , \cd[2] , \cd[1] , \cd[0] , ny, \U16/Z , nx, \U6/Z , \U15/Z ;
    chain_dr8bit_completion_32 U11 ( .o(\cd[3] ), .i({i[63], i[62], i[61], 
        i[60], i[59], i[58], i[57], i[56], i[31], i[30], i[29], i[28], i[27], 
        i[26], i[25], i[24]}) );
    chain_dr8bit_completion_35 U14 ( .o(\cd[2] ), .i({i[55], i[54], i[53], 
        i[52], i[51], i[50], i[49], i[48], i[23], i[22], i[21], i[20], i[19], 
        i[18], i[17], i[16]}) );
    chain_dr8bit_completion_34 U13 ( .o(\cd[1] ), .i({i[47], i[46], i[45], 
        i[44], i[43], i[42], i[41], i[40], i[15], i[14], i[13], i[12], i[11], 
        i[10], i[9], i[8]}) );
    chain_dr8bit_completion_33 U12 ( .o(\cd[0] ), .i({i[39], i[38], i[37], 
        i[36], i[35], i[34], i[33], i[32], i[7], i[6], i[5], i[4], i[3], i[2], 
        i[1], i[0]}) );
    aoi222_1 \U16/U30/U1  ( .x(ny), .a(\cd[0] ), .b(\cd[1] ), .c(\cd[0] ), .d(
        \U16/Z ), .e(\cd[1] ), .f(\U16/Z ) );
    inv_1 \U16/U30/Uinv  ( .x(\U16/Z ), .a(ny) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(ny), .b(nx), .c(ny), .d(\U6/Z ), .e(nx), 
        .f(\U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U15/U30/U1  ( .x(nx), .a(\cd[3] ), .b(\cd[2] ), .c(\cd[3] ), .d(
        \U15/Z ), .e(\cd[2] ), .f(\U15/Z ) );
    inv_1 \U15/U30/Uinv  ( .x(\U15/Z ), .a(nx) );
endmodule


module chain_dr8bit_completion_36 ( o, i );
input  [15:0] i;
output o;
    wire \nx[0] , \nx[1] , \nx[2] , \nx[3] , \ny[0] , \ny[1] , \ny[2] , 
        \ny[3] , y, x, \U6/Z , \U3/net3 , \U3/U20/Z , \U3/net2 , \U3/U21/Z , 
        \U3/U19/Z , \U5/net3 , \U5/U20/Z , \U5/net2 , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_39 ( o, i );
input  [15:0] i;
output o;
    wire \nx[0] , \nx[1] , \nx[2] , \nx[3] , \ny[0] , \ny[1] , \ny[2] , 
        \ny[3] , y, x, \U6/Z , \U3/net3 , \U3/U20/Z , \U3/net2 , \U3/U21/Z , 
        \U3/U19/Z , \U5/net3 , \U5/U20/Z , \U5/net2 , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_38 ( o, i );
input  [15:0] i;
output o;
    wire \nx[0] , \nx[1] , \nx[2] , \nx[3] , \ny[0] , \ny[1] , \ny[2] , 
        \ny[3] , y, x, \U6/Z , \U3/net3 , \U3/U20/Z , \U3/net2 , \U3/U21/Z , 
        \U3/U19/Z , \U5/net3 , \U5/U20/Z , \U5/net2 , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_37 ( o, i );
input  [15:0] i;
output o;
    wire \nx[0] , \nx[1] , \nx[2] , \nx[3] , \ny[0] , \ny[1] , \ny[2] , 
        \ny[3] , y, x, \U6/Z , \U3/net3 , \U3/U20/Z , \U3/net2 , \U3/U21/Z , 
        \U3/U19/Z , \U5/net3 , \U5/U20/Z , \U5/net2 , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr32bit_completion_7 ( o, i );
input  [63:0] i;
output o;
    wire \cd[3] , \cd[2] , \cd[1] , \cd[0] , ny, \U16/Z , nx, \U6/Z , \U15/Z ;
    chain_dr8bit_completion_36 U11 ( .o(\cd[3] ), .i({i[63], i[62], i[61], 
        i[60], i[59], i[58], i[57], i[56], i[31], i[30], i[29], i[28], i[27], 
        i[26], i[25], i[24]}) );
    chain_dr8bit_completion_39 U14 ( .o(\cd[2] ), .i({i[55], i[54], i[53], 
        i[52], i[51], i[50], i[49], i[48], i[23], i[22], i[21], i[20], i[19], 
        i[18], i[17], i[16]}) );
    chain_dr8bit_completion_38 U13 ( .o(\cd[1] ), .i({i[47], i[46], i[45], 
        i[44], i[43], i[42], i[41], i[40], i[15], i[14], i[13], i[12], i[11], 
        i[10], i[9], i[8]}) );
    chain_dr8bit_completion_37 U12 ( .o(\cd[0] ), .i({i[39], i[38], i[37], 
        i[36], i[35], i[34], i[33], i[32], i[7], i[6], i[5], i[4], i[3], i[2], 
        i[1], i[0]}) );
    aoi222_1 \U16/U30/U1  ( .x(ny), .a(\cd[0] ), .b(\cd[1] ), .c(\cd[0] ), .d(
        \U16/Z ), .e(\cd[1] ), .f(\U16/Z ) );
    inv_1 \U16/U30/Uinv  ( .x(\U16/Z ), .a(ny) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(ny), .b(nx), .c(ny), .d(\U6/Z ), .e(nx), 
        .f(\U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U15/U30/U1  ( .x(nx), .a(\cd[3] ), .b(\cd[2] ), .c(\cd[3] ), .d(
        \U15/Z ), .e(\cd[2] ), .f(\U15/Z ) );
    inv_1 \U15/U30/Uinv  ( .x(\U15/Z ), .a(nx) );
endmodule


module chain_icmux_2 ( ack, chainh, chainl, sendack, addr, col, itag, lock, 
    nReset, nia, pred, rnw, sendreq, seq, size, wd );
output [7:0] chainh;
output [7:0] chainl;
input  [63:0] addr;
input  [5:0] col;
input  [9:0] itag;
input  [1:0] lock;
input  [1:0] pred;
input  [1:0] rnw;
input  [1:0] seq;
input  [3:0] size;
input  [63:0] wd;
input  nReset, nia, sendreq;
output ack, sendack;
    wire net152, net146, net148, n1, net156, \bs[1] , net138, net160, \bs[2] , 
        net168, \bs[3] , net172, \bs[7] , net164, net132, \bs[4] , net289, 
        \bs[8] , net180, \bs[5] , net176, \bs[6] , \bs[0] , \hdr[4] , net185, 
        net187, net189, net191, net293, net131, \net246[15] , net265, 
        \net246[14] , \net246[13] , \net246[12] , \net246[11] , \net246[10] , 
        \net246[9] , \net246[8] , \net246[7] , \net246[6] , \net246[5] , 
        \net246[4] , \net246[3] , \net246[2] , \net246[1] , \net246[0] , 
        \net243[15] , net263, \net243[14] , \net243[13] , \net243[12] , 
        \net243[11] , \net243[10] , \net243[9] , \net243[8] , \net243[7] , 
        \net243[6] , \net243[5] , \net243[4] , \net243[3] , \net243[2] , 
        \net243[1] , \net243[0] , \net240[15] , net267, \net240[14] , 
        \net240[13] , \net240[12] , \net240[11] , \net240[10] , \net240[9] , 
        \net240[8] , \net240[7] , \net240[6] , \net240[5] , \net240[4] , 
        \net240[3] , \net240[2] , \net240[1] , \net240[0] , \net237[15] , 
        net269, \net237[14] , \net237[13] , \net237[12] , \net237[11] , 
        \net237[10] , \net237[9] , \net237[8] , \net237[7] , \net237[6] , 
        \net237[5] , \net237[2] , \net237[1] , \net237[0] , \net234[15] , 
        net259, \net234[14] , \net234[13] , \net234[12] , \net234[11] , 
        \net234[10] , \net234[9] , \net234[8] , \net234[7] , \net234[6] , 
        \net234[5] , \net234[4] , \net234[3] , \net234[2] , \net234[1] , 
        \net234[0] , \net231[15] , net253, \net231[14] , \net231[13] , 
        \net231[12] , \net231[11] , \net231[10] , \net231[9] , \net231[8] , 
        \net231[7] , \net231[6] , \net231[5] , \net231[4] , \net231[3] , 
        \net231[2] , \net231[1] , \net231[0] , \net228[15] , net255, 
        \net228[14] , \net228[13] , \net228[12] , \net228[11] , \net228[10] , 
        \net228[9] , \net228[8] , \net228[7] , \net228[6] , \net228[5] , 
        \net228[4] , \net228[3] , \net228[2] , \net228[1] , \net228[0] , 
        \net225[15] , net251, \net225[14] , \net225[13] , \net225[12] , 
        \net225[11] , \net225[10] , \net225[9] , \net225[8] , \net225[7] , 
        \net225[6] , \net225[5] , \net225[4] , \net225[3] , \net225[2] , 
        \net225[1] , \net225[0] , \net222[15] , net261, \net222[14] , 
        \net222[13] , \net222[12] , \net222[11] , \net222[10] , \net222[9] , 
        \net222[8] , \net222[7] , \net222[6] , \net222[5] , \net222[4] , 
        \net222[3] , \net222[2] , \net222[1] , \net222[0] , \net219[15] , 
        net249, \net219[14] , \net219[13] , \net219[12] , \net219[11] , 
        \net219[10] , \net219[9] , \net219[8] , \net219[7] , \net219[6] , 
        \net219[5] , \net219[4] , \net219[3] , \net219[2] , \net219[1] , 
        \net219[0] , \U40_0_/n3 , \U40_0_/n4 , \net217[15] , \U40_0_/n5 , 
        \U40_1_/n3 , \U40_1_/n4 , \net217[14] , \U40_1_/n5 , \U40_2_/n3 , 
        \U40_2_/n4 , \net217[13] , \U40_2_/n5 , \U40_3_/n3 , \U40_3_/n4 , 
        \net217[12] , \U40_3_/n5 , \U40_4_/n3 , \U40_4_/n4 , \net217[11] , 
        \U40_4_/n5 , \U40_5_/n3 , \U40_5_/n4 , \net217[10] , \U40_5_/n5 , 
        \U40_6_/n3 , \U40_6_/n4 , \net217[9] , \U40_6_/n5 , \U40_7_/n3 , 
        \U40_7_/n4 , \net217[8] , \U40_7_/n5 , \U40_8_/n3 , \U40_8_/n4 , 
        \net217[7] , \U40_8_/n5 , \U40_9_/n3 , \U40_9_/n4 , \net217[6] , 
        \U40_9_/n5 , \U40_10_/n3 , \U40_10_/n4 , \net217[5] , \U40_10_/n5 , 
        \U40_11_/n3 , \U40_11_/n4 , \net217[4] , \U40_11_/n5 , \U40_12_/n3 , 
        \U40_12_/n4 , \net217[3] , \U40_12_/n5 , \U40_13_/n3 , \U40_13_/n4 , 
        \net217[2] , \U40_13_/n5 , \U40_14_/n3 , \U40_14_/n4 , \net217[1] , 
        \U40_14_/n5 , \U40_15_/n3 , \U40_15_/n4 , \net217[0] , \U40_15_/n5 , 
        \U14_0_/n5 , \U14_0_/n1 , \U14_0_/n2 , \U14_0_/n3 , \U14_0_/n4 , 
        \net212[15] , \U14_1_/n5 , \U14_1_/n1 , \U14_1_/n2 , \U14_1_/n3 , 
        \U14_1_/n4 , \net212[14] , \U14_2_/n5 , \U14_2_/n1 , \U14_2_/n2 , 
        \U14_2_/n3 , \U14_2_/n4 , \net212[13] , \U14_3_/n5 , \U14_3_/n1 , 
        \U14_3_/n2 , \U14_3_/n3 , \U14_3_/n4 , \net212[12] , \U14_4_/n5 , 
        \U14_4_/n1 , \U14_4_/n2 , \U14_4_/n3 , \U14_4_/n4 , \net212[11] , 
        \U14_5_/n5 , \U14_5_/n1 , \U14_5_/n2 , \U14_5_/n3 , \U14_5_/n4 , 
        \net212[10] , \U14_6_/n5 , \U14_6_/n1 , \U14_6_/n2 , \U14_6_/n3 , 
        \U14_6_/n4 , \net212[9] , \U14_7_/n5 , \U14_7_/n1 , \U14_7_/n2 , 
        \U14_7_/n3 , \U14_7_/n4 , \net212[8] , \U14_8_/n5 , \U14_8_/n1 , 
        \U14_8_/n2 , \U14_8_/n3 , \U14_8_/n4 , \net212[7] , \U14_9_/n5 , 
        \U14_9_/n1 , \U14_9_/n2 , \U14_9_/n3 , \U14_9_/n4 , \net212[6] , 
        \U14_10_/n5 , \U14_10_/n1 , \U14_10_/n2 , \U14_10_/n3 , \U14_10_/n4 , 
        \net212[5] , \U14_11_/n1 , \U14_11_/n2 , \U14_11_/n4 , \net212[4] , 
        \U14_11_/n5 , \U14_12_/n1 , \U14_12_/n2 , \U14_12_/n4 , \net212[3] , 
        \U14_12_/n5 , \U14_13_/n5 , \U14_13_/n1 , \U14_13_/n2 , \U14_13_/n3 , 
        \U14_13_/n4 , \net212[2] , \U14_14_/n5 , \U14_14_/n1 , \U14_14_/n2 , 
        \U14_14_/n3 , \U14_14_/n4 , \net212[1] , \U14_15_/n5 , \U14_15_/n1 , 
        \U14_15_/n2 , \U14_15_/n3 , \U14_15_/n4 , \net212[0] , \U91_0_/n5 , 
        \U91_0_/n1 , \U91_0_/n2 , \U91_0_/n3 , \U91_0_/n4 , \net207[15] , 
        \U91_1_/n5 , \U91_1_/n1 , \U91_1_/n2 , \U91_1_/n3 , \U91_1_/n4 , 
        \net207[14] , \U91_2_/n5 , \U91_2_/n1 , \U91_2_/n2 , \U91_2_/n3 , 
        \U91_2_/n4 , \net207[13] , \U91_3_/n5 , \U91_3_/n1 , \U91_3_/n2 , 
        \U91_3_/n3 , \U91_3_/n4 , \net207[12] , \U91_4_/n5 , \U91_4_/n1 , 
        \U91_4_/n2 , \U91_4_/n3 , \U91_4_/n4 , \net207[11] , \U91_5_/n5 , 
        \U91_5_/n1 , \U91_5_/n2 , \U91_5_/n3 , \U91_5_/n4 , \net207[10] , 
        \U91_6_/n5 , \U91_6_/n1 , \U91_6_/n2 , \U91_6_/n3 , \U91_6_/n4 , 
        \net207[9] , \U91_7_/n5 , \U91_7_/n1 , \U91_7_/n2 , \U91_7_/n3 , 
        \U91_7_/n4 , \net207[8] , \U91_8_/n5 , \U91_8_/n1 , \U91_8_/n2 , 
        \U91_8_/n3 , \U91_8_/n4 , \net207[7] , \U91_9_/n5 , \U91_9_/n1 , 
        \U91_9_/n2 , \U91_9_/n3 , \U91_9_/n4 , \net207[6] , \U91_10_/n5 , 
        \U91_10_/n1 , \U91_10_/n2 , \U91_10_/n3 , \U91_10_/n4 , \net207[5] , 
        \U91_11_/n5 , \U91_11_/n1 , \U91_11_/n2 , \U91_11_/n3 , \U91_11_/n4 , 
        \net207[4] , \U91_12_/n5 , \U91_12_/n1 , \U91_12_/n2 , \U91_12_/n3 , 
        \U91_12_/n4 , \net207[3] , \U91_13_/n5 , \U91_13_/n1 , \U91_13_/n2 , 
        \U91_13_/n3 , \U91_13_/n4 , \net207[2] , \U91_14_/n5 , \U91_14_/n1 , 
        \U91_14_/n2 , \U91_14_/n3 , \U91_14_/n4 , \net207[1] , \U91_15_/n5 , 
        \U91_15_/n1 , \U91_15_/n2 , \U91_15_/n3 , \U91_15_/n4 , \net207[0] , 
        net198, net136, \U151/Z , \U148/U21/nr , \U148/U21/nd , \U148/U21/n2 ;
    chain_selement_ga_53 U163 ( .Aa(net152), .Br(net146), .Ar(net148), .Ba(n1)
         );
    chain_selement_ga_54 U164 ( .Aa(net156), .Br(\bs[1] ), .Ar(net152), .Ba(
        net138) );
    chain_selement_ga_55 U165 ( .Aa(net160), .Br(\bs[2] ), .Ar(net156), .Ba(n1
        ) );
    chain_selement_ga_56 U166 ( .Aa(net168), .Br(\bs[3] ), .Ar(net160), .Ba(
        net138) );
    chain_selement_ga_60 U170 ( .Aa(net172), .Br(\bs[7] ), .Ar(net164), .Ba(
        net138) );
    chain_selement_ga_57 U167 ( .Aa(net132), .Br(\bs[4] ), .Ar(net168), .Ba(
        net138) );
    chain_selement_ga_61 U171 ( .Aa(net289), .Br(\bs[8] ), .Ar(net172), .Ba(
        net138) );
    chain_selement_ga_58 U168 ( .Aa(net180), .Br(\bs[5] ), .Ar(net176), .Ba(
        net138) );
    chain_selement_ga_59 U169 ( .Aa(net164), .Br(\bs[6] ), .Ar(net180), .Ba(n1
        ) );
    chain_selement_ga_52 U161 ( .Aa(net148), .Br(\bs[0] ), .Ar(\hdr[4] ), .Ba(
        n1) );
    chain_dr8bit_completion_54 U119 ( .o(net185), .i({col[5], col[4], col[3], 
        itag[9], itag[8], itag[7], itag[6], itag[5], col[2], col[1], col[0], 
        itag[4], itag[3], itag[2], itag[1], itag[0]}) );
    chain_dr8bit_completion_55 U147 ( .o(net187), .i({size[3], size[2], rnw[1], 
        1'b0, 1'b0, lock[1], pred[1], seq[1], size[1], size[0], rnw[0], 
        \hdr[4] , \hdr[4] , lock[0], pred[0], seq[0]}) );
    chain_dr32bit_completion_6 U117 ( .o(net189), .i(wd) );
    chain_dr32bit_completion_7 U118 ( .o(net191), .i(addr) );
    or2_4 \U122/U12  ( .x(net293), .a(net189), .b(net131) );
    or2_4 \U53/U12  ( .x(sendack), .a(net131), .b(net289) );
    and2_1 \U32_0_/U8  ( .x(\net246[15] ), .a(itag[0]), .b(net265) );
    and2_1 \U32_1_/U8  ( .x(\net246[14] ), .a(itag[1]), .b(net265) );
    and2_1 \U32_2_/U8  ( .x(\net246[13] ), .a(itag[2]), .b(net265) );
    and2_1 \U32_3_/U8  ( .x(\net246[12] ), .a(itag[3]), .b(net265) );
    and2_1 \U32_4_/U8  ( .x(\net246[11] ), .a(itag[4]), .b(net265) );
    and2_1 \U32_5_/U8  ( .x(\net246[10] ), .a(col[0]), .b(net265) );
    and2_1 \U32_6_/U8  ( .x(\net246[9] ), .a(col[1]), .b(net265) );
    and2_1 \U32_7_/U8  ( .x(\net246[8] ), .a(col[2]), .b(net265) );
    and2_1 \U32_8_/U8  ( .x(\net246[7] ), .a(itag[5]), .b(net265) );
    and2_1 \U32_9_/U8  ( .x(\net246[6] ), .a(itag[6]), .b(net265) );
    and2_1 \U32_10_/U8  ( .x(\net246[5] ), .a(itag[7]), .b(net265) );
    and2_1 \U32_11_/U8  ( .x(\net246[4] ), .a(itag[8]), .b(net265) );
    and2_1 \U32_12_/U8  ( .x(\net246[3] ), .a(itag[9]), .b(net265) );
    and2_1 \U32_13_/U8  ( .x(\net246[2] ), .a(col[3]), .b(net265) );
    and2_1 \U32_14_/U8  ( .x(\net246[1] ), .a(col[4]), .b(net265) );
    and2_1 \U32_15_/U8  ( .x(\net246[0] ), .a(col[5]), .b(net265) );
    and2_1 \U76_0_/U8  ( .x(\net243[15] ), .a(wd[8]), .b(net263) );
    and2_1 \U76_1_/U8  ( .x(\net243[14] ), .a(wd[9]), .b(net263) );
    and2_1 \U76_2_/U8  ( .x(\net243[13] ), .a(wd[10]), .b(net263) );
    and2_1 \U76_3_/U8  ( .x(\net243[12] ), .a(wd[11]), .b(net263) );
    and2_1 \U76_4_/U8  ( .x(\net243[11] ), .a(wd[12]), .b(net263) );
    and2_1 \U76_5_/U8  ( .x(\net243[10] ), .a(wd[13]), .b(net263) );
    and2_1 \U76_6_/U8  ( .x(\net243[9] ), .a(wd[14]), .b(net263) );
    and2_1 \U76_7_/U8  ( .x(\net243[8] ), .a(wd[15]), .b(net263) );
    and2_1 \U76_8_/U8  ( .x(\net243[7] ), .a(wd[40]), .b(net263) );
    and2_1 \U76_9_/U8  ( .x(\net243[6] ), .a(wd[41]), .b(net263) );
    and2_1 \U76_10_/U8  ( .x(\net243[5] ), .a(wd[42]), .b(net263) );
    and2_1 \U76_11_/U8  ( .x(\net243[4] ), .a(wd[43]), .b(net263) );
    and2_1 \U76_12_/U8  ( .x(\net243[3] ), .a(wd[44]), .b(net263) );
    and2_1 \U76_13_/U8  ( .x(\net243[2] ), .a(wd[45]), .b(net263) );
    and2_1 \U76_14_/U8  ( .x(\net243[1] ), .a(wd[46]), .b(net263) );
    and2_1 \U76_15_/U8  ( .x(\net243[0] ), .a(wd[47]), .b(net263) );
    and2_1 \U80_0_/U8  ( .x(\net240[15] ), .a(wd[16]), .b(net267) );
    and2_1 \U80_1_/U8  ( .x(\net240[14] ), .a(wd[17]), .b(net267) );
    and2_1 \U80_2_/U8  ( .x(\net240[13] ), .a(wd[18]), .b(net267) );
    and2_1 \U80_3_/U8  ( .x(\net240[12] ), .a(wd[19]), .b(net267) );
    and2_1 \U80_4_/U8  ( .x(\net240[11] ), .a(wd[20]), .b(net267) );
    and2_1 \U80_5_/U8  ( .x(\net240[10] ), .a(wd[21]), .b(net267) );
    and2_1 \U80_6_/U8  ( .x(\net240[9] ), .a(wd[22]), .b(net267) );
    and2_1 \U80_7_/U8  ( .x(\net240[8] ), .a(wd[23]), .b(net267) );
    and2_1 \U80_8_/U8  ( .x(\net240[7] ), .a(wd[48]), .b(net267) );
    and2_1 \U80_9_/U8  ( .x(\net240[6] ), .a(wd[49]), .b(net267) );
    and2_1 \U80_10_/U8  ( .x(\net240[5] ), .a(wd[50]), .b(net267) );
    and2_1 \U80_11_/U8  ( .x(\net240[4] ), .a(wd[51]), .b(net267) );
    and2_1 \U80_12_/U8  ( .x(\net240[3] ), .a(wd[52]), .b(net267) );
    and2_1 \U80_13_/U8  ( .x(\net240[2] ), .a(wd[53]), .b(net267) );
    and2_1 \U80_14_/U8  ( .x(\net240[1] ), .a(wd[54]), .b(net267) );
    and2_1 \U80_15_/U8  ( .x(\net240[0] ), .a(wd[55]), .b(net267) );
    and2_1 \U128_0_/U8  ( .x(\net237[15] ), .a(seq[0]), .b(net269) );
    and2_1 \U128_1_/U8  ( .x(\net237[14] ), .a(pred[0]), .b(net269) );
    and2_1 \U128_2_/U8  ( .x(\net237[13] ), .a(lock[0]), .b(net269) );
    and2_1 \U128_3_/U8  ( .x(\net237[12] ), .a(\hdr[4] ), .b(net269) );
    and2_1 \U128_4_/U8  ( .x(\net237[11] ), .a(\hdr[4] ), .b(net269) );
    and2_1 \U128_5_/U8  ( .x(\net237[10] ), .a(rnw[0]), .b(net269) );
    and2_1 \U128_6_/U8  ( .x(\net237[9] ), .a(size[0]), .b(net269) );
    and2_1 \U128_7_/U8  ( .x(\net237[8] ), .a(size[1]), .b(net269) );
    and2_1 \U128_8_/U8  ( .x(\net237[7] ), .a(seq[1]), .b(net269) );
    and2_1 \U128_9_/U8  ( .x(\net237[6] ), .a(pred[1]), .b(net269) );
    and2_1 \U128_10_/U8  ( .x(\net237[5] ), .a(lock[1]), .b(net269) );
    and2_1 \U128_13_/U8  ( .x(\net237[2] ), .a(rnw[1]), .b(net269) );
    and2_1 \U128_14_/U8  ( .x(\net237[1] ), .a(size[2]), .b(net269) );
    and2_1 \U128_15_/U8  ( .x(\net237[0] ), .a(size[3]), .b(net269) );
    and2_1 \U37_0_/U8  ( .x(\net234[15] ), .a(addr[8]), .b(net259) );
    and2_1 \U37_1_/U8  ( .x(\net234[14] ), .a(addr[9]), .b(net259) );
    and2_1 \U37_2_/U8  ( .x(\net234[13] ), .a(addr[10]), .b(net259) );
    and2_1 \U37_3_/U8  ( .x(\net234[12] ), .a(addr[11]), .b(net259) );
    and2_1 \U37_4_/U8  ( .x(\net234[11] ), .a(addr[12]), .b(net259) );
    and2_1 \U37_5_/U8  ( .x(\net234[10] ), .a(addr[13]), .b(net259) );
    and2_1 \U37_6_/U8  ( .x(\net234[9] ), .a(addr[14]), .b(net259) );
    and2_1 \U37_7_/U8  ( .x(\net234[8] ), .a(addr[15]), .b(net259) );
    and2_1 \U37_8_/U8  ( .x(\net234[7] ), .a(addr[40]), .b(net259) );
    and2_1 \U37_9_/U8  ( .x(\net234[6] ), .a(addr[41]), .b(net259) );
    and2_1 \U37_10_/U8  ( .x(\net234[5] ), .a(addr[42]), .b(net259) );
    and2_1 \U37_11_/U8  ( .x(\net234[4] ), .a(addr[43]), .b(net259) );
    and2_1 \U37_12_/U8  ( .x(\net234[3] ), .a(addr[44]), .b(net259) );
    and2_1 \U37_13_/U8  ( .x(\net234[2] ), .a(addr[45]), .b(net259) );
    and2_1 \U37_14_/U8  ( .x(\net234[1] ), .a(addr[46]), .b(net259) );
    and2_1 \U37_15_/U8  ( .x(\net234[0] ), .a(addr[47]), .b(net259) );
    and2_1 \U33_0_/U8  ( .x(\net231[15] ), .a(addr[16]), .b(net253) );
    and2_1 \U33_1_/U8  ( .x(\net231[14] ), .a(addr[17]), .b(net253) );
    and2_1 \U33_2_/U8  ( .x(\net231[13] ), .a(addr[18]), .b(net253) );
    and2_1 \U33_3_/U8  ( .x(\net231[12] ), .a(addr[19]), .b(net253) );
    and2_1 \U33_4_/U8  ( .x(\net231[11] ), .a(addr[20]), .b(net253) );
    and2_1 \U33_5_/U8  ( .x(\net231[10] ), .a(addr[21]), .b(net253) );
    and2_1 \U33_6_/U8  ( .x(\net231[9] ), .a(addr[22]), .b(net253) );
    and2_1 \U33_7_/U8  ( .x(\net231[8] ), .a(addr[23]), .b(net253) );
    and2_1 \U33_8_/U8  ( .x(\net231[7] ), .a(addr[48]), .b(net253) );
    and2_1 \U33_9_/U8  ( .x(\net231[6] ), .a(addr[49]), .b(net253) );
    and2_1 \U33_10_/U8  ( .x(\net231[5] ), .a(addr[50]), .b(net253) );
    and2_1 \U33_11_/U8  ( .x(\net231[4] ), .a(addr[51]), .b(net253) );
    and2_1 \U33_12_/U8  ( .x(\net231[3] ), .a(addr[52]), .b(net253) );
    and2_1 \U33_13_/U8  ( .x(\net231[2] ), .a(addr[53]), .b(net253) );
    and2_1 \U33_14_/U8  ( .x(\net231[1] ), .a(addr[54]), .b(net253) );
    and2_1 \U33_15_/U8  ( .x(\net231[0] ), .a(addr[55]), .b(net253) );
    and2_1 \U81_0_/U8  ( .x(\net228[15] ), .a(wd[24]), .b(net255) );
    and2_1 \U81_1_/U8  ( .x(\net228[14] ), .a(wd[25]), .b(net255) );
    and2_1 \U81_2_/U8  ( .x(\net228[13] ), .a(wd[26]), .b(net255) );
    and2_1 \U81_3_/U8  ( .x(\net228[12] ), .a(wd[27]), .b(net255) );
    and2_1 \U81_4_/U8  ( .x(\net228[11] ), .a(wd[28]), .b(net255) );
    and2_1 \U81_5_/U8  ( .x(\net228[10] ), .a(wd[29]), .b(net255) );
    and2_1 \U81_6_/U8  ( .x(\net228[9] ), .a(wd[30]), .b(net255) );
    and2_1 \U81_7_/U8  ( .x(\net228[8] ), .a(wd[31]), .b(net255) );
    and2_1 \U81_8_/U8  ( .x(\net228[7] ), .a(wd[56]), .b(net255) );
    and2_1 \U81_9_/U8  ( .x(\net228[6] ), .a(wd[57]), .b(net255) );
    and2_1 \U81_10_/U8  ( .x(\net228[5] ), .a(wd[58]), .b(net255) );
    and2_1 \U81_11_/U8  ( .x(\net228[4] ), .a(wd[59]), .b(net255) );
    and2_1 \U81_12_/U8  ( .x(\net228[3] ), .a(wd[60]), .b(net255) );
    and2_1 \U81_13_/U8  ( .x(\net228[2] ), .a(wd[61]), .b(net255) );
    and2_1 \U81_14_/U8  ( .x(\net228[1] ), .a(wd[62]), .b(net255) );
    and2_1 \U81_15_/U8  ( .x(\net228[0] ), .a(wd[63]), .b(net255) );
    and2_1 \U34_0_/U8  ( .x(\net225[15] ), .a(addr[0]), .b(net251) );
    and2_1 \U34_1_/U8  ( .x(\net225[14] ), .a(addr[1]), .b(net251) );
    and2_1 \U34_2_/U8  ( .x(\net225[13] ), .a(addr[2]), .b(net251) );
    and2_1 \U34_3_/U8  ( .x(\net225[12] ), .a(addr[3]), .b(net251) );
    and2_1 \U34_4_/U8  ( .x(\net225[11] ), .a(addr[4]), .b(net251) );
    and2_1 \U34_5_/U8  ( .x(\net225[10] ), .a(addr[5]), .b(net251) );
    and2_1 \U34_6_/U8  ( .x(\net225[9] ), .a(addr[6]), .b(net251) );
    and2_1 \U34_7_/U8  ( .x(\net225[8] ), .a(addr[7]), .b(net251) );
    and2_1 \U34_8_/U8  ( .x(\net225[7] ), .a(addr[32]), .b(net251) );
    and2_1 \U34_9_/U8  ( .x(\net225[6] ), .a(addr[33]), .b(net251) );
    and2_1 \U34_10_/U8  ( .x(\net225[5] ), .a(addr[34]), .b(net251) );
    and2_1 \U34_11_/U8  ( .x(\net225[4] ), .a(addr[35]), .b(net251) );
    and2_1 \U34_12_/U8  ( .x(\net225[3] ), .a(addr[36]), .b(net251) );
    and2_1 \U34_13_/U8  ( .x(\net225[2] ), .a(addr[37]), .b(net251) );
    and2_1 \U34_14_/U8  ( .x(\net225[1] ), .a(addr[38]), .b(net251) );
    and2_1 \U34_15_/U8  ( .x(\net225[0] ), .a(addr[39]), .b(net251) );
    and2_1 \U30_0_/U8  ( .x(\net222[15] ), .a(addr[24]), .b(net261) );
    and2_1 \U30_1_/U8  ( .x(\net222[14] ), .a(addr[25]), .b(net261) );
    and2_1 \U30_2_/U8  ( .x(\net222[13] ), .a(addr[26]), .b(net261) );
    and2_1 \U30_3_/U8  ( .x(\net222[12] ), .a(addr[27]), .b(net261) );
    and2_1 \U30_4_/U8  ( .x(\net222[11] ), .a(addr[28]), .b(net261) );
    and2_1 \U30_5_/U8  ( .x(\net222[10] ), .a(addr[29]), .b(net261) );
    and2_1 \U30_6_/U8  ( .x(\net222[9] ), .a(addr[30]), .b(net261) );
    and2_1 \U30_7_/U8  ( .x(\net222[8] ), .a(addr[31]), .b(net261) );
    and2_1 \U30_8_/U8  ( .x(\net222[7] ), .a(addr[56]), .b(net261) );
    and2_1 \U30_9_/U8  ( .x(\net222[6] ), .a(addr[57]), .b(net261) );
    and2_1 \U30_10_/U8  ( .x(\net222[5] ), .a(addr[58]), .b(net261) );
    and2_1 \U30_11_/U8  ( .x(\net222[4] ), .a(addr[59]), .b(net261) );
    and2_1 \U30_12_/U8  ( .x(\net222[3] ), .a(addr[60]), .b(net261) );
    and2_1 \U30_13_/U8  ( .x(\net222[2] ), .a(addr[61]), .b(net261) );
    and2_1 \U30_14_/U8  ( .x(\net222[1] ), .a(addr[62]), .b(net261) );
    and2_1 \U30_15_/U8  ( .x(\net222[0] ), .a(addr[63]), .b(net261) );
    and2_1 \U82_0_/U8  ( .x(\net219[15] ), .a(wd[0]), .b(net249) );
    and2_1 \U82_1_/U8  ( .x(\net219[14] ), .a(wd[1]), .b(net249) );
    and2_1 \U82_2_/U8  ( .x(\net219[13] ), .a(wd[2]), .b(net249) );
    and2_1 \U82_3_/U8  ( .x(\net219[12] ), .a(wd[3]), .b(net249) );
    and2_1 \U82_4_/U8  ( .x(\net219[11] ), .a(wd[4]), .b(net249) );
    and2_1 \U82_5_/U8  ( .x(\net219[10] ), .a(wd[5]), .b(net249) );
    and2_1 \U82_6_/U8  ( .x(\net219[9] ), .a(wd[6]), .b(net249) );
    and2_1 \U82_7_/U8  ( .x(\net219[8] ), .a(wd[7]), .b(net249) );
    and2_1 \U82_8_/U8  ( .x(\net219[7] ), .a(wd[32]), .b(net249) );
    and2_1 \U82_9_/U8  ( .x(\net219[6] ), .a(wd[33]), .b(net249) );
    and2_1 \U82_10_/U8  ( .x(\net219[5] ), .a(wd[34]), .b(net249) );
    and2_1 \U82_11_/U8  ( .x(\net219[4] ), .a(wd[35]), .b(net249) );
    and2_1 \U82_12_/U8  ( .x(\net219[3] ), .a(wd[36]), .b(net249) );
    and2_1 \U82_13_/U8  ( .x(\net219[2] ), .a(wd[37]), .b(net249) );
    and2_1 \U82_14_/U8  ( .x(\net219[1] ), .a(wd[38]), .b(net249) );
    and2_1 \U82_15_/U8  ( .x(\net219[0] ), .a(wd[39]), .b(net249) );
    inv_1 \U40_0_/U3  ( .x(\U40_0_/n3 ), .a(\net225[15] ) );
    inv_1 \U40_0_/U4  ( .x(\U40_0_/n4 ), .a(\net234[15] ) );
    inv_1 \U40_0_/U5  ( .x(\net217[15] ), .a(\U40_0_/n5 ) );
    inv_1 \U40_1_/U3  ( .x(\U40_1_/n3 ), .a(\net225[14] ) );
    inv_1 \U40_1_/U4  ( .x(\U40_1_/n4 ), .a(\net234[14] ) );
    inv_1 \U40_1_/U5  ( .x(\net217[14] ), .a(\U40_1_/n5 ) );
    inv_1 \U40_2_/U3  ( .x(\U40_2_/n3 ), .a(\net225[13] ) );
    inv_1 \U40_2_/U4  ( .x(\U40_2_/n4 ), .a(\net234[13] ) );
    inv_1 \U40_2_/U5  ( .x(\net217[13] ), .a(\U40_2_/n5 ) );
    inv_1 \U40_3_/U3  ( .x(\U40_3_/n3 ), .a(\net225[12] ) );
    inv_1 \U40_3_/U4  ( .x(\U40_3_/n4 ), .a(\net234[12] ) );
    inv_1 \U40_3_/U5  ( .x(\net217[12] ), .a(\U40_3_/n5 ) );
    inv_1 \U40_4_/U3  ( .x(\U40_4_/n3 ), .a(\net225[11] ) );
    inv_1 \U40_4_/U4  ( .x(\U40_4_/n4 ), .a(\net234[11] ) );
    inv_1 \U40_4_/U5  ( .x(\net217[11] ), .a(\U40_4_/n5 ) );
    inv_1 \U40_5_/U3  ( .x(\U40_5_/n3 ), .a(\net225[10] ) );
    inv_1 \U40_5_/U4  ( .x(\U40_5_/n4 ), .a(\net234[10] ) );
    inv_1 \U40_5_/U5  ( .x(\net217[10] ), .a(\U40_5_/n5 ) );
    inv_1 \U40_6_/U3  ( .x(\U40_6_/n3 ), .a(\net225[9] ) );
    inv_1 \U40_6_/U4  ( .x(\U40_6_/n4 ), .a(\net234[9] ) );
    inv_1 \U40_6_/U5  ( .x(\net217[9] ), .a(\U40_6_/n5 ) );
    inv_1 \U40_7_/U3  ( .x(\U40_7_/n3 ), .a(\net225[8] ) );
    inv_1 \U40_7_/U4  ( .x(\U40_7_/n4 ), .a(\net234[8] ) );
    inv_1 \U40_7_/U5  ( .x(\net217[8] ), .a(\U40_7_/n5 ) );
    inv_1 \U40_8_/U3  ( .x(\U40_8_/n3 ), .a(\net225[7] ) );
    inv_1 \U40_8_/U4  ( .x(\U40_8_/n4 ), .a(\net234[7] ) );
    inv_1 \U40_8_/U5  ( .x(\net217[7] ), .a(\U40_8_/n5 ) );
    inv_1 \U40_9_/U3  ( .x(\U40_9_/n3 ), .a(\net225[6] ) );
    inv_1 \U40_9_/U4  ( .x(\U40_9_/n4 ), .a(\net234[6] ) );
    inv_1 \U40_9_/U5  ( .x(\net217[6] ), .a(\U40_9_/n5 ) );
    inv_1 \U40_10_/U3  ( .x(\U40_10_/n3 ), .a(\net225[5] ) );
    inv_1 \U40_10_/U4  ( .x(\U40_10_/n4 ), .a(\net234[5] ) );
    inv_1 \U40_10_/U5  ( .x(\net217[5] ), .a(\U40_10_/n5 ) );
    inv_1 \U40_11_/U3  ( .x(\U40_11_/n3 ), .a(\net225[4] ) );
    inv_1 \U40_11_/U4  ( .x(\U40_11_/n4 ), .a(\net234[4] ) );
    inv_1 \U40_11_/U5  ( .x(\net217[4] ), .a(\U40_11_/n5 ) );
    inv_1 \U40_12_/U3  ( .x(\U40_12_/n3 ), .a(\net225[3] ) );
    inv_1 \U40_12_/U4  ( .x(\U40_12_/n4 ), .a(\net234[3] ) );
    inv_1 \U40_12_/U5  ( .x(\net217[3] ), .a(\U40_12_/n5 ) );
    inv_1 \U40_13_/U3  ( .x(\U40_13_/n3 ), .a(\net225[2] ) );
    inv_1 \U40_13_/U4  ( .x(\U40_13_/n4 ), .a(\net234[2] ) );
    inv_1 \U40_13_/U5  ( .x(\net217[2] ), .a(\U40_13_/n5 ) );
    inv_1 \U40_14_/U3  ( .x(\U40_14_/n3 ), .a(\net225[1] ) );
    inv_1 \U40_14_/U4  ( .x(\U40_14_/n4 ), .a(\net234[1] ) );
    inv_1 \U40_14_/U5  ( .x(\net217[1] ), .a(\U40_14_/n5 ) );
    inv_1 \U40_15_/U3  ( .x(\U40_15_/n3 ), .a(\net225[0] ) );
    inv_1 \U40_15_/U4  ( .x(\U40_15_/n4 ), .a(\net234[0] ) );
    inv_1 \U40_15_/U5  ( .x(\net217[0] ), .a(\U40_15_/n5 ) );
    and4_1 \U14_0_/U16  ( .x(\U14_0_/n5 ), .a(\U14_0_/n1 ), .b(\U14_0_/n2 ), 
        .c(\U14_0_/n3 ), .d(\U14_0_/n4 ) );
    inv_1 \U14_0_/U1  ( .x(\U14_0_/n1 ), .a(\net231[15] ) );
    inv_1 \U14_0_/U2  ( .x(\U14_0_/n2 ), .a(\net222[15] ) );
    inv_1 \U14_0_/U3  ( .x(\U14_0_/n3 ), .a(\net237[15] ) );
    inv_1 \U14_0_/U4  ( .x(\U14_0_/n4 ), .a(\net246[15] ) );
    inv_1 \U14_0_/U5  ( .x(\net212[15] ), .a(\U14_0_/n5 ) );
    and4_1 \U14_1_/U16  ( .x(\U14_1_/n5 ), .a(\U14_1_/n1 ), .b(\U14_1_/n2 ), 
        .c(\U14_1_/n3 ), .d(\U14_1_/n4 ) );
    inv_1 \U14_1_/U1  ( .x(\U14_1_/n1 ), .a(\net231[14] ) );
    inv_1 \U14_1_/U2  ( .x(\U14_1_/n2 ), .a(\net222[14] ) );
    inv_1 \U14_1_/U3  ( .x(\U14_1_/n3 ), .a(\net237[14] ) );
    inv_1 \U14_1_/U4  ( .x(\U14_1_/n4 ), .a(\net246[14] ) );
    inv_1 \U14_1_/U5  ( .x(\net212[14] ), .a(\U14_1_/n5 ) );
    and4_1 \U14_2_/U16  ( .x(\U14_2_/n5 ), .a(\U14_2_/n1 ), .b(\U14_2_/n2 ), 
        .c(\U14_2_/n3 ), .d(\U14_2_/n4 ) );
    inv_1 \U14_2_/U1  ( .x(\U14_2_/n1 ), .a(\net231[13] ) );
    inv_1 \U14_2_/U2  ( .x(\U14_2_/n2 ), .a(\net222[13] ) );
    inv_1 \U14_2_/U3  ( .x(\U14_2_/n3 ), .a(\net237[13] ) );
    inv_1 \U14_2_/U4  ( .x(\U14_2_/n4 ), .a(\net246[13] ) );
    inv_1 \U14_2_/U5  ( .x(\net212[13] ), .a(\U14_2_/n5 ) );
    and4_1 \U14_3_/U16  ( .x(\U14_3_/n5 ), .a(\U14_3_/n1 ), .b(\U14_3_/n2 ), 
        .c(\U14_3_/n3 ), .d(\U14_3_/n4 ) );
    inv_1 \U14_3_/U1  ( .x(\U14_3_/n1 ), .a(\net231[12] ) );
    inv_1 \U14_3_/U2  ( .x(\U14_3_/n2 ), .a(\net222[12] ) );
    inv_1 \U14_3_/U3  ( .x(\U14_3_/n3 ), .a(\net237[12] ) );
    inv_1 \U14_3_/U4  ( .x(\U14_3_/n4 ), .a(\net246[12] ) );
    inv_1 \U14_3_/U5  ( .x(\net212[12] ), .a(\U14_3_/n5 ) );
    and4_1 \U14_4_/U16  ( .x(\U14_4_/n5 ), .a(\U14_4_/n1 ), .b(\U14_4_/n2 ), 
        .c(\U14_4_/n3 ), .d(\U14_4_/n4 ) );
    inv_1 \U14_4_/U1  ( .x(\U14_4_/n1 ), .a(\net231[11] ) );
    inv_1 \U14_4_/U2  ( .x(\U14_4_/n2 ), .a(\net222[11] ) );
    inv_1 \U14_4_/U3  ( .x(\U14_4_/n3 ), .a(\net237[11] ) );
    inv_1 \U14_4_/U4  ( .x(\U14_4_/n4 ), .a(\net246[11] ) );
    inv_1 \U14_4_/U5  ( .x(\net212[11] ), .a(\U14_4_/n5 ) );
    and4_1 \U14_5_/U16  ( .x(\U14_5_/n5 ), .a(\U14_5_/n1 ), .b(\U14_5_/n2 ), 
        .c(\U14_5_/n3 ), .d(\U14_5_/n4 ) );
    inv_1 \U14_5_/U1  ( .x(\U14_5_/n1 ), .a(\net231[10] ) );
    inv_1 \U14_5_/U2  ( .x(\U14_5_/n2 ), .a(\net222[10] ) );
    inv_1 \U14_5_/U3  ( .x(\U14_5_/n3 ), .a(\net237[10] ) );
    inv_1 \U14_5_/U4  ( .x(\U14_5_/n4 ), .a(\net246[10] ) );
    inv_1 \U14_5_/U5  ( .x(\net212[10] ), .a(\U14_5_/n5 ) );
    and4_1 \U14_6_/U16  ( .x(\U14_6_/n5 ), .a(\U14_6_/n1 ), .b(\U14_6_/n2 ), 
        .c(\U14_6_/n3 ), .d(\U14_6_/n4 ) );
    inv_1 \U14_6_/U1  ( .x(\U14_6_/n1 ), .a(\net231[9] ) );
    inv_1 \U14_6_/U2  ( .x(\U14_6_/n2 ), .a(\net222[9] ) );
    inv_1 \U14_6_/U3  ( .x(\U14_6_/n3 ), .a(\net237[9] ) );
    inv_1 \U14_6_/U4  ( .x(\U14_6_/n4 ), .a(\net246[9] ) );
    inv_1 \U14_6_/U5  ( .x(\net212[9] ), .a(\U14_6_/n5 ) );
    and4_1 \U14_7_/U16  ( .x(\U14_7_/n5 ), .a(\U14_7_/n1 ), .b(\U14_7_/n2 ), 
        .c(\U14_7_/n3 ), .d(\U14_7_/n4 ) );
    inv_1 \U14_7_/U1  ( .x(\U14_7_/n1 ), .a(\net231[8] ) );
    inv_1 \U14_7_/U2  ( .x(\U14_7_/n2 ), .a(\net222[8] ) );
    inv_1 \U14_7_/U3  ( .x(\U14_7_/n3 ), .a(\net237[8] ) );
    inv_1 \U14_7_/U4  ( .x(\U14_7_/n4 ), .a(\net246[8] ) );
    inv_1 \U14_7_/U5  ( .x(\net212[8] ), .a(\U14_7_/n5 ) );
    and4_1 \U14_8_/U16  ( .x(\U14_8_/n5 ), .a(\U14_8_/n1 ), .b(\U14_8_/n2 ), 
        .c(\U14_8_/n3 ), .d(\U14_8_/n4 ) );
    inv_1 \U14_8_/U1  ( .x(\U14_8_/n1 ), .a(\net231[7] ) );
    inv_1 \U14_8_/U2  ( .x(\U14_8_/n2 ), .a(\net222[7] ) );
    inv_1 \U14_8_/U3  ( .x(\U14_8_/n3 ), .a(\net237[7] ) );
    inv_1 \U14_8_/U4  ( .x(\U14_8_/n4 ), .a(\net246[7] ) );
    inv_1 \U14_8_/U5  ( .x(\net212[7] ), .a(\U14_8_/n5 ) );
    and4_1 \U14_9_/U16  ( .x(\U14_9_/n5 ), .a(\U14_9_/n1 ), .b(\U14_9_/n2 ), 
        .c(\U14_9_/n3 ), .d(\U14_9_/n4 ) );
    inv_1 \U14_9_/U1  ( .x(\U14_9_/n1 ), .a(\net231[6] ) );
    inv_1 \U14_9_/U2  ( .x(\U14_9_/n2 ), .a(\net222[6] ) );
    inv_1 \U14_9_/U3  ( .x(\U14_9_/n3 ), .a(\net237[6] ) );
    inv_1 \U14_9_/U4  ( .x(\U14_9_/n4 ), .a(\net246[6] ) );
    inv_1 \U14_9_/U5  ( .x(\net212[6] ), .a(\U14_9_/n5 ) );
    and4_1 \U14_10_/U16  ( .x(\U14_10_/n5 ), .a(\U14_10_/n1 ), .b(\U14_10_/n2 
        ), .c(\U14_10_/n3 ), .d(\U14_10_/n4 ) );
    inv_1 \U14_10_/U1  ( .x(\U14_10_/n1 ), .a(\net231[5] ) );
    inv_1 \U14_10_/U2  ( .x(\U14_10_/n2 ), .a(\net222[5] ) );
    inv_1 \U14_10_/U3  ( .x(\U14_10_/n3 ), .a(\net237[5] ) );
    inv_1 \U14_10_/U4  ( .x(\U14_10_/n4 ), .a(\net246[5] ) );
    inv_1 \U14_10_/U5  ( .x(\net212[5] ), .a(\U14_10_/n5 ) );
    inv_1 \U14_11_/U1  ( .x(\U14_11_/n1 ), .a(\net231[4] ) );
    inv_1 \U14_11_/U2  ( .x(\U14_11_/n2 ), .a(\net222[4] ) );
    inv_1 \U14_11_/U4  ( .x(\U14_11_/n4 ), .a(\net246[4] ) );
    inv_1 \U14_11_/U5  ( .x(\net212[4] ), .a(\U14_11_/n5 ) );
    inv_1 \U14_12_/U1  ( .x(\U14_12_/n1 ), .a(\net231[3] ) );
    inv_1 \U14_12_/U2  ( .x(\U14_12_/n2 ), .a(\net222[3] ) );
    inv_1 \U14_12_/U4  ( .x(\U14_12_/n4 ), .a(\net246[3] ) );
    inv_1 \U14_12_/U5  ( .x(\net212[3] ), .a(\U14_12_/n5 ) );
    and4_1 \U14_13_/U16  ( .x(\U14_13_/n5 ), .a(\U14_13_/n1 ), .b(\U14_13_/n2 
        ), .c(\U14_13_/n3 ), .d(\U14_13_/n4 ) );
    inv_1 \U14_13_/U1  ( .x(\U14_13_/n1 ), .a(\net231[2] ) );
    inv_1 \U14_13_/U2  ( .x(\U14_13_/n2 ), .a(\net222[2] ) );
    inv_1 \U14_13_/U3  ( .x(\U14_13_/n3 ), .a(\net237[2] ) );
    inv_1 \U14_13_/U4  ( .x(\U14_13_/n4 ), .a(\net246[2] ) );
    inv_1 \U14_13_/U5  ( .x(\net212[2] ), .a(\U14_13_/n5 ) );
    and4_1 \U14_14_/U16  ( .x(\U14_14_/n5 ), .a(\U14_14_/n1 ), .b(\U14_14_/n2 
        ), .c(\U14_14_/n3 ), .d(\U14_14_/n4 ) );
    inv_1 \U14_14_/U1  ( .x(\U14_14_/n1 ), .a(\net231[1] ) );
    inv_1 \U14_14_/U2  ( .x(\U14_14_/n2 ), .a(\net222[1] ) );
    inv_1 \U14_14_/U3  ( .x(\U14_14_/n3 ), .a(\net237[1] ) );
    inv_1 \U14_14_/U4  ( .x(\U14_14_/n4 ), .a(\net246[1] ) );
    inv_1 \U14_14_/U5  ( .x(\net212[1] ), .a(\U14_14_/n5 ) );
    and4_1 \U14_15_/U16  ( .x(\U14_15_/n5 ), .a(\U14_15_/n1 ), .b(\U14_15_/n2 
        ), .c(\U14_15_/n3 ), .d(\U14_15_/n4 ) );
    inv_1 \U14_15_/U1  ( .x(\U14_15_/n1 ), .a(\net231[0] ) );
    inv_1 \U14_15_/U2  ( .x(\U14_15_/n2 ), .a(\net222[0] ) );
    inv_1 \U14_15_/U3  ( .x(\U14_15_/n3 ), .a(\net237[0] ) );
    inv_1 \U14_15_/U4  ( .x(\U14_15_/n4 ), .a(\net246[0] ) );
    inv_1 \U14_15_/U5  ( .x(\net212[0] ), .a(\U14_15_/n5 ) );
    and4_1 \U91_0_/U16  ( .x(\U91_0_/n5 ), .a(\U91_0_/n1 ), .b(\U91_0_/n2 ), 
        .c(\U91_0_/n3 ), .d(\U91_0_/n4 ) );
    inv_1 \U91_0_/U1  ( .x(\U91_0_/n1 ), .a(\net219[15] ) );
    inv_1 \U91_0_/U2  ( .x(\U91_0_/n2 ), .a(\net243[15] ) );
    inv_1 \U91_0_/U3  ( .x(\U91_0_/n3 ), .a(\net240[15] ) );
    inv_1 \U91_0_/U4  ( .x(\U91_0_/n4 ), .a(\net228[15] ) );
    inv_1 \U91_0_/U5  ( .x(\net207[15] ), .a(\U91_0_/n5 ) );
    and4_1 \U91_1_/U16  ( .x(\U91_1_/n5 ), .a(\U91_1_/n1 ), .b(\U91_1_/n2 ), 
        .c(\U91_1_/n3 ), .d(\U91_1_/n4 ) );
    inv_1 \U91_1_/U1  ( .x(\U91_1_/n1 ), .a(\net219[14] ) );
    inv_1 \U91_1_/U2  ( .x(\U91_1_/n2 ), .a(\net243[14] ) );
    inv_1 \U91_1_/U3  ( .x(\U91_1_/n3 ), .a(\net240[14] ) );
    inv_1 \U91_1_/U4  ( .x(\U91_1_/n4 ), .a(\net228[14] ) );
    inv_1 \U91_1_/U5  ( .x(\net207[14] ), .a(\U91_1_/n5 ) );
    and4_1 \U91_2_/U16  ( .x(\U91_2_/n5 ), .a(\U91_2_/n1 ), .b(\U91_2_/n2 ), 
        .c(\U91_2_/n3 ), .d(\U91_2_/n4 ) );
    inv_1 \U91_2_/U1  ( .x(\U91_2_/n1 ), .a(\net219[13] ) );
    inv_1 \U91_2_/U2  ( .x(\U91_2_/n2 ), .a(\net243[13] ) );
    inv_1 \U91_2_/U3  ( .x(\U91_2_/n3 ), .a(\net240[13] ) );
    inv_1 \U91_2_/U4  ( .x(\U91_2_/n4 ), .a(\net228[13] ) );
    inv_1 \U91_2_/U5  ( .x(\net207[13] ), .a(\U91_2_/n5 ) );
    and4_1 \U91_3_/U16  ( .x(\U91_3_/n5 ), .a(\U91_3_/n1 ), .b(\U91_3_/n2 ), 
        .c(\U91_3_/n3 ), .d(\U91_3_/n4 ) );
    inv_1 \U91_3_/U1  ( .x(\U91_3_/n1 ), .a(\net219[12] ) );
    inv_1 \U91_3_/U2  ( .x(\U91_3_/n2 ), .a(\net243[12] ) );
    inv_1 \U91_3_/U3  ( .x(\U91_3_/n3 ), .a(\net240[12] ) );
    inv_1 \U91_3_/U4  ( .x(\U91_3_/n4 ), .a(\net228[12] ) );
    inv_1 \U91_3_/U5  ( .x(\net207[12] ), .a(\U91_3_/n5 ) );
    and4_1 \U91_4_/U16  ( .x(\U91_4_/n5 ), .a(\U91_4_/n1 ), .b(\U91_4_/n2 ), 
        .c(\U91_4_/n3 ), .d(\U91_4_/n4 ) );
    inv_1 \U91_4_/U1  ( .x(\U91_4_/n1 ), .a(\net219[11] ) );
    inv_1 \U91_4_/U2  ( .x(\U91_4_/n2 ), .a(\net243[11] ) );
    inv_1 \U91_4_/U3  ( .x(\U91_4_/n3 ), .a(\net240[11] ) );
    inv_1 \U91_4_/U4  ( .x(\U91_4_/n4 ), .a(\net228[11] ) );
    inv_1 \U91_4_/U5  ( .x(\net207[11] ), .a(\U91_4_/n5 ) );
    and4_1 \U91_5_/U16  ( .x(\U91_5_/n5 ), .a(\U91_5_/n1 ), .b(\U91_5_/n2 ), 
        .c(\U91_5_/n3 ), .d(\U91_5_/n4 ) );
    inv_1 \U91_5_/U1  ( .x(\U91_5_/n1 ), .a(\net219[10] ) );
    inv_1 \U91_5_/U2  ( .x(\U91_5_/n2 ), .a(\net243[10] ) );
    inv_1 \U91_5_/U3  ( .x(\U91_5_/n3 ), .a(\net240[10] ) );
    inv_1 \U91_5_/U4  ( .x(\U91_5_/n4 ), .a(\net228[10] ) );
    inv_1 \U91_5_/U5  ( .x(\net207[10] ), .a(\U91_5_/n5 ) );
    and4_1 \U91_6_/U16  ( .x(\U91_6_/n5 ), .a(\U91_6_/n1 ), .b(\U91_6_/n2 ), 
        .c(\U91_6_/n3 ), .d(\U91_6_/n4 ) );
    inv_1 \U91_6_/U1  ( .x(\U91_6_/n1 ), .a(\net219[9] ) );
    inv_1 \U91_6_/U2  ( .x(\U91_6_/n2 ), .a(\net243[9] ) );
    inv_1 \U91_6_/U3  ( .x(\U91_6_/n3 ), .a(\net240[9] ) );
    inv_1 \U91_6_/U4  ( .x(\U91_6_/n4 ), .a(\net228[9] ) );
    inv_1 \U91_6_/U5  ( .x(\net207[9] ), .a(\U91_6_/n5 ) );
    and4_1 \U91_7_/U16  ( .x(\U91_7_/n5 ), .a(\U91_7_/n1 ), .b(\U91_7_/n2 ), 
        .c(\U91_7_/n3 ), .d(\U91_7_/n4 ) );
    inv_1 \U91_7_/U1  ( .x(\U91_7_/n1 ), .a(\net219[8] ) );
    inv_1 \U91_7_/U2  ( .x(\U91_7_/n2 ), .a(\net243[8] ) );
    inv_1 \U91_7_/U3  ( .x(\U91_7_/n3 ), .a(\net240[8] ) );
    inv_1 \U91_7_/U4  ( .x(\U91_7_/n4 ), .a(\net228[8] ) );
    inv_1 \U91_7_/U5  ( .x(\net207[8] ), .a(\U91_7_/n5 ) );
    and4_1 \U91_8_/U16  ( .x(\U91_8_/n5 ), .a(\U91_8_/n1 ), .b(\U91_8_/n2 ), 
        .c(\U91_8_/n3 ), .d(\U91_8_/n4 ) );
    inv_1 \U91_8_/U1  ( .x(\U91_8_/n1 ), .a(\net219[7] ) );
    inv_1 \U91_8_/U2  ( .x(\U91_8_/n2 ), .a(\net243[7] ) );
    inv_1 \U91_8_/U3  ( .x(\U91_8_/n3 ), .a(\net240[7] ) );
    inv_1 \U91_8_/U4  ( .x(\U91_8_/n4 ), .a(\net228[7] ) );
    inv_1 \U91_8_/U5  ( .x(\net207[7] ), .a(\U91_8_/n5 ) );
    and4_1 \U91_9_/U16  ( .x(\U91_9_/n5 ), .a(\U91_9_/n1 ), .b(\U91_9_/n2 ), 
        .c(\U91_9_/n3 ), .d(\U91_9_/n4 ) );
    inv_1 \U91_9_/U1  ( .x(\U91_9_/n1 ), .a(\net219[6] ) );
    inv_1 \U91_9_/U2  ( .x(\U91_9_/n2 ), .a(\net243[6] ) );
    inv_1 \U91_9_/U3  ( .x(\U91_9_/n3 ), .a(\net240[6] ) );
    inv_1 \U91_9_/U4  ( .x(\U91_9_/n4 ), .a(\net228[6] ) );
    inv_1 \U91_9_/U5  ( .x(\net207[6] ), .a(\U91_9_/n5 ) );
    and4_1 \U91_10_/U16  ( .x(\U91_10_/n5 ), .a(\U91_10_/n1 ), .b(\U91_10_/n2 
        ), .c(\U91_10_/n3 ), .d(\U91_10_/n4 ) );
    inv_1 \U91_10_/U1  ( .x(\U91_10_/n1 ), .a(\net219[5] ) );
    inv_1 \U91_10_/U2  ( .x(\U91_10_/n2 ), .a(\net243[5] ) );
    inv_1 \U91_10_/U3  ( .x(\U91_10_/n3 ), .a(\net240[5] ) );
    inv_1 \U91_10_/U4  ( .x(\U91_10_/n4 ), .a(\net228[5] ) );
    inv_1 \U91_10_/U5  ( .x(\net207[5] ), .a(\U91_10_/n5 ) );
    and4_1 \U91_11_/U16  ( .x(\U91_11_/n5 ), .a(\U91_11_/n1 ), .b(\U91_11_/n2 
        ), .c(\U91_11_/n3 ), .d(\U91_11_/n4 ) );
    inv_1 \U91_11_/U1  ( .x(\U91_11_/n1 ), .a(\net219[4] ) );
    inv_1 \U91_11_/U2  ( .x(\U91_11_/n2 ), .a(\net243[4] ) );
    inv_1 \U91_11_/U3  ( .x(\U91_11_/n3 ), .a(\net240[4] ) );
    inv_1 \U91_11_/U4  ( .x(\U91_11_/n4 ), .a(\net228[4] ) );
    inv_1 \U91_11_/U5  ( .x(\net207[4] ), .a(\U91_11_/n5 ) );
    and4_1 \U91_12_/U16  ( .x(\U91_12_/n5 ), .a(\U91_12_/n1 ), .b(\U91_12_/n2 
        ), .c(\U91_12_/n3 ), .d(\U91_12_/n4 ) );
    inv_1 \U91_12_/U1  ( .x(\U91_12_/n1 ), .a(\net219[3] ) );
    inv_1 \U91_12_/U2  ( .x(\U91_12_/n2 ), .a(\net243[3] ) );
    inv_1 \U91_12_/U3  ( .x(\U91_12_/n3 ), .a(\net240[3] ) );
    inv_1 \U91_12_/U4  ( .x(\U91_12_/n4 ), .a(\net228[3] ) );
    inv_1 \U91_12_/U5  ( .x(\net207[3] ), .a(\U91_12_/n5 ) );
    and4_1 \U91_13_/U16  ( .x(\U91_13_/n5 ), .a(\U91_13_/n1 ), .b(\U91_13_/n2 
        ), .c(\U91_13_/n3 ), .d(\U91_13_/n4 ) );
    inv_1 \U91_13_/U1  ( .x(\U91_13_/n1 ), .a(\net219[2] ) );
    inv_1 \U91_13_/U2  ( .x(\U91_13_/n2 ), .a(\net243[2] ) );
    inv_1 \U91_13_/U3  ( .x(\U91_13_/n3 ), .a(\net240[2] ) );
    inv_1 \U91_13_/U4  ( .x(\U91_13_/n4 ), .a(\net228[2] ) );
    inv_1 \U91_13_/U5  ( .x(\net207[2] ), .a(\U91_13_/n5 ) );
    and4_1 \U91_14_/U16  ( .x(\U91_14_/n5 ), .a(\U91_14_/n1 ), .b(\U91_14_/n2 
        ), .c(\U91_14_/n3 ), .d(\U91_14_/n4 ) );
    inv_1 \U91_14_/U1  ( .x(\U91_14_/n1 ), .a(\net219[1] ) );
    inv_1 \U91_14_/U2  ( .x(\U91_14_/n2 ), .a(\net243[1] ) );
    inv_1 \U91_14_/U3  ( .x(\U91_14_/n3 ), .a(\net240[1] ) );
    inv_1 \U91_14_/U4  ( .x(\U91_14_/n4 ), .a(\net228[1] ) );
    inv_1 \U91_14_/U5  ( .x(\net207[1] ), .a(\U91_14_/n5 ) );
    and4_1 \U91_15_/U16  ( .x(\U91_15_/n5 ), .a(\U91_15_/n1 ), .b(\U91_15_/n2 
        ), .c(\U91_15_/n3 ), .d(\U91_15_/n4 ) );
    inv_1 \U91_15_/U1  ( .x(\U91_15_/n1 ), .a(\net219[0] ) );
    inv_1 \U91_15_/U2  ( .x(\U91_15_/n2 ), .a(\net243[0] ) );
    inv_1 \U91_15_/U3  ( .x(\U91_15_/n3 ), .a(\net240[0] ) );
    inv_1 \U91_15_/U4  ( .x(\U91_15_/n4 ), .a(\net228[0] ) );
    inv_1 \U91_15_/U5  ( .x(\net207[0] ), .a(\U91_15_/n5 ) );
    or3_2 \U93_0_/U12  ( .x(chainl[0]), .a(\net207[15] ), .b(\net217[15] ), 
        .c(\net212[15] ) );
    or3_2 \U93_1_/U12  ( .x(chainl[1]), .a(\net207[14] ), .b(\net217[14] ), 
        .c(\net212[14] ) );
    or3_2 \U93_2_/U12  ( .x(chainl[2]), .a(\net207[13] ), .b(\net217[13] ), 
        .c(\net212[13] ) );
    or3_2 \U93_3_/U12  ( .x(chainl[3]), .a(\net207[12] ), .b(\net217[12] ), 
        .c(\net212[12] ) );
    or3_2 \U93_4_/U12  ( .x(chainl[4]), .a(\net207[11] ), .b(\net217[11] ), 
        .c(\net212[11] ) );
    or3_2 \U93_5_/U12  ( .x(chainl[5]), .a(\net207[10] ), .b(\net217[10] ), 
        .c(\net212[10] ) );
    or3_2 \U93_6_/U12  ( .x(chainl[6]), .a(\net207[9] ), .b(\net217[9] ), .c(
        \net212[9] ) );
    or3_2 \U93_7_/U12  ( .x(chainl[7]), .a(\net207[8] ), .b(\net217[8] ), .c(
        \net212[8] ) );
    or3_2 \U93_8_/U12  ( .x(chainh[0]), .a(\net207[7] ), .b(\net217[7] ), .c(
        \net212[7] ) );
    or3_2 \U93_9_/U12  ( .x(chainh[1]), .a(\net207[6] ), .b(\net217[6] ), .c(
        \net212[6] ) );
    or3_2 \U93_10_/U12  ( .x(chainh[2]), .a(\net207[5] ), .b(\net217[5] ), .c(
        \net212[5] ) );
    or3_2 \U93_11_/U12  ( .x(chainh[3]), .a(\net207[4] ), .b(\net217[4] ), .c(
        \net212[4] ) );
    or3_2 \U93_12_/U12  ( .x(chainh[4]), .a(\net207[3] ), .b(\net217[3] ), .c(
        \net212[3] ) );
    or3_2 \U93_13_/U12  ( .x(chainh[5]), .a(\net207[2] ), .b(\net217[2] ), .c(
        \net212[2] ) );
    or3_2 \U93_14_/U12  ( .x(chainh[6]), .a(\net207[1] ), .b(\net217[1] ), .c(
        \net212[1] ) );
    or3_2 \U93_15_/U12  ( .x(chainh[7]), .a(\net207[0] ), .b(\net217[0] ), .c(
        \net212[0] ) );
    inv_1 \U152/U3  ( .x(net198), .a(sendreq) );
    ao23_1 \U158/U19/U21/U1/U1  ( .x(net131), .a(net132), .b(net131), .c(
        net132), .d(rnw[1]), .e(rnw[1]) );
    ao23_1 \U157/U19/U21/U1/U1  ( .x(net176), .a(net132), .b(net176), .c(
        net132), .d(rnw[0]), .e(rnw[0]) );
    ao222_1 \U123/U18/U1/U1  ( .x(net136), .a(net185), .b(net187), .c(net185), 
        .d(net136), .e(net187), .f(net136) );
    aoi21_1 \U151/U30/U1/U1  ( .x(\hdr[4] ), .a(\U151/Z ), .b(net138), .c(
        net198) );
    inv_1 \U151/U30/U1/U2  ( .x(\U151/Z ), .a(\hdr[4] ) );
    nor3_1 \U148/U21/Unr  ( .x(\U148/U21/nr ), .a(net191), .b(net136), .c(
        net293) );
    nand3_1 \U148/U21/Und  ( .x(\U148/U21/nd ), .a(net191), .b(net136), .c(
        net293) );
    oa21_1 \U148/U21/U1  ( .x(\U148/U21/n2 ), .a(\U148/U21/n2 ), .b(
        \U148/U21/nr ), .c(\U148/U21/nd ) );
    inv_1 \U148/U21/U3  ( .x(ack), .a(\U148/U21/n2 ) );
    buf_3 U1 ( .x(n1), .a(net138) );
    buf_3 U2 ( .x(net138), .a(nia) );
    buf_3 U3 ( .x(net269), .a(net146) );
    buf_3 U4 ( .x(net255), .a(\bs[5] ) );
    buf_3 U5 ( .x(net267), .a(\bs[6] ) );
    buf_3 U6 ( .x(net253), .a(\bs[2] ) );
    buf_3 U7 ( .x(net249), .a(\bs[8] ) );
    buf_3 U8 ( .x(net263), .a(\bs[7] ) );
    buf_3 U9 ( .x(net259), .a(\bs[3] ) );
    buf_3 U10 ( .x(net251), .a(\bs[4] ) );
    buf_3 U11 ( .x(net261), .a(\bs[1] ) );
    buf_3 U12 ( .x(net265), .a(\bs[0] ) );
    and2_1 U13 ( .x(\U40_2_/n5 ), .a(\U40_2_/n3 ), .b(\U40_2_/n4 ) );
    and2_1 U14 ( .x(\U40_1_/n5 ), .a(\U40_1_/n3 ), .b(\U40_1_/n4 ) );
    and2_1 U15 ( .x(\U40_9_/n5 ), .a(\U40_9_/n3 ), .b(\U40_9_/n4 ) );
    and2_1 U16 ( .x(\U40_8_/n5 ), .a(\U40_8_/n3 ), .b(\U40_8_/n4 ) );
    and2_1 U17 ( .x(\U40_13_/n5 ), .a(\U40_13_/n3 ), .b(\U40_13_/n4 ) );
    and2_1 U18 ( .x(\U40_0_/n5 ), .a(\U40_0_/n3 ), .b(\U40_0_/n4 ) );
    and2_1 U19 ( .x(\U40_5_/n5 ), .a(\U40_5_/n3 ), .b(\U40_5_/n4 ) );
    and2_1 U20 ( .x(\U40_4_/n5 ), .a(\U40_4_/n3 ), .b(\U40_4_/n4 ) );
    and3_1 U21 ( .x(\U14_12_/n5 ), .a(\U14_12_/n2 ), .b(\U14_12_/n4 ), .c(
        \U14_12_/n1 ) );
    and2_1 U22 ( .x(\U40_12_/n5 ), .a(\U40_12_/n3 ), .b(\U40_12_/n4 ) );
    and2_1 U23 ( .x(\U40_3_/n5 ), .a(\U40_3_/n3 ), .b(\U40_3_/n4 ) );
    and3_1 U24 ( .x(\U14_11_/n5 ), .a(\U14_11_/n2 ), .b(\U14_11_/n4 ), .c(
        \U14_11_/n1 ) );
    and2_1 U25 ( .x(\U40_11_/n5 ), .a(\U40_11_/n3 ), .b(\U40_11_/n4 ) );
    and2_1 U26 ( .x(\U40_10_/n5 ), .a(\U40_10_/n3 ), .b(\U40_10_/n4 ) );
    and2_1 U27 ( .x(\U40_15_/n5 ), .a(\U40_15_/n3 ), .b(\U40_15_/n4 ) );
    and2_1 U28 ( .x(\U40_7_/n5 ), .a(\U40_7_/n3 ), .b(\U40_7_/n4 ) );
    and2_1 U29 ( .x(\U40_6_/n5 ), .a(\U40_6_/n3 ), .b(\U40_6_/n4 ) );
    and2_1 U30 ( .x(\U40_14_/n5 ), .a(\U40_14_/n3 ), .b(\U40_14_/n4 ) );
endmodule


module chain_dr2fr_byte_2 ( eop_ack, ia, o, eop, ih, il, nReset, noa );
output [4:0] o;
input  [7:0] ih;
input  [7:0] il;
input  eop, nReset, noa;
output eop_ack, ia;
    wire eop_ack_wire, nbReset, eop_pass, nxa, naa, nlowack, \twobitack[0] , 
        \twobitack[1] , nhighack, \twobitack[2] , \twobitack[3] , \U1018/Z , 
        \U1270/net189 , \U1270/net192 , \U1270/net191 , net199, \U1270/net190 , 
        \U1270/U1141/Z , \U1268/net189 , \U1268/net192 , \U1268/net191 , 
        net194, \U1268/net190 , \U1268/U1141/Z , \U1224/nack[0] , \x[3] , 
        \x[2] , \U1224/nack[1] , \x[1] , \U1224/net4 , \x[0] , 
        \U1224/U1125/U28/U1/clr , asel, \U1224/U1125/U28/U1/set , 
        \U1224/U1122/U28/U1/clr , csel, nca, \U1224/U1122/U28/U1/set , 
        \U1224/U916_0_/U25/U1/clr , \a[0] , \c[0] , \U1224/U916_0_/U25/U1/ob , 
        \U1224/U916_1_/U25/U1/clr , \a[1] , \c[1] , \U1224/U916_1_/U25/U1/ob , 
        \U1224/U916_2_/U25/U1/clr , \a[2] , \c[2] , \U1224/U916_2_/U25/U1/ob , 
        \U1224/U916_3_/U25/U1/clr , \a[3] , \c[3] , \U1224/U916_3_/U25/U1/ob , 
        \U1209/nack[0] , \U1209/nack[1] , \U1209/net4 , 
        \U1209/U1125/U28/U1/clr , xsel, \U1209/U1125/U28/U1/set , 
        \U1209/U1122/U28/U1/clr , ysel, nyla, \U1209/U1122/U28/U1/set , 
        \U1209/U916_0_/U25/U1/clr , \yl[0] , \U1209/U916_0_/U25/U1/ob , 
        \U1209/U916_1_/U25/U1/clr , \yl[1] , \U1209/U916_1_/U25/U1/ob , 
        \U1209/U916_2_/U25/U1/clr , \yl[2] , \U1209/U916_2_/U25/U1/ob , 
        \U1209/U916_3_/U25/U1/clr , \yl[3] , \U1209/U916_3_/U25/U1/ob , 
        \U1213/nack[0] , \y[3] , \y[2] , \U1213/nack[1] , \y[1] , \U1213/net4 , 
        \y[0] , \U1213/U1125/U28/U1/clr , bsel, nba, \U1213/U1125/U28/U1/set , 
        \U1213/U1122/U28/U1/clr , dsel, nda, \U1213/U1122/U28/U1/set , 
        \U1213/U916_0_/U25/U1/clr , nya, \b[0] , \d[0] , 
        \U1213/U916_0_/U25/U1/ob , \U1213/U916_1_/U25/U1/clr , \b[1] , \d[1] , 
        \U1213/U916_1_/U25/U1/ob , \U1213/U916_2_/U25/U1/clr , \b[2] , \d[2] , 
        \U1213/U916_2_/U25/U1/ob , \U1213/U916_3_/U25/U1/clr , \b[3] , \d[3] , 
        \U1213/U916_3_/U25/U1/ob , \cdh[0] , \cdh[1] , \cdl[0] , \cdl[1] , 
        \cdh[2] , \cdh[3] , \cdl[2] , \cdl[3] , cg, \U1296/ng , net195, 
        \U1296/U1384/Z , \U1296/U1386/U25/U1/clr , \U1296/U1386/U25/U1/ob , dg, 
        \U1298/ng , net193, \U1298/U1384/Z , \U1298/U1386/U25/U1/clr , 
        \U1298/U1386/U25/U1/ob , bg, \U1306/ng , \U1306/U1384/Z , 
        \U1306/U1386/U25/U1/clr , \U1306/U1386/U25/U1/ob , ag, \U1295/ng , 
        \U1295/U1384/Z , \U1295/U1386/U25/U1/clr , \U1295/U1386/U25/U1/ob , 
        \U1297/s , \U1297/r , \U1297/nback , \U1297/naack , \U1297/reset , 
        \U1297/U1128/U28/U1/clr , \U1297/U1128/U28/U1/set , 
        \U1297/U1127/U28/U1/clr , \U1297/U1127/U28/U1/set , \U1300/s , 
        \U1300/r , \U1300/nback , \U1300/naack , \U1300/reset , 
        \U1300/U1128/U28/U1/clr , \U1300/U1128/U28/U1/set , 
        \U1300/U1127/U28/U1/clr , \U1300/U1127/U28/U1/set , 
        \U1289/U1150/U28/U1/clr , \U1289/bnreset , \U1289/U1150/U28/U1/set , 
        \U1289/U1152/U28/U1/clr , \U1289/U1152/U28/U1/set , 
        \U1289/U1149/U28/U1/clr , \U1289/U1149/U28/U1/set , 
        \U1289/U1151/U28/U1/clr , \U1289/U1151/U28/U1/set , 
        \U1289/U1148/net189 , \U1289/U1148/net192 , \U1289/U1148/net191 , 
        \U1289/U1148/net190 , \U1289/U1148/U1141/Z , \U1271/U1150/U28/U1/clr , 
        \U1271/bnreset , \U1271/U1150/U28/U1/set , \U1271/U1152/U28/U1/clr , 
        \U1271/U1152/U28/U1/set , \U1271/U1149/U28/U1/clr , 
        \U1271/U1149/U28/U1/set , \U1271/U1151/U28/U1/clr , 
        \U1271/U1151/U28/U1/set , \U1271/U1148/net189 , \U1271/U1148/net192 , 
        \U1271/U1148/net191 , \U1271/U1148/net190 , \U1271/U1148/U1141/Z , 
        \U1225/s , \U1225/r , \U1225/nback , \U1225/naack , \U1225/reset , 
        \U1308/nack[1] , \U1308/nack[0] ;
    assign eop_ack = eop_ack_wire;
    assign o[4] = eop_ack_wire;
    buf_2 U1231 ( .x(nbReset), .a(nReset) );
    and3_1 \U1194/U9  ( .x(eop_pass), .a(nxa), .b(naa), .c(eop) );
    ao222_1 \U1301/U18/U1/U1  ( .x(nlowack), .a(\twobitack[0] ), .b(
        \twobitack[1] ), .c(\twobitack[0] ), .d(nlowack), .e(\twobitack[1] ), 
        .f(nlowack) );
    ao222_1 \U1302/U18/U1/U1  ( .x(nhighack), .a(\twobitack[2] ), .b(
        \twobitack[3] ), .c(\twobitack[2] ), .d(nhighack), .e(\twobitack[3] ), 
        .f(nhighack) );
    aoi222_1 \U1018/U30/U1  ( .x(ia), .a(nhighack), .b(nlowack), .c(nhighack), 
        .d(\U1018/Z ), .e(nlowack), .f(\U1018/Z ) );
    inv_1 \U1018/U30/Uinv  ( .x(\U1018/Z ), .a(ia) );
    ao222_2 \U1038/U19/U1/U1  ( .x(eop_ack_wire), .a(eop_pass), .b(noa), .c(
        eop_pass), .d(eop_ack_wire), .e(noa), .f(eop_ack_wire) );
    inv_1 \U1270/U1147/U3  ( .x(\U1270/net189 ), .a(nbReset) );
    nor2_1 \U1270/U582/U5  ( .x(\U1270/net192 ), .a(il[4]), .b(ih[4]) );
    nor2_1 \U1270/U580/U5  ( .x(\U1270/net191 ), .a(il[5]), .b(ih[5]) );
    nor2_2 \U1270/U1146/U6  ( .x(net199), .a(\U1270/net190 ), .b(
        \U1270/net189 ) );
    aoi222_1 \U1270/U1141/U30/U1  ( .x(\U1270/net190 ), .a(\U1270/net191 ), 
        .b(\U1270/net192 ), .c(\U1270/net191 ), .d(\U1270/U1141/Z ), .e(
        \U1270/net192 ), .f(\U1270/U1141/Z ) );
    inv_1 \U1270/U1141/U30/Uinv  ( .x(\U1270/U1141/Z ), .a(\U1270/net190 ) );
    inv_1 \U1268/U1147/U3  ( .x(\U1268/net189 ), .a(nbReset) );
    nor2_1 \U1268/U582/U5  ( .x(\U1268/net192 ), .a(il[6]), .b(ih[6]) );
    nor2_1 \U1268/U580/U5  ( .x(\U1268/net191 ), .a(il[7]), .b(ih[7]) );
    nor2_2 \U1268/U1146/U6  ( .x(net194), .a(\U1268/net190 ), .b(
        \U1268/net189 ) );
    aoi222_1 \U1268/U1141/U30/U1  ( .x(\U1268/net190 ), .a(\U1268/net191 ), 
        .b(\U1268/net192 ), .c(\U1268/net191 ), .d(\U1268/U1141/Z ), .e(
        \U1268/net192 ), .f(\U1268/U1141/Z ) );
    inv_1 \U1268/U1141/U30/Uinv  ( .x(\U1268/U1141/Z ), .a(\U1268/net190 ) );
    nor2_1 \U1224/U1128/U5  ( .x(\U1224/nack[0] ), .a(\x[3] ), .b(\x[2] ) );
    nor3_1 \U1224/U1127/U7  ( .x(\U1224/nack[1] ), .a(\x[1] ), .b(\U1224/net4 
        ), .c(\x[0] ) );
    inv_1 \U1224/U907/U3  ( .x(\U1224/net4 ), .a(nbReset) );
    aoai211_1 \U1224/U1125/U28/U1/U1  ( .x(\U1224/U1125/U28/U1/clr ), .a(
        \U1224/nack[1] ), .b(\U1224/nack[0] ), .c(asel), .d(naa) );
    nand3_1 \U1224/U1125/U28/U1/U2  ( .x(\U1224/U1125/U28/U1/set ), .a(asel), 
        .b(\U1224/nack[1] ), .c(\U1224/nack[0] ) );
    nand2_2 \U1224/U1125/U28/U1/U3  ( .x(naa), .a(\U1224/U1125/U28/U1/clr ), 
        .b(\U1224/U1125/U28/U1/set ) );
    aoai211_1 \U1224/U1122/U28/U1/U1  ( .x(\U1224/U1122/U28/U1/clr ), .a(
        \U1224/nack[0] ), .b(\U1224/nack[1] ), .c(csel), .d(nca) );
    nand3_1 \U1224/U1122/U28/U1/U2  ( .x(\U1224/U1122/U28/U1/set ), .a(csel), 
        .b(\U1224/nack[0] ), .c(\U1224/nack[1] ) );
    nand2_2 \U1224/U1122/U28/U1/U3  ( .x(nca), .a(\U1224/U1122/U28/U1/clr ), 
        .b(\U1224/U1122/U28/U1/set ) );
    oa31_1 \U1224/U916_0_/U25/U1/Uclr  ( .x(\U1224/U916_0_/U25/U1/clr ), .a(
        nxa), .b(\a[0] ), .c(\c[0] ), .d(\x[0] ) );
    oaoi211_1 \U1224/U916_0_/U25/U1/Uaoi  ( .x(\U1224/U916_0_/U25/U1/ob ), .a(
        \a[0] ), .b(\c[0] ), .c(nxa), .d(\U1224/U916_0_/U25/U1/clr ) );
    inv_2 \U1224/U916_0_/U25/U1/Ui  ( .x(\x[0] ), .a(\U1224/U916_0_/U25/U1/ob 
        ) );
    oa31_1 \U1224/U916_1_/U25/U1/Uclr  ( .x(\U1224/U916_1_/U25/U1/clr ), .a(
        nxa), .b(\a[1] ), .c(\c[1] ), .d(\x[1] ) );
    oaoi211_1 \U1224/U916_1_/U25/U1/Uaoi  ( .x(\U1224/U916_1_/U25/U1/ob ), .a(
        \a[1] ), .b(\c[1] ), .c(nxa), .d(\U1224/U916_1_/U25/U1/clr ) );
    inv_2 \U1224/U916_1_/U25/U1/Ui  ( .x(\x[1] ), .a(\U1224/U916_1_/U25/U1/ob 
        ) );
    oa31_1 \U1224/U916_2_/U25/U1/Uclr  ( .x(\U1224/U916_2_/U25/U1/clr ), .a(
        nxa), .b(\a[2] ), .c(\c[2] ), .d(\x[2] ) );
    oaoi211_1 \U1224/U916_2_/U25/U1/Uaoi  ( .x(\U1224/U916_2_/U25/U1/ob ), .a(
        \a[2] ), .b(\c[2] ), .c(nxa), .d(\U1224/U916_2_/U25/U1/clr ) );
    inv_2 \U1224/U916_2_/U25/U1/Ui  ( .x(\x[2] ), .a(\U1224/U916_2_/U25/U1/ob 
        ) );
    oa31_1 \U1224/U916_3_/U25/U1/Uclr  ( .x(\U1224/U916_3_/U25/U1/clr ), .a(
        nxa), .b(\a[3] ), .c(\c[3] ), .d(\x[3] ) );
    oaoi211_1 \U1224/U916_3_/U25/U1/Uaoi  ( .x(\U1224/U916_3_/U25/U1/ob ), .a(
        \a[3] ), .b(\c[3] ), .c(nxa), .d(\U1224/U916_3_/U25/U1/clr ) );
    inv_2 \U1224/U916_3_/U25/U1/Ui  ( .x(\x[3] ), .a(\U1224/U916_3_/U25/U1/ob 
        ) );
    nor2_1 \U1209/U1128/U5  ( .x(\U1209/nack[0] ), .a(o[3]), .b(o[2]) );
    nor3_1 \U1209/U1127/U7  ( .x(\U1209/nack[1] ), .a(o[1]), .b(\U1209/net4 ), 
        .c(o[0]) );
    inv_1 \U1209/U907/U3  ( .x(\U1209/net4 ), .a(nbReset) );
    aoai211_1 \U1209/U1125/U28/U1/U1  ( .x(\U1209/U1125/U28/U1/clr ), .a(
        \U1209/nack[1] ), .b(\U1209/nack[0] ), .c(xsel), .d(nxa) );
    nand3_1 \U1209/U1125/U28/U1/U2  ( .x(\U1209/U1125/U28/U1/set ), .a(xsel), 
        .b(\U1209/nack[1] ), .c(\U1209/nack[0] ) );
    nand2_2 \U1209/U1125/U28/U1/U3  ( .x(nxa), .a(\U1209/U1125/U28/U1/clr ), 
        .b(\U1209/U1125/U28/U1/set ) );
    aoai211_1 \U1209/U1122/U28/U1/U1  ( .x(\U1209/U1122/U28/U1/clr ), .a(
        \U1209/nack[0] ), .b(\U1209/nack[1] ), .c(ysel), .d(nyla) );
    nand3_1 \U1209/U1122/U28/U1/U2  ( .x(\U1209/U1122/U28/U1/set ), .a(ysel), 
        .b(\U1209/nack[0] ), .c(\U1209/nack[1] ) );
    nand2_2 \U1209/U1122/U28/U1/U3  ( .x(nyla), .a(\U1209/U1122/U28/U1/clr ), 
        .b(\U1209/U1122/U28/U1/set ) );
    oa31_1 \U1209/U916_0_/U25/U1/Uclr  ( .x(\U1209/U916_0_/U25/U1/clr ), .a(
        noa), .b(\x[0] ), .c(\yl[0] ), .d(o[0]) );
    oaoi211_1 \U1209/U916_0_/U25/U1/Uaoi  ( .x(\U1209/U916_0_/U25/U1/ob ), .a(
        \x[0] ), .b(\yl[0] ), .c(noa), .d(\U1209/U916_0_/U25/U1/clr ) );
    inv_2 \U1209/U916_0_/U25/U1/Ui  ( .x(o[0]), .a(\U1209/U916_0_/U25/U1/ob )
         );
    oa31_1 \U1209/U916_1_/U25/U1/Uclr  ( .x(\U1209/U916_1_/U25/U1/clr ), .a(
        noa), .b(\x[1] ), .c(\yl[1] ), .d(o[1]) );
    oaoi211_1 \U1209/U916_1_/U25/U1/Uaoi  ( .x(\U1209/U916_1_/U25/U1/ob ), .a(
        \x[1] ), .b(\yl[1] ), .c(noa), .d(\U1209/U916_1_/U25/U1/clr ) );
    inv_2 \U1209/U916_1_/U25/U1/Ui  ( .x(o[1]), .a(\U1209/U916_1_/U25/U1/ob )
         );
    oa31_1 \U1209/U916_2_/U25/U1/Uclr  ( .x(\U1209/U916_2_/U25/U1/clr ), .a(
        noa), .b(\x[2] ), .c(\yl[2] ), .d(o[2]) );
    oaoi211_1 \U1209/U916_2_/U25/U1/Uaoi  ( .x(\U1209/U916_2_/U25/U1/ob ), .a(
        \x[2] ), .b(\yl[2] ), .c(noa), .d(\U1209/U916_2_/U25/U1/clr ) );
    inv_2 \U1209/U916_2_/U25/U1/Ui  ( .x(o[2]), .a(\U1209/U916_2_/U25/U1/ob )
         );
    oa31_1 \U1209/U916_3_/U25/U1/Uclr  ( .x(\U1209/U916_3_/U25/U1/clr ), .a(
        noa), .b(\x[3] ), .c(\yl[3] ), .d(o[3]) );
    oaoi211_1 \U1209/U916_3_/U25/U1/Uaoi  ( .x(\U1209/U916_3_/U25/U1/ob ), .a(
        \x[3] ), .b(\yl[3] ), .c(noa), .d(\U1209/U916_3_/U25/U1/clr ) );
    inv_2 \U1209/U916_3_/U25/U1/Ui  ( .x(o[3]), .a(\U1209/U916_3_/U25/U1/ob )
         );
    nor2_1 \U1213/U1128/U5  ( .x(\U1213/nack[0] ), .a(\y[3] ), .b(\y[2] ) );
    nor3_1 \U1213/U1127/U7  ( .x(\U1213/nack[1] ), .a(\y[1] ), .b(\U1213/net4 
        ), .c(\y[0] ) );
    inv_1 \U1213/U907/U3  ( .x(\U1213/net4 ), .a(nbReset) );
    aoai211_1 \U1213/U1125/U28/U1/U1  ( .x(\U1213/U1125/U28/U1/clr ), .a(
        \U1213/nack[1] ), .b(\U1213/nack[0] ), .c(bsel), .d(nba) );
    nand3_1 \U1213/U1125/U28/U1/U2  ( .x(\U1213/U1125/U28/U1/set ), .a(bsel), 
        .b(\U1213/nack[1] ), .c(\U1213/nack[0] ) );
    nand2_2 \U1213/U1125/U28/U1/U3  ( .x(nba), .a(\U1213/U1125/U28/U1/clr ), 
        .b(\U1213/U1125/U28/U1/set ) );
    aoai211_1 \U1213/U1122/U28/U1/U1  ( .x(\U1213/U1122/U28/U1/clr ), .a(
        \U1213/nack[0] ), .b(\U1213/nack[1] ), .c(dsel), .d(nda) );
    nand3_1 \U1213/U1122/U28/U1/U2  ( .x(\U1213/U1122/U28/U1/set ), .a(dsel), 
        .b(\U1213/nack[0] ), .c(\U1213/nack[1] ) );
    nand2_2 \U1213/U1122/U28/U1/U3  ( .x(nda), .a(\U1213/U1122/U28/U1/clr ), 
        .b(\U1213/U1122/U28/U1/set ) );
    oa31_1 \U1213/U916_0_/U25/U1/Uclr  ( .x(\U1213/U916_0_/U25/U1/clr ), .a(
        nya), .b(\b[0] ), .c(\d[0] ), .d(\y[0] ) );
    oaoi211_1 \U1213/U916_0_/U25/U1/Uaoi  ( .x(\U1213/U916_0_/U25/U1/ob ), .a(
        \b[0] ), .b(\d[0] ), .c(nya), .d(\U1213/U916_0_/U25/U1/clr ) );
    inv_2 \U1213/U916_0_/U25/U1/Ui  ( .x(\y[0] ), .a(\U1213/U916_0_/U25/U1/ob 
        ) );
    oa31_1 \U1213/U916_1_/U25/U1/Uclr  ( .x(\U1213/U916_1_/U25/U1/clr ), .a(
        nya), .b(\b[1] ), .c(\d[1] ), .d(\y[1] ) );
    oaoi211_1 \U1213/U916_1_/U25/U1/Uaoi  ( .x(\U1213/U916_1_/U25/U1/ob ), .a(
        \b[1] ), .b(\d[1] ), .c(nya), .d(\U1213/U916_1_/U25/U1/clr ) );
    inv_2 \U1213/U916_1_/U25/U1/Ui  ( .x(\y[1] ), .a(\U1213/U916_1_/U25/U1/ob 
        ) );
    oa31_1 \U1213/U916_2_/U25/U1/Uclr  ( .x(\U1213/U916_2_/U25/U1/clr ), .a(
        nya), .b(\b[2] ), .c(\d[2] ), .d(\y[2] ) );
    oaoi211_1 \U1213/U916_2_/U25/U1/Uaoi  ( .x(\U1213/U916_2_/U25/U1/ob ), .a(
        \b[2] ), .b(\d[2] ), .c(nya), .d(\U1213/U916_2_/U25/U1/clr ) );
    inv_2 \U1213/U916_2_/U25/U1/Ui  ( .x(\y[2] ), .a(\U1213/U916_2_/U25/U1/ob 
        ) );
    oa31_1 \U1213/U916_3_/U25/U1/Uclr  ( .x(\U1213/U916_3_/U25/U1/clr ), .a(
        nya), .b(\b[3] ), .c(\d[3] ), .d(\y[3] ) );
    oaoi211_1 \U1213/U916_3_/U25/U1/Uaoi  ( .x(\U1213/U916_3_/U25/U1/ob ), .a(
        \b[3] ), .b(\d[3] ), .c(nya), .d(\U1213/U916_3_/U25/U1/clr ) );
    inv_2 \U1213/U916_3_/U25/U1/Ui  ( .x(\y[3] ), .a(\U1213/U916_3_/U25/U1/ob 
        ) );
    and3_2 \U1210/U1138/U9  ( .x(\d[3] ), .a(\cdh[0] ), .b(nda), .c(\cdh[1] )
         );
    and3_2 \U1210/U1137/U9  ( .x(\d[2] ), .a(\cdl[0] ), .b(nda), .c(\cdh[1] )
         );
    and3_2 \U1210/U1139/U9  ( .x(\d[1] ), .a(\cdh[0] ), .b(nda), .c(\cdl[1] )
         );
    and3_2 \U1210/U1136/U9  ( .x(\d[0] ), .a(\cdl[0] ), .b(nda), .c(\cdl[1] )
         );
    and3_2 \U1162/U1138/U9  ( .x(\a[3] ), .a(ih[6]), .b(naa), .c(ih[7]) );
    and3_2 \U1162/U1137/U9  ( .x(\a[2] ), .a(il[6]), .b(naa), .c(ih[7]) );
    and3_2 \U1162/U1139/U9  ( .x(\a[1] ), .a(ih[6]), .b(naa), .c(il[7]) );
    and3_2 \U1162/U1136/U9  ( .x(\a[0] ), .a(il[6]), .b(naa), .c(il[7]) );
    and3_2 \U1211/U1138/U9  ( .x(\b[3] ), .a(ih[4]), .b(nba), .c(ih[5]) );
    and3_2 \U1211/U1137/U9  ( .x(\b[2] ), .a(il[4]), .b(nba), .c(ih[5]) );
    and3_2 \U1211/U1139/U9  ( .x(\b[1] ), .a(ih[4]), .b(nba), .c(il[5]) );
    and3_2 \U1211/U1136/U9  ( .x(\b[0] ), .a(il[4]), .b(nba), .c(il[5]) );
    and3_2 \U1163/U1138/U9  ( .x(\c[3] ), .a(\cdh[2] ), .b(nca), .c(\cdh[3] )
         );
    and3_2 \U1163/U1137/U9  ( .x(\c[2] ), .a(\cdl[2] ), .b(nca), .c(\cdh[3] )
         );
    and3_2 \U1163/U1139/U9  ( .x(\c[1] ), .a(\cdh[2] ), .b(nca), .c(\cdl[3] )
         );
    and3_2 \U1163/U1136/U9  ( .x(\c[0] ), .a(\cdl[2] ), .b(nca), .c(\cdl[3] )
         );
    and2_1 \U1296/U1385/U8  ( .x(cg), .a(nbReset), .b(\U1296/ng ) );
    aoi222_1 \U1296/U1384/U30/U1  ( .x(\U1296/ng ), .a(nca), .b(net195), .c(
        nca), .d(\U1296/U1384/Z ), .e(net195), .f(\U1296/U1384/Z ) );
    inv_1 \U1296/U1384/U30/Uinv  ( .x(\U1296/U1384/Z ), .a(\U1296/ng ) );
    oa31_1 \U1296/U1386/U25/U1/Uclr  ( .x(\U1296/U1386/U25/U1/clr ), .a(
        \twobitack[2] ), .b(cg), .c(nca), .d(net195) );
    oaoi211_1 \U1296/U1386/U25/U1/Uaoi  ( .x(\U1296/U1386/U25/U1/ob ), .a(cg), 
        .b(nca), .c(\twobitack[2] ), .d(\U1296/U1386/U25/U1/clr ) );
    inv_2 \U1296/U1386/U25/U1/Ui  ( .x(net195), .a(\U1296/U1386/U25/U1/ob ) );
    and2_1 \U1298/U1385/U8  ( .x(dg), .a(nbReset), .b(\U1298/ng ) );
    aoi222_1 \U1298/U1384/U30/U1  ( .x(\U1298/ng ), .a(nda), .b(net193), .c(
        nda), .d(\U1298/U1384/Z ), .e(net193), .f(\U1298/U1384/Z ) );
    inv_1 \U1298/U1384/U30/Uinv  ( .x(\U1298/U1384/Z ), .a(\U1298/ng ) );
    oa31_1 \U1298/U1386/U25/U1/Uclr  ( .x(\U1298/U1386/U25/U1/clr ), .a(
        \twobitack[0] ), .b(dg), .c(nda), .d(net193) );
    oaoi211_1 \U1298/U1386/U25/U1/Uaoi  ( .x(\U1298/U1386/U25/U1/ob ), .a(dg), 
        .b(nda), .c(\twobitack[0] ), .d(\U1298/U1386/U25/U1/clr ) );
    inv_2 \U1298/U1386/U25/U1/Ui  ( .x(net193), .a(\U1298/U1386/U25/U1/ob ) );
    and2_1 \U1306/U1385/U8  ( .x(bg), .a(nbReset), .b(\U1306/ng ) );
    aoi222_1 \U1306/U1384/U30/U1  ( .x(\U1306/ng ), .a(nba), .b(\twobitack[1] 
        ), .c(nba), .d(\U1306/U1384/Z ), .e(\twobitack[1] ), .f(
        \U1306/U1384/Z ) );
    inv_1 \U1306/U1384/U30/Uinv  ( .x(\U1306/U1384/Z ), .a(\U1306/ng ) );
    oa31_1 \U1306/U1386/U25/U1/Uclr  ( .x(\U1306/U1386/U25/U1/clr ), .a(net199
        ), .b(bg), .c(nba), .d(\twobitack[1] ) );
    oaoi211_1 \U1306/U1386/U25/U1/Uaoi  ( .x(\U1306/U1386/U25/U1/ob ), .a(bg), 
        .b(nba), .c(net199), .d(\U1306/U1386/U25/U1/clr ) );
    inv_2 \U1306/U1386/U25/U1/Ui  ( .x(\twobitack[1] ), .a(
        \U1306/U1386/U25/U1/ob ) );
    and2_1 \U1295/U1385/U8  ( .x(ag), .a(nbReset), .b(\U1295/ng ) );
    aoi222_1 \U1295/U1384/U30/U1  ( .x(\U1295/ng ), .a(naa), .b(\twobitack[3] 
        ), .c(naa), .d(\U1295/U1384/Z ), .e(\twobitack[3] ), .f(
        \U1295/U1384/Z ) );
    inv_1 \U1295/U1384/U30/Uinv  ( .x(\U1295/U1384/Z ), .a(\U1295/ng ) );
    oa31_1 \U1295/U1386/U25/U1/Uclr  ( .x(\U1295/U1386/U25/U1/clr ), .a(net194
        ), .b(ag), .c(naa), .d(\twobitack[3] ) );
    oaoi211_1 \U1295/U1386/U25/U1/Uaoi  ( .x(\U1295/U1386/U25/U1/ob ), .a(ag), 
        .b(naa), .c(net194), .d(\U1295/U1386/U25/U1/clr ) );
    inv_2 \U1295/U1386/U25/U1/Ui  ( .x(\twobitack[3] ), .a(
        \U1295/U1386/U25/U1/ob ) );
    nand2_1 \U1297/U1131/U5  ( .x(\U1297/s ), .a(\U1297/r ), .b(\U1297/nback )
         );
    nand2_1 \U1297/U1103/U5  ( .x(\U1297/r ), .a(\U1297/naack ), .b(\U1297/s )
         );
    inv_1 \U1297/U1111/U3  ( .x(\U1297/reset ), .a(nbReset) );
    inv_1 \U1297/U1112/U3  ( .x(\U1297/naack ), .a(naa) );
    nor2_1 \U1297/U1130/U5  ( .x(\U1297/nback ), .a(nca), .b(\U1297/reset ) );
    aoai211_1 \U1297/U1128/U28/U1/U1  ( .x(\U1297/U1128/U28/U1/clr ), .a(
        \U1297/r ), .b(\U1297/naack ), .c(cg), .d(csel) );
    nand3_1 \U1297/U1128/U28/U1/U2  ( .x(\U1297/U1128/U28/U1/set ), .a(cg), 
        .b(\U1297/r ), .c(\U1297/naack ) );
    nand2_2 \U1297/U1128/U28/U1/U3  ( .x(csel), .a(\U1297/U1128/U28/U1/clr ), 
        .b(\U1297/U1128/U28/U1/set ) );
    aoai211_1 \U1297/U1127/U28/U1/U1  ( .x(\U1297/U1127/U28/U1/clr ), .a(
        \U1297/s ), .b(\U1297/nback ), .c(ag), .d(asel) );
    nand3_1 \U1297/U1127/U28/U1/U2  ( .x(\U1297/U1127/U28/U1/set ), .a(ag), 
        .b(\U1297/s ), .c(\U1297/nback ) );
    nand2_2 \U1297/U1127/U28/U1/U3  ( .x(asel), .a(\U1297/U1127/U28/U1/clr ), 
        .b(\U1297/U1127/U28/U1/set ) );
    nand2_1 \U1300/U1131/U5  ( .x(\U1300/s ), .a(\U1300/r ), .b(\U1300/nback )
         );
    nand2_1 \U1300/U1103/U5  ( .x(\U1300/r ), .a(\U1300/naack ), .b(\U1300/s )
         );
    inv_1 \U1300/U1111/U3  ( .x(\U1300/reset ), .a(nbReset) );
    inv_1 \U1300/U1112/U3  ( .x(\U1300/naack ), .a(nba) );
    nor2_1 \U1300/U1130/U5  ( .x(\U1300/nback ), .a(nda), .b(\U1300/reset ) );
    aoai211_1 \U1300/U1128/U28/U1/U1  ( .x(\U1300/U1128/U28/U1/clr ), .a(
        \U1300/r ), .b(\U1300/naack ), .c(dg), .d(dsel) );
    nand3_1 \U1300/U1128/U28/U1/U2  ( .x(\U1300/U1128/U28/U1/set ), .a(dg), 
        .b(\U1300/r ), .c(\U1300/naack ) );
    nand2_2 \U1300/U1128/U28/U1/U3  ( .x(dsel), .a(\U1300/U1128/U28/U1/clr ), 
        .b(\U1300/U1128/U28/U1/set ) );
    aoai211_1 \U1300/U1127/U28/U1/U1  ( .x(\U1300/U1127/U28/U1/clr ), .a(
        \U1300/s ), .b(\U1300/nback ), .c(bg), .d(bsel) );
    nand3_1 \U1300/U1127/U28/U1/U2  ( .x(\U1300/U1127/U28/U1/set ), .a(bg), 
        .b(\U1300/s ), .c(\U1300/nback ) );
    nand2_2 \U1300/U1127/U28/U1/U3  ( .x(bsel), .a(\U1300/U1127/U28/U1/clr ), 
        .b(\U1300/U1127/U28/U1/set ) );
    aoai211_1 \U1289/U1150/U28/U1/U1  ( .x(\U1289/U1150/U28/U1/clr ), .a(il[2]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdl[2] ) );
    nand3_1 \U1289/U1150/U28/U1/U2  ( .x(\U1289/U1150/U28/U1/set ), .a(net195), 
        .b(il[2]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1150/U28/U1/U3  ( .x(\cdl[2] ), .a(
        \U1289/U1150/U28/U1/clr ), .b(\U1289/U1150/U28/U1/set ) );
    aoai211_1 \U1289/U1152/U28/U1/U1  ( .x(\U1289/U1152/U28/U1/clr ), .a(il[3]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdl[3] ) );
    nand3_1 \U1289/U1152/U28/U1/U2  ( .x(\U1289/U1152/U28/U1/set ), .a(net195), 
        .b(il[3]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1152/U28/U1/U3  ( .x(\cdl[3] ), .a(
        \U1289/U1152/U28/U1/clr ), .b(\U1289/U1152/U28/U1/set ) );
    aoai211_1 \U1289/U1149/U28/U1/U1  ( .x(\U1289/U1149/U28/U1/clr ), .a(ih[2]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdh[2] ) );
    nand3_1 \U1289/U1149/U28/U1/U2  ( .x(\U1289/U1149/U28/U1/set ), .a(net195), 
        .b(ih[2]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1149/U28/U1/U3  ( .x(\cdh[2] ), .a(
        \U1289/U1149/U28/U1/clr ), .b(\U1289/U1149/U28/U1/set ) );
    aoai211_1 \U1289/U1151/U28/U1/U1  ( .x(\U1289/U1151/U28/U1/clr ), .a(ih[3]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdh[3] ) );
    nand3_1 \U1289/U1151/U28/U1/U2  ( .x(\U1289/U1151/U28/U1/set ), .a(net195), 
        .b(ih[3]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1151/U28/U1/U3  ( .x(\cdh[3] ), .a(
        \U1289/U1151/U28/U1/clr ), .b(\U1289/U1151/U28/U1/set ) );
    inv_1 \U1289/U1148/U1147/U3  ( .x(\U1289/U1148/net189 ), .a(
        \U1289/bnreset ) );
    nor2_1 \U1289/U1148/U582/U5  ( .x(\U1289/U1148/net192 ), .a(\cdl[3] ), .b(
        \cdh[3] ) );
    nor2_1 \U1289/U1148/U580/U5  ( .x(\U1289/U1148/net191 ), .a(\cdl[2] ), .b(
        \cdh[2] ) );
    nor2_2 \U1289/U1148/U1146/U6  ( .x(\twobitack[2] ), .a(
        \U1289/U1148/net190 ), .b(\U1289/U1148/net189 ) );
    aoi222_1 \U1289/U1148/U1141/U30/U1  ( .x(\U1289/U1148/net190 ), .a(
        \U1289/U1148/net191 ), .b(\U1289/U1148/net192 ), .c(
        \U1289/U1148/net191 ), .d(\U1289/U1148/U1141/Z ), .e(
        \U1289/U1148/net192 ), .f(\U1289/U1148/U1141/Z ) );
    inv_1 \U1289/U1148/U1141/U30/Uinv  ( .x(\U1289/U1148/U1141/Z ), .a(
        \U1289/U1148/net190 ) );
    aoai211_1 \U1271/U1150/U28/U1/U1  ( .x(\U1271/U1150/U28/U1/clr ), .a(il[0]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdl[0] ) );
    nand3_1 \U1271/U1150/U28/U1/U2  ( .x(\U1271/U1150/U28/U1/set ), .a(net193), 
        .b(il[0]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1150/U28/U1/U3  ( .x(\cdl[0] ), .a(
        \U1271/U1150/U28/U1/clr ), .b(\U1271/U1150/U28/U1/set ) );
    aoai211_1 \U1271/U1152/U28/U1/U1  ( .x(\U1271/U1152/U28/U1/clr ), .a(il[1]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdl[1] ) );
    nand3_1 \U1271/U1152/U28/U1/U2  ( .x(\U1271/U1152/U28/U1/set ), .a(net193), 
        .b(il[1]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1152/U28/U1/U3  ( .x(\cdl[1] ), .a(
        \U1271/U1152/U28/U1/clr ), .b(\U1271/U1152/U28/U1/set ) );
    aoai211_1 \U1271/U1149/U28/U1/U1  ( .x(\U1271/U1149/U28/U1/clr ), .a(ih[0]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdh[0] ) );
    nand3_1 \U1271/U1149/U28/U1/U2  ( .x(\U1271/U1149/U28/U1/set ), .a(net193), 
        .b(ih[0]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1149/U28/U1/U3  ( .x(\cdh[0] ), .a(
        \U1271/U1149/U28/U1/clr ), .b(\U1271/U1149/U28/U1/set ) );
    aoai211_1 \U1271/U1151/U28/U1/U1  ( .x(\U1271/U1151/U28/U1/clr ), .a(ih[1]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdh[1] ) );
    nand3_1 \U1271/U1151/U28/U1/U2  ( .x(\U1271/U1151/U28/U1/set ), .a(net193), 
        .b(ih[1]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1151/U28/U1/U3  ( .x(\cdh[1] ), .a(
        \U1271/U1151/U28/U1/clr ), .b(\U1271/U1151/U28/U1/set ) );
    inv_1 \U1271/U1148/U1147/U3  ( .x(\U1271/U1148/net189 ), .a(
        \U1271/bnreset ) );
    nor2_1 \U1271/U1148/U582/U5  ( .x(\U1271/U1148/net192 ), .a(\cdl[1] ), .b(
        \cdh[1] ) );
    nor2_1 \U1271/U1148/U580/U5  ( .x(\U1271/U1148/net191 ), .a(\cdl[0] ), .b(
        \cdh[0] ) );
    nor2_2 \U1271/U1148/U1146/U6  ( .x(\twobitack[0] ), .a(
        \U1271/U1148/net190 ), .b(\U1271/U1148/net189 ) );
    aoi222_1 \U1271/U1148/U1141/U30/U1  ( .x(\U1271/U1148/net190 ), .a(
        \U1271/U1148/net191 ), .b(\U1271/U1148/net192 ), .c(
        \U1271/U1148/net191 ), .d(\U1271/U1148/U1141/Z ), .e(
        \U1271/U1148/net192 ), .f(\U1271/U1148/U1141/Z ) );
    inv_1 \U1271/U1148/U1141/U30/Uinv  ( .x(\U1271/U1148/U1141/Z ), .a(
        \U1271/U1148/net190 ) );
    nand2_1 \U1225/U1128/U5  ( .x(\U1225/s ), .a(\U1225/r ), .b(\U1225/nback )
         );
    nand2_1 \U1225/U1103/U5  ( .x(\U1225/r ), .a(\U1225/naack ), .b(\U1225/s )
         );
    inv_1 \U1225/U1111/U3  ( .x(\U1225/reset ), .a(nbReset) );
    inv_1 \U1225/U1112/U3  ( .x(\U1225/naack ), .a(nxa) );
    nor2_1 \U1225/U1127/U5  ( .x(\U1225/nback ), .a(nyla), .b(\U1225/reset )
         );
    and2_2 \U1225/U1129/U8  ( .x(xsel), .a(\U1225/nback ), .b(\U1225/s ) );
    and2_2 \U1225/U1124/U8  ( .x(ysel), .a(\U1225/r ), .b(\U1225/naack ) );
    and3_4 \U1308/U20/U9  ( .x(nya), .a(\U1308/nack[1] ), .b(\U1308/nack[0] ), 
        .c(nbReset) );
    nor2_1 \U1308/U18/U5  ( .x(\U1308/nack[0] ), .a(\yl[3] ), .b(\yl[0] ) );
    nor2_1 \U1308/U19/U5  ( .x(\U1308/nack[1] ), .a(\yl[1] ), .b(\yl[2] ) );
    ao222_2 \U1308/U15_0_/U19/U1/U1  ( .x(\yl[0] ), .a(\y[0] ), .b(nyla), .c(
        \y[0] ), .d(\yl[0] ), .e(nyla), .f(\yl[0] ) );
    ao222_2 \U1308/U15_1_/U19/U1/U1  ( .x(\yl[1] ), .a(\y[1] ), .b(nyla), .c(
        \y[1] ), .d(\yl[1] ), .e(nyla), .f(\yl[1] ) );
    ao222_2 \U1308/U15_2_/U19/U1/U1  ( .x(\yl[2] ), .a(\y[2] ), .b(nyla), .c(
        \y[2] ), .d(\yl[2] ), .e(nyla), .f(\yl[2] ) );
    ao222_2 \U1308/U15_3_/U19/U1/U1  ( .x(\yl[3] ), .a(\y[3] ), .b(nyla), .c(
        \y[3] ), .d(\yl[3] ), .e(nyla), .f(\yl[3] ) );
    buf_3 U1 ( .x(\U1289/bnreset ), .a(nbReset) );
    buf_3 U2 ( .x(\U1271/bnreset ), .a(nbReset) );
endmodule


module chain_mergepackets_2 ( naa, nba, o, a, b, nReset, noa );
output [4:0] o;
input  [4:0] a;
input  [4:0] b;
input  nReset, noa;
output naa, nba;
    wire as, seta, asel, bsel, setb, reset, \noack[1] , \noack[0] , 
        \U916_0_/U25/U1/clr , \U916_0_/U25/U1/ob , \U916_1_/U25/U1/clr , 
        \U916_1_/U25/U1/ob , \U916_2_/U25/U1/clr , \U916_2_/U25/U1/ob , 
        \U916_3_/U25/U1/clr , \U916_3_/U25/U1/ob ;
    and2_1 \U1155/U8  ( .x(as), .a(seta), .b(asel) );
    nand2_1 \U1145/U5  ( .x(asel), .a(bsel), .b(seta) );
    nand2_1 \U1103/U5  ( .x(bsel), .a(setb), .b(asel) );
    inv_1 \U1135/U3  ( .x(reset), .a(nReset) );
    inv_1 \U1134/U3  ( .x(setb), .a(a[4]) );
    and3_2 \U1154/U9  ( .x(naa), .a(\noack[1] ), .b(\noack[0] ), .c(as) );
    nor3_1 \U1127/U7  ( .x(\noack[0] ), .a(o[1]), .b(reset), .c(o[0]) );
    nor2_1 \U1132/U5  ( .x(\noack[1] ), .a(o[3]), .b(o[2]) );
    oa31_1 \U916_0_/U25/U1/Uclr  ( .x(\U916_0_/U25/U1/clr ), .a(noa), .b(a[0]), 
        .c(b[0]), .d(o[0]) );
    oaoi211_1 \U916_0_/U25/U1/Uaoi  ( .x(\U916_0_/U25/U1/ob ), .a(a[0]), .b(b
        [0]), .c(noa), .d(\U916_0_/U25/U1/clr ) );
    inv_2 \U916_0_/U25/U1/Ui  ( .x(o[0]), .a(\U916_0_/U25/U1/ob ) );
    oa31_1 \U916_1_/U25/U1/Uclr  ( .x(\U916_1_/U25/U1/clr ), .a(noa), .b(a[1]), 
        .c(b[1]), .d(o[1]) );
    oaoi211_1 \U916_1_/U25/U1/Uaoi  ( .x(\U916_1_/U25/U1/ob ), .a(a[1]), .b(b
        [1]), .c(noa), .d(\U916_1_/U25/U1/clr ) );
    inv_2 \U916_1_/U25/U1/Ui  ( .x(o[1]), .a(\U916_1_/U25/U1/ob ) );
    oa31_1 \U916_2_/U25/U1/Uclr  ( .x(\U916_2_/U25/U1/clr ), .a(noa), .b(a[2]), 
        .c(b[2]), .d(o[2]) );
    oaoi211_1 \U916_2_/U25/U1/Uaoi  ( .x(\U916_2_/U25/U1/ob ), .a(a[2]), .b(b
        [2]), .c(noa), .d(\U916_2_/U25/U1/clr ) );
    inv_2 \U916_2_/U25/U1/Ui  ( .x(o[2]), .a(\U916_2_/U25/U1/ob ) );
    oa31_1 \U916_3_/U25/U1/Uclr  ( .x(\U916_3_/U25/U1/clr ), .a(noa), .b(a[3]), 
        .c(b[3]), .d(o[3]) );
    oaoi211_1 \U916_3_/U25/U1/Uaoi  ( .x(\U916_3_/U25/U1/ob ), .a(a[3]), .b(b
        [3]), .c(noa), .d(\U916_3_/U25/U1/clr ) );
    inv_2 \U916_3_/U25/U1/Ui  ( .x(o[3]), .a(\U916_3_/U25/U1/ob ) );
    ao222_2 \U1148/U19/U1/U1  ( .x(o[4]), .a(noa), .b(b[4]), .c(noa), .d(o[4]), 
        .e(b[4]), .f(o[4]) );
    aoi21_1 \U1153/U11  ( .x(seta), .a(o[4]), .b(setb), .c(reset) );
    and3_3 U1 ( .x(nba), .a(bsel), .b(\noack[0] ), .c(\noack[1] ) );
endmodule


module initiator_tic ( cack, chaincommand, err, nchainresponseack, nrouteack, 
    rd, routetxreq, rrnw, a, chainresponse, col, crnw, itag, lock, nReset, 
    nchaincommandack, pred, rack, route, routetxack, seq, size, wd );
output [4:0] chaincommand;
output [1:0] err;
output [63:0] rd;
output [1:0] rrnw;
input  [63:0] a;
input  [4:0] chainresponse;
input  [5:0] col;
input  [1:0] crnw;
input  [9:0] itag;
input  [1:0] lock;
input  [1:0] pred;
input  [4:0] route;
input  [1:0] seq;
input  [3:0] size;
input  [63:0] wd;
input  nReset, nchaincommandack, rack, routetxack;
output cack, nchainresponseack, nrouteack, routetxreq;
    wire nircba, nResetb, responseack, rstatusack, \irbl[7] , \irbl[6] , 
        \irbl[5] , \irbl[4] , \irbl[3] , \irbl[2] , \irbl[1] , \irbl[0] , 
        \irbh[7] , \irbh[6] , \irbh[5] , \irbh[4] , \irbh[3] , \irbh[2] , 
        \irbh[1] , \irbh[0] , \rstatus[1] , \rstatus[0] , ictrlack, 
        \can_defer[0] , net116, ncstatusack, pltxreq, tok_ack, \cstatus[0] , 
        \cstatus[1] , net115, net128, pltxack, icmdack, nicba, \icbl[7] , 
        \icbl[6] , \icbl[5] , \icbl[4] , \icbl[3] , \icbl[2] , \icbl[1] , 
        \icbl[0] , \icbh[7] , \icbh[6] , \icbh[5] , \icbh[4] , \icbh[3] , 
        \icbh[2] , \icbh[1] , \icbh[0] , nipayloadack, \ipayload[4] , 
        \ipayload[3] , \ipayload[2] , \ipayload[1] , \ipayload[0] , net170, 
        reset, net165, \U1662/U28/U1/clr , \U1662/U28/U1/set ;
    chain_irdemuxNew_2 U1442 ( .err(err), .ncback(nircba), .rd(rd), .rnw(rrnw), 
        .status({\rstatus[1] , \rstatus[0] }), .cbh({\irbh[7] , \irbh[6] , 
        \irbh[5] , \irbh[4] , \irbh[3] , \irbh[2] , \irbh[1] , \irbh[0] }), 
        .cbl({\irbl[7] , \irbl[6] , \irbl[5] , \irbl[4] , \irbl[3] , \irbl[2] , 
        \irbl[1] , \irbl[0] }), .nReset(nResetb), .nack(responseack), 
        .statusack(rstatusack) );
    chain_fr2dr_byte_5 chain_decoder ( .nia(nchainresponseack), .oh({\irbh[7] , 
        \irbh[6] , \irbh[5] , \irbh[4] , \irbh[3] , \irbh[2] , \irbh[1] , 
        \irbh[0] }), .ol({\irbl[7] , \irbl[6] , \irbl[5] , \irbl[4] , 
        \irbl[3] , \irbl[2] , \irbl[1] , \irbl[0] }), .i(chainresponse), 
        .nReset(nResetb), .noa(nircba) );
    chain_ic_ctrl_2 cmd_ctrl ( .ack(ictrlack), .candefer(\can_defer[0] ), 
        .eop(net116), .nstatack(ncstatusack), .pltxreq(pltxreq), .routetxreq(
        routetxreq), .tok_ack(tok_ack), .accept(\cstatus[0] ), .candefer_ack({
        1'b0, \can_defer[0] }), .defer(\cstatus[1] ), .eopack(net115), .lock(
        lock), .nReset(net128), .pltxack(pltxack), .routetxack(routetxack), 
        .tok_err(err[1]), .tok_ok(err[0]) );
    chain_icmux_2 cmd_mux ( .ack(icmdack), .chainh({\icbh[7] , \icbh[6] , 
        \icbh[5] , \icbh[4] , \icbh[3] , \icbh[2] , \icbh[1] , \icbh[0] }), 
        .chainl({\icbl[7] , \icbl[6] , \icbl[5] , \icbl[4] , \icbl[3] , 
        \icbl[2] , \icbl[1] , \icbl[0] }), .sendack(pltxack), .addr(a), .col(
        col), .itag(itag), .lock(lock), .nReset(net128), .nia(nicba), .pred(
        pred), .rnw(crnw), .sendreq(pltxreq), .seq(seq), .size(size), .wd(wd)
         );
    chain_dr2fr_byte_2 U1604 ( .eop_ack(net115), .ia(nicba), .o({\ipayload[4] , 
        \ipayload[3] , \ipayload[2] , \ipayload[1] , \ipayload[0] }), .eop(
        net116), .ih({\icbh[7] , \icbh[6] , \icbh[5] , \icbh[4] , \icbh[3] , 
        \icbh[2] , \icbh[1] , \icbh[0] }), .il({\icbl[7] , \icbl[6] , 
        \icbl[5] , \icbl[4] , \icbl[3] , \icbl[2] , \icbl[1] , \icbl[0] }), 
        .nReset(net128), .noa(nipayloadack) );
    chain_mergepackets_2 U1605 ( .naa(nrouteack), .nba(nipayloadack), .o(
        chaincommand), .a(route), .b({\ipayload[4] , \ipayload[3] , 
        \ipayload[2] , \ipayload[1] , \ipayload[0] }), .nReset(net128), .noa(
        nchaincommandack) );
    and2_1 U1676 ( .x(cack), .a(net170), .b(nResetb) );
    inv_4 \U1643/U3  ( .x(net128), .a(reset) );
    or2_4 \U1660/U12  ( .x(net165), .a(\cstatus[0] ), .b(\cstatus[1] ) );
    or2_1 \U1661/U12  ( .x(rstatusack), .a(net165), .b(reset) );
    ao222_2 \status_pipe_0_/U19/U1/U1  ( .x(\cstatus[0] ), .a(\rstatus[0] ), 
        .b(ncstatusack), .c(\rstatus[0] ), .d(\cstatus[0] ), .e(ncstatusack), 
        .f(\cstatus[0] ) );
    ao222_2 \status_pipe_1_/U19/U1/U1  ( .x(\cstatus[1] ), .a(\rstatus[1] ), 
        .b(ncstatusack), .c(\rstatus[1] ), .d(\cstatus[1] ), .e(ncstatusack), 
        .f(\cstatus[1] ) );
    ao222_1 \U1609/U18/U1/U1  ( .x(net170), .a(ictrlack), .b(icmdack), .c(
        ictrlack), .d(net170), .e(icmdack), .f(net170) );
    aoai211_1 \U1662/U28/U1/U1  ( .x(\U1662/U28/U1/clr ), .a(rack), .b(nResetb
        ), .c(tok_ack), .d(responseack) );
    nand3_1 \U1662/U28/U1/U2  ( .x(\U1662/U28/U1/set ), .a(tok_ack), .b(rack), 
        .c(nResetb) );
    nand2_2 \U1662/U28/U1/U3  ( .x(responseack), .a(\U1662/U28/U1/clr ), .b(
        \U1662/U28/U1/set ) );
    inv_2 U1 ( .x(reset), .a(nResetb) );
    buf_3 U2 ( .x(nResetb), .a(nReset) );
endmodule


module master_if_tic ( nReset, mc_req, mc_we, mc_mult, mc_prd, mc_seq, mc_ts, 
    mc_sel, mc_adr, mc_dat, mc_ack, mr_req, mr_we, mr_err, mr_rty, mr_acc, 
    mr_ts, mr_sel, mr_dat, mr_ack, chaincommand, nchaincommandack, 
    chainresponse, nchainresponseack, e_bare, e_dm, e_im, e_wish, r_bare, r_dm, 
    r_im, r_wish, tag_id, force_bare );
input  [2:0] mc_ts;
input  [3:0] mc_sel;
input  [31:0] mc_adr;
input  [31:0] mc_dat;
output [2:0] mr_ts;
output [3:0] mr_sel;
output [31:0] mr_dat;
output [4:0] chaincommand;
input  [4:0] chainresponse;
input  [3:0] e_bare;
input  [3:0] e_dm;
input  [3:0] e_im;
input  [3:0] e_wish;
input  [3:0] r_bare;
input  [3:0] r_dm;
input  [3:0] r_im;
input  [3:0] r_wish;
input  [4:0] tag_id;
input  nReset, mc_req, mc_we, mc_mult, mc_prd, mc_seq, mr_ack, 
    nchaincommandack, force_bare;
output mc_ack, mr_req, mr_we, mr_err, mr_rty, mr_acc, nchainresponseack;
    wire reset, ci_ack, ri_ack, \ri_rnw[1] , \ri_rnw[0] , \ri_err[1] , 
        \ri_err[0] , \ri_rd[63] , \ri_rd[62] , \ri_rd[61] , \ri_rd[60] , 
        \ri_rd[59] , \ri_rd[58] , \ri_rd[57] , \ri_rd[56] , \ri_rd[55] , 
        \ri_rd[54] , \ri_rd[53] , \ri_rd[52] , \ri_rd[51] , \ri_rd[50] , 
        \ri_rd[49] , \ri_rd[48] , \ri_rd[47] , \ri_rd[46] , \ri_rd[45] , 
        \ri_rd[44] , \ri_rd[43] , \ri_rd[42] , \ri_rd[41] , \ri_rd[40] , 
        \ri_rd[39] , \ri_rd[38] , \ri_rd[37] , \ri_rd[36] , \ri_rd[35] , 
        \ri_rd[34] , \ri_rd[33] , \ri_rd[32] , \ri_rd[31] , \ri_rd[30] , 
        \ri_rd[29] , \ri_rd[28] , \ri_rd[27] , \ri_rd[26] , \ri_rd[25] , 
        \ri_rd[24] , \ri_rd[23] , \ri_rd[22] , \ri_rd[21] , \ri_rd[20] , 
        \ri_rd[19] , \ri_rd[18] , \ri_rd[17] , \ri_rd[16] , \ri_rd[15] , 
        \ri_rd[14] , \ri_rd[13] , \ri_rd[12] , \ri_rd[11] , \ri_rd[10] , 
        \ri_rd[9] , \ri_rd[8] , \ri_rd[7] , \ri_rd[6] , \ri_rd[5] , \ri_rd[4] , 
        \ri_rd[3] , \ri_rd[2] , \ri_rd[1] , \ri_rd[0] , \ci_col[5] , 
        \ci_col[4] , \ci_col[3] , \ci_col[2] , \ci_col[1] , \ci_col[0] , 
        \ci_rnw[1] , \ci_rnw[0] , \ci_a[63] , \ci_a[62] , \ci_a[61] , 
        \ci_a[60] , \ci_a[59] , \ci_a[58] , \ci_a[57] , \ci_a[56] , \ci_a[55] , 
        \ci_a[54] , \ci_a[53] , \ci_a[52] , \ci_a[51] , \ci_a[50] , \ci_a[49] , 
        \ci_a[48] , \ci_a[47] , \ci_a[46] , \ci_a[45] , \ci_a[44] , \ci_a[43] , 
        \ci_a[42] , \ci_a[41] , \ci_a[40] , \ci_a[39] , \ci_a[38] , \ci_a[37] , 
        \ci_a[36] , \ci_a[35] , \ci_a[34] , \ci_a[33] , \ci_a[32] , \ci_a[31] , 
        \ci_a[30] , \ci_a[29] , \ci_a[28] , \ci_a[27] , \ci_a[26] , \ci_a[25] , 
        \ci_a[24] , \ci_a[23] , \ci_a[22] , \ci_a[21] , \ci_a[20] , \ci_a[19] , 
        \ci_a[18] , \ci_a[17] , \ci_a[16] , \ci_a[15] , \ci_a[14] , \ci_a[13] , 
        \ci_a[12] , \ci_a[11] , \ci_a[10] , \ci_a[9] , \ci_a[8] , \ci_a[7] , 
        \ci_a[6] , \ci_a[5] , \ci_a[4] , \ci_a[3] , \ci_a[2] , \ci_a[1] , 
        \ci_a[0] , \ci_lock[1] , \ci_lock[0] , \ci_wd[63] , \ci_wd[62] , 
        \ci_wd[61] , \ci_wd[60] , \ci_wd[59] , \ci_wd[58] , \ci_wd[57] , 
        \ci_wd[56] , \ci_wd[55] , \ci_wd[54] , \ci_wd[53] , \ci_wd[52] , 
        \ci_wd[51] , \ci_wd[50] , \ci_wd[49] , \ci_wd[48] , \ci_wd[47] , 
        \ci_wd[46] , \ci_wd[45] , \ci_wd[44] , \ci_wd[43] , \ci_wd[42] , 
        \ci_wd[41] , \ci_wd[40] , \ci_wd[39] , \ci_wd[38] , \ci_wd[37] , 
        \ci_wd[36] , \ci_wd[35] , \ci_wd[34] , \ci_wd[33] , \ci_wd[32] , 
        \ci_wd[31] , \ci_wd[30] , \ci_wd[29] , \ci_wd[28] , \ci_wd[27] , 
        \ci_wd[26] , \ci_wd[25] , \ci_wd[24] , \ci_wd[23] , \ci_wd[22] , 
        \ci_wd[21] , \ci_wd[20] , \ci_wd[19] , \ci_wd[18] , \ci_wd[17] , 
        \ci_wd[16] , \ci_wd[15] , \ci_wd[14] , \ci_wd[13] , \ci_wd[12] , 
        \ci_wd[11] , \ci_wd[10] , \ci_wd[9] , \ci_wd[8] , \ci_wd[7] , 
        \ci_wd[6] , \ci_wd[5] , \ci_wd[4] , \ci_wd[3] , \ci_wd[2] , \ci_wd[1] , 
        \ci_wd[0] , \ci_itag[9] , \ci_itag[8] , \ci_itag[7] , \ci_itag[6] , 
        \ci_itag[5] , \ci_itag[4] , \ci_itag[3] , \ci_itag[2] , \ci_itag[1] , 
        \ci_itag[0] , \ci_size[3] , \ci_size[2] , \ci_size[1] , \ci_size[0] , 
        \ci_pred[1] , \ci_pred[0] , \ci_seq[1] , \ci_seq[0] , \i_rl[3] , 
        \i_rl[2] , \i_rl[1] , \i_rl[0] , \i_rh[3] , \i_rh[2] , \i_rh[1] , 
        SYNOPSYS_UNCONNECTED_2, \i_el[3] , \i_el[2] , \i_el[1] , \i_el[0] , 
        SYNOPSYS_UNCONNECTED_1, \i_eh[2] , \i_eh[1] , \i_eh[0] , routetx_ack, 
        nroute_ack, routetx_req, \route[4] , SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4, \route[1] , \route[0] ;
    assign mr_rty = 1'b0;
    assign mr_acc = 1'b0;
    assign mr_ts[2] = 1'b0;
    assign mr_ts[1] = 1'b0;
    assign mr_ts[0] = 1'b0;
    inv_2 U1 ( .x(reset), .a(nReset) );
    m2cp_tic master2chainif ( .req_in(mc_req), .ts_o(mc_ts), .sel_o(mc_sel), 
        .mult_o(mc_mult), .we_o(mc_we), .prd_o(mc_prd), .seq_o(mc_seq), 
        .adr_o(mc_adr), .dat_o(mc_dat), .ain(mc_ack), .ic_seq({\ci_seq[1] , 
        \ci_seq[0] }), .ic_pred({\ci_pred[1] , \ci_pred[0] }), .ic_size({
        \ci_size[3] , \ci_size[2] , \ci_size[1] , \ci_size[0] }), .ic_itag({
        \ci_itag[9] , \ci_itag[8] , \ci_itag[7] , \ci_itag[6] , \ci_itag[5] , 
        \ci_itag[4] , \ci_itag[3] , \ci_itag[2] , \ci_itag[1] , \ci_itag[0] }), 
        .ic_wd({\ci_wd[63] , \ci_wd[62] , \ci_wd[61] , \ci_wd[60] , 
        \ci_wd[59] , \ci_wd[58] , \ci_wd[57] , \ci_wd[56] , \ci_wd[55] , 
        \ci_wd[54] , \ci_wd[53] , \ci_wd[52] , \ci_wd[51] , \ci_wd[50] , 
        \ci_wd[49] , \ci_wd[48] , \ci_wd[47] , \ci_wd[46] , \ci_wd[45] , 
        \ci_wd[44] , \ci_wd[43] , \ci_wd[42] , \ci_wd[41] , \ci_wd[40] , 
        \ci_wd[39] , \ci_wd[38] , \ci_wd[37] , \ci_wd[36] , \ci_wd[35] , 
        \ci_wd[34] , \ci_wd[33] , \ci_wd[32] , \ci_wd[31] , \ci_wd[30] , 
        \ci_wd[29] , \ci_wd[28] , \ci_wd[27] , \ci_wd[26] , \ci_wd[25] , 
        \ci_wd[24] , \ci_wd[23] , \ci_wd[22] , \ci_wd[21] , \ci_wd[20] , 
        \ci_wd[19] , \ci_wd[18] , \ci_wd[17] , \ci_wd[16] , \ci_wd[15] , 
        \ci_wd[14] , \ci_wd[13] , \ci_wd[12] , \ci_wd[11] , \ci_wd[10] , 
        \ci_wd[9] , \ci_wd[8] , \ci_wd[7] , \ci_wd[6] , \ci_wd[5] , \ci_wd[4] , 
        \ci_wd[3] , \ci_wd[2] , \ci_wd[1] , \ci_wd[0] }), .ic_lock({
        \ci_lock[1] , \ci_lock[0] }), .ic_a({\ci_a[63] , \ci_a[62] , 
        \ci_a[61] , \ci_a[60] , \ci_a[59] , \ci_a[58] , \ci_a[57] , \ci_a[56] , 
        \ci_a[55] , \ci_a[54] , \ci_a[53] , \ci_a[52] , \ci_a[51] , \ci_a[50] , 
        \ci_a[49] , \ci_a[48] , \ci_a[47] , \ci_a[46] , \ci_a[45] , \ci_a[44] , 
        \ci_a[43] , \ci_a[42] , \ci_a[41] , \ci_a[40] , \ci_a[39] , \ci_a[38] , 
        \ci_a[37] , \ci_a[36] , \ci_a[35] , \ci_a[34] , \ci_a[33] , \ci_a[32] , 
        \ci_a[31] , \ci_a[30] , \ci_a[29] , \ci_a[28] , \ci_a[27] , \ci_a[26] , 
        \ci_a[25] , \ci_a[24] , \ci_a[23] , \ci_a[22] , \ci_a[21] , \ci_a[20] , 
        \ci_a[19] , \ci_a[18] , \ci_a[17] , \ci_a[16] , \ci_a[15] , \ci_a[14] , 
        \ci_a[13] , \ci_a[12] , \ci_a[11] , \ci_a[10] , \ci_a[9] , \ci_a[8] , 
        \ci_a[7] , \ci_a[6] , \ci_a[5] , \ci_a[4] , \ci_a[3] , \ci_a[2] , 
        \ci_a[1] , \ci_a[0] }), .ic_rnw({\ci_rnw[1] , \ci_rnw[0] }), .ic_col({
        \ci_col[5] , \ci_col[4] , \ci_col[3] , \ci_col[2] , \ci_col[1] , 
        \ci_col[0] }), .ic_ack(ci_ack), .req_out(mr_req), .we_i(mr_we), 
        .err_i(mr_err), .dat_i(mr_dat), .aout(mr_ack), .ir_rd({\ri_rd[63] , 
        \ri_rd[62] , \ri_rd[61] , \ri_rd[60] , \ri_rd[59] , \ri_rd[58] , 
        \ri_rd[57] , \ri_rd[56] , \ri_rd[55] , \ri_rd[54] , \ri_rd[53] , 
        \ri_rd[52] , \ri_rd[51] , \ri_rd[50] , \ri_rd[49] , \ri_rd[48] , 
        \ri_rd[47] , \ri_rd[46] , \ri_rd[45] , \ri_rd[44] , \ri_rd[43] , 
        \ri_rd[42] , \ri_rd[41] , \ri_rd[40] , \ri_rd[39] , \ri_rd[38] , 
        \ri_rd[37] , \ri_rd[36] , \ri_rd[35] , \ri_rd[34] , \ri_rd[33] , 
        \ri_rd[32] , \ri_rd[31] , \ri_rd[30] , \ri_rd[29] , \ri_rd[28] , 
        \ri_rd[27] , \ri_rd[26] , \ri_rd[25] , \ri_rd[24] , \ri_rd[23] , 
        \ri_rd[22] , \ri_rd[21] , \ri_rd[20] , \ri_rd[19] , \ri_rd[18] , 
        \ri_rd[17] , \ri_rd[16] , \ri_rd[15] , \ri_rd[14] , \ri_rd[13] , 
        \ri_rd[12] , \ri_rd[11] , \ri_rd[10] , \ri_rd[9] , \ri_rd[8] , 
        \ri_rd[7] , \ri_rd[6] , \ri_rd[5] , \ri_rd[4] , \ri_rd[3] , \ri_rd[2] , 
        \ri_rd[1] , \ri_rd[0] }), .ir_err({\ri_err[1] , \ri_err[0] }), 
        .ir_rnw({\ri_rnw[1] , \ri_rnw[0] }), .ir_ack(ri_ack), .tag_id(tag_id), 
        .reset(reset) );
    i_adec_tic dec ( .e_h({SYNOPSYS_UNCONNECTED_1, \i_eh[2] , \i_eh[1] , 
        \i_eh[0] }), .e_l({\i_el[3] , \i_el[2] , \i_el[1] , \i_el[0] }), .r_h(
        {\i_rh[3] , \i_rh[2] , \i_rh[1] , SYNOPSYS_UNCONNECTED_2}), .r_l({
        \i_rl[3] , \i_rl[2] , \i_rl[1] , \i_rl[0] }), .ah({\ci_a[63] , 
        \ci_a[62] , \ci_a[61] , \ci_a[60] , \ci_a[59] , \ci_a[58] , \ci_a[57] , 
        \ci_a[56] , \ci_a[55] , \ci_a[54] , \ci_a[53] , \ci_a[52] , \ci_a[51] , 
        \ci_a[50] , \ci_a[49] , \ci_a[48] , \ci_a[47] , \ci_a[46] , \ci_a[45] , 
        \ci_a[44] , \ci_a[43] , \ci_a[42] , \ci_a[41] , \ci_a[40] , \ci_a[39] , 
        \ci_a[38] , \ci_a[37] , \ci_a[36] , \ci_a[35] , \ci_a[34] , \ci_a[33] , 
        \ci_a[32] }), .al({\ci_a[31] , \ci_a[30] , \ci_a[29] , \ci_a[28] , 
        \ci_a[27] , \ci_a[26] , \ci_a[25] , \ci_a[24] , \ci_a[23] , \ci_a[22] , 
        \ci_a[21] , \ci_a[20] , \ci_a[19] , \ci_a[18] , \ci_a[17] , \ci_a[16] , 
        \ci_a[15] , \ci_a[14] , \ci_a[13] , \ci_a[12] , \ci_a[11] , \ci_a[10] , 
        \ci_a[9] , \ci_a[8] , \ci_a[7] , \ci_a[6] , \ci_a[5] , \ci_a[4] , 
        \ci_a[3] , \ci_a[2] , \ci_a[1] , \ci_a[0] }), .e_bare(e_bare), .e_dm(
        e_dm), .e_im(e_im), .e_wish(e_wish), .r_bare(r_bare), .r_dm(r_dm), 
        .r_im(r_im), .r_wish(r_wish), .force_bare(force_bare) );
    route_tx_tic rt ( .o({\route[4] , SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4, \route[1] , \route[0] }), .rtxack(routetx_ack), 
        .e_h({1'b0, \i_eh[2] , \i_eh[1] , \i_eh[0] }), .e_l({\i_el[3] , 
        \i_el[2] , \i_el[1] , \i_el[0] }), .noa(nroute_ack), .r_h({\i_rh[3] , 
        \i_rh[2] , \i_rh[1] , 1'b0}), .r_l({\i_rl[3] , \i_rl[2] , \i_rl[1] , 
        \i_rl[0] }), .rtxreq(routetx_req) );
    initiator_tic it ( .cack(ci_ack), .chaincommand(chaincommand), .err({
        \ri_err[1] , \ri_err[0] }), .nchainresponseack(nchainresponseack), 
        .nrouteack(nroute_ack), .rd({\ri_rd[63] , \ri_rd[62] , \ri_rd[61] , 
        \ri_rd[60] , \ri_rd[59] , \ri_rd[58] , \ri_rd[57] , \ri_rd[56] , 
        \ri_rd[55] , \ri_rd[54] , \ri_rd[53] , \ri_rd[52] , \ri_rd[51] , 
        \ri_rd[50] , \ri_rd[49] , \ri_rd[48] , \ri_rd[47] , \ri_rd[46] , 
        \ri_rd[45] , \ri_rd[44] , \ri_rd[43] , \ri_rd[42] , \ri_rd[41] , 
        \ri_rd[40] , \ri_rd[39] , \ri_rd[38] , \ri_rd[37] , \ri_rd[36] , 
        \ri_rd[35] , \ri_rd[34] , \ri_rd[33] , \ri_rd[32] , \ri_rd[31] , 
        \ri_rd[30] , \ri_rd[29] , \ri_rd[28] , \ri_rd[27] , \ri_rd[26] , 
        \ri_rd[25] , \ri_rd[24] , \ri_rd[23] , \ri_rd[22] , \ri_rd[21] , 
        \ri_rd[20] , \ri_rd[19] , \ri_rd[18] , \ri_rd[17] , \ri_rd[16] , 
        \ri_rd[15] , \ri_rd[14] , \ri_rd[13] , \ri_rd[12] , \ri_rd[11] , 
        \ri_rd[10] , \ri_rd[9] , \ri_rd[8] , \ri_rd[7] , \ri_rd[6] , 
        \ri_rd[5] , \ri_rd[4] , \ri_rd[3] , \ri_rd[2] , \ri_rd[1] , \ri_rd[0] 
        }), .routetxreq(routetx_req), .rrnw({\ri_rnw[1] , \ri_rnw[0] }), .a({
        \ci_a[63] , \ci_a[62] , \ci_a[61] , \ci_a[60] , \ci_a[59] , \ci_a[58] , 
        \ci_a[57] , \ci_a[56] , \ci_a[55] , \ci_a[54] , \ci_a[53] , \ci_a[52] , 
        \ci_a[51] , \ci_a[50] , \ci_a[49] , \ci_a[48] , \ci_a[47] , \ci_a[46] , 
        \ci_a[45] , \ci_a[44] , \ci_a[43] , \ci_a[42] , \ci_a[41] , \ci_a[40] , 
        \ci_a[39] , \ci_a[38] , \ci_a[37] , \ci_a[36] , \ci_a[35] , \ci_a[34] , 
        \ci_a[33] , \ci_a[32] , \ci_a[31] , \ci_a[30] , \ci_a[29] , \ci_a[28] , 
        \ci_a[27] , \ci_a[26] , \ci_a[25] , \ci_a[24] , \ci_a[23] , \ci_a[22] , 
        \ci_a[21] , \ci_a[20] , \ci_a[19] , \ci_a[18] , \ci_a[17] , \ci_a[16] , 
        \ci_a[15] , \ci_a[14] , \ci_a[13] , \ci_a[12] , \ci_a[11] , \ci_a[10] , 
        \ci_a[9] , \ci_a[8] , \ci_a[7] , \ci_a[6] , \ci_a[5] , \ci_a[4] , 
        \ci_a[3] , \ci_a[2] , \ci_a[1] , \ci_a[0] }), .chainresponse(
        chainresponse), .col({\ci_col[5] , \ci_col[4] , \ci_col[3] , 
        \ci_col[2] , \ci_col[1] , \ci_col[0] }), .crnw({\ci_rnw[1] , 
        \ci_rnw[0] }), .itag({\ci_itag[9] , \ci_itag[8] , \ci_itag[7] , 
        \ci_itag[6] , \ci_itag[5] , \ci_itag[4] , \ci_itag[3] , \ci_itag[2] , 
        \ci_itag[1] , \ci_itag[0] }), .lock({\ci_lock[1] , \ci_lock[0] }), 
        .nReset(nReset), .nchaincommandack(nchaincommandack), .pred({
        \ci_pred[1] , \ci_pred[0] }), .rack(ri_ack), .route({\route[4] , 1'b0, 
        1'b0, \route[1] , \route[0] }), .routetxack(routetx_ack), .seq({
        \ci_seq[1] , \ci_seq[0] }), .size({\ci_size[3] , \ci_size[2] , 
        \ci_size[1] , \ci_size[0] }), .wd({\ci_wd[63] , \ci_wd[62] , 
        \ci_wd[61] , \ci_wd[60] , \ci_wd[59] , \ci_wd[58] , \ci_wd[57] , 
        \ci_wd[56] , \ci_wd[55] , \ci_wd[54] , \ci_wd[53] , \ci_wd[52] , 
        \ci_wd[51] , \ci_wd[50] , \ci_wd[49] , \ci_wd[48] , \ci_wd[47] , 
        \ci_wd[46] , \ci_wd[45] , \ci_wd[44] , \ci_wd[43] , \ci_wd[42] , 
        \ci_wd[41] , \ci_wd[40] , \ci_wd[39] , \ci_wd[38] , \ci_wd[37] , 
        \ci_wd[36] , \ci_wd[35] , \ci_wd[34] , \ci_wd[33] , \ci_wd[32] , 
        \ci_wd[31] , \ci_wd[30] , \ci_wd[29] , \ci_wd[28] , \ci_wd[27] , 
        \ci_wd[26] , \ci_wd[25] , \ci_wd[24] , \ci_wd[23] , \ci_wd[22] , 
        \ci_wd[21] , \ci_wd[20] , \ci_wd[19] , \ci_wd[18] , \ci_wd[17] , 
        \ci_wd[16] , \ci_wd[15] , \ci_wd[14] , \ci_wd[13] , \ci_wd[12] , 
        \ci_wd[11] , \ci_wd[10] , \ci_wd[9] , \ci_wd[8] , \ci_wd[7] , 
        \ci_wd[6] , \ci_wd[5] , \ci_wd[4] , \ci_wd[3] , \ci_wd[2] , \ci_wd[1] , 
        \ci_wd[0] }) );
endmodule


module command4Cycle ( ri, ao, _reset, ai, ro, l0, l1, l2 );
input  ri, ao, _reset;
output ai, ro, l0, l1, l2;
    wire _X21, csc0, _X20, _X18, _X19, _X14, csc1, _X13, _X23, _X17, n6, _X16, 
        _X22, _X11, n1, n2, n3, n4;
    and2_1 _U29 ( .x(_X21), .a(ri), .b(csc0) );
    and2_1 _U28 ( .x(_X20), .a(_X18), .b(_X19) );
    and2_1 _U18 ( .x(_X14), .a(l1), .b(csc1) );
    and2_1 _U17 ( .x(_X13), .a(l1), .b(_X19) );
    and2_1 _U32 ( .x(_X23), .a(ri), .b(csc1) );
    and2_1 _U23 ( .x(_X17), .a(n6), .b(csc0) );
    and2_1 _U22 ( .x(_X16), .a(n6), .b(_X19) );
    or3_2 _U33 ( .x(csc1), .a(_X22), .b(l0), .c(_X23) );
    and2_1 _U13 ( .x(_X11), .a(_X19), .b(l0) );
    or3i_1 U1 ( .x(n6), .a(n1), .b(_X17), .c(_X16) );
    or3i_1 U2 ( .x(csc0), .a(_X22), .b(_X21), .c(_X20) );
    inv_0 U4 ( .x(_X19), .a(ri) );
    nor2_0 U6 ( .x(ro), .a(_X19), .b(n2) );
    aoi21_1 U7 ( .x(n2), .a(_X18), .b(csc0), .c(ao) );
    aoi31_1 U8 ( .x(n3), .a(csc0), .b(n4), .c(csc1), .d(ao) );
    aoi22_1 U10 ( .x(ai), .a(n3), .b(n6), .c(csc0), .d(_X18) );
    inv_0 U12 ( .x(_X22), .a(l1) );
    inv_0 U13 ( .x(n4), .a(l0) );
    nor2i_1 U14 ( .x(n1), .a(_reset), .b(ao) );
    or3i_2 U15 ( .x(l1), .a(n1), .b(_X14), .c(_X13) );
    inv_1 U16 ( .x(l2), .a(_X18) );
    inv_2 U17 ( .x(_X18), .a(n6) );
    nand2i_2 U18 ( .x(l0), .a(_X11), .b(n1) );
endmodule


module matched_delay_tic_com ( x, a );
input  a;
output x;
    assign x = a;
endmodule


module response4Cycle ( ri, ao, _reset, ai, ro, l0, l1, l2, l3 );
input  ri, ao, _reset;
output ai, ro, l0, l1, l2, l3;
    wire l3_csc0_reset, _reset__not, n4, n3, _X13, n2, csc0, csc2__reset, csc2, 
        _X26, _X25, csc1__reset, csc1, _X35, _X7, _X37, _X36, _X31, _X30, _X10, 
        _X9, _X8, _X14, _X11, _X18, _X16, _X20, _X21, csc0__reset, n5, n6, n7, 
        n10, n8, n9;
    or2_2 _U44 ( .x(l3_csc0_reset), .a(_reset__not), .b(l3) );
    and2_1 _U22_4 ( .x(n4), .a(n3), .b(_X13) );
    and2_1 _U22_3 ( .x(n3), .a(n2), .b(csc0) );
    and2_1 _U24 ( .x(csc2__reset), .a(_reset), .b(csc2) );
    and2_1 _U41 ( .x(_X26), .a(csc0), .b(_X25) );
    and2_1 _U57 ( .x(csc1__reset), .a(_reset), .b(csc1) );
    and2_1 _U53 ( .x(_X35), .a(_X7), .b(csc2) );
    and2_1 _U54 ( .x(_X37), .a(_X36), .b(csc2) );
    and2_1 _U47 ( .x(_X31), .a(csc1), .b(_X30) );
    and3_1 _U16 ( .x(_X10), .a(ri), .b(_X9), .c(csc1) );
    and2_1 _U15 ( .x(_X8), .a(_X7), .b(l0) );
    and2_1 _U22_5 ( .x(_X14), .a(n4), .b(csc1) );
    and2_1 _U21 ( .x(_X11), .a(l1), .b(csc2__reset) );
    and2_1 _U28 ( .x(_X18), .a(l2), .b(_X16) );
    and2_1 _U33 ( .x(_X20), .a(_X7), .b(l3) );
    and2_1 _U34 ( .x(_X21), .a(csc0__reset), .b(l3) );
    oai222_1 U1 ( .x(ro), .a(_X13), .b(n5), .c(_reset__not), .d(n6), .e(csc1), 
        .f(csc0) );
    inv_0 U2 ( .x(_reset__not), .a(_reset) );
    oai21_1 U3 ( .x(csc2), .a(csc1__reset), .b(_X7), .c(n7) );
    nor2_0 U4 ( .x(_X36), .a(_X14), .b(_X11) );
    ao21_1 U7 ( .x(csc0), .a(n10), .b(n8), .c(_X26) );
    inv_0 U9 ( .x(_X25), .a(l3_csc0_reset) );
    and3i_1 U11 ( .x(n2), .a(ao), .b(ri), .c(csc2__reset) );
    oa21_1 U12 ( .x(ai), .a(l3), .b(_X9), .c(ro) );
    nor3_0 U13 ( .x(n6), .a(l3), .b(l1), .c(l2) );
    nand2_0 U15 ( .x(n5), .a(csc0), .b(_reset) );
    nor2_0 U16 ( .x(n7), .a(_X35), .b(_X37) );
    inv_0 U17 ( .x(n8), .a(ao) );
    inv_0 U18 ( .x(csc0__reset), .a(n5) );
    inv_0 U20 ( .x(_X9), .a(csc0) );
    inv_0 U22 ( .x(_X16), .a(csc2) );
    inv_0 U23 ( .x(_X30), .a(l2) );
    nand3i_0 U24 ( .x(n9), .a(csc1), .b(_X30), .c(_X7) );
    nand2i_2 U25 ( .x(csc1), .a(_X31), .b(ri) );
    nor2_1 U26 ( .x(_X7), .a(ao), .b(_reset__not) );
    ao21_2 U27 ( .x(l2), .a(_X16), .b(n8), .c(_X18) );
    inv_2 U28 ( .x(l1), .a(_X36) );
    or3i_2 U29 ( .x(l3), .a(n9), .b(_X20), .c(_X21) );
    inv_0 U30 ( .x(n10), .a(_X13) );
    inv_1 U31 ( .x(l0), .a(_X13) );
    nor2_1 U32 ( .x(_X13), .a(_X10), .b(_X8) );
endmodule


module matched_delay_tic_resp ( x, a );
input  a;
output x;
    assign x = a;
endmodule


module tic ( c_req, c_ack, c_we, c_addr, r_req, r_ack, data_in, data_out, 
    reset_b, mc_req, mc_we, mc_adr, mc_dat, mc_ack, mr_req, mr_dat, mr_ack );
input  [10:0] c_addr;
input  [7:0] data_in;
output [7:0] data_out;
output [31:0] mc_adr;
output [31:0] mc_dat;
input  [31:0] mr_dat;
input  c_req, c_we, r_ack, reset_b, mc_ack, mr_req;
output c_ack, r_req, mc_req, mc_we, mr_ack;
    wire c_addr_10, c_addr_9, c_addr_8, c_addr_7, c_addr_6, c_addr_5, c_addr_4, 
        c_addr_3, c_addr_2, c_addr_1, c_addr_0, data_in_7, data_in_6, 
        data_in_5, data_in_4, data_in_3, data_in_2, data_in_1, data_in_0, cwr, 
        wr_ack, w_r, wl0, wl1, wl2, _66_net_, rrr, rd_ack, r_r, \s[0] , \s[1] , 
        \s[2] , \s[3] , _67_net_, \covResp/nh , rwr, \covResp/nl , 
        \convCom/nh , \convCom/nl , crr, \covResp/ni ;
    assign mc_we = c_we;
    assign c_addr_10 = c_addr[10];
    assign c_addr_9 = c_addr[9];
    assign c_addr_8 = c_addr[8];
    assign c_addr_7 = c_addr[7];
    assign c_addr_6 = c_addr[6];
    assign c_addr_5 = c_addr[5];
    assign c_addr_4 = c_addr[4];
    assign c_addr_3 = c_addr[3];
    assign c_addr_2 = c_addr[2];
    assign c_addr_1 = c_addr[1];
    assign c_addr_0 = c_addr[0];
    assign data_in_7 = data_in[7];
    assign data_in_6 = data_in[6];
    assign data_in_5 = data_in[5];
    assign data_in_4 = data_in[4];
    assign data_in_3 = data_in[3];
    assign data_in_2 = data_in[2];
    assign data_in_1 = data_in[1];
    assign data_in_0 = data_in[0];
    assign mc_adr[31] = c_addr_10;
    assign mc_adr[30] = c_addr_10;
    assign mc_adr[29] = 1'b0;
    assign mc_adr[28] = 1'b0;
    assign mc_adr[27] = 1'b0;
    assign mc_adr[26] = 1'b0;
    assign mc_adr[25] = 1'b0;
    assign mc_adr[24] = 1'b0;
    assign mc_adr[23] = 1'b0;
    assign mc_adr[22] = 1'b0;
    assign mc_adr[21] = 1'b0;
    assign mc_adr[20] = 1'b0;
    assign mc_adr[19] = 1'b0;
    assign mc_adr[18] = 1'b0;
    assign mc_adr[17] = 1'b0;
    assign mc_adr[16] = 1'b0;
    assign mc_adr[15] = 1'b0;
    assign mc_adr[14] = 1'b0;
    assign mc_adr[13] = 1'b0;
    assign mc_adr[12] = 1'b0;
    assign mc_adr[11] = c_addr_9;
    assign mc_adr[10] = c_addr_8;
    assign mc_adr[9] = c_addr_7;
    assign mc_adr[8] = c_addr_6;
    assign mc_adr[7] = c_addr_5;
    assign mc_adr[6] = c_addr_4;
    assign mc_adr[5] = c_addr_3;
    assign mc_adr[4] = c_addr_2;
    assign mc_adr[3] = c_addr_1;
    assign mc_adr[2] = c_addr_0;
    assign mc_adr[1] = 1'b0;
    assign mc_adr[0] = 1'b0;
    assign mc_dat[31] = data_in_7;
    assign mc_dat[30] = data_in_6;
    assign mc_dat[29] = data_in_5;
    assign mc_dat[28] = data_in_4;
    assign mc_dat[27] = data_in_3;
    assign mc_dat[26] = data_in_2;
    assign mc_dat[25] = data_in_1;
    assign mc_dat[24] = data_in_0;
    command4Cycle cc ( .ri(cwr), .ao(mc_ack), ._reset(reset_b), .ai(wr_ack), 
        .ro(w_r), .l0(wl0), .l1(wl1), .l2(wl2) );
    matched_delay_tic_com delCom ( .x(mc_req), .a(_66_net_) );
    response4Cycle rc ( .ri(rrr), .ao(r_ack), ._reset(reset_b), .ai(rd_ack), 
        .ro(r_r), .l0(\s[0] ), .l1(\s[1] ), .l2(\s[2] ), .l3(\s[3] ) );
    matched_delay_tic_resp delResp ( .x(r_req), .a(_67_net_) );
    inv_1 \covResp/Uih  ( .x(\covResp/nh ), .a(rwr) );
    inv_1 \covResp/Uil  ( .x(\covResp/nl ), .a(rrr) );
    inv_1 \convCom/Uih  ( .x(\convCom/nh ), .a(cwr) );
    inv_1 \convCom/Uil  ( .x(\convCom/nl ), .a(crr) );
    ao23_2 \covResp/Ucl/U1/U1  ( .x(rrr), .a(mr_req), .b(rrr), .c(mr_req), .d(
        \covResp/ni ), .e(\covResp/nh ) );
    ao23_2 \convCom/Ucl/U1/U1  ( .x(crr), .a(c_req), .b(crr), .c(c_req), .d(
        \covResp/ni ), .e(\convCom/nh ) );
    ao23_2 \convCom/Uch/U1/U1  ( .x(cwr), .a(c_req), .b(cwr), .c(c_req), .d(
        mc_we), .e(\convCom/nl ) );
    ao23_2 \covResp/Uch/U1/U1  ( .x(rwr), .a(mr_req), .b(rwr), .c(mr_req), .d(
        mc_we), .e(\covResp/nl ) );
    latn_2 \wd1_reg[7]  ( .q(mc_dat[15]), .d(data_in_7), .g(wl1) );
    latn_2 \wd1_reg[6]  ( .q(mc_dat[14]), .d(data_in_6), .g(wl1) );
    latn_2 \wd1_reg[5]  ( .q(mc_dat[13]), .d(data_in_5), .g(wl1) );
    latn_2 \wd1_reg[4]  ( .q(mc_dat[12]), .d(data_in_4), .g(wl1) );
    latn_2 \wd1_reg[3]  ( .q(mc_dat[11]), .d(data_in_3), .g(wl1) );
    latn_2 \wd1_reg[2]  ( .q(mc_dat[10]), .d(data_in_2), .g(wl1) );
    latn_2 \wd1_reg[1]  ( .q(mc_dat[9]), .d(data_in_1), .g(wl1) );
    latn_2 \wd1_reg[0]  ( .q(mc_dat[8]), .d(data_in_0), .g(wl1) );
    latn_1 \wd0_reg[6]  ( .q(mc_dat[6]), .d(data_in_6), .g(wl0) );
    latn_1 \wd0_reg[7]  ( .q(mc_dat[7]), .d(data_in_7), .g(wl0) );
    latn_1 \wd0_reg[2]  ( .q(mc_dat[2]), .d(data_in_2), .g(wl0) );
    latn_1 \wd0_reg[5]  ( .q(mc_dat[5]), .d(data_in_5), .g(wl0) );
    latn_1 \wd0_reg[1]  ( .q(mc_dat[1]), .d(data_in_1), .g(wl0) );
    latn_2 \wd0_reg[4]  ( .q(mc_dat[4]), .d(data_in_4), .g(wl0) );
    latn_2 \wd0_reg[3]  ( .q(mc_dat[3]), .d(data_in_3), .g(wl0) );
    latn_2 \wd0_reg[0]  ( .q(mc_dat[0]), .d(data_in_0), .g(wl0) );
    inv_0 U2 ( .x(\covResp/ni ), .a(mc_we) );
    or2_1 U3 ( .x(_67_net_), .a(r_r), .b(rwr) );
    ao21_1 U4 ( .x(mr_ack), .a(rwr), .b(r_ack), .c(rd_ack) );
    or2_1 U5 ( .x(_66_net_), .a(crr), .b(w_r) );
    ao21_1 U6 ( .x(c_ack), .a(crr), .b(mc_ack), .c(wr_ack) );
    mx4_1 U7 ( .x(data_out[0]), .d0(mr_dat[0]), .sl0(\s[0] ), .d1(mr_dat[8]), 
        .sl1(\s[1] ), .d2(mr_dat[16]), .sl2(\s[2] ), .d3(mr_dat[24]), .sl3(
        \s[3] ) );
    mx4_1 U8 ( .x(data_out[1]), .d0(mr_dat[1]), .sl0(\s[0] ), .d1(mr_dat[9]), 
        .sl1(\s[1] ), .d2(mr_dat[17]), .sl2(\s[2] ), .d3(mr_dat[25]), .sl3(
        \s[3] ) );
    mx4_1 U9 ( .x(data_out[2]), .d0(mr_dat[2]), .sl0(\s[0] ), .d1(mr_dat[10]), 
        .sl1(\s[1] ), .d2(mr_dat[18]), .sl2(\s[2] ), .d3(mr_dat[26]), .sl3(
        \s[3] ) );
    mx4_1 U10 ( .x(data_out[3]), .d0(mr_dat[3]), .sl0(\s[0] ), .d1(mr_dat[11]), 
        .sl1(\s[1] ), .d2(mr_dat[19]), .sl2(\s[2] ), .d3(mr_dat[27]), .sl3(
        \s[3] ) );
    mx4_1 U11 ( .x(data_out[4]), .d0(mr_dat[4]), .sl0(\s[0] ), .d1(mr_dat[12]), 
        .sl1(\s[1] ), .d2(mr_dat[20]), .sl2(\s[2] ), .d3(mr_dat[28]), .sl3(
        \s[3] ) );
    mx4_1 U12 ( .x(data_out[5]), .d0(mr_dat[5]), .sl0(\s[0] ), .d1(mr_dat[13]), 
        .sl1(\s[1] ), .d2(mr_dat[21]), .sl2(\s[2] ), .d3(mr_dat[29]), .sl3(
        \s[3] ) );
    mx4_1 U13 ( .x(data_out[6]), .d0(mr_dat[6]), .sl0(\s[0] ), .d1(mr_dat[14]), 
        .sl1(\s[1] ), .d2(mr_dat[22]), .sl2(\s[2] ), .d3(mr_dat[30]), .sl3(
        \s[3] ) );
    mx4_1 U14 ( .x(data_out[7]), .d0(\s[0] ), .sl0(mr_dat[7]), .d1(\s[1] ), 
        .sl1(mr_dat[15]), .d2(\s[2] ), .sl2(mr_dat[23]), .d3(\s[3] ), .sl3(
        mr_dat[31]) );
    latn_1 \wd2_reg[6]  ( .q(mc_dat[22]), .d(data_in_6), .g(wl2) );
    latn_1 \wd2_reg[7]  ( .q(mc_dat[23]), .d(data_in_7), .g(wl2) );
    latn_1 \wd2_reg[0]  ( .q(mc_dat[16]), .d(data_in_0), .g(wl2) );
    latn_1 \wd2_reg[1]  ( .q(mc_dat[17]), .d(data_in_1), .g(wl2) );
    latn_1 \wd2_reg[3]  ( .q(mc_dat[19]), .d(data_in_3), .g(wl2) );
    latn_1 \wd2_reg[2]  ( .q(mc_dat[18]), .d(data_in_2), .g(wl2) );
    latn_1 \wd2_reg[5]  ( .q(mc_dat[21]), .d(data_in_5), .g(wl2) );
    latn_1 \wd2_reg[4]  ( .q(mc_dat[20]), .d(data_in_4), .g(wl2) );
endmodule


module chain_arbiter0 ( eop_ix, d0_ix, d1_ix, d2_ix, d3_ix, ack_ix, eop_iy, 
    d0_iy, d1_iy, d2_iy, d3_iy, ack_iy, eop_ox, d0_ox, d1_ox, d2_ox, d3_ox, 
    eop_oy, d0_oy, d1_oy, d2_oy, d3_oy, ack_oxy, rst, test_si, test_se, 
    test_so, phi1, phi2, phi3 );
input  eop_ix, d0_ix, d1_ix, d2_ix, d3_ix, eop_iy, d0_iy, d1_iy, d2_iy, d3_iy, 
    ack_oxy, rst, test_si, test_se, phi1, phi2, phi3;
output ack_ix, ack_iy, eop_ox, d0_ox, d1_ox, d2_ox, d3_ox, eop_oy, d0_oy, 
    d1_oy, d2_oy, d3_oy, test_so;
    wire nack_x, ackx_l, n1x, n2x, nack_y, acky_l, n1y, n2y, req_x, n5x, n6x, 
        req_y, n5y, n6y, sx_pl, gx, sy_pl, gy, \cye/nr , sy, \cye/nd , 
        \cye/n2 , \cy3/__tmp99/loop , \cy2/__tmp99/loop , \cy1/__tmp99/loop , 
        \cy0/__tmp99/loop , \cxe/nr , sx, \cxe/nd , \cxe/n2 , 
        \cx3/__tmp99/loop , \cx2/__tmp99/loop , \cx1/__tmp99/loop , 
        \cx0/__tmp99/loop , \mtx/gr2 , mry, \mtx/gr1 , mrx, \sry/qz , \srx/qz , 
        \sl_sy/l1_q , \scan[1] , \sl_sy/mxl/muxout , \scan[0] , \sl_sx/l1_q , 
        \sl_sx/mxl/muxout , \slAcky/l1_q , \slAcky/mxl/muxout , \scan[2] , 
        \slAckx/l1_q , \slAckx/mxl/muxout ;
    nor2_2 U12 ( .x(nack_x), .a(ackx_l), .b(rst) );
    nand2_1 U4 ( .x(ack_ix), .a(n1x), .b(n2x) );
    nor3_1 U17 ( .x(n1x), .a(d2_ox), .b(d3_ox), .c(d1_ox) );
    nor2_1 U18 ( .x(n2x), .a(eop_ox), .b(d0_ox) );
    nor2_2 U11 ( .x(nack_y), .a(acky_l), .b(rst) );
    nand2_1 U3 ( .x(ack_iy), .a(n1y), .b(n2y) );
    nor3_1 U16 ( .x(n1y), .a(d2_oy), .b(d3_oy), .c(d1_oy) );
    nor2_1 U19 ( .x(n2y), .a(eop_oy), .b(d0_oy) );
    nand2_1 U15 ( .x(req_x), .a(n5x), .b(n6x) );
    nor3_1 U10 ( .x(n5x), .a(d2_ix), .b(d3_ix), .c(d1_ix) );
    nor2_1 U13 ( .x(n6x), .a(eop_ix), .b(d0_ix) );
    nand2_1 U14 ( .x(req_y), .a(n5y), .b(n6y) );
    nor3_1 U9 ( .x(n5y), .a(d2_iy), .b(d3_iy), .c(d1_iy) );
    nor2_1 U20 ( .x(n6y), .a(eop_iy), .b(d0_iy) );
    nor2i_1 U6 ( .x(sx_pl), .a(gx), .b(eop_oy) );
    nor2i_1 U5 ( .x(sy_pl), .a(gy), .b(eop_ox) );
    nor3_1 \cye/Unr  ( .x(\cye/nr ), .a(eop_iy), .b(nack_y), .c(sy) );
    nand3_1 \cye/Und  ( .x(\cye/nd ), .a(eop_iy), .b(nack_y), .c(sy) );
    oa21_1 \cye/U1  ( .x(\cye/n2 ), .a(\cye/n2 ), .b(\cye/nr ), .c(\cye/nd )
         );
    inv_1 \cye/U3  ( .x(eop_oy), .a(\cye/n2 ) );
    ao31_1 \cy3/__tmp99/aoi  ( .x(\cy3/__tmp99/loop ), .a(d3_iy), .b(nack_y), 
        .c(sy), .d(d3_oy) );
    oa21_1 \cy3/__tmp99/outGate  ( .x(d3_oy), .a(d3_iy), .b(nack_y), .c(
        \cy3/__tmp99/loop ) );
    ao31_1 \cy2/__tmp99/aoi  ( .x(\cy2/__tmp99/loop ), .a(d2_iy), .b(nack_y), 
        .c(sy), .d(d2_oy) );
    oa21_1 \cy2/__tmp99/outGate  ( .x(d2_oy), .a(d2_iy), .b(nack_y), .c(
        \cy2/__tmp99/loop ) );
    ao31_1 \cy1/__tmp99/aoi  ( .x(\cy1/__tmp99/loop ), .a(d1_iy), .b(nack_y), 
        .c(sy), .d(d1_oy) );
    oa21_1 \cy1/__tmp99/outGate  ( .x(d1_oy), .a(d1_iy), .b(nack_y), .c(
        \cy1/__tmp99/loop ) );
    ao31_1 \cy0/__tmp99/aoi  ( .x(\cy0/__tmp99/loop ), .a(d0_iy), .b(nack_y), 
        .c(sy), .d(d0_oy) );
    oa21_1 \cy0/__tmp99/outGate  ( .x(d0_oy), .a(d0_iy), .b(nack_y), .c(
        \cy0/__tmp99/loop ) );
    nor3_1 \cxe/Unr  ( .x(\cxe/nr ), .a(eop_ix), .b(nack_x), .c(sx) );
    nand3_1 \cxe/Und  ( .x(\cxe/nd ), .a(eop_ix), .b(nack_x), .c(sx) );
    oa21_1 \cxe/U1  ( .x(\cxe/n2 ), .a(\cxe/n2 ), .b(\cxe/nr ), .c(\cxe/nd )
         );
    inv_1 \cxe/U3  ( .x(eop_ox), .a(\cxe/n2 ) );
    ao31_1 \cx3/__tmp99/aoi  ( .x(\cx3/__tmp99/loop ), .a(d3_ix), .b(nack_x), 
        .c(sx), .d(d3_ox) );
    oa21_1 \cx3/__tmp99/outGate  ( .x(d3_ox), .a(d3_ix), .b(nack_x), .c(
        \cx3/__tmp99/loop ) );
    ao31_1 \cx2/__tmp99/aoi  ( .x(\cx2/__tmp99/loop ), .a(d2_ix), .b(nack_x), 
        .c(sx), .d(d2_ox) );
    oa21_1 \cx2/__tmp99/outGate  ( .x(d2_ox), .a(d2_ix), .b(nack_x), .c(
        \cx2/__tmp99/loop ) );
    ao31_1 \cx1/__tmp99/aoi  ( .x(\cx1/__tmp99/loop ), .a(d1_ix), .b(nack_x), 
        .c(sx), .d(d1_ox) );
    oa21_1 \cx1/__tmp99/outGate  ( .x(d1_ox), .a(d1_ix), .b(nack_x), .c(
        \cx1/__tmp99/loop ) );
    ao31_1 \cx0/__tmp99/aoi  ( .x(\cx0/__tmp99/loop ), .a(d0_ix), .b(nack_x), 
        .c(sx), .d(d0_ox) );
    oa21_1 \cx0/__tmp99/outGate  ( .x(d0_ox), .a(d0_ix), .b(nack_x), .c(
        \cx0/__tmp99/loop ) );
    nand2_1 \mtx/mg2  ( .x(\mtx/gr2 ), .a(mry), .b(\mtx/gr1 ) );
    nand2_1 \mtx/U1  ( .x(\mtx/gr1 ), .a(mrx), .b(\mtx/gr2 ) );
    nor3_1 \mtx/U2  ( .x(gy), .a(\mtx/gr2 ), .b(\mtx/gr2 ), .c(\mtx/gr2 ) );
    nor3_1 \mtx/U3  ( .x(gx), .a(\mtx/gr1 ), .b(\mtx/gr1 ), .c(\mtx/gr1 ) );
    nor2_1 \sry/i1  ( .x(\sry/qz ), .a(req_y), .b(mry) );
    nor2_1 \srx/i1  ( .x(\srx/qz ), .a(req_x), .b(mrx) );
    latn_1 \sl_sy/lph3  ( .q(sy), .d(\sl_sy/l1_q ), .g(phi3) );
    latn_1 \sl_sy/lph2  ( .q(\scan[1] ), .d(\sl_sy/l1_q ), .g(phi2) );
    mux2_1 \sl_sy/mxl/mux  ( .x(\sl_sy/mxl/muxout ), .d0(sy_pl), .sl(test_se), 
        .d1(\scan[0] ) );
    latn_1 \sl_sy/mxl/lph1  ( .q(\sl_sy/l1_q ), .d(\sl_sy/mxl/muxout ), .g(
        phi1) );
    latn_1 \sl_sx/lph3  ( .q(sx), .d(\sl_sx/l1_q ), .g(phi3) );
    latn_1 \sl_sx/lph2  ( .q(\scan[0] ), .d(\sl_sx/l1_q ), .g(phi2) );
    mux2_1 \sl_sx/mxl/mux  ( .x(\sl_sx/mxl/muxout ), .d0(sx_pl), .sl(test_se), 
        .d1(test_si) );
    latn_1 \sl_sx/mxl/lph1  ( .q(\sl_sx/l1_q ), .d(\sl_sx/mxl/muxout ), .g(
        phi1) );
    latn_1 \slAcky/lph3  ( .q(acky_l), .d(\slAcky/l1_q ), .g(phi3) );
    latn_1 \slAcky/lph2  ( .q(test_so), .d(\slAcky/l1_q ), .g(phi2) );
    mux2_1 \slAcky/mxl/mux  ( .x(\slAcky/mxl/muxout ), .d0(ack_oxy), .sl(
        test_se), .d1(\scan[2] ) );
    latn_1 \slAcky/mxl/lph1  ( .q(\slAcky/l1_q ), .d(\slAcky/mxl/muxout ), .g(
        phi1) );
    latn_1 \slAckx/lph3  ( .q(ackx_l), .d(\slAckx/l1_q ), .g(phi3) );
    latn_1 \slAckx/lph2  ( .q(\scan[2] ), .d(\slAckx/l1_q ), .g(phi2) );
    mux2_1 \slAckx/mxl/mux  ( .x(\slAckx/mxl/muxout ), .d0(ack_oxy), .sl(
        test_se), .d1(\scan[1] ) );
    latn_1 \slAckx/mxl/lph1  ( .q(\slAckx/l1_q ), .d(\slAckx/mxl/muxout ), .g(
        phi1) );
    nor3_0 U1 ( .x(mrx), .a(eop_ox), .b(rst), .c(\srx/qz ) );
    nor3_1 U2 ( .x(mry), .a(eop_oy), .b(rst), .c(\sry/qz ) );
endmodule


module chain_mux0 ( eop_ix, d0_ix, d1_ix, d2_ix, d3_ix, ack_ixy, eop_iy, d0_iy, 
    d1_iy, d2_iy, d3_iy, eop_o, d0_o, d1_o, d2_o, d3_o, ack_o, rst, test_si, 
    test_se, test_so, phi1, phi2, phi3 );
input  eop_ix, d0_ix, d1_ix, d2_ix, d3_ix, eop_iy, d0_iy, d1_iy, d2_iy, d3_iy, 
    ack_o, rst, test_si, test_se, phi1, phi2, phi3;
output ack_ixy, eop_o, d0_o, d1_o, d2_o, d3_o, test_so;
    wire d3_i, d2_i, d1_i, d0_i, eop_i, n1, n2, \ce/ob , ack, \c3/ob , \c2/ob , 
        \c1/ob , \c0/ob , ack_l, \slAck/l1_q , \slAck/mxl/muxout ;
    nor2_1 U2 ( .x(d3_i), .a(d3_iy), .b(d3_ix) );
    nor2_1 U3 ( .x(d2_i), .a(d2_iy), .b(d2_ix) );
    nor2_1 U4 ( .x(d1_i), .a(d1_iy), .b(d1_ix) );
    nor2_1 U5 ( .x(d0_i), .a(d0_iy), .b(d0_ix) );
    nor2_1 U6 ( .x(eop_i), .a(eop_iy), .b(eop_ix) );
    nand2_1 U1 ( .x(ack_ixy), .a(n1), .b(n2) );
    nor3_1 U9 ( .x(n1), .a(d2_o), .b(d3_o), .c(d1_o) );
    nor2_1 U8 ( .x(n2), .a(eop_o), .b(d0_o) );
    inv_1 \ce/Ui  ( .x(\ce/ob ), .a(eop_o) );
    aoi222_1 \ce/__tmp99/U1  ( .x(eop_o), .a(eop_i), .b(ack), .c(eop_i), .d(
        \ce/ob ), .e(ack), .f(\ce/ob ) );
    inv_1 \c3/Ui  ( .x(\c3/ob ), .a(d3_o) );
    aoi222_1 \c3/__tmp99/U1  ( .x(d3_o), .a(d3_i), .b(ack), .c(d3_i), .d(
        \c3/ob ), .e(ack), .f(\c3/ob ) );
    inv_1 \c2/Ui  ( .x(\c2/ob ), .a(d2_o) );
    aoi222_1 \c2/__tmp99/U1  ( .x(d2_o), .a(d2_i), .b(ack), .c(d2_i), .d(
        \c2/ob ), .e(ack), .f(\c2/ob ) );
    inv_1 \c1/Ui  ( .x(\c1/ob ), .a(d1_o) );
    aoi222_1 \c1/__tmp99/U1  ( .x(d1_o), .a(d1_i), .b(ack), .c(d1_i), .d(
        \c1/ob ), .e(ack), .f(\c1/ob ) );
    inv_1 \c0/Ui  ( .x(\c0/ob ), .a(d0_o) );
    aoi222_1 \c0/__tmp99/U1  ( .x(d0_o), .a(d0_i), .b(ack), .c(d0_i), .d(
        \c0/ob ), .e(ack), .f(\c0/ob ) );
    latn_1 \slAck/lph3  ( .q(ack_l), .d(\slAck/l1_q ), .g(phi3) );
    latn_1 \slAck/lph2  ( .q(test_so), .d(\slAck/l1_q ), .g(phi2) );
    mux2_1 \slAck/mxl/mux  ( .x(\slAck/mxl/muxout ), .d0(ack_o), .sl(test_se), 
        .d1(test_si) );
    latn_1 \slAck/mxl/lph1  ( .q(\slAck/l1_q ), .d(\slAck/mxl/muxout ), .g(
        phi1) );
    or2_3 U7 ( .x(ack), .a(ack_l), .b(rst) );
endmodule


module chain_arbiter1 ( eop_ix, d0_ix, d1_ix, d2_ix, d3_ix, ack_ix, eop_iy, 
    d0_iy, d1_iy, d2_iy, d3_iy, ack_iy, eop_ox, d0_ox, d1_ox, d2_ox, d3_ox, 
    eop_oy, d0_oy, d1_oy, d2_oy, d3_oy, ack_oxy, rst, test_si, test_se, 
    test_so, phi1, phi2, phi3 );
input  eop_ix, d0_ix, d1_ix, d2_ix, d3_ix, eop_iy, d0_iy, d1_iy, d2_iy, d3_iy, 
    ack_oxy, rst, test_si, test_se, phi1, phi2, phi3;
output ack_ix, ack_iy, eop_ox, d0_ox, d1_ox, d2_ox, d3_ox, eop_oy, d0_oy, 
    d1_oy, d2_oy, d3_oy, test_so;
    wire nack_x, ackx_l, n1x, n2x, nack_y, acky_l, n1y, n2y, req_x, n5x, n6x, 
        req_y, n5y, n6y, sx_pl, gx, sy_pl, gy, \cye/nr , sy, \cye/nd , 
        \cye/n2 , \cy3/__tmp99/loop , \cy2/__tmp99/loop , \cy1/__tmp99/loop , 
        \cy0/__tmp99/loop , \cxe/nr , sx, \cxe/nd , \cxe/n2 , 
        \cx3/__tmp99/loop , \cx2/__tmp99/loop , \cx1/__tmp99/loop , 
        \cx0/__tmp99/loop , \mtx/gr2 , mry, \mtx/gr1 , mrx, \sry/qz , \srx/qz , 
        \sl_sy/l1_q , \scan[1] , \sl_sy/mxl/muxout , \scan[0] , \sl_sx/l1_q , 
        \sl_sx/mxl/muxout , \slAcky/l1_q , \slAcky/mxl/muxout , \scan[2] , 
        \slAckx/l1_q , \slAckx/mxl/muxout ;
    nor2_2 U12 ( .x(nack_x), .a(ackx_l), .b(rst) );
    nand2_1 U4 ( .x(ack_ix), .a(n1x), .b(n2x) );
    nor3_1 U17 ( .x(n1x), .a(d2_ox), .b(d3_ox), .c(d1_ox) );
    nor2_1 U18 ( .x(n2x), .a(eop_ox), .b(d0_ox) );
    nor2_2 U11 ( .x(nack_y), .a(acky_l), .b(rst) );
    nand2_1 U3 ( .x(ack_iy), .a(n1y), .b(n2y) );
    nor3_1 U16 ( .x(n1y), .a(d2_oy), .b(d3_oy), .c(d1_oy) );
    nor2_1 U19 ( .x(n2y), .a(eop_oy), .b(d0_oy) );
    nand2_1 U15 ( .x(req_x), .a(n5x), .b(n6x) );
    nor3_1 U10 ( .x(n5x), .a(d2_ix), .b(d3_ix), .c(d1_ix) );
    nor2_1 U13 ( .x(n6x), .a(eop_ix), .b(d0_ix) );
    nand2_1 U14 ( .x(req_y), .a(n5y), .b(n6y) );
    nor3_1 U9 ( .x(n5y), .a(d2_iy), .b(d3_iy), .c(d1_iy) );
    nor2_1 U20 ( .x(n6y), .a(eop_iy), .b(d0_iy) );
    nor2i_1 U6 ( .x(sx_pl), .a(gx), .b(eop_oy) );
    nor2i_1 U5 ( .x(sy_pl), .a(gy), .b(eop_ox) );
    nor3_1 \cye/Unr  ( .x(\cye/nr ), .a(eop_iy), .b(nack_y), .c(sy) );
    nand3_1 \cye/Und  ( .x(\cye/nd ), .a(eop_iy), .b(nack_y), .c(sy) );
    oa21_1 \cye/U1  ( .x(\cye/n2 ), .a(\cye/n2 ), .b(\cye/nr ), .c(\cye/nd )
         );
    inv_1 \cye/U3  ( .x(eop_oy), .a(\cye/n2 ) );
    ao31_1 \cy3/__tmp99/aoi  ( .x(\cy3/__tmp99/loop ), .a(d3_iy), .b(nack_y), 
        .c(sy), .d(d3_oy) );
    oa21_1 \cy3/__tmp99/outGate  ( .x(d3_oy), .a(d3_iy), .b(nack_y), .c(
        \cy3/__tmp99/loop ) );
    ao31_1 \cy2/__tmp99/aoi  ( .x(\cy2/__tmp99/loop ), .a(d2_iy), .b(nack_y), 
        .c(sy), .d(d2_oy) );
    oa21_1 \cy2/__tmp99/outGate  ( .x(d2_oy), .a(d2_iy), .b(nack_y), .c(
        \cy2/__tmp99/loop ) );
    ao31_1 \cy1/__tmp99/aoi  ( .x(\cy1/__tmp99/loop ), .a(d1_iy), .b(nack_y), 
        .c(sy), .d(d1_oy) );
    oa21_1 \cy1/__tmp99/outGate  ( .x(d1_oy), .a(d1_iy), .b(nack_y), .c(
        \cy1/__tmp99/loop ) );
    ao31_1 \cy0/__tmp99/aoi  ( .x(\cy0/__tmp99/loop ), .a(d0_iy), .b(nack_y), 
        .c(sy), .d(d0_oy) );
    oa21_1 \cy0/__tmp99/outGate  ( .x(d0_oy), .a(d0_iy), .b(nack_y), .c(
        \cy0/__tmp99/loop ) );
    nor3_1 \cxe/Unr  ( .x(\cxe/nr ), .a(eop_ix), .b(nack_x), .c(sx) );
    nand3_1 \cxe/Und  ( .x(\cxe/nd ), .a(eop_ix), .b(nack_x), .c(sx) );
    oa21_1 \cxe/U1  ( .x(\cxe/n2 ), .a(\cxe/n2 ), .b(\cxe/nr ), .c(\cxe/nd )
         );
    inv_1 \cxe/U3  ( .x(eop_ox), .a(\cxe/n2 ) );
    ao31_1 \cx3/__tmp99/aoi  ( .x(\cx3/__tmp99/loop ), .a(d3_ix), .b(nack_x), 
        .c(sx), .d(d3_ox) );
    oa21_1 \cx3/__tmp99/outGate  ( .x(d3_ox), .a(d3_ix), .b(nack_x), .c(
        \cx3/__tmp99/loop ) );
    ao31_1 \cx2/__tmp99/aoi  ( .x(\cx2/__tmp99/loop ), .a(d2_ix), .b(nack_x), 
        .c(sx), .d(d2_ox) );
    oa21_1 \cx2/__tmp99/outGate  ( .x(d2_ox), .a(d2_ix), .b(nack_x), .c(
        \cx2/__tmp99/loop ) );
    ao31_1 \cx1/__tmp99/aoi  ( .x(\cx1/__tmp99/loop ), .a(d1_ix), .b(nack_x), 
        .c(sx), .d(d1_ox) );
    oa21_1 \cx1/__tmp99/outGate  ( .x(d1_ox), .a(d1_ix), .b(nack_x), .c(
        \cx1/__tmp99/loop ) );
    ao31_1 \cx0/__tmp99/aoi  ( .x(\cx0/__tmp99/loop ), .a(d0_ix), .b(nack_x), 
        .c(sx), .d(d0_ox) );
    oa21_1 \cx0/__tmp99/outGate  ( .x(d0_ox), .a(d0_ix), .b(nack_x), .c(
        \cx0/__tmp99/loop ) );
    nand2_1 \mtx/mg2  ( .x(\mtx/gr2 ), .a(mry), .b(\mtx/gr1 ) );
    nand2_1 \mtx/U1  ( .x(\mtx/gr1 ), .a(mrx), .b(\mtx/gr2 ) );
    nor3_1 \mtx/U2  ( .x(gy), .a(\mtx/gr2 ), .b(\mtx/gr2 ), .c(\mtx/gr2 ) );
    nor3_1 \mtx/U3  ( .x(gx), .a(\mtx/gr1 ), .b(\mtx/gr1 ), .c(\mtx/gr1 ) );
    nor2_1 \sry/i1  ( .x(\sry/qz ), .a(req_y), .b(mry) );
    nor2_1 \srx/i1  ( .x(\srx/qz ), .a(req_x), .b(mrx) );
    latn_1 \sl_sy/lph3  ( .q(sy), .d(\sl_sy/l1_q ), .g(phi3) );
    latn_1 \sl_sy/lph2  ( .q(\scan[1] ), .d(\sl_sy/l1_q ), .g(phi2) );
    mux2_1 \sl_sy/mxl/mux  ( .x(\sl_sy/mxl/muxout ), .d0(sy_pl), .sl(test_se), 
        .d1(\scan[0] ) );
    latn_1 \sl_sy/mxl/lph1  ( .q(\sl_sy/l1_q ), .d(\sl_sy/mxl/muxout ), .g(
        phi1) );
    latn_1 \sl_sx/lph3  ( .q(sx), .d(\sl_sx/l1_q ), .g(phi3) );
    latn_1 \sl_sx/lph2  ( .q(\scan[0] ), .d(\sl_sx/l1_q ), .g(phi2) );
    mux2_1 \sl_sx/mxl/mux  ( .x(\sl_sx/mxl/muxout ), .d0(sx_pl), .sl(test_se), 
        .d1(test_si) );
    latn_1 \sl_sx/mxl/lph1  ( .q(\sl_sx/l1_q ), .d(\sl_sx/mxl/muxout ), .g(
        phi1) );
    latn_1 \slAcky/lph3  ( .q(acky_l), .d(\slAcky/l1_q ), .g(phi3) );
    latn_1 \slAcky/lph2  ( .q(test_so), .d(\slAcky/l1_q ), .g(phi2) );
    mux2_1 \slAcky/mxl/mux  ( .x(\slAcky/mxl/muxout ), .d0(ack_oxy), .sl(
        test_se), .d1(\scan[2] ) );
    latn_1 \slAcky/mxl/lph1  ( .q(\slAcky/l1_q ), .d(\slAcky/mxl/muxout ), .g(
        phi1) );
    latn_1 \slAckx/lph3  ( .q(ackx_l), .d(\slAckx/l1_q ), .g(phi3) );
    latn_1 \slAckx/lph2  ( .q(\scan[2] ), .d(\slAckx/l1_q ), .g(phi2) );
    mux2_1 \slAckx/mxl/mux  ( .x(\slAckx/mxl/muxout ), .d0(ack_oxy), .sl(
        test_se), .d1(\scan[1] ) );
    latn_1 \slAckx/mxl/lph1  ( .q(\slAckx/l1_q ), .d(\slAckx/mxl/muxout ), .g(
        phi1) );
    nor3_1 U1 ( .x(mrx), .a(eop_ox), .b(rst), .c(\srx/qz ) );
    nor3_1 U2 ( .x(mry), .a(eop_oy), .b(rst), .c(\sry/qz ) );
endmodule


module chain_mux1 ( eop_ix, d0_ix, d1_ix, d2_ix, d3_ix, ack_ixy, eop_iy, d0_iy, 
    d1_iy, d2_iy, d3_iy, eop_o, d0_o, d1_o, d2_o, d3_o, ack_o, rst, test_si, 
    test_se, test_so, phi1, phi2, phi3 );
input  eop_ix, d0_ix, d1_ix, d2_ix, d3_ix, eop_iy, d0_iy, d1_iy, d2_iy, d3_iy, 
    ack_o, rst, test_si, test_se, phi1, phi2, phi3;
output ack_ixy, eop_o, d0_o, d1_o, d2_o, d3_o, test_so;
    wire d3_i, d2_i, d1_i, d0_i, eop_i, n1, n2, \ce/ob , ack, \c3/ob , \c2/ob , 
        \c1/ob , \c0/ob , ack_l, \slAck/l1_q , \slAck/mxl/muxout ;
    nor2_1 U2 ( .x(d3_i), .a(d3_iy), .b(d3_ix) );
    nor2_1 U3 ( .x(d2_i), .a(d2_iy), .b(d2_ix) );
    nor2_1 U4 ( .x(d1_i), .a(d1_iy), .b(d1_ix) );
    nor2_1 U5 ( .x(d0_i), .a(d0_iy), .b(d0_ix) );
    nor2_1 U6 ( .x(eop_i), .a(eop_iy), .b(eop_ix) );
    nand2_1 U1 ( .x(ack_ixy), .a(n1), .b(n2) );
    nor3_1 U9 ( .x(n1), .a(d2_o), .b(d3_o), .c(d1_o) );
    nor2_1 U8 ( .x(n2), .a(eop_o), .b(d0_o) );
    inv_1 \ce/Ui  ( .x(\ce/ob ), .a(eop_o) );
    aoi222_1 \ce/__tmp99/U1  ( .x(eop_o), .a(eop_i), .b(ack), .c(eop_i), .d(
        \ce/ob ), .e(ack), .f(\ce/ob ) );
    inv_1 \c3/Ui  ( .x(\c3/ob ), .a(d3_o) );
    aoi222_1 \c3/__tmp99/U1  ( .x(d3_o), .a(d3_i), .b(ack), .c(d3_i), .d(
        \c3/ob ), .e(ack), .f(\c3/ob ) );
    inv_1 \c2/Ui  ( .x(\c2/ob ), .a(d2_o) );
    aoi222_1 \c2/__tmp99/U1  ( .x(d2_o), .a(d2_i), .b(ack), .c(d2_i), .d(
        \c2/ob ), .e(ack), .f(\c2/ob ) );
    inv_1 \c1/Ui  ( .x(\c1/ob ), .a(d1_o) );
    aoi222_1 \c1/__tmp99/U1  ( .x(d1_o), .a(d1_i), .b(ack), .c(d1_i), .d(
        \c1/ob ), .e(ack), .f(\c1/ob ) );
    inv_1 \c0/Ui  ( .x(\c0/ob ), .a(d0_o) );
    aoi222_1 \c0/__tmp99/U1  ( .x(d0_o), .a(d0_i), .b(ack), .c(d0_i), .d(
        \c0/ob ), .e(ack), .f(\c0/ob ) );
    latn_1 \slAck/lph3  ( .q(ack_l), .d(\slAck/l1_q ), .g(phi3) );
    latn_1 \slAck/lph2  ( .q(test_so), .d(\slAck/l1_q ), .g(phi2) );
    mux2_1 \slAck/mxl/mux  ( .x(\slAck/mxl/muxout ), .d0(ack_o), .sl(test_se), 
        .d1(test_si) );
    latn_1 \slAck/mxl/lph1  ( .q(\slAck/l1_q ), .d(\slAck/mxl/muxout ), .g(
        phi1) );
    or2_3 U7 ( .x(ack), .a(ack_l), .b(rst) );
endmodule


module chain_router0 ( eop_i, d0_i, d1_i, d2_i, d3_i, ack_i, eop_ox, d0_ox, 
    d1_ox, d2_ox, d3_ox, ack_ox, eop_oy, d0_oy, d1_oy, d2_oy, d3_oy, ack_oy, 
    nrst, test_si, test_se, test_so, phi1, phi2, phi3 );
input  eop_i, d0_i, d1_i, d2_i, d3_i, ack_ox, ack_oy, nrst, test_si, test_se, 
    phi1, phi2, phi3;
output ack_i, eop_ox, d0_ox, d1_ox, d2_ox, d3_ox, eop_oy, d0_oy, d1_oy, d2_oy, 
    d3_oy, test_so;
    wire rst, nack_x, ackx_l, nack_y, acky_l, n10, n11, n12, neopxy, n1, n2, 
        n3, n4, n5, n6, n7, n8, nrouteAckx, nrouteAcky, nroutex, nroutey, qa, 
        nqx, nqy, sx_pl, qx, sy_pl, qy, routeAcky, \cy/__tmp99/nr , qa_l, 
        \cy/__tmp99/nd , routeAckx, \cx/__tmp99/nr , \cx/__tmp99/nd , \cye/nr , 
        sy, \cye/nd , \cye/n2 , \cy3/__tmp99/loop , \cy2/__tmp99/loop , 
        \cy1/__tmp99/loop , \cy0/__tmp99/loop , \cxe/nr , sx, \cxe/nd , 
        \cxe/n2 , \cx3/__tmp99/loop , \cx2/__tmp99/loop , \cx1/__tmp99/loop , 
        \cx0/__tmp99/loop , \sl_sy/l1_q , \scan[2] , \sl_sy/mxl/muxout , 
        \scan[1] , \sl_sx/l1_q , \sl_sx/mxl/muxout , \scan[0] , \sl_qa/l1_q , 
        \sl_qa/mxl/muxout , \slAcky/l1_q , \slAcky/mxl/muxout , \scan[3] , 
        \slAckx/l1_q , \slAckx/mxl/muxout ;
    inv_1 U0 ( .x(rst), .a(nrst) );
    nor2_2 U5 ( .x(nack_x), .a(ackx_l), .b(rst) );
    nor2_2 U4 ( .x(nack_y), .a(acky_l), .b(rst) );
    nand4_1 U1 ( .x(ack_i), .a(n10), .b(n11), .c(n12), .d(neopxy) );
    and4_1 U8 ( .x(n10), .a(n1), .b(n2), .c(n3), .d(n4) );
    inv_1 U10 ( .x(n1), .a(d0_oy) );
    inv_1 U11 ( .x(n2), .a(d1_oy) );
    inv_1 U14 ( .x(n3), .a(d2_oy) );
    inv_1 U16 ( .x(n4), .a(d3_oy) );
    and4_1 U9 ( .x(n11), .a(n5), .b(n6), .c(n7), .d(n8) );
    inv_1 U17 ( .x(n5), .a(d0_ox) );
    inv_1 U18 ( .x(n6), .a(d1_ox) );
    inv_1 U19 ( .x(n7), .a(d2_ox) );
    inv_1 U20 ( .x(n8), .a(d3_ox) );
    nor2_1 U7 ( .x(n12), .a(nrouteAckx), .b(nrouteAcky) );
    nor2_1 U6 ( .x(neopxy), .a(eop_oy), .b(eop_ox) );
    nor2_1 U3 ( .x(nroutex), .a(d3_i), .b(d1_i) );
    nor2_1 U2 ( .x(nroutey), .a(d2_i), .b(d0_i) );
    nand2_1 U12 ( .x(qa), .a(nqx), .b(nqy) );
    nor2i_1 U15 ( .x(sx_pl), .a(qx), .b(nrouteAckx) );
    nor2i_1 U13 ( .x(sy_pl), .a(qy), .b(nrouteAcky) );
    inv_1 \cy/U1  ( .x(nrouteAcky), .a(routeAcky) );
    nor2_1 \cy/__tmp99/U1  ( .x(\cy/__tmp99/nr ), .a(nroutey), .b(qa_l) );
    nand2_1 \cy/__tmp99/U2  ( .x(\cy/__tmp99/nd ), .a(nroutey), .b(qa_l) );
    oai211_1 \cy/__tmp99/U3  ( .x(routeAcky), .a(nrouteAcky), .b(
        \cy/__tmp99/nr ), .c(\cy/__tmp99/nd ), .d(nrst) );
    inv_1 \cx/U1  ( .x(nrouteAckx), .a(routeAckx) );
    nor2_1 \cx/__tmp99/U1  ( .x(\cx/__tmp99/nr ), .a(nroutex), .b(qa_l) );
    nand2_1 \cx/__tmp99/U2  ( .x(\cx/__tmp99/nd ), .a(nroutex), .b(qa_l) );
    oai211_1 \cx/__tmp99/U3  ( .x(routeAckx), .a(nrouteAckx), .b(
        \cx/__tmp99/nr ), .c(\cx/__tmp99/nd ), .d(nrst) );
    nor3_1 \cye/Unr  ( .x(\cye/nr ), .a(eop_i), .b(nack_y), .c(sy) );
    nand3_1 \cye/Und  ( .x(\cye/nd ), .a(eop_i), .b(nack_y), .c(sy) );
    oa21_1 \cye/U1  ( .x(\cye/n2 ), .a(\cye/n2 ), .b(\cye/nr ), .c(\cye/nd )
         );
    inv_1 \cye/U3  ( .x(eop_oy), .a(\cye/n2 ) );
    ao31_1 \cy3/__tmp99/aoi  ( .x(\cy3/__tmp99/loop ), .a(d3_i), .b(nack_y), 
        .c(sy), .d(d3_oy) );
    ao31_1 \cy2/__tmp99/aoi  ( .x(\cy2/__tmp99/loop ), .a(d2_i), .b(nack_y), 
        .c(sy), .d(d2_oy) );
    ao31_1 \cy1/__tmp99/aoi  ( .x(\cy1/__tmp99/loop ), .a(d1_i), .b(nack_y), 
        .c(sy), .d(d1_oy) );
    ao31_1 \cy0/__tmp99/aoi  ( .x(\cy0/__tmp99/loop ), .a(d0_i), .b(nack_y), 
        .c(sy), .d(d0_oy) );
    nor3_1 \cxe/Unr  ( .x(\cxe/nr ), .a(eop_i), .b(nack_x), .c(sx) );
    nand3_1 \cxe/Und  ( .x(\cxe/nd ), .a(eop_i), .b(nack_x), .c(sx) );
    oa21_1 \cxe/U1  ( .x(\cxe/n2 ), .a(\cxe/n2 ), .b(\cxe/nr ), .c(\cxe/nd )
         );
    inv_1 \cxe/U3  ( .x(eop_ox), .a(\cxe/n2 ) );
    ao31_1 \cx3/__tmp99/aoi  ( .x(\cx3/__tmp99/loop ), .a(d3_i), .b(nack_x), 
        .c(sx), .d(d3_ox) );
    oa21_1 \cx3/__tmp99/outGate  ( .x(d3_ox), .a(d3_i), .b(nack_x), .c(
        \cx3/__tmp99/loop ) );
    ao31_1 \cx2/__tmp99/aoi  ( .x(\cx2/__tmp99/loop ), .a(d2_i), .b(nack_x), 
        .c(sx), .d(d2_ox) );
    oa21_1 \cx2/__tmp99/outGate  ( .x(d2_ox), .a(d2_i), .b(nack_x), .c(
        \cx2/__tmp99/loop ) );
    ao31_1 \cx1/__tmp99/aoi  ( .x(\cx1/__tmp99/loop ), .a(d1_i), .b(nack_x), 
        .c(sx), .d(d1_ox) );
    oa21_1 \cx1/__tmp99/outGate  ( .x(d1_ox), .a(d1_i), .b(nack_x), .c(
        \cx1/__tmp99/loop ) );
    ao31_1 \cx0/__tmp99/aoi  ( .x(\cx0/__tmp99/loop ), .a(d0_i), .b(nack_x), 
        .c(sx), .d(d0_ox) );
    oa21_1 \cx0/__tmp99/outGate  ( .x(d0_ox), .a(d0_i), .b(nack_x), .c(
        \cx0/__tmp99/loop ) );
    nand3_1 \sry/i0  ( .x(nqy), .a(neopxy), .b(nrst), .c(qy) );
    nand2_1 \sry/i1  ( .x(qy), .a(routeAcky), .b(nqy) );
    nand3_1 \srx/i0  ( .x(nqx), .a(neopxy), .b(nrst), .c(qx) );
    nand2_1 \srx/i1  ( .x(qx), .a(routeAckx), .b(nqx) );
    latn_1 \sl_sy/lph3  ( .q(sy), .d(\sl_sy/l1_q ), .g(phi3) );
    latn_1 \sl_sy/lph2  ( .q(\scan[2] ), .d(\sl_sy/l1_q ), .g(phi2) );
    mux2_1 \sl_sy/mxl/mux  ( .x(\sl_sy/mxl/muxout ), .d0(sy_pl), .sl(test_se), 
        .d1(\scan[1] ) );
    latn_1 \sl_sy/mxl/lph1  ( .q(\sl_sy/l1_q ), .d(\sl_sy/mxl/muxout ), .g(
        phi1) );
    latn_1 \sl_sx/lph3  ( .q(sx), .d(\sl_sx/l1_q ), .g(phi3) );
    latn_1 \sl_sx/lph2  ( .q(\scan[1] ), .d(\sl_sx/l1_q ), .g(phi2) );
    mux2_1 \sl_sx/mxl/mux  ( .x(\sl_sx/mxl/muxout ), .d0(sx_pl), .sl(test_se), 
        .d1(\scan[0] ) );
    latn_1 \sl_sx/mxl/lph1  ( .q(\sl_sx/l1_q ), .d(\sl_sx/mxl/muxout ), .g(
        phi1) );
    latn_1 \sl_qa/lph3  ( .q(qa_l), .d(\sl_qa/l1_q ), .g(phi3) );
    latn_1 \sl_qa/lph2  ( .q(\scan[0] ), .d(\sl_qa/l1_q ), .g(phi2) );
    mux2_1 \sl_qa/mxl/mux  ( .x(\sl_qa/mxl/muxout ), .d0(qa), .sl(test_se), 
        .d1(test_si) );
    latn_1 \sl_qa/mxl/lph1  ( .q(\sl_qa/l1_q ), .d(\sl_qa/mxl/muxout ), .g(
        phi1) );
    latn_1 \slAcky/lph3  ( .q(acky_l), .d(\slAcky/l1_q ), .g(phi3) );
    latn_1 \slAcky/lph2  ( .q(test_so), .d(\slAcky/l1_q ), .g(phi2) );
    mux2_1 \slAcky/mxl/mux  ( .x(\slAcky/mxl/muxout ), .d0(ack_oy), .sl(
        test_se), .d1(\scan[3] ) );
    latn_1 \slAcky/mxl/lph1  ( .q(\slAcky/l1_q ), .d(\slAcky/mxl/muxout ), .g(
        phi1) );
    latn_1 \slAckx/lph3  ( .q(ackx_l), .d(\slAckx/l1_q ), .g(phi3) );
    latn_1 \slAckx/lph2  ( .q(\scan[3] ), .d(\slAckx/l1_q ), .g(phi2) );
    mux2_1 \slAckx/mxl/mux  ( .x(\slAckx/mxl/muxout ), .d0(ack_ox), .sl(
        test_se), .d1(\scan[2] ) );
    latn_1 \slAckx/mxl/lph1  ( .q(\slAckx/l1_q ), .d(\slAckx/mxl/muxout ), .g(
        phi1) );
    oa21_2 U21 ( .x(d2_oy), .a(d2_i), .b(nack_y), .c(\cy2/__tmp99/loop ) );
    oa21_2 U22 ( .x(d1_oy), .a(d1_i), .b(nack_y), .c(\cy1/__tmp99/loop ) );
    oa21_2 U23 ( .x(d3_oy), .a(d3_i), .b(nack_y), .c(\cy3/__tmp99/loop ) );
    oa21_2 U24 ( .x(d0_oy), .a(d0_i), .b(nack_y), .c(\cy0/__tmp99/loop ) );
endmodule


module chain_router1 ( eop_i, d0_i, d1_i, d2_i, d3_i, ack_i, eop_ox, d0_ox, 
    d1_ox, d2_ox, d3_ox, ack_ox, eop_oy, d0_oy, d1_oy, d2_oy, d3_oy, ack_oy, 
    nrst, test_si, test_se, test_so, phi1, phi2, phi3 );
input  eop_i, d0_i, d1_i, d2_i, d3_i, ack_ox, ack_oy, nrst, test_si, test_se, 
    phi1, phi2, phi3;
output ack_i, eop_ox, d0_ox, d1_ox, d2_ox, d3_ox, eop_oy, d0_oy, d1_oy, d2_oy, 
    d3_oy, test_so;
    wire rst, nack_x, ackx_l, nack_y, acky_l, n10, n11, n12, neopxy, n1, n2, 
        n3, n4, n5, n6, n7, n8, nrouteAckx, nrouteAcky, nroutex, nroutey, qa, 
        nqx, nqy, sx_pl, qx, sy_pl, qy, routeAcky, \cy/__tmp99/nr , qa_l, 
        \cy/__tmp99/nd , routeAckx, \cx/__tmp99/nr , \cx/__tmp99/nd , \cye/nr , 
        sy, \cye/nd , \cye/n2 , \cy3/__tmp99/loop , \cy2/__tmp99/loop , 
        \cy1/__tmp99/loop , \cy0/__tmp99/loop , \cxe/nr , sx, \cxe/nd , 
        \cxe/n2 , \cx3/__tmp99/loop , \cx2/__tmp99/loop , \cx1/__tmp99/loop , 
        \cx0/__tmp99/loop , \sl_sy/l1_q , \scan[2] , \sl_sy/mxl/muxout , 
        \scan[1] , \sl_sx/l1_q , \sl_sx/mxl/muxout , \scan[0] , \sl_qa/l1_q , 
        \sl_qa/mxl/muxout , \slAcky/l1_q , \slAcky/mxl/muxout , \scan[3] , 
        \slAckx/l1_q , \slAckx/mxl/muxout ;
    inv_1 U0 ( .x(rst), .a(nrst) );
    nor2_2 U5 ( .x(nack_x), .a(ackx_l), .b(rst) );
    nor2_2 U4 ( .x(nack_y), .a(acky_l), .b(rst) );
    nand4_1 U1 ( .x(ack_i), .a(n10), .b(n11), .c(n12), .d(neopxy) );
    and4_1 U8 ( .x(n10), .a(n1), .b(n2), .c(n3), .d(n4) );
    inv_1 U10 ( .x(n1), .a(d0_oy) );
    inv_1 U11 ( .x(n2), .a(d1_oy) );
    inv_1 U14 ( .x(n3), .a(d2_oy) );
    inv_1 U16 ( .x(n4), .a(d3_oy) );
    and4_1 U9 ( .x(n11), .a(n5), .b(n6), .c(n7), .d(n8) );
    inv_1 U17 ( .x(n5), .a(d0_ox) );
    inv_1 U18 ( .x(n6), .a(d1_ox) );
    inv_1 U19 ( .x(n7), .a(d2_ox) );
    inv_1 U20 ( .x(n8), .a(d3_ox) );
    nor2_1 U7 ( .x(n12), .a(nrouteAckx), .b(nrouteAcky) );
    nor2_1 U6 ( .x(neopxy), .a(eop_oy), .b(eop_ox) );
    nor2_1 U3 ( .x(nroutex), .a(d3_i), .b(d1_i) );
    nor2_1 U2 ( .x(nroutey), .a(d2_i), .b(d0_i) );
    nand2_1 U12 ( .x(qa), .a(nqx), .b(nqy) );
    nor2i_1 U15 ( .x(sx_pl), .a(qx), .b(nrouteAckx) );
    nor2i_1 U13 ( .x(sy_pl), .a(qy), .b(nrouteAcky) );
    inv_1 \cy/U1  ( .x(nrouteAcky), .a(routeAcky) );
    nor2_1 \cy/__tmp99/U1  ( .x(\cy/__tmp99/nr ), .a(nroutey), .b(qa_l) );
    nand2_1 \cy/__tmp99/U2  ( .x(\cy/__tmp99/nd ), .a(nroutey), .b(qa_l) );
    oai211_1 \cy/__tmp99/U3  ( .x(routeAcky), .a(nrouteAcky), .b(
        \cy/__tmp99/nr ), .c(\cy/__tmp99/nd ), .d(nrst) );
    inv_1 \cx/U1  ( .x(nrouteAckx), .a(routeAckx) );
    nor2_1 \cx/__tmp99/U1  ( .x(\cx/__tmp99/nr ), .a(nroutex), .b(qa_l) );
    nand2_1 \cx/__tmp99/U2  ( .x(\cx/__tmp99/nd ), .a(nroutex), .b(qa_l) );
    oai211_1 \cx/__tmp99/U3  ( .x(routeAckx), .a(nrouteAckx), .b(
        \cx/__tmp99/nr ), .c(\cx/__tmp99/nd ), .d(nrst) );
    nor3_1 \cye/Unr  ( .x(\cye/nr ), .a(eop_i), .b(nack_y), .c(sy) );
    nand3_1 \cye/Und  ( .x(\cye/nd ), .a(eop_i), .b(nack_y), .c(sy) );
    oa21_1 \cye/U1  ( .x(\cye/n2 ), .a(\cye/n2 ), .b(\cye/nr ), .c(\cye/nd )
         );
    inv_1 \cye/U3  ( .x(eop_oy), .a(\cye/n2 ) );
    ao31_1 \cy3/__tmp99/aoi  ( .x(\cy3/__tmp99/loop ), .a(d3_i), .b(nack_y), 
        .c(sy), .d(d3_oy) );
    oa21_1 \cy3/__tmp99/outGate  ( .x(d3_oy), .a(d3_i), .b(nack_y), .c(
        \cy3/__tmp99/loop ) );
    ao31_1 \cy2/__tmp99/aoi  ( .x(\cy2/__tmp99/loop ), .a(d2_i), .b(nack_y), 
        .c(sy), .d(d2_oy) );
    oa21_1 \cy2/__tmp99/outGate  ( .x(d2_oy), .a(d2_i), .b(nack_y), .c(
        \cy2/__tmp99/loop ) );
    ao31_1 \cy1/__tmp99/aoi  ( .x(\cy1/__tmp99/loop ), .a(d1_i), .b(nack_y), 
        .c(sy), .d(d1_oy) );
    oa21_1 \cy1/__tmp99/outGate  ( .x(d1_oy), .a(d1_i), .b(nack_y), .c(
        \cy1/__tmp99/loop ) );
    ao31_1 \cy0/__tmp99/aoi  ( .x(\cy0/__tmp99/loop ), .a(d0_i), .b(nack_y), 
        .c(sy), .d(d0_oy) );
    oa21_1 \cy0/__tmp99/outGate  ( .x(d0_oy), .a(d0_i), .b(nack_y), .c(
        \cy0/__tmp99/loop ) );
    nor3_1 \cxe/Unr  ( .x(\cxe/nr ), .a(eop_i), .b(nack_x), .c(sx) );
    nand3_1 \cxe/Und  ( .x(\cxe/nd ), .a(eop_i), .b(nack_x), .c(sx) );
    oa21_1 \cxe/U1  ( .x(\cxe/n2 ), .a(\cxe/n2 ), .b(\cxe/nr ), .c(\cxe/nd )
         );
    inv_1 \cxe/U3  ( .x(eop_ox), .a(\cxe/n2 ) );
    ao31_1 \cx3/__tmp99/aoi  ( .x(\cx3/__tmp99/loop ), .a(d3_i), .b(nack_x), 
        .c(sx), .d(d3_ox) );
    oa21_1 \cx3/__tmp99/outGate  ( .x(d3_ox), .a(d3_i), .b(nack_x), .c(
        \cx3/__tmp99/loop ) );
    ao31_1 \cx2/__tmp99/aoi  ( .x(\cx2/__tmp99/loop ), .a(d2_i), .b(nack_x), 
        .c(sx), .d(d2_ox) );
    oa21_1 \cx2/__tmp99/outGate  ( .x(d2_ox), .a(d2_i), .b(nack_x), .c(
        \cx2/__tmp99/loop ) );
    ao31_1 \cx1/__tmp99/aoi  ( .x(\cx1/__tmp99/loop ), .a(d1_i), .b(nack_x), 
        .c(sx), .d(d1_ox) );
    oa21_1 \cx1/__tmp99/outGate  ( .x(d1_ox), .a(d1_i), .b(nack_x), .c(
        \cx1/__tmp99/loop ) );
    ao31_1 \cx0/__tmp99/aoi  ( .x(\cx0/__tmp99/loop ), .a(d0_i), .b(nack_x), 
        .c(sx), .d(d0_ox) );
    oa21_1 \cx0/__tmp99/outGate  ( .x(d0_ox), .a(d0_i), .b(nack_x), .c(
        \cx0/__tmp99/loop ) );
    nand3_1 \sry/i0  ( .x(nqy), .a(neopxy), .b(nrst), .c(qy) );
    nand2_1 \sry/i1  ( .x(qy), .a(routeAcky), .b(nqy) );
    nand3_1 \srx/i0  ( .x(nqx), .a(neopxy), .b(nrst), .c(qx) );
    nand2_1 \srx/i1  ( .x(qx), .a(routeAckx), .b(nqx) );
    latn_1 \sl_sy/lph3  ( .q(sy), .d(\sl_sy/l1_q ), .g(phi3) );
    latn_1 \sl_sy/lph2  ( .q(\scan[2] ), .d(\sl_sy/l1_q ), .g(phi2) );
    mux2_1 \sl_sy/mxl/mux  ( .x(\sl_sy/mxl/muxout ), .d0(sy_pl), .sl(test_se), 
        .d1(\scan[1] ) );
    latn_1 \sl_sy/mxl/lph1  ( .q(\sl_sy/l1_q ), .d(\sl_sy/mxl/muxout ), .g(
        phi1) );
    latn_1 \sl_sx/lph3  ( .q(sx), .d(\sl_sx/l1_q ), .g(phi3) );
    latn_1 \sl_sx/lph2  ( .q(\scan[1] ), .d(\sl_sx/l1_q ), .g(phi2) );
    mux2_1 \sl_sx/mxl/mux  ( .x(\sl_sx/mxl/muxout ), .d0(sx_pl), .sl(test_se), 
        .d1(\scan[0] ) );
    latn_1 \sl_sx/mxl/lph1  ( .q(\sl_sx/l1_q ), .d(\sl_sx/mxl/muxout ), .g(
        phi1) );
    latn_1 \sl_qa/lph3  ( .q(qa_l), .d(\sl_qa/l1_q ), .g(phi3) );
    latn_1 \sl_qa/lph2  ( .q(\scan[0] ), .d(\sl_qa/l1_q ), .g(phi2) );
    mux2_1 \sl_qa/mxl/mux  ( .x(\sl_qa/mxl/muxout ), .d0(qa), .sl(test_se), 
        .d1(test_si) );
    latn_1 \sl_qa/mxl/lph1  ( .q(\sl_qa/l1_q ), .d(\sl_qa/mxl/muxout ), .g(
        phi1) );
    latn_1 \slAcky/lph3  ( .q(acky_l), .d(\slAcky/l1_q ), .g(phi3) );
    latn_1 \slAcky/lph2  ( .q(test_so), .d(\slAcky/l1_q ), .g(phi2) );
    mux2_1 \slAcky/mxl/mux  ( .x(\slAcky/mxl/muxout ), .d0(ack_oy), .sl(
        test_se), .d1(\scan[3] ) );
    latn_1 \slAcky/mxl/lph1  ( .q(\slAcky/l1_q ), .d(\slAcky/mxl/muxout ), .g(
        phi1) );
    latn_1 \slAckx/lph3  ( .q(ackx_l), .d(\slAckx/l1_q ), .g(phi3) );
    latn_1 \slAckx/lph2  ( .q(\scan[3] ), .d(\slAckx/l1_q ), .g(phi2) );
    mux2_1 \slAckx/mxl/mux  ( .x(\slAckx/mxl/muxout ), .d0(ack_ox), .sl(
        test_se), .d1(\scan[2] ) );
    latn_1 \slAckx/mxl/lph1  ( .q(\slAckx/l1_q ), .d(\slAckx/mxl/muxout ), .g(
        phi1) );
endmodule


module chain_router2 ( eop_i, d0_i, d1_i, d2_i, d3_i, ack_i, eop_ox, d0_ox, 
    d1_ox, d2_ox, d3_ox, ack_ox, eop_oy, d0_oy, d1_oy, d2_oy, d3_oy, ack_oy, 
    nrst, test_si, test_se, test_so, phi1, phi2, phi3 );
input  eop_i, d0_i, d1_i, d2_i, d3_i, ack_ox, ack_oy, nrst, test_si, test_se, 
    phi1, phi2, phi3;
output ack_i, eop_ox, d0_ox, d1_ox, d2_ox, d3_ox, eop_oy, d0_oy, d1_oy, d2_oy, 
    d3_oy, test_so;
    wire rst, nack_x, ackx_l, nack_y, acky_l, n10, n11, n12, neopxy, n1, n2, 
        n3, n4, n5, n6, n7, n8, nrouteAckx, nrouteAcky, nroutex, nroutey, qa, 
        nqx, nqy, sx_pl, qx, sy_pl, qy, routeAcky, \cy/__tmp99/nr , qa_l, 
        \cy/__tmp99/nd , routeAckx, \cx/__tmp99/nr , \cx/__tmp99/nd , \cye/nr , 
        sy, \cye/nd , \cye/n2 , \cy3/__tmp99/loop , \cy2/__tmp99/loop , 
        \cy1/__tmp99/loop , \cy0/__tmp99/loop , \cxe/nr , sx, \cxe/nd , 
        \cxe/n2 , \cx3/__tmp99/loop , \cx2/__tmp99/loop , \cx1/__tmp99/loop , 
        \cx0/__tmp99/loop , \sl_sy/l1_q , \scan[2] , \sl_sy/mxl/muxout , 
        \scan[1] , \sl_sx/l1_q , \sl_sx/mxl/muxout , \scan[0] , \sl_qa/l1_q , 
        \sl_qa/mxl/muxout , \slAcky/l1_q , \slAcky/mxl/muxout , \scan[3] , 
        \slAckx/l1_q , \slAckx/mxl/muxout ;
    inv_1 U0 ( .x(rst), .a(nrst) );
    nor2_2 U5 ( .x(nack_x), .a(ackx_l), .b(rst) );
    nor2_2 U4 ( .x(nack_y), .a(acky_l), .b(rst) );
    nand4_1 U1 ( .x(ack_i), .a(n10), .b(n11), .c(n12), .d(neopxy) );
    and4_1 U8 ( .x(n10), .a(n1), .b(n2), .c(n3), .d(n4) );
    inv_1 U10 ( .x(n1), .a(d0_oy) );
    inv_1 U11 ( .x(n2), .a(d1_oy) );
    inv_1 U14 ( .x(n3), .a(d2_oy) );
    inv_1 U16 ( .x(n4), .a(d3_oy) );
    and4_1 U9 ( .x(n11), .a(n5), .b(n6), .c(n7), .d(n8) );
    inv_1 U17 ( .x(n5), .a(d0_ox) );
    inv_1 U18 ( .x(n6), .a(d1_ox) );
    inv_1 U19 ( .x(n7), .a(d2_ox) );
    inv_1 U20 ( .x(n8), .a(d3_ox) );
    nor2_1 U7 ( .x(n12), .a(nrouteAckx), .b(nrouteAcky) );
    nor2_1 U6 ( .x(neopxy), .a(eop_oy), .b(eop_ox) );
    nor2_1 U3 ( .x(nroutex), .a(d3_i), .b(d1_i) );
    nor2_1 U2 ( .x(nroutey), .a(d2_i), .b(d0_i) );
    nand2_1 U12 ( .x(qa), .a(nqx), .b(nqy) );
    nor2i_1 U15 ( .x(sx_pl), .a(qx), .b(nrouteAckx) );
    nor2i_1 U13 ( .x(sy_pl), .a(qy), .b(nrouteAcky) );
    inv_1 \cy/U1  ( .x(nrouteAcky), .a(routeAcky) );
    nor2_1 \cy/__tmp99/U1  ( .x(\cy/__tmp99/nr ), .a(nroutey), .b(qa_l) );
    nand2_1 \cy/__tmp99/U2  ( .x(\cy/__tmp99/nd ), .a(nroutey), .b(qa_l) );
    oai211_1 \cy/__tmp99/U3  ( .x(routeAcky), .a(nrouteAcky), .b(
        \cy/__tmp99/nr ), .c(\cy/__tmp99/nd ), .d(nrst) );
    inv_1 \cx/U1  ( .x(nrouteAckx), .a(routeAckx) );
    nor2_1 \cx/__tmp99/U1  ( .x(\cx/__tmp99/nr ), .a(nroutex), .b(qa_l) );
    nand2_1 \cx/__tmp99/U2  ( .x(\cx/__tmp99/nd ), .a(nroutex), .b(qa_l) );
    oai211_1 \cx/__tmp99/U3  ( .x(routeAckx), .a(nrouteAckx), .b(
        \cx/__tmp99/nr ), .c(\cx/__tmp99/nd ), .d(nrst) );
    nor3_1 \cye/Unr  ( .x(\cye/nr ), .a(eop_i), .b(nack_y), .c(sy) );
    nand3_1 \cye/Und  ( .x(\cye/nd ), .a(eop_i), .b(nack_y), .c(sy) );
    oa21_1 \cye/U1  ( .x(\cye/n2 ), .a(\cye/n2 ), .b(\cye/nr ), .c(\cye/nd )
         );
    inv_1 \cye/U3  ( .x(eop_oy), .a(\cye/n2 ) );
    ao31_1 \cy3/__tmp99/aoi  ( .x(\cy3/__tmp99/loop ), .a(d3_i), .b(nack_y), 
        .c(sy), .d(d3_oy) );
    ao31_1 \cy2/__tmp99/aoi  ( .x(\cy2/__tmp99/loop ), .a(d2_i), .b(nack_y), 
        .c(sy), .d(d2_oy) );
    ao31_1 \cy1/__tmp99/aoi  ( .x(\cy1/__tmp99/loop ), .a(d1_i), .b(nack_y), 
        .c(sy), .d(d1_oy) );
    ao31_1 \cy0/__tmp99/aoi  ( .x(\cy0/__tmp99/loop ), .a(d0_i), .b(nack_y), 
        .c(sy), .d(d0_oy) );
    nor3_1 \cxe/Unr  ( .x(\cxe/nr ), .a(eop_i), .b(nack_x), .c(sx) );
    nand3_1 \cxe/Und  ( .x(\cxe/nd ), .a(eop_i), .b(nack_x), .c(sx) );
    oa21_1 \cxe/U1  ( .x(\cxe/n2 ), .a(\cxe/n2 ), .b(\cxe/nr ), .c(\cxe/nd )
         );
    inv_1 \cxe/U3  ( .x(eop_ox), .a(\cxe/n2 ) );
    ao31_1 \cx3/__tmp99/aoi  ( .x(\cx3/__tmp99/loop ), .a(d3_i), .b(nack_x), 
        .c(sx), .d(d3_ox) );
    ao31_1 \cx2/__tmp99/aoi  ( .x(\cx2/__tmp99/loop ), .a(d2_i), .b(nack_x), 
        .c(sx), .d(d2_ox) );
    ao31_1 \cx1/__tmp99/aoi  ( .x(\cx1/__tmp99/loop ), .a(d1_i), .b(nack_x), 
        .c(sx), .d(d1_ox) );
    ao31_1 \cx0/__tmp99/aoi  ( .x(\cx0/__tmp99/loop ), .a(d0_i), .b(nack_x), 
        .c(sx), .d(d0_ox) );
    nand3_1 \sry/i0  ( .x(nqy), .a(neopxy), .b(nrst), .c(qy) );
    nand2_1 \sry/i1  ( .x(qy), .a(routeAcky), .b(nqy) );
    nand3_1 \srx/i0  ( .x(nqx), .a(neopxy), .b(nrst), .c(qx) );
    nand2_1 \srx/i1  ( .x(qx), .a(routeAckx), .b(nqx) );
    latn_1 \sl_sy/lph3  ( .q(sy), .d(\sl_sy/l1_q ), .g(phi3) );
    latn_1 \sl_sy/lph2  ( .q(\scan[2] ), .d(\sl_sy/l1_q ), .g(phi2) );
    mux2_1 \sl_sy/mxl/mux  ( .x(\sl_sy/mxl/muxout ), .d0(sy_pl), .sl(test_se), 
        .d1(\scan[1] ) );
    latn_1 \sl_sy/mxl/lph1  ( .q(\sl_sy/l1_q ), .d(\sl_sy/mxl/muxout ), .g(
        phi1) );
    latn_1 \sl_sx/lph3  ( .q(sx), .d(\sl_sx/l1_q ), .g(phi3) );
    latn_1 \sl_sx/lph2  ( .q(\scan[1] ), .d(\sl_sx/l1_q ), .g(phi2) );
    mux2_1 \sl_sx/mxl/mux  ( .x(\sl_sx/mxl/muxout ), .d0(sx_pl), .sl(test_se), 
        .d1(\scan[0] ) );
    latn_1 \sl_sx/mxl/lph1  ( .q(\sl_sx/l1_q ), .d(\sl_sx/mxl/muxout ), .g(
        phi1) );
    latn_1 \sl_qa/lph3  ( .q(qa_l), .d(\sl_qa/l1_q ), .g(phi3) );
    latn_1 \sl_qa/lph2  ( .q(\scan[0] ), .d(\sl_qa/l1_q ), .g(phi2) );
    mux2_1 \sl_qa/mxl/mux  ( .x(\sl_qa/mxl/muxout ), .d0(qa), .sl(test_se), 
        .d1(test_si) );
    latn_1 \sl_qa/mxl/lph1  ( .q(\sl_qa/l1_q ), .d(\sl_qa/mxl/muxout ), .g(
        phi1) );
    latn_1 \slAcky/lph3  ( .q(acky_l), .d(\slAcky/l1_q ), .g(phi3) );
    latn_1 \slAcky/lph2  ( .q(test_so), .d(\slAcky/l1_q ), .g(phi2) );
    mux2_1 \slAcky/mxl/mux  ( .x(\slAcky/mxl/muxout ), .d0(ack_oy), .sl(
        test_se), .d1(\scan[3] ) );
    latn_1 \slAcky/mxl/lph1  ( .q(\slAcky/l1_q ), .d(\slAcky/mxl/muxout ), .g(
        phi1) );
    latn_1 \slAckx/lph3  ( .q(ackx_l), .d(\slAckx/l1_q ), .g(phi3) );
    latn_1 \slAckx/lph2  ( .q(\scan[3] ), .d(\slAckx/l1_q ), .g(phi2) );
    mux2_1 \slAckx/mxl/mux  ( .x(\slAckx/mxl/muxout ), .d0(ack_ox), .sl(
        test_se), .d1(\scan[2] ) );
    latn_1 \slAckx/mxl/lph1  ( .q(\slAckx/l1_q ), .d(\slAckx/mxl/muxout ), .g(
        phi1) );
    oa21_2 U21 ( .x(d3_oy), .a(d3_i), .b(nack_y), .c(\cy3/__tmp99/loop ) );
    oa21_2 U22 ( .x(d2_oy), .a(d2_i), .b(nack_y), .c(\cy2/__tmp99/loop ) );
    oa21_2 U23 ( .x(d1_ox), .a(d1_i), .b(nack_x), .c(\cx1/__tmp99/loop ) );
    oa21_2 U24 ( .x(d3_ox), .a(d3_i), .b(nack_x), .c(\cx3/__tmp99/loop ) );
    oa21_2 U25 ( .x(d2_ox), .a(d2_i), .b(nack_x), .c(\cx2/__tmp99/loop ) );
    oa21_2 U26 ( .x(d0_oy), .a(d0_i), .b(nack_y), .c(\cy0/__tmp99/loop ) );
    oa21_2 U27 ( .x(d0_ox), .a(d0_i), .b(nack_x), .c(\cx0/__tmp99/loop ) );
    oa21_2 U28 ( .x(d1_oy), .a(d1_i), .b(nack_y), .c(\cy1/__tmp99/loop ) );
endmodule


module comm_fab ( nrst, I_port_eop_i, I_port_d0_i, I_port_d1_i, I_port_d2_i, 
    I_port_d3_i, I_port_ack, TIC_eop_i, TIC_d0_i, TIC_d1_i, TIC_d2_i, TIC_d3_i, 
    TIC_ack, D_port_eop_i, D_port_d0_i, D_port_d1_i, D_port_d2_i, D_port_d3_i, 
    D_port_ack, BC_eop_i, BC_d0_i, BC_d1_i, BC_d2_i, BC_d3_i, BC_ack, WB_eop_i, 
    WB_d0_i, WB_d1_i, WB_d2_i, WB_d3_i, WB_ack, IMEM_eop_i, IMEM_d0_i, 
    IMEM_d1_i, IMEM_d2_i, IMEM_d3_i, IMEM_ack, DMEM_eop_i, DMEM_d0_i, 
    DMEM_d1_i, DMEM_d2_i, DMEM_d3_i, DMEM_ack, test_si, test_so, test_se, phi1, 
    phi2, phi3 );
input  nrst, I_port_eop_i, I_port_d0_i, I_port_d1_i, I_port_d2_i, I_port_d3_i, 
    TIC_eop_i, TIC_d0_i, TIC_d1_i, TIC_d2_i, TIC_d3_i, D_port_eop_i, 
    D_port_d0_i, D_port_d1_i, D_port_d2_i, D_port_d3_i, BC_ack, WB_ack, 
    IMEM_ack, DMEM_ack, test_si, test_se, phi1, phi2, phi3;
output I_port_ack, TIC_ack, D_port_ack, BC_eop_i, BC_d0_i, BC_d1_i, BC_d2_i, 
    BC_d3_i, WB_eop_i, WB_d0_i, WB_d1_i, WB_d2_i, WB_d3_i, IMEM_eop_i, 
    IMEM_d0_i, IMEM_d1_i, IMEM_d2_i, IMEM_d3_i, DMEM_eop_i, DMEM_d0_i, 
    DMEM_d1_i, DMEM_d2_i, DMEM_d3_i, test_so;
    wire rst, A0_eop_o0, A0_d0_o0, A0_d1_o0, A0_d2_o0, A0_d3_o0, A0_eop_o1, 
        A0_d0_o1, A0_d1_o1, A0_d2_o1, A0_d3_o1, A0_ack, n4, \scan[1] , M0_eop, 
        M0_d0, M0_d1, M0_d2, M0_d3, M0_ack, \scan[2] , n2, n1, n3, A1_eop_o0, 
        A1_d0_o0, A1_d1_o0, A1_d2_o0, A1_d3_o0, A1_eop_o1, A1_d0_o1, A1_d1_o1, 
        A1_d2_o1, A1_d3_o1, A1_ack, \scan[3] , M1_eop, M1_d0, M1_d1, M1_d2, 
        M1_d3, M1_ack, \scan[4] , R0_odd_eop, R0_odd_d0, R0_odd_d1, R0_odd_d2, 
        R0_odd_d3, R0_odd_ack, \scan[5] , R1_odd_eop, R1_odd_d0, R1_odd_d1, 
        R1_odd_d2, R1_odd_d3, R1_odd_ack, \scan[6] ;
    inv_2 U1 ( .x(rst), .a(nrst) );
    chain_arbiter0 arb0 ( .eop_ix(I_port_eop_i), .d0_ix(I_port_d0_i), .d1_ix(
        I_port_d1_i), .d2_ix(I_port_d2_i), .d3_ix(I_port_d3_i), .ack_ix(
        I_port_ack), .eop_iy(D_port_eop_i), .d0_iy(D_port_d0_i), .d1_iy(
        D_port_d1_i), .d2_iy(D_port_d2_i), .d3_iy(D_port_d3_i), .ack_iy(
        D_port_ack), .eop_ox(A0_eop_o0), .d0_ox(A0_d0_o0), .d1_ox(A0_d1_o0), 
        .d2_ox(A0_d2_o0), .d3_ox(A0_d3_o0), .eop_oy(A0_eop_o1), .d0_oy(
        A0_d0_o1), .d1_oy(A0_d1_o1), .d2_oy(A0_d2_o1), .d3_oy(A0_d3_o1), 
        .ack_oxy(A0_ack), .rst(rst), .test_si(test_si), .test_se(n4), 
        .test_so(\scan[1] ), .phi1(phi1), .phi2(phi2), .phi3(phi3) );
    chain_mux0 mux0 ( .eop_ix(A0_eop_o0), .d0_ix(A0_d0_o0), .d1_ix(A0_d1_o0), 
        .d2_ix(A0_d2_o0), .d3_ix(A0_d3_o0), .ack_ixy(A0_ack), .eop_iy(
        A0_eop_o1), .d0_iy(A0_d0_o1), .d1_iy(A0_d1_o1), .d2_iy(A0_d2_o1), 
        .d3_iy(A0_d3_o1), .eop_o(M0_eop), .d0_o(M0_d0), .d1_o(M0_d1), .d2_o(
        M0_d2), .d3_o(M0_d3), .ack_o(M0_ack), .rst(rst), .test_si(\scan[1] ), 
        .test_se(n4), .test_so(\scan[2] ), .phi1(n2), .phi2(n1), .phi3(n3) );
    chain_arbiter1 arb1 ( .eop_ix(M0_eop), .d0_ix(M0_d0), .d1_ix(M0_d1), 
        .d2_ix(M0_d2), .d3_ix(M0_d3), .ack_ix(M0_ack), .eop_iy(TIC_eop_i), 
        .d0_iy(TIC_d0_i), .d1_iy(TIC_d1_i), .d2_iy(TIC_d2_i), .d3_iy(TIC_d3_i), 
        .ack_iy(TIC_ack), .eop_ox(A1_eop_o0), .d0_ox(A1_d0_o0), .d1_ox(
        A1_d1_o0), .d2_ox(A1_d2_o0), .d3_ox(A1_d3_o0), .eop_oy(A1_eop_o1), 
        .d0_oy(A1_d0_o1), .d1_oy(A1_d1_o1), .d2_oy(A1_d2_o1), .d3_oy(A1_d3_o1), 
        .ack_oxy(A1_ack), .rst(rst), .test_si(\scan[2] ), .test_se(n4), 
        .test_so(\scan[3] ), .phi1(n2), .phi2(n1), .phi3(n3) );
    chain_mux1 mux1 ( .eop_ix(A1_eop_o0), .d0_ix(A1_d0_o0), .d1_ix(A1_d1_o0), 
        .d2_ix(A1_d2_o0), .d3_ix(A1_d3_o0), .ack_ixy(A1_ack), .eop_iy(
        A1_eop_o1), .d0_iy(A1_d0_o1), .d1_iy(A1_d1_o1), .d2_iy(A1_d2_o1), 
        .d3_iy(A1_d3_o1), .eop_o(M1_eop), .d0_o(M1_d0), .d1_o(M1_d1), .d2_o(
        M1_d2), .d3_o(M1_d3), .ack_o(M1_ack), .rst(rst), .test_si(\scan[3] ), 
        .test_se(test_se), .test_so(\scan[4] ), .phi1(phi1), .phi2(phi2), 
        .phi3(phi3) );
    chain_router0 router0 ( .eop_i(M1_eop), .d0_i(M1_d0), .d1_i(M1_d1), .d2_i(
        M1_d2), .d3_i(M1_d3), .ack_i(M1_ack), .eop_ox(R0_odd_eop), .d0_ox(
        R0_odd_d0), .d1_ox(R0_odd_d1), .d2_ox(R0_odd_d2), .d3_ox(R0_odd_d3), 
        .ack_ox(R0_odd_ack), .eop_oy(WB_eop_i), .d0_oy(WB_d0_i), .d1_oy(
        WB_d1_i), .d2_oy(WB_d2_i), .d3_oy(WB_d3_i), .ack_oy(WB_ack), .nrst(
        nrst), .test_si(\scan[4] ), .test_se(test_se), .test_so(\scan[5] ), 
        .phi1(phi1), .phi2(phi2), .phi3(phi3) );
    chain_router1 router1 ( .eop_i(R0_odd_eop), .d0_i(R0_odd_d0), .d1_i(
        R0_odd_d1), .d2_i(R0_odd_d2), .d3_i(R0_odd_d3), .ack_i(R0_odd_ack), 
        .eop_ox(R1_odd_eop), .d0_ox(R1_odd_d0), .d1_ox(R1_odd_d1), .d2_ox(
        R1_odd_d2), .d3_ox(R1_odd_d3), .ack_ox(R1_odd_ack), .eop_oy(BC_eop_i), 
        .d0_oy(BC_d0_i), .d1_oy(BC_d1_i), .d2_oy(BC_d2_i), .d3_oy(BC_d3_i), 
        .ack_oy(BC_ack), .nrst(nrst), .test_si(\scan[5] ), .test_se(n4), 
        .test_so(\scan[6] ), .phi1(n2), .phi2(n1), .phi3(n3) );
    chain_router2 router2 ( .eop_i(R1_odd_eop), .d0_i(R1_odd_d0), .d1_i(
        R1_odd_d1), .d2_i(R1_odd_d2), .d3_i(R1_odd_d3), .ack_i(R1_odd_ack), 
        .eop_ox(DMEM_eop_i), .d0_ox(DMEM_d0_i), .d1_ox(DMEM_d1_i), .d2_ox(
        DMEM_d2_i), .d3_ox(DMEM_d3_i), .ack_ox(DMEM_ack), .eop_oy(IMEM_eop_i), 
        .d0_oy(IMEM_d0_i), .d1_oy(IMEM_d1_i), .d2_oy(IMEM_d2_i), .d3_oy(
        IMEM_d3_i), .ack_oy(IMEM_ack), .nrst(nrst), .test_si(\scan[6] ), 
        .test_se(test_se), .test_so(test_so), .phi1(phi1), .phi2(phi2), .phi3(
        phi3) );
    buf_1 U2 ( .x(n1), .a(phi2) );
    buf_1 U3 ( .x(n2), .a(phi1) );
    buf_1 U4 ( .x(n3), .a(phi3) );
    buf_3 U5 ( .x(n4), .a(test_se) );
endmodule


module comm_fab_scan ( nrst, I_port_eop_i, I_port_d0_i, I_port_d1_i, 
    I_port_d2_i, I_port_d3_i, I_port_ack, TIC_eop_i, TIC_d0_i, TIC_d1_i, 
    TIC_d2_i, TIC_d3_i, TIC_ack, D_port_eop_i, D_port_d0_i, D_port_d1_i, 
    D_port_d2_i, D_port_d3_i, D_port_ack, BC_eop_i, BC_d0_i, BC_d1_i, BC_d2_i, 
    BC_d3_i, BC_ack, WB_eop_i, WB_d0_i, WB_d1_i, WB_d2_i, WB_d3_i, WB_ack, 
    IMEM_eop_i, IMEM_d0_i, IMEM_d1_i, IMEM_d2_i, IMEM_d3_i, IMEM_ack, 
    DMEM_eop_i, DMEM_d0_i, DMEM_d1_i, DMEM_d2_i, DMEM_d3_i, DMEM_ack, test_si, 
    test_so, test_se, phi1, phi2, phi3 );
input  nrst, I_port_eop_i, I_port_d0_i, I_port_d1_i, I_port_d2_i, I_port_d3_i, 
    TIC_eop_i, TIC_d0_i, TIC_d1_i, TIC_d2_i, TIC_d3_i, D_port_eop_i, 
    D_port_d0_i, D_port_d1_i, D_port_d2_i, D_port_d3_i, BC_ack, WB_ack, 
    IMEM_ack, DMEM_ack, test_si, test_se, phi1, phi2, phi3;
output I_port_ack, TIC_ack, D_port_ack, BC_eop_i, BC_d0_i, BC_d1_i, BC_d2_i, 
    BC_d3_i, WB_eop_i, WB_d0_i, WB_d1_i, WB_d2_i, WB_d3_i, IMEM_eop_i, 
    IMEM_d0_i, IMEM_d1_i, IMEM_d2_i, IMEM_d3_i, DMEM_eop_i, DMEM_d0_i, 
    DMEM_d1_i, DMEM_d2_i, DMEM_d3_i, test_so;
    wire I_port_eop_i_sc, I_port_d0_i_sc, I_port_d1_i_sc, I_port_d2_i_sc, 
        I_port_d3_i_sc, TIC_eop_i_sc, TIC_d0_i_sc, TIC_d1_i_sc, TIC_d2_i_sc, 
        TIC_d3_i_sc, D_port_eop_i_sc, D_port_d0_i_sc, D_port_d1_i_sc, 
        D_port_d2_i_sc, D_port_d3_i_sc, WB_ack_sc, IMEM_ack_sc, DMEM_ack_sc, 
        \scan[6] , \scan[7] , n13, n9, n5, n2, \scan[11] , scan_m10, n7, 
        \scan[12] , scan_m11, n4, scan_m12, n6, \sc12_m_dpAck/muxout , n15, 
        n11, \sc11_m_ticAck/muxout , n14, n8, \sc10_m_ipAck/muxout , 
        \scan[10] , n10, \sc5_dmAck/l1_q , n1, \sc5_dmAck/mxl/muxout , 
        \scan[5] , \sc4_imAck/l1_q , \sc4_imAck/mxl/muxout , n12, \scan[4] , 
        \sc3_wbAck/l1_q , \sc3_wbAck/mxl/muxout , \scan[3] , \sc_dm/intI4 , 
        \sc_dm/scn3 , \sc_dm/intI3 , \sc_dm/scn2 , \sc_dm/intI2 , \sc_dm/scn1 , 
        \sc_dm/intI1 , \sc_dm/scn0 , \sc_dm/intI0 , \sc_dm/l4_m/muxout , 
        \sc_dm/l3_m/muxout , \sc_dm/l2_m/muxout , \sc_dm/l1_m/muxout , 
        \sc_dm/l0_m/muxout , \scan[9] , \sc_im/intI4 , \sc_im/scn3 , 
        \sc_im/intI3 , \sc_im/scn2 , \sc_im/intI2 , \sc_im/scn1 , 
        \sc_im/intI1 , \sc_im/scn0 , \sc_im/intI0 , \sc_im/l4_m/muxout , 
        \sc_im/l3_m/muxout , \sc_im/l2_m/muxout , \sc_im/l1_m/muxout , 
        \sc_im/l0_m/muxout , \scan[8] , \sc_wb/intI4 , \sc_wb/scn3 , 
        \sc_wb/intI3 , \sc_wb/scn2 , \sc_wb/intI2 , \sc_wb/scn1 , 
        \sc_wb/intI1 , \sc_wb/scn0 , \sc_wb/intI0 , \sc_wb/l4_m/muxout , 
        \sc_wb/l3_m/muxout , \sc_wb/l2_m/muxout , \sc_wb/l1_m/muxout , 
        \sc_wb/l0_m/muxout , \sc_dp/sl4/l1_q , n3, \sc_dp/sl4/mxl/muxout , 
        \sc_dp/scn4 , \sc_dp/sl3/l1_q , \sc_dp/sl3/mxl/muxout , \sc_dp/scn3 , 
        \sc_dp/sl2/l1_q , \sc_dp/sl2/mxl/muxout , \sc_dp/scn2 , 
        \sc_dp/sl1/l1_q , \sc_dp/sl1/mxl/muxout , \sc_dp/scn1 , 
        \sc_dp/sl0/l1_q , \sc_dp/sl0/mxl/muxout , \scan[2] , \sc_tic/sl4/l1_q , 
        \sc_tic/sl4/mxl/muxout , \sc_tic/scn4 , \sc_tic/sl3/l1_q , 
        \sc_tic/sl3/mxl/muxout , \sc_tic/scn3 , \sc_tic/sl2/l1_q , 
        \sc_tic/sl2/mxl/muxout , \sc_tic/scn2 , \sc_tic/sl1/l1_q , 
        \sc_tic/sl1/mxl/muxout , \sc_tic/scn1 , \sc_tic/sl0/l1_q , 
        \sc_tic/sl0/mxl/muxout , \scan[1] , \sc_ip/sl4/l1_q , 
        \sc_ip/sl4/mxl/muxout , \sc_ip/scn4 , \sc_ip/sl3/l1_q , 
        \sc_ip/sl3/mxl/muxout , \sc_ip/scn3 , \sc_ip/sl2/l1_q , 
        \sc_ip/sl2/mxl/muxout , \sc_ip/scn2 , \sc_ip/sl1/l1_q , 
        \sc_ip/sl1/mxl/muxout , \sc_ip/scn1 , \sc_ip/sl0/l1_q , 
        \sc_ip/sl0/mxl/muxout ;
    comm_fab fab1 ( .nrst(nrst), .I_port_eop_i(I_port_eop_i_sc), .I_port_d0_i(
        I_port_d0_i_sc), .I_port_d1_i(I_port_d1_i_sc), .I_port_d2_i(
        I_port_d2_i_sc), .I_port_d3_i(I_port_d3_i_sc), .I_port_ack(I_port_ack), 
        .TIC_eop_i(TIC_eop_i_sc), .TIC_d0_i(TIC_d0_i_sc), .TIC_d1_i(
        TIC_d1_i_sc), .TIC_d2_i(TIC_d2_i_sc), .TIC_d3_i(TIC_d3_i_sc), 
        .TIC_ack(TIC_ack), .D_port_eop_i(D_port_eop_i_sc), .D_port_d0_i(
        D_port_d0_i_sc), .D_port_d1_i(D_port_d1_i_sc), .D_port_d2_i(
        D_port_d2_i_sc), .D_port_d3_i(D_port_d3_i_sc), .D_port_ack(D_port_ack), 
        .BC_eop_i(BC_eop_i), .BC_d0_i(BC_d0_i), .BC_d1_i(BC_d1_i), .BC_d2_i(
        BC_d2_i), .BC_d3_i(BC_d3_i), .BC_ack(BC_ack), .WB_eop_i(WB_eop_i), 
        .WB_d0_i(WB_d0_i), .WB_d1_i(WB_d1_i), .WB_d2_i(WB_d2_i), .WB_d3_i(
        WB_d3_i), .WB_ack(WB_ack_sc), .IMEM_eop_i(IMEM_eop_i), .IMEM_d0_i(
        IMEM_d0_i), .IMEM_d1_i(IMEM_d1_i), .IMEM_d2_i(IMEM_d2_i), .IMEM_d3_i(
        IMEM_d3_i), .IMEM_ack(IMEM_ack_sc), .DMEM_eop_i(DMEM_eop_i), 
        .DMEM_d0_i(DMEM_d0_i), .DMEM_d1_i(DMEM_d1_i), .DMEM_d2_i(DMEM_d2_i), 
        .DMEM_d3_i(DMEM_d3_i), .DMEM_ack(DMEM_ack_sc), .test_si(\scan[6] ), 
        .test_so(\scan[7] ), .test_se(n13), .phi1(n9), .phi2(n5), .phi3(n2) );
    latn_1 sc10_s_ipAck ( .q(\scan[11] ), .d(scan_m10), .g(n7) );
    latn_1 sc11_s_ticAck ( .q(\scan[12] ), .d(scan_m11), .g(n4) );
    latn_1 sc12_s_dpAck ( .q(test_so), .d(scan_m12), .g(n6) );
    mux2_1 \sc12_m_dpAck/mux  ( .x(\sc12_m_dpAck/muxout ), .d0(D_port_ack), 
        .sl(n15), .d1(\scan[12] ) );
    latn_1 \sc12_m_dpAck/lph1  ( .q(scan_m12), .d(\sc12_m_dpAck/muxout ), .g(
        n11) );
    mux2_1 \sc11_m_ticAck/mux  ( .x(\sc11_m_ticAck/muxout ), .d0(TIC_ack), 
        .sl(n14), .d1(\scan[11] ) );
    latn_1 \sc11_m_ticAck/lph1  ( .q(scan_m11), .d(\sc11_m_ticAck/muxout ), 
        .g(n8) );
    mux2_1 \sc10_m_ipAck/mux  ( .x(\sc10_m_ipAck/muxout ), .d0(I_port_ack), 
        .sl(n14), .d1(\scan[10] ) );
    latn_1 \sc10_m_ipAck/lph1  ( .q(scan_m10), .d(\sc10_m_ipAck/muxout ), .g(
        n10) );
    latn_1 \sc5_dmAck/lph3  ( .q(DMEM_ack_sc), .d(\sc5_dmAck/l1_q ), .g(n1) );
    latn_1 \sc5_dmAck/lph2  ( .q(\scan[6] ), .d(\sc5_dmAck/l1_q ), .g(n7) );
    mux2_1 \sc5_dmAck/mxl/mux  ( .x(\sc5_dmAck/mxl/muxout ), .d0(DMEM_ack), 
        .sl(n15), .d1(\scan[5] ) );
    latn_1 \sc5_dmAck/mxl/lph1  ( .q(\sc5_dmAck/l1_q ), .d(
        \sc5_dmAck/mxl/muxout ), .g(n10) );
    latn_1 \sc4_imAck/lph3  ( .q(IMEM_ack_sc), .d(\sc4_imAck/l1_q ), .g(n1) );
    latn_1 \sc4_imAck/lph2  ( .q(\scan[5] ), .d(\sc4_imAck/l1_q ), .g(n4) );
    mux2_1 \sc4_imAck/mxl/mux  ( .x(\sc4_imAck/mxl/muxout ), .d0(IMEM_ack), 
        .sl(n12), .d1(\scan[4] ) );
    latn_1 \sc4_imAck/mxl/lph1  ( .q(\sc4_imAck/l1_q ), .d(
        \sc4_imAck/mxl/muxout ), .g(n8) );
    latn_1 \sc3_wbAck/lph3  ( .q(WB_ack_sc), .d(\sc3_wbAck/l1_q ), .g(n1) );
    latn_1 \sc3_wbAck/lph2  ( .q(\scan[4] ), .d(\sc3_wbAck/l1_q ), .g(n6) );
    mux2_1 \sc3_wbAck/mxl/mux  ( .x(\sc3_wbAck/mxl/muxout ), .d0(WB_ack), .sl(
        n12), .d1(\scan[3] ) );
    latn_1 \sc3_wbAck/mxl/lph1  ( .q(\sc3_wbAck/l1_q ), .d(
        \sc3_wbAck/mxl/muxout ), .g(n11) );
    latn_1 \sc_dm/l4_s  ( .q(\scan[10] ), .d(\sc_dm/intI4 ), .g(n7) );
    latn_1 \sc_dm/l3_s  ( .q(\sc_dm/scn3 ), .d(\sc_dm/intI3 ), .g(n4) );
    latn_1 \sc_dm/l2_s  ( .q(\sc_dm/scn2 ), .d(\sc_dm/intI2 ), .g(n6) );
    latn_1 \sc_dm/l1_s  ( .q(\sc_dm/scn1 ), .d(\sc_dm/intI1 ), .g(n7) );
    latn_1 \sc_dm/l0_s  ( .q(\sc_dm/scn0 ), .d(\sc_dm/intI0 ), .g(n4) );
    mux2_1 \sc_dm/l4_m/mux  ( .x(\sc_dm/l4_m/muxout ), .d0(DMEM_d3_i), .sl(n12
        ), .d1(\sc_dm/scn3 ) );
    latn_1 \sc_dm/l4_m/lph1  ( .q(\sc_dm/intI4 ), .d(\sc_dm/l4_m/muxout ), .g(
        n8) );
    mux2_1 \sc_dm/l3_m/mux  ( .x(\sc_dm/l3_m/muxout ), .d0(DMEM_d2_i), .sl(n15
        ), .d1(\sc_dm/scn2 ) );
    latn_1 \sc_dm/l3_m/lph1  ( .q(\sc_dm/intI3 ), .d(\sc_dm/l3_m/muxout ), .g(
        n11) );
    mux2_1 \sc_dm/l2_m/mux  ( .x(\sc_dm/l2_m/muxout ), .d0(DMEM_d1_i), .sl(n14
        ), .d1(\sc_dm/scn1 ) );
    latn_1 \sc_dm/l2_m/lph1  ( .q(\sc_dm/intI2 ), .d(\sc_dm/l2_m/muxout ), .g(
        n10) );
    mux2_1 \sc_dm/l1_m/mux  ( .x(\sc_dm/l1_m/muxout ), .d0(DMEM_d0_i), .sl(n12
        ), .d1(\sc_dm/scn0 ) );
    latn_1 \sc_dm/l1_m/lph1  ( .q(\sc_dm/intI1 ), .d(\sc_dm/l1_m/muxout ), .g(
        n8) );
    mux2_1 \sc_dm/l0_m/mux  ( .x(\sc_dm/l0_m/muxout ), .d0(DMEM_eop_i), .sl(
        n15), .d1(\scan[9] ) );
    latn_1 \sc_dm/l0_m/lph1  ( .q(\sc_dm/intI0 ), .d(\sc_dm/l0_m/muxout ), .g(
        n11) );
    latn_1 \sc_im/l4_s  ( .q(\scan[9] ), .d(\sc_im/intI4 ), .g(n4) );
    latn_1 \sc_im/l3_s  ( .q(\sc_im/scn3 ), .d(\sc_im/intI3 ), .g(n6) );
    latn_1 \sc_im/l2_s  ( .q(\sc_im/scn2 ), .d(\sc_im/intI2 ), .g(n7) );
    latn_1 \sc_im/l1_s  ( .q(\sc_im/scn1 ), .d(\sc_im/intI1 ), .g(n4) );
    latn_1 \sc_im/l0_s  ( .q(\sc_im/scn0 ), .d(\sc_im/intI0 ), .g(n6) );
    mux2_1 \sc_im/l4_m/mux  ( .x(\sc_im/l4_m/muxout ), .d0(IMEM_d3_i), .sl(n14
        ), .d1(\sc_im/scn3 ) );
    latn_1 \sc_im/l4_m/lph1  ( .q(\sc_im/intI4 ), .d(\sc_im/l4_m/muxout ), .g(
        n10) );
    mux2_1 \sc_im/l3_m/mux  ( .x(\sc_im/l3_m/muxout ), .d0(IMEM_d2_i), .sl(n12
        ), .d1(\sc_im/scn2 ) );
    latn_1 \sc_im/l3_m/lph1  ( .q(\sc_im/intI3 ), .d(\sc_im/l3_m/muxout ), .g(
        n8) );
    mux2_1 \sc_im/l2_m/mux  ( .x(\sc_im/l2_m/muxout ), .d0(IMEM_d1_i), .sl(n15
        ), .d1(\sc_im/scn1 ) );
    latn_1 \sc_im/l2_m/lph1  ( .q(\sc_im/intI2 ), .d(\sc_im/l2_m/muxout ), .g(
        n11) );
    mux2_1 \sc_im/l1_m/mux  ( .x(\sc_im/l1_m/muxout ), .d0(IMEM_d0_i), .sl(n14
        ), .d1(\sc_im/scn0 ) );
    latn_1 \sc_im/l1_m/lph1  ( .q(\sc_im/intI1 ), .d(\sc_im/l1_m/muxout ), .g(
        n10) );
    mux2_1 \sc_im/l0_m/mux  ( .x(\sc_im/l0_m/muxout ), .d0(IMEM_eop_i), .sl(
        n12), .d1(\scan[8] ) );
    latn_1 \sc_im/l0_m/lph1  ( .q(\sc_im/intI0 ), .d(\sc_im/l0_m/muxout ), .g(
        n8) );
    latn_1 \sc_wb/l4_s  ( .q(\scan[8] ), .d(\sc_wb/intI4 ), .g(n6) );
    latn_1 \sc_wb/l3_s  ( .q(\sc_wb/scn3 ), .d(\sc_wb/intI3 ), .g(n7) );
    latn_1 \sc_wb/l2_s  ( .q(\sc_wb/scn2 ), .d(\sc_wb/intI2 ), .g(n4) );
    latn_1 \sc_wb/l1_s  ( .q(\sc_wb/scn1 ), .d(\sc_wb/intI1 ), .g(n6) );
    latn_1 \sc_wb/l0_s  ( .q(\sc_wb/scn0 ), .d(\sc_wb/intI0 ), .g(n7) );
    mux2_1 \sc_wb/l4_m/mux  ( .x(\sc_wb/l4_m/muxout ), .d0(WB_d3_i), .sl(n15), 
        .d1(\sc_wb/scn3 ) );
    latn_1 \sc_wb/l4_m/lph1  ( .q(\sc_wb/intI4 ), .d(\sc_wb/l4_m/muxout ), .g(
        n11) );
    mux2_1 \sc_wb/l3_m/mux  ( .x(\sc_wb/l3_m/muxout ), .d0(WB_d2_i), .sl(n15), 
        .d1(\sc_wb/scn2 ) );
    latn_1 \sc_wb/l3_m/lph1  ( .q(\sc_wb/intI3 ), .d(\sc_wb/l3_m/muxout ), .g(
        n10) );
    mux2_1 \sc_wb/l2_m/mux  ( .x(\sc_wb/l2_m/muxout ), .d0(WB_d1_i), .sl(n14), 
        .d1(\sc_wb/scn1 ) );
    latn_1 \sc_wb/l2_m/lph1  ( .q(\sc_wb/intI2 ), .d(\sc_wb/l2_m/muxout ), .g(
        n8) );
    mux2_1 \sc_wb/l1_m/mux  ( .x(\sc_wb/l1_m/muxout ), .d0(WB_d0_i), .sl(n12), 
        .d1(\sc_wb/scn0 ) );
    latn_1 \sc_wb/l1_m/lph1  ( .q(\sc_wb/intI1 ), .d(\sc_wb/l1_m/muxout ), .g(
        n11) );
    mux2_1 \sc_wb/l0_m/mux  ( .x(\sc_wb/l0_m/muxout ), .d0(WB_eop_i), .sl(n15), 
        .d1(\scan[7] ) );
    latn_1 \sc_wb/l0_m/lph1  ( .q(\sc_wb/intI0 ), .d(\sc_wb/l0_m/muxout ), .g(
        n10) );
    latn_1 \sc_dp/sl4/lph3  ( .q(D_port_d3_i_sc), .d(\sc_dp/sl4/l1_q ), .g(n3)
         );
    latn_1 \sc_dp/sl4/lph2  ( .q(\scan[3] ), .d(\sc_dp/sl4/l1_q ), .g(n4) );
    mux2_1 \sc_dp/sl4/mxl/mux  ( .x(\sc_dp/sl4/mxl/muxout ), .d0(D_port_d3_i), 
        .sl(n14), .d1(\sc_dp/scn4 ) );
    latn_1 \sc_dp/sl4/mxl/lph1  ( .q(\sc_dp/sl4/l1_q ), .d(
        \sc_dp/sl4/mxl/muxout ), .g(n8) );
    latn_1 \sc_dp/sl3/lph3  ( .q(D_port_d2_i_sc), .d(\sc_dp/sl3/l1_q ), .g(n3)
         );
    latn_1 \sc_dp/sl3/lph2  ( .q(\sc_dp/scn4 ), .d(\sc_dp/sl3/l1_q ), .g(n7)
         );
    mux2_1 \sc_dp/sl3/mxl/mux  ( .x(\sc_dp/sl3/mxl/muxout ), .d0(D_port_d2_i), 
        .sl(n12), .d1(\sc_dp/scn3 ) );
    latn_1 \sc_dp/sl3/mxl/lph1  ( .q(\sc_dp/sl3/l1_q ), .d(
        \sc_dp/sl3/mxl/muxout ), .g(n11) );
    latn_1 \sc_dp/sl2/lph3  ( .q(D_port_d1_i_sc), .d(\sc_dp/sl2/l1_q ), .g(n3)
         );
    latn_1 \sc_dp/sl2/lph2  ( .q(\sc_dp/scn3 ), .d(\sc_dp/sl2/l1_q ), .g(n6)
         );
    mux2_1 \sc_dp/sl2/mxl/mux  ( .x(\sc_dp/sl2/mxl/muxout ), .d0(D_port_d1_i), 
        .sl(n15), .d1(\sc_dp/scn2 ) );
    latn_1 \sc_dp/sl2/mxl/lph1  ( .q(\sc_dp/sl2/l1_q ), .d(
        \sc_dp/sl2/mxl/muxout ), .g(n10) );
    latn_1 \sc_dp/sl1/lph3  ( .q(D_port_d0_i_sc), .d(\sc_dp/sl1/l1_q ), .g(n3)
         );
    latn_1 \sc_dp/sl1/lph2  ( .q(\sc_dp/scn2 ), .d(\sc_dp/sl1/l1_q ), .g(n7)
         );
    mux2_1 \sc_dp/sl1/mxl/mux  ( .x(\sc_dp/sl1/mxl/muxout ), .d0(D_port_d0_i), 
        .sl(n12), .d1(\sc_dp/scn1 ) );
    latn_1 \sc_dp/sl1/mxl/lph1  ( .q(\sc_dp/sl1/l1_q ), .d(
        \sc_dp/sl1/mxl/muxout ), .g(n11) );
    latn_1 \sc_dp/sl0/lph3  ( .q(D_port_eop_i_sc), .d(\sc_dp/sl0/l1_q ), .g(n3
        ) );
    latn_1 \sc_dp/sl0/lph2  ( .q(\sc_dp/scn1 ), .d(\sc_dp/sl0/l1_q ), .g(n4)
         );
    mux2_1 \sc_dp/sl0/mxl/mux  ( .x(\sc_dp/sl0/mxl/muxout ), .d0(D_port_eop_i), 
        .sl(n12), .d1(\scan[2] ) );
    latn_1 \sc_dp/sl0/mxl/lph1  ( .q(\sc_dp/sl0/l1_q ), .d(
        \sc_dp/sl0/mxl/muxout ), .g(n8) );
    latn_1 \sc_tic/sl4/lph3  ( .q(TIC_d3_i_sc), .d(\sc_tic/sl4/l1_q ), .g(n3)
         );
    latn_1 \sc_tic/sl4/lph2  ( .q(\scan[2] ), .d(\sc_tic/sl4/l1_q ), .g(n6) );
    mux2_1 \sc_tic/sl4/mxl/mux  ( .x(\sc_tic/sl4/mxl/muxout ), .d0(TIC_d3_i), 
        .sl(n14), .d1(\sc_tic/scn4 ) );
    latn_1 \sc_tic/sl4/mxl/lph1  ( .q(\sc_tic/sl4/l1_q ), .d(
        \sc_tic/sl4/mxl/muxout ), .g(n10) );
    latn_1 \sc_tic/sl3/lph3  ( .q(TIC_d2_i_sc), .d(\sc_tic/sl3/l1_q ), .g(n3)
         );
    latn_1 \sc_tic/sl3/lph2  ( .q(\sc_tic/scn4 ), .d(\sc_tic/sl3/l1_q ), .g(n7
        ) );
    mux2_1 \sc_tic/sl3/mxl/mux  ( .x(\sc_tic/sl3/mxl/muxout ), .d0(TIC_d2_i), 
        .sl(n15), .d1(\sc_tic/scn3 ) );
    latn_1 \sc_tic/sl3/mxl/lph1  ( .q(\sc_tic/sl3/l1_q ), .d(
        \sc_tic/sl3/mxl/muxout ), .g(n11) );
    latn_1 \sc_tic/sl2/lph3  ( .q(TIC_d1_i_sc), .d(\sc_tic/sl2/l1_q ), .g(n3)
         );
    latn_1 \sc_tic/sl2/lph2  ( .q(\sc_tic/scn3 ), .d(\sc_tic/sl2/l1_q ), .g(n4
        ) );
    mux2_1 \sc_tic/sl2/mxl/mux  ( .x(\sc_tic/sl2/mxl/muxout ), .d0(TIC_d1_i), 
        .sl(n14), .d1(\sc_tic/scn2 ) );
    latn_1 \sc_tic/sl2/mxl/lph1  ( .q(\sc_tic/sl2/l1_q ), .d(
        \sc_tic/sl2/mxl/muxout ), .g(n8) );
    latn_1 \sc_tic/sl1/lph3  ( .q(TIC_d0_i_sc), .d(\sc_tic/sl1/l1_q ), .g(n3)
         );
    latn_1 \sc_tic/sl1/lph2  ( .q(\sc_tic/scn2 ), .d(\sc_tic/sl1/l1_q ), .g(n7
        ) );
    mux2_1 \sc_tic/sl1/mxl/mux  ( .x(\sc_tic/sl1/mxl/muxout ), .d0(TIC_d0_i), 
        .sl(n15), .d1(\sc_tic/scn1 ) );
    latn_1 \sc_tic/sl1/mxl/lph1  ( .q(\sc_tic/sl1/l1_q ), .d(
        \sc_tic/sl1/mxl/muxout ), .g(n11) );
    latn_1 \sc_tic/sl0/lph3  ( .q(TIC_eop_i_sc), .d(\sc_tic/sl0/l1_q ), .g(n1)
         );
    latn_1 \sc_tic/sl0/lph2  ( .q(\sc_tic/scn1 ), .d(\sc_tic/sl0/l1_q ), .g(n7
        ) );
    mux2_1 \sc_tic/sl0/mxl/mux  ( .x(\sc_tic/sl0/mxl/muxout ), .d0(TIC_eop_i), 
        .sl(n12), .d1(\scan[1] ) );
    latn_1 \sc_tic/sl0/mxl/lph1  ( .q(\sc_tic/sl0/l1_q ), .d(
        \sc_tic/sl0/mxl/muxout ), .g(n11) );
    latn_1 \sc_ip/sl4/lph3  ( .q(I_port_d3_i_sc), .d(\sc_ip/sl4/l1_q ), .g(n1)
         );
    latn_1 \sc_ip/sl4/lph2  ( .q(\scan[1] ), .d(\sc_ip/sl4/l1_q ), .g(n4) );
    mux2_1 \sc_ip/sl4/mxl/mux  ( .x(\sc_ip/sl4/mxl/muxout ), .d0(I_port_d3_i), 
        .sl(n12), .d1(\sc_ip/scn4 ) );
    latn_1 \sc_ip/sl4/mxl/lph1  ( .q(\sc_ip/sl4/l1_q ), .d(
        \sc_ip/sl4/mxl/muxout ), .g(n8) );
    latn_1 \sc_ip/sl3/lph3  ( .q(I_port_d2_i_sc), .d(\sc_ip/sl3/l1_q ), .g(n1)
         );
    latn_1 \sc_ip/sl3/lph2  ( .q(\sc_ip/scn4 ), .d(\sc_ip/sl3/l1_q ), .g(n6)
         );
    mux2_1 \sc_ip/sl3/mxl/mux  ( .x(\sc_ip/sl3/mxl/muxout ), .d0(I_port_d2_i), 
        .sl(n15), .d1(\sc_ip/scn3 ) );
    latn_1 \sc_ip/sl3/mxl/lph1  ( .q(\sc_ip/sl3/l1_q ), .d(
        \sc_ip/sl3/mxl/muxout ), .g(n10) );
    latn_1 \sc_ip/sl2/lph3  ( .q(I_port_d1_i_sc), .d(\sc_ip/sl2/l1_q ), .g(n1)
         );
    latn_1 \sc_ip/sl2/lph2  ( .q(\sc_ip/scn3 ), .d(\sc_ip/sl2/l1_q ), .g(n6)
         );
    mux2_1 \sc_ip/sl2/mxl/mux  ( .x(\sc_ip/sl2/mxl/muxout ), .d0(I_port_d1_i), 
        .sl(n14), .d1(\sc_ip/scn2 ) );
    latn_1 \sc_ip/sl2/mxl/lph1  ( .q(\sc_ip/sl2/l1_q ), .d(
        \sc_ip/sl2/mxl/muxout ), .g(n10) );
    latn_1 \sc_ip/sl1/lph3  ( .q(I_port_d0_i_sc), .d(\sc_ip/sl1/l1_q ), .g(n1)
         );
    latn_1 \sc_ip/sl1/lph2  ( .q(\sc_ip/scn2 ), .d(\sc_ip/sl1/l1_q ), .g(n4)
         );
    mux2_1 \sc_ip/sl1/mxl/mux  ( .x(\sc_ip/sl1/mxl/muxout ), .d0(I_port_d0_i), 
        .sl(n14), .d1(\sc_ip/scn1 ) );
    latn_1 \sc_ip/sl1/mxl/lph1  ( .q(\sc_ip/sl1/l1_q ), .d(
        \sc_ip/sl1/mxl/muxout ), .g(n8) );
    latn_1 \sc_ip/sl0/lph3  ( .q(I_port_eop_i_sc), .d(\sc_ip/sl0/l1_q ), .g(n1
        ) );
    latn_1 \sc_ip/sl0/lph2  ( .q(\sc_ip/scn1 ), .d(\sc_ip/sl0/l1_q ), .g(n6)
         );
    mux2_1 \sc_ip/sl0/mxl/mux  ( .x(\sc_ip/sl0/mxl/muxout ), .d0(I_port_eop_i), 
        .sl(n14), .d1(test_si) );
    latn_1 \sc_ip/sl0/mxl/lph1  ( .q(\sc_ip/sl0/l1_q ), .d(
        \sc_ip/sl0/mxl/muxout ), .g(n10) );
    buf_3 U1 ( .x(n13), .a(test_se) );
    buf_1 U2 ( .x(n1), .a(phi3) );
    buf_1 U3 ( .x(n3), .a(phi3) );
    buf_3 U4 ( .x(n2), .a(phi3) );
    buf_3 U5 ( .x(n4), .a(phi2) );
    buf_3 U6 ( .x(n7), .a(phi2) );
    buf_3 U7 ( .x(n5), .a(phi2) );
    buf_3 U8 ( .x(n6), .a(phi2) );
    buf_3 U9 ( .x(n8), .a(phi1) );
    buf_3 U10 ( .x(n11), .a(phi1) );
    buf_3 U11 ( .x(n9), .a(phi1) );
    buf_3 U12 ( .x(n10), .a(phi1) );
    buf_3 U13 ( .x(n12), .a(test_se) );
    buf_3 U14 ( .x(n15), .a(test_se) );
    buf_3 U15 ( .x(n14), .a(test_se) );
endmodule


module chain_arbiter10 ( eop_ix, d0_ix, d1_ix, d2_ix, d3_ix, ack_ix, eop_iy, 
    d0_iy, d1_iy, d2_iy, d3_iy, ack_iy, eop_ox, d0_ox, d1_ox, d2_ox, d3_ox, 
    eop_oy, d0_oy, d1_oy, d2_oy, d3_oy, ack_oxy, rst, test_si, test_se, 
    test_so, phi1, phi2, phi3 );
input  eop_ix, d0_ix, d1_ix, d2_ix, d3_ix, eop_iy, d0_iy, d1_iy, d2_iy, d3_iy, 
    ack_oxy, rst, test_si, test_se, phi1, phi2, phi3;
output ack_ix, ack_iy, eop_ox, d0_ox, d1_ox, d2_ox, d3_ox, eop_oy, d0_oy, 
    d1_oy, d2_oy, d3_oy, test_so;
    wire nack_x, ackx_l, n1x, n2x, nack_y, acky_l, n1y, n2y, req_x, n5x, n6x, 
        req_y, n5y, n6y, sx_pl, gx, sy_pl, gy, \cye/nr , sy, \cye/nd , 
        \cye/n2 , \cy3/__tmp99/loop , \cy2/__tmp99/loop , \cy1/__tmp99/loop , 
        \cy0/__tmp99/loop , \cxe/nr , sx, \cxe/nd , \cxe/n2 , 
        \cx3/__tmp99/loop , \cx2/__tmp99/loop , \cx1/__tmp99/loop , 
        \cx0/__tmp99/loop , \mtx/gr2 , mry, \mtx/gr1 , mrx, \sry/qz , \srx/qz , 
        \sl_sy/l1_q , \scan[1] , \sl_sy/mxl/muxout , \scan[0] , \sl_sx/l1_q , 
        \sl_sx/mxl/muxout , \slAcky/l1_q , \slAcky/mxl/muxout , \scan[2] , 
        \slAckx/l1_q , \slAckx/mxl/muxout ;
    nor2_2 U12 ( .x(nack_x), .a(ackx_l), .b(rst) );
    nand2_1 U4 ( .x(ack_ix), .a(n1x), .b(n2x) );
    nor3_1 U17 ( .x(n1x), .a(d2_ox), .b(d3_ox), .c(d1_ox) );
    nor2_1 U18 ( .x(n2x), .a(eop_ox), .b(d0_ox) );
    nor2_2 U11 ( .x(nack_y), .a(acky_l), .b(rst) );
    nand2_1 U3 ( .x(ack_iy), .a(n1y), .b(n2y) );
    nor3_1 U16 ( .x(n1y), .a(d2_oy), .b(d3_oy), .c(d1_oy) );
    nor2_1 U19 ( .x(n2y), .a(eop_oy), .b(d0_oy) );
    nand2_1 U15 ( .x(req_x), .a(n5x), .b(n6x) );
    nor3_1 U10 ( .x(n5x), .a(d2_ix), .b(d3_ix), .c(d1_ix) );
    nor2_1 U13 ( .x(n6x), .a(eop_ix), .b(d0_ix) );
    nand2_1 U14 ( .x(req_y), .a(n5y), .b(n6y) );
    nor3_1 U9 ( .x(n5y), .a(d2_iy), .b(d3_iy), .c(d1_iy) );
    nor2_1 U20 ( .x(n6y), .a(eop_iy), .b(d0_iy) );
    nor2i_1 U6 ( .x(sx_pl), .a(gx), .b(eop_oy) );
    nor2i_1 U5 ( .x(sy_pl), .a(gy), .b(eop_ox) );
    nor3_1 \cye/Unr  ( .x(\cye/nr ), .a(eop_iy), .b(nack_y), .c(sy) );
    nand3_1 \cye/Und  ( .x(\cye/nd ), .a(eop_iy), .b(nack_y), .c(sy) );
    oa21_1 \cye/U1  ( .x(\cye/n2 ), .a(\cye/n2 ), .b(\cye/nr ), .c(\cye/nd )
         );
    inv_1 \cye/U3  ( .x(eop_oy), .a(\cye/n2 ) );
    ao31_1 \cy3/__tmp99/aoi  ( .x(\cy3/__tmp99/loop ), .a(d3_iy), .b(nack_y), 
        .c(sy), .d(d3_oy) );
    oa21_1 \cy3/__tmp99/outGate  ( .x(d3_oy), .a(d3_iy), .b(nack_y), .c(
        \cy3/__tmp99/loop ) );
    ao31_1 \cy2/__tmp99/aoi  ( .x(\cy2/__tmp99/loop ), .a(d2_iy), .b(nack_y), 
        .c(sy), .d(d2_oy) );
    oa21_1 \cy2/__tmp99/outGate  ( .x(d2_oy), .a(d2_iy), .b(nack_y), .c(
        \cy2/__tmp99/loop ) );
    ao31_1 \cy1/__tmp99/aoi  ( .x(\cy1/__tmp99/loop ), .a(d1_iy), .b(nack_y), 
        .c(sy), .d(d1_oy) );
    oa21_1 \cy1/__tmp99/outGate  ( .x(d1_oy), .a(d1_iy), .b(nack_y), .c(
        \cy1/__tmp99/loop ) );
    ao31_1 \cy0/__tmp99/aoi  ( .x(\cy0/__tmp99/loop ), .a(d0_iy), .b(nack_y), 
        .c(sy), .d(d0_oy) );
    oa21_1 \cy0/__tmp99/outGate  ( .x(d0_oy), .a(d0_iy), .b(nack_y), .c(
        \cy0/__tmp99/loop ) );
    nor3_1 \cxe/Unr  ( .x(\cxe/nr ), .a(eop_ix), .b(nack_x), .c(sx) );
    nand3_1 \cxe/Und  ( .x(\cxe/nd ), .a(eop_ix), .b(nack_x), .c(sx) );
    oa21_1 \cxe/U1  ( .x(\cxe/n2 ), .a(\cxe/n2 ), .b(\cxe/nr ), .c(\cxe/nd )
         );
    inv_1 \cxe/U3  ( .x(eop_ox), .a(\cxe/n2 ) );
    ao31_1 \cx3/__tmp99/aoi  ( .x(\cx3/__tmp99/loop ), .a(d3_ix), .b(nack_x), 
        .c(sx), .d(d3_ox) );
    oa21_1 \cx3/__tmp99/outGate  ( .x(d3_ox), .a(d3_ix), .b(nack_x), .c(
        \cx3/__tmp99/loop ) );
    ao31_1 \cx2/__tmp99/aoi  ( .x(\cx2/__tmp99/loop ), .a(d2_ix), .b(nack_x), 
        .c(sx), .d(d2_ox) );
    oa21_1 \cx2/__tmp99/outGate  ( .x(d2_ox), .a(d2_ix), .b(nack_x), .c(
        \cx2/__tmp99/loop ) );
    ao31_1 \cx1/__tmp99/aoi  ( .x(\cx1/__tmp99/loop ), .a(d1_ix), .b(nack_x), 
        .c(sx), .d(d1_ox) );
    oa21_1 \cx1/__tmp99/outGate  ( .x(d1_ox), .a(d1_ix), .b(nack_x), .c(
        \cx1/__tmp99/loop ) );
    ao31_1 \cx0/__tmp99/aoi  ( .x(\cx0/__tmp99/loop ), .a(d0_ix), .b(nack_x), 
        .c(sx), .d(d0_ox) );
    oa21_1 \cx0/__tmp99/outGate  ( .x(d0_ox), .a(d0_ix), .b(nack_x), .c(
        \cx0/__tmp99/loop ) );
    nand2_1 \mtx/mg2  ( .x(\mtx/gr2 ), .a(mry), .b(\mtx/gr1 ) );
    nand2_1 \mtx/U1  ( .x(\mtx/gr1 ), .a(mrx), .b(\mtx/gr2 ) );
    nor3_1 \mtx/U2  ( .x(gy), .a(\mtx/gr2 ), .b(\mtx/gr2 ), .c(\mtx/gr2 ) );
    nor3_1 \mtx/U3  ( .x(gx), .a(\mtx/gr1 ), .b(\mtx/gr1 ), .c(\mtx/gr1 ) );
    nor2_1 \sry/i1  ( .x(\sry/qz ), .a(req_y), .b(mry) );
    nor2_1 \srx/i1  ( .x(\srx/qz ), .a(req_x), .b(mrx) );
    latn_1 \sl_sy/lph3  ( .q(sy), .d(\sl_sy/l1_q ), .g(phi3) );
    latn_1 \sl_sy/lph2  ( .q(\scan[1] ), .d(\sl_sy/l1_q ), .g(phi2) );
    mux2_1 \sl_sy/mxl/mux  ( .x(\sl_sy/mxl/muxout ), .d0(sy_pl), .sl(test_se), 
        .d1(\scan[0] ) );
    latn_1 \sl_sy/mxl/lph1  ( .q(\sl_sy/l1_q ), .d(\sl_sy/mxl/muxout ), .g(
        phi1) );
    latn_1 \sl_sx/lph3  ( .q(sx), .d(\sl_sx/l1_q ), .g(phi3) );
    latn_1 \sl_sx/lph2  ( .q(\scan[0] ), .d(\sl_sx/l1_q ), .g(phi2) );
    mux2_1 \sl_sx/mxl/mux  ( .x(\sl_sx/mxl/muxout ), .d0(sx_pl), .sl(test_se), 
        .d1(test_si) );
    latn_1 \sl_sx/mxl/lph1  ( .q(\sl_sx/l1_q ), .d(\sl_sx/mxl/muxout ), .g(
        phi1) );
    latn_1 \slAcky/lph3  ( .q(acky_l), .d(\slAcky/l1_q ), .g(phi3) );
    latn_1 \slAcky/lph2  ( .q(test_so), .d(\slAcky/l1_q ), .g(phi2) );
    mux2_1 \slAcky/mxl/mux  ( .x(\slAcky/mxl/muxout ), .d0(ack_oxy), .sl(
        test_se), .d1(\scan[2] ) );
    latn_1 \slAcky/mxl/lph1  ( .q(\slAcky/l1_q ), .d(\slAcky/mxl/muxout ), .g(
        phi1) );
    latn_1 \slAckx/lph3  ( .q(ackx_l), .d(\slAckx/l1_q ), .g(phi3) );
    latn_1 \slAckx/lph2  ( .q(\scan[2] ), .d(\slAckx/l1_q ), .g(phi2) );
    mux2_1 \slAckx/mxl/mux  ( .x(\slAckx/mxl/muxout ), .d0(ack_oxy), .sl(
        test_se), .d1(\scan[1] ) );
    latn_1 \slAckx/mxl/lph1  ( .q(\slAckx/l1_q ), .d(\slAckx/mxl/muxout ), .g(
        phi1) );
    nor3_1 U1 ( .x(mry), .a(eop_oy), .b(rst), .c(\sry/qz ) );
    nor3_1 U2 ( .x(mrx), .a(eop_ox), .b(rst), .c(\srx/qz ) );
endmodule


module chain_mux10 ( eop_ix, d0_ix, d1_ix, d2_ix, d3_ix, ack_ixy, eop_iy, 
    d0_iy, d1_iy, d2_iy, d3_iy, eop_o, d0_o, d1_o, d2_o, d3_o, ack_o, rst, 
    test_si, test_se, test_so, phi1, phi2, phi3 );
input  eop_ix, d0_ix, d1_ix, d2_ix, d3_ix, eop_iy, d0_iy, d1_iy, d2_iy, d3_iy, 
    ack_o, rst, test_si, test_se, phi1, phi2, phi3;
output ack_ixy, eop_o, d0_o, d1_o, d2_o, d3_o, test_so;
    wire d3_i, d2_i, d1_i, d0_i, eop_i, n1, n2, \ce/ob , ack, \c3/ob , \c2/ob , 
        \c1/ob , \c0/ob , ack_l, \slAck/l1_q , \slAck/mxl/muxout ;
    nor2_1 U2 ( .x(d3_i), .a(d3_iy), .b(d3_ix) );
    nor2_1 U3 ( .x(d2_i), .a(d2_iy), .b(d2_ix) );
    nor2_1 U4 ( .x(d1_i), .a(d1_iy), .b(d1_ix) );
    nor2_1 U5 ( .x(d0_i), .a(d0_iy), .b(d0_ix) );
    nor2_1 U6 ( .x(eop_i), .a(eop_iy), .b(eop_ix) );
    nand2_1 U1 ( .x(ack_ixy), .a(n1), .b(n2) );
    nor3_1 U9 ( .x(n1), .a(d2_o), .b(d3_o), .c(d1_o) );
    nor2_1 U8 ( .x(n2), .a(eop_o), .b(d0_o) );
    inv_1 \ce/Ui  ( .x(\ce/ob ), .a(eop_o) );
    aoi222_1 \ce/__tmp99/U1  ( .x(eop_o), .a(eop_i), .b(ack), .c(eop_i), .d(
        \ce/ob ), .e(ack), .f(\ce/ob ) );
    inv_1 \c3/Ui  ( .x(\c3/ob ), .a(d3_o) );
    aoi222_1 \c3/__tmp99/U1  ( .x(d3_o), .a(d3_i), .b(ack), .c(d3_i), .d(
        \c3/ob ), .e(ack), .f(\c3/ob ) );
    inv_1 \c2/Ui  ( .x(\c2/ob ), .a(d2_o) );
    aoi222_1 \c2/__tmp99/U1  ( .x(d2_o), .a(d2_i), .b(ack), .c(d2_i), .d(
        \c2/ob ), .e(ack), .f(\c2/ob ) );
    inv_1 \c1/Ui  ( .x(\c1/ob ), .a(d1_o) );
    aoi222_1 \c1/__tmp99/U1  ( .x(d1_o), .a(d1_i), .b(ack), .c(d1_i), .d(
        \c1/ob ), .e(ack), .f(\c1/ob ) );
    inv_1 \c0/Ui  ( .x(\c0/ob ), .a(d0_o) );
    aoi222_1 \c0/__tmp99/U1  ( .x(d0_o), .a(d0_i), .b(ack), .c(d0_i), .d(
        \c0/ob ), .e(ack), .f(\c0/ob ) );
    latn_1 \slAck/lph3  ( .q(ack_l), .d(\slAck/l1_q ), .g(phi3) );
    latn_1 \slAck/lph2  ( .q(test_so), .d(\slAck/l1_q ), .g(phi2) );
    mux2_1 \slAck/mxl/mux  ( .x(\slAck/mxl/muxout ), .d0(ack_o), .sl(test_se), 
        .d1(test_si) );
    latn_1 \slAck/mxl/lph1  ( .q(\slAck/l1_q ), .d(\slAck/mxl/muxout ), .g(
        phi1) );
    or2_4 U7 ( .x(ack), .a(ack_l), .b(rst) );
endmodule


module chain_arbiter11 ( eop_ix, d0_ix, d1_ix, d2_ix, d3_ix, ack_ix, eop_iy, 
    d0_iy, d1_iy, d2_iy, d3_iy, ack_iy, eop_ox, d0_ox, d1_ox, d2_ox, d3_ox, 
    eop_oy, d0_oy, d1_oy, d2_oy, d3_oy, ack_oxy, rst, test_si, test_se, 
    test_so, phi1, phi2, phi3 );
input  eop_ix, d0_ix, d1_ix, d2_ix, d3_ix, eop_iy, d0_iy, d1_iy, d2_iy, d3_iy, 
    ack_oxy, rst, test_si, test_se, phi1, phi2, phi3;
output ack_ix, ack_iy, eop_ox, d0_ox, d1_ox, d2_ox, d3_ox, eop_oy, d0_oy, 
    d1_oy, d2_oy, d3_oy, test_so;
    wire nack_x, ackx_l, n1x, n2x, nack_y, acky_l, n1y, n2y, req_x, n5x, n6x, 
        req_y, n5y, n6y, sx_pl, gx, sy_pl, gy, \cye/nr , sy, \cye/nd , 
        \cye/n2 , \cy3/__tmp99/loop , \cy2/__tmp99/loop , \cy1/__tmp99/loop , 
        \cy0/__tmp99/loop , \cxe/nr , sx, \cxe/nd , \cxe/n2 , 
        \cx3/__tmp99/loop , \cx2/__tmp99/loop , \cx1/__tmp99/loop , 
        \cx0/__tmp99/loop , \mtx/gr2 , mry, \mtx/gr1 , mrx, \sry/qz , \srx/qz , 
        \sl_sy/l1_q , \scan[1] , \sl_sy/mxl/muxout , \scan[0] , \sl_sx/l1_q , 
        \sl_sx/mxl/muxout , \slAcky/l1_q , \slAcky/mxl/muxout , \scan[2] , 
        \slAckx/l1_q , \slAckx/mxl/muxout ;
    nor2_2 U12 ( .x(nack_x), .a(ackx_l), .b(rst) );
    nand2_1 U4 ( .x(ack_ix), .a(n1x), .b(n2x) );
    nor3_1 U17 ( .x(n1x), .a(d2_ox), .b(d3_ox), .c(d1_ox) );
    nor2_1 U18 ( .x(n2x), .a(eop_ox), .b(d0_ox) );
    nor2_2 U11 ( .x(nack_y), .a(acky_l), .b(rst) );
    nand2_1 U3 ( .x(ack_iy), .a(n1y), .b(n2y) );
    nor3_1 U16 ( .x(n1y), .a(d2_oy), .b(d3_oy), .c(d1_oy) );
    nor2_1 U19 ( .x(n2y), .a(eop_oy), .b(d0_oy) );
    nand2_1 U15 ( .x(req_x), .a(n5x), .b(n6x) );
    nor3_1 U10 ( .x(n5x), .a(d2_ix), .b(d3_ix), .c(d1_ix) );
    nor2_1 U13 ( .x(n6x), .a(eop_ix), .b(d0_ix) );
    nand2_1 U14 ( .x(req_y), .a(n5y), .b(n6y) );
    nor3_1 U9 ( .x(n5y), .a(d2_iy), .b(d3_iy), .c(d1_iy) );
    nor2_1 U20 ( .x(n6y), .a(eop_iy), .b(d0_iy) );
    nor2i_1 U6 ( .x(sx_pl), .a(gx), .b(eop_oy) );
    nor2i_1 U5 ( .x(sy_pl), .a(gy), .b(eop_ox) );
    nor3_1 \cye/Unr  ( .x(\cye/nr ), .a(eop_iy), .b(nack_y), .c(sy) );
    nand3_1 \cye/Und  ( .x(\cye/nd ), .a(eop_iy), .b(nack_y), .c(sy) );
    oa21_1 \cye/U1  ( .x(\cye/n2 ), .a(\cye/n2 ), .b(\cye/nr ), .c(\cye/nd )
         );
    inv_1 \cye/U3  ( .x(eop_oy), .a(\cye/n2 ) );
    ao31_1 \cy3/__tmp99/aoi  ( .x(\cy3/__tmp99/loop ), .a(d3_iy), .b(nack_y), 
        .c(sy), .d(d3_oy) );
    oa21_1 \cy3/__tmp99/outGate  ( .x(d3_oy), .a(d3_iy), .b(nack_y), .c(
        \cy3/__tmp99/loop ) );
    ao31_1 \cy2/__tmp99/aoi  ( .x(\cy2/__tmp99/loop ), .a(d2_iy), .b(nack_y), 
        .c(sy), .d(d2_oy) );
    oa21_1 \cy2/__tmp99/outGate  ( .x(d2_oy), .a(d2_iy), .b(nack_y), .c(
        \cy2/__tmp99/loop ) );
    ao31_1 \cy1/__tmp99/aoi  ( .x(\cy1/__tmp99/loop ), .a(d1_iy), .b(nack_y), 
        .c(sy), .d(d1_oy) );
    oa21_1 \cy1/__tmp99/outGate  ( .x(d1_oy), .a(d1_iy), .b(nack_y), .c(
        \cy1/__tmp99/loop ) );
    ao31_1 \cy0/__tmp99/aoi  ( .x(\cy0/__tmp99/loop ), .a(d0_iy), .b(nack_y), 
        .c(sy), .d(d0_oy) );
    oa21_1 \cy0/__tmp99/outGate  ( .x(d0_oy), .a(d0_iy), .b(nack_y), .c(
        \cy0/__tmp99/loop ) );
    nor3_1 \cxe/Unr  ( .x(\cxe/nr ), .a(eop_ix), .b(nack_x), .c(sx) );
    nand3_1 \cxe/Und  ( .x(\cxe/nd ), .a(eop_ix), .b(nack_x), .c(sx) );
    oa21_1 \cxe/U1  ( .x(\cxe/n2 ), .a(\cxe/n2 ), .b(\cxe/nr ), .c(\cxe/nd )
         );
    inv_1 \cxe/U3  ( .x(eop_ox), .a(\cxe/n2 ) );
    ao31_1 \cx3/__tmp99/aoi  ( .x(\cx3/__tmp99/loop ), .a(d3_ix), .b(nack_x), 
        .c(sx), .d(d3_ox) );
    oa21_1 \cx3/__tmp99/outGate  ( .x(d3_ox), .a(d3_ix), .b(nack_x), .c(
        \cx3/__tmp99/loop ) );
    ao31_1 \cx2/__tmp99/aoi  ( .x(\cx2/__tmp99/loop ), .a(d2_ix), .b(nack_x), 
        .c(sx), .d(d2_ox) );
    oa21_1 \cx2/__tmp99/outGate  ( .x(d2_ox), .a(d2_ix), .b(nack_x), .c(
        \cx2/__tmp99/loop ) );
    ao31_1 \cx1/__tmp99/aoi  ( .x(\cx1/__tmp99/loop ), .a(d1_ix), .b(nack_x), 
        .c(sx), .d(d1_ox) );
    oa21_1 \cx1/__tmp99/outGate  ( .x(d1_ox), .a(d1_ix), .b(nack_x), .c(
        \cx1/__tmp99/loop ) );
    ao31_1 \cx0/__tmp99/aoi  ( .x(\cx0/__tmp99/loop ), .a(d0_ix), .b(nack_x), 
        .c(sx), .d(d0_ox) );
    oa21_1 \cx0/__tmp99/outGate  ( .x(d0_ox), .a(d0_ix), .b(nack_x), .c(
        \cx0/__tmp99/loop ) );
    nand2_1 \mtx/mg2  ( .x(\mtx/gr2 ), .a(mry), .b(\mtx/gr1 ) );
    nand2_1 \mtx/U1  ( .x(\mtx/gr1 ), .a(mrx), .b(\mtx/gr2 ) );
    nor3_1 \mtx/U2  ( .x(gy), .a(\mtx/gr2 ), .b(\mtx/gr2 ), .c(\mtx/gr2 ) );
    nor3_1 \mtx/U3  ( .x(gx), .a(\mtx/gr1 ), .b(\mtx/gr1 ), .c(\mtx/gr1 ) );
    nor2_1 \sry/i1  ( .x(\sry/qz ), .a(req_y), .b(mry) );
    nor2_1 \srx/i1  ( .x(\srx/qz ), .a(req_x), .b(mrx) );
    latn_1 \sl_sy/lph3  ( .q(sy), .d(\sl_sy/l1_q ), .g(phi3) );
    latn_1 \sl_sy/lph2  ( .q(\scan[1] ), .d(\sl_sy/l1_q ), .g(phi2) );
    mux2_1 \sl_sy/mxl/mux  ( .x(\sl_sy/mxl/muxout ), .d0(sy_pl), .sl(test_se), 
        .d1(\scan[0] ) );
    latn_1 \sl_sy/mxl/lph1  ( .q(\sl_sy/l1_q ), .d(\sl_sy/mxl/muxout ), .g(
        phi1) );
    latn_1 \sl_sx/lph3  ( .q(sx), .d(\sl_sx/l1_q ), .g(phi3) );
    latn_1 \sl_sx/lph2  ( .q(\scan[0] ), .d(\sl_sx/l1_q ), .g(phi2) );
    mux2_1 \sl_sx/mxl/mux  ( .x(\sl_sx/mxl/muxout ), .d0(sx_pl), .sl(test_se), 
        .d1(test_si) );
    latn_1 \sl_sx/mxl/lph1  ( .q(\sl_sx/l1_q ), .d(\sl_sx/mxl/muxout ), .g(
        phi1) );
    latn_1 \slAcky/lph3  ( .q(acky_l), .d(\slAcky/l1_q ), .g(phi3) );
    latn_1 \slAcky/lph2  ( .q(test_so), .d(\slAcky/l1_q ), .g(phi2) );
    mux2_1 \slAcky/mxl/mux  ( .x(\slAcky/mxl/muxout ), .d0(ack_oxy), .sl(
        test_se), .d1(\scan[2] ) );
    latn_1 \slAcky/mxl/lph1  ( .q(\slAcky/l1_q ), .d(\slAcky/mxl/muxout ), .g(
        phi1) );
    latn_1 \slAckx/lph3  ( .q(ackx_l), .d(\slAckx/l1_q ), .g(phi3) );
    latn_1 \slAckx/lph2  ( .q(\scan[2] ), .d(\slAckx/l1_q ), .g(phi2) );
    mux2_1 \slAckx/mxl/mux  ( .x(\slAckx/mxl/muxout ), .d0(ack_oxy), .sl(
        test_se), .d1(\scan[1] ) );
    latn_1 \slAckx/mxl/lph1  ( .q(\slAckx/l1_q ), .d(\slAckx/mxl/muxout ), .g(
        phi1) );
    nor3_1 U1 ( .x(mrx), .a(eop_ox), .b(rst), .c(\srx/qz ) );
    nor3_1 U2 ( .x(mry), .a(eop_oy), .b(rst), .c(\sry/qz ) );
endmodule


module chain_mux11 ( eop_ix, d0_ix, d1_ix, d2_ix, d3_ix, ack_ixy, eop_iy, 
    d0_iy, d1_iy, d2_iy, d3_iy, eop_o, d0_o, d1_o, d2_o, d3_o, ack_o, rst, 
    test_si, test_se, test_so, phi1, phi2, phi3 );
input  eop_ix, d0_ix, d1_ix, d2_ix, d3_ix, eop_iy, d0_iy, d1_iy, d2_iy, d3_iy, 
    ack_o, rst, test_si, test_se, phi1, phi2, phi3;
output ack_ixy, eop_o, d0_o, d1_o, d2_o, d3_o, test_so;
    wire d3_i, d2_i, d1_i, d0_i, eop_i, n1, n2, \ce/ob , ack, \c3/ob , \c2/ob , 
        \c1/ob , \c0/ob , ack_l, \slAck/l1_q , \slAck/mxl/muxout ;
    nor2_1 U2 ( .x(d3_i), .a(d3_iy), .b(d3_ix) );
    nor2_1 U3 ( .x(d2_i), .a(d2_iy), .b(d2_ix) );
    nor2_1 U4 ( .x(d1_i), .a(d1_iy), .b(d1_ix) );
    nor2_1 U5 ( .x(d0_i), .a(d0_iy), .b(d0_ix) );
    nor2_1 U6 ( .x(eop_i), .a(eop_iy), .b(eop_ix) );
    nand2_1 U1 ( .x(ack_ixy), .a(n1), .b(n2) );
    nor3_1 U9 ( .x(n1), .a(d2_o), .b(d3_o), .c(d1_o) );
    nor2_1 U8 ( .x(n2), .a(eop_o), .b(d0_o) );
    inv_1 \ce/Ui  ( .x(\ce/ob ), .a(eop_o) );
    aoi222_1 \ce/__tmp99/U1  ( .x(eop_o), .a(eop_i), .b(ack), .c(eop_i), .d(
        \ce/ob ), .e(ack), .f(\ce/ob ) );
    inv_1 \c3/Ui  ( .x(\c3/ob ), .a(d3_o) );
    aoi222_1 \c3/__tmp99/U1  ( .x(d3_o), .a(d3_i), .b(ack), .c(d3_i), .d(
        \c3/ob ), .e(ack), .f(\c3/ob ) );
    inv_1 \c2/Ui  ( .x(\c2/ob ), .a(d2_o) );
    aoi222_1 \c2/__tmp99/U1  ( .x(d2_o), .a(d2_i), .b(ack), .c(d2_i), .d(
        \c2/ob ), .e(ack), .f(\c2/ob ) );
    inv_1 \c1/Ui  ( .x(\c1/ob ), .a(d1_o) );
    aoi222_1 \c1/__tmp99/U1  ( .x(d1_o), .a(d1_i), .b(ack), .c(d1_i), .d(
        \c1/ob ), .e(ack), .f(\c1/ob ) );
    inv_1 \c0/Ui  ( .x(\c0/ob ), .a(d0_o) );
    aoi222_1 \c0/__tmp99/U1  ( .x(d0_o), .a(d0_i), .b(ack), .c(d0_i), .d(
        \c0/ob ), .e(ack), .f(\c0/ob ) );
    latn_1 \slAck/lph3  ( .q(ack_l), .d(\slAck/l1_q ), .g(phi3) );
    latn_1 \slAck/lph2  ( .q(test_so), .d(\slAck/l1_q ), .g(phi2) );
    mux2_1 \slAck/mxl/mux  ( .x(\slAck/mxl/muxout ), .d0(ack_o), .sl(test_se), 
        .d1(test_si) );
    latn_1 \slAck/mxl/lph1  ( .q(\slAck/l1_q ), .d(\slAck/mxl/muxout ), .g(
        phi1) );
    or2_4 U7 ( .x(ack), .a(ack_l), .b(rst) );
endmodule


module chain_arbiter12 ( eop_ix, d0_ix, d1_ix, d2_ix, d3_ix, ack_ix, eop_iy, 
    d0_iy, d1_iy, d2_iy, d3_iy, ack_iy, eop_ox, d0_ox, d1_ox, d2_ox, d3_ox, 
    eop_oy, d0_oy, d1_oy, d2_oy, d3_oy, ack_oxy, rst, test_si, test_se, 
    test_so, phi1, phi2, phi3 );
input  eop_ix, d0_ix, d1_ix, d2_ix, d3_ix, eop_iy, d0_iy, d1_iy, d2_iy, d3_iy, 
    ack_oxy, rst, test_si, test_se, phi1, phi2, phi3;
output ack_ix, ack_iy, eop_ox, d0_ox, d1_ox, d2_ox, d3_ox, eop_oy, d0_oy, 
    d1_oy, d2_oy, d3_oy, test_so;
    wire nack_x, ackx_l, n1x, n2x, nack_y, acky_l, n1y, n2y, req_x, n5x, n6x, 
        req_y, n5y, n6y, sx_pl, gx, sy_pl, gy, \cye/nr , sy, \cye/nd , 
        \cye/n2 , \cy3/__tmp99/loop , \cy2/__tmp99/loop , \cy1/__tmp99/loop , 
        \cy0/__tmp99/loop , \cxe/nr , sx, \cxe/nd , \cxe/n2 , 
        \cx3/__tmp99/loop , \cx2/__tmp99/loop , \cx1/__tmp99/loop , 
        \cx0/__tmp99/loop , \mtx/gr2 , mry, \mtx/gr1 , mrx, \sry/qz , \srx/qz , 
        \sl_sy/l1_q , \scan[1] , \sl_sy/mxl/muxout , \scan[0] , \sl_sx/l1_q , 
        \sl_sx/mxl/muxout , \slAcky/l1_q , \slAcky/mxl/muxout , \scan[2] , 
        \slAckx/l1_q , \slAckx/mxl/muxout ;
    nor2_2 U12 ( .x(nack_x), .a(ackx_l), .b(rst) );
    nand2_1 U4 ( .x(ack_ix), .a(n1x), .b(n2x) );
    nor3_1 U17 ( .x(n1x), .a(d2_ox), .b(d3_ox), .c(d1_ox) );
    nor2_1 U18 ( .x(n2x), .a(eop_ox), .b(d0_ox) );
    nor2_2 U11 ( .x(nack_y), .a(acky_l), .b(rst) );
    nand2_1 U3 ( .x(ack_iy), .a(n1y), .b(n2y) );
    nor3_1 U16 ( .x(n1y), .a(d2_oy), .b(d3_oy), .c(d1_oy) );
    nor2_1 U19 ( .x(n2y), .a(eop_oy), .b(d0_oy) );
    nand2_1 U15 ( .x(req_x), .a(n5x), .b(n6x) );
    nor3_1 U10 ( .x(n5x), .a(d2_ix), .b(d3_ix), .c(d1_ix) );
    nor2_1 U13 ( .x(n6x), .a(eop_ix), .b(d0_ix) );
    nand2_1 U14 ( .x(req_y), .a(n5y), .b(n6y) );
    nor3_1 U9 ( .x(n5y), .a(d2_iy), .b(d3_iy), .c(d1_iy) );
    nor2_1 U20 ( .x(n6y), .a(eop_iy), .b(d0_iy) );
    nor2i_1 U6 ( .x(sx_pl), .a(gx), .b(eop_oy) );
    nor2i_1 U5 ( .x(sy_pl), .a(gy), .b(eop_ox) );
    nor3_1 \cye/Unr  ( .x(\cye/nr ), .a(eop_iy), .b(nack_y), .c(sy) );
    nand3_1 \cye/Und  ( .x(\cye/nd ), .a(eop_iy), .b(nack_y), .c(sy) );
    oa21_1 \cye/U1  ( .x(\cye/n2 ), .a(\cye/n2 ), .b(\cye/nr ), .c(\cye/nd )
         );
    inv_1 \cye/U3  ( .x(eop_oy), .a(\cye/n2 ) );
    ao31_1 \cy3/__tmp99/aoi  ( .x(\cy3/__tmp99/loop ), .a(d3_iy), .b(nack_y), 
        .c(sy), .d(d3_oy) );
    oa21_1 \cy3/__tmp99/outGate  ( .x(d3_oy), .a(d3_iy), .b(nack_y), .c(
        \cy3/__tmp99/loop ) );
    ao31_1 \cy2/__tmp99/aoi  ( .x(\cy2/__tmp99/loop ), .a(d2_iy), .b(nack_y), 
        .c(sy), .d(d2_oy) );
    oa21_1 \cy2/__tmp99/outGate  ( .x(d2_oy), .a(d2_iy), .b(nack_y), .c(
        \cy2/__tmp99/loop ) );
    ao31_1 \cy1/__tmp99/aoi  ( .x(\cy1/__tmp99/loop ), .a(d1_iy), .b(nack_y), 
        .c(sy), .d(d1_oy) );
    oa21_1 \cy1/__tmp99/outGate  ( .x(d1_oy), .a(d1_iy), .b(nack_y), .c(
        \cy1/__tmp99/loop ) );
    ao31_1 \cy0/__tmp99/aoi  ( .x(\cy0/__tmp99/loop ), .a(d0_iy), .b(nack_y), 
        .c(sy), .d(d0_oy) );
    oa21_1 \cy0/__tmp99/outGate  ( .x(d0_oy), .a(d0_iy), .b(nack_y), .c(
        \cy0/__tmp99/loop ) );
    nor3_1 \cxe/Unr  ( .x(\cxe/nr ), .a(eop_ix), .b(nack_x), .c(sx) );
    nand3_1 \cxe/Und  ( .x(\cxe/nd ), .a(eop_ix), .b(nack_x), .c(sx) );
    oa21_1 \cxe/U1  ( .x(\cxe/n2 ), .a(\cxe/n2 ), .b(\cxe/nr ), .c(\cxe/nd )
         );
    inv_1 \cxe/U3  ( .x(eop_ox), .a(\cxe/n2 ) );
    ao31_1 \cx3/__tmp99/aoi  ( .x(\cx3/__tmp99/loop ), .a(d3_ix), .b(nack_x), 
        .c(sx), .d(d3_ox) );
    oa21_1 \cx3/__tmp99/outGate  ( .x(d3_ox), .a(d3_ix), .b(nack_x), .c(
        \cx3/__tmp99/loop ) );
    ao31_1 \cx2/__tmp99/aoi  ( .x(\cx2/__tmp99/loop ), .a(d2_ix), .b(nack_x), 
        .c(sx), .d(d2_ox) );
    oa21_1 \cx2/__tmp99/outGate  ( .x(d2_ox), .a(d2_ix), .b(nack_x), .c(
        \cx2/__tmp99/loop ) );
    ao31_1 \cx1/__tmp99/aoi  ( .x(\cx1/__tmp99/loop ), .a(d1_ix), .b(nack_x), 
        .c(sx), .d(d1_ox) );
    oa21_1 \cx1/__tmp99/outGate  ( .x(d1_ox), .a(d1_ix), .b(nack_x), .c(
        \cx1/__tmp99/loop ) );
    ao31_1 \cx0/__tmp99/aoi  ( .x(\cx0/__tmp99/loop ), .a(d0_ix), .b(nack_x), 
        .c(sx), .d(d0_ox) );
    oa21_1 \cx0/__tmp99/outGate  ( .x(d0_ox), .a(d0_ix), .b(nack_x), .c(
        \cx0/__tmp99/loop ) );
    nand2_1 \mtx/mg2  ( .x(\mtx/gr2 ), .a(mry), .b(\mtx/gr1 ) );
    nand2_1 \mtx/U1  ( .x(\mtx/gr1 ), .a(mrx), .b(\mtx/gr2 ) );
    nor3_1 \mtx/U2  ( .x(gy), .a(\mtx/gr2 ), .b(\mtx/gr2 ), .c(\mtx/gr2 ) );
    nor3_1 \mtx/U3  ( .x(gx), .a(\mtx/gr1 ), .b(\mtx/gr1 ), .c(\mtx/gr1 ) );
    nor2_1 \sry/i1  ( .x(\sry/qz ), .a(req_y), .b(mry) );
    nor2_1 \srx/i1  ( .x(\srx/qz ), .a(req_x), .b(mrx) );
    latn_1 \sl_sy/lph3  ( .q(sy), .d(\sl_sy/l1_q ), .g(phi3) );
    latn_1 \sl_sy/lph2  ( .q(\scan[1] ), .d(\sl_sy/l1_q ), .g(phi2) );
    mux2_1 \sl_sy/mxl/mux  ( .x(\sl_sy/mxl/muxout ), .d0(sy_pl), .sl(test_se), 
        .d1(\scan[0] ) );
    latn_1 \sl_sy/mxl/lph1  ( .q(\sl_sy/l1_q ), .d(\sl_sy/mxl/muxout ), .g(
        phi1) );
    latn_1 \sl_sx/lph3  ( .q(sx), .d(\sl_sx/l1_q ), .g(phi3) );
    latn_1 \sl_sx/lph2  ( .q(\scan[0] ), .d(\sl_sx/l1_q ), .g(phi2) );
    mux2_1 \sl_sx/mxl/mux  ( .x(\sl_sx/mxl/muxout ), .d0(sx_pl), .sl(test_se), 
        .d1(test_si) );
    latn_1 \sl_sx/mxl/lph1  ( .q(\sl_sx/l1_q ), .d(\sl_sx/mxl/muxout ), .g(
        phi1) );
    latn_1 \slAcky/lph3  ( .q(acky_l), .d(\slAcky/l1_q ), .g(phi3) );
    latn_1 \slAcky/lph2  ( .q(test_so), .d(\slAcky/l1_q ), .g(phi2) );
    mux2_1 \slAcky/mxl/mux  ( .x(\slAcky/mxl/muxout ), .d0(ack_oxy), .sl(
        test_se), .d1(\scan[2] ) );
    latn_1 \slAcky/mxl/lph1  ( .q(\slAcky/l1_q ), .d(\slAcky/mxl/muxout ), .g(
        phi1) );
    latn_1 \slAckx/lph3  ( .q(ackx_l), .d(\slAckx/l1_q ), .g(phi3) );
    latn_1 \slAckx/lph2  ( .q(\scan[2] ), .d(\slAckx/l1_q ), .g(phi2) );
    mux2_1 \slAckx/mxl/mux  ( .x(\slAckx/mxl/muxout ), .d0(ack_oxy), .sl(
        test_se), .d1(\scan[1] ) );
    latn_1 \slAckx/mxl/lph1  ( .q(\slAckx/l1_q ), .d(\slAckx/mxl/muxout ), .g(
        phi1) );
    nor3_1 U1 ( .x(mry), .a(eop_oy), .b(rst), .c(\sry/qz ) );
    nor3_1 U2 ( .x(mrx), .a(eop_ox), .b(rst), .c(\srx/qz ) );
endmodule


module chain_mux12 ( eop_ix, d0_ix, d1_ix, d2_ix, d3_ix, ack_ixy, eop_iy, 
    d0_iy, d1_iy, d2_iy, d3_iy, eop_o, d0_o, d1_o, d2_o, d3_o, ack_o, rst, 
    test_si, test_se, test_so, phi1, phi2, phi3 );
input  eop_ix, d0_ix, d1_ix, d2_ix, d3_ix, eop_iy, d0_iy, d1_iy, d2_iy, d3_iy, 
    ack_o, rst, test_si, test_se, phi1, phi2, phi3;
output ack_ixy, eop_o, d0_o, d1_o, d2_o, d3_o, test_so;
    wire d3_i, d2_i, d1_i, d0_i, eop_i, n1, n2, \ce/ob , ack, \c3/ob , \c2/ob , 
        \c1/ob , \c0/ob , ack_l, \slAck/l1_q , \slAck/mxl/muxout ;
    nor2_1 U2 ( .x(d3_i), .a(d3_iy), .b(d3_ix) );
    nor2_1 U3 ( .x(d2_i), .a(d2_iy), .b(d2_ix) );
    nor2_1 U4 ( .x(d1_i), .a(d1_iy), .b(d1_ix) );
    nor2_1 U5 ( .x(d0_i), .a(d0_iy), .b(d0_ix) );
    nor2_1 U6 ( .x(eop_i), .a(eop_iy), .b(eop_ix) );
    nand2_1 U1 ( .x(ack_ixy), .a(n1), .b(n2) );
    nor3_1 U9 ( .x(n1), .a(d2_o), .b(d3_o), .c(d1_o) );
    nor2_1 U8 ( .x(n2), .a(eop_o), .b(d0_o) );
    inv_1 \ce/Ui  ( .x(\ce/ob ), .a(eop_o) );
    aoi222_1 \ce/__tmp99/U1  ( .x(eop_o), .a(eop_i), .b(ack), .c(eop_i), .d(
        \ce/ob ), .e(ack), .f(\ce/ob ) );
    inv_1 \c3/Ui  ( .x(\c3/ob ), .a(d3_o) );
    aoi222_1 \c3/__tmp99/U1  ( .x(d3_o), .a(d3_i), .b(ack), .c(d3_i), .d(
        \c3/ob ), .e(ack), .f(\c3/ob ) );
    inv_1 \c2/Ui  ( .x(\c2/ob ), .a(d2_o) );
    aoi222_1 \c2/__tmp99/U1  ( .x(d2_o), .a(d2_i), .b(ack), .c(d2_i), .d(
        \c2/ob ), .e(ack), .f(\c2/ob ) );
    inv_1 \c1/Ui  ( .x(\c1/ob ), .a(d1_o) );
    aoi222_1 \c1/__tmp99/U1  ( .x(d1_o), .a(d1_i), .b(ack), .c(d1_i), .d(
        \c1/ob ), .e(ack), .f(\c1/ob ) );
    inv_1 \c0/Ui  ( .x(\c0/ob ), .a(d0_o) );
    aoi222_1 \c0/__tmp99/U1  ( .x(d0_o), .a(d0_i), .b(ack), .c(d0_i), .d(
        \c0/ob ), .e(ack), .f(\c0/ob ) );
    latn_1 \slAck/lph3  ( .q(ack_l), .d(\slAck/l1_q ), .g(phi3) );
    latn_1 \slAck/lph2  ( .q(test_so), .d(\slAck/l1_q ), .g(phi2) );
    mux2_1 \slAck/mxl/mux  ( .x(\slAck/mxl/muxout ), .d0(ack_o), .sl(test_se), 
        .d1(test_si) );
    latn_1 \slAck/mxl/lph1  ( .q(\slAck/l1_q ), .d(\slAck/mxl/muxout ), .g(
        phi1) );
    or2_4 U7 ( .x(ack), .a(ack_l), .b(rst) );
endmodule


module chain_router10 ( eop_i, d0_i, d1_i, d2_i, d3_i, ack_i, eop_ox, d0_ox, 
    d1_ox, d2_ox, d3_ox, ack_ox, eop_oy, d0_oy, d1_oy, d2_oy, d3_oy, ack_oy, 
    nrst, test_si, test_se, test_so, phi1, phi2, phi3 );
input  eop_i, d0_i, d1_i, d2_i, d3_i, ack_ox, ack_oy, nrst, test_si, test_se, 
    phi1, phi2, phi3;
output ack_i, eop_ox, d0_ox, d1_ox, d2_ox, d3_ox, eop_oy, d0_oy, d1_oy, d2_oy, 
    d3_oy, test_so;
    wire rst, nack_x, ackx_l, nack_y, acky_l, n10, n11, n12, neopxy, n1, n2, 
        n3, n4, n5, n6, n7, n8, nrouteAckx, nrouteAcky, nroutex, nroutey, qa, 
        nqx, nqy, sx_pl, qx, sy_pl, qy, routeAcky, \cy/__tmp99/nr , qa_l, 
        \cy/__tmp99/nd , routeAckx, \cx/__tmp99/nr , \cx/__tmp99/nd , \cye/nr , 
        sy, \cye/nd , \cye/n2 , \cy3/__tmp99/loop , \cy2/__tmp99/loop , 
        \cy1/__tmp99/loop , \cy0/__tmp99/loop , \cxe/nr , sx, \cxe/nd , 
        \cxe/n2 , \cx3/__tmp99/loop , \cx2/__tmp99/loop , \cx1/__tmp99/loop , 
        \cx0/__tmp99/loop , \sl_sy/l1_q , \scan[2] , \sl_sy/mxl/muxout , 
        \scan[1] , \sl_sx/l1_q , \sl_sx/mxl/muxout , \scan[0] , \sl_qa/l1_q , 
        \sl_qa/mxl/muxout , \slAcky/l1_q , \slAcky/mxl/muxout , \scan[3] , 
        \slAckx/l1_q , \slAckx/mxl/muxout ;
    inv_1 U0 ( .x(rst), .a(nrst) );
    nor2_2 U5 ( .x(nack_x), .a(ackx_l), .b(rst) );
    nor2_2 U4 ( .x(nack_y), .a(acky_l), .b(rst) );
    nand4_1 U1 ( .x(ack_i), .a(n10), .b(n11), .c(n12), .d(neopxy) );
    and4_1 U8 ( .x(n10), .a(n1), .b(n2), .c(n3), .d(n4) );
    inv_1 U10 ( .x(n1), .a(d0_oy) );
    inv_1 U11 ( .x(n2), .a(d1_oy) );
    inv_1 U14 ( .x(n3), .a(d2_oy) );
    inv_1 U16 ( .x(n4), .a(d3_oy) );
    and4_1 U9 ( .x(n11), .a(n5), .b(n6), .c(n7), .d(n8) );
    inv_1 U17 ( .x(n5), .a(d0_ox) );
    inv_1 U18 ( .x(n6), .a(d1_ox) );
    inv_1 U19 ( .x(n7), .a(d2_ox) );
    inv_1 U20 ( .x(n8), .a(d3_ox) );
    nor2_1 U7 ( .x(n12), .a(nrouteAckx), .b(nrouteAcky) );
    nor2_1 U6 ( .x(neopxy), .a(eop_oy), .b(eop_ox) );
    nor2_1 U3 ( .x(nroutex), .a(d3_i), .b(d1_i) );
    nor2_1 U2 ( .x(nroutey), .a(d2_i), .b(d0_i) );
    nand2_1 U12 ( .x(qa), .a(nqx), .b(nqy) );
    nor2i_1 U15 ( .x(sx_pl), .a(qx), .b(nrouteAckx) );
    nor2i_1 U13 ( .x(sy_pl), .a(qy), .b(nrouteAcky) );
    inv_1 \cy/U1  ( .x(nrouteAcky), .a(routeAcky) );
    nor2_1 \cy/__tmp99/U1  ( .x(\cy/__tmp99/nr ), .a(nroutey), .b(qa_l) );
    nand2_1 \cy/__tmp99/U2  ( .x(\cy/__tmp99/nd ), .a(nroutey), .b(qa_l) );
    oai211_1 \cy/__tmp99/U3  ( .x(routeAcky), .a(nrouteAcky), .b(
        \cy/__tmp99/nr ), .c(\cy/__tmp99/nd ), .d(nrst) );
    inv_1 \cx/U1  ( .x(nrouteAckx), .a(routeAckx) );
    nor2_1 \cx/__tmp99/U1  ( .x(\cx/__tmp99/nr ), .a(nroutex), .b(qa_l) );
    nand2_1 \cx/__tmp99/U2  ( .x(\cx/__tmp99/nd ), .a(nroutex), .b(qa_l) );
    oai211_1 \cx/__tmp99/U3  ( .x(routeAckx), .a(nrouteAckx), .b(
        \cx/__tmp99/nr ), .c(\cx/__tmp99/nd ), .d(nrst) );
    nor3_1 \cye/Unr  ( .x(\cye/nr ), .a(eop_i), .b(nack_y), .c(sy) );
    nand3_1 \cye/Und  ( .x(\cye/nd ), .a(eop_i), .b(nack_y), .c(sy) );
    oa21_1 \cye/U1  ( .x(\cye/n2 ), .a(\cye/n2 ), .b(\cye/nr ), .c(\cye/nd )
         );
    inv_1 \cye/U3  ( .x(eop_oy), .a(\cye/n2 ) );
    ao31_1 \cy3/__tmp99/aoi  ( .x(\cy3/__tmp99/loop ), .a(d3_i), .b(nack_y), 
        .c(sy), .d(d3_oy) );
    ao31_1 \cy2/__tmp99/aoi  ( .x(\cy2/__tmp99/loop ), .a(d2_i), .b(nack_y), 
        .c(sy), .d(d2_oy) );
    ao31_1 \cy1/__tmp99/aoi  ( .x(\cy1/__tmp99/loop ), .a(d1_i), .b(nack_y), 
        .c(sy), .d(d1_oy) );
    ao31_1 \cy0/__tmp99/aoi  ( .x(\cy0/__tmp99/loop ), .a(d0_i), .b(nack_y), 
        .c(sy), .d(d0_oy) );
    nor3_1 \cxe/Unr  ( .x(\cxe/nr ), .a(eop_i), .b(nack_x), .c(sx) );
    nand3_1 \cxe/Und  ( .x(\cxe/nd ), .a(eop_i), .b(nack_x), .c(sx) );
    oa21_1 \cxe/U1  ( .x(\cxe/n2 ), .a(\cxe/n2 ), .b(\cxe/nr ), .c(\cxe/nd )
         );
    inv_1 \cxe/U3  ( .x(eop_ox), .a(\cxe/n2 ) );
    ao31_1 \cx3/__tmp99/aoi  ( .x(\cx3/__tmp99/loop ), .a(d3_i), .b(nack_x), 
        .c(sx), .d(d3_ox) );
    oa21_1 \cx3/__tmp99/outGate  ( .x(d3_ox), .a(d3_i), .b(nack_x), .c(
        \cx3/__tmp99/loop ) );
    ao31_1 \cx2/__tmp99/aoi  ( .x(\cx2/__tmp99/loop ), .a(d2_i), .b(nack_x), 
        .c(sx), .d(d2_ox) );
    oa21_1 \cx2/__tmp99/outGate  ( .x(d2_ox), .a(d2_i), .b(nack_x), .c(
        \cx2/__tmp99/loop ) );
    ao31_1 \cx1/__tmp99/aoi  ( .x(\cx1/__tmp99/loop ), .a(d1_i), .b(nack_x), 
        .c(sx), .d(d1_ox) );
    oa21_1 \cx1/__tmp99/outGate  ( .x(d1_ox), .a(d1_i), .b(nack_x), .c(
        \cx1/__tmp99/loop ) );
    ao31_1 \cx0/__tmp99/aoi  ( .x(\cx0/__tmp99/loop ), .a(d0_i), .b(nack_x), 
        .c(sx), .d(d0_ox) );
    oa21_1 \cx0/__tmp99/outGate  ( .x(d0_ox), .a(d0_i), .b(nack_x), .c(
        \cx0/__tmp99/loop ) );
    nand3_1 \sry/i0  ( .x(nqy), .a(neopxy), .b(nrst), .c(qy) );
    nand2_1 \sry/i1  ( .x(qy), .a(routeAcky), .b(nqy) );
    nand3_1 \srx/i0  ( .x(nqx), .a(neopxy), .b(nrst), .c(qx) );
    nand2_1 \srx/i1  ( .x(qx), .a(routeAckx), .b(nqx) );
    latn_1 \sl_sy/lph3  ( .q(sy), .d(\sl_sy/l1_q ), .g(phi3) );
    latn_1 \sl_sy/lph2  ( .q(\scan[2] ), .d(\sl_sy/l1_q ), .g(phi2) );
    mux2_1 \sl_sy/mxl/mux  ( .x(\sl_sy/mxl/muxout ), .d0(sy_pl), .sl(test_se), 
        .d1(\scan[1] ) );
    latn_1 \sl_sy/mxl/lph1  ( .q(\sl_sy/l1_q ), .d(\sl_sy/mxl/muxout ), .g(
        phi1) );
    latn_1 \sl_sx/lph3  ( .q(sx), .d(\sl_sx/l1_q ), .g(phi3) );
    latn_1 \sl_sx/lph2  ( .q(\scan[1] ), .d(\sl_sx/l1_q ), .g(phi2) );
    mux2_1 \sl_sx/mxl/mux  ( .x(\sl_sx/mxl/muxout ), .d0(sx_pl), .sl(test_se), 
        .d1(\scan[0] ) );
    latn_1 \sl_sx/mxl/lph1  ( .q(\sl_sx/l1_q ), .d(\sl_sx/mxl/muxout ), .g(
        phi1) );
    latn_1 \sl_qa/lph3  ( .q(qa_l), .d(\sl_qa/l1_q ), .g(phi3) );
    latn_1 \sl_qa/lph2  ( .q(\scan[0] ), .d(\sl_qa/l1_q ), .g(phi2) );
    mux2_1 \sl_qa/mxl/mux  ( .x(\sl_qa/mxl/muxout ), .d0(qa), .sl(test_se), 
        .d1(test_si) );
    latn_1 \sl_qa/mxl/lph1  ( .q(\sl_qa/l1_q ), .d(\sl_qa/mxl/muxout ), .g(
        phi1) );
    latn_1 \slAcky/lph3  ( .q(acky_l), .d(\slAcky/l1_q ), .g(phi3) );
    latn_1 \slAcky/lph2  ( .q(test_so), .d(\slAcky/l1_q ), .g(phi2) );
    mux2_1 \slAcky/mxl/mux  ( .x(\slAcky/mxl/muxout ), .d0(ack_oy), .sl(
        test_se), .d1(\scan[3] ) );
    latn_1 \slAcky/mxl/lph1  ( .q(\slAcky/l1_q ), .d(\slAcky/mxl/muxout ), .g(
        phi1) );
    latn_1 \slAckx/lph3  ( .q(ackx_l), .d(\slAckx/l1_q ), .g(phi3) );
    latn_1 \slAckx/lph2  ( .q(\scan[3] ), .d(\slAckx/l1_q ), .g(phi2) );
    mux2_1 \slAckx/mxl/mux  ( .x(\slAckx/mxl/muxout ), .d0(ack_ox), .sl(
        test_se), .d1(\scan[2] ) );
    latn_1 \slAckx/mxl/lph1  ( .q(\slAckx/l1_q ), .d(\slAckx/mxl/muxout ), .g(
        phi1) );
    oa21_2 U21 ( .x(d1_oy), .a(d1_i), .b(nack_y), .c(\cy1/__tmp99/loop ) );
    oa21_2 U22 ( .x(d2_oy), .a(d2_i), .b(nack_y), .c(\cy2/__tmp99/loop ) );
    oa21_2 U23 ( .x(d0_oy), .a(d0_i), .b(nack_y), .c(\cy0/__tmp99/loop ) );
    oa21_2 U24 ( .x(d3_oy), .a(d3_i), .b(nack_y), .c(\cy3/__tmp99/loop ) );
endmodule


module chain_router11 ( eop_i, d0_i, d1_i, d2_i, d3_i, ack_i, eop_ox, d0_ox, 
    d1_ox, d2_ox, d3_ox, ack_ox, eop_oy, d0_oy, d1_oy, d2_oy, d3_oy, ack_oy, 
    nrst, test_si, test_se, test_so, phi1, phi2, phi3 );
input  eop_i, d0_i, d1_i, d2_i, d3_i, ack_ox, ack_oy, nrst, test_si, test_se, 
    phi1, phi2, phi3;
output ack_i, eop_ox, d0_ox, d1_ox, d2_ox, d3_ox, eop_oy, d0_oy, d1_oy, d2_oy, 
    d3_oy, test_so;
    wire rst, nack_x, ackx_l, nack_y, acky_l, n10, n11, n12, neopxy, n1, n2, 
        n3, n4, n5, n6, n7, n8, nrouteAckx, nrouteAcky, nroutex, nroutey, qa, 
        nqx, nqy, sx_pl, qx, sy_pl, qy, routeAcky, \cy/__tmp99/nr , qa_l, 
        \cy/__tmp99/nd , routeAckx, \cx/__tmp99/nr , \cx/__tmp99/nd , \cye/nr , 
        sy, \cye/nd , \cye/n2 , \cy3/__tmp99/loop , \cy2/__tmp99/loop , 
        \cy1/__tmp99/loop , \cy0/__tmp99/loop , \cxe/nr , sx, \cxe/nd , 
        \cxe/n2 , \cx3/__tmp99/loop , \cx2/__tmp99/loop , \cx1/__tmp99/loop , 
        \cx0/__tmp99/loop , \sl_sy/l1_q , \scan[2] , \sl_sy/mxl/muxout , 
        \scan[1] , \sl_sx/l1_q , \sl_sx/mxl/muxout , \scan[0] , \sl_qa/l1_q , 
        \sl_qa/mxl/muxout , \slAcky/l1_q , \slAcky/mxl/muxout , \scan[3] , 
        \slAckx/l1_q , \slAckx/mxl/muxout ;
    inv_1 U0 ( .x(rst), .a(nrst) );
    nor2_2 U5 ( .x(nack_x), .a(ackx_l), .b(rst) );
    nor2_2 U4 ( .x(nack_y), .a(acky_l), .b(rst) );
    nand4_1 U1 ( .x(ack_i), .a(n10), .b(n11), .c(n12), .d(neopxy) );
    and4_1 U8 ( .x(n10), .a(n1), .b(n2), .c(n3), .d(n4) );
    inv_1 U10 ( .x(n1), .a(d0_oy) );
    inv_1 U11 ( .x(n2), .a(d1_oy) );
    inv_1 U14 ( .x(n3), .a(d2_oy) );
    inv_1 U16 ( .x(n4), .a(d3_oy) );
    and4_1 U9 ( .x(n11), .a(n5), .b(n6), .c(n7), .d(n8) );
    inv_1 U17 ( .x(n5), .a(d0_ox) );
    inv_1 U18 ( .x(n6), .a(d1_ox) );
    inv_1 U19 ( .x(n7), .a(d2_ox) );
    inv_1 U20 ( .x(n8), .a(d3_ox) );
    nor2_1 U7 ( .x(n12), .a(nrouteAckx), .b(nrouteAcky) );
    nor2_1 U6 ( .x(neopxy), .a(eop_oy), .b(eop_ox) );
    nor2_1 U3 ( .x(nroutex), .a(d3_i), .b(d1_i) );
    nor2_1 U2 ( .x(nroutey), .a(d2_i), .b(d0_i) );
    nand2_1 U12 ( .x(qa), .a(nqx), .b(nqy) );
    nor2i_1 U15 ( .x(sx_pl), .a(qx), .b(nrouteAckx) );
    nor2i_1 U13 ( .x(sy_pl), .a(qy), .b(nrouteAcky) );
    inv_1 \cy/U1  ( .x(nrouteAcky), .a(routeAcky) );
    nor2_1 \cy/__tmp99/U1  ( .x(\cy/__tmp99/nr ), .a(nroutey), .b(qa_l) );
    nand2_1 \cy/__tmp99/U2  ( .x(\cy/__tmp99/nd ), .a(nroutey), .b(qa_l) );
    oai211_1 \cy/__tmp99/U3  ( .x(routeAcky), .a(nrouteAcky), .b(
        \cy/__tmp99/nr ), .c(\cy/__tmp99/nd ), .d(nrst) );
    inv_1 \cx/U1  ( .x(nrouteAckx), .a(routeAckx) );
    nor2_1 \cx/__tmp99/U1  ( .x(\cx/__tmp99/nr ), .a(nroutex), .b(qa_l) );
    nand2_1 \cx/__tmp99/U2  ( .x(\cx/__tmp99/nd ), .a(nroutex), .b(qa_l) );
    oai211_1 \cx/__tmp99/U3  ( .x(routeAckx), .a(nrouteAckx), .b(
        \cx/__tmp99/nr ), .c(\cx/__tmp99/nd ), .d(nrst) );
    nor3_1 \cye/Unr  ( .x(\cye/nr ), .a(eop_i), .b(nack_y), .c(sy) );
    nand3_1 \cye/Und  ( .x(\cye/nd ), .a(eop_i), .b(nack_y), .c(sy) );
    oa21_1 \cye/U1  ( .x(\cye/n2 ), .a(\cye/n2 ), .b(\cye/nr ), .c(\cye/nd )
         );
    inv_1 \cye/U3  ( .x(eop_oy), .a(\cye/n2 ) );
    ao31_1 \cy3/__tmp99/aoi  ( .x(\cy3/__tmp99/loop ), .a(d3_i), .b(nack_y), 
        .c(sy), .d(d3_oy) );
    ao31_1 \cy2/__tmp99/aoi  ( .x(\cy2/__tmp99/loop ), .a(d2_i), .b(nack_y), 
        .c(sy), .d(d2_oy) );
    ao31_1 \cy1/__tmp99/aoi  ( .x(\cy1/__tmp99/loop ), .a(d1_i), .b(nack_y), 
        .c(sy), .d(d1_oy) );
    ao31_1 \cy0/__tmp99/aoi  ( .x(\cy0/__tmp99/loop ), .a(d0_i), .b(nack_y), 
        .c(sy), .d(d0_oy) );
    nor3_1 \cxe/Unr  ( .x(\cxe/nr ), .a(eop_i), .b(nack_x), .c(sx) );
    nand3_1 \cxe/Und  ( .x(\cxe/nd ), .a(eop_i), .b(nack_x), .c(sx) );
    oa21_1 \cxe/U1  ( .x(\cxe/n2 ), .a(\cxe/n2 ), .b(\cxe/nr ), .c(\cxe/nd )
         );
    inv_1 \cxe/U3  ( .x(eop_ox), .a(\cxe/n2 ) );
    ao31_1 \cx3/__tmp99/aoi  ( .x(\cx3/__tmp99/loop ), .a(d3_i), .b(nack_x), 
        .c(sx), .d(d3_ox) );
    ao31_1 \cx2/__tmp99/aoi  ( .x(\cx2/__tmp99/loop ), .a(d2_i), .b(nack_x), 
        .c(sx), .d(d2_ox) );
    ao31_1 \cx1/__tmp99/aoi  ( .x(\cx1/__tmp99/loop ), .a(d1_i), .b(nack_x), 
        .c(sx), .d(d1_ox) );
    ao31_1 \cx0/__tmp99/aoi  ( .x(\cx0/__tmp99/loop ), .a(d0_i), .b(nack_x), 
        .c(sx), .d(d0_ox) );
    nand3_1 \sry/i0  ( .x(nqy), .a(neopxy), .b(nrst), .c(qy) );
    nand2_1 \sry/i1  ( .x(qy), .a(routeAcky), .b(nqy) );
    nand3_1 \srx/i0  ( .x(nqx), .a(neopxy), .b(nrst), .c(qx) );
    nand2_1 \srx/i1  ( .x(qx), .a(routeAckx), .b(nqx) );
    latn_1 \sl_sy/lph3  ( .q(sy), .d(\sl_sy/l1_q ), .g(phi3) );
    latn_1 \sl_sy/lph2  ( .q(\scan[2] ), .d(\sl_sy/l1_q ), .g(phi2) );
    mux2_1 \sl_sy/mxl/mux  ( .x(\sl_sy/mxl/muxout ), .d0(sy_pl), .sl(test_se), 
        .d1(\scan[1] ) );
    latn_1 \sl_sy/mxl/lph1  ( .q(\sl_sy/l1_q ), .d(\sl_sy/mxl/muxout ), .g(
        phi1) );
    latn_1 \sl_sx/lph3  ( .q(sx), .d(\sl_sx/l1_q ), .g(phi3) );
    latn_1 \sl_sx/lph2  ( .q(\scan[1] ), .d(\sl_sx/l1_q ), .g(phi2) );
    mux2_1 \sl_sx/mxl/mux  ( .x(\sl_sx/mxl/muxout ), .d0(sx_pl), .sl(test_se), 
        .d1(\scan[0] ) );
    latn_1 \sl_sx/mxl/lph1  ( .q(\sl_sx/l1_q ), .d(\sl_sx/mxl/muxout ), .g(
        phi1) );
    latn_1 \sl_qa/lph3  ( .q(qa_l), .d(\sl_qa/l1_q ), .g(phi3) );
    latn_1 \sl_qa/lph2  ( .q(\scan[0] ), .d(\sl_qa/l1_q ), .g(phi2) );
    mux2_1 \sl_qa/mxl/mux  ( .x(\sl_qa/mxl/muxout ), .d0(qa), .sl(test_se), 
        .d1(test_si) );
    latn_1 \sl_qa/mxl/lph1  ( .q(\sl_qa/l1_q ), .d(\sl_qa/mxl/muxout ), .g(
        phi1) );
    latn_1 \slAcky/lph3  ( .q(acky_l), .d(\slAcky/l1_q ), .g(phi3) );
    latn_1 \slAcky/lph2  ( .q(test_so), .d(\slAcky/l1_q ), .g(phi2) );
    mux2_1 \slAcky/mxl/mux  ( .x(\slAcky/mxl/muxout ), .d0(ack_oy), .sl(
        test_se), .d1(\scan[3] ) );
    latn_1 \slAcky/mxl/lph1  ( .q(\slAcky/l1_q ), .d(\slAcky/mxl/muxout ), .g(
        phi1) );
    latn_1 \slAckx/lph3  ( .q(ackx_l), .d(\slAckx/l1_q ), .g(phi3) );
    latn_1 \slAckx/lph2  ( .q(\scan[3] ), .d(\slAckx/l1_q ), .g(phi2) );
    mux2_1 \slAckx/mxl/mux  ( .x(\slAckx/mxl/muxout ), .d0(ack_ox), .sl(
        test_se), .d1(\scan[2] ) );
    latn_1 \slAckx/mxl/lph1  ( .q(\slAckx/l1_q ), .d(\slAckx/mxl/muxout ), .g(
        phi1) );
    oa21_2 U21 ( .x(d3_oy), .a(d3_i), .b(nack_y), .c(\cy3/__tmp99/loop ) );
    oa21_2 U22 ( .x(d2_oy), .a(d2_i), .b(nack_y), .c(\cy2/__tmp99/loop ) );
    oa21_2 U23 ( .x(d1_oy), .a(d1_i), .b(nack_y), .c(\cy1/__tmp99/loop ) );
    oa21_2 U24 ( .x(d0_ox), .a(d0_i), .b(nack_x), .c(\cx0/__tmp99/loop ) );
    oa21_2 U25 ( .x(d2_ox), .a(d2_i), .b(nack_x), .c(\cx2/__tmp99/loop ) );
    oa21_2 U26 ( .x(d3_ox), .a(d3_i), .b(nack_x), .c(\cx3/__tmp99/loop ) );
    oa21_2 U27 ( .x(d1_ox), .a(d1_i), .b(nack_x), .c(\cx1/__tmp99/loop ) );
    oa21_2 U28 ( .x(d0_oy), .a(d0_i), .b(nack_y), .c(\cy0/__tmp99/loop ) );
endmodule


module resp_fab ( nrst, IMEM_eop_i, IMEM_d0_i, IMEM_d1_i, IMEM_d2_i, IMEM_d3_i, 
    IMEM_ack, DMEM_eop_i, DMEM_d0_i, DMEM_d1_i, DMEM_d2_i, DMEM_d3_i, DMEM_ack, 
    WB_eop_i, WB_d0_i, WB_d1_i, WB_d2_i, WB_d3_i, WB_ack, BC_eop_i, BC_d0_i, 
    BC_d1_i, BC_d2_i, BC_d3_i, BC_ack, I_port_eop_i, I_port_d0_i, I_port_d1_i, 
    I_port_d2_i, I_port_d3_i, I_port_ack, TIC_eop_i, TIC_d0_i, TIC_d1_i, 
    TIC_d2_i, TIC_d3_i, TIC_ack, D_port_eop_i, D_port_d0_i, D_port_d1_i, 
    D_port_d2_i, D_port_d3_i, D_port_ack, test_si, test_so, test_se, phi1, 
    phi2, phi3 );
input  nrst, IMEM_eop_i, IMEM_d0_i, IMEM_d1_i, IMEM_d2_i, IMEM_d3_i, 
    DMEM_eop_i, DMEM_d0_i, DMEM_d1_i, DMEM_d2_i, DMEM_d3_i, WB_eop_i, WB_d0_i, 
    WB_d1_i, WB_d2_i, WB_d3_i, BC_eop_i, BC_d0_i, BC_d1_i, BC_d2_i, BC_d3_i, 
    I_port_ack, TIC_ack, D_port_ack, test_si, test_se, phi1, phi2, phi3;
output IMEM_ack, DMEM_ack, WB_ack, BC_ack, I_port_eop_i, I_port_d0_i, 
    I_port_d1_i, I_port_d2_i, I_port_d3_i, TIC_eop_i, TIC_d0_i, TIC_d1_i, 
    TIC_d2_i, TIC_d3_i, D_port_eop_i, D_port_d0_i, D_port_d1_i, D_port_d2_i, 
    D_port_d3_i, test_so;
    wire A10_eop_o0, A10_d0_o0, A10_d1_o0, A10_d2_o0, A10_d3_o0, A10_eop_o1, 
        A10_d0_o1, A10_d1_o1, A10_d2_o1, A10_d3_o1, A10_ack, rst, \scan[1] , 
        M10_eop, M10_d0, M10_d1, M10_d2, M10_d3, M10_ack, n4, \scan[2] , n2, 
        n1, n3, A11_eop_o0, A11_d0_o0, A11_d1_o0, A11_d2_o0, A11_d3_o0, 
        A11_eop_o1, A11_d0_o1, A11_d1_o1, A11_d2_o1, A11_d3_o1, A11_ack, 
        \scan[3] , M11_eop, M11_d0, M11_d1, M11_d2, M11_d3, M11_ack, \scan[4] , 
        A12_eop_o0, A12_d0_o0, A12_d1_o0, A12_d2_o0, A12_d3_o0, A12_eop_o1, 
        A12_d0_o1, A12_d1_o1, A12_d2_o1, A12_d3_o1, A12_ack, \scan[5] , 
        M12_eop, M12_d0, M12_d1, M12_d2, M12_d3, M12_ack, \scan[6] , 
        R10_odd_eop, R10_odd_d0, R10_odd_d1, R10_odd_d2, R10_odd_d3, 
        R10_odd_ack, \scan[7] ;
    chain_arbiter10 arb10 ( .eop_ix(IMEM_eop_i), .d0_ix(IMEM_d0_i), .d1_ix(
        IMEM_d1_i), .d2_ix(IMEM_d2_i), .d3_ix(IMEM_d3_i), .ack_ix(IMEM_ack), 
        .eop_iy(DMEM_eop_i), .d0_iy(DMEM_d0_i), .d1_iy(DMEM_d1_i), .d2_iy(
        DMEM_d2_i), .d3_iy(DMEM_d3_i), .ack_iy(DMEM_ack), .eop_ox(A10_eop_o0), 
        .d0_ox(A10_d0_o0), .d1_ox(A10_d1_o0), .d2_ox(A10_d2_o0), .d3_ox(
        A10_d3_o0), .eop_oy(A10_eop_o1), .d0_oy(A10_d0_o1), .d1_oy(A10_d1_o1), 
        .d2_oy(A10_d2_o1), .d3_oy(A10_d3_o1), .ack_oxy(A10_ack), .rst(rst), 
        .test_si(test_si), .test_se(test_se), .test_so(\scan[1] ), .phi1(phi1), 
        .phi2(phi2), .phi3(phi3) );
    chain_mux10 mux10 ( .eop_ix(A10_eop_o0), .d0_ix(A10_d0_o0), .d1_ix(
        A10_d1_o0), .d2_ix(A10_d2_o0), .d3_ix(A10_d3_o0), .ack_ixy(A10_ack), 
        .eop_iy(A10_eop_o1), .d0_iy(A10_d0_o1), .d1_iy(A10_d1_o1), .d2_iy(
        A10_d2_o1), .d3_iy(A10_d3_o1), .eop_o(M10_eop), .d0_o(M10_d0), .d1_o(
        M10_d1), .d2_o(M10_d2), .d3_o(M10_d3), .ack_o(M10_ack), .rst(rst), 
        .test_si(\scan[1] ), .test_se(n4), .test_so(\scan[2] ), .phi1(n2), 
        .phi2(n1), .phi3(n3) );
    chain_arbiter11 arb11 ( .eop_ix(M10_eop), .d0_ix(M10_d0), .d1_ix(M10_d1), 
        .d2_ix(M10_d2), .d3_ix(M10_d3), .ack_ix(M10_ack), .eop_iy(BC_eop_i), 
        .d0_iy(BC_d0_i), .d1_iy(BC_d1_i), .d2_iy(BC_d2_i), .d3_iy(BC_d3_i), 
        .ack_iy(BC_ack), .eop_ox(A11_eop_o0), .d0_ox(A11_d0_o0), .d1_ox(
        A11_d1_o0), .d2_ox(A11_d2_o0), .d3_ox(A11_d3_o0), .eop_oy(A11_eop_o1), 
        .d0_oy(A11_d0_o1), .d1_oy(A11_d1_o1), .d2_oy(A11_d2_o1), .d3_oy(
        A11_d3_o1), .ack_oxy(A11_ack), .rst(rst), .test_si(\scan[2] ), 
        .test_se(n4), .test_so(\scan[3] ), .phi1(n2), .phi2(n1), .phi3(n3) );
    chain_mux11 mux11 ( .eop_ix(A11_eop_o0), .d0_ix(A11_d0_o0), .d1_ix(
        A11_d1_o0), .d2_ix(A11_d2_o0), .d3_ix(A11_d3_o0), .ack_ixy(A11_ack), 
        .eop_iy(A11_eop_o1), .d0_iy(A11_d0_o1), .d1_iy(A11_d1_o1), .d2_iy(
        A11_d2_o1), .d3_iy(A11_d3_o1), .eop_o(M11_eop), .d0_o(M11_d0), .d1_o(
        M11_d1), .d2_o(M11_d2), .d3_o(M11_d3), .ack_o(M11_ack), .rst(rst), 
        .test_si(\scan[3] ), .test_se(test_se), .test_so(\scan[4] ), .phi1(
        phi1), .phi2(phi2), .phi3(phi3) );
    chain_arbiter12 arb12 ( .eop_ix(M11_eop), .d0_ix(M11_d0), .d1_ix(M11_d1), 
        .d2_ix(M11_d2), .d3_ix(M11_d3), .ack_ix(M11_ack), .eop_iy(WB_eop_i), 
        .d0_iy(WB_d0_i), .d1_iy(WB_d1_i), .d2_iy(WB_d2_i), .d3_iy(WB_d3_i), 
        .ack_iy(WB_ack), .eop_ox(A12_eop_o0), .d0_ox(A12_d0_o0), .d1_ox(
        A12_d1_o0), .d2_ox(A12_d2_o0), .d3_ox(A12_d3_o0), .eop_oy(A12_eop_o1), 
        .d0_oy(A12_d0_o1), .d1_oy(A12_d1_o1), .d2_oy(A12_d2_o1), .d3_oy(
        A12_d3_o1), .ack_oxy(A12_ack), .rst(rst), .test_si(\scan[4] ), 
        .test_se(n4), .test_so(\scan[5] ), .phi1(n2), .phi2(n1), .phi3(n3) );
    chain_mux12 mux12 ( .eop_ix(A12_eop_o0), .d0_ix(A12_d0_o0), .d1_ix(
        A12_d1_o0), .d2_ix(A12_d2_o0), .d3_ix(A12_d3_o0), .ack_ixy(A12_ack), 
        .eop_iy(A12_eop_o1), .d0_iy(A12_d0_o1), .d1_iy(A12_d1_o1), .d2_iy(
        A12_d2_o1), .d3_iy(A12_d3_o1), .eop_o(M12_eop), .d0_o(M12_d0), .d1_o(
        M12_d1), .d2_o(M12_d2), .d3_o(M12_d3), .ack_o(M12_ack), .rst(rst), 
        .test_si(\scan[5] ), .test_se(n4), .test_so(\scan[6] ), .phi1(n2), 
        .phi2(n1), .phi3(n3) );
    chain_router10 router10 ( .eop_i(M12_eop), .d0_i(M12_d0), .d1_i(M12_d1), 
        .d2_i(M12_d2), .d3_i(M12_d3), .ack_i(M12_ack), .eop_ox(R10_odd_eop), 
        .d0_ox(R10_odd_d0), .d1_ox(R10_odd_d1), .d2_ox(R10_odd_d2), .d3_ox(
        R10_odd_d3), .ack_ox(R10_odd_ack), .eop_oy(TIC_eop_i), .d0_oy(TIC_d0_i
        ), .d1_oy(TIC_d1_i), .d2_oy(TIC_d2_i), .d3_oy(TIC_d3_i), .ack_oy(
        TIC_ack), .nrst(nrst), .test_si(\scan[6] ), .test_se(n4), .test_so(
        \scan[7] ), .phi1(phi1), .phi2(phi2), .phi3(phi3) );
    chain_router11 router11 ( .eop_i(R10_odd_eop), .d0_i(R10_odd_d0), .d1_i(
        R10_odd_d1), .d2_i(R10_odd_d2), .d3_i(R10_odd_d3), .ack_i(R10_odd_ack), 
        .eop_ox(I_port_eop_i), .d0_ox(I_port_d0_i), .d1_ox(I_port_d1_i), 
        .d2_ox(I_port_d2_i), .d3_ox(I_port_d3_i), .ack_ox(I_port_ack), 
        .eop_oy(D_port_eop_i), .d0_oy(D_port_d0_i), .d1_oy(D_port_d1_i), 
        .d2_oy(D_port_d2_i), .d3_oy(D_port_d3_i), .ack_oy(D_port_ack), .nrst(
        nrst), .test_si(\scan[7] ), .test_se(test_se), .test_so(test_so), 
        .phi1(phi1), .phi2(phi2), .phi3(phi3) );
    buf_1 U1 ( .x(n1), .a(phi2) );
    buf_1 U2 ( .x(n2), .a(phi1) );
    buf_1 U3 ( .x(n3), .a(phi3) );
    buf_3 U4 ( .x(n4), .a(test_se) );
    inv_5 U5 ( .x(rst), .a(nrst) );
endmodule


module resp_fab_scan ( nrst, IMEM_eop_i, IMEM_d0_i, IMEM_d1_i, IMEM_d2_i, 
    IMEM_d3_i, IMEM_ack, DMEM_eop_i, DMEM_d0_i, DMEM_d1_i, DMEM_d2_i, 
    DMEM_d3_i, DMEM_ack, WB_eop_i, WB_d0_i, WB_d1_i, WB_d2_i, WB_d3_i, WB_ack, 
    BC_eop_i, BC_d0_i, BC_d1_i, BC_d2_i, BC_d3_i, BC_ack, I_port_eop_i, 
    I_port_d0_i, I_port_d1_i, I_port_d2_i, I_port_d3_i, I_port_ack, TIC_eop_i, 
    TIC_d0_i, TIC_d1_i, TIC_d2_i, TIC_d3_i, TIC_ack, D_port_eop_i, D_port_d0_i, 
    D_port_d1_i, D_port_d2_i, D_port_d3_i, D_port_ack, test_si, test_so, 
    test_se, phi1, phi2, phi3 );
input  nrst, IMEM_eop_i, IMEM_d0_i, IMEM_d1_i, IMEM_d2_i, IMEM_d3_i, 
    DMEM_eop_i, DMEM_d0_i, DMEM_d1_i, DMEM_d2_i, DMEM_d3_i, WB_eop_i, WB_d0_i, 
    WB_d1_i, WB_d2_i, WB_d3_i, BC_eop_i, BC_d0_i, BC_d1_i, BC_d2_i, BC_d3_i, 
    I_port_ack, TIC_ack, D_port_ack, test_si, test_se, phi1, phi2, phi3;
output IMEM_ack, DMEM_ack, WB_ack, BC_ack, I_port_eop_i, I_port_d0_i, 
    I_port_d1_i, I_port_d2_i, I_port_d3_i, TIC_eop_i, TIC_d0_i, TIC_d1_i, 
    TIC_d2_i, TIC_d3_i, D_port_eop_i, D_port_d0_i, D_port_d1_i, D_port_d2_i, 
    D_port_d3_i, test_so;
    wire IMEM_eop_i_sc, IMEM_d0_i_sc, IMEM_d1_i_sc, IMEM_d2_i_sc, IMEM_d3_i_sc, 
        DMEM_eop_i_sc, DMEM_d0_i_sc, DMEM_d1_i_sc, DMEM_d2_i_sc, DMEM_d3_i_sc, 
        WB_eop_i_sc, WB_d0_i_sc, WB_d1_i_sc, WB_d2_i_sc, WB_d3_i_sc, 
        I_port_ack_sc, TIC_ack_sc, D_port_ack_sc, \scan[6] , \scan[7] , n5, n9, 
        n13, n2, \scan[11] , scan_m10, n15, \scan[12] , scan_m11, n12, 
        scan_m12, n14, \sc12_m_wbAck/muxout , n7, n11, \sc11_m_dmAck/muxout , 
        n6, n8, \sc10_m_imAck/muxout , \scan[10] , n10, \sc6_dpAck/l1_q , n1, 
        \sc6_dpAck/mxl/muxout , \scan[5] , \sc5_ticAck/l1_q , 
        \sc5_ticAck/mxl/muxout , n4, \scan[4] , \sc4_ipAck/l1_q , 
        \sc4_ipAck/mxl/muxout , \scan[3] , \sc_dp/intI4 , \sc_dp/scn3 , 
        \sc_dp/intI3 , \sc_dp/scn2 , \sc_dp/intI2 , \sc_dp/scn1 , 
        \sc_dp/intI1 , \sc_dp/scn0 , \sc_dp/intI0 , \sc_dp/l4_m/muxout , 
        \sc_dp/l3_m/muxout , \sc_dp/l2_m/muxout , \sc_dp/l1_m/muxout , 
        \sc_dp/l0_m/muxout , \scan[9] , \sc_tic/intI4 , \sc_tic/scn3 , 
        \sc_tic/intI3 , \sc_tic/scn2 , \sc_tic/intI2 , \sc_tic/scn1 , 
        \sc_tic/intI1 , \sc_tic/scn0 , \sc_tic/intI0 , \sc_tic/l4_m/muxout , 
        \sc_tic/l3_m/muxout , \sc_tic/l2_m/muxout , \sc_tic/l1_m/muxout , 
        \sc_tic/l0_m/muxout , \scan[8] , \sc_ip/intI4 , \sc_ip/scn3 , 
        \sc_ip/intI3 , \sc_ip/scn2 , \sc_ip/intI2 , \sc_ip/scn1 , 
        \sc_ip/intI1 , \sc_ip/scn0 , \sc_ip/intI0 , \sc_ip/l4_m/muxout , 
        \sc_ip/l3_m/muxout , \sc_ip/l2_m/muxout , \sc_ip/l1_m/muxout , 
        \sc_ip/l0_m/muxout , \sc_wb/sl4/l1_q , n3, \sc_wb/sl4/mxl/muxout , 
        \sc_wb/scn4 , \sc_wb/sl3/l1_q , \sc_wb/sl3/mxl/muxout , \sc_wb/scn3 , 
        \sc_wb/sl2/l1_q , \sc_wb/sl2/mxl/muxout , \sc_wb/scn2 , 
        \sc_wb/sl1/l1_q , \sc_wb/sl1/mxl/muxout , \sc_wb/scn1 , 
        \sc_wb/sl0/l1_q , \sc_wb/sl0/mxl/muxout , \scan[2] , \sc_dm/sl4/l1_q , 
        \sc_dm/sl4/mxl/muxout , \sc_dm/scn4 , \sc_dm/sl3/l1_q , 
        \sc_dm/sl3/mxl/muxout , \sc_dm/scn3 , \sc_dm/sl2/l1_q , 
        \sc_dm/sl2/mxl/muxout , \sc_dm/scn2 , \sc_dm/sl1/l1_q , 
        \sc_dm/sl1/mxl/muxout , \sc_dm/scn1 , \sc_dm/sl0/l1_q , 
        \sc_dm/sl0/mxl/muxout , \scan[1] , \sc_im/sl4/l1_q , 
        \sc_im/sl4/mxl/muxout , \sc_im/scn4 , \sc_im/sl3/l1_q , 
        \sc_im/sl3/mxl/muxout , \sc_im/scn3 , \sc_im/sl2/l1_q , 
        \sc_im/sl2/mxl/muxout , \sc_im/scn2 , \sc_im/sl1/l1_q , 
        \sc_im/sl1/mxl/muxout , \sc_im/scn1 , \sc_im/sl0/l1_q , 
        \sc_im/sl0/mxl/muxout ;
    resp_fab fab2 ( .nrst(nrst), .IMEM_eop_i(IMEM_eop_i_sc), .IMEM_d0_i(
        IMEM_d0_i_sc), .IMEM_d1_i(IMEM_d1_i_sc), .IMEM_d2_i(IMEM_d2_i_sc), 
        .IMEM_d3_i(IMEM_d3_i_sc), .IMEM_ack(IMEM_ack), .DMEM_eop_i(
        DMEM_eop_i_sc), .DMEM_d0_i(DMEM_d0_i_sc), .DMEM_d1_i(DMEM_d1_i_sc), 
        .DMEM_d2_i(DMEM_d2_i_sc), .DMEM_d3_i(DMEM_d3_i_sc), .DMEM_ack(DMEM_ack
        ), .WB_eop_i(WB_eop_i_sc), .WB_d0_i(WB_d0_i_sc), .WB_d1_i(WB_d1_i_sc), 
        .WB_d2_i(WB_d2_i_sc), .WB_d3_i(WB_d3_i_sc), .WB_ack(WB_ack), 
        .BC_eop_i(BC_eop_i), .BC_d0_i(BC_d0_i), .BC_d1_i(BC_d1_i), .BC_d2_i(
        BC_d2_i), .BC_d3_i(BC_d3_i), .BC_ack(BC_ack), .I_port_eop_i(
        I_port_eop_i), .I_port_d0_i(I_port_d0_i), .I_port_d1_i(I_port_d1_i), 
        .I_port_d2_i(I_port_d2_i), .I_port_d3_i(I_port_d3_i), .I_port_ack(
        I_port_ack_sc), .TIC_eop_i(TIC_eop_i), .TIC_d0_i(TIC_d0_i), .TIC_d1_i(
        TIC_d1_i), .TIC_d2_i(TIC_d2_i), .TIC_d3_i(TIC_d3_i), .TIC_ack(
        TIC_ack_sc), .D_port_eop_i(D_port_eop_i), .D_port_d0_i(D_port_d0_i), 
        .D_port_d1_i(D_port_d1_i), .D_port_d2_i(D_port_d2_i), .D_port_d3_i(
        D_port_d3_i), .D_port_ack(D_port_ack_sc), .test_si(\scan[6] ), 
        .test_so(\scan[7] ), .test_se(n5), .phi1(n9), .phi2(n13), .phi3(n2) );
    latn_1 sc10_s_imAck ( .q(\scan[11] ), .d(scan_m10), .g(n15) );
    latn_1 sc11_s_dmAck ( .q(\scan[12] ), .d(scan_m11), .g(n12) );
    latn_1 sc12_s_wbAck ( .q(test_so), .d(scan_m12), .g(n14) );
    mux2_1 \sc12_m_wbAck/mux  ( .x(\sc12_m_wbAck/muxout ), .d0(WB_ack), .sl(n7
        ), .d1(\scan[12] ) );
    latn_1 \sc12_m_wbAck/lph1  ( .q(scan_m12), .d(\sc12_m_wbAck/muxout ), .g(
        n11) );
    mux2_1 \sc11_m_dmAck/mux  ( .x(\sc11_m_dmAck/muxout ), .d0(DMEM_ack), .sl(
        n6), .d1(\scan[11] ) );
    latn_1 \sc11_m_dmAck/lph1  ( .q(scan_m11), .d(\sc11_m_dmAck/muxout ), .g(
        n8) );
    mux2_1 \sc10_m_imAck/mux  ( .x(\sc10_m_imAck/muxout ), .d0(IMEM_ack), .sl(
        n6), .d1(\scan[10] ) );
    latn_1 \sc10_m_imAck/lph1  ( .q(scan_m10), .d(\sc10_m_imAck/muxout ), .g(
        n10) );
    latn_1 \sc6_dpAck/lph3  ( .q(D_port_ack_sc), .d(\sc6_dpAck/l1_q ), .g(n1)
         );
    latn_1 \sc6_dpAck/lph2  ( .q(\scan[6] ), .d(\sc6_dpAck/l1_q ), .g(n15) );
    mux2_1 \sc6_dpAck/mxl/mux  ( .x(\sc6_dpAck/mxl/muxout ), .d0(D_port_ack), 
        .sl(n7), .d1(\scan[5] ) );
    latn_1 \sc6_dpAck/mxl/lph1  ( .q(\sc6_dpAck/l1_q ), .d(
        \sc6_dpAck/mxl/muxout ), .g(n10) );
    latn_1 \sc5_ticAck/lph3  ( .q(TIC_ack_sc), .d(\sc5_ticAck/l1_q ), .g(n1)
         );
    latn_1 \sc5_ticAck/lph2  ( .q(\scan[5] ), .d(\sc5_ticAck/l1_q ), .g(n12)
         );
    mux2_1 \sc5_ticAck/mxl/mux  ( .x(\sc5_ticAck/mxl/muxout ), .d0(TIC_ack), 
        .sl(n4), .d1(\scan[4] ) );
    latn_1 \sc5_ticAck/mxl/lph1  ( .q(\sc5_ticAck/l1_q ), .d(
        \sc5_ticAck/mxl/muxout ), .g(n8) );
    latn_1 \sc4_ipAck/lph3  ( .q(I_port_ack_sc), .d(\sc4_ipAck/l1_q ), .g(n1)
         );
    latn_1 \sc4_ipAck/lph2  ( .q(\scan[4] ), .d(\sc4_ipAck/l1_q ), .g(n14) );
    mux2_1 \sc4_ipAck/mxl/mux  ( .x(\sc4_ipAck/mxl/muxout ), .d0(I_port_ack), 
        .sl(n4), .d1(\scan[3] ) );
    latn_1 \sc4_ipAck/mxl/lph1  ( .q(\sc4_ipAck/l1_q ), .d(
        \sc4_ipAck/mxl/muxout ), .g(n11) );
    latn_1 \sc_dp/l4_s  ( .q(\scan[10] ), .d(\sc_dp/intI4 ), .g(n15) );
    latn_1 \sc_dp/l3_s  ( .q(\sc_dp/scn3 ), .d(\sc_dp/intI3 ), .g(n12) );
    latn_1 \sc_dp/l2_s  ( .q(\sc_dp/scn2 ), .d(\sc_dp/intI2 ), .g(n14) );
    latn_1 \sc_dp/l1_s  ( .q(\sc_dp/scn1 ), .d(\sc_dp/intI1 ), .g(n15) );
    latn_1 \sc_dp/l0_s  ( .q(\sc_dp/scn0 ), .d(\sc_dp/intI0 ), .g(n12) );
    mux2_1 \sc_dp/l4_m/mux  ( .x(\sc_dp/l4_m/muxout ), .d0(D_port_d3_i), .sl(
        n4), .d1(\sc_dp/scn3 ) );
    latn_1 \sc_dp/l4_m/lph1  ( .q(\sc_dp/intI4 ), .d(\sc_dp/l4_m/muxout ), .g(
        n8) );
    mux2_1 \sc_dp/l3_m/mux  ( .x(\sc_dp/l3_m/muxout ), .d0(D_port_d2_i), .sl(
        n7), .d1(\sc_dp/scn2 ) );
    latn_1 \sc_dp/l3_m/lph1  ( .q(\sc_dp/intI3 ), .d(\sc_dp/l3_m/muxout ), .g(
        n11) );
    mux2_1 \sc_dp/l2_m/mux  ( .x(\sc_dp/l2_m/muxout ), .d0(D_port_d1_i), .sl(
        n6), .d1(\sc_dp/scn1 ) );
    latn_1 \sc_dp/l2_m/lph1  ( .q(\sc_dp/intI2 ), .d(\sc_dp/l2_m/muxout ), .g(
        n10) );
    mux2_1 \sc_dp/l1_m/mux  ( .x(\sc_dp/l1_m/muxout ), .d0(D_port_d0_i), .sl(
        n4), .d1(\sc_dp/scn0 ) );
    latn_1 \sc_dp/l1_m/lph1  ( .q(\sc_dp/intI1 ), .d(\sc_dp/l1_m/muxout ), .g(
        n8) );
    mux2_1 \sc_dp/l0_m/mux  ( .x(\sc_dp/l0_m/muxout ), .d0(D_port_eop_i), .sl(
        n7), .d1(\scan[9] ) );
    latn_1 \sc_dp/l0_m/lph1  ( .q(\sc_dp/intI0 ), .d(\sc_dp/l0_m/muxout ), .g(
        n11) );
    latn_1 \sc_tic/l4_s  ( .q(\scan[9] ), .d(\sc_tic/intI4 ), .g(n12) );
    latn_1 \sc_tic/l3_s  ( .q(\sc_tic/scn3 ), .d(\sc_tic/intI3 ), .g(n14) );
    latn_1 \sc_tic/l2_s  ( .q(\sc_tic/scn2 ), .d(\sc_tic/intI2 ), .g(n15) );
    latn_1 \sc_tic/l1_s  ( .q(\sc_tic/scn1 ), .d(\sc_tic/intI1 ), .g(n12) );
    latn_1 \sc_tic/l0_s  ( .q(\sc_tic/scn0 ), .d(\sc_tic/intI0 ), .g(n14) );
    mux2_1 \sc_tic/l4_m/mux  ( .x(\sc_tic/l4_m/muxout ), .d0(TIC_d3_i), .sl(n6
        ), .d1(\sc_tic/scn3 ) );
    latn_1 \sc_tic/l4_m/lph1  ( .q(\sc_tic/intI4 ), .d(\sc_tic/l4_m/muxout ), 
        .g(n10) );
    mux2_1 \sc_tic/l3_m/mux  ( .x(\sc_tic/l3_m/muxout ), .d0(TIC_d2_i), .sl(n4
        ), .d1(\sc_tic/scn2 ) );
    latn_1 \sc_tic/l3_m/lph1  ( .q(\sc_tic/intI3 ), .d(\sc_tic/l3_m/muxout ), 
        .g(n8) );
    mux2_1 \sc_tic/l2_m/mux  ( .x(\sc_tic/l2_m/muxout ), .d0(TIC_d1_i), .sl(n7
        ), .d1(\sc_tic/scn1 ) );
    latn_1 \sc_tic/l2_m/lph1  ( .q(\sc_tic/intI2 ), .d(\sc_tic/l2_m/muxout ), 
        .g(n11) );
    mux2_1 \sc_tic/l1_m/mux  ( .x(\sc_tic/l1_m/muxout ), .d0(TIC_d0_i), .sl(n6
        ), .d1(\sc_tic/scn0 ) );
    latn_1 \sc_tic/l1_m/lph1  ( .q(\sc_tic/intI1 ), .d(\sc_tic/l1_m/muxout ), 
        .g(n10) );
    mux2_1 \sc_tic/l0_m/mux  ( .x(\sc_tic/l0_m/muxout ), .d0(TIC_eop_i), .sl(
        n4), .d1(\scan[8] ) );
    latn_1 \sc_tic/l0_m/lph1  ( .q(\sc_tic/intI0 ), .d(\sc_tic/l0_m/muxout ), 
        .g(n8) );
    latn_1 \sc_ip/l4_s  ( .q(\scan[8] ), .d(\sc_ip/intI4 ), .g(n14) );
    latn_1 \sc_ip/l3_s  ( .q(\sc_ip/scn3 ), .d(\sc_ip/intI3 ), .g(n15) );
    latn_1 \sc_ip/l2_s  ( .q(\sc_ip/scn2 ), .d(\sc_ip/intI2 ), .g(n12) );
    latn_1 \sc_ip/l1_s  ( .q(\sc_ip/scn1 ), .d(\sc_ip/intI1 ), .g(n14) );
    latn_1 \sc_ip/l0_s  ( .q(\sc_ip/scn0 ), .d(\sc_ip/intI0 ), .g(n15) );
    mux2_1 \sc_ip/l4_m/mux  ( .x(\sc_ip/l4_m/muxout ), .d0(I_port_d3_i), .sl(
        n7), .d1(\sc_ip/scn3 ) );
    latn_1 \sc_ip/l4_m/lph1  ( .q(\sc_ip/intI4 ), .d(\sc_ip/l4_m/muxout ), .g(
        n11) );
    mux2_1 \sc_ip/l3_m/mux  ( .x(\sc_ip/l3_m/muxout ), .d0(I_port_d2_i), .sl(
        n7), .d1(\sc_ip/scn2 ) );
    latn_1 \sc_ip/l3_m/lph1  ( .q(\sc_ip/intI3 ), .d(\sc_ip/l3_m/muxout ), .g(
        n10) );
    mux2_1 \sc_ip/l2_m/mux  ( .x(\sc_ip/l2_m/muxout ), .d0(I_port_d1_i), .sl(
        n6), .d1(\sc_ip/scn1 ) );
    latn_1 \sc_ip/l2_m/lph1  ( .q(\sc_ip/intI2 ), .d(\sc_ip/l2_m/muxout ), .g(
        n8) );
    mux2_1 \sc_ip/l1_m/mux  ( .x(\sc_ip/l1_m/muxout ), .d0(I_port_d0_i), .sl(
        n4), .d1(\sc_ip/scn0 ) );
    latn_1 \sc_ip/l1_m/lph1  ( .q(\sc_ip/intI1 ), .d(\sc_ip/l1_m/muxout ), .g(
        n11) );
    mux2_1 \sc_ip/l0_m/mux  ( .x(\sc_ip/l0_m/muxout ), .d0(I_port_eop_i), .sl(
        n7), .d1(\scan[7] ) );
    latn_1 \sc_ip/l0_m/lph1  ( .q(\sc_ip/intI0 ), .d(\sc_ip/l0_m/muxout ), .g(
        n10) );
    latn_1 \sc_wb/sl4/lph3  ( .q(WB_d3_i_sc), .d(\sc_wb/sl4/l1_q ), .g(n3) );
    latn_1 \sc_wb/sl4/lph2  ( .q(\scan[3] ), .d(\sc_wb/sl4/l1_q ), .g(n12) );
    mux2_1 \sc_wb/sl4/mxl/mux  ( .x(\sc_wb/sl4/mxl/muxout ), .d0(WB_d3_i), 
        .sl(n6), .d1(\sc_wb/scn4 ) );
    latn_1 \sc_wb/sl4/mxl/lph1  ( .q(\sc_wb/sl4/l1_q ), .d(
        \sc_wb/sl4/mxl/muxout ), .g(n8) );
    latn_1 \sc_wb/sl3/lph3  ( .q(WB_d2_i_sc), .d(\sc_wb/sl3/l1_q ), .g(n3) );
    latn_1 \sc_wb/sl3/lph2  ( .q(\sc_wb/scn4 ), .d(\sc_wb/sl3/l1_q ), .g(n15)
         );
    mux2_1 \sc_wb/sl3/mxl/mux  ( .x(\sc_wb/sl3/mxl/muxout ), .d0(WB_d2_i), 
        .sl(n4), .d1(\sc_wb/scn3 ) );
    latn_1 \sc_wb/sl3/mxl/lph1  ( .q(\sc_wb/sl3/l1_q ), .d(
        \sc_wb/sl3/mxl/muxout ), .g(n11) );
    latn_1 \sc_wb/sl2/lph3  ( .q(WB_d1_i_sc), .d(\sc_wb/sl2/l1_q ), .g(n3) );
    latn_1 \sc_wb/sl2/lph2  ( .q(\sc_wb/scn3 ), .d(\sc_wb/sl2/l1_q ), .g(n14)
         );
    mux2_1 \sc_wb/sl2/mxl/mux  ( .x(\sc_wb/sl2/mxl/muxout ), .d0(WB_d1_i), 
        .sl(n7), .d1(\sc_wb/scn2 ) );
    latn_1 \sc_wb/sl2/mxl/lph1  ( .q(\sc_wb/sl2/l1_q ), .d(
        \sc_wb/sl2/mxl/muxout ), .g(n10) );
    latn_1 \sc_wb/sl1/lph3  ( .q(WB_d0_i_sc), .d(\sc_wb/sl1/l1_q ), .g(n3) );
    latn_1 \sc_wb/sl1/lph2  ( .q(\sc_wb/scn2 ), .d(\sc_wb/sl1/l1_q ), .g(n15)
         );
    mux2_1 \sc_wb/sl1/mxl/mux  ( .x(\sc_wb/sl1/mxl/muxout ), .d0(WB_d0_i), 
        .sl(n4), .d1(\sc_wb/scn1 ) );
    latn_1 \sc_wb/sl1/mxl/lph1  ( .q(\sc_wb/sl1/l1_q ), .d(
        \sc_wb/sl1/mxl/muxout ), .g(n11) );
    latn_1 \sc_wb/sl0/lph3  ( .q(WB_eop_i_sc), .d(\sc_wb/sl0/l1_q ), .g(n3) );
    latn_1 \sc_wb/sl0/lph2  ( .q(\sc_wb/scn1 ), .d(\sc_wb/sl0/l1_q ), .g(n12)
         );
    mux2_1 \sc_wb/sl0/mxl/mux  ( .x(\sc_wb/sl0/mxl/muxout ), .d0(WB_eop_i), 
        .sl(n4), .d1(\scan[2] ) );
    latn_1 \sc_wb/sl0/mxl/lph1  ( .q(\sc_wb/sl0/l1_q ), .d(
        \sc_wb/sl0/mxl/muxout ), .g(n8) );
    latn_1 \sc_dm/sl4/lph3  ( .q(DMEM_d3_i_sc), .d(\sc_dm/sl4/l1_q ), .g(n3)
         );
    latn_1 \sc_dm/sl4/lph2  ( .q(\scan[2] ), .d(\sc_dm/sl4/l1_q ), .g(n14) );
    mux2_1 \sc_dm/sl4/mxl/mux  ( .x(\sc_dm/sl4/mxl/muxout ), .d0(DMEM_d3_i), 
        .sl(n6), .d1(\sc_dm/scn4 ) );
    latn_1 \sc_dm/sl4/mxl/lph1  ( .q(\sc_dm/sl4/l1_q ), .d(
        \sc_dm/sl4/mxl/muxout ), .g(n10) );
    latn_1 \sc_dm/sl3/lph3  ( .q(DMEM_d2_i_sc), .d(\sc_dm/sl3/l1_q ), .g(n3)
         );
    latn_1 \sc_dm/sl3/lph2  ( .q(\sc_dm/scn4 ), .d(\sc_dm/sl3/l1_q ), .g(n15)
         );
    mux2_1 \sc_dm/sl3/mxl/mux  ( .x(\sc_dm/sl3/mxl/muxout ), .d0(DMEM_d2_i), 
        .sl(n7), .d1(\sc_dm/scn3 ) );
    latn_1 \sc_dm/sl3/mxl/lph1  ( .q(\sc_dm/sl3/l1_q ), .d(
        \sc_dm/sl3/mxl/muxout ), .g(n11) );
    latn_1 \sc_dm/sl2/lph3  ( .q(DMEM_d1_i_sc), .d(\sc_dm/sl2/l1_q ), .g(n3)
         );
    latn_1 \sc_dm/sl2/lph2  ( .q(\sc_dm/scn3 ), .d(\sc_dm/sl2/l1_q ), .g(n12)
         );
    mux2_1 \sc_dm/sl2/mxl/mux  ( .x(\sc_dm/sl2/mxl/muxout ), .d0(DMEM_d1_i), 
        .sl(n6), .d1(\sc_dm/scn2 ) );
    latn_1 \sc_dm/sl2/mxl/lph1  ( .q(\sc_dm/sl2/l1_q ), .d(
        \sc_dm/sl2/mxl/muxout ), .g(n8) );
    latn_1 \sc_dm/sl1/lph3  ( .q(DMEM_d0_i_sc), .d(\sc_dm/sl1/l1_q ), .g(n3)
         );
    latn_1 \sc_dm/sl1/lph2  ( .q(\sc_dm/scn2 ), .d(\sc_dm/sl1/l1_q ), .g(n15)
         );
    mux2_1 \sc_dm/sl1/mxl/mux  ( .x(\sc_dm/sl1/mxl/muxout ), .d0(DMEM_d0_i), 
        .sl(n7), .d1(\sc_dm/scn1 ) );
    latn_1 \sc_dm/sl1/mxl/lph1  ( .q(\sc_dm/sl1/l1_q ), .d(
        \sc_dm/sl1/mxl/muxout ), .g(n11) );
    latn_1 \sc_dm/sl0/lph3  ( .q(DMEM_eop_i_sc), .d(\sc_dm/sl0/l1_q ), .g(n1)
         );
    latn_1 \sc_dm/sl0/lph2  ( .q(\sc_dm/scn1 ), .d(\sc_dm/sl0/l1_q ), .g(n15)
         );
    mux2_1 \sc_dm/sl0/mxl/mux  ( .x(\sc_dm/sl0/mxl/muxout ), .d0(DMEM_eop_i), 
        .sl(n4), .d1(\scan[1] ) );
    latn_1 \sc_dm/sl0/mxl/lph1  ( .q(\sc_dm/sl0/l1_q ), .d(
        \sc_dm/sl0/mxl/muxout ), .g(n11) );
    latn_1 \sc_im/sl4/lph3  ( .q(IMEM_d3_i_sc), .d(\sc_im/sl4/l1_q ), .g(n1)
         );
    latn_1 \sc_im/sl4/lph2  ( .q(\scan[1] ), .d(\sc_im/sl4/l1_q ), .g(n12) );
    mux2_1 \sc_im/sl4/mxl/mux  ( .x(\sc_im/sl4/mxl/muxout ), .d0(IMEM_d3_i), 
        .sl(n4), .d1(\sc_im/scn4 ) );
    latn_1 \sc_im/sl4/mxl/lph1  ( .q(\sc_im/sl4/l1_q ), .d(
        \sc_im/sl4/mxl/muxout ), .g(n8) );
    latn_1 \sc_im/sl3/lph3  ( .q(IMEM_d2_i_sc), .d(\sc_im/sl3/l1_q ), .g(n1)
         );
    latn_1 \sc_im/sl3/lph2  ( .q(\sc_im/scn4 ), .d(\sc_im/sl3/l1_q ), .g(n14)
         );
    mux2_1 \sc_im/sl3/mxl/mux  ( .x(\sc_im/sl3/mxl/muxout ), .d0(IMEM_d2_i), 
        .sl(n7), .d1(\sc_im/scn3 ) );
    latn_1 \sc_im/sl3/mxl/lph1  ( .q(\sc_im/sl3/l1_q ), .d(
        \sc_im/sl3/mxl/muxout ), .g(n10) );
    latn_1 \sc_im/sl2/lph3  ( .q(IMEM_d1_i_sc), .d(\sc_im/sl2/l1_q ), .g(n1)
         );
    latn_1 \sc_im/sl2/lph2  ( .q(\sc_im/scn3 ), .d(\sc_im/sl2/l1_q ), .g(n14)
         );
    mux2_1 \sc_im/sl2/mxl/mux  ( .x(\sc_im/sl2/mxl/muxout ), .d0(IMEM_d1_i), 
        .sl(n6), .d1(\sc_im/scn2 ) );
    latn_1 \sc_im/sl2/mxl/lph1  ( .q(\sc_im/sl2/l1_q ), .d(
        \sc_im/sl2/mxl/muxout ), .g(n10) );
    latn_1 \sc_im/sl1/lph3  ( .q(IMEM_d0_i_sc), .d(\sc_im/sl1/l1_q ), .g(n1)
         );
    latn_1 \sc_im/sl1/lph2  ( .q(\sc_im/scn2 ), .d(\sc_im/sl1/l1_q ), .g(n12)
         );
    mux2_1 \sc_im/sl1/mxl/mux  ( .x(\sc_im/sl1/mxl/muxout ), .d0(IMEM_d0_i), 
        .sl(n6), .d1(\sc_im/scn1 ) );
    latn_1 \sc_im/sl1/mxl/lph1  ( .q(\sc_im/sl1/l1_q ), .d(
        \sc_im/sl1/mxl/muxout ), .g(n8) );
    latn_1 \sc_im/sl0/lph3  ( .q(IMEM_eop_i_sc), .d(\sc_im/sl0/l1_q ), .g(n1)
         );
    latn_1 \sc_im/sl0/lph2  ( .q(\sc_im/scn1 ), .d(\sc_im/sl0/l1_q ), .g(n14)
         );
    mux2_1 \sc_im/sl0/mxl/mux  ( .x(\sc_im/sl0/mxl/muxout ), .d0(IMEM_eop_i), 
        .sl(n6), .d1(test_si) );
    latn_1 \sc_im/sl0/mxl/lph1  ( .q(\sc_im/sl0/l1_q ), .d(
        \sc_im/sl0/mxl/muxout ), .g(n10) );
    buf_3 U1 ( .x(n5), .a(test_se) );
    buf_1 U2 ( .x(n1), .a(phi3) );
    buf_1 U3 ( .x(n3), .a(phi3) );
    buf_3 U4 ( .x(n2), .a(phi3) );
    buf_3 U5 ( .x(n4), .a(test_se) );
    buf_3 U6 ( .x(n7), .a(test_se) );
    buf_3 U7 ( .x(n6), .a(test_se) );
    buf_3 U8 ( .x(n8), .a(phi1) );
    buf_3 U9 ( .x(n11), .a(phi1) );
    buf_3 U10 ( .x(n9), .a(phi1) );
    buf_3 U11 ( .x(n10), .a(phi1) );
    buf_3 U12 ( .x(n12), .a(phi2) );
    buf_3 U13 ( .x(n15), .a(phi2) );
    buf_3 U14 ( .x(n13), .a(phi2) );
    buf_3 U15 ( .x(n14), .a(phi2) );
endmodule


module chain_sendmux8_6 ( ctrlack, oh, ol, i_h, i_l, ctrlreq, oa );
output [7:0] oh;
output [7:0] ol;
input  [7:0] i_h;
input  [7:0] i_l;
input  ctrlreq, oa;
output ctrlack;
    wire \drive[1] , \drive[0] , \U1693/drivemonitor , \U1693/naa , 
        \U1693/net2 , \U1693/net3 , \U1693/bdone , \U1693/U1702/Z ;
    and2_1 \U33_0_/U8  ( .x(oh[0]), .a(i_h[0]), .b(\drive[1] ) );
    and2_1 \U33_1_/U8  ( .x(oh[1]), .a(i_h[1]), .b(\drive[1] ) );
    and2_1 \U33_2_/U8  ( .x(oh[2]), .a(i_h[2]), .b(\drive[1] ) );
    and2_1 \U33_3_/U8  ( .x(oh[3]), .a(i_h[3]), .b(\drive[1] ) );
    and2_1 \U33_4_/U8  ( .x(oh[4]), .a(i_h[4]), .b(\drive[1] ) );
    and2_1 \U33_5_/U8  ( .x(oh[5]), .a(i_h[5]), .b(\drive[1] ) );
    and2_1 \U33_6_/U8  ( .x(oh[6]), .a(i_h[6]), .b(\drive[1] ) );
    and2_1 \U33_7_/U8  ( .x(oh[7]), .a(i_h[7]), .b(\drive[1] ) );
    and2_1 \U1670_0_/U8  ( .x(ol[0]), .a(\drive[0] ), .b(i_l[0]) );
    and2_1 \U1670_1_/U8  ( .x(ol[1]), .a(\drive[0] ), .b(i_l[1]) );
    and2_1 \U1670_2_/U8  ( .x(ol[2]), .a(\drive[0] ), .b(i_l[2]) );
    and2_1 \U1670_3_/U8  ( .x(ol[3]), .a(\drive[0] ), .b(i_l[3]) );
    and2_1 \U1670_4_/U8  ( .x(ol[4]), .a(\drive[0] ), .b(i_l[4]) );
    and2_1 \U1670_5_/U8  ( .x(ol[5]), .a(\drive[0] ), .b(i_l[5]) );
    and2_1 \U1670_6_/U8  ( .x(ol[6]), .a(\drive[0] ), .b(i_l[6]) );
    and2_1 \U1670_7_/U8  ( .x(ol[7]), .a(\drive[0] ), .b(i_l[7]) );
    nor2_2 \U1693/U1703/U6  ( .x(ctrlack), .a(\U1693/drivemonitor ), .b(
        \U1693/naa ) );
    inv_2 \U1693/U1699/U3  ( .x(\U1693/net2 ), .a(\U1693/net3 ) );
    and2_4 \U1693/U2_0_/U8  ( .x(\drive[0] ), .a(ctrlreq), .b(\U1693/net2 ) );
    and2_4 \U1693/U2_1_/U8  ( .x(\drive[1] ), .a(ctrlreq), .b(\U1693/net2 ) );
    inv_1 \U1693/U1701/U3  ( .x(\U1693/naa ), .a(\U1693/bdone ) );
    ao222_1 \U1693/U13/U18/U1/U1  ( .x(\U1693/drivemonitor ), .a(\drive[1] ), 
        .b(\drive[0] ), .c(\drive[1] ), .d(\U1693/drivemonitor ), .e(
        \drive[0] ), .f(\U1693/drivemonitor ) );
    aoi21_1 \U1693/U1702/U30/U1/U1  ( .x(\U1693/bdone ), .a(\U1693/U1702/Z ), 
        .b(oa), .c(\U1693/net2 ) );
    inv_1 \U1693/U1702/U30/U1/U2  ( .x(\U1693/U1702/Z ), .a(\U1693/bdone ) );
    ao23_1 \U1693/U1693/U21/U1/U1  ( .x(\U1693/net3 ), .a(ctrlreq), .b(
        \U1693/net3 ), .c(ctrlreq), .d(\U1693/drivemonitor ), .e(oa) );
endmodule


module chain_sendmux8_5 ( ctrlack, oh, ol, i_h, i_l, ctrlreq, oa );
output [7:0] oh;
output [7:0] ol;
input  [7:0] i_h;
input  [7:0] i_l;
input  ctrlreq, oa;
output ctrlack;
    wire \drive[1] , \drive[0] , \U1693/drivemonitor , \U1693/naa , 
        \U1693/net2 , \U1693/net3 , \U1693/bdone , \U1693/U1702/Z ;
    and2_1 \U33_0_/U8  ( .x(oh[0]), .a(i_h[0]), .b(\drive[1] ) );
    and2_1 \U33_1_/U8  ( .x(oh[1]), .a(i_h[1]), .b(\drive[1] ) );
    and2_1 \U33_2_/U8  ( .x(oh[2]), .a(i_h[2]), .b(\drive[1] ) );
    and2_1 \U33_3_/U8  ( .x(oh[3]), .a(i_h[3]), .b(\drive[1] ) );
    and2_1 \U33_4_/U8  ( .x(oh[4]), .a(i_h[4]), .b(\drive[1] ) );
    and2_1 \U33_5_/U8  ( .x(oh[5]), .a(i_h[5]), .b(\drive[1] ) );
    and2_1 \U33_6_/U8  ( .x(oh[6]), .a(i_h[6]), .b(\drive[1] ) );
    and2_1 \U33_7_/U8  ( .x(oh[7]), .a(i_h[7]), .b(\drive[1] ) );
    and2_1 \U1670_0_/U8  ( .x(ol[0]), .a(\drive[0] ), .b(i_l[0]) );
    and2_1 \U1670_1_/U8  ( .x(ol[1]), .a(\drive[0] ), .b(i_l[1]) );
    and2_1 \U1670_2_/U8  ( .x(ol[2]), .a(\drive[0] ), .b(i_l[2]) );
    and2_1 \U1670_3_/U8  ( .x(ol[3]), .a(\drive[0] ), .b(i_l[3]) );
    and2_1 \U1670_4_/U8  ( .x(ol[4]), .a(\drive[0] ), .b(i_l[4]) );
    and2_1 \U1670_5_/U8  ( .x(ol[5]), .a(\drive[0] ), .b(i_l[5]) );
    and2_1 \U1670_6_/U8  ( .x(ol[6]), .a(\drive[0] ), .b(i_l[6]) );
    and2_1 \U1670_7_/U8  ( .x(ol[7]), .a(\drive[0] ), .b(i_l[7]) );
    nor2_2 \U1693/U1703/U6  ( .x(ctrlack), .a(\U1693/drivemonitor ), .b(
        \U1693/naa ) );
    inv_2 \U1693/U1699/U3  ( .x(\U1693/net2 ), .a(\U1693/net3 ) );
    and2_4 \U1693/U2_0_/U8  ( .x(\drive[0] ), .a(ctrlreq), .b(\U1693/net2 ) );
    and2_4 \U1693/U2_1_/U8  ( .x(\drive[1] ), .a(ctrlreq), .b(\U1693/net2 ) );
    inv_1 \U1693/U1701/U3  ( .x(\U1693/naa ), .a(\U1693/bdone ) );
    ao222_1 \U1693/U13/U18/U1/U1  ( .x(\U1693/drivemonitor ), .a(\drive[1] ), 
        .b(\drive[0] ), .c(\drive[1] ), .d(\U1693/drivemonitor ), .e(
        \drive[0] ), .f(\U1693/drivemonitor ) );
    aoi21_1 \U1693/U1702/U30/U1/U1  ( .x(\U1693/bdone ), .a(\U1693/U1702/Z ), 
        .b(oa), .c(\U1693/net2 ) );
    inv_1 \U1693/U1702/U30/U1/U2  ( .x(\U1693/U1702/Z ), .a(\U1693/bdone ) );
    ao23_1 \U1693/U1693/U21/U1/U1  ( .x(\U1693/net3 ), .a(ctrlreq), .b(
        \U1693/net3 ), .c(ctrlreq), .d(\U1693/drivemonitor ), .e(oa) );
endmodule


module chain_sendmux8_4 ( ctrlack, oh, ol, i_h, i_l, ctrlreq, oa );
output [7:0] oh;
output [7:0] ol;
input  [7:0] i_h;
input  [7:0] i_l;
input  ctrlreq, oa;
output ctrlack;
    wire \drive[1] , \drive[0] , \U1693/drivemonitor , \U1693/naa , 
        \U1693/net2 , \U1693/net3 , \U1693/bdone , \U1693/U1702/Z ;
    and2_1 \U33_0_/U8  ( .x(oh[0]), .a(i_h[0]), .b(\drive[1] ) );
    and2_1 \U33_1_/U8  ( .x(oh[1]), .a(i_h[1]), .b(\drive[1] ) );
    and2_1 \U33_2_/U8  ( .x(oh[2]), .a(i_h[2]), .b(\drive[1] ) );
    and2_1 \U33_3_/U8  ( .x(oh[3]), .a(i_h[3]), .b(\drive[1] ) );
    and2_1 \U33_4_/U8  ( .x(oh[4]), .a(i_h[4]), .b(\drive[1] ) );
    and2_1 \U33_5_/U8  ( .x(oh[5]), .a(i_h[5]), .b(\drive[1] ) );
    and2_1 \U33_6_/U8  ( .x(oh[6]), .a(i_h[6]), .b(\drive[1] ) );
    and2_1 \U33_7_/U8  ( .x(oh[7]), .a(i_h[7]), .b(\drive[1] ) );
    and2_1 \U1670_0_/U8  ( .x(ol[0]), .a(\drive[0] ), .b(i_l[0]) );
    and2_1 \U1670_1_/U8  ( .x(ol[1]), .a(\drive[0] ), .b(i_l[1]) );
    and2_1 \U1670_2_/U8  ( .x(ol[2]), .a(\drive[0] ), .b(i_l[2]) );
    and2_1 \U1670_3_/U8  ( .x(ol[3]), .a(\drive[0] ), .b(i_l[3]) );
    and2_1 \U1670_4_/U8  ( .x(ol[4]), .a(\drive[0] ), .b(i_l[4]) );
    and2_1 \U1670_5_/U8  ( .x(ol[5]), .a(\drive[0] ), .b(i_l[5]) );
    and2_1 \U1670_6_/U8  ( .x(ol[6]), .a(\drive[0] ), .b(i_l[6]) );
    and2_1 \U1670_7_/U8  ( .x(ol[7]), .a(\drive[0] ), .b(i_l[7]) );
    nor2_2 \U1693/U1703/U6  ( .x(ctrlack), .a(\U1693/drivemonitor ), .b(
        \U1693/naa ) );
    inv_2 \U1693/U1699/U3  ( .x(\U1693/net2 ), .a(\U1693/net3 ) );
    and2_4 \U1693/U2_0_/U8  ( .x(\drive[0] ), .a(ctrlreq), .b(\U1693/net2 ) );
    and2_4 \U1693/U2_1_/U8  ( .x(\drive[1] ), .a(ctrlreq), .b(\U1693/net2 ) );
    inv_1 \U1693/U1701/U3  ( .x(\U1693/naa ), .a(\U1693/bdone ) );
    ao222_1 \U1693/U13/U18/U1/U1  ( .x(\U1693/drivemonitor ), .a(\drive[1] ), 
        .b(\drive[0] ), .c(\drive[1] ), .d(\U1693/drivemonitor ), .e(
        \drive[0] ), .f(\U1693/drivemonitor ) );
    aoi21_1 \U1693/U1702/U30/U1/U1  ( .x(\U1693/bdone ), .a(\U1693/U1702/Z ), 
        .b(oa), .c(\U1693/net2 ) );
    inv_1 \U1693/U1702/U30/U1/U2  ( .x(\U1693/U1702/Z ), .a(\U1693/bdone ) );
    ao23_1 \U1693/U1693/U21/U1/U1  ( .x(\U1693/net3 ), .a(ctrlreq), .b(
        \U1693/net3 ), .c(ctrlreq), .d(\U1693/drivemonitor ), .e(oa) );
endmodule


module chain_sendmux8_7 ( ctrlack, oh, ol, i_h, i_l, ctrlreq, oa );
output [7:0] oh;
output [7:0] ol;
input  [7:0] i_h;
input  [7:0] i_l;
input  ctrlreq, oa;
output ctrlack;
    wire \drive[1] , \drive[0] , \U1693/drivemonitor , \U1693/naa , 
        \U1693/net2 , \U1693/net3 , \U1693/bdone , \U1693/U1702/Z ;
    and2_1 \U33_0_/U8  ( .x(oh[0]), .a(i_h[0]), .b(\drive[1] ) );
    and2_1 \U33_1_/U8  ( .x(oh[1]), .a(i_h[1]), .b(\drive[1] ) );
    and2_1 \U33_2_/U8  ( .x(oh[2]), .a(i_h[2]), .b(\drive[1] ) );
    and2_1 \U33_3_/U8  ( .x(oh[3]), .a(i_h[3]), .b(\drive[1] ) );
    and2_1 \U33_4_/U8  ( .x(oh[4]), .a(i_h[4]), .b(\drive[1] ) );
    and2_1 \U33_5_/U8  ( .x(oh[5]), .a(i_h[5]), .b(\drive[1] ) );
    and2_1 \U33_6_/U8  ( .x(oh[6]), .a(i_h[6]), .b(\drive[1] ) );
    and2_1 \U33_7_/U8  ( .x(oh[7]), .a(i_h[7]), .b(\drive[1] ) );
    and2_1 \U1670_0_/U8  ( .x(ol[0]), .a(\drive[0] ), .b(i_l[0]) );
    and2_1 \U1670_1_/U8  ( .x(ol[1]), .a(\drive[0] ), .b(i_l[1]) );
    and2_1 \U1670_2_/U8  ( .x(ol[2]), .a(\drive[0] ), .b(i_l[2]) );
    and2_1 \U1670_3_/U8  ( .x(ol[3]), .a(\drive[0] ), .b(i_l[3]) );
    and2_1 \U1670_4_/U8  ( .x(ol[4]), .a(\drive[0] ), .b(i_l[4]) );
    and2_1 \U1670_5_/U8  ( .x(ol[5]), .a(\drive[0] ), .b(i_l[5]) );
    and2_1 \U1670_6_/U8  ( .x(ol[6]), .a(\drive[0] ), .b(i_l[6]) );
    and2_1 \U1670_7_/U8  ( .x(ol[7]), .a(\drive[0] ), .b(i_l[7]) );
    nor2_2 \U1693/U1703/U6  ( .x(ctrlack), .a(\U1693/drivemonitor ), .b(
        \U1693/naa ) );
    inv_2 \U1693/U1699/U3  ( .x(\U1693/net2 ), .a(\U1693/net3 ) );
    and2_4 \U1693/U2_0_/U8  ( .x(\drive[0] ), .a(ctrlreq), .b(\U1693/net2 ) );
    and2_4 \U1693/U2_1_/U8  ( .x(\drive[1] ), .a(ctrlreq), .b(\U1693/net2 ) );
    inv_1 \U1693/U1701/U3  ( .x(\U1693/naa ), .a(\U1693/bdone ) );
    ao222_1 \U1693/U13/U18/U1/U1  ( .x(\U1693/drivemonitor ), .a(\drive[1] ), 
        .b(\drive[0] ), .c(\drive[1] ), .d(\U1693/drivemonitor ), .e(
        \drive[0] ), .f(\U1693/drivemonitor ) );
    aoi21_1 \U1693/U1702/U30/U1/U1  ( .x(\U1693/bdone ), .a(\U1693/U1702/Z ), 
        .b(oa), .c(\U1693/net2 ) );
    inv_1 \U1693/U1702/U30/U1/U2  ( .x(\U1693/U1702/Z ), .a(\U1693/bdone ) );
    ao23_1 \U1693/U1693/U21/U1/U1  ( .x(\U1693/net3 ), .a(ctrlreq), .b(
        \U1693/net3 ), .c(ctrlreq), .d(\U1693/drivemonitor ), .e(oa) );
endmodule


module chain_sendword_0 ( ctrlack, oh, ol, chainackff, ctrlreq, ih, il );
output [7:0] oh;
output [7:0] ol;
input  [31:0] ih;
input  [31:0] il;
input  chainackff, ctrlreq;
output ctrlack;
    wire net44, \fourth_ol[7] , \fourth_ol[6] , \fourth_ol[5] , \fourth_ol[4] , 
        \fourth_ol[3] , \fourth_ol[2] , \fourth_ol[1] , \fourth_ol[0] , 
        \fourth_oh[7] , \fourth_oh[6] , \fourth_oh[5] , \fourth_oh[4] , 
        \fourth_oh[3] , \fourth_oh[2] , \fourth_oh[1] , \fourth_oh[0] , net51, 
        \third_ol[7] , \third_ol[6] , \third_ol[5] , \third_ol[4] , 
        \third_ol[3] , \third_ol[2] , \third_ol[1] , \third_ol[0] , 
        \third_oh[7] , \third_oh[6] , \third_oh[5] , \third_oh[4] , 
        \third_oh[3] , \third_oh[2] , \third_oh[1] , \third_oh[0] , net58, 
        \second_ol[7] , \second_ol[6] , \second_ol[5] , \second_ol[4] , 
        \second_ol[3] , \second_ol[2] , \second_ol[1] , \second_ol[0] , 
        \second_oh[7] , \second_oh[6] , \second_oh[5] , \second_oh[4] , 
        \second_oh[3] , \second_oh[2] , \second_oh[1] , \second_oh[0] , 
        bctrlreq, \first_ol[7] , \first_ol[6] , \first_ol[5] , \first_ol[4] , 
        \first_ol[3] , \first_ol[2] , \first_ol[1] , \first_ol[0] , 
        \first_oh[7] , \first_oh[6] , \first_oh[5] , \first_oh[4] , 
        \first_oh[3] , \first_oh[2] , \first_oh[1] , \first_oh[0] , 
        \U309_0_/n5 , \U309_0_/n1 , \U309_0_/n2 , \U309_0_/n3 , \U309_0_/n4 , 
        \U309_1_/n5 , \U309_1_/n1 , \U309_1_/n2 , \U309_1_/n3 , \U309_1_/n4 , 
        \U309_2_/n5 , \U309_2_/n1 , \U309_2_/n2 , \U309_2_/n3 , \U309_2_/n4 , 
        \U309_3_/n5 , \U309_3_/n1 , \U309_3_/n2 , \U309_3_/n3 , \U309_3_/n4 , 
        \U309_4_/n5 , \U309_4_/n1 , \U309_4_/n2 , \U309_4_/n3 , \U309_4_/n4 , 
        \U309_5_/n5 , \U309_5_/n1 , \U309_5_/n2 , \U309_5_/n3 , \U309_5_/n4 , 
        \U309_6_/n5 , \U309_6_/n1 , \U309_6_/n2 , \U309_6_/n3 , \U309_6_/n4 , 
        \U309_7_/n5 , \U309_7_/n1 , \U309_7_/n2 , \U309_7_/n3 , \U309_7_/n4 , 
        \U310_0_/n5 , \U310_0_/n1 , \U310_0_/n2 , \U310_0_/n3 , \U310_0_/n4 , 
        \U310_1_/n5 , \U310_1_/n1 , \U310_1_/n2 , \U310_1_/n3 , \U310_1_/n4 , 
        \U310_2_/n5 , \U310_2_/n1 , \U310_2_/n2 , \U310_2_/n3 , \U310_2_/n4 , 
        \U310_3_/n5 , \U310_3_/n1 , \U310_3_/n2 , \U310_3_/n3 , \U310_3_/n4 , 
        \U310_4_/n5 , \U310_4_/n1 , \U310_4_/n2 , \U310_4_/n3 , \U310_4_/n4 , 
        \U310_5_/n5 , \U310_5_/n1 , \U310_5_/n2 , \U310_5_/n3 , \U310_5_/n4 , 
        \U310_6_/n5 , \U310_6_/n1 , \U310_6_/n2 , \U310_6_/n3 , \U310_6_/n4 , 
        \U310_7_/n5 , \U310_7_/n1 , \U310_7_/n2 , \U310_7_/n3 , \U310_7_/n4 ;
    chain_sendmux8_6 I4 ( .ctrlack(ctrlack), .oh({\fourth_oh[7] , 
        \fourth_oh[6] , \fourth_oh[5] , \fourth_oh[4] , \fourth_oh[3] , 
        \fourth_oh[2] , \fourth_oh[1] , \fourth_oh[0] }), .ol({\fourth_ol[7] , 
        \fourth_ol[6] , \fourth_ol[5] , \fourth_ol[4] , \fourth_ol[3] , 
        \fourth_ol[2] , \fourth_ol[1] , \fourth_ol[0] }), .i_h(ih[7:0]), .i_l(
        il[7:0]), .ctrlreq(net44), .oa(chainackff) );
    chain_sendmux8_5 I3 ( .ctrlack(net44), .oh({\third_oh[7] , \third_oh[6] , 
        \third_oh[5] , \third_oh[4] , \third_oh[3] , \third_oh[2] , 
        \third_oh[1] , \third_oh[0] }), .ol({\third_ol[7] , \third_ol[6] , 
        \third_ol[5] , \third_ol[4] , \third_ol[3] , \third_ol[2] , 
        \third_ol[1] , \third_ol[0] }), .i_h(ih[15:8]), .i_l(il[15:8]), 
        .ctrlreq(net51), .oa(chainackff) );
    chain_sendmux8_4 I2 ( .ctrlack(net51), .oh({\second_oh[7] , \second_oh[6] , 
        \second_oh[5] , \second_oh[4] , \second_oh[3] , \second_oh[2] , 
        \second_oh[1] , \second_oh[0] }), .ol({\second_ol[7] , \second_ol[6] , 
        \second_ol[5] , \second_ol[4] , \second_ol[3] , \second_ol[2] , 
        \second_ol[1] , \second_ol[0] }), .i_h(ih[23:16]), .i_l(il[23:16]), 
        .ctrlreq(net58), .oa(chainackff) );
    chain_sendmux8_7 U320 ( .ctrlack(net58), .oh({\first_oh[7] , \first_oh[6] , 
        \first_oh[5] , \first_oh[4] , \first_oh[3] , \first_oh[2] , 
        \first_oh[1] , \first_oh[0] }), .ol({\first_ol[7] , \first_ol[6] , 
        \first_ol[5] , \first_ol[4] , \first_ol[3] , \first_ol[2] , 
        \first_ol[1] , \first_ol[0] }), .i_h(ih[31:24]), .i_l(il[31:24]), 
        .ctrlreq(bctrlreq), .oa(chainackff) );
    buf_2 \U328/U7  ( .x(bctrlreq), .a(ctrlreq) );
    and4_2 \U309_0_/U24  ( .x(\U309_0_/n5 ), .a(\U309_0_/n1 ), .b(\U309_0_/n2 
        ), .c(\U309_0_/n3 ), .d(\U309_0_/n4 ) );
    inv_1 \U309_0_/U1  ( .x(\U309_0_/n1 ), .a(\fourth_oh[0] ) );
    inv_1 \U309_0_/U2  ( .x(\U309_0_/n2 ), .a(\third_oh[0] ) );
    inv_1 \U309_0_/U3  ( .x(\U309_0_/n3 ), .a(\second_oh[0] ) );
    inv_1 \U309_0_/U4  ( .x(\U309_0_/n4 ), .a(\first_oh[0] ) );
    inv_4 \U309_0_/U5  ( .x(oh[0]), .a(\U309_0_/n5 ) );
    and4_2 \U309_1_/U24  ( .x(\U309_1_/n5 ), .a(\U309_1_/n1 ), .b(\U309_1_/n2 
        ), .c(\U309_1_/n3 ), .d(\U309_1_/n4 ) );
    inv_1 \U309_1_/U1  ( .x(\U309_1_/n1 ), .a(\fourth_oh[1] ) );
    inv_1 \U309_1_/U2  ( .x(\U309_1_/n2 ), .a(\third_oh[1] ) );
    inv_1 \U309_1_/U3  ( .x(\U309_1_/n3 ), .a(\second_oh[1] ) );
    inv_1 \U309_1_/U4  ( .x(\U309_1_/n4 ), .a(\first_oh[1] ) );
    inv_4 \U309_1_/U5  ( .x(oh[1]), .a(\U309_1_/n5 ) );
    and4_2 \U309_2_/U24  ( .x(\U309_2_/n5 ), .a(\U309_2_/n1 ), .b(\U309_2_/n2 
        ), .c(\U309_2_/n3 ), .d(\U309_2_/n4 ) );
    inv_1 \U309_2_/U1  ( .x(\U309_2_/n1 ), .a(\fourth_oh[2] ) );
    inv_1 \U309_2_/U2  ( .x(\U309_2_/n2 ), .a(\third_oh[2] ) );
    inv_1 \U309_2_/U3  ( .x(\U309_2_/n3 ), .a(\second_oh[2] ) );
    inv_1 \U309_2_/U4  ( .x(\U309_2_/n4 ), .a(\first_oh[2] ) );
    inv_4 \U309_2_/U5  ( .x(oh[2]), .a(\U309_2_/n5 ) );
    and4_2 \U309_3_/U24  ( .x(\U309_3_/n5 ), .a(\U309_3_/n1 ), .b(\U309_3_/n2 
        ), .c(\U309_3_/n3 ), .d(\U309_3_/n4 ) );
    inv_1 \U309_3_/U1  ( .x(\U309_3_/n1 ), .a(\fourth_oh[3] ) );
    inv_1 \U309_3_/U2  ( .x(\U309_3_/n2 ), .a(\third_oh[3] ) );
    inv_1 \U309_3_/U3  ( .x(\U309_3_/n3 ), .a(\second_oh[3] ) );
    inv_1 \U309_3_/U4  ( .x(\U309_3_/n4 ), .a(\first_oh[3] ) );
    inv_4 \U309_3_/U5  ( .x(oh[3]), .a(\U309_3_/n5 ) );
    and4_2 \U309_4_/U24  ( .x(\U309_4_/n5 ), .a(\U309_4_/n1 ), .b(\U309_4_/n2 
        ), .c(\U309_4_/n3 ), .d(\U309_4_/n4 ) );
    inv_1 \U309_4_/U1  ( .x(\U309_4_/n1 ), .a(\fourth_oh[4] ) );
    inv_1 \U309_4_/U2  ( .x(\U309_4_/n2 ), .a(\third_oh[4] ) );
    inv_1 \U309_4_/U3  ( .x(\U309_4_/n3 ), .a(\second_oh[4] ) );
    inv_1 \U309_4_/U4  ( .x(\U309_4_/n4 ), .a(\first_oh[4] ) );
    inv_4 \U309_4_/U5  ( .x(oh[4]), .a(\U309_4_/n5 ) );
    and4_2 \U309_5_/U24  ( .x(\U309_5_/n5 ), .a(\U309_5_/n1 ), .b(\U309_5_/n2 
        ), .c(\U309_5_/n3 ), .d(\U309_5_/n4 ) );
    inv_1 \U309_5_/U1  ( .x(\U309_5_/n1 ), .a(\fourth_oh[5] ) );
    inv_1 \U309_5_/U2  ( .x(\U309_5_/n2 ), .a(\third_oh[5] ) );
    inv_1 \U309_5_/U3  ( .x(\U309_5_/n3 ), .a(\second_oh[5] ) );
    inv_1 \U309_5_/U4  ( .x(\U309_5_/n4 ), .a(\first_oh[5] ) );
    inv_4 \U309_5_/U5  ( .x(oh[5]), .a(\U309_5_/n5 ) );
    and4_2 \U309_6_/U24  ( .x(\U309_6_/n5 ), .a(\U309_6_/n1 ), .b(\U309_6_/n2 
        ), .c(\U309_6_/n3 ), .d(\U309_6_/n4 ) );
    inv_1 \U309_6_/U1  ( .x(\U309_6_/n1 ), .a(\fourth_oh[6] ) );
    inv_1 \U309_6_/U2  ( .x(\U309_6_/n2 ), .a(\third_oh[6] ) );
    inv_1 \U309_6_/U3  ( .x(\U309_6_/n3 ), .a(\second_oh[6] ) );
    inv_1 \U309_6_/U4  ( .x(\U309_6_/n4 ), .a(\first_oh[6] ) );
    inv_4 \U309_6_/U5  ( .x(oh[6]), .a(\U309_6_/n5 ) );
    and4_2 \U309_7_/U24  ( .x(\U309_7_/n5 ), .a(\U309_7_/n1 ), .b(\U309_7_/n2 
        ), .c(\U309_7_/n3 ), .d(\U309_7_/n4 ) );
    inv_1 \U309_7_/U1  ( .x(\U309_7_/n1 ), .a(\fourth_oh[7] ) );
    inv_1 \U309_7_/U2  ( .x(\U309_7_/n2 ), .a(\third_oh[7] ) );
    inv_1 \U309_7_/U3  ( .x(\U309_7_/n3 ), .a(\second_oh[7] ) );
    inv_1 \U309_7_/U4  ( .x(\U309_7_/n4 ), .a(\first_oh[7] ) );
    inv_4 \U309_7_/U5  ( .x(oh[7]), .a(\U309_7_/n5 ) );
    and4_2 \U310_0_/U24  ( .x(\U310_0_/n5 ), .a(\U310_0_/n1 ), .b(\U310_0_/n2 
        ), .c(\U310_0_/n3 ), .d(\U310_0_/n4 ) );
    inv_1 \U310_0_/U1  ( .x(\U310_0_/n1 ), .a(\fourth_ol[0] ) );
    inv_1 \U310_0_/U2  ( .x(\U310_0_/n2 ), .a(\third_ol[0] ) );
    inv_1 \U310_0_/U3  ( .x(\U310_0_/n3 ), .a(\second_ol[0] ) );
    inv_1 \U310_0_/U4  ( .x(\U310_0_/n4 ), .a(\first_ol[0] ) );
    inv_4 \U310_0_/U5  ( .x(ol[0]), .a(\U310_0_/n5 ) );
    and4_2 \U310_1_/U24  ( .x(\U310_1_/n5 ), .a(\U310_1_/n1 ), .b(\U310_1_/n2 
        ), .c(\U310_1_/n3 ), .d(\U310_1_/n4 ) );
    inv_1 \U310_1_/U1  ( .x(\U310_1_/n1 ), .a(\fourth_ol[1] ) );
    inv_1 \U310_1_/U2  ( .x(\U310_1_/n2 ), .a(\third_ol[1] ) );
    inv_1 \U310_1_/U3  ( .x(\U310_1_/n3 ), .a(\second_ol[1] ) );
    inv_1 \U310_1_/U4  ( .x(\U310_1_/n4 ), .a(\first_ol[1] ) );
    inv_4 \U310_1_/U5  ( .x(ol[1]), .a(\U310_1_/n5 ) );
    and4_2 \U310_2_/U24  ( .x(\U310_2_/n5 ), .a(\U310_2_/n1 ), .b(\U310_2_/n2 
        ), .c(\U310_2_/n3 ), .d(\U310_2_/n4 ) );
    inv_1 \U310_2_/U1  ( .x(\U310_2_/n1 ), .a(\fourth_ol[2] ) );
    inv_1 \U310_2_/U2  ( .x(\U310_2_/n2 ), .a(\third_ol[2] ) );
    inv_1 \U310_2_/U3  ( .x(\U310_2_/n3 ), .a(\second_ol[2] ) );
    inv_1 \U310_2_/U4  ( .x(\U310_2_/n4 ), .a(\first_ol[2] ) );
    inv_4 \U310_2_/U5  ( .x(ol[2]), .a(\U310_2_/n5 ) );
    and4_2 \U310_3_/U24  ( .x(\U310_3_/n5 ), .a(\U310_3_/n1 ), .b(\U310_3_/n2 
        ), .c(\U310_3_/n3 ), .d(\U310_3_/n4 ) );
    inv_1 \U310_3_/U1  ( .x(\U310_3_/n1 ), .a(\fourth_ol[3] ) );
    inv_1 \U310_3_/U2  ( .x(\U310_3_/n2 ), .a(\third_ol[3] ) );
    inv_1 \U310_3_/U3  ( .x(\U310_3_/n3 ), .a(\second_ol[3] ) );
    inv_1 \U310_3_/U4  ( .x(\U310_3_/n4 ), .a(\first_ol[3] ) );
    inv_4 \U310_3_/U5  ( .x(ol[3]), .a(\U310_3_/n5 ) );
    and4_2 \U310_4_/U24  ( .x(\U310_4_/n5 ), .a(\U310_4_/n1 ), .b(\U310_4_/n2 
        ), .c(\U310_4_/n3 ), .d(\U310_4_/n4 ) );
    inv_1 \U310_4_/U1  ( .x(\U310_4_/n1 ), .a(\fourth_ol[4] ) );
    inv_1 \U310_4_/U2  ( .x(\U310_4_/n2 ), .a(\third_ol[4] ) );
    inv_1 \U310_4_/U3  ( .x(\U310_4_/n3 ), .a(\second_ol[4] ) );
    inv_1 \U310_4_/U4  ( .x(\U310_4_/n4 ), .a(\first_ol[4] ) );
    inv_4 \U310_4_/U5  ( .x(ol[4]), .a(\U310_4_/n5 ) );
    and4_2 \U310_5_/U24  ( .x(\U310_5_/n5 ), .a(\U310_5_/n1 ), .b(\U310_5_/n2 
        ), .c(\U310_5_/n3 ), .d(\U310_5_/n4 ) );
    inv_1 \U310_5_/U1  ( .x(\U310_5_/n1 ), .a(\fourth_ol[5] ) );
    inv_1 \U310_5_/U2  ( .x(\U310_5_/n2 ), .a(\third_ol[5] ) );
    inv_1 \U310_5_/U3  ( .x(\U310_5_/n3 ), .a(\second_ol[5] ) );
    inv_1 \U310_5_/U4  ( .x(\U310_5_/n4 ), .a(\first_ol[5] ) );
    inv_4 \U310_5_/U5  ( .x(ol[5]), .a(\U310_5_/n5 ) );
    and4_2 \U310_6_/U24  ( .x(\U310_6_/n5 ), .a(\U310_6_/n1 ), .b(\U310_6_/n2 
        ), .c(\U310_6_/n3 ), .d(\U310_6_/n4 ) );
    inv_1 \U310_6_/U1  ( .x(\U310_6_/n1 ), .a(\fourth_ol[6] ) );
    inv_1 \U310_6_/U2  ( .x(\U310_6_/n2 ), .a(\third_ol[6] ) );
    inv_1 \U310_6_/U3  ( .x(\U310_6_/n3 ), .a(\second_ol[6] ) );
    inv_1 \U310_6_/U4  ( .x(\U310_6_/n4 ), .a(\first_ol[6] ) );
    inv_4 \U310_6_/U5  ( .x(ol[6]), .a(\U310_6_/n5 ) );
    and4_2 \U310_7_/U24  ( .x(\U310_7_/n5 ), .a(\U310_7_/n1 ), .b(\U310_7_/n2 
        ), .c(\U310_7_/n3 ), .d(\U310_7_/n4 ) );
    inv_1 \U310_7_/U1  ( .x(\U310_7_/n1 ), .a(\fourth_ol[7] ) );
    inv_1 \U310_7_/U2  ( .x(\U310_7_/n2 ), .a(\third_ol[7] ) );
    inv_1 \U310_7_/U3  ( .x(\U310_7_/n3 ), .a(\second_ol[7] ) );
    inv_1 \U310_7_/U4  ( .x(\U310_7_/n4 ), .a(\first_ol[7] ) );
    inv_4 \U310_7_/U5  ( .x(ol[7]), .a(\U310_7_/n5 ) );
endmodule


module chain_dr8bit_completion_12 ( o, i );
input  [15:0] i;
output o;
    wire \nx[0] , \nx[1] , \nx[2] , \nx[3] , \ny[0] , \ny[1] , \ny[2] , 
        \ny[3] , y, x, \U6/Z , \U3/net3 , \U3/U20/Z , \U3/net2 , \U3/U21/Z , 
        \U3/U19/Z , \U5/net3 , \U5/U20/Z , \U5/net2 , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_15 ( o, i );
input  [15:0] i;
output o;
    wire \nx[0] , \nx[1] , \nx[2] , \nx[3] , \ny[0] , \ny[1] , \ny[2] , 
        \ny[3] , y, x, \U6/Z , \U3/net3 , \U3/U20/Z , \U3/net2 , \U3/U21/Z , 
        \U3/U19/Z , \U5/net3 , \U5/U20/Z , \U5/net2 , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_14 ( o, i );
input  [15:0] i;
output o;
    wire \nx[0] , \nx[1] , \nx[2] , \nx[3] , \ny[0] , \ny[1] , \ny[2] , 
        \ny[3] , y, x, \U6/Z , \U3/net3 , \U3/U20/Z , \U3/net2 , \U3/U21/Z , 
        \U3/U19/Z , \U5/net3 , \U5/U20/Z , \U5/net2 , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_13 ( o, i );
input  [15:0] i;
output o;
    wire \nx[0] , \nx[1] , \nx[2] , \nx[3] , \ny[0] , \ny[1] , \ny[2] , 
        \ny[3] , y, x, \U6/Z , \U3/net3 , \U3/U20/Z , \U3/net2 , \U3/U21/Z , 
        \U3/U19/Z , \U5/net3 , \U5/U20/Z , \U5/net2 , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr32bit_completion_8 ( o, i );
input  [63:0] i;
output o;
    wire \cd[3] , \cd[2] , \cd[1] , \cd[0] , ny, \U16/Z , nx, \U6/Z , \U15/Z ;
    chain_dr8bit_completion_12 U11 ( .o(\cd[3] ), .i({i[63], i[62], i[61], 
        i[60], i[59], i[58], i[57], i[56], i[31], i[30], i[29], i[28], i[27], 
        i[26], i[25], i[24]}) );
    chain_dr8bit_completion_15 U14 ( .o(\cd[2] ), .i({i[55], i[54], i[53], 
        i[52], i[51], i[50], i[49], i[48], i[23], i[22], i[21], i[20], i[19], 
        i[18], i[17], i[16]}) );
    chain_dr8bit_completion_14 U13 ( .o(\cd[1] ), .i({i[47], i[46], i[45], 
        i[44], i[43], i[42], i[41], i[40], i[15], i[14], i[13], i[12], i[11], 
        i[10], i[9], i[8]}) );
    chain_dr8bit_completion_13 U12 ( .o(\cd[0] ), .i({i[39], i[38], i[37], 
        i[36], i[35], i[34], i[33], i[32], i[7], i[6], i[5], i[4], i[3], i[2], 
        i[1], i[0]}) );
    aoi222_1 \U16/U30/U1  ( .x(ny), .a(\cd[0] ), .b(\cd[1] ), .c(\cd[0] ), .d(
        \U16/Z ), .e(\cd[1] ), .f(\U16/Z ) );
    inv_1 \U16/U30/Uinv  ( .x(\U16/Z ), .a(ny) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(ny), .b(nx), .c(ny), .d(\U6/Z ), .e(nx), 
        .f(\U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U15/U30/U1  ( .x(nx), .a(\cd[3] ), .b(\cd[2] ), .c(\cd[3] ), .d(
        \U15/Z ), .e(\cd[2] ), .f(\U15/Z ) );
    inv_1 \U15/U30/Uinv  ( .x(\U15/Z ), .a(nx) );
endmodule


module chain_selement_ga_63 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_trhdr_0 ( chainff_ack, chainh, chainl, eop, hdrack, normal_ack, 
    notify_ack, read_req, routereq, chain_ff_h, chainack, chainff_l, eopack, 
    err, nReset, normal_response, notify_accept, notify_defer, rcol_h, rcol_l, 
    read_ack, rnw_h, rnw_l, routeack, rsize_h, rsize_l, rtag_h, rtag_l );
output [7:0] chainh;
output [7:0] chainl;
input  [7:0] chain_ff_h;
input  [7:0] chainff_l;
input  [1:0] err;
input  [2:0] rcol_h;
input  [2:0] rcol_l;
input  [1:0] rsize_h;
input  [1:0] rsize_l;
input  [4:0] rtag_h;
input  [4:0] rtag_l;
input  chainack, eopack, nReset, normal_response, notify_accept, notify_defer, 
    read_ack, rnw_h, rnw_l, routeack;
output chainff_ack, eop, hdrack, normal_ack, notify_ack, read_req, routereq;
    wire done_eop, done_pl, \net413[15] , \hdr[16] , \hdr[0] , \net413[14] , 
        \hdr[17] , \hdr[1] , \net413[13] , \net413[12] , \net413[11] , 
        \net413[10] , \net413[9] , \net413[8] , \net413[7] , \net413[6] , 
        \net413[5] , \net413[4] , \net413[3] , \net413[2] , \net413[1] , 
        \net413[0] , net364, donotify, dowrite, net383, done_defer, done_write, 
        done_read, \net343[7] , \drive_l[0] , \net343[6] , \net343[5] , 
        \net343[3] , \net343[2] , \net343[1] , \net343[0] , net340, net337, 
        \net334[7] , \drive_l[1] , \net334[6] , \net334[4] , \net334[2] , 
        \net334[1] , \net334[0] , \net284[7] , \drive_h[1] , \net284[6] , 
        \net284[5] , \net284[4] , \net284[3] , \net284[2] , \net284[1] , 
        \net284[0] , \net288[7] , \drive_h[0] , \net288[6] , \net288[5] , 
        \net288[4] , \net288[3] , \net288[2] , \net288[1] , \net288[0] , 
        net332, done_accept, net321, net359, net362, ctrl_cd, \U311/nz[0] , 
        \U311/nz[1] , \U311/x[3] , \U311/U28/Z , \U311/x[0] , \U311/U32/Z , 
        \U311/x[5] , \U311/U20/Z , \U311/x[2] , \U311/U29/Z , \U311/x[7] , 
        \U311/U25/Z , \U311/y[0] , \U311/x[1] , \U311/U33/Z , \U311/y[2] , 
        \U311/x[4] , \U311/U21/Z , \U311/x[6] , \U311/U26/Z , \U311/y[1] , 
        \U311/U34/Z , \U311/U30/Z , \U311/U19/Z , \U311/y[3] , \U311/U27/Z , 
        \U311/U35/Z , \U311/U31/Z , net407, \U151/Z , done_hdr, 
        \U319/U21/U1/loop , \U323/U21/U1/loop , \U320/U21/U1/loop , 
        \U321/U21/U1/loop , \U322/U21/U1/loop , \U210/drivemonitor , 
        \U210/naa , \U210/net2 , \U210/net3 , net0230, \U210/bdone , 
        \U210/U1702/Z , \I0/drivemonitor , \I0/naa , \I0/net2 , \I0/net3 , 
        \I0/bdone , \I0/U1702/Z ;
    chain_selement_ga_63 U215 ( .Aa(done_eop), .Br(eop), .Ar(done_pl), .Ba(
        eopack) );
    nor2_1 \U308_0_/U5  ( .x(\net413[15] ), .a(\hdr[16] ), .b(\hdr[0] ) );
    nor2_1 \U308_1_/U5  ( .x(\net413[14] ), .a(\hdr[17] ), .b(\hdr[1] ) );
    nor2_1 \U308_2_/U5  ( .x(\net413[13] ), .a(1'b0), .b(routereq) );
    nor2_1 \U308_3_/U5  ( .x(\net413[12] ), .a(routereq), .b(1'b0) );
    nor2_1 \U308_4_/U5  ( .x(\net413[11] ), .a(1'b0), .b(routereq) );
    nor2_1 \U308_5_/U5  ( .x(\net413[10] ), .a(rnw_h), .b(rnw_l) );
    nor2_1 \U308_6_/U5  ( .x(\net413[9] ), .a(rsize_h[0]), .b(rsize_l[0]) );
    nor2_1 \U308_7_/U5  ( .x(\net413[8] ), .a(rsize_h[1]), .b(rsize_l[1]) );
    nor2_1 \U308_8_/U5  ( .x(\net413[7] ), .a(rtag_h[0]), .b(rtag_l[0]) );
    nor2_1 \U308_9_/U5  ( .x(\net413[6] ), .a(rtag_h[1]), .b(rtag_l[1]) );
    nor2_1 \U308_10_/U5  ( .x(\net413[5] ), .a(rtag_h[2]), .b(rtag_l[2]) );
    nor2_1 \U308_11_/U5  ( .x(\net413[4] ), .a(rtag_h[3]), .b(rtag_l[3]) );
    nor2_1 \U308_12_/U5  ( .x(\net413[3] ), .a(rtag_h[4]), .b(rtag_l[4]) );
    nor2_1 \U308_13_/U5  ( .x(\net413[2] ), .a(rcol_h[0]), .b(rcol_l[0]) );
    nor2_1 \U308_14_/U5  ( .x(\net413[1] ), .a(rcol_h[1]), .b(rcol_l[1]) );
    nor2_1 \U308_15_/U5  ( .x(\net413[0] ), .a(rcol_h[2]), .b(rcol_l[2]) );
    or3_1 \U257/U12  ( .x(net364), .a(donotify), .b(dowrite), .c(read_ack) );
    or3_1 \U297/U12  ( .x(net383), .a(done_defer), .b(done_write), .c(
        done_read) );
    and2_2 \U237/U8  ( .x(\hdr[1] ), .a(nReset), .b(normal_response) );
    and2_1 \U307_0_/U8  ( .x(\net343[7] ), .a(\drive_l[0] ), .b(\hdr[0] ) );
    and2_1 \U307_1_/U8  ( .x(\net343[6] ), .a(\drive_l[0] ), .b(\hdr[1] ) );
    and2_1 \U307_2_/U8  ( .x(\net343[5] ), .a(\drive_l[0] ), .b(routereq) );
    and2_1 \U307_4_/U8  ( .x(\net343[3] ), .a(\drive_l[0] ), .b(routereq) );
    and2_1 \U307_5_/U8  ( .x(\net343[2] ), .a(\drive_l[0] ), .b(rnw_l) );
    and2_1 \U307_6_/U8  ( .x(\net343[1] ), .a(\drive_l[0] ), .b(rsize_l[0]) );
    and2_1 \U307_7_/U8  ( .x(\net343[0] ), .a(\drive_l[0] ), .b(rsize_l[1]) );
    and2_1 \U235/U8  ( .x(net340), .a(err[1]), .b(nReset) );
    and2_1 \U236/U8  ( .x(net337), .a(nReset), .b(err[0]) );
    and2_1 \U306_0_/U8  ( .x(\net334[7] ), .a(\hdr[16] ), .b(\drive_l[1] ) );
    and2_1 \U306_1_/U8  ( .x(\net334[6] ), .a(\hdr[17] ), .b(\drive_l[1] ) );
    and2_1 \U306_3_/U8  ( .x(\net334[4] ), .a(routereq), .b(\drive_l[1] ) );
    and2_1 \U306_5_/U8  ( .x(\net334[2] ), .a(rnw_h), .b(\drive_l[1] ) );
    and2_1 \U306_6_/U8  ( .x(\net334[1] ), .a(rsize_h[0]), .b(\drive_l[1] ) );
    and2_1 \U306_7_/U8  ( .x(\net334[0] ), .a(rsize_h[1]), .b(\drive_l[1] ) );
    and2_1 \I1_0_/U8  ( .x(\net284[7] ), .a(rtag_h[0]), .b(\drive_h[1] ) );
    and2_1 \I1_1_/U8  ( .x(\net284[6] ), .a(rtag_h[1]), .b(\drive_h[1] ) );
    and2_1 \I1_2_/U8  ( .x(\net284[5] ), .a(rtag_h[2]), .b(\drive_h[1] ) );
    and2_1 \I1_3_/U8  ( .x(\net284[4] ), .a(rtag_h[3]), .b(\drive_h[1] ) );
    and2_1 \I1_4_/U8  ( .x(\net284[3] ), .a(rtag_h[4]), .b(\drive_h[1] ) );
    and2_1 \I1_5_/U8  ( .x(\net284[2] ), .a(rcol_h[0]), .b(\drive_h[1] ) );
    and2_1 \I1_6_/U8  ( .x(\net284[1] ), .a(rcol_h[1]), .b(\drive_h[1] ) );
    and2_1 \I1_7_/U8  ( .x(\net284[0] ), .a(rcol_h[2]), .b(\drive_h[1] ) );
    and2_1 \I2_0_/U8  ( .x(\net288[7] ), .a(\drive_h[0] ), .b(rtag_l[0]) );
    and2_1 \I2_1_/U8  ( .x(\net288[6] ), .a(\drive_h[0] ), .b(rtag_l[1]) );
    and2_1 \I2_2_/U8  ( .x(\net288[5] ), .a(\drive_h[0] ), .b(rtag_l[2]) );
    and2_1 \I2_3_/U8  ( .x(\net288[4] ), .a(\drive_h[0] ), .b(rtag_l[3]) );
    and2_1 \I2_4_/U8  ( .x(\net288[3] ), .a(\drive_h[0] ), .b(rtag_l[4]) );
    and2_1 \I2_5_/U8  ( .x(\net288[2] ), .a(\drive_h[0] ), .b(rcol_l[0]) );
    and2_1 \I2_6_/U8  ( .x(\net288[1] ), .a(\drive_h[0] ), .b(rcol_l[1]) );
    and2_1 \I2_7_/U8  ( .x(\net288[0] ), .a(\drive_h[0] ), .b(rcol_l[2]) );
    inv_1 \U318/U3  ( .x(net332), .a(routereq) );
    or2_4 \U255/U12  ( .x(notify_ack), .a(done_accept), .b(done_defer) );
    or2_4 \U228/U12  ( .x(\hdr[17] ), .a(notify_defer), .b(notify_accept) );
    or2_4 \U204/U12  ( .x(net321), .a(net359), .b(net362) );
    or2_4 \U221/U12  ( .x(\hdr[16] ), .a(net359), .b(notify_defer) );
    or2_4 \U252/U12  ( .x(normal_ack), .a(done_write), .b(done_read) );
    or2_4 \U280/U12  ( .x(\hdr[0] ), .a(net362), .b(notify_accept) );
    or2_4 \U317/U12  ( .x(routereq), .a(\hdr[17] ), .b(net321) );
    or3_4 \U309_0_/U12  ( .x(chainh[0]), .a(\net334[7] ), .b(\net284[7] ), .c(
        chain_ff_h[0]) );
    or3_4 \U309_1_/U12  ( .x(chainh[1]), .a(\net334[6] ), .b(\net284[6] ), .c(
        chain_ff_h[1]) );
    or3_4 \U309_3_/U12  ( .x(chainh[3]), .a(\net334[4] ), .b(\net284[4] ), .c(
        chain_ff_h[3]) );
    or3_4 \U309_5_/U12  ( .x(chainh[5]), .a(\net334[2] ), .b(\net284[2] ), .c(
        chain_ff_h[5]) );
    or3_4 \U309_6_/U12  ( .x(chainh[6]), .a(\net334[1] ), .b(\net284[1] ), .c(
        chain_ff_h[6]) );
    or3_4 \U309_7_/U12  ( .x(chainh[7]), .a(\net334[0] ), .b(\net284[0] ), .c(
        chain_ff_h[7]) );
    or3_4 \U310_0_/U12  ( .x(chainl[0]), .a(\net343[7] ), .b(\net288[7] ), .c(
        chainff_l[0]) );
    or3_4 \U310_1_/U12  ( .x(chainl[1]), .a(\net343[6] ), .b(\net288[6] ), .c(
        chainff_l[1]) );
    or3_4 \U310_2_/U12  ( .x(chainl[2]), .a(\net343[5] ), .b(\net288[5] ), .c(
        chainff_l[2]) );
    or3_4 \U310_4_/U12  ( .x(chainl[4]), .a(\net343[3] ), .b(\net288[3] ), .c(
        chainff_l[4]) );
    or3_4 \U310_5_/U12  ( .x(chainl[5]), .a(\net343[2] ), .b(\net288[2] ), .c(
        chainff_l[5]) );
    or3_4 \U310_6_/U12  ( .x(chainl[6]), .a(\net343[1] ), .b(\net288[1] ), .c(
        chainff_l[6]) );
    or3_4 \U310_7_/U12  ( .x(chainl[7]), .a(\net343[0] ), .b(\net288[0] ), .c(
        chainff_l[7]) );
    ao222_1 \U311/U37/U18/U1/U1  ( .x(ctrl_cd), .a(\U311/nz[0] ), .b(
        \U311/nz[1] ), .c(\U311/nz[0] ), .d(ctrl_cd), .e(\U311/nz[1] ), .f(
        ctrl_cd) );
    aoi222_1 \U311/U28/U30/U1  ( .x(\U311/x[3] ), .a(\net413[8] ), .b(
        \net413[9] ), .c(\net413[8] ), .d(\U311/U28/Z ), .e(\net413[9] ), .f(
        \U311/U28/Z ) );
    inv_1 \U311/U28/U30/Uinv  ( .x(\U311/U28/Z ), .a(\U311/x[3] ) );
    aoi222_1 \U311/U32/U30/U1  ( .x(\U311/x[0] ), .a(\net413[14] ), .b(
        \net413[15] ), .c(\net413[14] ), .d(\U311/U32/Z ), .e(\net413[15] ), 
        .f(\U311/U32/Z ) );
    inv_1 \U311/U32/U30/Uinv  ( .x(\U311/U32/Z ), .a(\U311/x[0] ) );
    aoi222_1 \U311/U20/U30/U1  ( .x(\U311/x[5] ), .a(\net413[4] ), .b(
        \net413[5] ), .c(\net413[4] ), .d(\U311/U20/Z ), .e(\net413[5] ), .f(
        \U311/U20/Z ) );
    inv_1 \U311/U20/U30/Uinv  ( .x(\U311/U20/Z ), .a(\U311/x[5] ) );
    aoi222_1 \U311/U29/U30/U1  ( .x(\U311/x[2] ), .a(\net413[10] ), .b(
        \net413[11] ), .c(\net413[10] ), .d(\U311/U29/Z ), .e(\net413[11] ), 
        .f(\U311/U29/Z ) );
    inv_1 \U311/U29/U30/Uinv  ( .x(\U311/U29/Z ), .a(\U311/x[2] ) );
    aoi222_1 \U311/U25/U30/U1  ( .x(\U311/x[7] ), .a(\net413[0] ), .b(
        \net413[1] ), .c(\net413[0] ), .d(\U311/U25/Z ), .e(\net413[1] ), .f(
        \U311/U25/Z ) );
    inv_1 \U311/U25/U30/Uinv  ( .x(\U311/U25/Z ), .a(\U311/x[7] ) );
    aoi222_1 \U311/U33/U30/U1  ( .x(\U311/y[0] ), .a(\U311/x[1] ), .b(
        \U311/x[0] ), .c(\U311/x[1] ), .d(\U311/U33/Z ), .e(\U311/x[0] ), .f(
        \U311/U33/Z ) );
    inv_1 \U311/U33/U30/Uinv  ( .x(\U311/U33/Z ), .a(\U311/y[0] ) );
    aoi222_1 \U311/U21/U30/U1  ( .x(\U311/y[2] ), .a(\U311/x[5] ), .b(
        \U311/x[4] ), .c(\U311/x[5] ), .d(\U311/U21/Z ), .e(\U311/x[4] ), .f(
        \U311/U21/Z ) );
    inv_1 \U311/U21/U30/Uinv  ( .x(\U311/U21/Z ), .a(\U311/y[2] ) );
    aoi222_1 \U311/U26/U30/U1  ( .x(\U311/x[6] ), .a(\net413[2] ), .b(
        \net413[3] ), .c(\net413[2] ), .d(\U311/U26/Z ), .e(\net413[3] ), .f(
        \U311/U26/Z ) );
    inv_1 \U311/U26/U30/Uinv  ( .x(\U311/U26/Z ), .a(\U311/x[6] ) );
    aoi222_1 \U311/U34/U30/U1  ( .x(\U311/nz[0] ), .a(\U311/y[1] ), .b(
        \U311/y[0] ), .c(\U311/y[1] ), .d(\U311/U34/Z ), .e(\U311/y[0] ), .f(
        \U311/U34/Z ) );
    inv_1 \U311/U34/U30/Uinv  ( .x(\U311/U34/Z ), .a(\U311/nz[0] ) );
    aoi222_1 \U311/U30/U30/U1  ( .x(\U311/y[1] ), .a(\U311/x[3] ), .b(
        \U311/x[2] ), .c(\U311/x[3] ), .d(\U311/U30/Z ), .e(\U311/x[2] ), .f(
        \U311/U30/Z ) );
    inv_1 \U311/U30/U30/Uinv  ( .x(\U311/U30/Z ), .a(\U311/y[1] ) );
    aoi222_1 \U311/U19/U30/U1  ( .x(\U311/x[4] ), .a(\net413[6] ), .b(
        \net413[7] ), .c(\net413[6] ), .d(\U311/U19/Z ), .e(\net413[7] ), .f(
        \U311/U19/Z ) );
    inv_1 \U311/U19/U30/Uinv  ( .x(\U311/U19/Z ), .a(\U311/x[4] ) );
    aoi222_1 \U311/U27/U30/U1  ( .x(\U311/y[3] ), .a(\U311/x[7] ), .b(
        \U311/x[6] ), .c(\U311/x[7] ), .d(\U311/U27/Z ), .e(\U311/x[6] ), .f(
        \U311/U27/Z ) );
    inv_1 \U311/U27/U30/Uinv  ( .x(\U311/U27/Z ), .a(\U311/y[3] ) );
    aoi222_1 \U311/U35/U30/U1  ( .x(\U311/nz[1] ), .a(\U311/y[3] ), .b(
        \U311/y[2] ), .c(\U311/y[3] ), .d(\U311/U35/Z ), .e(\U311/y[2] ), .f(
        \U311/U35/Z ) );
    inv_1 \U311/U35/U30/Uinv  ( .x(\U311/U35/Z ), .a(\U311/nz[1] ) );
    aoi222_1 \U311/U31/U30/U1  ( .x(\U311/x[1] ), .a(\net413[12] ), .b(
        \net413[13] ), .c(\net413[12] ), .d(\U311/U31/Z ), .e(\net413[13] ), 
        .f(\U311/U31/Z ) );
    inv_1 \U311/U31/U30/Uinv  ( .x(\U311/U31/Z ), .a(\U311/x[1] ) );
    aoi21_1 \U151/U30/U1/U1  ( .x(net407), .a(\U151/Z ), .b(chainff_ack), .c(
        net332) );
    inv_1 \U151/U30/U1/U2  ( .x(\U151/Z ), .a(net407) );
    ao222_1 \U324/U18/U1/U1  ( .x(hdrack), .a(ctrl_cd), .b(net383), .c(ctrl_cd
        ), .d(hdrack), .e(net383), .f(hdrack) );
    ao222_1 \U244/U18/U1/U1  ( .x(donotify), .a(done_hdr), .b(\hdr[17] ), .c(
        done_hdr), .d(donotify), .e(\hdr[17] ), .f(donotify) );
    ao222_1 \U260/U18/U1/U1  ( .x(net362), .a(net337), .b(\hdr[1] ), .c(net337
        ), .d(net362), .e(\hdr[1] ), .f(net362) );
    ao222_1 \U296/U18/U1/U1  ( .x(done_accept), .a(done_eop), .b(notify_accept
        ), .c(done_eop), .d(done_accept), .e(notify_accept), .f(done_accept)
         );
    ao222_1 \U261/U18/U1/U1  ( .x(net359), .a(net340), .b(\hdr[1] ), .c(net340
        ), .d(net359), .e(\hdr[1] ), .f(net359) );
    ao222_1 \U316/U18/U1/U1  ( .x(done_pl), .a(net364), .b(routeack), .c(
        net364), .d(done_pl), .e(routeack), .f(done_pl) );
    ao31_1 \U319/U21/U1/aoi  ( .x(\U319/U21/U1/loop ), .a(\hdr[1] ), .b(
        done_hdr), .c(rnw_h), .d(read_req) );
    oa21_1 \U319/U21/U1/outGate  ( .x(read_req), .a(\hdr[1] ), .b(done_hdr), 
        .c(\U319/U21/U1/loop ) );
    ao31_1 \U323/U21/U1/aoi  ( .x(\U323/U21/U1/loop ), .a(done_eop), .b(
        notify_defer), .c(ctrl_cd), .d(done_defer) );
    oa21_1 \U323/U21/U1/outGate  ( .x(done_defer), .a(done_eop), .b(
        notify_defer), .c(\U323/U21/U1/loop ) );
    ao31_1 \U320/U21/U1/aoi  ( .x(\U320/U21/U1/loop ), .a(\hdr[1] ), .b(
        done_hdr), .c(rnw_l), .d(dowrite) );
    oa21_1 \U320/U21/U1/outGate  ( .x(dowrite), .a(\hdr[1] ), .b(done_hdr), 
        .c(\U320/U21/U1/loop ) );
    ao31_1 \U321/U21/U1/aoi  ( .x(\U321/U21/U1/loop ), .a(read_req), .b(
        done_eop), .c(ctrl_cd), .d(done_read) );
    oa21_1 \U321/U21/U1/outGate  ( .x(done_read), .a(read_req), .b(done_eop), 
        .c(\U321/U21/U1/loop ) );
    ao31_1 \U322/U21/U1/aoi  ( .x(\U322/U21/U1/loop ), .a(dowrite), .b(
        done_eop), .c(ctrl_cd), .d(done_write) );
    oa21_1 \U322/U21/U1/outGate  ( .x(done_write), .a(dowrite), .b(done_eop), 
        .c(\U322/U21/U1/loop ) );
    nor2_2 \U210/U1703/U6  ( .x(done_hdr), .a(\U210/drivemonitor ), .b(
        \U210/naa ) );
    inv_2 \U210/U1699/U3  ( .x(\U210/net2 ), .a(\U210/net3 ) );
    and2_4 \U210/U2_0_/U8  ( .x(\drive_l[0] ), .a(net0230), .b(\U210/net2 ) );
    and2_4 \U210/U2_1_/U8  ( .x(\drive_l[1] ), .a(net0230), .b(\U210/net2 ) );
    inv_1 \U210/U1701/U3  ( .x(\U210/naa ), .a(\U210/bdone ) );
    ao222_1 \U210/U13/U18/U1/U1  ( .x(\U210/drivemonitor ), .a(\drive_l[1] ), 
        .b(\drive_l[0] ), .c(\drive_l[1] ), .d(\U210/drivemonitor ), .e(
        \drive_l[0] ), .f(\U210/drivemonitor ) );
    aoi21_1 \U210/U1702/U30/U1/U1  ( .x(\U210/bdone ), .a(\U210/U1702/Z ), .b(
        chainff_ack), .c(\U210/net2 ) );
    inv_1 \U210/U1702/U30/U1/U2  ( .x(\U210/U1702/Z ), .a(\U210/bdone ) );
    ao23_1 \U210/U1693/U21/U1/U1  ( .x(\U210/net3 ), .a(net0230), .b(
        \U210/net3 ), .c(net0230), .d(\U210/drivemonitor ), .e(chainff_ack) );
    nor2_2 \I0/U1703/U6  ( .x(net0230), .a(\I0/drivemonitor ), .b(\I0/naa ) );
    inv_2 \I0/U1699/U3  ( .x(\I0/net2 ), .a(\I0/net3 ) );
    and2_4 \I0/U2_0_/U8  ( .x(\drive_h[0] ), .a(net407), .b(\I0/net2 ) );
    and2_4 \I0/U2_1_/U8  ( .x(\drive_h[1] ), .a(net407), .b(\I0/net2 ) );
    inv_1 \I0/U1701/U3  ( .x(\I0/naa ), .a(\I0/bdone ) );
    ao222_1 \I0/U13/U18/U1/U1  ( .x(\I0/drivemonitor ), .a(\drive_h[1] ), .b(
        \drive_h[0] ), .c(\drive_h[1] ), .d(\I0/drivemonitor ), .e(
        \drive_h[0] ), .f(\I0/drivemonitor ) );
    aoi21_1 \I0/U1702/U30/U1/U1  ( .x(\I0/bdone ), .a(\I0/U1702/Z ), .b(
        chainff_ack), .c(\I0/net2 ) );
    inv_1 \I0/U1702/U30/U1/U2  ( .x(\I0/U1702/Z ), .a(\I0/bdone ) );
    ao23_1 \I0/U1693/U21/U1/U1  ( .x(\I0/net3 ), .a(net407), .b(\I0/net3 ), 
        .c(net407), .d(\I0/drivemonitor ), .e(chainff_ack) );
    buf_3 U1 ( .x(chainff_ack), .a(chainack) );
    or2_1 U2 ( .x(chainh[4]), .a(chain_ff_h[4]), .b(\net284[3] ) );
    or2_1 U3 ( .x(chainh[2]), .a(chain_ff_h[2]), .b(\net284[5] ) );
    or2_1 U4 ( .x(chainl[3]), .a(chainff_l[3]), .b(\net288[4] ) );
endmodule


module chain_dr2fr_byte_3 ( eop_ack, ia, o, eop, ih, il, nReset, noa );
output [4:0] o;
input  [7:0] ih;
input  [7:0] il;
input  eop, nReset, noa;
output eop_ack, ia;
    wire eop_ack_wire, nbReset, eop_pass, nxa, naa, nlowack, \twobitack[0] , 
        \twobitack[1] , nhighack, \twobitack[2] , \twobitack[3] , \U1018/Z , 
        \U1270/net189 , \U1270/net192 , \U1270/net191 , net199, \U1270/net190 , 
        \U1270/U1141/Z , \U1268/net189 , \U1268/net192 , \U1268/net191 , 
        net194, \U1268/net190 , \U1268/U1141/Z , \U1224/nack[0] , \x[3] , 
        \x[2] , \U1224/nack[1] , \x[1] , \U1224/net4 , \x[0] , 
        \U1224/U1125/U28/U1/clr , asel, \U1224/U1125/U28/U1/set , 
        \U1224/U1122/U28/U1/clr , csel, nca, \U1224/U1122/U28/U1/set , 
        \U1224/U916_0_/U25/U1/clr , \a[0] , \c[0] , \U1224/U916_0_/U25/U1/ob , 
        \U1224/U916_1_/U25/U1/clr , \a[1] , \c[1] , \U1224/U916_1_/U25/U1/ob , 
        \U1224/U916_2_/U25/U1/clr , \a[2] , \c[2] , \U1224/U916_2_/U25/U1/ob , 
        \U1224/U916_3_/U25/U1/clr , \a[3] , \c[3] , \U1224/U916_3_/U25/U1/ob , 
        \U1209/nack[0] , \U1209/nack[1] , \U1209/net4 , 
        \U1209/U1125/U28/U1/clr , xsel, \U1209/U1125/U28/U1/set , 
        \U1209/U1122/U28/U1/clr , ysel, nyla, \U1209/U1122/U28/U1/set , 
        \U1209/U916_0_/U25/U1/clr , \yl[0] , \U1209/U916_0_/U25/U1/ob , 
        \U1209/U916_1_/U25/U1/clr , \yl[1] , \U1209/U916_1_/U25/U1/ob , 
        \U1209/U916_2_/U25/U1/clr , \yl[2] , \U1209/U916_2_/U25/U1/ob , 
        \U1209/U916_3_/U25/U1/clr , \yl[3] , \U1209/U916_3_/U25/U1/ob , 
        \U1213/nack[0] , \y[3] , \y[2] , \U1213/nack[1] , \y[1] , \U1213/net4 , 
        \y[0] , \U1213/U1125/U28/U1/clr , bsel, nba, \U1213/U1125/U28/U1/set , 
        \U1213/U1122/U28/U1/clr , dsel, nda, \U1213/U1122/U28/U1/set , 
        \U1213/U916_0_/U25/U1/clr , nya, \b[0] , \d[0] , 
        \U1213/U916_0_/U25/U1/ob , \U1213/U916_1_/U25/U1/clr , \b[1] , \d[1] , 
        \U1213/U916_1_/U25/U1/ob , \U1213/U916_2_/U25/U1/clr , \b[2] , \d[2] , 
        \U1213/U916_2_/U25/U1/ob , \U1213/U916_3_/U25/U1/clr , \b[3] , \d[3] , 
        \U1213/U916_3_/U25/U1/ob , \cdh[0] , \cdh[1] , \cdl[0] , \cdl[1] , 
        \cdh[2] , \cdh[3] , \cdl[2] , \cdl[3] , cg, \U1296/ng , net195, 
        \U1296/U1384/Z , \U1296/U1386/U25/U1/clr , \U1296/U1386/U25/U1/ob , dg, 
        \U1298/ng , net193, \U1298/U1384/Z , \U1298/U1386/U25/U1/clr , 
        \U1298/U1386/U25/U1/ob , bg, \U1306/ng , \U1306/U1384/Z , 
        \U1306/U1386/U25/U1/clr , \U1306/U1386/U25/U1/ob , ag, \U1295/ng , 
        \U1295/U1384/Z , \U1295/U1386/U25/U1/clr , \U1295/U1386/U25/U1/ob , 
        \U1297/s , \U1297/r , \U1297/nback , \U1297/naack , \U1297/reset , 
        \U1297/U1128/U28/U1/clr , \U1297/U1128/U28/U1/set , 
        \U1297/U1127/U28/U1/clr , \U1297/U1127/U28/U1/set , \U1300/s , 
        \U1300/r , \U1300/nback , \U1300/naack , \U1300/reset , 
        \U1300/U1128/U28/U1/clr , \U1300/U1128/U28/U1/set , 
        \U1300/U1127/U28/U1/clr , \U1300/U1127/U28/U1/set , 
        \U1289/U1150/U28/U1/clr , \U1289/bnreset , \U1289/U1150/U28/U1/set , 
        \U1289/U1152/U28/U1/clr , \U1289/U1152/U28/U1/set , 
        \U1289/U1149/U28/U1/clr , \U1289/U1149/U28/U1/set , 
        \U1289/U1151/U28/U1/clr , \U1289/U1151/U28/U1/set , 
        \U1289/U1148/net189 , \U1289/U1148/net192 , \U1289/U1148/net191 , 
        \U1289/U1148/net190 , \U1289/U1148/U1141/Z , \U1271/U1150/U28/U1/clr , 
        \U1271/bnreset , \U1271/U1150/U28/U1/set , \U1271/U1152/U28/U1/clr , 
        \U1271/U1152/U28/U1/set , \U1271/U1149/U28/U1/clr , 
        \U1271/U1149/U28/U1/set , \U1271/U1151/U28/U1/clr , 
        \U1271/U1151/U28/U1/set , \U1271/U1148/net189 , \U1271/U1148/net192 , 
        \U1271/U1148/net191 , \U1271/U1148/net190 , \U1271/U1148/U1141/Z , 
        \U1225/s , \U1225/r , \U1225/nback , \U1225/naack , \U1225/reset , 
        \U1308/nack[1] , \U1308/nack[0] ;
    assign eop_ack = eop_ack_wire;
    assign o[4] = eop_ack_wire;
    buf_2 U1231 ( .x(nbReset), .a(nReset) );
    and3_1 \U1194/U9  ( .x(eop_pass), .a(nxa), .b(naa), .c(eop) );
    ao222_1 \U1301/U18/U1/U1  ( .x(nlowack), .a(\twobitack[0] ), .b(
        \twobitack[1] ), .c(\twobitack[0] ), .d(nlowack), .e(\twobitack[1] ), 
        .f(nlowack) );
    ao222_1 \U1302/U18/U1/U1  ( .x(nhighack), .a(\twobitack[2] ), .b(
        \twobitack[3] ), .c(\twobitack[2] ), .d(nhighack), .e(\twobitack[3] ), 
        .f(nhighack) );
    aoi222_1 \U1018/U30/U1  ( .x(ia), .a(nhighack), .b(nlowack), .c(nhighack), 
        .d(\U1018/Z ), .e(nlowack), .f(\U1018/Z ) );
    inv_1 \U1018/U30/Uinv  ( .x(\U1018/Z ), .a(ia) );
    ao222_2 \U1038/U19/U1/U1  ( .x(eop_ack_wire), .a(eop_pass), .b(noa), .c(
        eop_pass), .d(eop_ack_wire), .e(noa), .f(eop_ack_wire) );
    inv_1 \U1270/U1147/U3  ( .x(\U1270/net189 ), .a(nbReset) );
    nor2_1 \U1270/U582/U5  ( .x(\U1270/net192 ), .a(il[4]), .b(ih[4]) );
    nor2_1 \U1270/U580/U5  ( .x(\U1270/net191 ), .a(il[5]), .b(ih[5]) );
    nor2_2 \U1270/U1146/U6  ( .x(net199), .a(\U1270/net190 ), .b(
        \U1270/net189 ) );
    aoi222_1 \U1270/U1141/U30/U1  ( .x(\U1270/net190 ), .a(\U1270/net191 ), 
        .b(\U1270/net192 ), .c(\U1270/net191 ), .d(\U1270/U1141/Z ), .e(
        \U1270/net192 ), .f(\U1270/U1141/Z ) );
    inv_1 \U1270/U1141/U30/Uinv  ( .x(\U1270/U1141/Z ), .a(\U1270/net190 ) );
    inv_1 \U1268/U1147/U3  ( .x(\U1268/net189 ), .a(nbReset) );
    nor2_1 \U1268/U582/U5  ( .x(\U1268/net192 ), .a(il[6]), .b(ih[6]) );
    nor2_1 \U1268/U580/U5  ( .x(\U1268/net191 ), .a(il[7]), .b(ih[7]) );
    nor2_2 \U1268/U1146/U6  ( .x(net194), .a(\U1268/net190 ), .b(
        \U1268/net189 ) );
    aoi222_1 \U1268/U1141/U30/U1  ( .x(\U1268/net190 ), .a(\U1268/net191 ), 
        .b(\U1268/net192 ), .c(\U1268/net191 ), .d(\U1268/U1141/Z ), .e(
        \U1268/net192 ), .f(\U1268/U1141/Z ) );
    inv_1 \U1268/U1141/U30/Uinv  ( .x(\U1268/U1141/Z ), .a(\U1268/net190 ) );
    nor2_1 \U1224/U1128/U5  ( .x(\U1224/nack[0] ), .a(\x[3] ), .b(\x[2] ) );
    nor3_1 \U1224/U1127/U7  ( .x(\U1224/nack[1] ), .a(\x[1] ), .b(\U1224/net4 
        ), .c(\x[0] ) );
    inv_1 \U1224/U907/U3  ( .x(\U1224/net4 ), .a(nbReset) );
    aoai211_1 \U1224/U1125/U28/U1/U1  ( .x(\U1224/U1125/U28/U1/clr ), .a(
        \U1224/nack[1] ), .b(\U1224/nack[0] ), .c(asel), .d(naa) );
    nand3_1 \U1224/U1125/U28/U1/U2  ( .x(\U1224/U1125/U28/U1/set ), .a(asel), 
        .b(\U1224/nack[1] ), .c(\U1224/nack[0] ) );
    nand2_2 \U1224/U1125/U28/U1/U3  ( .x(naa), .a(\U1224/U1125/U28/U1/clr ), 
        .b(\U1224/U1125/U28/U1/set ) );
    aoai211_1 \U1224/U1122/U28/U1/U1  ( .x(\U1224/U1122/U28/U1/clr ), .a(
        \U1224/nack[0] ), .b(\U1224/nack[1] ), .c(csel), .d(nca) );
    nand3_1 \U1224/U1122/U28/U1/U2  ( .x(\U1224/U1122/U28/U1/set ), .a(csel), 
        .b(\U1224/nack[0] ), .c(\U1224/nack[1] ) );
    nand2_2 \U1224/U1122/U28/U1/U3  ( .x(nca), .a(\U1224/U1122/U28/U1/clr ), 
        .b(\U1224/U1122/U28/U1/set ) );
    oa31_1 \U1224/U916_0_/U25/U1/Uclr  ( .x(\U1224/U916_0_/U25/U1/clr ), .a(
        nxa), .b(\a[0] ), .c(\c[0] ), .d(\x[0] ) );
    oaoi211_1 \U1224/U916_0_/U25/U1/Uaoi  ( .x(\U1224/U916_0_/U25/U1/ob ), .a(
        \a[0] ), .b(\c[0] ), .c(nxa), .d(\U1224/U916_0_/U25/U1/clr ) );
    inv_2 \U1224/U916_0_/U25/U1/Ui  ( .x(\x[0] ), .a(\U1224/U916_0_/U25/U1/ob 
        ) );
    oa31_1 \U1224/U916_1_/U25/U1/Uclr  ( .x(\U1224/U916_1_/U25/U1/clr ), .a(
        nxa), .b(\a[1] ), .c(\c[1] ), .d(\x[1] ) );
    oaoi211_1 \U1224/U916_1_/U25/U1/Uaoi  ( .x(\U1224/U916_1_/U25/U1/ob ), .a(
        \a[1] ), .b(\c[1] ), .c(nxa), .d(\U1224/U916_1_/U25/U1/clr ) );
    inv_2 \U1224/U916_1_/U25/U1/Ui  ( .x(\x[1] ), .a(\U1224/U916_1_/U25/U1/ob 
        ) );
    oa31_1 \U1224/U916_2_/U25/U1/Uclr  ( .x(\U1224/U916_2_/U25/U1/clr ), .a(
        nxa), .b(\a[2] ), .c(\c[2] ), .d(\x[2] ) );
    oaoi211_1 \U1224/U916_2_/U25/U1/Uaoi  ( .x(\U1224/U916_2_/U25/U1/ob ), .a(
        \a[2] ), .b(\c[2] ), .c(nxa), .d(\U1224/U916_2_/U25/U1/clr ) );
    inv_2 \U1224/U916_2_/U25/U1/Ui  ( .x(\x[2] ), .a(\U1224/U916_2_/U25/U1/ob 
        ) );
    oa31_1 \U1224/U916_3_/U25/U1/Uclr  ( .x(\U1224/U916_3_/U25/U1/clr ), .a(
        nxa), .b(\a[3] ), .c(\c[3] ), .d(\x[3] ) );
    oaoi211_1 \U1224/U916_3_/U25/U1/Uaoi  ( .x(\U1224/U916_3_/U25/U1/ob ), .a(
        \a[3] ), .b(\c[3] ), .c(nxa), .d(\U1224/U916_3_/U25/U1/clr ) );
    inv_2 \U1224/U916_3_/U25/U1/Ui  ( .x(\x[3] ), .a(\U1224/U916_3_/U25/U1/ob 
        ) );
    nor2_1 \U1209/U1128/U5  ( .x(\U1209/nack[0] ), .a(o[3]), .b(o[2]) );
    nor3_1 \U1209/U1127/U7  ( .x(\U1209/nack[1] ), .a(o[1]), .b(\U1209/net4 ), 
        .c(o[0]) );
    inv_1 \U1209/U907/U3  ( .x(\U1209/net4 ), .a(nbReset) );
    aoai211_1 \U1209/U1125/U28/U1/U1  ( .x(\U1209/U1125/U28/U1/clr ), .a(
        \U1209/nack[1] ), .b(\U1209/nack[0] ), .c(xsel), .d(nxa) );
    nand3_1 \U1209/U1125/U28/U1/U2  ( .x(\U1209/U1125/U28/U1/set ), .a(xsel), 
        .b(\U1209/nack[1] ), .c(\U1209/nack[0] ) );
    nand2_2 \U1209/U1125/U28/U1/U3  ( .x(nxa), .a(\U1209/U1125/U28/U1/clr ), 
        .b(\U1209/U1125/U28/U1/set ) );
    aoai211_1 \U1209/U1122/U28/U1/U1  ( .x(\U1209/U1122/U28/U1/clr ), .a(
        \U1209/nack[0] ), .b(\U1209/nack[1] ), .c(ysel), .d(nyla) );
    nand3_1 \U1209/U1122/U28/U1/U2  ( .x(\U1209/U1122/U28/U1/set ), .a(ysel), 
        .b(\U1209/nack[0] ), .c(\U1209/nack[1] ) );
    nand2_2 \U1209/U1122/U28/U1/U3  ( .x(nyla), .a(\U1209/U1122/U28/U1/clr ), 
        .b(\U1209/U1122/U28/U1/set ) );
    oa31_1 \U1209/U916_0_/U25/U1/Uclr  ( .x(\U1209/U916_0_/U25/U1/clr ), .a(
        noa), .b(\x[0] ), .c(\yl[0] ), .d(o[0]) );
    oaoi211_1 \U1209/U916_0_/U25/U1/Uaoi  ( .x(\U1209/U916_0_/U25/U1/ob ), .a(
        \x[0] ), .b(\yl[0] ), .c(noa), .d(\U1209/U916_0_/U25/U1/clr ) );
    inv_2 \U1209/U916_0_/U25/U1/Ui  ( .x(o[0]), .a(\U1209/U916_0_/U25/U1/ob )
         );
    oa31_1 \U1209/U916_1_/U25/U1/Uclr  ( .x(\U1209/U916_1_/U25/U1/clr ), .a(
        noa), .b(\x[1] ), .c(\yl[1] ), .d(o[1]) );
    oaoi211_1 \U1209/U916_1_/U25/U1/Uaoi  ( .x(\U1209/U916_1_/U25/U1/ob ), .a(
        \x[1] ), .b(\yl[1] ), .c(noa), .d(\U1209/U916_1_/U25/U1/clr ) );
    inv_2 \U1209/U916_1_/U25/U1/Ui  ( .x(o[1]), .a(\U1209/U916_1_/U25/U1/ob )
         );
    oa31_1 \U1209/U916_2_/U25/U1/Uclr  ( .x(\U1209/U916_2_/U25/U1/clr ), .a(
        noa), .b(\x[2] ), .c(\yl[2] ), .d(o[2]) );
    oaoi211_1 \U1209/U916_2_/U25/U1/Uaoi  ( .x(\U1209/U916_2_/U25/U1/ob ), .a(
        \x[2] ), .b(\yl[2] ), .c(noa), .d(\U1209/U916_2_/U25/U1/clr ) );
    inv_2 \U1209/U916_2_/U25/U1/Ui  ( .x(o[2]), .a(\U1209/U916_2_/U25/U1/ob )
         );
    oa31_1 \U1209/U916_3_/U25/U1/Uclr  ( .x(\U1209/U916_3_/U25/U1/clr ), .a(
        noa), .b(\x[3] ), .c(\yl[3] ), .d(o[3]) );
    oaoi211_1 \U1209/U916_3_/U25/U1/Uaoi  ( .x(\U1209/U916_3_/U25/U1/ob ), .a(
        \x[3] ), .b(\yl[3] ), .c(noa), .d(\U1209/U916_3_/U25/U1/clr ) );
    inv_2 \U1209/U916_3_/U25/U1/Ui  ( .x(o[3]), .a(\U1209/U916_3_/U25/U1/ob )
         );
    nor2_1 \U1213/U1128/U5  ( .x(\U1213/nack[0] ), .a(\y[3] ), .b(\y[2] ) );
    nor3_1 \U1213/U1127/U7  ( .x(\U1213/nack[1] ), .a(\y[1] ), .b(\U1213/net4 
        ), .c(\y[0] ) );
    inv_1 \U1213/U907/U3  ( .x(\U1213/net4 ), .a(nbReset) );
    aoai211_1 \U1213/U1125/U28/U1/U1  ( .x(\U1213/U1125/U28/U1/clr ), .a(
        \U1213/nack[1] ), .b(\U1213/nack[0] ), .c(bsel), .d(nba) );
    nand3_1 \U1213/U1125/U28/U1/U2  ( .x(\U1213/U1125/U28/U1/set ), .a(bsel), 
        .b(\U1213/nack[1] ), .c(\U1213/nack[0] ) );
    nand2_2 \U1213/U1125/U28/U1/U3  ( .x(nba), .a(\U1213/U1125/U28/U1/clr ), 
        .b(\U1213/U1125/U28/U1/set ) );
    aoai211_1 \U1213/U1122/U28/U1/U1  ( .x(\U1213/U1122/U28/U1/clr ), .a(
        \U1213/nack[0] ), .b(\U1213/nack[1] ), .c(dsel), .d(nda) );
    nand3_1 \U1213/U1122/U28/U1/U2  ( .x(\U1213/U1122/U28/U1/set ), .a(dsel), 
        .b(\U1213/nack[0] ), .c(\U1213/nack[1] ) );
    nand2_2 \U1213/U1122/U28/U1/U3  ( .x(nda), .a(\U1213/U1122/U28/U1/clr ), 
        .b(\U1213/U1122/U28/U1/set ) );
    oa31_1 \U1213/U916_0_/U25/U1/Uclr  ( .x(\U1213/U916_0_/U25/U1/clr ), .a(
        nya), .b(\b[0] ), .c(\d[0] ), .d(\y[0] ) );
    oaoi211_1 \U1213/U916_0_/U25/U1/Uaoi  ( .x(\U1213/U916_0_/U25/U1/ob ), .a(
        \b[0] ), .b(\d[0] ), .c(nya), .d(\U1213/U916_0_/U25/U1/clr ) );
    inv_2 \U1213/U916_0_/U25/U1/Ui  ( .x(\y[0] ), .a(\U1213/U916_0_/U25/U1/ob 
        ) );
    oa31_1 \U1213/U916_1_/U25/U1/Uclr  ( .x(\U1213/U916_1_/U25/U1/clr ), .a(
        nya), .b(\b[1] ), .c(\d[1] ), .d(\y[1] ) );
    oaoi211_1 \U1213/U916_1_/U25/U1/Uaoi  ( .x(\U1213/U916_1_/U25/U1/ob ), .a(
        \b[1] ), .b(\d[1] ), .c(nya), .d(\U1213/U916_1_/U25/U1/clr ) );
    inv_2 \U1213/U916_1_/U25/U1/Ui  ( .x(\y[1] ), .a(\U1213/U916_1_/U25/U1/ob 
        ) );
    oa31_1 \U1213/U916_2_/U25/U1/Uclr  ( .x(\U1213/U916_2_/U25/U1/clr ), .a(
        nya), .b(\b[2] ), .c(\d[2] ), .d(\y[2] ) );
    oaoi211_1 \U1213/U916_2_/U25/U1/Uaoi  ( .x(\U1213/U916_2_/U25/U1/ob ), .a(
        \b[2] ), .b(\d[2] ), .c(nya), .d(\U1213/U916_2_/U25/U1/clr ) );
    inv_2 \U1213/U916_2_/U25/U1/Ui  ( .x(\y[2] ), .a(\U1213/U916_2_/U25/U1/ob 
        ) );
    oa31_1 \U1213/U916_3_/U25/U1/Uclr  ( .x(\U1213/U916_3_/U25/U1/clr ), .a(
        nya), .b(\b[3] ), .c(\d[3] ), .d(\y[3] ) );
    oaoi211_1 \U1213/U916_3_/U25/U1/Uaoi  ( .x(\U1213/U916_3_/U25/U1/ob ), .a(
        \b[3] ), .b(\d[3] ), .c(nya), .d(\U1213/U916_3_/U25/U1/clr ) );
    inv_2 \U1213/U916_3_/U25/U1/Ui  ( .x(\y[3] ), .a(\U1213/U916_3_/U25/U1/ob 
        ) );
    and3_2 \U1210/U1138/U9  ( .x(\d[3] ), .a(\cdh[0] ), .b(nda), .c(\cdh[1] )
         );
    and3_2 \U1210/U1137/U9  ( .x(\d[2] ), .a(\cdl[0] ), .b(nda), .c(\cdh[1] )
         );
    and3_2 \U1210/U1139/U9  ( .x(\d[1] ), .a(\cdh[0] ), .b(nda), .c(\cdl[1] )
         );
    and3_2 \U1210/U1136/U9  ( .x(\d[0] ), .a(\cdl[0] ), .b(nda), .c(\cdl[1] )
         );
    and3_2 \U1162/U1138/U9  ( .x(\a[3] ), .a(ih[6]), .b(naa), .c(ih[7]) );
    and3_2 \U1162/U1137/U9  ( .x(\a[2] ), .a(il[6]), .b(naa), .c(ih[7]) );
    and3_2 \U1162/U1139/U9  ( .x(\a[1] ), .a(ih[6]), .b(naa), .c(il[7]) );
    and3_2 \U1162/U1136/U9  ( .x(\a[0] ), .a(il[6]), .b(naa), .c(il[7]) );
    and3_2 \U1211/U1138/U9  ( .x(\b[3] ), .a(ih[4]), .b(nba), .c(ih[5]) );
    and3_2 \U1211/U1137/U9  ( .x(\b[2] ), .a(il[4]), .b(nba), .c(ih[5]) );
    and3_2 \U1211/U1139/U9  ( .x(\b[1] ), .a(ih[4]), .b(nba), .c(il[5]) );
    and3_2 \U1211/U1136/U9  ( .x(\b[0] ), .a(il[4]), .b(nba), .c(il[5]) );
    and3_2 \U1163/U1138/U9  ( .x(\c[3] ), .a(\cdh[2] ), .b(nca), .c(\cdh[3] )
         );
    and3_2 \U1163/U1137/U9  ( .x(\c[2] ), .a(\cdl[2] ), .b(nca), .c(\cdh[3] )
         );
    and3_2 \U1163/U1139/U9  ( .x(\c[1] ), .a(\cdh[2] ), .b(nca), .c(\cdl[3] )
         );
    and3_2 \U1163/U1136/U9  ( .x(\c[0] ), .a(\cdl[2] ), .b(nca), .c(\cdl[3] )
         );
    and2_1 \U1296/U1385/U8  ( .x(cg), .a(nbReset), .b(\U1296/ng ) );
    aoi222_1 \U1296/U1384/U30/U1  ( .x(\U1296/ng ), .a(nca), .b(net195), .c(
        nca), .d(\U1296/U1384/Z ), .e(net195), .f(\U1296/U1384/Z ) );
    inv_1 \U1296/U1384/U30/Uinv  ( .x(\U1296/U1384/Z ), .a(\U1296/ng ) );
    oa31_1 \U1296/U1386/U25/U1/Uclr  ( .x(\U1296/U1386/U25/U1/clr ), .a(
        \twobitack[2] ), .b(cg), .c(nca), .d(net195) );
    oaoi211_1 \U1296/U1386/U25/U1/Uaoi  ( .x(\U1296/U1386/U25/U1/ob ), .a(cg), 
        .b(nca), .c(\twobitack[2] ), .d(\U1296/U1386/U25/U1/clr ) );
    inv_2 \U1296/U1386/U25/U1/Ui  ( .x(net195), .a(\U1296/U1386/U25/U1/ob ) );
    and2_1 \U1298/U1385/U8  ( .x(dg), .a(nbReset), .b(\U1298/ng ) );
    aoi222_1 \U1298/U1384/U30/U1  ( .x(\U1298/ng ), .a(nda), .b(net193), .c(
        nda), .d(\U1298/U1384/Z ), .e(net193), .f(\U1298/U1384/Z ) );
    inv_1 \U1298/U1384/U30/Uinv  ( .x(\U1298/U1384/Z ), .a(\U1298/ng ) );
    oa31_1 \U1298/U1386/U25/U1/Uclr  ( .x(\U1298/U1386/U25/U1/clr ), .a(
        \twobitack[0] ), .b(dg), .c(nda), .d(net193) );
    oaoi211_1 \U1298/U1386/U25/U1/Uaoi  ( .x(\U1298/U1386/U25/U1/ob ), .a(dg), 
        .b(nda), .c(\twobitack[0] ), .d(\U1298/U1386/U25/U1/clr ) );
    inv_2 \U1298/U1386/U25/U1/Ui  ( .x(net193), .a(\U1298/U1386/U25/U1/ob ) );
    and2_1 \U1306/U1385/U8  ( .x(bg), .a(nbReset), .b(\U1306/ng ) );
    aoi222_1 \U1306/U1384/U30/U1  ( .x(\U1306/ng ), .a(nba), .b(\twobitack[1] 
        ), .c(nba), .d(\U1306/U1384/Z ), .e(\twobitack[1] ), .f(
        \U1306/U1384/Z ) );
    inv_1 \U1306/U1384/U30/Uinv  ( .x(\U1306/U1384/Z ), .a(\U1306/ng ) );
    oa31_1 \U1306/U1386/U25/U1/Uclr  ( .x(\U1306/U1386/U25/U1/clr ), .a(net199
        ), .b(bg), .c(nba), .d(\twobitack[1] ) );
    oaoi211_1 \U1306/U1386/U25/U1/Uaoi  ( .x(\U1306/U1386/U25/U1/ob ), .a(bg), 
        .b(nba), .c(net199), .d(\U1306/U1386/U25/U1/clr ) );
    inv_2 \U1306/U1386/U25/U1/Ui  ( .x(\twobitack[1] ), .a(
        \U1306/U1386/U25/U1/ob ) );
    and2_1 \U1295/U1385/U8  ( .x(ag), .a(nbReset), .b(\U1295/ng ) );
    aoi222_1 \U1295/U1384/U30/U1  ( .x(\U1295/ng ), .a(naa), .b(\twobitack[3] 
        ), .c(naa), .d(\U1295/U1384/Z ), .e(\twobitack[3] ), .f(
        \U1295/U1384/Z ) );
    inv_1 \U1295/U1384/U30/Uinv  ( .x(\U1295/U1384/Z ), .a(\U1295/ng ) );
    oa31_1 \U1295/U1386/U25/U1/Uclr  ( .x(\U1295/U1386/U25/U1/clr ), .a(net194
        ), .b(ag), .c(naa), .d(\twobitack[3] ) );
    oaoi211_1 \U1295/U1386/U25/U1/Uaoi  ( .x(\U1295/U1386/U25/U1/ob ), .a(ag), 
        .b(naa), .c(net194), .d(\U1295/U1386/U25/U1/clr ) );
    inv_2 \U1295/U1386/U25/U1/Ui  ( .x(\twobitack[3] ), .a(
        \U1295/U1386/U25/U1/ob ) );
    nand2_1 \U1297/U1131/U5  ( .x(\U1297/s ), .a(\U1297/r ), .b(\U1297/nback )
         );
    nand2_1 \U1297/U1103/U5  ( .x(\U1297/r ), .a(\U1297/naack ), .b(\U1297/s )
         );
    inv_1 \U1297/U1111/U3  ( .x(\U1297/reset ), .a(nbReset) );
    inv_1 \U1297/U1112/U3  ( .x(\U1297/naack ), .a(naa) );
    nor2_1 \U1297/U1130/U5  ( .x(\U1297/nback ), .a(nca), .b(\U1297/reset ) );
    aoai211_1 \U1297/U1128/U28/U1/U1  ( .x(\U1297/U1128/U28/U1/clr ), .a(
        \U1297/r ), .b(\U1297/naack ), .c(cg), .d(csel) );
    nand3_1 \U1297/U1128/U28/U1/U2  ( .x(\U1297/U1128/U28/U1/set ), .a(cg), 
        .b(\U1297/r ), .c(\U1297/naack ) );
    nand2_2 \U1297/U1128/U28/U1/U3  ( .x(csel), .a(\U1297/U1128/U28/U1/clr ), 
        .b(\U1297/U1128/U28/U1/set ) );
    aoai211_1 \U1297/U1127/U28/U1/U1  ( .x(\U1297/U1127/U28/U1/clr ), .a(
        \U1297/s ), .b(\U1297/nback ), .c(ag), .d(asel) );
    nand3_1 \U1297/U1127/U28/U1/U2  ( .x(\U1297/U1127/U28/U1/set ), .a(ag), 
        .b(\U1297/s ), .c(\U1297/nback ) );
    nand2_2 \U1297/U1127/U28/U1/U3  ( .x(asel), .a(\U1297/U1127/U28/U1/clr ), 
        .b(\U1297/U1127/U28/U1/set ) );
    nand2_1 \U1300/U1131/U5  ( .x(\U1300/s ), .a(\U1300/r ), .b(\U1300/nback )
         );
    nand2_1 \U1300/U1103/U5  ( .x(\U1300/r ), .a(\U1300/naack ), .b(\U1300/s )
         );
    inv_1 \U1300/U1111/U3  ( .x(\U1300/reset ), .a(nbReset) );
    inv_1 \U1300/U1112/U3  ( .x(\U1300/naack ), .a(nba) );
    nor2_1 \U1300/U1130/U5  ( .x(\U1300/nback ), .a(nda), .b(\U1300/reset ) );
    aoai211_1 \U1300/U1128/U28/U1/U1  ( .x(\U1300/U1128/U28/U1/clr ), .a(
        \U1300/r ), .b(\U1300/naack ), .c(dg), .d(dsel) );
    nand3_1 \U1300/U1128/U28/U1/U2  ( .x(\U1300/U1128/U28/U1/set ), .a(dg), 
        .b(\U1300/r ), .c(\U1300/naack ) );
    nand2_2 \U1300/U1128/U28/U1/U3  ( .x(dsel), .a(\U1300/U1128/U28/U1/clr ), 
        .b(\U1300/U1128/U28/U1/set ) );
    aoai211_1 \U1300/U1127/U28/U1/U1  ( .x(\U1300/U1127/U28/U1/clr ), .a(
        \U1300/s ), .b(\U1300/nback ), .c(bg), .d(bsel) );
    nand3_1 \U1300/U1127/U28/U1/U2  ( .x(\U1300/U1127/U28/U1/set ), .a(bg), 
        .b(\U1300/s ), .c(\U1300/nback ) );
    nand2_2 \U1300/U1127/U28/U1/U3  ( .x(bsel), .a(\U1300/U1127/U28/U1/clr ), 
        .b(\U1300/U1127/U28/U1/set ) );
    aoai211_1 \U1289/U1150/U28/U1/U1  ( .x(\U1289/U1150/U28/U1/clr ), .a(il[2]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdl[2] ) );
    nand3_1 \U1289/U1150/U28/U1/U2  ( .x(\U1289/U1150/U28/U1/set ), .a(net195), 
        .b(il[2]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1150/U28/U1/U3  ( .x(\cdl[2] ), .a(
        \U1289/U1150/U28/U1/clr ), .b(\U1289/U1150/U28/U1/set ) );
    aoai211_1 \U1289/U1152/U28/U1/U1  ( .x(\U1289/U1152/U28/U1/clr ), .a(il[3]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdl[3] ) );
    nand3_1 \U1289/U1152/U28/U1/U2  ( .x(\U1289/U1152/U28/U1/set ), .a(net195), 
        .b(il[3]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1152/U28/U1/U3  ( .x(\cdl[3] ), .a(
        \U1289/U1152/U28/U1/clr ), .b(\U1289/U1152/U28/U1/set ) );
    aoai211_1 \U1289/U1149/U28/U1/U1  ( .x(\U1289/U1149/U28/U1/clr ), .a(ih[2]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdh[2] ) );
    nand3_1 \U1289/U1149/U28/U1/U2  ( .x(\U1289/U1149/U28/U1/set ), .a(net195), 
        .b(ih[2]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1149/U28/U1/U3  ( .x(\cdh[2] ), .a(
        \U1289/U1149/U28/U1/clr ), .b(\U1289/U1149/U28/U1/set ) );
    aoai211_1 \U1289/U1151/U28/U1/U1  ( .x(\U1289/U1151/U28/U1/clr ), .a(ih[3]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdh[3] ) );
    nand3_1 \U1289/U1151/U28/U1/U2  ( .x(\U1289/U1151/U28/U1/set ), .a(net195), 
        .b(ih[3]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1151/U28/U1/U3  ( .x(\cdh[3] ), .a(
        \U1289/U1151/U28/U1/clr ), .b(\U1289/U1151/U28/U1/set ) );
    inv_1 \U1289/U1148/U1147/U3  ( .x(\U1289/U1148/net189 ), .a(
        \U1289/bnreset ) );
    nor2_1 \U1289/U1148/U582/U5  ( .x(\U1289/U1148/net192 ), .a(\cdl[3] ), .b(
        \cdh[3] ) );
    nor2_1 \U1289/U1148/U580/U5  ( .x(\U1289/U1148/net191 ), .a(\cdl[2] ), .b(
        \cdh[2] ) );
    nor2_2 \U1289/U1148/U1146/U6  ( .x(\twobitack[2] ), .a(
        \U1289/U1148/net190 ), .b(\U1289/U1148/net189 ) );
    aoi222_1 \U1289/U1148/U1141/U30/U1  ( .x(\U1289/U1148/net190 ), .a(
        \U1289/U1148/net191 ), .b(\U1289/U1148/net192 ), .c(
        \U1289/U1148/net191 ), .d(\U1289/U1148/U1141/Z ), .e(
        \U1289/U1148/net192 ), .f(\U1289/U1148/U1141/Z ) );
    inv_1 \U1289/U1148/U1141/U30/Uinv  ( .x(\U1289/U1148/U1141/Z ), .a(
        \U1289/U1148/net190 ) );
    aoai211_1 \U1271/U1150/U28/U1/U1  ( .x(\U1271/U1150/U28/U1/clr ), .a(il[0]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdl[0] ) );
    nand3_1 \U1271/U1150/U28/U1/U2  ( .x(\U1271/U1150/U28/U1/set ), .a(net193), 
        .b(il[0]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1150/U28/U1/U3  ( .x(\cdl[0] ), .a(
        \U1271/U1150/U28/U1/clr ), .b(\U1271/U1150/U28/U1/set ) );
    aoai211_1 \U1271/U1152/U28/U1/U1  ( .x(\U1271/U1152/U28/U1/clr ), .a(il[1]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdl[1] ) );
    nand3_1 \U1271/U1152/U28/U1/U2  ( .x(\U1271/U1152/U28/U1/set ), .a(net193), 
        .b(il[1]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1152/U28/U1/U3  ( .x(\cdl[1] ), .a(
        \U1271/U1152/U28/U1/clr ), .b(\U1271/U1152/U28/U1/set ) );
    aoai211_1 \U1271/U1149/U28/U1/U1  ( .x(\U1271/U1149/U28/U1/clr ), .a(ih[0]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdh[0] ) );
    nand3_1 \U1271/U1149/U28/U1/U2  ( .x(\U1271/U1149/U28/U1/set ), .a(net193), 
        .b(ih[0]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1149/U28/U1/U3  ( .x(\cdh[0] ), .a(
        \U1271/U1149/U28/U1/clr ), .b(\U1271/U1149/U28/U1/set ) );
    aoai211_1 \U1271/U1151/U28/U1/U1  ( .x(\U1271/U1151/U28/U1/clr ), .a(ih[1]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdh[1] ) );
    nand3_1 \U1271/U1151/U28/U1/U2  ( .x(\U1271/U1151/U28/U1/set ), .a(net193), 
        .b(ih[1]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1151/U28/U1/U3  ( .x(\cdh[1] ), .a(
        \U1271/U1151/U28/U1/clr ), .b(\U1271/U1151/U28/U1/set ) );
    inv_1 \U1271/U1148/U1147/U3  ( .x(\U1271/U1148/net189 ), .a(
        \U1271/bnreset ) );
    nor2_1 \U1271/U1148/U582/U5  ( .x(\U1271/U1148/net192 ), .a(\cdl[1] ), .b(
        \cdh[1] ) );
    nor2_1 \U1271/U1148/U580/U5  ( .x(\U1271/U1148/net191 ), .a(\cdl[0] ), .b(
        \cdh[0] ) );
    nor2_2 \U1271/U1148/U1146/U6  ( .x(\twobitack[0] ), .a(
        \U1271/U1148/net190 ), .b(\U1271/U1148/net189 ) );
    aoi222_1 \U1271/U1148/U1141/U30/U1  ( .x(\U1271/U1148/net190 ), .a(
        \U1271/U1148/net191 ), .b(\U1271/U1148/net192 ), .c(
        \U1271/U1148/net191 ), .d(\U1271/U1148/U1141/Z ), .e(
        \U1271/U1148/net192 ), .f(\U1271/U1148/U1141/Z ) );
    inv_1 \U1271/U1148/U1141/U30/Uinv  ( .x(\U1271/U1148/U1141/Z ), .a(
        \U1271/U1148/net190 ) );
    nand2_1 \U1225/U1128/U5  ( .x(\U1225/s ), .a(\U1225/r ), .b(\U1225/nback )
         );
    nand2_1 \U1225/U1103/U5  ( .x(\U1225/r ), .a(\U1225/naack ), .b(\U1225/s )
         );
    inv_1 \U1225/U1111/U3  ( .x(\U1225/reset ), .a(nbReset) );
    inv_1 \U1225/U1112/U3  ( .x(\U1225/naack ), .a(nxa) );
    nor2_1 \U1225/U1127/U5  ( .x(\U1225/nback ), .a(nyla), .b(\U1225/reset )
         );
    and2_2 \U1225/U1129/U8  ( .x(xsel), .a(\U1225/nback ), .b(\U1225/s ) );
    and2_2 \U1225/U1124/U8  ( .x(ysel), .a(\U1225/r ), .b(\U1225/naack ) );
    and3_4 \U1308/U20/U9  ( .x(nya), .a(\U1308/nack[1] ), .b(\U1308/nack[0] ), 
        .c(nbReset) );
    nor2_1 \U1308/U18/U5  ( .x(\U1308/nack[0] ), .a(\yl[3] ), .b(\yl[0] ) );
    nor2_1 \U1308/U19/U5  ( .x(\U1308/nack[1] ), .a(\yl[1] ), .b(\yl[2] ) );
    ao222_2 \U1308/U15_0_/U19/U1/U1  ( .x(\yl[0] ), .a(\y[0] ), .b(nyla), .c(
        \y[0] ), .d(\yl[0] ), .e(nyla), .f(\yl[0] ) );
    ao222_2 \U1308/U15_1_/U19/U1/U1  ( .x(\yl[1] ), .a(\y[1] ), .b(nyla), .c(
        \y[1] ), .d(\yl[1] ), .e(nyla), .f(\yl[1] ) );
    ao222_2 \U1308/U15_2_/U19/U1/U1  ( .x(\yl[2] ), .a(\y[2] ), .b(nyla), .c(
        \y[2] ), .d(\yl[2] ), .e(nyla), .f(\yl[2] ) );
    ao222_2 \U1308/U15_3_/U19/U1/U1  ( .x(\yl[3] ), .a(\y[3] ), .b(nyla), .c(
        \y[3] ), .d(\yl[3] ), .e(nyla), .f(\yl[3] ) );
    buf_3 U1 ( .x(\U1271/bnreset ), .a(nbReset) );
    buf_3 U2 ( .x(\U1289/bnreset ), .a(nbReset) );
endmodule


module chain_mergepackets_3 ( naa, nba, o, a, b, nReset, noa );
output [4:0] o;
input  [4:0] a;
input  [4:0] b;
input  nReset, noa;
output naa, nba;
    wire as, seta, asel, bsel, setb, reset, \noack[1] , \noack[0] , 
        \U916_0_/U25/U1/clr , \U916_0_/U25/U1/ob , \U916_1_/U25/U1/clr , 
        \U916_1_/U25/U1/ob , \U916_2_/U25/U1/clr , \U916_2_/U25/U1/ob , 
        \U916_3_/U25/U1/clr , \U916_3_/U25/U1/ob ;
    and2_1 \U1155/U8  ( .x(as), .a(seta), .b(asel) );
    nand2_1 \U1145/U5  ( .x(asel), .a(bsel), .b(seta) );
    nand2_1 \U1103/U5  ( .x(bsel), .a(setb), .b(asel) );
    inv_1 \U1135/U3  ( .x(reset), .a(nReset) );
    inv_1 \U1134/U3  ( .x(setb), .a(a[4]) );
    and3_2 \U1154/U9  ( .x(naa), .a(\noack[1] ), .b(\noack[0] ), .c(as) );
    nor3_1 \U1127/U7  ( .x(\noack[0] ), .a(o[1]), .b(reset), .c(o[0]) );
    nor2_1 \U1132/U5  ( .x(\noack[1] ), .a(o[3]), .b(o[2]) );
    oa31_1 \U916_0_/U25/U1/Uclr  ( .x(\U916_0_/U25/U1/clr ), .a(noa), .b(a[0]), 
        .c(b[0]), .d(o[0]) );
    oaoi211_1 \U916_0_/U25/U1/Uaoi  ( .x(\U916_0_/U25/U1/ob ), .a(a[0]), .b(b
        [0]), .c(noa), .d(\U916_0_/U25/U1/clr ) );
    inv_2 \U916_0_/U25/U1/Ui  ( .x(o[0]), .a(\U916_0_/U25/U1/ob ) );
    oa31_1 \U916_1_/U25/U1/Uclr  ( .x(\U916_1_/U25/U1/clr ), .a(noa), .b(a[1]), 
        .c(b[1]), .d(o[1]) );
    oaoi211_1 \U916_1_/U25/U1/Uaoi  ( .x(\U916_1_/U25/U1/ob ), .a(a[1]), .b(b
        [1]), .c(noa), .d(\U916_1_/U25/U1/clr ) );
    inv_2 \U916_1_/U25/U1/Ui  ( .x(o[1]), .a(\U916_1_/U25/U1/ob ) );
    oa31_1 \U916_2_/U25/U1/Uclr  ( .x(\U916_2_/U25/U1/clr ), .a(noa), .b(a[2]), 
        .c(b[2]), .d(o[2]) );
    oaoi211_1 \U916_2_/U25/U1/Uaoi  ( .x(\U916_2_/U25/U1/ob ), .a(a[2]), .b(b
        [2]), .c(noa), .d(\U916_2_/U25/U1/clr ) );
    inv_2 \U916_2_/U25/U1/Ui  ( .x(o[2]), .a(\U916_2_/U25/U1/ob ) );
    oa31_1 \U916_3_/U25/U1/Uclr  ( .x(\U916_3_/U25/U1/clr ), .a(noa), .b(a[3]), 
        .c(b[3]), .d(o[3]) );
    oaoi211_1 \U916_3_/U25/U1/Uaoi  ( .x(\U916_3_/U25/U1/ob ), .a(a[3]), .b(b
        [3]), .c(noa), .d(\U916_3_/U25/U1/clr ) );
    inv_2 \U916_3_/U25/U1/Ui  ( .x(o[3]), .a(\U916_3_/U25/U1/ob ) );
    ao222_2 \U1148/U19/U1/U1  ( .x(o[4]), .a(noa), .b(b[4]), .c(noa), .d(o[4]), 
        .e(b[4]), .f(o[4]) );
    aoi21_1 \U1153/U11  ( .x(seta), .a(o[4]), .b(setb), .c(reset) );
    and3_3 U1 ( .x(nba), .a(bsel), .b(\noack[0] ), .c(\noack[1] ) );
endmodule


module chain_tchdr_0 ( addr_req, col_h, col_l, itag_h, itag_l, lock, ncback, 
    neop, pred, pullcd, reset, rnw_h, rnw_l, seq, size_h, size_l, write_req, 
    chwh, chwl, addr_ack, addr_pull, nReset, nack, write_ack, write_pull );
output [2:0] col_h;
output [2:0] col_l;
output [4:0] itag_h;
output [4:0] itag_l;
output [1:0] lock;
output [1:0] pred;
output [1:0] seq;
output [1:0] size_h;
output [1:0] size_l;
input  [7:0] chwh;
input  [7:0] chwl;
input  addr_ack, addr_pull, nReset, nack, write_ack, write_pull;
output addr_req, ncback, neop, pullcd, reset, rnw_h, rnw_l, write_req;
    wire n9, pullcdwk, net94, net88, \ncd[0] , \ncd[1] , \ncd[2] , \ncd[3] , 
        \ncd[4] , \ncd[5] , \ncd[6] , \ncd[7] , read, ack, net83, \U1664/x[3] , 
        \U1664/U28/Z , \U1664/x[0] , \U1664/U32/Z , \U1664/x[2] , 
        \U1664/U29/Z , \U1664/y[0] , \U1664/x[1] , \U1664/U33/Z , \U1664/y[1] , 
        \U1664/U30/Z , \U1664/U31/Z , \U1664/U37/Z , receive, \U473/Z , 
        \hdr_hld/net32 , \hdr_hld/net33 , \hdr_hld/low/latch , 
        \hdr_hld/low/nlocalcd , \hdr_hld/low/localcd , \hdr_hld/low/ncd[0] , 
        \hdr_hld/low/ncd[1] , \hdr_hld/low/ncd[2] , \hdr_hld/low/ncd[3] , 
        \hdr_hld/ol[3] , \hdr_hld/oh[3] , \hdr_hld/low/ncd[4] , 
        \hdr_hld/ol[4] , \hdr_hld/oh[4] , \hdr_hld/low/ncd[5] , 
        \hdr_hld/low/ncd[6] , \hdr_hld/low/ncd[7] , 
        \hdr_hld/low/ctrlack_internal , \hdr_hld/low/acb , \hdr_hld/low/ba , 
        \hdr_hld/low/driveh , \hdr_hld/net20 , \hdr_hld/low/drivel , n7, n5, 
        n6, \hdr_hld/low/U4/U28/U1/clr , \hdr_hld/low/U4/U28/U1/set , 
        \hdr_hld/low/U1/Z , \hdr_hld/low/U1664/x[3] , 
        \hdr_hld/low/U1664/U28/Z , \hdr_hld/low/U1664/x[0] , 
        \hdr_hld/low/U1664/U32/Z , \hdr_hld/low/U1664/x[2] , 
        \hdr_hld/low/U1664/U29/Z , \hdr_hld/low/U1664/y[0] , 
        \hdr_hld/low/U1664/x[1] , \hdr_hld/low/U1664/U33/Z , 
        \hdr_hld/low/U1664/y[1] , \hdr_hld/low/U1664/U30/Z , 
        \hdr_hld/low/U1664/U31/Z , \hdr_hld/low/U1664/U37/Z , 
        \hdr_hld/low/U1669/nr , \hdr_hld/low/U1669/nd , \hdr_hld/low/U1669/n2 , 
        \hdr_hld/high/latch , \hdr_hld/high/nlocalcd , \hdr_hld/high/localcd , 
        \hdr_hld/high/ncd[0] , \hdr_hld/high/ncd[1] , \hdr_hld/high/ncd[2] , 
        \hdr_hld/high/ncd[3] , \hdr_hld/high/ncd[4] , \hdr_hld/high/ncd[5] , 
        \hdr_hld/high/ncd[6] , \hdr_hld/high/ncd[7] , 
        \hdr_hld/high/ctrlack_internal , \hdr_hld/high/acb , \hdr_hld/high/ba , 
        \hdr_hld/high/driveh , \hdr_hld/high/drivel , n1, n4, n2, n3, 
        \hdr_hld/high/U4/U28/U1/clr , \hdr_hld/high/U4/U28/U1/set , 
        \hdr_hld/high/U1/Z , \hdr_hld/high/U1664/x[3] , 
        \hdr_hld/high/U1664/U28/Z , \hdr_hld/high/U1664/x[0] , 
        \hdr_hld/high/U1664/U32/Z , \hdr_hld/high/U1664/x[2] , 
        \hdr_hld/high/U1664/U29/Z , \hdr_hld/high/U1664/y[0] , 
        \hdr_hld/high/U1664/x[1] , \hdr_hld/high/U1664/U33/Z , 
        \hdr_hld/high/U1664/y[1] , \hdr_hld/high/U1664/U30/Z , 
        \hdr_hld/high/U1664/U31/Z , \hdr_hld/high/U1664/U37/Z , 
        \hdr_hld/high/U1669/nr , \hdr_hld/high/U1669/nd , 
        \hdr_hld/high/U1669/n2 ;
    buf_1 U262 ( .x(n9), .a(pullcdwk) );
    or3_2 \U1668/U12  ( .x(ncback), .a(net94), .b(addr_pull), .c(write_pull)
         );
    inv_1 \I0/U3  ( .x(net94), .a(net88) );
    nor2_1 \U514_0_/U5  ( .x(\ncd[0] ), .a(chwh[0]), .b(chwl[0]) );
    nor2_1 \U514_1_/U5  ( .x(\ncd[1] ), .a(chwh[1]), .b(chwl[1]) );
    nor2_1 \U514_2_/U5  ( .x(\ncd[2] ), .a(chwh[2]), .b(chwl[2]) );
    nor2_1 \U514_3_/U5  ( .x(\ncd[3] ), .a(chwh[3]), .b(chwl[3]) );
    nor2_1 \U514_4_/U5  ( .x(\ncd[4] ), .a(chwh[4]), .b(chwl[4]) );
    nor2_1 \U514_5_/U5  ( .x(\ncd[5] ), .a(chwh[5]), .b(chwl[5]) );
    nor2_1 \U514_6_/U5  ( .x(\ncd[6] ), .a(chwh[6]), .b(chwl[6]) );
    nor2_1 \U514_7_/U5  ( .x(\ncd[7] ), .a(chwh[7]), .b(chwl[7]) );
    nor2_1 \U1669/U5  ( .x(neop), .a(read), .b(write_ack) );
    nand2_1 \U303/U5  ( .x(ack), .a(nack), .b(nReset) );
    nand2_1 \U1670/U5  ( .x(net83), .a(neop), .b(nReset) );
    ao222_1 \U47/U18/U1/U1  ( .x(read), .a(addr_ack), .b(rnw_h), .c(addr_ack), 
        .d(read), .e(rnw_h), .f(read) );
    ao222_1 \U48/U18/U1/U1  ( .x(write_req), .a(rnw_l), .b(addr_ack), .c(rnw_l
        ), .d(write_req), .e(addr_ack), .f(write_req) );
    aoi222_1 \U1664/U28/U30/U1  ( .x(\U1664/x[3] ), .a(\ncd[7] ), .b(\ncd[6] ), 
        .c(\ncd[7] ), .d(\U1664/U28/Z ), .e(\ncd[6] ), .f(\U1664/U28/Z ) );
    inv_1 \U1664/U28/U30/Uinv  ( .x(\U1664/U28/Z ), .a(\U1664/x[3] ) );
    aoi222_1 \U1664/U32/U30/U1  ( .x(\U1664/x[0] ), .a(\ncd[1] ), .b(\ncd[0] ), 
        .c(\ncd[1] ), .d(\U1664/U32/Z ), .e(\ncd[0] ), .f(\U1664/U32/Z ) );
    inv_1 \U1664/U32/U30/Uinv  ( .x(\U1664/U32/Z ), .a(\U1664/x[0] ) );
    aoi222_1 \U1664/U29/U30/U1  ( .x(\U1664/x[2] ), .a(\ncd[5] ), .b(\ncd[4] ), 
        .c(\ncd[5] ), .d(\U1664/U29/Z ), .e(\ncd[4] ), .f(\U1664/U29/Z ) );
    inv_1 \U1664/U29/U30/Uinv  ( .x(\U1664/U29/Z ), .a(\U1664/x[2] ) );
    aoi222_1 \U1664/U33/U30/U1  ( .x(\U1664/y[0] ), .a(\U1664/x[1] ), .b(
        \U1664/x[0] ), .c(\U1664/x[1] ), .d(\U1664/U33/Z ), .e(\U1664/x[0] ), 
        .f(\U1664/U33/Z ) );
    inv_1 \U1664/U33/U30/Uinv  ( .x(\U1664/U33/Z ), .a(\U1664/y[0] ) );
    aoi222_1 \U1664/U30/U30/U1  ( .x(\U1664/y[1] ), .a(\U1664/x[3] ), .b(
        \U1664/x[2] ), .c(\U1664/x[3] ), .d(\U1664/U30/Z ), .e(\U1664/x[2] ), 
        .f(\U1664/U30/Z ) );
    inv_1 \U1664/U30/U30/Uinv  ( .x(\U1664/U30/Z ), .a(\U1664/y[1] ) );
    aoi222_1 \U1664/U31/U30/U1  ( .x(\U1664/x[1] ), .a(\ncd[3] ), .b(\ncd[2] ), 
        .c(\ncd[3] ), .d(\U1664/U31/Z ), .e(\ncd[2] ), .f(\U1664/U31/Z ) );
    inv_1 \U1664/U31/U30/Uinv  ( .x(\U1664/U31/Z ), .a(\U1664/x[1] ) );
    aoi222_1 \U1664/U37/U30/U1  ( .x(pullcdwk), .a(\U1664/y[0] ), .b(
        \U1664/y[1] ), .c(\U1664/y[0] ), .d(\U1664/U37/Z ), .e(\U1664/y[1] ), 
        .f(\U1664/U37/Z ) );
    inv_1 \U1664/U37/U30/Uinv  ( .x(\U1664/U37/Z ), .a(pullcdwk) );
    aoi222_1 \U473/U30/U1  ( .x(receive), .a(net83), .b(ack), .c(net83), .d(
        \U473/Z ), .e(ack), .f(\U473/Z ) );
    inv_1 \U473/U30/Uinv  ( .x(\U473/Z ), .a(receive) );
    nor2_1 \hdr_hld/U3/U5  ( .x(net88), .a(\hdr_hld/net32 ), .b(
        \hdr_hld/net33 ) );
    buf_2 \hdr_hld/low/U1653  ( .x(\hdr_hld/low/latch ), .a(\hdr_hld/net32 )
         );
    nor2_1 \hdr_hld/low/U264/U5  ( .x(\hdr_hld/low/nlocalcd ), .a(reset), .b(
        \hdr_hld/low/localcd ) );
    nor2_1 \hdr_hld/low/U1659_0_/U5  ( .x(\hdr_hld/low/ncd[0] ), .a(seq[0]), 
        .b(seq[1]) );
    nor2_1 \hdr_hld/low/U1659_1_/U5  ( .x(\hdr_hld/low/ncd[1] ), .a(pred[0]), 
        .b(pred[1]) );
    nor2_1 \hdr_hld/low/U1659_2_/U5  ( .x(\hdr_hld/low/ncd[2] ), .a(lock[0]), 
        .b(lock[1]) );
    nor2_1 \hdr_hld/low/U1659_3_/U5  ( .x(\hdr_hld/low/ncd[3] ), .a(
        \hdr_hld/ol[3] ), .b(\hdr_hld/oh[3] ) );
    nor2_1 \hdr_hld/low/U1659_4_/U5  ( .x(\hdr_hld/low/ncd[4] ), .a(
        \hdr_hld/ol[4] ), .b(\hdr_hld/oh[4] ) );
    nor2_1 \hdr_hld/low/U1659_5_/U5  ( .x(\hdr_hld/low/ncd[5] ), .a(rnw_l), 
        .b(rnw_h) );
    nor2_1 \hdr_hld/low/U1659_6_/U5  ( .x(\hdr_hld/low/ncd[6] ), .a(size_l[0]), 
        .b(size_h[0]) );
    nor2_1 \hdr_hld/low/U1659_7_/U5  ( .x(\hdr_hld/low/ncd[7] ), .a(size_l[1]), 
        .b(size_h[1]) );
    nor2_1 \hdr_hld/low/U3/U5  ( .x(\hdr_hld/low/ctrlack_internal ), .a(
        \hdr_hld/low/acb ), .b(\hdr_hld/low/ba ) );
    buf_2 \hdr_hld/low/U1665/U7  ( .x(\hdr_hld/low/driveh ), .a(
        \hdr_hld/net20 ) );
    buf_2 \hdr_hld/low/U1666/U7  ( .x(\hdr_hld/low/drivel ), .a(
        \hdr_hld/net20 ) );
    ao23_1 \hdr_hld/low/U1658_0_/U21/U1/U1  ( .x(seq[0]), .a(n7), .b(seq[0]), 
        .c(n7), .d(chwl[0]), .e(n5) );
    ao23_1 \hdr_hld/low/U1658_1_/U21/U1/U1  ( .x(pred[0]), .a(
        \hdr_hld/low/drivel ), .b(pred[0]), .c(\hdr_hld/low/drivel ), .d(chwl
        [1]), .e(n5) );
    ao23_1 \hdr_hld/low/U1658_2_/U21/U1/U1  ( .x(lock[0]), .a(n6), .b(lock[0]), 
        .c(n7), .d(chwl[2]), .e(n5) );
    ao23_1 \hdr_hld/low/U1658_3_/U21/U1/U1  ( .x(\hdr_hld/ol[3] ), .a(
        \hdr_hld/low/drivel ), .b(\hdr_hld/ol[3] ), .c(n6), .d(chwl[3]), .e(
        \hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1658_4_/U21/U1/U1  ( .x(\hdr_hld/ol[4] ), .a(n7), .b(
        \hdr_hld/ol[4] ), .c(n6), .d(chwl[4]), .e(\hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1658_5_/U21/U1/U1  ( .x(rnw_l), .a(n7), .b(rnw_l), 
        .c(n7), .d(chwl[5]), .e(\hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1658_6_/U21/U1/U1  ( .x(size_l[0]), .a(
        \hdr_hld/low/driveh ), .b(size_l[0]), .c(n6), .d(chwl[6]), .e(
        \hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1658_7_/U21/U1/U1  ( .x(size_l[1]), .a(
        \hdr_hld/low/driveh ), .b(size_l[1]), .c(n7), .d(chwl[7]), .e(
        \hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1651_0_/U21/U1/U1  ( .x(seq[1]), .a(
        \hdr_hld/low/driveh ), .b(seq[1]), .c(n6), .d(chwh[0]), .e(
        \hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1651_1_/U21/U1/U1  ( .x(pred[1]), .a(
        \hdr_hld/low/drivel ), .b(pred[1]), .c(\hdr_hld/low/drivel ), .d(chwh
        [1]), .e(\hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1651_2_/U21/U1/U1  ( .x(lock[1]), .a(n6), .b(lock[1]), 
        .c(\hdr_hld/low/driveh ), .d(chwh[2]), .e(\hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1651_3_/U21/U1/U1  ( .x(\hdr_hld/oh[3] ), .a(
        \hdr_hld/low/drivel ), .b(\hdr_hld/oh[3] ), .c(\hdr_hld/low/driveh ), 
        .d(chwh[3]), .e(\hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1651_4_/U21/U1/U1  ( .x(\hdr_hld/oh[4] ), .a(n7), .b(
        \hdr_hld/oh[4] ), .c(\hdr_hld/low/drivel ), .d(chwh[4]), .e(
        \hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1651_5_/U21/U1/U1  ( .x(rnw_h), .a(
        \hdr_hld/low/driveh ), .b(rnw_h), .c(\hdr_hld/low/driveh ), .d(chwh[5]
        ), .e(\hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1651_6_/U21/U1/U1  ( .x(size_h[0]), .a(n6), .b(size_h
        [0]), .c(\hdr_hld/low/drivel ), .d(chwh[6]), .e(\hdr_hld/low/latch )
         );
    ao23_1 \hdr_hld/low/U1651_7_/U21/U1/U1  ( .x(size_h[1]), .a(n6), .b(size_h
        [1]), .c(\hdr_hld/low/driveh ), .d(chwh[7]), .e(\hdr_hld/low/latch )
         );
    aoai211_1 \hdr_hld/low/U4/U28/U1/U1  ( .x(\hdr_hld/low/U4/U28/U1/clr ), 
        .a(\hdr_hld/net20 ), .b(\hdr_hld/low/acb ), .c(\hdr_hld/low/nlocalcd ), 
        .d(\hdr_hld/net32 ) );
    nand3_1 \hdr_hld/low/U4/U28/U1/U2  ( .x(\hdr_hld/low/U4/U28/U1/set ), .a(
        \hdr_hld/low/nlocalcd ), .b(\hdr_hld/net20 ), .c(\hdr_hld/low/acb ) );
    nand2_2 \hdr_hld/low/U4/U28/U1/U3  ( .x(\hdr_hld/net32 ), .a(
        \hdr_hld/low/U4/U28/U1/clr ), .b(\hdr_hld/low/U4/U28/U1/set ) );
    oai21_1 \hdr_hld/low/U1/U30/U1/U1  ( .x(\hdr_hld/low/acb ), .a(
        \hdr_hld/low/U1/Z ), .b(\hdr_hld/low/ba ), .c(\hdr_hld/net20 ) );
    inv_1 \hdr_hld/low/U1/U30/U1/U2  ( .x(\hdr_hld/low/U1/Z ), .a(
        \hdr_hld/low/acb ) );
    ao222_1 \hdr_hld/low/U5/U18/U1/U1  ( .x(\hdr_hld/low/ba ), .a(
        \hdr_hld/low/latch ), .b(n9), .c(\hdr_hld/low/latch ), .d(
        \hdr_hld/low/ba ), .e(n9), .f(\hdr_hld/low/ba ) );
    aoi222_1 \hdr_hld/low/U1664/U28/U30/U1  ( .x(\hdr_hld/low/U1664/x[3] ), 
        .a(\hdr_hld/low/ncd[7] ), .b(\hdr_hld/low/ncd[6] ), .c(
        \hdr_hld/low/ncd[7] ), .d(\hdr_hld/low/U1664/U28/Z ), .e(
        \hdr_hld/low/ncd[6] ), .f(\hdr_hld/low/U1664/U28/Z ) );
    inv_1 \hdr_hld/low/U1664/U28/U30/Uinv  ( .x(\hdr_hld/low/U1664/U28/Z ), 
        .a(\hdr_hld/low/U1664/x[3] ) );
    aoi222_1 \hdr_hld/low/U1664/U32/U30/U1  ( .x(\hdr_hld/low/U1664/x[0] ), 
        .a(\hdr_hld/low/ncd[1] ), .b(\hdr_hld/low/ncd[0] ), .c(
        \hdr_hld/low/ncd[1] ), .d(\hdr_hld/low/U1664/U32/Z ), .e(
        \hdr_hld/low/ncd[0] ), .f(\hdr_hld/low/U1664/U32/Z ) );
    inv_1 \hdr_hld/low/U1664/U32/U30/Uinv  ( .x(\hdr_hld/low/U1664/U32/Z ), 
        .a(\hdr_hld/low/U1664/x[0] ) );
    aoi222_1 \hdr_hld/low/U1664/U29/U30/U1  ( .x(\hdr_hld/low/U1664/x[2] ), 
        .a(\hdr_hld/low/ncd[5] ), .b(\hdr_hld/low/ncd[4] ), .c(
        \hdr_hld/low/ncd[5] ), .d(\hdr_hld/low/U1664/U29/Z ), .e(
        \hdr_hld/low/ncd[4] ), .f(\hdr_hld/low/U1664/U29/Z ) );
    inv_1 \hdr_hld/low/U1664/U29/U30/Uinv  ( .x(\hdr_hld/low/U1664/U29/Z ), 
        .a(\hdr_hld/low/U1664/x[2] ) );
    aoi222_1 \hdr_hld/low/U1664/U33/U30/U1  ( .x(\hdr_hld/low/U1664/y[0] ), 
        .a(\hdr_hld/low/U1664/x[1] ), .b(\hdr_hld/low/U1664/x[0] ), .c(
        \hdr_hld/low/U1664/x[1] ), .d(\hdr_hld/low/U1664/U33/Z ), .e(
        \hdr_hld/low/U1664/x[0] ), .f(\hdr_hld/low/U1664/U33/Z ) );
    inv_1 \hdr_hld/low/U1664/U33/U30/Uinv  ( .x(\hdr_hld/low/U1664/U33/Z ), 
        .a(\hdr_hld/low/U1664/y[0] ) );
    aoi222_1 \hdr_hld/low/U1664/U30/U30/U1  ( .x(\hdr_hld/low/U1664/y[1] ), 
        .a(\hdr_hld/low/U1664/x[3] ), .b(\hdr_hld/low/U1664/x[2] ), .c(
        \hdr_hld/low/U1664/x[3] ), .d(\hdr_hld/low/U1664/U30/Z ), .e(
        \hdr_hld/low/U1664/x[2] ), .f(\hdr_hld/low/U1664/U30/Z ) );
    inv_1 \hdr_hld/low/U1664/U30/U30/Uinv  ( .x(\hdr_hld/low/U1664/U30/Z ), 
        .a(\hdr_hld/low/U1664/y[1] ) );
    aoi222_1 \hdr_hld/low/U1664/U31/U30/U1  ( .x(\hdr_hld/low/U1664/x[1] ), 
        .a(\hdr_hld/low/ncd[3] ), .b(\hdr_hld/low/ncd[2] ), .c(
        \hdr_hld/low/ncd[3] ), .d(\hdr_hld/low/U1664/U31/Z ), .e(
        \hdr_hld/low/ncd[2] ), .f(\hdr_hld/low/U1664/U31/Z ) );
    inv_1 \hdr_hld/low/U1664/U31/U30/Uinv  ( .x(\hdr_hld/low/U1664/U31/Z ), 
        .a(\hdr_hld/low/U1664/x[1] ) );
    aoi222_1 \hdr_hld/low/U1664/U37/U30/U1  ( .x(\hdr_hld/low/localcd ), .a(
        \hdr_hld/low/U1664/y[0] ), .b(\hdr_hld/low/U1664/y[1] ), .c(
        \hdr_hld/low/U1664/y[0] ), .d(\hdr_hld/low/U1664/U37/Z ), .e(
        \hdr_hld/low/U1664/y[1] ), .f(\hdr_hld/low/U1664/U37/Z ) );
    inv_1 \hdr_hld/low/U1664/U37/U30/Uinv  ( .x(\hdr_hld/low/U1664/U37/Z ), 
        .a(\hdr_hld/low/localcd ) );
    nor3_1 \hdr_hld/low/U1669/Unr  ( .x(\hdr_hld/low/U1669/nr ), .a(
        \hdr_hld/low/ctrlack_internal ), .b(\hdr_hld/low/drivel ), .c(n6) );
    nand3_1 \hdr_hld/low/U1669/Und  ( .x(\hdr_hld/low/U1669/nd ), .a(
        \hdr_hld/low/ctrlack_internal ), .b(n7), .c(\hdr_hld/low/driveh ) );
    oa21_1 \hdr_hld/low/U1669/U1  ( .x(\hdr_hld/low/U1669/n2 ), .a(
        \hdr_hld/low/U1669/n2 ), .b(\hdr_hld/low/U1669/nr ), .c(
        \hdr_hld/low/U1669/nd ) );
    inv_2 \hdr_hld/low/U1669/U3  ( .x(addr_req), .a(\hdr_hld/low/U1669/n2 ) );
    buf_2 \hdr_hld/high/U1653  ( .x(\hdr_hld/high/latch ), .a(\hdr_hld/net33 )
         );
    nor2_1 \hdr_hld/high/U264/U5  ( .x(\hdr_hld/high/nlocalcd ), .a(reset), 
        .b(\hdr_hld/high/localcd ) );
    nor2_1 \hdr_hld/high/U1659_0_/U5  ( .x(\hdr_hld/high/ncd[0] ), .a(itag_l
        [0]), .b(itag_h[0]) );
    nor2_1 \hdr_hld/high/U1659_1_/U5  ( .x(\hdr_hld/high/ncd[1] ), .a(itag_l
        [1]), .b(itag_h[1]) );
    nor2_1 \hdr_hld/high/U1659_2_/U5  ( .x(\hdr_hld/high/ncd[2] ), .a(itag_l
        [2]), .b(itag_h[2]) );
    nor2_1 \hdr_hld/high/U1659_3_/U5  ( .x(\hdr_hld/high/ncd[3] ), .a(itag_l
        [3]), .b(itag_h[3]) );
    nor2_1 \hdr_hld/high/U1659_4_/U5  ( .x(\hdr_hld/high/ncd[4] ), .a(itag_l
        [4]), .b(itag_h[4]) );
    nor2_1 \hdr_hld/high/U1659_5_/U5  ( .x(\hdr_hld/high/ncd[5] ), .a(col_l[0]
        ), .b(col_h[0]) );
    nor2_1 \hdr_hld/high/U1659_6_/U5  ( .x(\hdr_hld/high/ncd[6] ), .a(col_l[1]
        ), .b(col_h[1]) );
    nor2_1 \hdr_hld/high/U1659_7_/U5  ( .x(\hdr_hld/high/ncd[7] ), .a(col_l[2]
        ), .b(col_h[2]) );
    nor2_1 \hdr_hld/high/U3/U5  ( .x(\hdr_hld/high/ctrlack_internal ), .a(
        \hdr_hld/high/acb ), .b(\hdr_hld/high/ba ) );
    buf_2 \hdr_hld/high/U1665/U7  ( .x(\hdr_hld/high/driveh ), .a(receive) );
    buf_2 \hdr_hld/high/U1666/U7  ( .x(\hdr_hld/high/drivel ), .a(receive) );
    ao23_1 \hdr_hld/high/U1658_0_/U21/U1/U1  ( .x(itag_l[0]), .a(
        \hdr_hld/high/drivel ), .b(itag_l[0]), .c(\hdr_hld/high/drivel ), .d(
        chwl[0]), .e(n1) );
    ao23_1 \hdr_hld/high/U1658_1_/U21/U1/U1  ( .x(itag_l[1]), .a(
        \hdr_hld/high/drivel ), .b(itag_l[1]), .c(\hdr_hld/high/drivel ), .d(
        chwl[1]), .e(n1) );
    ao23_1 \hdr_hld/high/U1658_2_/U21/U1/U1  ( .x(itag_l[2]), .a(
        \hdr_hld/high/drivel ), .b(itag_l[2]), .c(\hdr_hld/high/drivel ), .d(
        chwl[2]), .e(n1) );
    ao23_1 \hdr_hld/high/U1658_3_/U21/U1/U1  ( .x(itag_l[3]), .a(
        \hdr_hld/high/drivel ), .b(itag_l[3]), .c(\hdr_hld/high/drivel ), .d(
        chwl[3]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1658_4_/U21/U1/U1  ( .x(itag_l[4]), .a(n4), .b(
        itag_l[4]), .c(\hdr_hld/high/drivel ), .d(chwl[4]), .e(
        \hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1658_5_/U21/U1/U1  ( .x(col_l[0]), .a(n4), .b(col_l
        [0]), .c(\hdr_hld/high/drivel ), .d(chwl[5]), .e(\hdr_hld/high/latch )
         );
    ao23_1 \hdr_hld/high/U1658_6_/U21/U1/U1  ( .x(col_l[1]), .a(
        \hdr_hld/high/drivel ), .b(col_l[1]), .c(\hdr_hld/high/drivel ), .d(
        chwl[6]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1658_7_/U21/U1/U1  ( .x(col_l[2]), .a(n4), .b(col_l
        [2]), .c(\hdr_hld/high/drivel ), .d(chwl[7]), .e(\hdr_hld/high/latch )
         );
    ao23_1 \hdr_hld/high/U1651_0_/U21/U1/U1  ( .x(itag_h[0]), .a(n2), .b(
        itag_h[0]), .c(n2), .d(chwh[0]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1651_1_/U21/U1/U1  ( .x(itag_h[1]), .a(n2), .b(
        itag_h[1]), .c(n3), .d(chwh[1]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1651_2_/U21/U1/U1  ( .x(itag_h[2]), .a(n2), .b(
        itag_h[2]), .c(n3), .d(chwh[2]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1651_3_/U21/U1/U1  ( .x(itag_h[3]), .a(n2), .b(
        itag_h[3]), .c(n3), .d(chwh[3]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1651_4_/U21/U1/U1  ( .x(itag_h[4]), .a(n2), .b(
        itag_h[4]), .c(n3), .d(chwh[4]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1651_5_/U21/U1/U1  ( .x(col_h[0]), .a(n2), .b(col_h
        [0]), .c(n3), .d(chwh[5]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1651_6_/U21/U1/U1  ( .x(col_h[1]), .a(n2), .b(col_h
        [1]), .c(n2), .d(chwh[6]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1651_7_/U21/U1/U1  ( .x(col_h[2]), .a(n2), .b(col_h
        [2]), .c(n2), .d(chwh[7]), .e(\hdr_hld/high/latch ) );
    aoai211_1 \hdr_hld/high/U4/U28/U1/U1  ( .x(\hdr_hld/high/U4/U28/U1/clr ), 
        .a(receive), .b(\hdr_hld/high/acb ), .c(\hdr_hld/high/nlocalcd ), .d(
        \hdr_hld/net33 ) );
    nand3_1 \hdr_hld/high/U4/U28/U1/U2  ( .x(\hdr_hld/high/U4/U28/U1/set ), 
        .a(\hdr_hld/high/nlocalcd ), .b(receive), .c(\hdr_hld/high/acb ) );
    nand2_2 \hdr_hld/high/U4/U28/U1/U3  ( .x(\hdr_hld/net33 ), .a(
        \hdr_hld/high/U4/U28/U1/clr ), .b(\hdr_hld/high/U4/U28/U1/set ) );
    oai21_1 \hdr_hld/high/U1/U30/U1/U1  ( .x(\hdr_hld/high/acb ), .a(
        \hdr_hld/high/U1/Z ), .b(\hdr_hld/high/ba ), .c(receive) );
    inv_1 \hdr_hld/high/U1/U30/U1/U2  ( .x(\hdr_hld/high/U1/Z ), .a(
        \hdr_hld/high/acb ) );
    ao222_1 \hdr_hld/high/U5/U18/U1/U1  ( .x(\hdr_hld/high/ba ), .a(
        \hdr_hld/high/latch ), .b(n9), .c(\hdr_hld/high/latch ), .d(
        \hdr_hld/high/ba ), .e(n9), .f(\hdr_hld/high/ba ) );
    aoi222_1 \hdr_hld/high/U1664/U28/U30/U1  ( .x(\hdr_hld/high/U1664/x[3] ), 
        .a(\hdr_hld/high/ncd[7] ), .b(\hdr_hld/high/ncd[6] ), .c(
        \hdr_hld/high/ncd[7] ), .d(\hdr_hld/high/U1664/U28/Z ), .e(
        \hdr_hld/high/ncd[6] ), .f(\hdr_hld/high/U1664/U28/Z ) );
    inv_1 \hdr_hld/high/U1664/U28/U30/Uinv  ( .x(\hdr_hld/high/U1664/U28/Z ), 
        .a(\hdr_hld/high/U1664/x[3] ) );
    aoi222_1 \hdr_hld/high/U1664/U32/U30/U1  ( .x(\hdr_hld/high/U1664/x[0] ), 
        .a(\hdr_hld/high/ncd[1] ), .b(\hdr_hld/high/ncd[0] ), .c(
        \hdr_hld/high/ncd[1] ), .d(\hdr_hld/high/U1664/U32/Z ), .e(
        \hdr_hld/high/ncd[0] ), .f(\hdr_hld/high/U1664/U32/Z ) );
    inv_1 \hdr_hld/high/U1664/U32/U30/Uinv  ( .x(\hdr_hld/high/U1664/U32/Z ), 
        .a(\hdr_hld/high/U1664/x[0] ) );
    aoi222_1 \hdr_hld/high/U1664/U29/U30/U1  ( .x(\hdr_hld/high/U1664/x[2] ), 
        .a(\hdr_hld/high/ncd[5] ), .b(\hdr_hld/high/ncd[4] ), .c(
        \hdr_hld/high/ncd[5] ), .d(\hdr_hld/high/U1664/U29/Z ), .e(
        \hdr_hld/high/ncd[4] ), .f(\hdr_hld/high/U1664/U29/Z ) );
    inv_1 \hdr_hld/high/U1664/U29/U30/Uinv  ( .x(\hdr_hld/high/U1664/U29/Z ), 
        .a(\hdr_hld/high/U1664/x[2] ) );
    aoi222_1 \hdr_hld/high/U1664/U33/U30/U1  ( .x(\hdr_hld/high/U1664/y[0] ), 
        .a(\hdr_hld/high/U1664/x[1] ), .b(\hdr_hld/high/U1664/x[0] ), .c(
        \hdr_hld/high/U1664/x[1] ), .d(\hdr_hld/high/U1664/U33/Z ), .e(
        \hdr_hld/high/U1664/x[0] ), .f(\hdr_hld/high/U1664/U33/Z ) );
    inv_1 \hdr_hld/high/U1664/U33/U30/Uinv  ( .x(\hdr_hld/high/U1664/U33/Z ), 
        .a(\hdr_hld/high/U1664/y[0] ) );
    aoi222_1 \hdr_hld/high/U1664/U30/U30/U1  ( .x(\hdr_hld/high/U1664/y[1] ), 
        .a(\hdr_hld/high/U1664/x[3] ), .b(\hdr_hld/high/U1664/x[2] ), .c(
        \hdr_hld/high/U1664/x[3] ), .d(\hdr_hld/high/U1664/U30/Z ), .e(
        \hdr_hld/high/U1664/x[2] ), .f(\hdr_hld/high/U1664/U30/Z ) );
    inv_1 \hdr_hld/high/U1664/U30/U30/Uinv  ( .x(\hdr_hld/high/U1664/U30/Z ), 
        .a(\hdr_hld/high/U1664/y[1] ) );
    aoi222_1 \hdr_hld/high/U1664/U31/U30/U1  ( .x(\hdr_hld/high/U1664/x[1] ), 
        .a(\hdr_hld/high/ncd[3] ), .b(\hdr_hld/high/ncd[2] ), .c(
        \hdr_hld/high/ncd[3] ), .d(\hdr_hld/high/U1664/U31/Z ), .e(
        \hdr_hld/high/ncd[2] ), .f(\hdr_hld/high/U1664/U31/Z ) );
    inv_1 \hdr_hld/high/U1664/U31/U30/Uinv  ( .x(\hdr_hld/high/U1664/U31/Z ), 
        .a(\hdr_hld/high/U1664/x[1] ) );
    aoi222_1 \hdr_hld/high/U1664/U37/U30/U1  ( .x(\hdr_hld/high/localcd ), .a(
        \hdr_hld/high/U1664/y[0] ), .b(\hdr_hld/high/U1664/y[1] ), .c(
        \hdr_hld/high/U1664/y[0] ), .d(\hdr_hld/high/U1664/U37/Z ), .e(
        \hdr_hld/high/U1664/y[1] ), .f(\hdr_hld/high/U1664/U37/Z ) );
    inv_1 \hdr_hld/high/U1664/U37/U30/Uinv  ( .x(\hdr_hld/high/U1664/U37/Z ), 
        .a(\hdr_hld/high/localcd ) );
    nor3_1 \hdr_hld/high/U1669/Unr  ( .x(\hdr_hld/high/U1669/nr ), .a(
        \hdr_hld/high/ctrlack_internal ), .b(\hdr_hld/high/drivel ), .c(n3) );
    nand3_1 \hdr_hld/high/U1669/Und  ( .x(\hdr_hld/high/U1669/nd ), .a(
        \hdr_hld/high/ctrlack_internal ), .b(\hdr_hld/high/drivel ), .c(n3) );
    oa21_1 \hdr_hld/high/U1669/U1  ( .x(\hdr_hld/high/U1669/n2 ), .a(
        \hdr_hld/high/U1669/n2 ), .b(\hdr_hld/high/U1669/nr ), .c(
        \hdr_hld/high/U1669/nd ) );
    inv_2 \hdr_hld/high/U1669/U3  ( .x(\hdr_hld/net20 ), .a(
        \hdr_hld/high/U1669/n2 ) );
    buf_1 U1 ( .x(n1), .a(\hdr_hld/high/latch ) );
    buf_3 U2 ( .x(n2), .a(\hdr_hld/high/driveh ) );
    buf_3 U3 ( .x(n3), .a(\hdr_hld/high/driveh ) );
    buf_1 U4 ( .x(n4), .a(\hdr_hld/high/drivel ) );
    buf_1 U5 ( .x(n5), .a(\hdr_hld/low/latch ) );
    buf_2 U6 ( .x(n7), .a(\hdr_hld/net20 ) );
    buf_2 U7 ( .x(n6), .a(\hdr_hld/net20 ) );
    inv_2 U8 ( .x(reset), .a(nReset) );
    buf_3 U9 ( .x(pullcd), .a(n9) );
endmodule


module chain_irdemux_32new_1 ( ctrlack, oh, ol, pullreq, pull_h, pull_l, 
    pullcd, reset, ctrlreq );
output [31:0] oh;
output [31:0] ol;
input  [7:0] pull_h;
input  [7:0] pull_l;
input  pullcd, reset, ctrlreq;
output ctrlack, pullreq;
    wire net30, net31, \I0/net32 , \I0/net33 , \I0/low/latch , 
        \I0/low/nlocalcd , \I0/low/localcd , \I0/low/ncd[0] , \I0/low/ncd[1] , 
        \I0/low/ncd[2] , \I0/low/ncd[3] , \I0/low/ncd[4] , \I0/low/ncd[5] , 
        \I0/low/ncd[6] , \I0/low/ncd[7] , \I0/low/ctrlack_internal , 
        \I0/low/acb , \I0/low/ba , \I0/low/driveh , \I0/net20 , 
        \I0/low/drivel , n12, n11, \I0/low/U4/U28/U1/clr , 
        \I0/low/U4/U28/U1/set , \I0/low/U1/Z , \I0/low/U1664/x[3] , 
        \I0/low/U1664/U28/Z , \I0/low/U1664/x[0] , \I0/low/U1664/U32/Z , 
        \I0/low/U1664/x[2] , \I0/low/U1664/U29/Z , \I0/low/U1664/y[0] , 
        \I0/low/U1664/x[1] , \I0/low/U1664/U33/Z , \I0/low/U1664/y[1] , 
        \I0/low/U1664/U30/Z , \I0/low/U1664/U31/Z , \I0/low/U1664/U37/Z , 
        \I0/low/U1669/nr , \I0/low/U1669/nd , \I0/low/U1669/n2 , 
        \I0/high/latch , \I0/high/nlocalcd , \I0/high/localcd , 
        \I0/high/ncd[0] , \I0/high/ncd[1] , \I0/high/ncd[2] , \I0/high/ncd[3] , 
        \I0/high/ncd[4] , \I0/high/ncd[5] , \I0/high/ncd[6] , \I0/high/ncd[7] , 
        \I0/high/ctrlack_internal , \I0/high/acb , \I0/high/ba , 
        \I0/high/driveh , net17, \I0/high/drivel , n10, n9, 
        \I0/high/U4/U28/U1/clr , \I0/high/U4/U28/U1/set , \I0/high/U1/Z , 
        \I0/high/U1664/x[3] , \I0/high/U1664/U28/Z , \I0/high/U1664/x[0] , 
        \I0/high/U1664/U32/Z , \I0/high/U1664/x[2] , \I0/high/U1664/U29/Z , 
        \I0/high/U1664/y[0] , \I0/high/U1664/x[1] , \I0/high/U1664/U33/Z , 
        \I0/high/U1664/y[1] , \I0/high/U1664/U30/Z , \I0/high/U1664/U31/Z , 
        \I0/high/U1664/U37/Z , \I0/high/U1669/nr , \I0/high/U1669/nd , 
        \I0/high/U1669/n2 , \I1/net32 , \I1/net33 , \I1/low/latch , 
        \I1/low/nlocalcd , \I1/low/localcd , \I1/low/ncd[0] , \I1/low/ncd[1] , 
        \I1/low/ncd[2] , \I1/low/ncd[3] , \I1/low/ncd[4] , \I1/low/ncd[5] , 
        \I1/low/ncd[6] , \I1/low/ncd[7] , \I1/low/ctrlack_internal , 
        \I1/low/acb , \I1/low/ba , \I1/low/driveh , \I1/net20 , 
        \I1/low/drivel , n8, n7, \I1/low/U4/U28/U1/clr , 
        \I1/low/U4/U28/U1/set , \I1/low/U1/Z , \I1/low/U1664/x[3] , 
        \I1/low/U1664/U28/Z , \I1/low/U1664/x[0] , \I1/low/U1664/U32/Z , 
        \I1/low/U1664/x[2] , \I1/low/U1664/U29/Z , \I1/low/U1664/y[0] , 
        \I1/low/U1664/x[1] , \I1/low/U1664/U33/Z , \I1/low/U1664/y[1] , 
        \I1/low/U1664/U30/Z , \I1/low/U1664/U31/Z , \I1/low/U1664/U37/Z , 
        \I1/low/U1669/nr , \I1/low/U1669/nd , \I1/low/U1669/n2 , 
        \I1/high/latch , \I1/high/nlocalcd , \I1/high/localcd , 
        \I1/high/ncd[0] , \I1/high/ncd[1] , \I1/high/ncd[2] , \I1/high/ncd[3] , 
        \I1/high/ncd[4] , \I1/high/ncd[5] , \I1/high/ncd[6] , \I1/high/ncd[7] , 
        \I1/high/ctrlack_internal , \I1/high/acb , \I1/high/ba , n5, n6, n1, 
        n2, n3, \I1/high/U4/U28/U1/clr , \I1/high/U4/U28/U1/set , 
        \I1/high/U1/Z , \I1/high/U1664/x[3] , \I1/high/U1664/U28/Z , 
        \I1/high/U1664/x[0] , \I1/high/U1664/U32/Z , \I1/high/U1664/x[2] , 
        \I1/high/U1664/U29/Z , \I1/high/U1664/y[0] , \I1/high/U1664/x[1] , 
        \I1/high/U1664/U33/Z , \I1/high/U1664/y[1] , \I1/high/U1664/U30/Z , 
        \I1/high/U1664/U31/Z , \I1/high/U1664/U37/Z , \I1/high/U1669/nr , 
        \I1/high/U1669/nd , \I1/high/U1669/n2 , n4;
    nand2_1 \U3/U5  ( .x(pullreq), .a(net30), .b(net31) );
    nor2_1 \I0/U3/U5  ( .x(net30), .a(\I0/net32 ), .b(\I0/net33 ) );
    buf_2 \I0/low/U1653  ( .x(\I0/low/latch ), .a(\I0/net32 ) );
    nor2_1 \I0/low/U264/U5  ( .x(\I0/low/nlocalcd ), .a(reset), .b(
        \I0/low/localcd ) );
    nor2_1 \I0/low/U1659_0_/U5  ( .x(\I0/low/ncd[0] ), .a(ol[0]), .b(oh[0]) );
    nor2_1 \I0/low/U1659_1_/U5  ( .x(\I0/low/ncd[1] ), .a(ol[1]), .b(oh[1]) );
    nor2_1 \I0/low/U1659_2_/U5  ( .x(\I0/low/ncd[2] ), .a(ol[2]), .b(oh[2]) );
    nor2_1 \I0/low/U1659_3_/U5  ( .x(\I0/low/ncd[3] ), .a(ol[3]), .b(oh[3]) );
    nor2_1 \I0/low/U1659_4_/U5  ( .x(\I0/low/ncd[4] ), .a(ol[4]), .b(oh[4]) );
    nor2_1 \I0/low/U1659_5_/U5  ( .x(\I0/low/ncd[5] ), .a(ol[5]), .b(oh[5]) );
    nor2_1 \I0/low/U1659_6_/U5  ( .x(\I0/low/ncd[6] ), .a(ol[6]), .b(oh[6]) );
    nor2_1 \I0/low/U1659_7_/U5  ( .x(\I0/low/ncd[7] ), .a(ol[7]), .b(oh[7]) );
    nor2_1 \I0/low/U3/U5  ( .x(\I0/low/ctrlack_internal ), .a(\I0/low/acb ), 
        .b(\I0/low/ba ) );
    buf_2 \I0/low/U1665/U7  ( .x(\I0/low/driveh ), .a(\I0/net20 ) );
    buf_2 \I0/low/U1666/U7  ( .x(\I0/low/drivel ), .a(\I0/net20 ) );
    ao23_1 \I0/low/U1658_0_/U21/U1/U1  ( .x(ol[0]), .a(n12), .b(ol[0]), .c(
        \I0/low/drivel ), .d(pull_l[0]), .e(n11) );
    ao23_1 \I0/low/U1658_1_/U21/U1/U1  ( .x(ol[1]), .a(n12), .b(ol[1]), .c(
        \I0/low/driveh ), .d(pull_l[1]), .e(n11) );
    ao23_1 \I0/low/U1658_2_/U21/U1/U1  ( .x(ol[2]), .a(\I0/low/driveh ), .b(ol
        [2]), .c(n12), .d(pull_l[2]), .e(n11) );
    ao23_1 \I0/low/U1658_3_/U21/U1/U1  ( .x(ol[3]), .a(n12), .b(ol[3]), .c(
        \I0/low/driveh ), .d(pull_l[3]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_4_/U21/U1/U1  ( .x(ol[4]), .a(\I0/low/drivel ), .b(ol
        [4]), .c(n12), .d(pull_l[4]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_5_/U21/U1/U1  ( .x(ol[5]), .a(\I0/low/drivel ), .b(ol
        [5]), .c(n12), .d(pull_l[5]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_6_/U21/U1/U1  ( .x(ol[6]), .a(\I0/low/driveh ), .b(ol
        [6]), .c(\I0/low/drivel ), .d(pull_l[6]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_7_/U21/U1/U1  ( .x(ol[7]), .a(\I0/low/driveh ), .b(ol
        [7]), .c(\I0/low/driveh ), .d(pull_l[7]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_0_/U21/U1/U1  ( .x(oh[0]), .a(\I0/low/drivel ), .b(oh
        [0]), .c(n12), .d(pull_h[0]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_1_/U21/U1/U1  ( .x(oh[1]), .a(\I0/low/driveh ), .b(oh
        [1]), .c(\I0/low/drivel ), .d(pull_h[1]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_2_/U21/U1/U1  ( .x(oh[2]), .a(\I0/low/drivel ), .b(oh
        [2]), .c(\I0/low/drivel ), .d(pull_h[2]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_3_/U21/U1/U1  ( .x(oh[3]), .a(\I0/low/driveh ), .b(oh
        [3]), .c(\I0/low/driveh ), .d(pull_h[3]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_4_/U21/U1/U1  ( .x(oh[4]), .a(\I0/low/drivel ), .b(oh
        [4]), .c(\I0/low/driveh ), .d(pull_h[4]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_5_/U21/U1/U1  ( .x(oh[5]), .a(\I0/low/driveh ), .b(oh
        [5]), .c(n12), .d(pull_h[5]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_6_/U21/U1/U1  ( .x(oh[6]), .a(n12), .b(oh[6]), .c(
        \I0/low/drivel ), .d(pull_h[6]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_7_/U21/U1/U1  ( .x(oh[7]), .a(n12), .b(oh[7]), .c(n12
        ), .d(pull_h[7]), .e(\I0/low/latch ) );
    aoai211_1 \I0/low/U4/U28/U1/U1  ( .x(\I0/low/U4/U28/U1/clr ), .a(
        \I0/net20 ), .b(\I0/low/acb ), .c(\I0/low/nlocalcd ), .d(\I0/net32 )
         );
    nand3_1 \I0/low/U4/U28/U1/U2  ( .x(\I0/low/U4/U28/U1/set ), .a(
        \I0/low/nlocalcd ), .b(\I0/net20 ), .c(\I0/low/acb ) );
    nand2_2 \I0/low/U4/U28/U1/U3  ( .x(\I0/net32 ), .a(\I0/low/U4/U28/U1/clr ), 
        .b(\I0/low/U4/U28/U1/set ) );
    oai21_1 \I0/low/U1/U30/U1/U1  ( .x(\I0/low/acb ), .a(\I0/low/U1/Z ), .b(
        \I0/low/ba ), .c(\I0/net20 ) );
    inv_1 \I0/low/U1/U30/U1/U2  ( .x(\I0/low/U1/Z ), .a(\I0/low/acb ) );
    ao222_1 \I0/low/U5/U18/U1/U1  ( .x(\I0/low/ba ), .a(\I0/low/latch ), .b(
        pullcd), .c(\I0/low/latch ), .d(\I0/low/ba ), .e(pullcd), .f(
        \I0/low/ba ) );
    aoi222_1 \I0/low/U1664/U28/U30/U1  ( .x(\I0/low/U1664/x[3] ), .a(
        \I0/low/ncd[7] ), .b(\I0/low/ncd[6] ), .c(\I0/low/ncd[7] ), .d(
        \I0/low/U1664/U28/Z ), .e(\I0/low/ncd[6] ), .f(\I0/low/U1664/U28/Z )
         );
    inv_1 \I0/low/U1664/U28/U30/Uinv  ( .x(\I0/low/U1664/U28/Z ), .a(
        \I0/low/U1664/x[3] ) );
    aoi222_1 \I0/low/U1664/U32/U30/U1  ( .x(\I0/low/U1664/x[0] ), .a(
        \I0/low/ncd[1] ), .b(\I0/low/ncd[0] ), .c(\I0/low/ncd[1] ), .d(
        \I0/low/U1664/U32/Z ), .e(\I0/low/ncd[0] ), .f(\I0/low/U1664/U32/Z )
         );
    inv_1 \I0/low/U1664/U32/U30/Uinv  ( .x(\I0/low/U1664/U32/Z ), .a(
        \I0/low/U1664/x[0] ) );
    aoi222_1 \I0/low/U1664/U29/U30/U1  ( .x(\I0/low/U1664/x[2] ), .a(
        \I0/low/ncd[5] ), .b(\I0/low/ncd[4] ), .c(\I0/low/ncd[5] ), .d(
        \I0/low/U1664/U29/Z ), .e(\I0/low/ncd[4] ), .f(\I0/low/U1664/U29/Z )
         );
    inv_1 \I0/low/U1664/U29/U30/Uinv  ( .x(\I0/low/U1664/U29/Z ), .a(
        \I0/low/U1664/x[2] ) );
    aoi222_1 \I0/low/U1664/U33/U30/U1  ( .x(\I0/low/U1664/y[0] ), .a(
        \I0/low/U1664/x[1] ), .b(\I0/low/U1664/x[0] ), .c(\I0/low/U1664/x[1] ), 
        .d(\I0/low/U1664/U33/Z ), .e(\I0/low/U1664/x[0] ), .f(
        \I0/low/U1664/U33/Z ) );
    inv_1 \I0/low/U1664/U33/U30/Uinv  ( .x(\I0/low/U1664/U33/Z ), .a(
        \I0/low/U1664/y[0] ) );
    aoi222_1 \I0/low/U1664/U30/U30/U1  ( .x(\I0/low/U1664/y[1] ), .a(
        \I0/low/U1664/x[3] ), .b(\I0/low/U1664/x[2] ), .c(\I0/low/U1664/x[3] ), 
        .d(\I0/low/U1664/U30/Z ), .e(\I0/low/U1664/x[2] ), .f(
        \I0/low/U1664/U30/Z ) );
    inv_1 \I0/low/U1664/U30/U30/Uinv  ( .x(\I0/low/U1664/U30/Z ), .a(
        \I0/low/U1664/y[1] ) );
    aoi222_1 \I0/low/U1664/U31/U30/U1  ( .x(\I0/low/U1664/x[1] ), .a(
        \I0/low/ncd[3] ), .b(\I0/low/ncd[2] ), .c(\I0/low/ncd[3] ), .d(
        \I0/low/U1664/U31/Z ), .e(\I0/low/ncd[2] ), .f(\I0/low/U1664/U31/Z )
         );
    inv_1 \I0/low/U1664/U31/U30/Uinv  ( .x(\I0/low/U1664/U31/Z ), .a(
        \I0/low/U1664/x[1] ) );
    aoi222_1 \I0/low/U1664/U37/U30/U1  ( .x(\I0/low/localcd ), .a(
        \I0/low/U1664/y[0] ), .b(\I0/low/U1664/y[1] ), .c(\I0/low/U1664/y[0] ), 
        .d(\I0/low/U1664/U37/Z ), .e(\I0/low/U1664/y[1] ), .f(
        \I0/low/U1664/U37/Z ) );
    inv_1 \I0/low/U1664/U37/U30/Uinv  ( .x(\I0/low/U1664/U37/Z ), .a(
        \I0/low/localcd ) );
    nor3_1 \I0/low/U1669/Unr  ( .x(\I0/low/U1669/nr ), .a(
        \I0/low/ctrlack_internal ), .b(n12), .c(\I0/low/drivel ) );
    nand3_1 \I0/low/U1669/Und  ( .x(\I0/low/U1669/nd ), .a(
        \I0/low/ctrlack_internal ), .b(\I0/low/driveh ), .c(\I0/low/drivel )
         );
    oa21_1 \I0/low/U1669/U1  ( .x(\I0/low/U1669/n2 ), .a(\I0/low/U1669/n2 ), 
        .b(\I0/low/U1669/nr ), .c(\I0/low/U1669/nd ) );
    inv_2 \I0/low/U1669/U3  ( .x(ctrlack), .a(\I0/low/U1669/n2 ) );
    buf_2 \I0/high/U1653  ( .x(\I0/high/latch ), .a(\I0/net33 ) );
    nor2_1 \I0/high/U264/U5  ( .x(\I0/high/nlocalcd ), .a(reset), .b(
        \I0/high/localcd ) );
    nor2_1 \I0/high/U1659_0_/U5  ( .x(\I0/high/ncd[0] ), .a(ol[8]), .b(oh[8])
         );
    nor2_1 \I0/high/U1659_1_/U5  ( .x(\I0/high/ncd[1] ), .a(ol[9]), .b(oh[9])
         );
    nor2_1 \I0/high/U1659_2_/U5  ( .x(\I0/high/ncd[2] ), .a(ol[10]), .b(oh[10]
        ) );
    nor2_1 \I0/high/U1659_3_/U5  ( .x(\I0/high/ncd[3] ), .a(ol[11]), .b(oh[11]
        ) );
    nor2_1 \I0/high/U1659_4_/U5  ( .x(\I0/high/ncd[4] ), .a(ol[12]), .b(oh[12]
        ) );
    nor2_1 \I0/high/U1659_5_/U5  ( .x(\I0/high/ncd[5] ), .a(ol[13]), .b(oh[13]
        ) );
    nor2_1 \I0/high/U1659_6_/U5  ( .x(\I0/high/ncd[6] ), .a(ol[14]), .b(oh[14]
        ) );
    nor2_1 \I0/high/U1659_7_/U5  ( .x(\I0/high/ncd[7] ), .a(ol[15]), .b(oh[15]
        ) );
    nor2_1 \I0/high/U3/U5  ( .x(\I0/high/ctrlack_internal ), .a(\I0/high/acb ), 
        .b(\I0/high/ba ) );
    buf_2 \I0/high/U1665/U7  ( .x(\I0/high/driveh ), .a(net17) );
    buf_2 \I0/high/U1666/U7  ( .x(\I0/high/drivel ), .a(net17) );
    ao23_1 \I0/high/U1658_0_/U21/U1/U1  ( .x(ol[8]), .a(n10), .b(ol[8]), .c(
        \I0/high/drivel ), .d(pull_l[0]), .e(n9) );
    ao23_1 \I0/high/U1658_1_/U21/U1/U1  ( .x(ol[9]), .a(n10), .b(ol[9]), .c(
        \I0/high/driveh ), .d(pull_l[1]), .e(n9) );
    ao23_1 \I0/high/U1658_2_/U21/U1/U1  ( .x(ol[10]), .a(\I0/high/driveh ), 
        .b(ol[10]), .c(n10), .d(pull_l[2]), .e(n9) );
    ao23_1 \I0/high/U1658_3_/U21/U1/U1  ( .x(ol[11]), .a(n10), .b(ol[11]), .c(
        \I0/high/driveh ), .d(pull_l[3]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1658_4_/U21/U1/U1  ( .x(ol[12]), .a(\I0/high/drivel ), 
        .b(ol[12]), .c(n10), .d(pull_l[4]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1658_5_/U21/U1/U1  ( .x(ol[13]), .a(\I0/high/drivel ), 
        .b(ol[13]), .c(n10), .d(pull_l[5]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1658_6_/U21/U1/U1  ( .x(ol[14]), .a(\I0/high/driveh ), 
        .b(ol[14]), .c(\I0/high/drivel ), .d(pull_l[6]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1658_7_/U21/U1/U1  ( .x(ol[15]), .a(\I0/high/driveh ), 
        .b(ol[15]), .c(\I0/high/driveh ), .d(pull_l[7]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1651_0_/U21/U1/U1  ( .x(oh[8]), .a(\I0/high/drivel ), .b(
        oh[8]), .c(n10), .d(pull_h[0]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_1_/U21/U1/U1  ( .x(oh[9]), .a(\I0/high/driveh ), .b(
        oh[9]), .c(\I0/high/drivel ), .d(pull_h[1]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_2_/U21/U1/U1  ( .x(oh[10]), .a(\I0/high/drivel ), 
        .b(oh[10]), .c(\I0/high/drivel ), .d(pull_h[2]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1651_3_/U21/U1/U1  ( .x(oh[11]), .a(\I0/high/driveh ), 
        .b(oh[11]), .c(\I0/high/driveh ), .d(pull_h[3]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1651_4_/U21/U1/U1  ( .x(oh[12]), .a(\I0/high/drivel ), 
        .b(oh[12]), .c(\I0/high/driveh ), .d(pull_h[4]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1651_5_/U21/U1/U1  ( .x(oh[13]), .a(\I0/high/driveh ), 
        .b(oh[13]), .c(n10), .d(pull_h[5]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_6_/U21/U1/U1  ( .x(oh[14]), .a(n10), .b(oh[14]), .c(
        \I0/high/drivel ), .d(pull_h[6]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_7_/U21/U1/U1  ( .x(oh[15]), .a(n10), .b(oh[15]), .c(
        n10), .d(pull_h[7]), .e(\I0/high/latch ) );
    aoai211_1 \I0/high/U4/U28/U1/U1  ( .x(\I0/high/U4/U28/U1/clr ), .a(net17), 
        .b(\I0/high/acb ), .c(\I0/high/nlocalcd ), .d(\I0/net33 ) );
    nand3_1 \I0/high/U4/U28/U1/U2  ( .x(\I0/high/U4/U28/U1/set ), .a(
        \I0/high/nlocalcd ), .b(net17), .c(\I0/high/acb ) );
    nand2_2 \I0/high/U4/U28/U1/U3  ( .x(\I0/net33 ), .a(
        \I0/high/U4/U28/U1/clr ), .b(\I0/high/U4/U28/U1/set ) );
    oai21_1 \I0/high/U1/U30/U1/U1  ( .x(\I0/high/acb ), .a(\I0/high/U1/Z ), 
        .b(\I0/high/ba ), .c(net17) );
    inv_1 \I0/high/U1/U30/U1/U2  ( .x(\I0/high/U1/Z ), .a(\I0/high/acb ) );
    ao222_1 \I0/high/U5/U18/U1/U1  ( .x(\I0/high/ba ), .a(\I0/high/latch ), 
        .b(pullcd), .c(\I0/high/latch ), .d(\I0/high/ba ), .e(pullcd), .f(
        \I0/high/ba ) );
    aoi222_1 \I0/high/U1664/U28/U30/U1  ( .x(\I0/high/U1664/x[3] ), .a(
        \I0/high/ncd[7] ), .b(\I0/high/ncd[6] ), .c(\I0/high/ncd[7] ), .d(
        \I0/high/U1664/U28/Z ), .e(\I0/high/ncd[6] ), .f(\I0/high/U1664/U28/Z 
        ) );
    inv_1 \I0/high/U1664/U28/U30/Uinv  ( .x(\I0/high/U1664/U28/Z ), .a(
        \I0/high/U1664/x[3] ) );
    aoi222_1 \I0/high/U1664/U32/U30/U1  ( .x(\I0/high/U1664/x[0] ), .a(
        \I0/high/ncd[1] ), .b(\I0/high/ncd[0] ), .c(\I0/high/ncd[1] ), .d(
        \I0/high/U1664/U32/Z ), .e(\I0/high/ncd[0] ), .f(\I0/high/U1664/U32/Z 
        ) );
    inv_1 \I0/high/U1664/U32/U30/Uinv  ( .x(\I0/high/U1664/U32/Z ), .a(
        \I0/high/U1664/x[0] ) );
    aoi222_1 \I0/high/U1664/U29/U30/U1  ( .x(\I0/high/U1664/x[2] ), .a(
        \I0/high/ncd[5] ), .b(\I0/high/ncd[4] ), .c(\I0/high/ncd[5] ), .d(
        \I0/high/U1664/U29/Z ), .e(\I0/high/ncd[4] ), .f(\I0/high/U1664/U29/Z 
        ) );
    inv_1 \I0/high/U1664/U29/U30/Uinv  ( .x(\I0/high/U1664/U29/Z ), .a(
        \I0/high/U1664/x[2] ) );
    aoi222_1 \I0/high/U1664/U33/U30/U1  ( .x(\I0/high/U1664/y[0] ), .a(
        \I0/high/U1664/x[1] ), .b(\I0/high/U1664/x[0] ), .c(
        \I0/high/U1664/x[1] ), .d(\I0/high/U1664/U33/Z ), .e(
        \I0/high/U1664/x[0] ), .f(\I0/high/U1664/U33/Z ) );
    inv_1 \I0/high/U1664/U33/U30/Uinv  ( .x(\I0/high/U1664/U33/Z ), .a(
        \I0/high/U1664/y[0] ) );
    aoi222_1 \I0/high/U1664/U30/U30/U1  ( .x(\I0/high/U1664/y[1] ), .a(
        \I0/high/U1664/x[3] ), .b(\I0/high/U1664/x[2] ), .c(
        \I0/high/U1664/x[3] ), .d(\I0/high/U1664/U30/Z ), .e(
        \I0/high/U1664/x[2] ), .f(\I0/high/U1664/U30/Z ) );
    inv_1 \I0/high/U1664/U30/U30/Uinv  ( .x(\I0/high/U1664/U30/Z ), .a(
        \I0/high/U1664/y[1] ) );
    aoi222_1 \I0/high/U1664/U31/U30/U1  ( .x(\I0/high/U1664/x[1] ), .a(
        \I0/high/ncd[3] ), .b(\I0/high/ncd[2] ), .c(\I0/high/ncd[3] ), .d(
        \I0/high/U1664/U31/Z ), .e(\I0/high/ncd[2] ), .f(\I0/high/U1664/U31/Z 
        ) );
    inv_1 \I0/high/U1664/U31/U30/Uinv  ( .x(\I0/high/U1664/U31/Z ), .a(
        \I0/high/U1664/x[1] ) );
    aoi222_1 \I0/high/U1664/U37/U30/U1  ( .x(\I0/high/localcd ), .a(
        \I0/high/U1664/y[0] ), .b(\I0/high/U1664/y[1] ), .c(
        \I0/high/U1664/y[0] ), .d(\I0/high/U1664/U37/Z ), .e(
        \I0/high/U1664/y[1] ), .f(\I0/high/U1664/U37/Z ) );
    inv_1 \I0/high/U1664/U37/U30/Uinv  ( .x(\I0/high/U1664/U37/Z ), .a(
        \I0/high/localcd ) );
    nor3_1 \I0/high/U1669/Unr  ( .x(\I0/high/U1669/nr ), .a(
        \I0/high/ctrlack_internal ), .b(n10), .c(\I0/high/drivel ) );
    nand3_1 \I0/high/U1669/Und  ( .x(\I0/high/U1669/nd ), .a(
        \I0/high/ctrlack_internal ), .b(\I0/high/driveh ), .c(\I0/high/drivel 
        ) );
    oa21_1 \I0/high/U1669/U1  ( .x(\I0/high/U1669/n2 ), .a(\I0/high/U1669/n2 ), 
        .b(\I0/high/U1669/nr ), .c(\I0/high/U1669/nd ) );
    inv_2 \I0/high/U1669/U3  ( .x(\I0/net20 ), .a(\I0/high/U1669/n2 ) );
    nor2_1 \I1/U3/U5  ( .x(net31), .a(\I1/net32 ), .b(\I1/net33 ) );
    buf_2 \I1/low/U1653  ( .x(\I1/low/latch ), .a(\I1/net32 ) );
    nor2_1 \I1/low/U264/U5  ( .x(\I1/low/nlocalcd ), .a(reset), .b(
        \I1/low/localcd ) );
    nor2_1 \I1/low/U1659_0_/U5  ( .x(\I1/low/ncd[0] ), .a(ol[16]), .b(oh[16])
         );
    nor2_1 \I1/low/U1659_1_/U5  ( .x(\I1/low/ncd[1] ), .a(ol[17]), .b(oh[17])
         );
    nor2_1 \I1/low/U1659_2_/U5  ( .x(\I1/low/ncd[2] ), .a(ol[18]), .b(oh[18])
         );
    nor2_1 \I1/low/U1659_3_/U5  ( .x(\I1/low/ncd[3] ), .a(ol[19]), .b(oh[19])
         );
    nor2_1 \I1/low/U1659_4_/U5  ( .x(\I1/low/ncd[4] ), .a(ol[20]), .b(oh[20])
         );
    nor2_1 \I1/low/U1659_5_/U5  ( .x(\I1/low/ncd[5] ), .a(ol[21]), .b(oh[21])
         );
    nor2_1 \I1/low/U1659_6_/U5  ( .x(\I1/low/ncd[6] ), .a(ol[22]), .b(oh[22])
         );
    nor2_1 \I1/low/U1659_7_/U5  ( .x(\I1/low/ncd[7] ), .a(ol[23]), .b(oh[23])
         );
    nor2_1 \I1/low/U3/U5  ( .x(\I1/low/ctrlack_internal ), .a(\I1/low/acb ), 
        .b(\I1/low/ba ) );
    buf_2 \I1/low/U1665/U7  ( .x(\I1/low/driveh ), .a(\I1/net20 ) );
    buf_2 \I1/low/U1666/U7  ( .x(\I1/low/drivel ), .a(\I1/net20 ) );
    ao23_1 \I1/low/U1658_0_/U21/U1/U1  ( .x(ol[16]), .a(n8), .b(ol[16]), .c(
        \I1/low/drivel ), .d(pull_l[0]), .e(n7) );
    ao23_1 \I1/low/U1658_1_/U21/U1/U1  ( .x(ol[17]), .a(n8), .b(ol[17]), .c(
        \I1/low/driveh ), .d(pull_l[1]), .e(n7) );
    ao23_1 \I1/low/U1658_2_/U21/U1/U1  ( .x(ol[18]), .a(\I1/low/driveh ), .b(
        ol[18]), .c(n8), .d(pull_l[2]), .e(n7) );
    ao23_1 \I1/low/U1658_3_/U21/U1/U1  ( .x(ol[19]), .a(n8), .b(ol[19]), .c(
        \I1/low/driveh ), .d(pull_l[3]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_4_/U21/U1/U1  ( .x(ol[20]), .a(\I1/low/drivel ), .b(
        ol[20]), .c(n8), .d(pull_l[4]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_5_/U21/U1/U1  ( .x(ol[21]), .a(\I1/low/drivel ), .b(
        ol[21]), .c(n8), .d(pull_l[5]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_6_/U21/U1/U1  ( .x(ol[22]), .a(\I1/low/driveh ), .b(
        ol[22]), .c(\I1/low/drivel ), .d(pull_l[6]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_7_/U21/U1/U1  ( .x(ol[23]), .a(\I1/low/driveh ), .b(
        ol[23]), .c(\I1/low/driveh ), .d(pull_l[7]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_0_/U21/U1/U1  ( .x(oh[16]), .a(\I1/low/drivel ), .b(
        oh[16]), .c(n8), .d(pull_h[0]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_1_/U21/U1/U1  ( .x(oh[17]), .a(\I1/low/driveh ), .b(
        oh[17]), .c(\I1/low/drivel ), .d(pull_h[1]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_2_/U21/U1/U1  ( .x(oh[18]), .a(\I1/low/drivel ), .b(
        oh[18]), .c(\I1/low/drivel ), .d(pull_h[2]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_3_/U21/U1/U1  ( .x(oh[19]), .a(\I1/low/driveh ), .b(
        oh[19]), .c(\I1/low/driveh ), .d(pull_h[3]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_4_/U21/U1/U1  ( .x(oh[20]), .a(\I1/low/drivel ), .b(
        oh[20]), .c(\I1/low/driveh ), .d(pull_h[4]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_5_/U21/U1/U1  ( .x(oh[21]), .a(\I1/low/driveh ), .b(
        oh[21]), .c(n8), .d(pull_h[5]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_6_/U21/U1/U1  ( .x(oh[22]), .a(n8), .b(oh[22]), .c(
        \I1/low/drivel ), .d(pull_h[6]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_7_/U21/U1/U1  ( .x(oh[23]), .a(n8), .b(oh[23]), .c(n8
        ), .d(pull_h[7]), .e(\I1/low/latch ) );
    aoai211_1 \I1/low/U4/U28/U1/U1  ( .x(\I1/low/U4/U28/U1/clr ), .a(
        \I1/net20 ), .b(\I1/low/acb ), .c(\I1/low/nlocalcd ), .d(\I1/net32 )
         );
    nand3_1 \I1/low/U4/U28/U1/U2  ( .x(\I1/low/U4/U28/U1/set ), .a(
        \I1/low/nlocalcd ), .b(\I1/net20 ), .c(\I1/low/acb ) );
    nand2_2 \I1/low/U4/U28/U1/U3  ( .x(\I1/net32 ), .a(\I1/low/U4/U28/U1/clr ), 
        .b(\I1/low/U4/U28/U1/set ) );
    oai21_1 \I1/low/U1/U30/U1/U1  ( .x(\I1/low/acb ), .a(\I1/low/U1/Z ), .b(
        \I1/low/ba ), .c(\I1/net20 ) );
    inv_1 \I1/low/U1/U30/U1/U2  ( .x(\I1/low/U1/Z ), .a(\I1/low/acb ) );
    ao222_1 \I1/low/U5/U18/U1/U1  ( .x(\I1/low/ba ), .a(\I1/low/latch ), .b(
        pullcd), .c(\I1/low/latch ), .d(\I1/low/ba ), .e(pullcd), .f(
        \I1/low/ba ) );
    aoi222_1 \I1/low/U1664/U28/U30/U1  ( .x(\I1/low/U1664/x[3] ), .a(
        \I1/low/ncd[7] ), .b(\I1/low/ncd[6] ), .c(\I1/low/ncd[7] ), .d(
        \I1/low/U1664/U28/Z ), .e(\I1/low/ncd[6] ), .f(\I1/low/U1664/U28/Z )
         );
    inv_1 \I1/low/U1664/U28/U30/Uinv  ( .x(\I1/low/U1664/U28/Z ), .a(
        \I1/low/U1664/x[3] ) );
    aoi222_1 \I1/low/U1664/U32/U30/U1  ( .x(\I1/low/U1664/x[0] ), .a(
        \I1/low/ncd[1] ), .b(\I1/low/ncd[0] ), .c(\I1/low/ncd[1] ), .d(
        \I1/low/U1664/U32/Z ), .e(\I1/low/ncd[0] ), .f(\I1/low/U1664/U32/Z )
         );
    inv_1 \I1/low/U1664/U32/U30/Uinv  ( .x(\I1/low/U1664/U32/Z ), .a(
        \I1/low/U1664/x[0] ) );
    aoi222_1 \I1/low/U1664/U29/U30/U1  ( .x(\I1/low/U1664/x[2] ), .a(
        \I1/low/ncd[5] ), .b(\I1/low/ncd[4] ), .c(\I1/low/ncd[5] ), .d(
        \I1/low/U1664/U29/Z ), .e(\I1/low/ncd[4] ), .f(\I1/low/U1664/U29/Z )
         );
    inv_1 \I1/low/U1664/U29/U30/Uinv  ( .x(\I1/low/U1664/U29/Z ), .a(
        \I1/low/U1664/x[2] ) );
    aoi222_1 \I1/low/U1664/U33/U30/U1  ( .x(\I1/low/U1664/y[0] ), .a(
        \I1/low/U1664/x[1] ), .b(\I1/low/U1664/x[0] ), .c(\I1/low/U1664/x[1] ), 
        .d(\I1/low/U1664/U33/Z ), .e(\I1/low/U1664/x[0] ), .f(
        \I1/low/U1664/U33/Z ) );
    inv_1 \I1/low/U1664/U33/U30/Uinv  ( .x(\I1/low/U1664/U33/Z ), .a(
        \I1/low/U1664/y[0] ) );
    aoi222_1 \I1/low/U1664/U30/U30/U1  ( .x(\I1/low/U1664/y[1] ), .a(
        \I1/low/U1664/x[3] ), .b(\I1/low/U1664/x[2] ), .c(\I1/low/U1664/x[3] ), 
        .d(\I1/low/U1664/U30/Z ), .e(\I1/low/U1664/x[2] ), .f(
        \I1/low/U1664/U30/Z ) );
    inv_1 \I1/low/U1664/U30/U30/Uinv  ( .x(\I1/low/U1664/U30/Z ), .a(
        \I1/low/U1664/y[1] ) );
    aoi222_1 \I1/low/U1664/U31/U30/U1  ( .x(\I1/low/U1664/x[1] ), .a(
        \I1/low/ncd[3] ), .b(\I1/low/ncd[2] ), .c(\I1/low/ncd[3] ), .d(
        \I1/low/U1664/U31/Z ), .e(\I1/low/ncd[2] ), .f(\I1/low/U1664/U31/Z )
         );
    inv_1 \I1/low/U1664/U31/U30/Uinv  ( .x(\I1/low/U1664/U31/Z ), .a(
        \I1/low/U1664/x[1] ) );
    aoi222_1 \I1/low/U1664/U37/U30/U1  ( .x(\I1/low/localcd ), .a(
        \I1/low/U1664/y[0] ), .b(\I1/low/U1664/y[1] ), .c(\I1/low/U1664/y[0] ), 
        .d(\I1/low/U1664/U37/Z ), .e(\I1/low/U1664/y[1] ), .f(
        \I1/low/U1664/U37/Z ) );
    inv_1 \I1/low/U1664/U37/U30/Uinv  ( .x(\I1/low/U1664/U37/Z ), .a(
        \I1/low/localcd ) );
    nor3_1 \I1/low/U1669/Unr  ( .x(\I1/low/U1669/nr ), .a(
        \I1/low/ctrlack_internal ), .b(n8), .c(\I1/low/drivel ) );
    nand3_1 \I1/low/U1669/Und  ( .x(\I1/low/U1669/nd ), .a(
        \I1/low/ctrlack_internal ), .b(\I1/low/driveh ), .c(\I1/low/drivel )
         );
    oa21_1 \I1/low/U1669/U1  ( .x(\I1/low/U1669/n2 ), .a(\I1/low/U1669/n2 ), 
        .b(\I1/low/U1669/nr ), .c(\I1/low/U1669/nd ) );
    inv_2 \I1/low/U1669/U3  ( .x(net17), .a(\I1/low/U1669/n2 ) );
    buf_2 \I1/high/U1653  ( .x(\I1/high/latch ), .a(\I1/net33 ) );
    nor2_1 \I1/high/U264/U5  ( .x(\I1/high/nlocalcd ), .a(reset), .b(
        \I1/high/localcd ) );
    nor2_1 \I1/high/U1659_0_/U5  ( .x(\I1/high/ncd[0] ), .a(ol[24]), .b(oh[24]
        ) );
    nor2_1 \I1/high/U1659_1_/U5  ( .x(\I1/high/ncd[1] ), .a(ol[25]), .b(oh[25]
        ) );
    nor2_1 \I1/high/U1659_2_/U5  ( .x(\I1/high/ncd[2] ), .a(ol[26]), .b(oh[26]
        ) );
    nor2_1 \I1/high/U1659_3_/U5  ( .x(\I1/high/ncd[3] ), .a(ol[27]), .b(oh[27]
        ) );
    nor2_1 \I1/high/U1659_4_/U5  ( .x(\I1/high/ncd[4] ), .a(ol[28]), .b(oh[28]
        ) );
    nor2_1 \I1/high/U1659_5_/U5  ( .x(\I1/high/ncd[5] ), .a(ol[29]), .b(oh[29]
        ) );
    nor2_1 \I1/high/U1659_6_/U5  ( .x(\I1/high/ncd[6] ), .a(ol[30]), .b(oh[30]
        ) );
    nor2_1 \I1/high/U1659_7_/U5  ( .x(\I1/high/ncd[7] ), .a(ol[31]), .b(oh[31]
        ) );
    nor2_1 \I1/high/U3/U5  ( .x(\I1/high/ctrlack_internal ), .a(\I1/high/acb ), 
        .b(\I1/high/ba ) );
    ao23_1 \I1/high/U1658_0_/U21/U1/U1  ( .x(ol[24]), .a(n5), .b(ol[24]), .c(
        n6), .d(pull_l[0]), .e(n1) );
    ao23_1 \I1/high/U1658_1_/U21/U1/U1  ( .x(ol[25]), .a(n5), .b(ol[25]), .c(
        n6), .d(pull_l[1]), .e(n1) );
    ao23_1 \I1/high/U1658_2_/U21/U1/U1  ( .x(ol[26]), .a(n5), .b(ol[26]), .c(
        n6), .d(pull_l[2]), .e(n1) );
    ao23_1 \I1/high/U1658_3_/U21/U1/U1  ( .x(ol[27]), .a(n5), .b(ol[27]), .c(
        n5), .d(pull_l[3]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1658_4_/U21/U1/U1  ( .x(ol[28]), .a(n5), .b(ol[28]), .c(
        n6), .d(pull_l[4]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1658_5_/U21/U1/U1  ( .x(ol[29]), .a(n5), .b(ol[29]), .c(
        n6), .d(pull_l[5]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1658_6_/U21/U1/U1  ( .x(ol[30]), .a(n5), .b(ol[30]), .c(
        n5), .d(pull_l[6]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1658_7_/U21/U1/U1  ( .x(ol[31]), .a(n5), .b(ol[31]), .c(
        n5), .d(pull_l[7]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_0_/U21/U1/U1  ( .x(oh[24]), .a(n2), .b(oh[24]), .c(
        n3), .d(pull_h[0]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_1_/U21/U1/U1  ( .x(oh[25]), .a(n2), .b(oh[25]), .c(
        n2), .d(pull_h[1]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_2_/U21/U1/U1  ( .x(oh[26]), .a(n2), .b(oh[26]), .c(
        n3), .d(pull_h[2]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_3_/U21/U1/U1  ( .x(oh[27]), .a(n2), .b(oh[27]), .c(
        n2), .d(pull_h[3]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_4_/U21/U1/U1  ( .x(oh[28]), .a(n2), .b(oh[28]), .c(
        n3), .d(pull_h[4]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_5_/U21/U1/U1  ( .x(oh[29]), .a(n2), .b(oh[29]), .c(
        n2), .d(pull_h[5]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_6_/U21/U1/U1  ( .x(oh[30]), .a(n2), .b(oh[30]), .c(
        n3), .d(pull_h[6]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_7_/U21/U1/U1  ( .x(oh[31]), .a(n2), .b(oh[31]), .c(
        n3), .d(pull_h[7]), .e(\I1/high/latch ) );
    aoai211_1 \I1/high/U4/U28/U1/U1  ( .x(\I1/high/U4/U28/U1/clr ), .a(ctrlreq
        ), .b(\I1/high/acb ), .c(\I1/high/nlocalcd ), .d(\I1/net33 ) );
    nand3_1 \I1/high/U4/U28/U1/U2  ( .x(\I1/high/U4/U28/U1/set ), .a(
        \I1/high/nlocalcd ), .b(ctrlreq), .c(\I1/high/acb ) );
    nand2_2 \I1/high/U4/U28/U1/U3  ( .x(\I1/net33 ), .a(
        \I1/high/U4/U28/U1/clr ), .b(\I1/high/U4/U28/U1/set ) );
    oai21_1 \I1/high/U1/U30/U1/U1  ( .x(\I1/high/acb ), .a(\I1/high/U1/Z ), 
        .b(\I1/high/ba ), .c(ctrlreq) );
    inv_1 \I1/high/U1/U30/U1/U2  ( .x(\I1/high/U1/Z ), .a(\I1/high/acb ) );
    ao222_1 \I1/high/U5/U18/U1/U1  ( .x(\I1/high/ba ), .a(\I1/high/latch ), 
        .b(pullcd), .c(\I1/high/latch ), .d(\I1/high/ba ), .e(pullcd), .f(
        \I1/high/ba ) );
    aoi222_1 \I1/high/U1664/U28/U30/U1  ( .x(\I1/high/U1664/x[3] ), .a(
        \I1/high/ncd[7] ), .b(\I1/high/ncd[6] ), .c(\I1/high/ncd[7] ), .d(
        \I1/high/U1664/U28/Z ), .e(\I1/high/ncd[6] ), .f(\I1/high/U1664/U28/Z 
        ) );
    inv_1 \I1/high/U1664/U28/U30/Uinv  ( .x(\I1/high/U1664/U28/Z ), .a(
        \I1/high/U1664/x[3] ) );
    aoi222_1 \I1/high/U1664/U32/U30/U1  ( .x(\I1/high/U1664/x[0] ), .a(
        \I1/high/ncd[1] ), .b(\I1/high/ncd[0] ), .c(\I1/high/ncd[1] ), .d(
        \I1/high/U1664/U32/Z ), .e(\I1/high/ncd[0] ), .f(\I1/high/U1664/U32/Z 
        ) );
    inv_1 \I1/high/U1664/U32/U30/Uinv  ( .x(\I1/high/U1664/U32/Z ), .a(
        \I1/high/U1664/x[0] ) );
    aoi222_1 \I1/high/U1664/U29/U30/U1  ( .x(\I1/high/U1664/x[2] ), .a(
        \I1/high/ncd[5] ), .b(\I1/high/ncd[4] ), .c(\I1/high/ncd[5] ), .d(
        \I1/high/U1664/U29/Z ), .e(\I1/high/ncd[4] ), .f(\I1/high/U1664/U29/Z 
        ) );
    inv_1 \I1/high/U1664/U29/U30/Uinv  ( .x(\I1/high/U1664/U29/Z ), .a(
        \I1/high/U1664/x[2] ) );
    aoi222_1 \I1/high/U1664/U33/U30/U1  ( .x(\I1/high/U1664/y[0] ), .a(
        \I1/high/U1664/x[1] ), .b(\I1/high/U1664/x[0] ), .c(
        \I1/high/U1664/x[1] ), .d(\I1/high/U1664/U33/Z ), .e(
        \I1/high/U1664/x[0] ), .f(\I1/high/U1664/U33/Z ) );
    inv_1 \I1/high/U1664/U33/U30/Uinv  ( .x(\I1/high/U1664/U33/Z ), .a(
        \I1/high/U1664/y[0] ) );
    aoi222_1 \I1/high/U1664/U30/U30/U1  ( .x(\I1/high/U1664/y[1] ), .a(
        \I1/high/U1664/x[3] ), .b(\I1/high/U1664/x[2] ), .c(
        \I1/high/U1664/x[3] ), .d(\I1/high/U1664/U30/Z ), .e(
        \I1/high/U1664/x[2] ), .f(\I1/high/U1664/U30/Z ) );
    inv_1 \I1/high/U1664/U30/U30/Uinv  ( .x(\I1/high/U1664/U30/Z ), .a(
        \I1/high/U1664/y[1] ) );
    aoi222_1 \I1/high/U1664/U31/U30/U1  ( .x(\I1/high/U1664/x[1] ), .a(
        \I1/high/ncd[3] ), .b(\I1/high/ncd[2] ), .c(\I1/high/ncd[3] ), .d(
        \I1/high/U1664/U31/Z ), .e(\I1/high/ncd[2] ), .f(\I1/high/U1664/U31/Z 
        ) );
    inv_1 \I1/high/U1664/U31/U30/Uinv  ( .x(\I1/high/U1664/U31/Z ), .a(
        \I1/high/U1664/x[1] ) );
    aoi222_1 \I1/high/U1664/U37/U30/U1  ( .x(\I1/high/localcd ), .a(
        \I1/high/U1664/y[0] ), .b(\I1/high/U1664/y[1] ), .c(
        \I1/high/U1664/y[0] ), .d(\I1/high/U1664/U37/Z ), .e(
        \I1/high/U1664/y[1] ), .f(\I1/high/U1664/U37/Z ) );
    inv_1 \I1/high/U1664/U37/U30/Uinv  ( .x(\I1/high/U1664/U37/Z ), .a(
        \I1/high/localcd ) );
    nor3_1 \I1/high/U1669/Unr  ( .x(\I1/high/U1669/nr ), .a(
        \I1/high/ctrlack_internal ), .b(n6), .c(n3) );
    nand3_1 \I1/high/U1669/Und  ( .x(\I1/high/U1669/nd ), .a(
        \I1/high/ctrlack_internal ), .b(n6), .c(n3) );
    oa21_1 \I1/high/U1669/U1  ( .x(\I1/high/U1669/n2 ), .a(\I1/high/U1669/n2 ), 
        .b(\I1/high/U1669/nr ), .c(\I1/high/U1669/nd ) );
    inv_2 \I1/high/U1669/U3  ( .x(\I1/net20 ), .a(\I1/high/U1669/n2 ) );
    buf_1 U1 ( .x(n1), .a(\I1/high/latch ) );
    inv_2 U2 ( .x(n2), .a(n4) );
    inv_1 U3 ( .x(n3), .a(n4) );
    inv_0 U4 ( .x(n4), .a(ctrlreq) );
    inv_2 U5 ( .x(n5), .a(n4) );
    inv_1 U6 ( .x(n6), .a(n4) );
    buf_1 U7 ( .x(n7), .a(\I1/low/latch ) );
    buf_2 U8 ( .x(n8), .a(\I1/net20 ) );
    buf_1 U9 ( .x(n9), .a(\I0/high/latch ) );
    buf_2 U10 ( .x(n10), .a(net17) );
    buf_1 U11 ( .x(n11), .a(\I0/low/latch ) );
    buf_2 U12 ( .x(n12), .a(\I0/net20 ) );
endmodule


module chain_irdemux_32new_0 ( ctrlack, oh, ol, pullreq, pull_h, pull_l, 
    pullcd, reset, ctrlreq );
output [31:0] oh;
output [31:0] ol;
input  [7:0] pull_h;
input  [7:0] pull_l;
input  pullcd, reset, ctrlreq;
output ctrlack, pullreq;
    wire net30, net31, \I0/net32 , \I0/net33 , \I0/low/latch , 
        \I0/low/nlocalcd , \I0/low/localcd , \I0/low/ncd[0] , \I0/low/ncd[1] , 
        \I0/low/ncd[2] , \I0/low/ncd[3] , \I0/low/ncd[4] , \I0/low/ncd[5] , 
        \I0/low/ncd[6] , \I0/low/ncd[7] , \I0/low/ctrlack_internal , 
        \I0/low/acb , \I0/low/ba , \I0/low/driveh , \I0/net20 , 
        \I0/low/drivel , n1, n2, \I0/low/U4/U28/U1/clr , 
        \I0/low/U4/U28/U1/set , \I0/low/U1/Z , \I0/low/U1664/x[3] , 
        \I0/low/U1664/U28/Z , \I0/low/U1664/x[0] , \I0/low/U1664/U32/Z , 
        \I0/low/U1664/x[2] , \I0/low/U1664/U29/Z , \I0/low/U1664/y[0] , 
        \I0/low/U1664/x[1] , \I0/low/U1664/U33/Z , \I0/low/U1664/y[1] , 
        \I0/low/U1664/U30/Z , \I0/low/U1664/U31/Z , \I0/low/U1664/U37/Z , 
        \I0/low/U1669/nr , \I0/low/U1669/nd , \I0/low/U1669/n2 , 
        \I0/high/latch , \I0/high/nlocalcd , \I0/high/localcd , 
        \I0/high/ncd[0] , \I0/high/ncd[1] , \I0/high/ncd[2] , \I0/high/ncd[3] , 
        \I0/high/ncd[4] , \I0/high/ncd[5] , \I0/high/ncd[6] , \I0/high/ncd[7] , 
        \I0/high/ctrlack_internal , \I0/high/acb , \I0/high/ba , 
        \I0/high/driveh , net17, \I0/high/drivel , n3, n4, 
        \I0/high/U4/U28/U1/clr , \I0/high/U4/U28/U1/set , \I0/high/U1/Z , 
        \I0/high/U1664/x[3] , \I0/high/U1664/U28/Z , \I0/high/U1664/x[0] , 
        \I0/high/U1664/U32/Z , \I0/high/U1664/x[2] , \I0/high/U1664/U29/Z , 
        \I0/high/U1664/y[0] , \I0/high/U1664/x[1] , \I0/high/U1664/U33/Z , 
        \I0/high/U1664/y[1] , \I0/high/U1664/U30/Z , \I0/high/U1664/U31/Z , 
        \I0/high/U1664/U37/Z , \I0/high/U1669/nr , \I0/high/U1669/nd , 
        \I0/high/U1669/n2 , \I1/net32 , \I1/net33 , \I1/low/latch , 
        \I1/low/nlocalcd , \I1/low/localcd , \I1/low/ncd[0] , \I1/low/ncd[1] , 
        \I1/low/ncd[2] , \I1/low/ncd[3] , \I1/low/ncd[4] , \I1/low/ncd[5] , 
        \I1/low/ncd[6] , \I1/low/ncd[7] , \I1/low/ctrlack_internal , 
        \I1/low/acb , \I1/low/ba , \I1/low/driveh , \I1/net20 , 
        \I1/low/drivel , n5, n6, \I1/low/U4/U28/U1/clr , 
        \I1/low/U4/U28/U1/set , \I1/low/U1/Z , \I1/low/U1664/x[3] , 
        \I1/low/U1664/U28/Z , \I1/low/U1664/x[0] , \I1/low/U1664/U32/Z , 
        \I1/low/U1664/x[2] , \I1/low/U1664/U29/Z , \I1/low/U1664/y[0] , 
        \I1/low/U1664/x[1] , \I1/low/U1664/U33/Z , \I1/low/U1664/y[1] , 
        \I1/low/U1664/U30/Z , \I1/low/U1664/U31/Z , \I1/low/U1664/U37/Z , 
        \I1/low/U1669/nr , \I1/low/U1669/nd , \I1/low/U1669/n2 , 
        \I1/high/latch , \I1/high/nlocalcd , \I1/high/localcd , 
        \I1/high/ncd[0] , \I1/high/ncd[1] , \I1/high/ncd[2] , \I1/high/ncd[3] , 
        \I1/high/ncd[4] , \I1/high/ncd[5] , \I1/high/ncd[6] , \I1/high/ncd[7] , 
        \I1/high/ctrlack_internal , \I1/high/acb , \I1/high/ba , 
        \I1/high/driveh , \I1/high/drivel , n7, n8, \I1/high/U4/U28/U1/clr , 
        \I1/high/U4/U28/U1/set , \I1/high/U1/Z , \I1/high/U1664/x[3] , 
        \I1/high/U1664/U28/Z , \I1/high/U1664/x[0] , \I1/high/U1664/U32/Z , 
        \I1/high/U1664/x[2] , \I1/high/U1664/U29/Z , \I1/high/U1664/y[0] , 
        \I1/high/U1664/x[1] , \I1/high/U1664/U33/Z , \I1/high/U1664/y[1] , 
        \I1/high/U1664/U30/Z , \I1/high/U1664/U31/Z , \I1/high/U1664/U37/Z , 
        \I1/high/U1669/nr , \I1/high/U1669/nd , \I1/high/U1669/n2 ;
    nand2_1 \U3/U5  ( .x(pullreq), .a(net30), .b(net31) );
    nor2_1 \I0/U3/U5  ( .x(net30), .a(\I0/net32 ), .b(\I0/net33 ) );
    buf_2 \I0/low/U1653  ( .x(\I0/low/latch ), .a(\I0/net32 ) );
    nor2_1 \I0/low/U264/U5  ( .x(\I0/low/nlocalcd ), .a(reset), .b(
        \I0/low/localcd ) );
    nor2_1 \I0/low/U1659_0_/U5  ( .x(\I0/low/ncd[0] ), .a(ol[0]), .b(oh[0]) );
    nor2_1 \I0/low/U1659_1_/U5  ( .x(\I0/low/ncd[1] ), .a(ol[1]), .b(oh[1]) );
    nor2_1 \I0/low/U1659_2_/U5  ( .x(\I0/low/ncd[2] ), .a(ol[2]), .b(oh[2]) );
    nor2_1 \I0/low/U1659_3_/U5  ( .x(\I0/low/ncd[3] ), .a(ol[3]), .b(oh[3]) );
    nor2_1 \I0/low/U1659_4_/U5  ( .x(\I0/low/ncd[4] ), .a(ol[4]), .b(oh[4]) );
    nor2_1 \I0/low/U1659_5_/U5  ( .x(\I0/low/ncd[5] ), .a(ol[5]), .b(oh[5]) );
    nor2_1 \I0/low/U1659_6_/U5  ( .x(\I0/low/ncd[6] ), .a(ol[6]), .b(oh[6]) );
    nor2_1 \I0/low/U1659_7_/U5  ( .x(\I0/low/ncd[7] ), .a(ol[7]), .b(oh[7]) );
    nor2_1 \I0/low/U3/U5  ( .x(\I0/low/ctrlack_internal ), .a(\I0/low/acb ), 
        .b(\I0/low/ba ) );
    buf_2 \I0/low/U1665/U7  ( .x(\I0/low/driveh ), .a(\I0/net20 ) );
    buf_2 \I0/low/U1666/U7  ( .x(\I0/low/drivel ), .a(\I0/net20 ) );
    ao23_1 \I0/low/U1658_0_/U21/U1/U1  ( .x(ol[0]), .a(\I0/low/driveh ), .b(ol
        [0]), .c(n1), .d(pull_l[0]), .e(n2) );
    ao23_1 \I0/low/U1658_1_/U21/U1/U1  ( .x(ol[1]), .a(\I0/low/drivel ), .b(ol
        [1]), .c(\I0/low/driveh ), .d(pull_l[1]), .e(n2) );
    ao23_1 \I0/low/U1658_2_/U21/U1/U1  ( .x(ol[2]), .a(\I0/low/drivel ), .b(ol
        [2]), .c(\I0/low/driveh ), .d(pull_l[2]), .e(n2) );
    ao23_1 \I0/low/U1658_3_/U21/U1/U1  ( .x(ol[3]), .a(\I0/low/driveh ), .b(ol
        [3]), .c(\I0/low/drivel ), .d(pull_l[3]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_4_/U21/U1/U1  ( .x(ol[4]), .a(n1), .b(ol[4]), .c(
        \I0/low/drivel ), .d(pull_l[4]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_5_/U21/U1/U1  ( .x(ol[5]), .a(\I0/low/driveh ), .b(ol
        [5]), .c(n1), .d(pull_l[5]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_6_/U21/U1/U1  ( .x(ol[6]), .a(\I0/low/drivel ), .b(ol
        [6]), .c(\I0/low/driveh ), .d(pull_l[6]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_7_/U21/U1/U1  ( .x(ol[7]), .a(n1), .b(ol[7]), .c(n1), 
        .d(pull_l[7]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_0_/U21/U1/U1  ( .x(oh[0]), .a(\I0/low/driveh ), .b(oh
        [0]), .c(n1), .d(pull_h[0]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_1_/U21/U1/U1  ( .x(oh[1]), .a(n1), .b(oh[1]), .c(
        \I0/low/drivel ), .d(pull_h[1]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_2_/U21/U1/U1  ( .x(oh[2]), .a(\I0/low/drivel ), .b(oh
        [2]), .c(\I0/low/drivel ), .d(pull_h[2]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_3_/U21/U1/U1  ( .x(oh[3]), .a(n1), .b(oh[3]), .c(
        \I0/low/driveh ), .d(pull_h[3]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_4_/U21/U1/U1  ( .x(oh[4]), .a(n1), .b(oh[4]), .c(n1), 
        .d(pull_h[4]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_5_/U21/U1/U1  ( .x(oh[5]), .a(\I0/low/drivel ), .b(oh
        [5]), .c(n1), .d(pull_h[5]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_6_/U21/U1/U1  ( .x(oh[6]), .a(\I0/low/drivel ), .b(oh
        [6]), .c(\I0/low/driveh ), .d(pull_h[6]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_7_/U21/U1/U1  ( .x(oh[7]), .a(\I0/low/driveh ), .b(oh
        [7]), .c(\I0/low/drivel ), .d(pull_h[7]), .e(\I0/low/latch ) );
    aoai211_1 \I0/low/U4/U28/U1/U1  ( .x(\I0/low/U4/U28/U1/clr ), .a(
        \I0/net20 ), .b(\I0/low/acb ), .c(\I0/low/nlocalcd ), .d(\I0/net32 )
         );
    nand3_1 \I0/low/U4/U28/U1/U2  ( .x(\I0/low/U4/U28/U1/set ), .a(
        \I0/low/nlocalcd ), .b(\I0/net20 ), .c(\I0/low/acb ) );
    nand2_2 \I0/low/U4/U28/U1/U3  ( .x(\I0/net32 ), .a(\I0/low/U4/U28/U1/clr ), 
        .b(\I0/low/U4/U28/U1/set ) );
    oai21_1 \I0/low/U1/U30/U1/U1  ( .x(\I0/low/acb ), .a(\I0/low/U1/Z ), .b(
        \I0/low/ba ), .c(\I0/net20 ) );
    inv_1 \I0/low/U1/U30/U1/U2  ( .x(\I0/low/U1/Z ), .a(\I0/low/acb ) );
    ao222_1 \I0/low/U5/U18/U1/U1  ( .x(\I0/low/ba ), .a(\I0/low/latch ), .b(
        pullcd), .c(\I0/low/latch ), .d(\I0/low/ba ), .e(pullcd), .f(
        \I0/low/ba ) );
    aoi222_1 \I0/low/U1664/U28/U30/U1  ( .x(\I0/low/U1664/x[3] ), .a(
        \I0/low/ncd[7] ), .b(\I0/low/ncd[6] ), .c(\I0/low/ncd[7] ), .d(
        \I0/low/U1664/U28/Z ), .e(\I0/low/ncd[6] ), .f(\I0/low/U1664/U28/Z )
         );
    inv_1 \I0/low/U1664/U28/U30/Uinv  ( .x(\I0/low/U1664/U28/Z ), .a(
        \I0/low/U1664/x[3] ) );
    aoi222_1 \I0/low/U1664/U32/U30/U1  ( .x(\I0/low/U1664/x[0] ), .a(
        \I0/low/ncd[1] ), .b(\I0/low/ncd[0] ), .c(\I0/low/ncd[1] ), .d(
        \I0/low/U1664/U32/Z ), .e(\I0/low/ncd[0] ), .f(\I0/low/U1664/U32/Z )
         );
    inv_1 \I0/low/U1664/U32/U30/Uinv  ( .x(\I0/low/U1664/U32/Z ), .a(
        \I0/low/U1664/x[0] ) );
    aoi222_1 \I0/low/U1664/U29/U30/U1  ( .x(\I0/low/U1664/x[2] ), .a(
        \I0/low/ncd[5] ), .b(\I0/low/ncd[4] ), .c(\I0/low/ncd[5] ), .d(
        \I0/low/U1664/U29/Z ), .e(\I0/low/ncd[4] ), .f(\I0/low/U1664/U29/Z )
         );
    inv_1 \I0/low/U1664/U29/U30/Uinv  ( .x(\I0/low/U1664/U29/Z ), .a(
        \I0/low/U1664/x[2] ) );
    aoi222_1 \I0/low/U1664/U33/U30/U1  ( .x(\I0/low/U1664/y[0] ), .a(
        \I0/low/U1664/x[1] ), .b(\I0/low/U1664/x[0] ), .c(\I0/low/U1664/x[1] ), 
        .d(\I0/low/U1664/U33/Z ), .e(\I0/low/U1664/x[0] ), .f(
        \I0/low/U1664/U33/Z ) );
    inv_1 \I0/low/U1664/U33/U30/Uinv  ( .x(\I0/low/U1664/U33/Z ), .a(
        \I0/low/U1664/y[0] ) );
    aoi222_1 \I0/low/U1664/U30/U30/U1  ( .x(\I0/low/U1664/y[1] ), .a(
        \I0/low/U1664/x[3] ), .b(\I0/low/U1664/x[2] ), .c(\I0/low/U1664/x[3] ), 
        .d(\I0/low/U1664/U30/Z ), .e(\I0/low/U1664/x[2] ), .f(
        \I0/low/U1664/U30/Z ) );
    inv_1 \I0/low/U1664/U30/U30/Uinv  ( .x(\I0/low/U1664/U30/Z ), .a(
        \I0/low/U1664/y[1] ) );
    aoi222_1 \I0/low/U1664/U31/U30/U1  ( .x(\I0/low/U1664/x[1] ), .a(
        \I0/low/ncd[3] ), .b(\I0/low/ncd[2] ), .c(\I0/low/ncd[3] ), .d(
        \I0/low/U1664/U31/Z ), .e(\I0/low/ncd[2] ), .f(\I0/low/U1664/U31/Z )
         );
    inv_1 \I0/low/U1664/U31/U30/Uinv  ( .x(\I0/low/U1664/U31/Z ), .a(
        \I0/low/U1664/x[1] ) );
    aoi222_1 \I0/low/U1664/U37/U30/U1  ( .x(\I0/low/localcd ), .a(
        \I0/low/U1664/y[0] ), .b(\I0/low/U1664/y[1] ), .c(\I0/low/U1664/y[0] ), 
        .d(\I0/low/U1664/U37/Z ), .e(\I0/low/U1664/y[1] ), .f(
        \I0/low/U1664/U37/Z ) );
    inv_1 \I0/low/U1664/U37/U30/Uinv  ( .x(\I0/low/U1664/U37/Z ), .a(
        \I0/low/localcd ) );
    nor3_1 \I0/low/U1669/Unr  ( .x(\I0/low/U1669/nr ), .a(
        \I0/low/ctrlack_internal ), .b(n1), .c(\I0/low/driveh ) );
    nand3_1 \I0/low/U1669/Und  ( .x(\I0/low/U1669/nd ), .a(
        \I0/low/ctrlack_internal ), .b(\I0/low/drivel ), .c(\I0/low/driveh )
         );
    oa21_1 \I0/low/U1669/U1  ( .x(\I0/low/U1669/n2 ), .a(\I0/low/U1669/n2 ), 
        .b(\I0/low/U1669/nr ), .c(\I0/low/U1669/nd ) );
    inv_2 \I0/low/U1669/U3  ( .x(ctrlack), .a(\I0/low/U1669/n2 ) );
    buf_2 \I0/high/U1653  ( .x(\I0/high/latch ), .a(\I0/net33 ) );
    nor2_1 \I0/high/U264/U5  ( .x(\I0/high/nlocalcd ), .a(reset), .b(
        \I0/high/localcd ) );
    nor2_1 \I0/high/U1659_0_/U5  ( .x(\I0/high/ncd[0] ), .a(ol[8]), .b(oh[8])
         );
    nor2_1 \I0/high/U1659_1_/U5  ( .x(\I0/high/ncd[1] ), .a(ol[9]), .b(oh[9])
         );
    nor2_1 \I0/high/U1659_2_/U5  ( .x(\I0/high/ncd[2] ), .a(ol[10]), .b(oh[10]
        ) );
    nor2_1 \I0/high/U1659_3_/U5  ( .x(\I0/high/ncd[3] ), .a(ol[11]), .b(oh[11]
        ) );
    nor2_1 \I0/high/U1659_4_/U5  ( .x(\I0/high/ncd[4] ), .a(ol[12]), .b(oh[12]
        ) );
    nor2_1 \I0/high/U1659_5_/U5  ( .x(\I0/high/ncd[5] ), .a(ol[13]), .b(oh[13]
        ) );
    nor2_1 \I0/high/U1659_6_/U5  ( .x(\I0/high/ncd[6] ), .a(ol[14]), .b(oh[14]
        ) );
    nor2_1 \I0/high/U1659_7_/U5  ( .x(\I0/high/ncd[7] ), .a(ol[15]), .b(oh[15]
        ) );
    nor2_1 \I0/high/U3/U5  ( .x(\I0/high/ctrlack_internal ), .a(\I0/high/acb ), 
        .b(\I0/high/ba ) );
    buf_2 \I0/high/U1665/U7  ( .x(\I0/high/driveh ), .a(net17) );
    buf_2 \I0/high/U1666/U7  ( .x(\I0/high/drivel ), .a(net17) );
    ao23_1 \I0/high/U1658_0_/U21/U1/U1  ( .x(ol[8]), .a(\I0/high/driveh ), .b(
        ol[8]), .c(n3), .d(pull_l[0]), .e(n4) );
    ao23_1 \I0/high/U1658_1_/U21/U1/U1  ( .x(ol[9]), .a(\I0/high/drivel ), .b(
        ol[9]), .c(\I0/high/driveh ), .d(pull_l[1]), .e(n4) );
    ao23_1 \I0/high/U1658_2_/U21/U1/U1  ( .x(ol[10]), .a(\I0/high/drivel ), 
        .b(ol[10]), .c(\I0/high/driveh ), .d(pull_l[2]), .e(n4) );
    ao23_1 \I0/high/U1658_3_/U21/U1/U1  ( .x(ol[11]), .a(\I0/high/driveh ), 
        .b(ol[11]), .c(\I0/high/drivel ), .d(pull_l[3]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1658_4_/U21/U1/U1  ( .x(ol[12]), .a(n3), .b(ol[12]), .c(
        \I0/high/drivel ), .d(pull_l[4]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1658_5_/U21/U1/U1  ( .x(ol[13]), .a(\I0/high/driveh ), 
        .b(ol[13]), .c(n3), .d(pull_l[5]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1658_6_/U21/U1/U1  ( .x(ol[14]), .a(\I0/high/drivel ), 
        .b(ol[14]), .c(\I0/high/driveh ), .d(pull_l[6]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1658_7_/U21/U1/U1  ( .x(ol[15]), .a(n3), .b(ol[15]), .c(
        n3), .d(pull_l[7]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_0_/U21/U1/U1  ( .x(oh[8]), .a(\I0/high/driveh ), .b(
        oh[8]), .c(n3), .d(pull_h[0]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_1_/U21/U1/U1  ( .x(oh[9]), .a(n3), .b(oh[9]), .c(
        \I0/high/drivel ), .d(pull_h[1]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_2_/U21/U1/U1  ( .x(oh[10]), .a(\I0/high/drivel ), 
        .b(oh[10]), .c(\I0/high/drivel ), .d(pull_h[2]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1651_3_/U21/U1/U1  ( .x(oh[11]), .a(n3), .b(oh[11]), .c(
        \I0/high/driveh ), .d(pull_h[3]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_4_/U21/U1/U1  ( .x(oh[12]), .a(n3), .b(oh[12]), .c(
        n3), .d(pull_h[4]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_5_/U21/U1/U1  ( .x(oh[13]), .a(\I0/high/drivel ), 
        .b(oh[13]), .c(n3), .d(pull_h[5]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_6_/U21/U1/U1  ( .x(oh[14]), .a(\I0/high/drivel ), 
        .b(oh[14]), .c(\I0/high/driveh ), .d(pull_h[6]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1651_7_/U21/U1/U1  ( .x(oh[15]), .a(\I0/high/driveh ), 
        .b(oh[15]), .c(\I0/high/drivel ), .d(pull_h[7]), .e(\I0/high/latch )
         );
    aoai211_1 \I0/high/U4/U28/U1/U1  ( .x(\I0/high/U4/U28/U1/clr ), .a(net17), 
        .b(\I0/high/acb ), .c(\I0/high/nlocalcd ), .d(\I0/net33 ) );
    nand3_1 \I0/high/U4/U28/U1/U2  ( .x(\I0/high/U4/U28/U1/set ), .a(
        \I0/high/nlocalcd ), .b(net17), .c(\I0/high/acb ) );
    nand2_2 \I0/high/U4/U28/U1/U3  ( .x(\I0/net33 ), .a(
        \I0/high/U4/U28/U1/clr ), .b(\I0/high/U4/U28/U1/set ) );
    oai21_1 \I0/high/U1/U30/U1/U1  ( .x(\I0/high/acb ), .a(\I0/high/U1/Z ), 
        .b(\I0/high/ba ), .c(net17) );
    inv_1 \I0/high/U1/U30/U1/U2  ( .x(\I0/high/U1/Z ), .a(\I0/high/acb ) );
    ao222_1 \I0/high/U5/U18/U1/U1  ( .x(\I0/high/ba ), .a(\I0/high/latch ), 
        .b(pullcd), .c(\I0/high/latch ), .d(\I0/high/ba ), .e(pullcd), .f(
        \I0/high/ba ) );
    aoi222_1 \I0/high/U1664/U28/U30/U1  ( .x(\I0/high/U1664/x[3] ), .a(
        \I0/high/ncd[7] ), .b(\I0/high/ncd[6] ), .c(\I0/high/ncd[7] ), .d(
        \I0/high/U1664/U28/Z ), .e(\I0/high/ncd[6] ), .f(\I0/high/U1664/U28/Z 
        ) );
    inv_1 \I0/high/U1664/U28/U30/Uinv  ( .x(\I0/high/U1664/U28/Z ), .a(
        \I0/high/U1664/x[3] ) );
    aoi222_1 \I0/high/U1664/U32/U30/U1  ( .x(\I0/high/U1664/x[0] ), .a(
        \I0/high/ncd[1] ), .b(\I0/high/ncd[0] ), .c(\I0/high/ncd[1] ), .d(
        \I0/high/U1664/U32/Z ), .e(\I0/high/ncd[0] ), .f(\I0/high/U1664/U32/Z 
        ) );
    inv_1 \I0/high/U1664/U32/U30/Uinv  ( .x(\I0/high/U1664/U32/Z ), .a(
        \I0/high/U1664/x[0] ) );
    aoi222_1 \I0/high/U1664/U29/U30/U1  ( .x(\I0/high/U1664/x[2] ), .a(
        \I0/high/ncd[5] ), .b(\I0/high/ncd[4] ), .c(\I0/high/ncd[5] ), .d(
        \I0/high/U1664/U29/Z ), .e(\I0/high/ncd[4] ), .f(\I0/high/U1664/U29/Z 
        ) );
    inv_1 \I0/high/U1664/U29/U30/Uinv  ( .x(\I0/high/U1664/U29/Z ), .a(
        \I0/high/U1664/x[2] ) );
    aoi222_1 \I0/high/U1664/U33/U30/U1  ( .x(\I0/high/U1664/y[0] ), .a(
        \I0/high/U1664/x[1] ), .b(\I0/high/U1664/x[0] ), .c(
        \I0/high/U1664/x[1] ), .d(\I0/high/U1664/U33/Z ), .e(
        \I0/high/U1664/x[0] ), .f(\I0/high/U1664/U33/Z ) );
    inv_1 \I0/high/U1664/U33/U30/Uinv  ( .x(\I0/high/U1664/U33/Z ), .a(
        \I0/high/U1664/y[0] ) );
    aoi222_1 \I0/high/U1664/U30/U30/U1  ( .x(\I0/high/U1664/y[1] ), .a(
        \I0/high/U1664/x[3] ), .b(\I0/high/U1664/x[2] ), .c(
        \I0/high/U1664/x[3] ), .d(\I0/high/U1664/U30/Z ), .e(
        \I0/high/U1664/x[2] ), .f(\I0/high/U1664/U30/Z ) );
    inv_1 \I0/high/U1664/U30/U30/Uinv  ( .x(\I0/high/U1664/U30/Z ), .a(
        \I0/high/U1664/y[1] ) );
    aoi222_1 \I0/high/U1664/U31/U30/U1  ( .x(\I0/high/U1664/x[1] ), .a(
        \I0/high/ncd[3] ), .b(\I0/high/ncd[2] ), .c(\I0/high/ncd[3] ), .d(
        \I0/high/U1664/U31/Z ), .e(\I0/high/ncd[2] ), .f(\I0/high/U1664/U31/Z 
        ) );
    inv_1 \I0/high/U1664/U31/U30/Uinv  ( .x(\I0/high/U1664/U31/Z ), .a(
        \I0/high/U1664/x[1] ) );
    aoi222_1 \I0/high/U1664/U37/U30/U1  ( .x(\I0/high/localcd ), .a(
        \I0/high/U1664/y[0] ), .b(\I0/high/U1664/y[1] ), .c(
        \I0/high/U1664/y[0] ), .d(\I0/high/U1664/U37/Z ), .e(
        \I0/high/U1664/y[1] ), .f(\I0/high/U1664/U37/Z ) );
    inv_1 \I0/high/U1664/U37/U30/Uinv  ( .x(\I0/high/U1664/U37/Z ), .a(
        \I0/high/localcd ) );
    nor3_1 \I0/high/U1669/Unr  ( .x(\I0/high/U1669/nr ), .a(
        \I0/high/ctrlack_internal ), .b(n3), .c(\I0/high/driveh ) );
    nand3_1 \I0/high/U1669/Und  ( .x(\I0/high/U1669/nd ), .a(
        \I0/high/ctrlack_internal ), .b(\I0/high/drivel ), .c(\I0/high/driveh 
        ) );
    oa21_1 \I0/high/U1669/U1  ( .x(\I0/high/U1669/n2 ), .a(\I0/high/U1669/n2 ), 
        .b(\I0/high/U1669/nr ), .c(\I0/high/U1669/nd ) );
    inv_2 \I0/high/U1669/U3  ( .x(\I0/net20 ), .a(\I0/high/U1669/n2 ) );
    nor2_1 \I1/U3/U5  ( .x(net31), .a(\I1/net32 ), .b(\I1/net33 ) );
    buf_2 \I1/low/U1653  ( .x(\I1/low/latch ), .a(\I1/net32 ) );
    nor2_1 \I1/low/U264/U5  ( .x(\I1/low/nlocalcd ), .a(reset), .b(
        \I1/low/localcd ) );
    nor2_1 \I1/low/U1659_0_/U5  ( .x(\I1/low/ncd[0] ), .a(ol[16]), .b(oh[16])
         );
    nor2_1 \I1/low/U1659_1_/U5  ( .x(\I1/low/ncd[1] ), .a(ol[17]), .b(oh[17])
         );
    nor2_1 \I1/low/U1659_2_/U5  ( .x(\I1/low/ncd[2] ), .a(ol[18]), .b(oh[18])
         );
    nor2_1 \I1/low/U1659_3_/U5  ( .x(\I1/low/ncd[3] ), .a(ol[19]), .b(oh[19])
         );
    nor2_1 \I1/low/U1659_4_/U5  ( .x(\I1/low/ncd[4] ), .a(ol[20]), .b(oh[20])
         );
    nor2_1 \I1/low/U1659_5_/U5  ( .x(\I1/low/ncd[5] ), .a(ol[21]), .b(oh[21])
         );
    nor2_1 \I1/low/U1659_6_/U5  ( .x(\I1/low/ncd[6] ), .a(ol[22]), .b(oh[22])
         );
    nor2_1 \I1/low/U1659_7_/U5  ( .x(\I1/low/ncd[7] ), .a(ol[23]), .b(oh[23])
         );
    nor2_1 \I1/low/U3/U5  ( .x(\I1/low/ctrlack_internal ), .a(\I1/low/acb ), 
        .b(\I1/low/ba ) );
    buf_2 \I1/low/U1665/U7  ( .x(\I1/low/driveh ), .a(\I1/net20 ) );
    buf_2 \I1/low/U1666/U7  ( .x(\I1/low/drivel ), .a(\I1/net20 ) );
    ao23_1 \I1/low/U1658_0_/U21/U1/U1  ( .x(ol[16]), .a(\I1/low/driveh ), .b(
        ol[16]), .c(n5), .d(pull_l[0]), .e(n6) );
    ao23_1 \I1/low/U1658_1_/U21/U1/U1  ( .x(ol[17]), .a(\I1/low/drivel ), .b(
        ol[17]), .c(\I1/low/driveh ), .d(pull_l[1]), .e(n6) );
    ao23_1 \I1/low/U1658_2_/U21/U1/U1  ( .x(ol[18]), .a(\I1/low/drivel ), .b(
        ol[18]), .c(\I1/low/driveh ), .d(pull_l[2]), .e(n6) );
    ao23_1 \I1/low/U1658_3_/U21/U1/U1  ( .x(ol[19]), .a(\I1/low/driveh ), .b(
        ol[19]), .c(\I1/low/drivel ), .d(pull_l[3]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_4_/U21/U1/U1  ( .x(ol[20]), .a(n5), .b(ol[20]), .c(
        \I1/low/drivel ), .d(pull_l[4]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_5_/U21/U1/U1  ( .x(ol[21]), .a(\I1/low/driveh ), .b(
        ol[21]), .c(n5), .d(pull_l[5]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_6_/U21/U1/U1  ( .x(ol[22]), .a(\I1/low/drivel ), .b(
        ol[22]), .c(\I1/low/driveh ), .d(pull_l[6]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_7_/U21/U1/U1  ( .x(ol[23]), .a(n5), .b(ol[23]), .c(n5
        ), .d(pull_l[7]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_0_/U21/U1/U1  ( .x(oh[16]), .a(\I1/low/driveh ), .b(
        oh[16]), .c(n5), .d(pull_h[0]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_1_/U21/U1/U1  ( .x(oh[17]), .a(n5), .b(oh[17]), .c(
        \I1/low/drivel ), .d(pull_h[1]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_2_/U21/U1/U1  ( .x(oh[18]), .a(\I1/low/drivel ), .b(
        oh[18]), .c(\I1/low/drivel ), .d(pull_h[2]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_3_/U21/U1/U1  ( .x(oh[19]), .a(n5), .b(oh[19]), .c(
        \I1/low/driveh ), .d(pull_h[3]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_4_/U21/U1/U1  ( .x(oh[20]), .a(n5), .b(oh[20]), .c(n5
        ), .d(pull_h[4]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_5_/U21/U1/U1  ( .x(oh[21]), .a(\I1/low/drivel ), .b(
        oh[21]), .c(n5), .d(pull_h[5]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_6_/U21/U1/U1  ( .x(oh[22]), .a(\I1/low/drivel ), .b(
        oh[22]), .c(\I1/low/driveh ), .d(pull_h[6]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_7_/U21/U1/U1  ( .x(oh[23]), .a(\I1/low/driveh ), .b(
        oh[23]), .c(\I1/low/drivel ), .d(pull_h[7]), .e(\I1/low/latch ) );
    aoai211_1 \I1/low/U4/U28/U1/U1  ( .x(\I1/low/U4/U28/U1/clr ), .a(
        \I1/net20 ), .b(\I1/low/acb ), .c(\I1/low/nlocalcd ), .d(\I1/net32 )
         );
    nand3_1 \I1/low/U4/U28/U1/U2  ( .x(\I1/low/U4/U28/U1/set ), .a(
        \I1/low/nlocalcd ), .b(\I1/net20 ), .c(\I1/low/acb ) );
    nand2_2 \I1/low/U4/U28/U1/U3  ( .x(\I1/net32 ), .a(\I1/low/U4/U28/U1/clr ), 
        .b(\I1/low/U4/U28/U1/set ) );
    oai21_1 \I1/low/U1/U30/U1/U1  ( .x(\I1/low/acb ), .a(\I1/low/U1/Z ), .b(
        \I1/low/ba ), .c(\I1/net20 ) );
    inv_1 \I1/low/U1/U30/U1/U2  ( .x(\I1/low/U1/Z ), .a(\I1/low/acb ) );
    ao222_1 \I1/low/U5/U18/U1/U1  ( .x(\I1/low/ba ), .a(\I1/low/latch ), .b(
        pullcd), .c(\I1/low/latch ), .d(\I1/low/ba ), .e(pullcd), .f(
        \I1/low/ba ) );
    aoi222_1 \I1/low/U1664/U28/U30/U1  ( .x(\I1/low/U1664/x[3] ), .a(
        \I1/low/ncd[7] ), .b(\I1/low/ncd[6] ), .c(\I1/low/ncd[7] ), .d(
        \I1/low/U1664/U28/Z ), .e(\I1/low/ncd[6] ), .f(\I1/low/U1664/U28/Z )
         );
    inv_1 \I1/low/U1664/U28/U30/Uinv  ( .x(\I1/low/U1664/U28/Z ), .a(
        \I1/low/U1664/x[3] ) );
    aoi222_1 \I1/low/U1664/U32/U30/U1  ( .x(\I1/low/U1664/x[0] ), .a(
        \I1/low/ncd[1] ), .b(\I1/low/ncd[0] ), .c(\I1/low/ncd[1] ), .d(
        \I1/low/U1664/U32/Z ), .e(\I1/low/ncd[0] ), .f(\I1/low/U1664/U32/Z )
         );
    inv_1 \I1/low/U1664/U32/U30/Uinv  ( .x(\I1/low/U1664/U32/Z ), .a(
        \I1/low/U1664/x[0] ) );
    aoi222_1 \I1/low/U1664/U29/U30/U1  ( .x(\I1/low/U1664/x[2] ), .a(
        \I1/low/ncd[5] ), .b(\I1/low/ncd[4] ), .c(\I1/low/ncd[5] ), .d(
        \I1/low/U1664/U29/Z ), .e(\I1/low/ncd[4] ), .f(\I1/low/U1664/U29/Z )
         );
    inv_1 \I1/low/U1664/U29/U30/Uinv  ( .x(\I1/low/U1664/U29/Z ), .a(
        \I1/low/U1664/x[2] ) );
    aoi222_1 \I1/low/U1664/U33/U30/U1  ( .x(\I1/low/U1664/y[0] ), .a(
        \I1/low/U1664/x[1] ), .b(\I1/low/U1664/x[0] ), .c(\I1/low/U1664/x[1] ), 
        .d(\I1/low/U1664/U33/Z ), .e(\I1/low/U1664/x[0] ), .f(
        \I1/low/U1664/U33/Z ) );
    inv_1 \I1/low/U1664/U33/U30/Uinv  ( .x(\I1/low/U1664/U33/Z ), .a(
        \I1/low/U1664/y[0] ) );
    aoi222_1 \I1/low/U1664/U30/U30/U1  ( .x(\I1/low/U1664/y[1] ), .a(
        \I1/low/U1664/x[3] ), .b(\I1/low/U1664/x[2] ), .c(\I1/low/U1664/x[3] ), 
        .d(\I1/low/U1664/U30/Z ), .e(\I1/low/U1664/x[2] ), .f(
        \I1/low/U1664/U30/Z ) );
    inv_1 \I1/low/U1664/U30/U30/Uinv  ( .x(\I1/low/U1664/U30/Z ), .a(
        \I1/low/U1664/y[1] ) );
    aoi222_1 \I1/low/U1664/U31/U30/U1  ( .x(\I1/low/U1664/x[1] ), .a(
        \I1/low/ncd[3] ), .b(\I1/low/ncd[2] ), .c(\I1/low/ncd[3] ), .d(
        \I1/low/U1664/U31/Z ), .e(\I1/low/ncd[2] ), .f(\I1/low/U1664/U31/Z )
         );
    inv_1 \I1/low/U1664/U31/U30/Uinv  ( .x(\I1/low/U1664/U31/Z ), .a(
        \I1/low/U1664/x[1] ) );
    aoi222_1 \I1/low/U1664/U37/U30/U1  ( .x(\I1/low/localcd ), .a(
        \I1/low/U1664/y[0] ), .b(\I1/low/U1664/y[1] ), .c(\I1/low/U1664/y[0] ), 
        .d(\I1/low/U1664/U37/Z ), .e(\I1/low/U1664/y[1] ), .f(
        \I1/low/U1664/U37/Z ) );
    inv_1 \I1/low/U1664/U37/U30/Uinv  ( .x(\I1/low/U1664/U37/Z ), .a(
        \I1/low/localcd ) );
    nor3_1 \I1/low/U1669/Unr  ( .x(\I1/low/U1669/nr ), .a(
        \I1/low/ctrlack_internal ), .b(n5), .c(\I1/low/driveh ) );
    nand3_1 \I1/low/U1669/Und  ( .x(\I1/low/U1669/nd ), .a(
        \I1/low/ctrlack_internal ), .b(\I1/low/drivel ), .c(\I1/low/driveh )
         );
    oa21_1 \I1/low/U1669/U1  ( .x(\I1/low/U1669/n2 ), .a(\I1/low/U1669/n2 ), 
        .b(\I1/low/U1669/nr ), .c(\I1/low/U1669/nd ) );
    inv_2 \I1/low/U1669/U3  ( .x(net17), .a(\I1/low/U1669/n2 ) );
    buf_2 \I1/high/U1653  ( .x(\I1/high/latch ), .a(\I1/net33 ) );
    nor2_1 \I1/high/U264/U5  ( .x(\I1/high/nlocalcd ), .a(reset), .b(
        \I1/high/localcd ) );
    nor2_1 \I1/high/U1659_0_/U5  ( .x(\I1/high/ncd[0] ), .a(ol[24]), .b(oh[24]
        ) );
    nor2_1 \I1/high/U1659_1_/U5  ( .x(\I1/high/ncd[1] ), .a(ol[25]), .b(oh[25]
        ) );
    nor2_1 \I1/high/U1659_2_/U5  ( .x(\I1/high/ncd[2] ), .a(ol[26]), .b(oh[26]
        ) );
    nor2_1 \I1/high/U1659_3_/U5  ( .x(\I1/high/ncd[3] ), .a(ol[27]), .b(oh[27]
        ) );
    nor2_1 \I1/high/U1659_4_/U5  ( .x(\I1/high/ncd[4] ), .a(ol[28]), .b(oh[28]
        ) );
    nor2_1 \I1/high/U1659_5_/U5  ( .x(\I1/high/ncd[5] ), .a(ol[29]), .b(oh[29]
        ) );
    nor2_1 \I1/high/U1659_6_/U5  ( .x(\I1/high/ncd[6] ), .a(ol[30]), .b(oh[30]
        ) );
    nor2_1 \I1/high/U1659_7_/U5  ( .x(\I1/high/ncd[7] ), .a(ol[31]), .b(oh[31]
        ) );
    nor2_1 \I1/high/U3/U5  ( .x(\I1/high/ctrlack_internal ), .a(\I1/high/acb ), 
        .b(\I1/high/ba ) );
    buf_2 \I1/high/U1665/U7  ( .x(\I1/high/driveh ), .a(ctrlreq) );
    buf_2 \I1/high/U1666/U7  ( .x(\I1/high/drivel ), .a(ctrlreq) );
    ao23_1 \I1/high/U1658_0_/U21/U1/U1  ( .x(ol[24]), .a(\I1/high/driveh ), 
        .b(ol[24]), .c(n7), .d(pull_l[0]), .e(n8) );
    ao23_1 \I1/high/U1658_1_/U21/U1/U1  ( .x(ol[25]), .a(\I1/high/drivel ), 
        .b(ol[25]), .c(\I1/high/driveh ), .d(pull_l[1]), .e(n8) );
    ao23_1 \I1/high/U1658_2_/U21/U1/U1  ( .x(ol[26]), .a(\I1/high/drivel ), 
        .b(ol[26]), .c(\I1/high/driveh ), .d(pull_l[2]), .e(n8) );
    ao23_1 \I1/high/U1658_3_/U21/U1/U1  ( .x(ol[27]), .a(\I1/high/driveh ), 
        .b(ol[27]), .c(\I1/high/drivel ), .d(pull_l[3]), .e(\I1/high/latch )
         );
    ao23_1 \I1/high/U1658_4_/U21/U1/U1  ( .x(ol[28]), .a(n7), .b(ol[28]), .c(
        \I1/high/drivel ), .d(pull_l[4]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1658_5_/U21/U1/U1  ( .x(ol[29]), .a(\I1/high/driveh ), 
        .b(ol[29]), .c(n7), .d(pull_l[5]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1658_6_/U21/U1/U1  ( .x(ol[30]), .a(\I1/high/drivel ), 
        .b(ol[30]), .c(\I1/high/driveh ), .d(pull_l[6]), .e(\I1/high/latch )
         );
    ao23_1 \I1/high/U1658_7_/U21/U1/U1  ( .x(ol[31]), .a(n7), .b(ol[31]), .c(
        n7), .d(pull_l[7]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_0_/U21/U1/U1  ( .x(oh[24]), .a(\I1/high/driveh ), 
        .b(oh[24]), .c(n7), .d(pull_h[0]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_1_/U21/U1/U1  ( .x(oh[25]), .a(n7), .b(oh[25]), .c(
        \I1/high/drivel ), .d(pull_h[1]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_2_/U21/U1/U1  ( .x(oh[26]), .a(\I1/high/drivel ), 
        .b(oh[26]), .c(\I1/high/drivel ), .d(pull_h[2]), .e(\I1/high/latch )
         );
    ao23_1 \I1/high/U1651_3_/U21/U1/U1  ( .x(oh[27]), .a(n7), .b(oh[27]), .c(
        \I1/high/driveh ), .d(pull_h[3]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_4_/U21/U1/U1  ( .x(oh[28]), .a(n7), .b(oh[28]), .c(
        n7), .d(pull_h[4]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_5_/U21/U1/U1  ( .x(oh[29]), .a(\I1/high/drivel ), 
        .b(oh[29]), .c(n7), .d(pull_h[5]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_6_/U21/U1/U1  ( .x(oh[30]), .a(\I1/high/drivel ), 
        .b(oh[30]), .c(\I1/high/driveh ), .d(pull_h[6]), .e(\I1/high/latch )
         );
    ao23_1 \I1/high/U1651_7_/U21/U1/U1  ( .x(oh[31]), .a(\I1/high/driveh ), 
        .b(oh[31]), .c(\I1/high/drivel ), .d(pull_h[7]), .e(\I1/high/latch )
         );
    aoai211_1 \I1/high/U4/U28/U1/U1  ( .x(\I1/high/U4/U28/U1/clr ), .a(ctrlreq
        ), .b(\I1/high/acb ), .c(\I1/high/nlocalcd ), .d(\I1/net33 ) );
    nand3_1 \I1/high/U4/U28/U1/U2  ( .x(\I1/high/U4/U28/U1/set ), .a(
        \I1/high/nlocalcd ), .b(ctrlreq), .c(\I1/high/acb ) );
    nand2_2 \I1/high/U4/U28/U1/U3  ( .x(\I1/net33 ), .a(
        \I1/high/U4/U28/U1/clr ), .b(\I1/high/U4/U28/U1/set ) );
    oai21_1 \I1/high/U1/U30/U1/U1  ( .x(\I1/high/acb ), .a(\I1/high/U1/Z ), 
        .b(\I1/high/ba ), .c(ctrlreq) );
    inv_1 \I1/high/U1/U30/U1/U2  ( .x(\I1/high/U1/Z ), .a(\I1/high/acb ) );
    ao222_1 \I1/high/U5/U18/U1/U1  ( .x(\I1/high/ba ), .a(\I1/high/latch ), 
        .b(pullcd), .c(\I1/high/latch ), .d(\I1/high/ba ), .e(pullcd), .f(
        \I1/high/ba ) );
    aoi222_1 \I1/high/U1664/U28/U30/U1  ( .x(\I1/high/U1664/x[3] ), .a(
        \I1/high/ncd[7] ), .b(\I1/high/ncd[6] ), .c(\I1/high/ncd[7] ), .d(
        \I1/high/U1664/U28/Z ), .e(\I1/high/ncd[6] ), .f(\I1/high/U1664/U28/Z 
        ) );
    inv_1 \I1/high/U1664/U28/U30/Uinv  ( .x(\I1/high/U1664/U28/Z ), .a(
        \I1/high/U1664/x[3] ) );
    aoi222_1 \I1/high/U1664/U32/U30/U1  ( .x(\I1/high/U1664/x[0] ), .a(
        \I1/high/ncd[1] ), .b(\I1/high/ncd[0] ), .c(\I1/high/ncd[1] ), .d(
        \I1/high/U1664/U32/Z ), .e(\I1/high/ncd[0] ), .f(\I1/high/U1664/U32/Z 
        ) );
    inv_1 \I1/high/U1664/U32/U30/Uinv  ( .x(\I1/high/U1664/U32/Z ), .a(
        \I1/high/U1664/x[0] ) );
    aoi222_1 \I1/high/U1664/U29/U30/U1  ( .x(\I1/high/U1664/x[2] ), .a(
        \I1/high/ncd[5] ), .b(\I1/high/ncd[4] ), .c(\I1/high/ncd[5] ), .d(
        \I1/high/U1664/U29/Z ), .e(\I1/high/ncd[4] ), .f(\I1/high/U1664/U29/Z 
        ) );
    inv_1 \I1/high/U1664/U29/U30/Uinv  ( .x(\I1/high/U1664/U29/Z ), .a(
        \I1/high/U1664/x[2] ) );
    aoi222_1 \I1/high/U1664/U33/U30/U1  ( .x(\I1/high/U1664/y[0] ), .a(
        \I1/high/U1664/x[1] ), .b(\I1/high/U1664/x[0] ), .c(
        \I1/high/U1664/x[1] ), .d(\I1/high/U1664/U33/Z ), .e(
        \I1/high/U1664/x[0] ), .f(\I1/high/U1664/U33/Z ) );
    inv_1 \I1/high/U1664/U33/U30/Uinv  ( .x(\I1/high/U1664/U33/Z ), .a(
        \I1/high/U1664/y[0] ) );
    aoi222_1 \I1/high/U1664/U30/U30/U1  ( .x(\I1/high/U1664/y[1] ), .a(
        \I1/high/U1664/x[3] ), .b(\I1/high/U1664/x[2] ), .c(
        \I1/high/U1664/x[3] ), .d(\I1/high/U1664/U30/Z ), .e(
        \I1/high/U1664/x[2] ), .f(\I1/high/U1664/U30/Z ) );
    inv_1 \I1/high/U1664/U30/U30/Uinv  ( .x(\I1/high/U1664/U30/Z ), .a(
        \I1/high/U1664/y[1] ) );
    aoi222_1 \I1/high/U1664/U31/U30/U1  ( .x(\I1/high/U1664/x[1] ), .a(
        \I1/high/ncd[3] ), .b(\I1/high/ncd[2] ), .c(\I1/high/ncd[3] ), .d(
        \I1/high/U1664/U31/Z ), .e(\I1/high/ncd[2] ), .f(\I1/high/U1664/U31/Z 
        ) );
    inv_1 \I1/high/U1664/U31/U30/Uinv  ( .x(\I1/high/U1664/U31/Z ), .a(
        \I1/high/U1664/x[1] ) );
    aoi222_1 \I1/high/U1664/U37/U30/U1  ( .x(\I1/high/localcd ), .a(
        \I1/high/U1664/y[0] ), .b(\I1/high/U1664/y[1] ), .c(
        \I1/high/U1664/y[0] ), .d(\I1/high/U1664/U37/Z ), .e(
        \I1/high/U1664/y[1] ), .f(\I1/high/U1664/U37/Z ) );
    inv_1 \I1/high/U1664/U37/U30/Uinv  ( .x(\I1/high/U1664/U37/Z ), .a(
        \I1/high/localcd ) );
    nor3_1 \I1/high/U1669/Unr  ( .x(\I1/high/U1669/nr ), .a(
        \I1/high/ctrlack_internal ), .b(n7), .c(\I1/high/driveh ) );
    nand3_1 \I1/high/U1669/Und  ( .x(\I1/high/U1669/nd ), .a(
        \I1/high/ctrlack_internal ), .b(\I1/high/drivel ), .c(\I1/high/driveh 
        ) );
    oa21_1 \I1/high/U1669/U1  ( .x(\I1/high/U1669/n2 ), .a(\I1/high/U1669/n2 ), 
        .b(\I1/high/U1669/nr ), .c(\I1/high/U1669/nd ) );
    inv_2 \I1/high/U1669/U3  ( .x(\I1/net20 ), .a(\I1/high/U1669/n2 ) );
    buf_2 U1 ( .x(n1), .a(\I0/net20 ) );
    buf_1 U2 ( .x(n2), .a(\I0/low/latch ) );
    buf_2 U3 ( .x(n3), .a(net17) );
    buf_1 U4 ( .x(n4), .a(\I0/high/latch ) );
    buf_2 U5 ( .x(n5), .a(\I1/net20 ) );
    buf_1 U6 ( .x(n6), .a(\I1/low/latch ) );
    buf_2 U7 ( .x(n7), .a(ctrlreq) );
    buf_1 U8 ( .x(n8), .a(\I1/high/latch ) );
endmodule


module chain_fr2dr_byte_0 ( nia, oh, ol, i, nReset, noa );
output [7:0] oh;
output [7:0] ol;
input  [4:0] i;
input  nReset, noa;
output nia;
    wire nbReset, eop, ncla, csela, asela, \U891/reset , \U891/neopack , 
        \U891/iay , \U891/naack[0] , \U891/naack[1] , \U891/U1128/nb , \b[3] , 
        \b[2] , \U891/U1128/na , \b[1] , \b[0] , \U891/ackb , \a[3] , \a[2] , 
        \U891/nack , \U891/acka , \a[1] , \a[0] , bsela, bsel, asel, 
        \U891/U1118_0_/nr , naa, \U891/U1118_0_/nd , \U891/U1118_0_/n2 , 
        \U891/U1118_1_/nr , \U891/U1118_1_/nd , \U891/U1118_1_/n2 , 
        \U891/U1118_2_/nr , \U891/U1118_2_/nd , \U891/U1118_2_/n2 , 
        \U891/U1118_3_/nr , \U891/U1118_3_/nd , \U891/U1118_3_/n2 , 
        \U891/U1117_0_/nr , nba, \U891/U1117_0_/nd , \U891/U1117_0_/n2 , 
        \U891/U1117_1_/nr , \U891/U1117_1_/nd , \U891/U1117_1_/n2 , 
        \U891/U1117_2_/nr , \U891/U1117_2_/nd , \U891/U1117_2_/n2 , 
        \U891/U1117_3_/nr , \U891/U1117_3_/nd , \U891/U1117_3_/n2 , 
        \U886/reset , \U886/U1128/nb , \f[3] , \f[2] , \U886/U1128/na , \f[1] , 
        \f[0] , \U886/ackb , \U886/nack , \U886/acka , \U886/U1127/n5 , 
        \U886/U1127/n1 , \U886/U1127/n2 , \U886/U1127/n3 , \U886/U1127/n4 , 
        \e[3] , \e[2] , \e[1] , \e[0] , fsela, fsel, esela, esel, 
        \U886/U1118_0_/nr , nea, \U886/U1118_0_/nd , \U886/U1118_0_/n2 , 
        \U886/U1118_1_/nr , \U886/U1118_1_/nd , \U886/U1118_1_/n2 , 
        \U886/U1118_2_/nr , \U886/U1118_2_/nd , \U886/U1118_2_/n2 , 
        \U886/U1118_3_/nr , \U886/U1118_3_/nd , \U886/U1118_3_/n2 , 
        \U886/U1117_0_/nr , nfa, \U886/U1117_0_/nd , \U886/U1117_0_/n2 , 
        \U886/U1117_1_/nr , \U886/U1117_1_/nd , \U886/U1117_1_/n2 , 
        \U886/U1117_2_/nr , \U886/U1117_2_/nd , \U886/U1117_2_/n2 , 
        \U886/U1117_3_/nr , \U886/U1117_3_/nd , \U886/U1117_3_/n2 , 
        \U884/reset , \U884/U1128/nb , \d[3] , \d[2] , \U884/U1128/na , \d[1] , 
        \d[0] , \U884/ackb , \U884/nack , \U884/acka , \U884/U1127/n5 , 
        \U884/U1127/n1 , \U884/U1127/n2 , \U884/U1127/n3 , \U884/U1127/n4 , 
        \c[3] , \c[2] , \c[1] , \c[0] , dsela, dsel, csel, \U884/U1118_0_/nr , 
        nca, \U884/U1118_0_/nd , \U884/U1118_0_/n2 , \U884/U1118_1_/nr , 
        \U884/U1118_1_/nd , \U884/U1118_1_/n2 , \U884/U1118_2_/nr , 
        \U884/U1118_2_/nd , \U884/U1118_2_/n2 , \U884/U1118_3_/nr , 
        \U884/U1118_3_/nd , \U884/U1118_3_/n2 , \U884/U1117_0_/nr , nda, 
        \U884/U1117_0_/nd , \U884/U1117_0_/n2 , \U884/U1117_1_/nr , 
        \U884/U1117_1_/nd , \U884/U1117_1_/n2 , \U884/U1117_2_/nr , 
        \U884/U1117_2_/nd , \U884/U1117_2_/n2 , \U884/U1117_3_/nr , 
        \U884/U1117_3_/nd , \U884/U1117_3_/n2 , \U888/s , \U888/r , 
        \U888/nback , \U888/naack , \U888/reset , \U887/s , \U887/r , 
        \U887/nback , \U887/naack , \U887/reset , \U885/s , \U885/r , 
        \U885/nback , \U885/naack , \U885/reset , \U877/x , \U877/reset , 
        \U877/y , \U877/U590/U25/U1/clr , net135, \cl[3] , \cl[1] , 
        \U877/U590/U25/U1/ob , n1, \U877/U589/U25/U1/clr , \cl[0] , 
        \U877/U589/U25/U1/ob , \U877/U588/U25/U1/clr , \cl[2] , 
        \U877/U588/U25/U1/ob , \U877/U591/U25/U1/clr , \U877/U591/U25/U1/ob , 
        \U876/x , \U876/reset , \U876/y , \U876/U590/U25/U1/clr , 
        \U876/U590/U25/U1/ob , \U876/U589/U25/U1/clr , \U876/U589/U25/U1/ob , 
        \U876/U588/U25/U1/clr , \U876/U588/U25/U1/ob , \U876/U591/U25/U1/clr , 
        \U876/U591/U25/U1/ob , \U2/x , \U2/reset , \U2/y , 
        \U2/U590/U25/U1/clr , \U2/U590/U25/U1/ob , \U2/U589/U25/U1/clr , 
        \U2/U589/U25/U1/ob , \U2/U588/U25/U1/clr , \U2/U588/U25/U1/ob , 
        \U2/U591/U25/U1/clr , \U2/U591/U25/U1/ob , \U1/x , \U1/reset , \U1/y , 
        \U1/U590/U25/U1/clr , \U1/U590/U25/U1/ob , \U1/U589/U25/U1/clr , 
        \U1/U589/U25/U1/ob , \U1/U588/U25/U1/clr , \U1/U588/U25/U1/ob , 
        \U1/U591/U25/U1/clr , \U1/U591/U25/U1/ob , \U881/nack[1] , 
        \U881/nack[0] ;
    buf_2 U897 ( .x(nbReset), .a(nReset) );
    and4_1 \U894/U12  ( .x(eop), .a(ncla), .b(csela), .c(asela), .d(i[4]) );
    inv_1 \U891/U1126/U3  ( .x(\U891/reset ), .a(nbReset) );
    inv_1 \U891/U1139/U3  ( .x(\U891/neopack ), .a(eop) );
    nand3_1 \U891/U1131/U9  ( .x(\U891/iay ), .a(\U891/neopack ), .b(
        \U891/naack[0] ), .c(\U891/naack[1] ) );
    nor3_1 \U891/U1128/U27  ( .x(\U891/U1128/nb ), .a(\U891/reset ), .b(\b[3] 
        ), .c(\b[2] ) );
    nor2_1 \U891/U1128/U26  ( .x(\U891/U1128/na ), .a(\b[1] ), .b(\b[0] ) );
    nand2_2 \U891/U1128/U29  ( .x(\U891/ackb ), .a(\U891/U1128/nb ), .b(
        \U891/U1128/na ) );
    nor2_1 \U891/U1133/U5  ( .x(\U891/naack[0] ), .a(\a[3] ), .b(\a[2] ) );
    nor2_1 \U891/U1108/U5  ( .x(\U891/nack ), .a(\U891/acka ), .b(\U891/ackb )
         );
    nor2_1 \U891/U1134/U5  ( .x(\U891/naack[1] ), .a(\a[1] ), .b(\a[0] ) );
    nor2_2 \U891/U914/U6  ( .x(nia), .a(\U891/iay ), .b(\U891/ackb ) );
    nand2_1 \U891/U1130/U5  ( .x(\U891/acka ), .a(\U891/naack[0] ), .b(
        \U891/naack[1] ) );
    ao222_4 \U891/U1121/U1/U1  ( .x(bsela), .a(\U891/nack ), .b(bsel), .c(
        \U891/nack ), .d(bsela), .e(bsel), .f(bsela) );
    ao222_4 \U891/U1120/U1/U1  ( .x(asela), .a(asel), .b(\U891/nack ), .c(asel
        ), .d(asela), .e(\U891/nack ), .f(asela) );
    nor3_1 \U891/U1118_0_/Unr  ( .x(\U891/U1118_0_/nr ), .a(i[0]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_0_/Und  ( .x(\U891/U1118_0_/nd ), .a(i[0]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_0_/U1  ( .x(\U891/U1118_0_/n2 ), .a(\U891/U1118_0_/n2 ), 
        .b(\U891/U1118_0_/nr ), .c(\U891/U1118_0_/nd ) );
    inv_2 \U891/U1118_0_/U3  ( .x(\a[0] ), .a(\U891/U1118_0_/n2 ) );
    nor3_1 \U891/U1118_1_/Unr  ( .x(\U891/U1118_1_/nr ), .a(i[1]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_1_/Und  ( .x(\U891/U1118_1_/nd ), .a(i[1]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_1_/U1  ( .x(\U891/U1118_1_/n2 ), .a(\U891/U1118_1_/n2 ), 
        .b(\U891/U1118_1_/nr ), .c(\U891/U1118_1_/nd ) );
    inv_2 \U891/U1118_1_/U3  ( .x(\a[1] ), .a(\U891/U1118_1_/n2 ) );
    nor3_1 \U891/U1118_2_/Unr  ( .x(\U891/U1118_2_/nr ), .a(i[2]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_2_/Und  ( .x(\U891/U1118_2_/nd ), .a(i[2]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_2_/U1  ( .x(\U891/U1118_2_/n2 ), .a(\U891/U1118_2_/n2 ), 
        .b(\U891/U1118_2_/nr ), .c(\U891/U1118_2_/nd ) );
    inv_2 \U891/U1118_2_/U3  ( .x(\a[2] ), .a(\U891/U1118_2_/n2 ) );
    nor3_1 \U891/U1118_3_/Unr  ( .x(\U891/U1118_3_/nr ), .a(i[3]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_3_/Und  ( .x(\U891/U1118_3_/nd ), .a(i[3]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_3_/U1  ( .x(\U891/U1118_3_/n2 ), .a(\U891/U1118_3_/n2 ), 
        .b(\U891/U1118_3_/nr ), .c(\U891/U1118_3_/nd ) );
    inv_2 \U891/U1118_3_/U3  ( .x(\a[3] ), .a(\U891/U1118_3_/n2 ) );
    nor3_1 \U891/U1117_0_/Unr  ( .x(\U891/U1117_0_/nr ), .a(i[0]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_0_/Und  ( .x(\U891/U1117_0_/nd ), .a(i[0]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_0_/U1  ( .x(\U891/U1117_0_/n2 ), .a(\U891/U1117_0_/n2 ), 
        .b(\U891/U1117_0_/nr ), .c(\U891/U1117_0_/nd ) );
    inv_2 \U891/U1117_0_/U3  ( .x(\b[0] ), .a(\U891/U1117_0_/n2 ) );
    nor3_1 \U891/U1117_1_/Unr  ( .x(\U891/U1117_1_/nr ), .a(i[1]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_1_/Und  ( .x(\U891/U1117_1_/nd ), .a(i[1]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_1_/U1  ( .x(\U891/U1117_1_/n2 ), .a(\U891/U1117_1_/n2 ), 
        .b(\U891/U1117_1_/nr ), .c(\U891/U1117_1_/nd ) );
    inv_2 \U891/U1117_1_/U3  ( .x(\b[1] ), .a(\U891/U1117_1_/n2 ) );
    nor3_1 \U891/U1117_2_/Unr  ( .x(\U891/U1117_2_/nr ), .a(i[2]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_2_/Und  ( .x(\U891/U1117_2_/nd ), .a(i[2]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_2_/U1  ( .x(\U891/U1117_2_/n2 ), .a(\U891/U1117_2_/n2 ), 
        .b(\U891/U1117_2_/nr ), .c(\U891/U1117_2_/nd ) );
    inv_2 \U891/U1117_2_/U3  ( .x(\b[2] ), .a(\U891/U1117_2_/n2 ) );
    nor3_1 \U891/U1117_3_/Unr  ( .x(\U891/U1117_3_/nr ), .a(i[3]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_3_/Und  ( .x(\U891/U1117_3_/nd ), .a(i[3]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_3_/U1  ( .x(\U891/U1117_3_/n2 ), .a(\U891/U1117_3_/n2 ), 
        .b(\U891/U1117_3_/nr ), .c(\U891/U1117_3_/nd ) );
    inv_2 \U891/U1117_3_/U3  ( .x(\b[3] ), .a(\U891/U1117_3_/n2 ) );
    inv_1 \U886/U1126/U3  ( .x(\U886/reset ), .a(nbReset) );
    nor3_1 \U886/U1128/U27  ( .x(\U886/U1128/nb ), .a(\U886/reset ), .b(\f[3] 
        ), .c(\f[2] ) );
    nor2_1 \U886/U1128/U26  ( .x(\U886/U1128/na ), .a(\f[1] ), .b(\f[0] ) );
    nand2_2 \U886/U1128/U29  ( .x(\U886/ackb ), .a(\U886/U1128/nb ), .b(
        \U886/U1128/na ) );
    nor2_1 \U886/U1108/U5  ( .x(\U886/nack ), .a(\U886/acka ), .b(\U886/ackb )
         );
    nor2_2 \U886/U914/U6  ( .x(nba), .a(\U886/acka ), .b(\U886/ackb ) );
    and4_1 \U886/U1127/U25  ( .x(\U886/U1127/n5 ), .a(\U886/U1127/n1 ), .b(
        \U886/U1127/n2 ), .c(\U886/U1127/n3 ), .d(\U886/U1127/n4 ) );
    inv_1 \U886/U1127/U1  ( .x(\U886/U1127/n1 ), .a(\e[3] ) );
    inv_1 \U886/U1127/U2  ( .x(\U886/U1127/n2 ), .a(\e[2] ) );
    inv_1 \U886/U1127/U3  ( .x(\U886/U1127/n3 ), .a(\e[1] ) );
    inv_1 \U886/U1127/U4  ( .x(\U886/U1127/n4 ), .a(\e[0] ) );
    inv_2 \U886/U1127/U5  ( .x(\U886/acka ), .a(\U886/U1127/n5 ) );
    ao222_2 \U886/U1121/U19/U1/U1  ( .x(fsela), .a(\U886/nack ), .b(fsel), .c(
        \U886/nack ), .d(fsela), .e(fsel), .f(fsela) );
    ao222_2 \U886/U1120/U19/U1/U1  ( .x(esela), .a(esel), .b(\U886/nack ), .c(
        esel), .d(esela), .e(\U886/nack ), .f(esela) );
    nor3_1 \U886/U1118_0_/Unr  ( .x(\U886/U1118_0_/nr ), .a(\b[0] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_0_/Und  ( .x(\U886/U1118_0_/nd ), .a(\b[0] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_0_/U1  ( .x(\U886/U1118_0_/n2 ), .a(\U886/U1118_0_/n2 ), 
        .b(\U886/U1118_0_/nr ), .c(\U886/U1118_0_/nd ) );
    inv_2 \U886/U1118_0_/U3  ( .x(\e[0] ), .a(\U886/U1118_0_/n2 ) );
    nor3_1 \U886/U1118_1_/Unr  ( .x(\U886/U1118_1_/nr ), .a(\b[1] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_1_/Und  ( .x(\U886/U1118_1_/nd ), .a(\b[1] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_1_/U1  ( .x(\U886/U1118_1_/n2 ), .a(\U886/U1118_1_/n2 ), 
        .b(\U886/U1118_1_/nr ), .c(\U886/U1118_1_/nd ) );
    inv_2 \U886/U1118_1_/U3  ( .x(\e[1] ), .a(\U886/U1118_1_/n2 ) );
    nor3_1 \U886/U1118_2_/Unr  ( .x(\U886/U1118_2_/nr ), .a(\b[2] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_2_/Und  ( .x(\U886/U1118_2_/nd ), .a(\b[2] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_2_/U1  ( .x(\U886/U1118_2_/n2 ), .a(\U886/U1118_2_/n2 ), 
        .b(\U886/U1118_2_/nr ), .c(\U886/U1118_2_/nd ) );
    inv_2 \U886/U1118_2_/U3  ( .x(\e[2] ), .a(\U886/U1118_2_/n2 ) );
    nor3_1 \U886/U1118_3_/Unr  ( .x(\U886/U1118_3_/nr ), .a(\b[3] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_3_/Und  ( .x(\U886/U1118_3_/nd ), .a(\b[3] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_3_/U1  ( .x(\U886/U1118_3_/n2 ), .a(\U886/U1118_3_/n2 ), 
        .b(\U886/U1118_3_/nr ), .c(\U886/U1118_3_/nd ) );
    inv_2 \U886/U1118_3_/U3  ( .x(\e[3] ), .a(\U886/U1118_3_/n2 ) );
    nor3_1 \U886/U1117_0_/Unr  ( .x(\U886/U1117_0_/nr ), .a(\b[0] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_0_/Und  ( .x(\U886/U1117_0_/nd ), .a(\b[0] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_0_/U1  ( .x(\U886/U1117_0_/n2 ), .a(\U886/U1117_0_/n2 ), 
        .b(\U886/U1117_0_/nr ), .c(\U886/U1117_0_/nd ) );
    inv_2 \U886/U1117_0_/U3  ( .x(\f[0] ), .a(\U886/U1117_0_/n2 ) );
    nor3_1 \U886/U1117_1_/Unr  ( .x(\U886/U1117_1_/nr ), .a(\b[1] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_1_/Und  ( .x(\U886/U1117_1_/nd ), .a(\b[1] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_1_/U1  ( .x(\U886/U1117_1_/n2 ), .a(\U886/U1117_1_/n2 ), 
        .b(\U886/U1117_1_/nr ), .c(\U886/U1117_1_/nd ) );
    inv_2 \U886/U1117_1_/U3  ( .x(\f[1] ), .a(\U886/U1117_1_/n2 ) );
    nor3_1 \U886/U1117_2_/Unr  ( .x(\U886/U1117_2_/nr ), .a(\b[2] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_2_/Und  ( .x(\U886/U1117_2_/nd ), .a(\b[2] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_2_/U1  ( .x(\U886/U1117_2_/n2 ), .a(\U886/U1117_2_/n2 ), 
        .b(\U886/U1117_2_/nr ), .c(\U886/U1117_2_/nd ) );
    inv_2 \U886/U1117_2_/U3  ( .x(\f[2] ), .a(\U886/U1117_2_/n2 ) );
    nor3_1 \U886/U1117_3_/Unr  ( .x(\U886/U1117_3_/nr ), .a(\b[3] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_3_/Und  ( .x(\U886/U1117_3_/nd ), .a(\b[3] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_3_/U1  ( .x(\U886/U1117_3_/n2 ), .a(\U886/U1117_3_/n2 ), 
        .b(\U886/U1117_3_/nr ), .c(\U886/U1117_3_/nd ) );
    inv_2 \U886/U1117_3_/U3  ( .x(\f[3] ), .a(\U886/U1117_3_/n2 ) );
    inv_1 \U884/U1126/U3  ( .x(\U884/reset ), .a(nbReset) );
    nor3_1 \U884/U1128/U27  ( .x(\U884/U1128/nb ), .a(\U884/reset ), .b(\d[3] 
        ), .c(\d[2] ) );
    nor2_1 \U884/U1128/U26  ( .x(\U884/U1128/na ), .a(\d[1] ), .b(\d[0] ) );
    nand2_2 \U884/U1128/U29  ( .x(\U884/ackb ), .a(\U884/U1128/nb ), .b(
        \U884/U1128/na ) );
    nor2_1 \U884/U1108/U5  ( .x(\U884/nack ), .a(\U884/acka ), .b(\U884/ackb )
         );
    nor2_2 \U884/U914/U6  ( .x(naa), .a(\U884/acka ), .b(\U884/ackb ) );
    and4_1 \U884/U1127/U25  ( .x(\U884/U1127/n5 ), .a(\U884/U1127/n1 ), .b(
        \U884/U1127/n2 ), .c(\U884/U1127/n3 ), .d(\U884/U1127/n4 ) );
    inv_1 \U884/U1127/U1  ( .x(\U884/U1127/n1 ), .a(\c[3] ) );
    inv_1 \U884/U1127/U2  ( .x(\U884/U1127/n2 ), .a(\c[2] ) );
    inv_1 \U884/U1127/U3  ( .x(\U884/U1127/n3 ), .a(\c[1] ) );
    inv_1 \U884/U1127/U4  ( .x(\U884/U1127/n4 ), .a(\c[0] ) );
    inv_2 \U884/U1127/U5  ( .x(\U884/acka ), .a(\U884/U1127/n5 ) );
    ao222_2 \U884/U1121/U19/U1/U1  ( .x(dsela), .a(\U884/nack ), .b(dsel), .c(
        \U884/nack ), .d(dsela), .e(dsel), .f(dsela) );
    ao222_2 \U884/U1120/U19/U1/U1  ( .x(csela), .a(csel), .b(\U884/nack ), .c(
        csel), .d(csela), .e(\U884/nack ), .f(csela) );
    nor3_1 \U884/U1118_0_/Unr  ( .x(\U884/U1118_0_/nr ), .a(\a[0] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_0_/Und  ( .x(\U884/U1118_0_/nd ), .a(\a[0] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_0_/U1  ( .x(\U884/U1118_0_/n2 ), .a(\U884/U1118_0_/n2 ), 
        .b(\U884/U1118_0_/nr ), .c(\U884/U1118_0_/nd ) );
    inv_2 \U884/U1118_0_/U3  ( .x(\c[0] ), .a(\U884/U1118_0_/n2 ) );
    nor3_1 \U884/U1118_1_/Unr  ( .x(\U884/U1118_1_/nr ), .a(\a[1] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_1_/Und  ( .x(\U884/U1118_1_/nd ), .a(\a[1] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_1_/U1  ( .x(\U884/U1118_1_/n2 ), .a(\U884/U1118_1_/n2 ), 
        .b(\U884/U1118_1_/nr ), .c(\U884/U1118_1_/nd ) );
    inv_2 \U884/U1118_1_/U3  ( .x(\c[1] ), .a(\U884/U1118_1_/n2 ) );
    nor3_1 \U884/U1118_2_/Unr  ( .x(\U884/U1118_2_/nr ), .a(\a[2] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_2_/Und  ( .x(\U884/U1118_2_/nd ), .a(\a[2] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_2_/U1  ( .x(\U884/U1118_2_/n2 ), .a(\U884/U1118_2_/n2 ), 
        .b(\U884/U1118_2_/nr ), .c(\U884/U1118_2_/nd ) );
    inv_2 \U884/U1118_2_/U3  ( .x(\c[2] ), .a(\U884/U1118_2_/n2 ) );
    nor3_1 \U884/U1118_3_/Unr  ( .x(\U884/U1118_3_/nr ), .a(\a[3] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_3_/Und  ( .x(\U884/U1118_3_/nd ), .a(\a[3] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_3_/U1  ( .x(\U884/U1118_3_/n2 ), .a(\U884/U1118_3_/n2 ), 
        .b(\U884/U1118_3_/nr ), .c(\U884/U1118_3_/nd ) );
    inv_2 \U884/U1118_3_/U3  ( .x(\c[3] ), .a(\U884/U1118_3_/n2 ) );
    nor3_1 \U884/U1117_0_/Unr  ( .x(\U884/U1117_0_/nr ), .a(\a[0] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_0_/Und  ( .x(\U884/U1117_0_/nd ), .a(\a[0] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_0_/U1  ( .x(\U884/U1117_0_/n2 ), .a(\U884/U1117_0_/n2 ), 
        .b(\U884/U1117_0_/nr ), .c(\U884/U1117_0_/nd ) );
    inv_2 \U884/U1117_0_/U3  ( .x(\d[0] ), .a(\U884/U1117_0_/n2 ) );
    nor3_1 \U884/U1117_1_/Unr  ( .x(\U884/U1117_1_/nr ), .a(\a[1] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_1_/Und  ( .x(\U884/U1117_1_/nd ), .a(\a[1] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_1_/U1  ( .x(\U884/U1117_1_/n2 ), .a(\U884/U1117_1_/n2 ), 
        .b(\U884/U1117_1_/nr ), .c(\U884/U1117_1_/nd ) );
    inv_2 \U884/U1117_1_/U3  ( .x(\d[1] ), .a(\U884/U1117_1_/n2 ) );
    nor3_1 \U884/U1117_2_/Unr  ( .x(\U884/U1117_2_/nr ), .a(\a[2] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_2_/Und  ( .x(\U884/U1117_2_/nd ), .a(\a[2] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_2_/U1  ( .x(\U884/U1117_2_/n2 ), .a(\U884/U1117_2_/n2 ), 
        .b(\U884/U1117_2_/nr ), .c(\U884/U1117_2_/nd ) );
    inv_2 \U884/U1117_2_/U3  ( .x(\d[2] ), .a(\U884/U1117_2_/n2 ) );
    nor3_1 \U884/U1117_3_/Unr  ( .x(\U884/U1117_3_/nr ), .a(\a[3] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_3_/Und  ( .x(\U884/U1117_3_/nd ), .a(\a[3] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_3_/U1  ( .x(\U884/U1117_3_/n2 ), .a(\U884/U1117_3_/n2 ), 
        .b(\U884/U1117_3_/nr ), .c(\U884/U1117_3_/nd ) );
    inv_2 \U884/U1117_3_/U3  ( .x(\d[3] ), .a(\U884/U1117_3_/n2 ) );
    nand2_1 \U888/U1128/U5  ( .x(\U888/s ), .a(\U888/r ), .b(\U888/nback ) );
    nand2_1 \U888/U1103/U5  ( .x(\U888/r ), .a(\U888/naack ), .b(\U888/s ) );
    inv_1 \U888/U1111/U3  ( .x(\U888/reset ), .a(nbReset) );
    inv_1 \U888/U1112/U3  ( .x(\U888/naack ), .a(esela) );
    nor2_1 \U888/U1127/U5  ( .x(\U888/nback ), .a(fsela), .b(\U888/reset ) );
    and2_2 \U888/U1129/U8  ( .x(esel), .a(\U888/nback ), .b(\U888/s ) );
    and2_2 \U888/U1124/U8  ( .x(fsel), .a(\U888/r ), .b(\U888/naack ) );
    nand2_1 \U887/U1128/U5  ( .x(\U887/s ), .a(\U887/r ), .b(\U887/nback ) );
    nand2_1 \U887/U1103/U5  ( .x(\U887/r ), .a(\U887/naack ), .b(\U887/s ) );
    inv_1 \U887/U1111/U3  ( .x(\U887/reset ), .a(nbReset) );
    inv_1 \U887/U1112/U3  ( .x(\U887/naack ), .a(csela) );
    nor2_1 \U887/U1127/U5  ( .x(\U887/nback ), .a(dsela), .b(\U887/reset ) );
    and2_2 \U887/U1129/U8  ( .x(csel), .a(\U887/nback ), .b(\U887/s ) );
    and2_2 \U887/U1124/U8  ( .x(dsel), .a(\U887/r ), .b(\U887/naack ) );
    nand2_1 \U885/U1128/U5  ( .x(\U885/s ), .a(\U885/r ), .b(\U885/nback ) );
    nand2_1 \U885/U1103/U5  ( .x(\U885/r ), .a(\U885/naack ), .b(\U885/s ) );
    inv_1 \U885/U1111/U3  ( .x(\U885/reset ), .a(nbReset) );
    inv_1 \U885/U1112/U3  ( .x(\U885/naack ), .a(asela) );
    nor2_1 \U885/U1127/U5  ( .x(\U885/nback ), .a(bsela), .b(\U885/reset ) );
    and2_2 \U885/U1129/U8  ( .x(asel), .a(\U885/nback ), .b(\U885/s ) );
    and2_2 \U885/U1124/U8  ( .x(bsel), .a(\U885/r ), .b(\U885/naack ) );
    nor3_1 \U877/U594/U7  ( .x(\U877/x ), .a(ol[7]), .b(\U877/reset ), .c(oh
        [7]) );
    nor3_1 \U877/U593/U7  ( .x(\U877/y ), .a(ol[6]), .b(\U877/reset ), .c(oh
        [6]) );
    inv_1 \U877/U604/U3  ( .x(\U877/reset ), .a(nbReset) );
    oa31_1 \U877/U590/U25/U1/Uclr  ( .x(\U877/U590/U25/U1/clr ), .a(net135), 
        .b(\cl[3] ), .c(\cl[1] ), .d(oh[6]) );
    oaoi211_1 \U877/U590/U25/U1/Uaoi  ( .x(\U877/U590/U25/U1/ob ), .a(\cl[3] ), 
        .b(\cl[1] ), .c(n1), .d(\U877/U590/U25/U1/clr ) );
    inv_2 \U877/U590/U25/U1/Ui  ( .x(oh[6]), .a(\U877/U590/U25/U1/ob ) );
    oa31_1 \U877/U589/U25/U1/Uclr  ( .x(\U877/U589/U25/U1/clr ), .a(net135), 
        .b(\cl[1] ), .c(\cl[0] ), .d(ol[7]) );
    oaoi211_1 \U877/U589/U25/U1/Uaoi  ( .x(\U877/U589/U25/U1/ob ), .a(\cl[1] ), 
        .b(\cl[0] ), .c(n1), .d(\U877/U589/U25/U1/clr ) );
    inv_2 \U877/U589/U25/U1/Ui  ( .x(ol[7]), .a(\U877/U589/U25/U1/ob ) );
    oa31_1 \U877/U588/U25/U1/Uclr  ( .x(\U877/U588/U25/U1/clr ), .a(net135), 
        .b(\cl[3] ), .c(\cl[2] ), .d(oh[7]) );
    oaoi211_1 \U877/U588/U25/U1/Uaoi  ( .x(\U877/U588/U25/U1/ob ), .a(\cl[3] ), 
        .b(\cl[2] ), .c(n1), .d(\U877/U588/U25/U1/clr ) );
    inv_2 \U877/U588/U25/U1/Ui  ( .x(oh[7]), .a(\U877/U588/U25/U1/ob ) );
    oa31_1 \U877/U591/U25/U1/Uclr  ( .x(\U877/U591/U25/U1/clr ), .a(net135), 
        .b(\cl[2] ), .c(\cl[0] ), .d(ol[6]) );
    oaoi211_1 \U877/U591/U25/U1/Uaoi  ( .x(\U877/U591/U25/U1/ob ), .a(\cl[2] ), 
        .b(\cl[0] ), .c(n1), .d(\U877/U591/U25/U1/clr ) );
    inv_2 \U877/U591/U25/U1/Ui  ( .x(ol[6]), .a(\U877/U591/U25/U1/ob ) );
    ao222_2 \U877/U592/U19/U1/U1  ( .x(ncla), .a(\U877/x ), .b(\U877/y ), .c(
        \U877/x ), .d(ncla), .e(\U877/y ), .f(ncla) );
    nor3_1 \U876/U594/U7  ( .x(\U876/x ), .a(ol[3]), .b(\U876/reset ), .c(oh
        [3]) );
    nor3_1 \U876/U593/U7  ( .x(\U876/y ), .a(ol[2]), .b(\U876/reset ), .c(oh
        [2]) );
    inv_1 \U876/U604/U3  ( .x(\U876/reset ), .a(nbReset) );
    oa31_1 \U876/U590/U25/U1/Uclr  ( .x(\U876/U590/U25/U1/clr ), .a(net135), 
        .b(\d[3] ), .c(\d[1] ), .d(oh[2]) );
    oaoi211_1 \U876/U590/U25/U1/Uaoi  ( .x(\U876/U590/U25/U1/ob ), .a(\d[3] ), 
        .b(\d[1] ), .c(n1), .d(\U876/U590/U25/U1/clr ) );
    inv_2 \U876/U590/U25/U1/Ui  ( .x(oh[2]), .a(\U876/U590/U25/U1/ob ) );
    oa31_1 \U876/U589/U25/U1/Uclr  ( .x(\U876/U589/U25/U1/clr ), .a(net135), 
        .b(\d[1] ), .c(\d[0] ), .d(ol[3]) );
    oaoi211_1 \U876/U589/U25/U1/Uaoi  ( .x(\U876/U589/U25/U1/ob ), .a(\d[1] ), 
        .b(\d[0] ), .c(n1), .d(\U876/U589/U25/U1/clr ) );
    inv_2 \U876/U589/U25/U1/Ui  ( .x(ol[3]), .a(\U876/U589/U25/U1/ob ) );
    oa31_1 \U876/U588/U25/U1/Uclr  ( .x(\U876/U588/U25/U1/clr ), .a(net135), 
        .b(\d[3] ), .c(\d[2] ), .d(oh[3]) );
    oaoi211_1 \U876/U588/U25/U1/Uaoi  ( .x(\U876/U588/U25/U1/ob ), .a(\d[3] ), 
        .b(\d[2] ), .c(n1), .d(\U876/U588/U25/U1/clr ) );
    inv_2 \U876/U588/U25/U1/Ui  ( .x(oh[3]), .a(\U876/U588/U25/U1/ob ) );
    oa31_1 \U876/U591/U25/U1/Uclr  ( .x(\U876/U591/U25/U1/clr ), .a(net135), 
        .b(\d[2] ), .c(\d[0] ), .d(ol[2]) );
    oaoi211_1 \U876/U591/U25/U1/Uaoi  ( .x(\U876/U591/U25/U1/ob ), .a(\d[2] ), 
        .b(\d[0] ), .c(n1), .d(\U876/U591/U25/U1/clr ) );
    inv_2 \U876/U591/U25/U1/Ui  ( .x(ol[2]), .a(\U876/U591/U25/U1/ob ) );
    ao222_2 \U876/U592/U19/U1/U1  ( .x(nda), .a(\U876/x ), .b(\U876/y ), .c(
        \U876/x ), .d(nda), .e(\U876/y ), .f(nda) );
    nor3_1 \U2/U594/U7  ( .x(\U2/x ), .a(ol[1]), .b(\U2/reset ), .c(oh[1]) );
    nor3_1 \U2/U593/U7  ( .x(\U2/y ), .a(ol[0]), .b(\U2/reset ), .c(oh[0]) );
    inv_1 \U2/U604/U3  ( .x(\U2/reset ), .a(nbReset) );
    oa31_1 \U2/U590/U25/U1/Uclr  ( .x(\U2/U590/U25/U1/clr ), .a(net135), .b(
        \f[3] ), .c(\f[1] ), .d(oh[0]) );
    oaoi211_1 \U2/U590/U25/U1/Uaoi  ( .x(\U2/U590/U25/U1/ob ), .a(\f[3] ), .b(
        \f[1] ), .c(n1), .d(\U2/U590/U25/U1/clr ) );
    inv_2 \U2/U590/U25/U1/Ui  ( .x(oh[0]), .a(\U2/U590/U25/U1/ob ) );
    oa31_1 \U2/U589/U25/U1/Uclr  ( .x(\U2/U589/U25/U1/clr ), .a(net135), .b(
        \f[1] ), .c(\f[0] ), .d(ol[1]) );
    oaoi211_1 \U2/U589/U25/U1/Uaoi  ( .x(\U2/U589/U25/U1/ob ), .a(\f[1] ), .b(
        \f[0] ), .c(n1), .d(\U2/U589/U25/U1/clr ) );
    inv_2 \U2/U589/U25/U1/Ui  ( .x(ol[1]), .a(\U2/U589/U25/U1/ob ) );
    oa31_1 \U2/U588/U25/U1/Uclr  ( .x(\U2/U588/U25/U1/clr ), .a(net135), .b(
        \f[3] ), .c(\f[2] ), .d(oh[1]) );
    oaoi211_1 \U2/U588/U25/U1/Uaoi  ( .x(\U2/U588/U25/U1/ob ), .a(\f[3] ), .b(
        \f[2] ), .c(n1), .d(\U2/U588/U25/U1/clr ) );
    inv_2 \U2/U588/U25/U1/Ui  ( .x(oh[1]), .a(\U2/U588/U25/U1/ob ) );
    oa31_1 \U2/U591/U25/U1/Uclr  ( .x(\U2/U591/U25/U1/clr ), .a(net135), .b(
        \f[2] ), .c(\f[0] ), .d(ol[0]) );
    oaoi211_1 \U2/U591/U25/U1/Uaoi  ( .x(\U2/U591/U25/U1/ob ), .a(\f[2] ), .b(
        \f[0] ), .c(n1), .d(\U2/U591/U25/U1/clr ) );
    inv_2 \U2/U591/U25/U1/Ui  ( .x(ol[0]), .a(\U2/U591/U25/U1/ob ) );
    ao222_2 \U2/U592/U19/U1/U1  ( .x(nfa), .a(\U2/x ), .b(\U2/y ), .c(\U2/x ), 
        .d(nfa), .e(\U2/y ), .f(nfa) );
    nor3_1 \U1/U594/U7  ( .x(\U1/x ), .a(ol[5]), .b(\U1/reset ), .c(oh[5]) );
    nor3_1 \U1/U593/U7  ( .x(\U1/y ), .a(ol[4]), .b(\U1/reset ), .c(oh[4]) );
    inv_1 \U1/U604/U3  ( .x(\U1/reset ), .a(nbReset) );
    oa31_1 \U1/U590/U25/U1/Uclr  ( .x(\U1/U590/U25/U1/clr ), .a(net135), .b(
        \e[3] ), .c(\e[1] ), .d(oh[4]) );
    oaoi211_1 \U1/U590/U25/U1/Uaoi  ( .x(\U1/U590/U25/U1/ob ), .a(\e[3] ), .b(
        \e[1] ), .c(n1), .d(\U1/U590/U25/U1/clr ) );
    inv_2 \U1/U590/U25/U1/Ui  ( .x(oh[4]), .a(\U1/U590/U25/U1/ob ) );
    oa31_1 \U1/U589/U25/U1/Uclr  ( .x(\U1/U589/U25/U1/clr ), .a(net135), .b(
        \e[1] ), .c(\e[0] ), .d(ol[5]) );
    oaoi211_1 \U1/U589/U25/U1/Uaoi  ( .x(\U1/U589/U25/U1/ob ), .a(\e[1] ), .b(
        \e[0] ), .c(n1), .d(\U1/U589/U25/U1/clr ) );
    inv_2 \U1/U589/U25/U1/Ui  ( .x(ol[5]), .a(\U1/U589/U25/U1/ob ) );
    oa31_1 \U1/U588/U25/U1/Uclr  ( .x(\U1/U588/U25/U1/clr ), .a(net135), .b(
        \e[3] ), .c(\e[2] ), .d(oh[5]) );
    oaoi211_1 \U1/U588/U25/U1/Uaoi  ( .x(\U1/U588/U25/U1/ob ), .a(\e[3] ), .b(
        \e[2] ), .c(n1), .d(\U1/U588/U25/U1/clr ) );
    inv_2 \U1/U588/U25/U1/Ui  ( .x(oh[5]), .a(\U1/U588/U25/U1/ob ) );
    oa31_1 \U1/U591/U25/U1/Uclr  ( .x(\U1/U591/U25/U1/clr ), .a(net135), .b(
        \e[2] ), .c(\e[0] ), .d(ol[4]) );
    oaoi211_1 \U1/U591/U25/U1/Uaoi  ( .x(\U1/U591/U25/U1/ob ), .a(\e[2] ), .b(
        \e[0] ), .c(n1), .d(\U1/U591/U25/U1/clr ) );
    inv_2 \U1/U591/U25/U1/Ui  ( .x(ol[4]), .a(\U1/U591/U25/U1/ob ) );
    ao222_2 \U1/U592/U19/U1/U1  ( .x(nea), .a(\U1/x ), .b(\U1/y ), .c(\U1/x ), 
        .d(nea), .e(\U1/y ), .f(nea) );
    and3_4 \U881/U20/U9  ( .x(nca), .a(\U881/nack[1] ), .b(\U881/nack[0] ), 
        .c(nbReset) );
    nor2_1 \U881/U18/U5  ( .x(\U881/nack[0] ), .a(\cl[3] ), .b(\cl[0] ) );
    nor2_1 \U881/U19/U5  ( .x(\U881/nack[1] ), .a(\cl[1] ), .b(\cl[2] ) );
    ao222_2 \U881/U15_0_/U19/U1/U1  ( .x(\cl[0] ), .a(\c[0] ), .b(ncla), .c(
        \c[0] ), .d(\cl[0] ), .e(ncla), .f(\cl[0] ) );
    ao222_2 \U881/U15_1_/U19/U1/U1  ( .x(\cl[1] ), .a(\c[1] ), .b(ncla), .c(
        \c[1] ), .d(\cl[1] ), .e(ncla), .f(\cl[1] ) );
    ao222_2 \U881/U15_2_/U19/U1/U1  ( .x(\cl[2] ), .a(\c[2] ), .b(ncla), .c(
        \c[2] ), .d(\cl[2] ), .e(ncla), .f(\cl[2] ) );
    ao222_2 \U881/U15_3_/U19/U1/U1  ( .x(\cl[3] ), .a(\c[3] ), .b(ncla), .c(
        \c[3] ), .d(\cl[3] ), .e(ncla), .f(\cl[3] ) );
    and2_5 U1 ( .x(n1), .a(nbReset), .b(noa) );
    and2_3 U2 ( .x(net135), .a(nbReset), .b(noa) );
endmodule


module chain_selement_ga_69 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_68 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_t_ctrl_0 ( cack, fcdefer, fcslowack, screq, ack, defer, fcack, 
    nReset, scack, slowack );
input  ack, defer, fcack, nReset, scack, slowack;
output cack, fcdefer, fcslowack, screq;
    wire net269, net280, net275, net270, net268, net266, net274, net273, 
        net267, net264, net272, net271, net263, net277, net265, net278, net276, 
        net279, \U49/U28/U1/clr , \U49/U28/U1/set , \U50/U28/U1/clr , 
        \U50/U28/U1/set , \U51/U28/U1/clr , \U51/U28/U1/set , \U57/acb , 
        \U57/U1/Z ;
    chain_selement_ga_69 U55 ( .Aa(net269), .Br(fcdefer), .Ar(net280), .Ba(
        fcack) );
    chain_selement_ga_68 U54 ( .Aa(net275), .Br(fcslowack), .Ar(net270), .Ba(
        fcack) );
    or2_4 \U12/U12  ( .x(net268), .a(net266), .b(net270) );
    or2_4 \U56/U12  ( .x(net274), .a(net275), .b(net269) );
    or2_4 \U14/U12  ( .x(net273), .a(net274), .b(net266) );
    or3_1 \U36/U12  ( .x(cack), .a(net267), .b(net264), .c(net272) );
    nor3_1 \U21/U7  ( .x(net271), .a(net270), .b(net266), .c(net280) );
    and2_1 \U53/U8  ( .x(net263), .a(net271), .b(nReset) );
    and2_1 \U43/U8  ( .x(net277), .a(net265), .b(nReset) );
    nor2_1 \U22/U5  ( .x(net265), .a(net278), .b(net276) );
    ao222_2 \U44/U19/U1/U1  ( .x(net276), .a(net280), .b(net273), .c(net280), 
        .d(net276), .e(net273), .f(net276) );
    ao222_2 \U40/U19/U1/U1  ( .x(net280), .a(net272), .b(net277), .c(net272), 
        .d(net280), .e(net277), .f(net280) );
    ao222_2 \U45/U19/U1/U1  ( .x(net279), .a(net273), .b(net268), .c(net273), 
        .d(net279), .e(net268), .f(net279) );
    ao222_2 \U42/U19/U1/U1  ( .x(net266), .a(net277), .b(net267), .c(net277), 
        .d(net266), .e(net267), .f(net266) );
    ao222_2 \U39/U19/U1/U1  ( .x(net270), .a(net277), .b(net264), .c(net277), 
        .d(net270), .e(net264), .f(net270) );
    aoai211_1 \U49/U28/U1/U1  ( .x(\U49/U28/U1/clr ), .a(ack), .b(nReset), .c(
        net263), .d(net267) );
    nand3_1 \U49/U28/U1/U2  ( .x(\U49/U28/U1/set ), .a(net263), .b(ack), .c(
        nReset) );
    nand2_2 \U49/U28/U1/U3  ( .x(net267), .a(\U49/U28/U1/clr ), .b(
        \U49/U28/U1/set ) );
    aoai211_1 \U50/U28/U1/U1  ( .x(\U50/U28/U1/clr ), .a(slowack), .b(nReset), 
        .c(net263), .d(net264) );
    nand3_1 \U50/U28/U1/U2  ( .x(\U50/U28/U1/set ), .a(net263), .b(slowack), 
        .c(nReset) );
    nand2_2 \U50/U28/U1/U3  ( .x(net264), .a(\U50/U28/U1/clr ), .b(
        \U50/U28/U1/set ) );
    aoai211_1 \U51/U28/U1/U1  ( .x(\U51/U28/U1/clr ), .a(defer), .b(nReset), 
        .c(net263), .d(net272) );
    nand2_2 \U51/U28/U1/U3  ( .x(net272), .a(\U51/U28/U1/clr ), .b(
        \U51/U28/U1/set ) );
    and2_1 \U57/U2/U8  ( .x(screq), .a(net279), .b(\U57/acb ) );
    nor2_1 \U57/U3/U5  ( .x(net278), .a(\U57/acb ), .b(scack) );
    oai21_1 \U57/U1/U30/U1/U1  ( .x(\U57/acb ), .a(\U57/U1/Z ), .b(scack), .c(
        net279) );
    inv_1 \U57/U1/U30/U1/U2  ( .x(\U57/U1/Z ), .a(\U57/acb ) );
    nand3_0 U1 ( .x(\U51/U28/U1/set ), .a(net263), .b(defer), .c(nReset) );
endmodule


module target_wb ( addr, ccol, chainresponse, crnw, csize, ctag, lock, 
    nchaincommandack, nrouteack, pred, rack, routetxreq, seq, tag_h, tag_l, wd, 
    cack, cdefer, chaincommand, cndefer, cok, err, nReset, nchainresponseack, 
    rd, route, routetxack );
output [63:0] addr;
output [5:0] ccol;
output [4:0] chainresponse;
output [1:0] crnw;
output [3:0] csize;
output [9:0] ctag;
output [1:0] lock;
output [1:0] pred;
output [1:0] seq;
output [4:0] tag_h;
output [4:0] tag_l;
output [63:0] wd;
input  [4:0] chaincommand;
input  [1:0] err;
input  [63:0] rd;
input  [4:0] route;
input  cack, cdefer, cndefer, cok, nReset, nchainresponseack, routetxack;
output nchaincommandack, nrouteack, rack, routetxreq;
    wire read_ctrlack, chainff_ack, read_req, \chainff_l[7] , \chainff_l[6] , 
        \chainff_l[5] , \chainff_l[4] , \chainff_l[3] , \chainff_l[2] , 
        \chainff_l[1] , \chainff_l[0] , \chainff_h[7] , \chainff_h[6] , 
        \chainff_h[5] , \chainff_h[4] , \chainff_h[3] , \chainff_h[2] , 
        \chainff_h[1] , \chainff_h[0] , read_cd, teop, rhdrack, fcack, tcba, 
        net145, n7, screq, fcslowack, fcdefer, read_ack, \rhdr_h[7] , 
        \rhdr_l[7] , \rhdr_l[6] , \rhdr_l[5] , \rhdr_h[6] , \rhdr_h[5] , 
        \rhdr_l[15] , \rhdr_l[14] , \rhdr_l[13] , \rhdr_h[15] , \rhdr_h[14] , 
        \rhdr_h[13] , \tcbl[7] , \tcbl[6] , \tcbl[5] , \tcbl[4] , \tcbl[3] , 
        \tcbl[2] , \tcbl[1] , \tcbl[0] , \tcbh[7] , \tcbh[6] , \tcbh[5] , 
        \tcbh[4] , \tcbh[3] , \tcbh[2] , \tcbh[1] , \tcbh[0] , nbreset, 
        ntresponseack, \tresponse[4] , \tresponse[3] , \tresponse[2] , 
        \tresponse[1] , \tresponse[0] , net200, noba, pullcd, net168, n11, n12, 
        net188, net201, net194, net178, net189, net191, \obl[7] , \obl[6] , 
        \obl[5] , \obl[4] , \obl[3] , \obl[2] , \obl[1] , \obl[0] , \obh[7] , 
        \obh[6] , \obh[5] , \obh[4] , \obh[3] , \obh[2] , \obh[1] , \obh[0] , 
        n14, n15, n13, net284, net265, \chdrack[0] , \U1761/y[0] , 
        \U1761/y[1] , chdrctrlack, hdrcd, \U1761/x[3] , \nchdr_ack[7] , 
        \nchdr_ack[6] , \U1761/U28/Z , \U1761/x[0] , \nchdr_ack[1] , 
        \nchdr_ack[0] , \U1761/U32/Z , \U1761/x[2] , \nchdr_ack[5] , 
        \nchdr_ack[4] , \U1761/U29/Z , \U1761/x[1] , \U1761/U33/Z , 
        \U1761/U30/Z , \nchdr_ack[3] , \nchdr_ack[2] , \U1761/U31/Z , 
        \U1632/Z , \chdrack[1] , \U1676/Z , \U1770/U21/nr , \nchdr_ack[10] , 
        \nchdr_ack[9] , \nchdr_ack[8] , \U1770/U21/nd , \U1770/U21/n2 , 
        \net242[10] , \net244[10] , \net243[10] , \net242[9] , \net244[9] , 
        \net243[9] , \net242[8] , \net244[8] , \net243[8] , \net242[7] , 
        \net244[7] , \net243[7] , \net242[6] , \net244[6] , \net243[6] , 
        \net242[5] , \net244[5] , \net243[5] , \net242[4] , \net244[4] , 
        \net243[4] , \net242[3] , \net244[3] , \net243[3] , \net242[2] , 
        \net244[2] , \net243[2] , \net242[1] , \net244[1] , \net243[1] , 
        \net242[0] , \net244[0] , \net243[0] , \U1574_0_/net231 , n10, n9, 
        \U1574_1_/net231 , n8, \U1574_2_/net231 , \U1574_3_/net231 , 
        \U1574_4_/net231 , \U1574_5_/net231 , \U1574_6_/net231 , 
        \U1574_7_/net231 , \U1574_8_/net231 , \U1574_9_/net231 , 
        \U1574_10_/net231 , n4, net248;
    chain_sendword_0 U1765 ( .ctrlack(read_ctrlack), .oh({\chainff_h[7] , 
        \chainff_h[6] , \chainff_h[5] , \chainff_h[4] , \chainff_h[3] , 
        \chainff_h[2] , \chainff_h[1] , \chainff_h[0] }), .ol({\chainff_l[7] , 
        \chainff_l[6] , \chainff_l[5] , \chainff_l[4] , \chainff_l[3] , 
        \chainff_l[2] , \chainff_l[1] , \chainff_l[0] }), .chainackff(
        chainff_ack), .ctrlreq(read_req), .ih(rd[63:32]), .il(rd[31:0]) );
    chain_dr32bit_completion_8 rd_cd ( .o(read_cd), .i(rd) );
    chain_trhdr_0 xmitHdr ( .chainff_ack(chainff_ack), .chainh({\tcbh[7] , 
        \tcbh[6] , \tcbh[5] , \tcbh[4] , \tcbh[3] , \tcbh[2] , \tcbh[1] , 
        \tcbh[0] }), .chainl({\tcbl[7] , \tcbl[6] , \tcbl[5] , \tcbl[4] , 
        \tcbl[3] , \tcbl[2] , \tcbl[1] , \tcbl[0] }), .eop(teop), .hdrack(
        rhdrack), .normal_ack(rack), .notify_ack(fcack), .read_req(read_req), 
        .routereq(routetxreq), .chain_ff_h({\chainff_h[7] , \chainff_h[6] , 
        \chainff_h[5] , \chainff_h[4] , \chainff_h[3] , \chainff_h[2] , 
        \chainff_h[1] , \chainff_h[0] }), .chainack(tcba), .chainff_l({
        \chainff_l[7] , \chainff_l[6] , \chainff_l[5] , \chainff_l[4] , 
        \chainff_l[3] , \chainff_l[2] , \chainff_l[1] , \chainff_l[0] }), 
        .eopack(net145), .err(err), .nReset(n7), .normal_response(screq), 
        .notify_accept(fcslowack), .notify_defer(fcdefer), .rcol_h({
        \rhdr_h[15] , \rhdr_h[14] , \rhdr_h[13] }), .rcol_l({\rhdr_l[15] , 
        \rhdr_l[14] , \rhdr_l[13] }), .read_ack(read_ack), .rnw_h(\rhdr_h[7] ), 
        .rnw_l(\rhdr_l[7] ), .routeack(routetxack), .rsize_h({\rhdr_h[6] , 
        \rhdr_h[5] }), .rsize_l({\rhdr_l[6] , \rhdr_l[5] }), .rtag_h(tag_h), 
        .rtag_l(tag_l) );
    chain_dr2fr_byte_3 dr2fr ( .eop_ack(net145), .ia(tcba), .o({\tresponse[4] , 
        \tresponse[3] , \tresponse[2] , \tresponse[1] , \tresponse[0] }), 
        .eop(teop), .ih({\tcbh[7] , \tcbh[6] , \tcbh[5] , \tcbh[4] , \tcbh[3] , 
        \tcbh[2] , \tcbh[1] , \tcbh[0] }), .il({\tcbl[7] , \tcbl[6] , 
        \tcbl[5] , \tcbl[4] , \tcbl[3] , \tcbl[2] , \tcbl[1] , \tcbl[0] }), 
        .nReset(nbreset), .noa(ntresponseack) );
    chain_mergepackets_3 merger ( .naa(nrouteack), .nba(ntresponseack), .o(
        chainresponse), .a(route), .b({\tresponse[4] , \tresponse[3] , 
        \tresponse[2] , \tresponse[1] , \tresponse[0] }), .nReset(nbreset), 
        .noa(nchainresponseack) );
    chain_tchdr_0 header ( .addr_req(net200), .col_h(ccol[5:3]), .col_l(ccol
        [2:0]), .itag_h(ctag[9:5]), .itag_l(ctag[4:0]), .lock(lock), .ncback(
        noba), .pred(pred), .pullcd(pullcd), .reset(net168), .rnw_h(n11), 
        .rnw_l(n12), .seq(seq), .size_h({n13, csize[2]}), .size_l({n14, n15}), 
        .write_req(net188), .chwh({\obh[7] , \obh[6] , \obh[5] , \obh[4] , 
        \obh[3] , \obh[2] , \obh[1] , \obh[0] }), .chwl({\obl[7] , \obl[6] , 
        \obl[5] , \obl[4] , \obl[3] , \obl[2] , \obl[1] , \obl[0] }), 
        .addr_ack(net201), .addr_pull(net194), .nReset(n7), .nack(net178), 
        .write_ack(net189), .write_pull(net191) );
    chain_irdemux_32new_1 wd_hld ( .ctrlack(net189), .oh(wd[63:32]), .ol(wd
        [31:0]), .pullreq(net191), .pull_h({\obh[7] , \obh[6] , \obh[5] , 
        \obh[4] , \obh[3] , \obh[2] , \obh[1] , \obh[0] }), .pull_l({\obl[7] , 
        \obl[6] , \obl[5] , \obl[4] , \obl[3] , \obl[2] , \obl[1] , \obl[0] }), 
        .pullcd(pullcd), .reset(net168), .ctrlreq(net188) );
    chain_irdemux_32new_0 adr_hld ( .ctrlack(net201), .oh(addr[63:32]), .ol(
        addr[31:0]), .pullreq(net194), .pull_h({\obh[7] , \obh[6] , \obh[5] , 
        \obh[4] , \obh[3] , \obh[2] , \obh[1] , \obh[0] }), .pull_l({\obl[7] , 
        \obl[6] , \obl[5] , \obl[4] , \obl[3] , \obl[2] , \obl[1] , \obl[0] }), 
        .pullcd(pullcd), .reset(net168), .ctrlreq(net200) );
    chain_fr2dr_byte_0 chain_decoder ( .nia(nchaincommandack), .oh({\obh[7] , 
        \obh[6] , \obh[5] , \obh[4] , \obh[3] , \obh[2] , \obh[1] , \obh[0] }), 
        .ol({\obl[7] , \obl[6] , \obl[5] , \obl[4] , \obl[3] , \obl[2] , 
        \obl[1] , \obl[0] }), .i(chaincommand), .nReset(nbreset), .noa(noba)
         );
    chain_t_ctrl_0 cmd_ctrl ( .cack(net284), .fcdefer(fcdefer), .fcslowack(
        fcslowack), .screq(screq), .ack(cok), .defer(cdefer), .fcack(fcack), 
        .nReset(n7), .scack(rack), .slowack(cndefer) );
    inv_1 \I4/U3  ( .x(net265), .a(nbreset) );
    ao222_1 \U1761/U37/U18/U1/U1  ( .x(\chdrack[0] ), .a(\U1761/y[0] ), .b(
        \U1761/y[1] ), .c(\U1761/y[0] ), .d(\chdrack[0] ), .e(\U1761/y[1] ), 
        .f(\chdrack[0] ) );
    ao222_1 \U1762/U18/U1/U1  ( .x(chdrctrlack), .a(hdrcd), .b(net284), .c(
        hdrcd), .d(chdrctrlack), .e(net284), .f(chdrctrlack) );
    ao222_1 \U1769/U18/U1/U1  ( .x(read_ack), .a(read_ctrlack), .b(read_cd), 
        .c(read_ctrlack), .d(read_ack), .e(read_cd), .f(read_ack) );
    aoi222_1 \U1761/U28/U30/U1  ( .x(\U1761/x[3] ), .a(\nchdr_ack[7] ), .b(
        \nchdr_ack[6] ), .c(\nchdr_ack[7] ), .d(\U1761/U28/Z ), .e(
        \nchdr_ack[6] ), .f(\U1761/U28/Z ) );
    inv_1 \U1761/U28/U30/Uinv  ( .x(\U1761/U28/Z ), .a(\U1761/x[3] ) );
    aoi222_1 \U1761/U32/U30/U1  ( .x(\U1761/x[0] ), .a(\nchdr_ack[1] ), .b(
        \nchdr_ack[0] ), .c(\nchdr_ack[1] ), .d(\U1761/U32/Z ), .e(
        \nchdr_ack[0] ), .f(\U1761/U32/Z ) );
    inv_1 \U1761/U32/U30/Uinv  ( .x(\U1761/U32/Z ), .a(\U1761/x[0] ) );
    aoi222_1 \U1761/U29/U30/U1  ( .x(\U1761/x[2] ), .a(\nchdr_ack[5] ), .b(
        \nchdr_ack[4] ), .c(\nchdr_ack[5] ), .d(\U1761/U29/Z ), .e(
        \nchdr_ack[4] ), .f(\U1761/U29/Z ) );
    inv_1 \U1761/U29/U30/Uinv  ( .x(\U1761/U29/Z ), .a(\U1761/x[2] ) );
    aoi222_1 \U1761/U33/U30/U1  ( .x(\U1761/y[0] ), .a(\U1761/x[1] ), .b(
        \U1761/x[0] ), .c(\U1761/x[1] ), .d(\U1761/U33/Z ), .e(\U1761/x[0] ), 
        .f(\U1761/U33/Z ) );
    inv_1 \U1761/U33/U30/Uinv  ( .x(\U1761/U33/Z ), .a(\U1761/y[0] ) );
    aoi222_1 \U1761/U30/U30/U1  ( .x(\U1761/y[1] ), .a(\U1761/x[3] ), .b(
        \U1761/x[2] ), .c(\U1761/x[3] ), .d(\U1761/U30/Z ), .e(\U1761/x[2] ), 
        .f(\U1761/U30/Z ) );
    inv_1 \U1761/U30/U30/Uinv  ( .x(\U1761/U30/Z ), .a(\U1761/y[1] ) );
    aoi222_1 \U1761/U31/U30/U1  ( .x(\U1761/x[1] ), .a(\nchdr_ack[3] ), .b(
        \nchdr_ack[2] ), .c(\nchdr_ack[3] ), .d(\U1761/U31/Z ), .e(
        \nchdr_ack[2] ), .f(\U1761/U31/Z ) );
    inv_1 \U1761/U31/U30/Uinv  ( .x(\U1761/U31/Z ), .a(\U1761/x[1] ) );
    aoi222_1 \U1632/U30/U1  ( .x(net178), .a(cack), .b(chdrctrlack), .c(cack), 
        .d(\U1632/Z ), .e(chdrctrlack), .f(\U1632/Z ) );
    inv_1 \U1632/U30/Uinv  ( .x(\U1632/Z ), .a(net178) );
    aoi222_1 \U1676/U30/U1  ( .x(hdrcd), .a(\chdrack[0] ), .b(\chdrack[1] ), 
        .c(\chdrack[0] ), .d(\U1676/Z ), .e(\chdrack[1] ), .f(\U1676/Z ) );
    inv_1 \U1676/U30/Uinv  ( .x(\U1676/Z ), .a(hdrcd) );
    nor3_1 \U1770/U21/Unr  ( .x(\U1770/U21/nr ), .a(\nchdr_ack[10] ), .b(
        \nchdr_ack[9] ), .c(\nchdr_ack[8] ) );
    nand3_1 \U1770/U21/Und  ( .x(\U1770/U21/nd ), .a(\nchdr_ack[10] ), .b(
        \nchdr_ack[9] ), .c(\nchdr_ack[8] ) );
    oa21_1 \U1770/U21/U1  ( .x(\U1770/U21/n2 ), .a(\U1770/U21/n2 ), .b(
        \U1770/U21/nr ), .c(\U1770/U21/nd ) );
    inv_1 \U1770/U21/U3  ( .x(\chdrack[1] ), .a(\U1770/U21/n2 ) );
    nor2_1 \U1652_0_/U2/U5  ( .x(\nchdr_ack[0] ), .a(\net242[10] ), .b(
        \net244[10] ) );
    ao222_2 \U1652_0_/U12/U19/U1/U1  ( .x(\net244[10] ), .a(\net243[10] ), .b(
        csize[0]), .c(\net243[10] ), .d(\net244[10] ), .e(csize[0]), .f(
        \net244[10] ) );
    ao222_2 \U1652_0_/U11/U19/U1/U1  ( .x(\net242[10] ), .a(csize[2]), .b(
        \net243[10] ), .c(csize[2]), .d(\net242[10] ), .e(\net243[10] ), .f(
        \net242[10] ) );
    nor2_1 \U1652_1_/U2/U5  ( .x(\nchdr_ack[1] ), .a(\net242[9] ), .b(
        \net244[9] ) );
    ao222_2 \U1652_1_/U12/U19/U1/U1  ( .x(\net244[9] ), .a(\net243[9] ), .b(
        csize[1]), .c(\net243[9] ), .d(\net244[9] ), .e(csize[1]), .f(
        \net244[9] ) );
    ao222_2 \U1652_1_/U11/U19/U1/U1  ( .x(\net242[9] ), .a(csize[3]), .b(
        \net243[9] ), .c(csize[3]), .d(\net242[9] ), .e(\net243[9] ), .f(
        \net242[9] ) );
    nor2_1 \U1652_2_/U2/U5  ( .x(\nchdr_ack[2] ), .a(\net242[8] ), .b(
        \net244[8] ) );
    ao222_2 \U1652_2_/U12/U19/U1/U1  ( .x(\net244[8] ), .a(\net243[8] ), .b(
        crnw[0]), .c(\net243[8] ), .d(\net244[8] ), .e(crnw[0]), .f(
        \net244[8] ) );
    ao222_2 \U1652_2_/U11/U19/U1/U1  ( .x(\net242[8] ), .a(crnw[1]), .b(
        \net243[8] ), .c(crnw[1]), .d(\net242[8] ), .e(\net243[8] ), .f(
        \net242[8] ) );
    nor2_1 \U1652_3_/U2/U5  ( .x(\nchdr_ack[3] ), .a(\net242[7] ), .b(
        \net244[7] ) );
    ao222_2 \U1652_3_/U12/U19/U1/U1  ( .x(\net244[7] ), .a(\net243[7] ), .b(
        ctag[0]), .c(\net243[7] ), .d(\net244[7] ), .e(ctag[0]), .f(
        \net244[7] ) );
    ao222_2 \U1652_3_/U11/U19/U1/U1  ( .x(\net242[7] ), .a(ctag[5]), .b(
        \net243[7] ), .c(ctag[5]), .d(\net242[7] ), .e(\net243[7] ), .f(
        \net242[7] ) );
    nor2_1 \U1652_4_/U2/U5  ( .x(\nchdr_ack[4] ), .a(\net242[6] ), .b(
        \net244[6] ) );
    ao222_2 \U1652_4_/U12/U19/U1/U1  ( .x(\net244[6] ), .a(\net243[6] ), .b(
        ctag[1]), .c(\net243[6] ), .d(\net244[6] ), .e(ctag[1]), .f(
        \net244[6] ) );
    ao222_2 \U1652_4_/U11/U19/U1/U1  ( .x(\net242[6] ), .a(ctag[6]), .b(
        \net243[6] ), .c(ctag[6]), .d(\net242[6] ), .e(\net243[6] ), .f(
        \net242[6] ) );
    nor2_1 \U1652_5_/U2/U5  ( .x(\nchdr_ack[5] ), .a(\net242[5] ), .b(
        \net244[5] ) );
    ao222_2 \U1652_5_/U12/U19/U1/U1  ( .x(\net244[5] ), .a(\net243[5] ), .b(
        ctag[2]), .c(\net243[5] ), .d(\net244[5] ), .e(ctag[2]), .f(
        \net244[5] ) );
    ao222_2 \U1652_5_/U11/U19/U1/U1  ( .x(\net242[5] ), .a(ctag[7]), .b(
        \net243[5] ), .c(ctag[7]), .d(\net242[5] ), .e(\net243[5] ), .f(
        \net242[5] ) );
    nor2_1 \U1652_6_/U2/U5  ( .x(\nchdr_ack[6] ), .a(\net242[4] ), .b(
        \net244[4] ) );
    ao222_2 \U1652_6_/U12/U19/U1/U1  ( .x(\net244[4] ), .a(\net243[4] ), .b(
        ctag[3]), .c(\net243[4] ), .d(\net244[4] ), .e(ctag[3]), .f(
        \net244[4] ) );
    ao222_2 \U1652_6_/U11/U19/U1/U1  ( .x(\net242[4] ), .a(ctag[8]), .b(
        \net243[4] ), .c(ctag[8]), .d(\net242[4] ), .e(\net243[4] ), .f(
        \net242[4] ) );
    nor2_1 \U1652_7_/U2/U5  ( .x(\nchdr_ack[7] ), .a(\net242[3] ), .b(
        \net244[3] ) );
    ao222_2 \U1652_7_/U12/U19/U1/U1  ( .x(\net244[3] ), .a(\net243[3] ), .b(
        ctag[4]), .c(\net243[3] ), .d(\net244[3] ), .e(ctag[4]), .f(
        \net244[3] ) );
    ao222_2 \U1652_7_/U11/U19/U1/U1  ( .x(\net242[3] ), .a(ctag[9]), .b(
        \net243[3] ), .c(ctag[9]), .d(\net242[3] ), .e(\net243[3] ), .f(
        \net242[3] ) );
    nor2_1 \U1652_8_/U2/U5  ( .x(\nchdr_ack[8] ), .a(\net242[2] ), .b(
        \net244[2] ) );
    ao222_2 \U1652_8_/U12/U19/U1/U1  ( .x(\net244[2] ), .a(\net243[2] ), .b(
        ccol[0]), .c(\net243[2] ), .d(\net244[2] ), .e(ccol[0]), .f(
        \net244[2] ) );
    ao222_2 \U1652_8_/U11/U19/U1/U1  ( .x(\net242[2] ), .a(ccol[3]), .b(
        \net243[2] ), .c(ccol[3]), .d(\net242[2] ), .e(\net243[2] ), .f(
        \net242[2] ) );
    nor2_1 \U1652_9_/U2/U5  ( .x(\nchdr_ack[9] ), .a(\net242[1] ), .b(
        \net244[1] ) );
    ao222_2 \U1652_9_/U12/U19/U1/U1  ( .x(\net244[1] ), .a(\net243[1] ), .b(
        ccol[1]), .c(\net243[1] ), .d(\net244[1] ), .e(ccol[1]), .f(
        \net244[1] ) );
    ao222_2 \U1652_9_/U11/U19/U1/U1  ( .x(\net242[1] ), .a(ccol[4]), .b(
        \net243[1] ), .c(ccol[4]), .d(\net242[1] ), .e(\net243[1] ), .f(
        \net242[1] ) );
    nor2_1 \U1652_10_/U2/U5  ( .x(\nchdr_ack[10] ), .a(\net242[0] ), .b(
        \net244[0] ) );
    ao222_2 \U1652_10_/U12/U19/U1/U1  ( .x(\net244[0] ), .a(\net243[0] ), .b(
        ccol[2]), .c(\net243[0] ), .d(\net244[0] ), .e(ccol[2]), .f(
        \net244[0] ) );
    ao222_2 \U1652_10_/U11/U19/U1/U1  ( .x(\net242[0] ), .a(ccol[5]), .b(
        \net243[0] ), .c(ccol[5]), .d(\net242[0] ), .e(\net243[0] ), .f(
        \net242[0] ) );
    nor2_1 \U1574_0_/U2/U5  ( .x(\U1574_0_/net231 ), .a(\rhdr_l[5] ), .b(
        \rhdr_h[5] ) );
    and2_1 \U1574_0_/U13/U8  ( .x(\net243[10] ), .a(\U1574_0_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_0_/U12/U19/U1/U1  ( .x(\rhdr_h[5] ), .a(n10), .b(
        \net242[10] ), .c(n10), .d(\rhdr_h[5] ), .e(\net242[10] ), .f(
        \rhdr_h[5] ) );
    ao222_2 \U1574_0_/U11/U19/U1/U1  ( .x(\rhdr_l[5] ), .a(\net244[10] ), .b(
        n9), .c(\net244[10] ), .d(\rhdr_l[5] ), .e(n10), .f(\rhdr_l[5] ) );
    nor2_1 \U1574_1_/U2/U5  ( .x(\U1574_1_/net231 ), .a(\rhdr_l[6] ), .b(
        \rhdr_h[6] ) );
    and2_1 \U1574_1_/U13/U8  ( .x(\net243[9] ), .a(\U1574_1_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_1_/U12/U19/U1/U1  ( .x(\rhdr_h[6] ), .a(n9), .b(\net242[9] 
        ), .c(n8), .d(\rhdr_h[6] ), .e(\net242[9] ), .f(\rhdr_h[6] ) );
    ao222_2 \U1574_1_/U11/U19/U1/U1  ( .x(\rhdr_l[6] ), .a(\net244[9] ), .b(n9
        ), .c(\net244[9] ), .d(\rhdr_l[6] ), .e(n10), .f(\rhdr_l[6] ) );
    nor2_1 \U1574_2_/U2/U5  ( .x(\U1574_2_/net231 ), .a(\rhdr_l[7] ), .b(
        \rhdr_h[7] ) );
    and2_1 \U1574_2_/U13/U8  ( .x(\net243[8] ), .a(\U1574_2_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_2_/U12/U19/U1/U1  ( .x(\rhdr_h[7] ), .a(n8), .b(\net242[8] 
        ), .c(n8), .d(\rhdr_h[7] ), .e(\net242[8] ), .f(\rhdr_h[7] ) );
    ao222_2 \U1574_2_/U11/U19/U1/U1  ( .x(\rhdr_l[7] ), .a(\net244[8] ), .b(n9
        ), .c(\net244[8] ), .d(\rhdr_l[7] ), .e(n10), .f(\rhdr_l[7] ) );
    nor2_1 \U1574_3_/U2/U5  ( .x(\U1574_3_/net231 ), .a(tag_l[0]), .b(tag_h[0]
        ) );
    and2_1 \U1574_3_/U13/U8  ( .x(\net243[7] ), .a(\U1574_3_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_3_/U12/U19/U1/U1  ( .x(tag_h[0]), .a(n10), .b(\net242[7] ), 
        .c(n8), .d(tag_h[0]), .e(\net242[7] ), .f(tag_h[0]) );
    ao222_2 \U1574_3_/U11/U19/U1/U1  ( .x(tag_l[0]), .a(\net244[7] ), .b(n9), 
        .c(\net244[7] ), .d(tag_l[0]), .e(n8), .f(tag_l[0]) );
    nor2_1 \U1574_4_/U2/U5  ( .x(\U1574_4_/net231 ), .a(tag_l[1]), .b(tag_h[1]
        ) );
    and2_1 \U1574_4_/U13/U8  ( .x(\net243[6] ), .a(\U1574_4_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_4_/U12/U19/U1/U1  ( .x(tag_h[1]), .a(n8), .b(\net242[6] ), 
        .c(n8), .d(tag_h[1]), .e(\net242[6] ), .f(tag_h[1]) );
    ao222_2 \U1574_4_/U11/U19/U1/U1  ( .x(tag_l[1]), .a(\net244[6] ), .b(n9), 
        .c(\net244[6] ), .d(tag_l[1]), .e(n8), .f(tag_l[1]) );
    nor2_1 \U1574_5_/U2/U5  ( .x(\U1574_5_/net231 ), .a(tag_l[2]), .b(tag_h[2]
        ) );
    and2_1 \U1574_5_/U13/U8  ( .x(\net243[5] ), .a(\U1574_5_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_5_/U12/U19/U1/U1  ( .x(tag_h[2]), .a(n9), .b(\net242[5] ), 
        .c(n8), .d(tag_h[2]), .e(\net242[5] ), .f(tag_h[2]) );
    ao222_2 \U1574_5_/U11/U19/U1/U1  ( .x(tag_l[2]), .a(\net244[5] ), .b(n9), 
        .c(\net244[5] ), .d(tag_l[2]), .e(n10), .f(tag_l[2]) );
    nor2_1 \U1574_6_/U2/U5  ( .x(\U1574_6_/net231 ), .a(tag_l[3]), .b(tag_h[3]
        ) );
    and2_1 \U1574_6_/U13/U8  ( .x(\net243[4] ), .a(\U1574_6_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_6_/U12/U19/U1/U1  ( .x(tag_h[3]), .a(n8), .b(\net242[4] ), 
        .c(n10), .d(tag_h[3]), .e(\net242[4] ), .f(tag_h[3]) );
    ao222_2 \U1574_6_/U11/U19/U1/U1  ( .x(tag_l[3]), .a(\net244[4] ), .b(n9), 
        .c(\net244[4] ), .d(tag_l[3]), .e(n8), .f(tag_l[3]) );
    nor2_1 \U1574_7_/U2/U5  ( .x(\U1574_7_/net231 ), .a(tag_l[4]), .b(tag_h[4]
        ) );
    and2_1 \U1574_7_/U13/U8  ( .x(\net243[3] ), .a(\U1574_7_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_7_/U12/U19/U1/U1  ( .x(tag_h[4]), .a(n8), .b(\net242[3] ), 
        .c(n10), .d(tag_h[4]), .e(\net242[3] ), .f(tag_h[4]) );
    ao222_2 \U1574_7_/U11/U19/U1/U1  ( .x(tag_l[4]), .a(\net244[3] ), .b(n9), 
        .c(\net244[3] ), .d(tag_l[4]), .e(n8), .f(tag_l[4]) );
    nor2_1 \U1574_8_/U2/U5  ( .x(\U1574_8_/net231 ), .a(\rhdr_l[13] ), .b(
        \rhdr_h[13] ) );
    and2_1 \U1574_8_/U13/U8  ( .x(\net243[2] ), .a(\U1574_8_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_8_/U12/U19/U1/U1  ( .x(\rhdr_h[13] ), .a(n9), .b(
        \net242[2] ), .c(n10), .d(\rhdr_h[13] ), .e(\net242[2] ), .f(
        \rhdr_h[13] ) );
    ao222_2 \U1574_8_/U11/U19/U1/U1  ( .x(\rhdr_l[13] ), .a(\net244[2] ), .b(
        n9), .c(\net244[2] ), .d(\rhdr_l[13] ), .e(n8), .f(\rhdr_l[13] ) );
    nor2_1 \U1574_9_/U2/U5  ( .x(\U1574_9_/net231 ), .a(\rhdr_l[14] ), .b(
        \rhdr_h[14] ) );
    and2_1 \U1574_9_/U13/U8  ( .x(\net243[1] ), .a(\U1574_9_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_9_/U12/U19/U1/U1  ( .x(\rhdr_h[14] ), .a(n10), .b(
        \net242[1] ), .c(n8), .d(\rhdr_h[14] ), .e(\net242[1] ), .f(
        \rhdr_h[14] ) );
    ao222_2 \U1574_9_/U11/U19/U1/U1  ( .x(\rhdr_l[14] ), .a(\net244[1] ), .b(
        n9), .c(\net244[1] ), .d(\rhdr_l[14] ), .e(n10), .f(\rhdr_l[14] ) );
    nor2_1 \U1574_10_/U2/U5  ( .x(\U1574_10_/net231 ), .a(\rhdr_l[15] ), .b(
        \rhdr_h[15] ) );
    and2_1 \U1574_10_/U13/U8  ( .x(\net243[0] ), .a(\U1574_10_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_10_/U12/U19/U1/U1  ( .x(\rhdr_h[15] ), .a(n10), .b(
        \net242[0] ), .c(n10), .d(\rhdr_h[15] ), .e(\net242[0] ), .f(
        \rhdr_h[15] ) );
    ao222_2 \U1574_10_/U11/U19/U1/U1  ( .x(\rhdr_l[15] ), .a(\net244[0] ), .b(
        n9), .c(\net244[0] ), .d(\rhdr_l[15] ), .e(n10), .f(\rhdr_l[15] ) );
    buf_1 U1 ( .x(csize[0]), .a(n15) );
    buf_1 U2 ( .x(csize[1]), .a(n14) );
    buf_1 U3 ( .x(csize[3]), .a(n13) );
    inv_0 U4 ( .x(n4), .a(n12) );
    inv_2 U5 ( .x(crnw[0]), .a(n4) );
    buf_1 U6 ( .x(crnw[1]), .a(n11) );
    inv_5 U7 ( .x(n7), .a(net265) );
    buf_3 U8 ( .x(nbreset), .a(nReset) );
    buf_3 U9 ( .x(n8), .a(net248) );
    buf_3 U10 ( .x(n10), .a(net248) );
    buf_3 U11 ( .x(n9), .a(net248) );
    nor2_1 U12 ( .x(net248), .a(net265), .b(rhdrack) );
endmodule


module t_adec_wb ( e_h, e_l, r_h, r_l, e_dp, e_ip, e_tic, r_dp, r_ip, r_tic, 
    tag_h, tag_l );
output [2:0] e_h;
output [2:0] e_l;
output [2:0] r_h;
output [2:0] r_l;
input  [2:0] e_dp;
input  [2:0] e_ip;
input  [2:0] e_tic;
input  [2:0] r_dp;
input  [2:0] r_ip;
input  [2:0] r_tic;
input  [4:0] tag_h;
input  [4:0] tag_l;
    wire e_h_1, e_h_0, e_l_2, r_h_1;
    assign e_h[2] = 1'b0;
    assign e_h[1] = e_h_1;
    assign e_h[0] = e_h_0;
    assign e_l[2] = e_l_2;
    assign e_l[1] = e_h_0;
    assign e_l[0] = e_h_1;
    assign r_h[2] = e_h_0;
    assign r_h[1] = r_h_1;
    assign r_h[0] = 1'b0;
    assign r_l[2] = e_h_1;
    assign r_l[0] = e_l_2;
    assign r_h_1 = tag_h[4];
    or2_1 U3 ( .x(r_l[1]), .a(e_h_1), .b(tag_h[3]) );
    buf_3 U6 ( .x(e_h_1), .a(tag_h[2]) );
    or2_2 U7 ( .x(e_l_2), .a(r_h_1), .b(r_l[1]) );
    or2_2 U8 ( .x(e_h_0), .a(tag_h[3]), .b(r_h_1) );
endmodule


module chain_selement_ga_74 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_2 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_symbol_13 ( o, txack, txack_last, e, oa, r, txreq );
output [2:0] o;
input  [1:0] e;
input  [1:0] r;
input  oa, txreq;
output txack, txack_last;
    wire ack, net10, \c[0] , \c[1] ;
    chain_selement_ga_2 U1239 ( .Aa(ack), .Br(net10), .Ar(txreq), .Ba(oa) );
    and2_1 \U1229_0_/U8  ( .x(o[0]), .a(\c[0] ), .b(net10) );
    and2_1 \U1229_1_/U8  ( .x(o[1]), .a(\c[1] ), .b(net10) );
    and2_1 \U1229_2_/U8  ( .x(o[2]), .a(e[1]), .b(net10) );
    ao23_1 \U1251/U19/U21/U1/U1  ( .x(txack_last), .a(ack), .b(txack_last), 
        .c(ack), .d(e[1]), .e(e[1]) );
    ao23_1 \U1250/U19/U21/U1/U1  ( .x(txack), .a(ack), .b(txack), .c(ack), .d(
        e[0]), .e(e[0]) );
    ao222_1 \U1210/U18/U1/U1  ( .x(\c[0] ), .a(e[0]), .b(r[0]), .c(e[0]), .d(
        \c[0] ), .e(r[0]), .f(\c[0] ) );
    ao222_1 \U1209/U18/U1/U1  ( .x(\c[1] ), .a(e[0]), .b(r[1]), .c(e[0]), .d(
        \c[1] ), .e(r[1]), .f(\c[1] ) );
endmodule


module chain_selement_ga_3 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_symbol_14 ( o, txack, txack_last, e, oa, r, txreq );
output [2:0] o;
input  [1:0] e;
input  [1:0] r;
input  oa, txreq;
output txack, txack_last;
    wire ack, net10, \c[0] , \c[1] , n2, n1;
    chain_selement_ga_3 U1239 ( .Aa(ack), .Br(net10), .Ar(txreq), .Ba(oa) );
    and2_1 \U1229_0_/U8  ( .x(o[0]), .a(\c[0] ), .b(net10) );
    and2_1 \U1229_1_/U8  ( .x(o[1]), .a(\c[1] ), .b(net10) );
    and2_1 \U1229_2_/U8  ( .x(o[2]), .a(e[1]), .b(net10) );
    ao23_1 \U1251/U19/U21/U1/U1  ( .x(txack_last), .a(ack), .b(txack_last), 
        .c(ack), .d(e[1]), .e(e[1]) );
    ao23_1 \U1250/U19/U21/U1/U1  ( .x(txack), .a(ack), .b(txack), .c(ack), .d(
        n2), .e(n2) );
    ao222_1 \U1210/U18/U1/U1  ( .x(\c[0] ), .a(n2), .b(r[0]), .c(n2), .d(
        \c[0] ), .e(r[0]), .f(\c[0] ) );
    ao222_1 \U1209/U18/U1/U1  ( .x(\c[1] ), .a(n2), .b(r[1]), .c(n2), .d(
        \c[1] ), .e(r[1]), .f(\c[1] ) );
    inv_0 U1 ( .x(n1), .a(e[0]) );
    inv_2 U2 ( .x(n2), .a(n1) );
endmodule


module chain_selement_ga_1 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_symbol_12 ( o, txack, txack_last, e, oa, r, txreq );
output [2:0] o;
input  [1:0] e;
input  [1:0] r;
input  oa, txreq;
output txack, txack_last;
    wire ack, net10, \c[0] , \c[1] ;
    chain_selement_ga_1 U1239 ( .Aa(ack), .Br(net10), .Ar(txreq), .Ba(oa) );
    and2_1 \U1229_0_/U8  ( .x(o[0]), .a(\c[0] ), .b(net10) );
    and2_1 \U1229_1_/U8  ( .x(o[1]), .a(\c[1] ), .b(net10) );
    and2_1 \U1229_2_/U8  ( .x(o[2]), .a(e[1]), .b(net10) );
    ao23_1 \U1251/U19/U21/U1/U1  ( .x(txack_last), .a(ack), .b(txack_last), 
        .c(ack), .d(e[1]), .e(e[1]) );
    ao23_1 \U1250/U19/U21/U1/U1  ( .x(txack), .a(ack), .b(txack), .c(ack), .d(
        e[0]), .e(e[0]) );
    ao222_1 \U1210/U18/U1/U1  ( .x(\c[0] ), .a(e[0]), .b(r[0]), .c(e[0]), .d(
        \c[0] ), .e(r[0]), .f(\c[0] ) );
    ao222_1 \U1209/U18/U1/U1  ( .x(\c[1] ), .a(e[0]), .b(r[1]), .c(e[0]), .d(
        \c[1] ), .e(r[1]), .f(\c[1] ) );
endmodule


module resp_route_tx_wb ( o, rtxack, e_h, e_l, noa, r_h, r_l, rtxreq );
output [4:0] o;
input  [2:0] e_h;
input  [2:0] e_l;
input  [2:0] r_h;
input  [2:0] r_l;
input  noa, rtxreq;
output rtxack;
    wire \last[0] , eopsym, net87, net66, net84, \last[2] , net77, \r1[2] , 
        \r1[1] , \r1[0] , \last[1] , \r0[2] , \r0[1] , \r0[0] , \last[3] , 
        \r2[2] , \r2[1] , \r2[0] , net106, net103, \net72[1] , \net72[0] , 
        \I8/nb , \I8/na , \I11/n5 , \I11/n1 , \I11/n2 , \I11/n3 , \I11/n4 , 
        net56, \I7_0_/U25/U1/clr , \I7_0_/U25/U1/ob , \I7_1_/U25/U1/clr , 
        \I7_1_/U25/U1/ob ;
    assign o[3] = 1'b0;
    assign o[2] = 1'b0;
    chain_selement_ga_74 I9 ( .Aa(\last[0] ), .Br(eopsym), .Ar(net87), .Ba(
        net66) );
    route_symbol_13 I2 ( .o({\r1[2] , \r1[1] , \r1[0] }), .txack(net84), 
        .txack_last(\last[2] ), .e({e_h[1], e_l[1]}), .oa(net66), .r({r_h[1], 
        r_l[1]}), .txreq(net77) );
    route_symbol_14 I3 ( .o({\r0[2] , \r0[1] , \r0[0] }), .txack(net87), 
        .txack_last(\last[1] ), .e({e_h[0], e_l[0]}), .oa(net66), .r({r_h[0], 
        r_l[0]}), .txreq(net84) );
    route_symbol_12 I1 ( .o({\r2[2] , \r2[1] , \r2[0] }), .txack(net77), 
        .txack_last(\last[3] ), .e({e_h[2], e_l[2]}), .oa(net66), .r({r_h[2], 
        r_l[2]}), .txreq(rtxreq) );
    nor2_1 \I5/U5  ( .x(net106), .a(eopsym), .b(\r2[2] ) );
    nor2_1 \I16/U5  ( .x(net103), .a(\r1[2] ), .b(\r0[2] ) );
    or2_1 \I14_0_/U12  ( .x(\net72[1] ), .a(\r2[0] ), .b(\r1[0] ) );
    or2_1 \I14_1_/U12  ( .x(\net72[0] ), .a(\r2[1] ), .b(\r1[1] ) );
    nor3_1 \I8/U27  ( .x(\I8/nb ), .a(o[4]), .b(1'b0), .c(1'b0) );
    nor2_1 \I8/U26  ( .x(\I8/na ), .a(o[1]), .b(o[0]) );
    nand2_2 \I8/U29  ( .x(net66), .a(\I8/nb ), .b(\I8/na ) );
    and4_1 \I11/U16  ( .x(\I11/n5 ), .a(\I11/n1 ), .b(\I11/n2 ), .c(\I11/n3 ), 
        .d(\I11/n4 ) );
    inv_1 \I11/U1  ( .x(\I11/n1 ), .a(\last[3] ) );
    inv_1 \I11/U2  ( .x(\I11/n2 ), .a(\last[2] ) );
    inv_1 \I11/U3  ( .x(\I11/n3 ), .a(\last[1] ) );
    inv_1 \I11/U4  ( .x(\I11/n4 ), .a(\last[0] ) );
    inv_1 \I11/U5  ( .x(rtxack), .a(\I11/n5 ) );
    nand2_1 \I17/U5  ( .x(net56), .a(net106), .b(net103) );
    ao222_1 \I15/U18/U1/U1  ( .x(o[4]), .a(noa), .b(net56), .c(noa), .d(o[4]), 
        .e(net56), .f(o[4]) );
    oa31_1 \I7_0_/U25/U1/Uclr  ( .x(\I7_0_/U25/U1/clr ), .a(noa), .b(\r0[0] ), 
        .c(\net72[1] ), .d(o[0]) );
    oaoi211_1 \I7_0_/U25/U1/Uaoi  ( .x(\I7_0_/U25/U1/ob ), .a(\r0[0] ), .b(
        \net72[1] ), .c(noa), .d(\I7_0_/U25/U1/clr ) );
    inv_2 \I7_0_/U25/U1/Ui  ( .x(o[0]), .a(\I7_0_/U25/U1/ob ) );
    oa31_1 \I7_1_/U25/U1/Uclr  ( .x(\I7_1_/U25/U1/clr ), .a(noa), .b(\r0[1] ), 
        .c(\net72[0] ), .d(o[1]) );
    oaoi211_1 \I7_1_/U25/U1/Uaoi  ( .x(\I7_1_/U25/U1/ob ), .a(\r0[1] ), .b(
        \net72[0] ), .c(noa), .d(\I7_1_/U25/U1/clr ) );
    inv_2 \I7_1_/U25/U1/Ui  ( .x(o[1]), .a(\I7_1_/U25/U1/ob ) );
endmodule


module sr2dr_word_6 ( i, req, h, l );
input  [31:0] i;
output [31:0] h;
output [31:0] l;
input  req;
    wire \U31/ni , \U31/nh , \U31/nl , n9, n1, n2, \U30/ni , \U30/nh , 
        \U30/nl , n8, \U29/ni , \U29/nh , \U29/nl , \U28/ni , \U28/nh , 
        \U28/nl , \U27/ni , \U27/nh , \U27/nl , \U26/ni , \U26/nh , \U26/nl , 
        n7, n4, \U25/ni , \U25/nh , \U25/nl , \U24/ni , \U24/nh , \U24/nl , 
        \U23/ni , \U23/nh , \U23/nl , n3, \U22/ni , \U22/nh , \U22/nl , n6, 
        \U21/ni , \U21/nh , \U21/nl , \U20/ni , \U20/nh , \U20/nl , n5, 
        \U19/ni , \U19/nh , \U19/nl , \U18/ni , \U18/nh , \U18/nl , \U17/ni , 
        \U17/nh , \U17/nl , \U16/ni , \U16/nh , \U16/nl , \U15/ni , \U15/nh , 
        \U15/nl , \U14/ni , \U14/nh , \U14/nl , \U13/ni , \U13/nh , \U13/nl , 
        \U12/ni , \U12/nh , \U12/nl , \U11/ni , \U11/nh , \U11/nl , \U10/ni , 
        \U10/nh , \U10/nl , \U9/ni , \U9/nh , \U9/nl , \U8/ni , \U8/nh , 
        \U8/nl , \U7/ni , \U7/nh , \U7/nl , \U6/ni , \U6/nh , \U6/nl , \U5/ni , 
        \U5/nh , \U5/nl , \U4/ni , \U4/nh , \U4/nl , \U3/ni , \U3/nh , \U3/nl , 
        \U2/ni , \U2/nh , \U2/nl , \U1/ni , \U1/nh , \U1/nl , \U0/ni , \U0/nh , 
        \U0/nl , n12, n11, n10;
    inv_1 \U31/Uii  ( .x(\U31/ni ), .a(i[31]) );
    inv_1 \U31/Uih  ( .x(\U31/nh ), .a(h[31]) );
    inv_1 \U31/Uil  ( .x(\U31/nl ), .a(l[31]) );
    ao23_1 \U31/Ucl/U1/U1  ( .x(l[31]), .a(n9), .b(l[31]), .c(n1), .d(\U31/ni 
        ), .e(\U31/nh ) );
    ao23_1 \U31/Uch/U1/U1  ( .x(h[31]), .a(n9), .b(h[31]), .c(n2), .d(i[31]), 
        .e(\U31/nl ) );
    inv_1 \U30/Uii  ( .x(\U30/ni ), .a(i[30]) );
    inv_1 \U30/Uih  ( .x(\U30/nh ), .a(h[30]) );
    inv_1 \U30/Uil  ( .x(\U30/nl ), .a(l[30]) );
    ao23_1 \U30/Ucl/U1/U1  ( .x(l[30]), .a(n8), .b(l[30]), .c(n1), .d(\U30/ni 
        ), .e(\U30/nh ) );
    ao23_1 \U30/Uch/U1/U1  ( .x(h[30]), .a(n8), .b(h[30]), .c(n1), .d(i[30]), 
        .e(\U30/nl ) );
    inv_1 \U29/Uii  ( .x(\U29/ni ), .a(i[29]) );
    inv_1 \U29/Uih  ( .x(\U29/nh ), .a(h[29]) );
    inv_1 \U29/Uil  ( .x(\U29/nl ), .a(l[29]) );
    ao23_1 \U29/Ucl/U1/U1  ( .x(l[29]), .a(n8), .b(l[29]), .c(n1), .d(\U29/ni 
        ), .e(\U29/nh ) );
    ao23_1 \U29/Uch/U1/U1  ( .x(h[29]), .a(n8), .b(h[29]), .c(n2), .d(i[29]), 
        .e(\U29/nl ) );
    inv_1 \U28/Uii  ( .x(\U28/ni ), .a(i[28]) );
    inv_1 \U28/Uih  ( .x(\U28/nh ), .a(h[28]) );
    inv_1 \U28/Uil  ( .x(\U28/nl ), .a(l[28]) );
    ao23_1 \U28/Ucl/U1/U1  ( .x(l[28]), .a(n8), .b(l[28]), .c(n2), .d(\U28/ni 
        ), .e(\U28/nh ) );
    ao23_1 \U28/Uch/U1/U1  ( .x(h[28]), .a(n8), .b(h[28]), .c(n2), .d(i[28]), 
        .e(\U28/nl ) );
    inv_1 \U27/Uii  ( .x(\U27/ni ), .a(i[27]) );
    inv_1 \U27/Uih  ( .x(\U27/nh ), .a(h[27]) );
    inv_1 \U27/Uil  ( .x(\U27/nl ), .a(l[27]) );
    ao23_1 \U27/Ucl/U1/U1  ( .x(l[27]), .a(n8), .b(l[27]), .c(n2), .d(\U27/ni 
        ), .e(\U27/nh ) );
    ao23_1 \U27/Uch/U1/U1  ( .x(h[27]), .a(n8), .b(h[27]), .c(n2), .d(i[27]), 
        .e(\U27/nl ) );
    inv_1 \U26/Uii  ( .x(\U26/ni ), .a(i[26]) );
    inv_1 \U26/Uih  ( .x(\U26/nh ), .a(h[26]) );
    inv_1 \U26/Uil  ( .x(\U26/nl ), .a(l[26]) );
    ao23_1 \U26/Ucl/U1/U1  ( .x(l[26]), .a(n7), .b(l[26]), .c(n2), .d(\U26/ni 
        ), .e(\U26/nh ) );
    ao23_1 \U26/Uch/U1/U1  ( .x(h[26]), .a(n7), .b(h[26]), .c(n4), .d(i[26]), 
        .e(\U26/nl ) );
    inv_1 \U25/Uii  ( .x(\U25/ni ), .a(i[25]) );
    inv_1 \U25/Uih  ( .x(\U25/nh ), .a(h[25]) );
    inv_1 \U25/Uil  ( .x(\U25/nl ), .a(l[25]) );
    ao23_1 \U25/Ucl/U1/U1  ( .x(l[25]), .a(n7), .b(l[25]), .c(n4), .d(\U25/ni 
        ), .e(\U25/nh ) );
    ao23_1 \U25/Uch/U1/U1  ( .x(h[25]), .a(n7), .b(h[25]), .c(n4), .d(i[25]), 
        .e(\U25/nl ) );
    inv_1 \U24/Uii  ( .x(\U24/ni ), .a(i[24]) );
    inv_1 \U24/Uih  ( .x(\U24/nh ), .a(h[24]) );
    inv_1 \U24/Uil  ( .x(\U24/nl ), .a(l[24]) );
    ao23_1 \U24/Ucl/U1/U1  ( .x(l[24]), .a(n7), .b(l[24]), .c(n4), .d(\U24/ni 
        ), .e(\U24/nh ) );
    ao23_1 \U24/Uch/U1/U1  ( .x(h[24]), .a(n7), .b(h[24]), .c(n4), .d(i[24]), 
        .e(\U24/nl ) );
    inv_1 \U23/Uii  ( .x(\U23/ni ), .a(i[23]) );
    inv_1 \U23/Uih  ( .x(\U23/nh ), .a(h[23]) );
    inv_1 \U23/Uil  ( .x(\U23/nl ), .a(l[23]) );
    ao23_1 \U23/Ucl/U1/U1  ( .x(l[23]), .a(n7), .b(l[23]), .c(n3), .d(\U23/ni 
        ), .e(\U23/nh ) );
    ao23_1 \U23/Uch/U1/U1  ( .x(h[23]), .a(n7), .b(h[23]), .c(n3), .d(i[23]), 
        .e(\U23/nl ) );
    inv_1 \U22/Uii  ( .x(\U22/ni ), .a(i[22]) );
    inv_1 \U22/Uih  ( .x(\U22/nh ), .a(h[22]) );
    inv_1 \U22/Uil  ( .x(\U22/nl ), .a(l[22]) );
    ao23_1 \U22/Ucl/U1/U1  ( .x(l[22]), .a(n6), .b(l[22]), .c(n3), .d(\U22/ni 
        ), .e(\U22/nh ) );
    ao23_1 \U22/Uch/U1/U1  ( .x(h[22]), .a(n6), .b(h[22]), .c(n3), .d(i[22]), 
        .e(\U22/nl ) );
    inv_1 \U21/Uii  ( .x(\U21/ni ), .a(i[21]) );
    inv_1 \U21/Uih  ( .x(\U21/nh ), .a(h[21]) );
    inv_1 \U21/Uil  ( .x(\U21/nl ), .a(l[21]) );
    ao23_1 \U21/Ucl/U1/U1  ( .x(l[21]), .a(n6), .b(l[21]), .c(n3), .d(\U21/ni 
        ), .e(\U21/nh ) );
    ao23_1 \U21/Uch/U1/U1  ( .x(h[21]), .a(n6), .b(h[21]), .c(n3), .d(i[21]), 
        .e(\U21/nl ) );
    inv_1 \U20/Uii  ( .x(\U20/ni ), .a(i[20]) );
    inv_1 \U20/Uih  ( .x(\U20/nh ), .a(h[20]) );
    inv_1 \U20/Uil  ( .x(\U20/nl ), .a(l[20]) );
    ao23_1 \U20/Ucl/U1/U1  ( .x(l[20]), .a(n6), .b(l[20]), .c(n5), .d(\U20/ni 
        ), .e(\U20/nh ) );
    ao23_1 \U20/Uch/U1/U1  ( .x(h[20]), .a(n6), .b(h[20]), .c(n4), .d(i[20]), 
        .e(\U20/nl ) );
    inv_1 \U19/Uii  ( .x(\U19/ni ), .a(i[19]) );
    inv_1 \U19/Uih  ( .x(\U19/nh ), .a(h[19]) );
    inv_1 \U19/Uil  ( .x(\U19/nl ), .a(l[19]) );
    ao23_1 \U19/Ucl/U1/U1  ( .x(l[19]), .a(n6), .b(l[19]), .c(n4), .d(\U19/ni 
        ), .e(\U19/nh ) );
    ao23_1 \U19/Uch/U1/U1  ( .x(h[19]), .a(n6), .b(h[19]), .c(n4), .d(i[19]), 
        .e(\U19/nl ) );
    inv_1 \U18/Uii  ( .x(\U18/ni ), .a(i[18]) );
    inv_1 \U18/Uih  ( .x(\U18/nh ), .a(h[18]) );
    inv_1 \U18/Uil  ( .x(\U18/nl ), .a(l[18]) );
    ao23_1 \U18/Ucl/U1/U1  ( .x(l[18]), .a(n5), .b(l[18]), .c(n5), .d(\U18/ni 
        ), .e(\U18/nh ) );
    ao23_1 \U18/Uch/U1/U1  ( .x(h[18]), .a(n5), .b(h[18]), .c(n5), .d(i[18]), 
        .e(\U18/nl ) );
    inv_1 \U17/Uii  ( .x(\U17/ni ), .a(i[17]) );
    inv_1 \U17/Uih  ( .x(\U17/nh ), .a(h[17]) );
    inv_1 \U17/Uil  ( .x(\U17/nl ), .a(l[17]) );
    ao23_1 \U17/Ucl/U1/U1  ( .x(l[17]), .a(n6), .b(l[17]), .c(n5), .d(\U17/ni 
        ), .e(\U17/nh ) );
    ao23_1 \U17/Uch/U1/U1  ( .x(h[17]), .a(n7), .b(h[17]), .c(n4), .d(i[17]), 
        .e(\U17/nl ) );
    inv_1 \U16/Uii  ( .x(\U16/ni ), .a(i[16]) );
    inv_1 \U16/Uih  ( .x(\U16/nh ), .a(h[16]) );
    inv_1 \U16/Uil  ( .x(\U16/nl ), .a(l[16]) );
    ao23_1 \U16/Ucl/U1/U1  ( .x(l[16]), .a(n9), .b(l[16]), .c(n3), .d(\U16/ni 
        ), .e(\U16/nh ) );
    ao23_1 \U16/Uch/U1/U1  ( .x(h[16]), .a(n9), .b(h[16]), .c(n1), .d(i[16]), 
        .e(\U16/nl ) );
    inv_1 \U15/Uii  ( .x(\U15/ni ), .a(i[15]) );
    inv_1 \U15/Uih  ( .x(\U15/nh ), .a(h[15]) );
    inv_1 \U15/Uil  ( .x(\U15/nl ), .a(l[15]) );
    ao23_1 \U15/Ucl/U1/U1  ( .x(l[15]), .a(n8), .b(l[15]), .c(n1), .d(\U15/ni 
        ), .e(\U15/nh ) );
    ao23_1 \U15/Uch/U1/U1  ( .x(h[15]), .a(n7), .b(h[15]), .c(n1), .d(i[15]), 
        .e(\U15/nl ) );
    inv_1 \U14/Uii  ( .x(\U14/ni ), .a(i[14]) );
    inv_1 \U14/Uih  ( .x(\U14/nh ), .a(h[14]) );
    inv_1 \U14/Uil  ( .x(\U14/nl ), .a(l[14]) );
    ao23_1 \U14/Ucl/U1/U1  ( .x(l[14]), .a(n6), .b(l[14]), .c(n1), .d(\U14/ni 
        ), .e(\U14/nh ) );
    ao23_1 \U14/Uch/U1/U1  ( .x(h[14]), .a(n6), .b(h[14]), .c(n3), .d(i[14]), 
        .e(\U14/nl ) );
    inv_1 \U13/Uii  ( .x(\U13/ni ), .a(i[13]) );
    inv_1 \U13/Uih  ( .x(\U13/nh ), .a(h[13]) );
    inv_1 \U13/Uil  ( .x(\U13/nl ), .a(l[13]) );
    ao23_1 \U13/Ucl/U1/U1  ( .x(l[13]), .a(n6), .b(l[13]), .c(n4), .d(\U13/ni 
        ), .e(\U13/nh ) );
    ao23_1 \U13/Uch/U1/U1  ( .x(h[13]), .a(n6), .b(h[13]), .c(n4), .d(i[13]), 
        .e(\U13/nl ) );
    inv_1 \U12/Uii  ( .x(\U12/ni ), .a(i[12]) );
    inv_1 \U12/Uih  ( .x(\U12/nh ), .a(h[12]) );
    inv_1 \U12/Uil  ( .x(\U12/nl ), .a(l[12]) );
    ao23_1 \U12/Ucl/U1/U1  ( .x(l[12]), .a(n5), .b(l[12]), .c(n4), .d(\U12/ni 
        ), .e(\U12/nh ) );
    ao23_1 \U12/Uch/U1/U1  ( .x(h[12]), .a(n5), .b(h[12]), .c(n4), .d(i[12]), 
        .e(\U12/nl ) );
    inv_1 \U11/Uii  ( .x(\U11/ni ), .a(i[11]) );
    inv_1 \U11/Uih  ( .x(\U11/nh ), .a(h[11]) );
    inv_1 \U11/Uil  ( .x(\U11/nl ), .a(l[11]) );
    ao23_1 \U11/Ucl/U1/U1  ( .x(l[11]), .a(n5), .b(l[11]), .c(n4), .d(\U11/ni 
        ), .e(\U11/nh ) );
    ao23_1 \U11/Uch/U1/U1  ( .x(h[11]), .a(n5), .b(h[11]), .c(n4), .d(i[11]), 
        .e(\U11/nl ) );
    inv_1 \U10/Uii  ( .x(\U10/ni ), .a(i[10]) );
    inv_1 \U10/Uih  ( .x(\U10/nh ), .a(h[10]) );
    inv_1 \U10/Uil  ( .x(\U10/nl ), .a(l[10]) );
    ao23_1 \U10/Ucl/U1/U1  ( .x(l[10]), .a(n5), .b(l[10]), .c(n3), .d(\U10/ni 
        ), .e(\U10/nh ) );
    ao23_1 \U10/Uch/U1/U1  ( .x(h[10]), .a(n5), .b(h[10]), .c(n3), .d(i[10]), 
        .e(\U10/nl ) );
    inv_1 \U9/Uii  ( .x(\U9/ni ), .a(i[9]) );
    inv_1 \U9/Uih  ( .x(\U9/nh ), .a(h[9]) );
    inv_1 \U9/Uil  ( .x(\U9/nl ), .a(l[9]) );
    ao23_1 \U9/Ucl/U1/U1  ( .x(l[9]), .a(n5), .b(l[9]), .c(n3), .d(\U9/ni ), 
        .e(\U9/nh ) );
    ao23_1 \U9/Uch/U1/U1  ( .x(h[9]), .a(n5), .b(h[9]), .c(n3), .d(i[9]), .e(
        \U9/nl ) );
    inv_1 \U8/Uii  ( .x(\U8/ni ), .a(i[8]) );
    inv_1 \U8/Uih  ( .x(\U8/nh ), .a(h[8]) );
    inv_1 \U8/Uil  ( .x(\U8/nl ), .a(l[8]) );
    ao23_1 \U8/Ucl/U1/U1  ( .x(l[8]), .a(n5), .b(l[8]), .c(n3), .d(\U8/ni ), 
        .e(\U8/nh ) );
    ao23_1 \U8/Uch/U1/U1  ( .x(h[8]), .a(n5), .b(h[8]), .c(n3), .d(i[8]), .e(
        \U8/nl ) );
    inv_1 \U7/Uii  ( .x(\U7/ni ), .a(i[7]) );
    inv_1 \U7/Uih  ( .x(\U7/nh ), .a(h[7]) );
    inv_1 \U7/Uil  ( .x(\U7/nl ), .a(l[7]) );
    ao23_1 \U7/Ucl/U1/U1  ( .x(l[7]), .a(n7), .b(l[7]), .c(n3), .d(\U7/ni ), 
        .e(\U7/nh ) );
    ao23_1 \U7/Uch/U1/U1  ( .x(h[7]), .a(n7), .b(h[7]), .c(n2), .d(i[7]), .e(
        \U7/nl ) );
    inv_1 \U6/Uii  ( .x(\U6/ni ), .a(i[6]) );
    inv_1 \U6/Uih  ( .x(\U6/nh ), .a(h[6]) );
    inv_1 \U6/Uil  ( .x(\U6/nl ), .a(l[6]) );
    ao23_1 \U6/Ucl/U1/U1  ( .x(l[6]), .a(n7), .b(l[6]), .c(n2), .d(\U6/ni ), 
        .e(\U6/nh ) );
    ao23_1 \U6/Uch/U1/U1  ( .x(h[6]), .a(n7), .b(h[6]), .c(n2), .d(i[6]), .e(
        \U6/nl ) );
    inv_1 \U5/Uii  ( .x(\U5/ni ), .a(i[5]) );
    inv_1 \U5/Uih  ( .x(\U5/nh ), .a(h[5]) );
    inv_1 \U5/Uil  ( .x(\U5/nl ), .a(l[5]) );
    ao23_1 \U5/Ucl/U1/U1  ( .x(l[5]), .a(n7), .b(l[5]), .c(n2), .d(\U5/ni ), 
        .e(\U5/nh ) );
    ao23_1 \U5/Uch/U1/U1  ( .x(h[5]), .a(n7), .b(h[5]), .c(n2), .d(i[5]), .e(
        \U5/nl ) );
    inv_1 \U4/Uii  ( .x(\U4/ni ), .a(i[4]) );
    inv_1 \U4/Uih  ( .x(\U4/nh ), .a(h[4]) );
    inv_1 \U4/Uil  ( .x(\U4/nl ), .a(l[4]) );
    ao23_1 \U4/Ucl/U1/U1  ( .x(l[4]), .a(n6), .b(l[4]), .c(n2), .d(\U4/ni ), 
        .e(\U4/nh ) );
    ao23_1 \U4/Uch/U1/U1  ( .x(h[4]), .a(n6), .b(h[4]), .c(n2), .d(i[4]), .e(
        \U4/nl ) );
    inv_1 \U3/Uii  ( .x(\U3/ni ), .a(i[3]) );
    inv_1 \U3/Uih  ( .x(\U3/nh ), .a(h[3]) );
    inv_1 \U3/Uil  ( .x(\U3/nl ), .a(l[3]) );
    ao23_1 \U3/Ucl/U1/U1  ( .x(l[3]), .a(n6), .b(l[3]), .c(n2), .d(\U3/ni ), 
        .e(\U3/nh ) );
    ao23_1 \U3/Uch/U1/U1  ( .x(h[3]), .a(n8), .b(h[3]), .c(n1), .d(i[3]), .e(
        \U3/nl ) );
    inv_1 \U2/Uii  ( .x(\U2/ni ), .a(i[2]) );
    inv_1 \U2/Uih  ( .x(\U2/nh ), .a(h[2]) );
    inv_1 \U2/Uil  ( .x(\U2/nl ), .a(l[2]) );
    ao23_1 \U2/Ucl/U1/U1  ( .x(l[2]), .a(n8), .b(l[2]), .c(n1), .d(\U2/ni ), 
        .e(\U2/nh ) );
    ao23_1 \U2/Uch/U1/U1  ( .x(h[2]), .a(n8), .b(h[2]), .c(n1), .d(i[2]), .e(
        \U2/nl ) );
    inv_1 \U1/Uii  ( .x(\U1/ni ), .a(i[1]) );
    inv_1 \U1/Uih  ( .x(\U1/nh ), .a(h[1]) );
    inv_1 \U1/Uil  ( .x(\U1/nl ), .a(l[1]) );
    ao23_1 \U1/Ucl/U1/U1  ( .x(l[1]), .a(n8), .b(l[1]), .c(n1), .d(\U1/ni ), 
        .e(\U1/nh ) );
    ao23_1 \U1/Uch/U1/U1  ( .x(h[1]), .a(n8), .b(h[1]), .c(n1), .d(i[1]), .e(
        \U1/nl ) );
    inv_1 \U0/Uii  ( .x(\U0/ni ), .a(i[0]) );
    inv_1 \U0/Uih  ( .x(\U0/nh ), .a(h[0]) );
    inv_1 \U0/Uil  ( .x(\U0/nl ), .a(l[0]) );
    ao23_1 \U0/Ucl/U1/U1  ( .x(l[0]), .a(n8), .b(l[0]), .c(n1), .d(\U0/ni ), 
        .e(\U0/nh ) );
    ao23_1 \U0/Uch/U1/U1  ( .x(h[0]), .a(n8), .b(h[0]), .c(n1), .d(i[0]), .e(
        \U0/nl ) );
    buf_16 U1 ( .x(n1), .a(n12) );
    buf_16 U2 ( .x(n2), .a(n12) );
    buf_16 U3 ( .x(n3), .a(n12) );
    buf_16 U4 ( .x(n4), .a(n11) );
    buf_16 U5 ( .x(n5), .a(n11) );
    buf_16 U6 ( .x(n6), .a(n11) );
    buf_16 U7 ( .x(n7), .a(n10) );
    buf_16 U8 ( .x(n8), .a(n10) );
    buf_16 U9 ( .x(n9), .a(n10) );
    buf_16 U10 ( .x(n10), .a(req) );
    buf_16 U11 ( .x(n11), .a(req) );
    buf_16 U12 ( .x(n12), .a(req) );
endmodule


module matched_delay_cp2slave_resp_wb ( x, a );
input  a;
output x;
    buf_1 I1 ( .x(x), .a(a) );
endmodule


module matched_delay_cp2slave_com_wb ( x, a );
input  a;
output x;
    buf_1 I1 ( .x(x), .a(a) );
endmodule


module cp2slave_wb ( tc_seq, tc_size, tc_itag, tc_wd, tc_lock, tc_a, tc_rnw, 
    tc_ok, tc_defer, tc_slow, tc_ack, req_in, ts_i, st_i, we_i, mult_i, adr_i, 
    dat_i, seq_i, prd_i, sel_i, ack_in, tr_rd, tr_err, tr_size, tr_ack, tr_rnw, 
    req_out, dat_o, err_o, rty_o, acc_o, sel_o, mult_o, rt_o, ack_out, reset
     );
input  [1:0] tc_seq;
input  [3:0] tc_size;
input  [9:0] tc_itag;
input  [63:0] tc_wd;
input  [1:0] tc_lock;
input  [63:0] tc_a;
input  [1:0] tc_rnw;
output [2:0] ts_i;
output [4:0] st_i;
output [31:0] adr_i;
output [31:0] dat_i;
output [3:0] sel_i;
output [63:0] tr_rd;
output [1:0] tr_err;
output [3:0] tr_size;
output [1:0] tr_rnw;
input  [31:0] dat_o;
input  [3:0] sel_o;
input  [4:0] rt_o;
input  ack_in, tr_ack, req_out, err_o, rty_o, acc_o, mult_o, reset;
output tc_ok, tc_defer, tc_slow, tc_ack, req_in, we_i, mult_i, seq_i, prd_i, 
    ack_out;
    wire tc_wd_63, tc_wd_62, tc_wd_61, tc_wd_60, tc_wd_59, tc_wd_58, tc_wd_56, 
        tc_wd_55, tc_wd_54, tc_wd_53, tc_wd_52, tc_wd_51, tc_wd_50, tc_wd_49, 
        tc_wd_48, tc_wd_47, tc_wd_46, tc_wd_45, tc_wd_44, tc_wd_43, tc_wd_40, 
        tc_wd_39, tc_wd_38, tc_wd_36, tc_wd_32, tc_a_60, tc_a_58, sel_i_3, n1, 
        n334, n311, n129, n309, n310, n315, n348, n349, n350, n456, n336, n457, 
        n345, n303, n505, n193, n476, n479, n229, n226, n257, n263, n260, n268, 
        n269, n270, n265, n266, n267, n277, n252, n248, n249, n250, n245, n246, 
        n247, n242, n243, n244, n222, n223, n224, n220, n234, n235, n236, n231, 
        n232, n233, n205, n206, n207, n203, n199, n200, n201, n197, n218, n214, 
        n215, n216, n211, n212, n213, n208, n209, n210, n374, n375, n368, n251, 
        n280, n274, n271, n427, n196, n424, n202, n240, n237, n413, n219, n421, 
        n418, n416, n428, n425, n422, n414, n411, n408, n238, n272, n351, n366, 
        n335, n355, n531, n532, respond, n313, n121, n122, n359, n360, n123, 
        n337, n124, n125, n126, n127, n217, n128, n312, n130, n284, n285, n449, 
        n282, n283, n380, n279, n276, n397, n454, n463, n453, n395, n404, n383, 
        n443, n477, n455, n230, n135, n305, n487, n302, n445, n446, n442, n136, 
        n320, n400, n137, n340, n198, n386, n381, n478, n475, n407, n402, n204, 
        n221, n141, n321, n483, n484, n485, n480, n474, n227, n188, n517, n525, 
        n180, n401, n387, n394, n481, n482, n491, n195, n492, n369, n181, n429, 
        n415, n324, n343, n363, n319, n344, n354, n304, n330, n497, n496, n291, 
        n438, n373, n367, n439, n440, n333, n308, n297, n347, n301, n503, n499, 
        n502, n498, n288, n327, n316, n298, n294, n358, complb0, n189, n510, 
        n507, n192, n473, n508, n471, n488, n489, n490, complw0, n182, n183, 
        n184, n185, n364, n365, n391, n388, n430, n423, n426, n431, n417, n419, 
        n420, n432, n409, n410, n412, n433, n403, n405, n406, n434, n396, n398, 
        n399, n435, n389, n390, n392, n393, n436, n382, n384, n385, n437, n376, 
        n377, n378, n379, n441, n370, n444, n470, n472, n194, n486, n493, n494, 
        n495, n191, n500, n501, n504, n506, n509, n511, n465, n466, n468, n512, 
        n460, n513, n514, n462, n459, n515, n516, n518, n452, n519, n450, n520, 
        n522, n521, n523, n524, n371, complb1, n190, complw1, n447, n469, n5, 
        n3, n4, n448, n467, n461, n372, n451, n458, n464, n273, n262, n259, 
        n256, n253, n228, n225, n239, n361, n356, n331, n295, n275, n281, n278, 
        n264, n261, n258, n254, n255, n241, n341, n328, n325, n338, n362, n357, 
        n352, n299, n289, n286, n292, n317, n322, n306, n314, n332, n296, n342, 
        n346, n329, n326, n339, n353, n300, n290, n287, n293, n318, n323, n307, 
        req_out_delayed, _25_net_, n529, n530, _24_net_, _26_net_, n142, 
        req_in_i, n186, n187, all_w, all_r, comp_basic, 
        \cg_all_w/__tmp99/loop , comp_wd, \Usze1/ni , \Usze1/nh , \Usze1/nl , 
        n2, \Usze0/ni , \Usze0/nh , \Usze0/nl , \Urnw/ni , \Urnw/nh , 
        \Urnw/nl , \Uerr/ni , \Uerr/nh , \Uerr/nl ;
    assign tc_wd_63 = tc_wd[63];
    assign tc_wd_62 = tc_wd[62];
    assign tc_wd_61 = tc_wd[61];
    assign tc_wd_60 = tc_wd[60];
    assign tc_wd_59 = tc_wd[59];
    assign tc_wd_58 = tc_wd[58];
    assign tc_wd_56 = tc_wd[56];
    assign tc_wd_55 = tc_wd[55];
    assign tc_wd_54 = tc_wd[54];
    assign tc_wd_53 = tc_wd[53];
    assign tc_wd_52 = tc_wd[52];
    assign tc_wd_51 = tc_wd[51];
    assign tc_wd_50 = tc_wd[50];
    assign tc_wd_49 = tc_wd[49];
    assign tc_wd_48 = tc_wd[48];
    assign tc_wd_47 = tc_wd[47];
    assign tc_wd_46 = tc_wd[46];
    assign tc_wd_45 = tc_wd[45];
    assign tc_wd_44 = tc_wd[44];
    assign tc_wd_43 = tc_wd[43];
    assign tc_wd_40 = tc_wd[40];
    assign tc_wd_39 = tc_wd[39];
    assign tc_wd_38 = tc_wd[38];
    assign tc_wd_36 = tc_wd[36];
    assign tc_wd_32 = tc_wd[32];
    assign tc_a_60 = tc_a[60];
    assign tc_a_58 = tc_a[58];
    assign ts_i[2] = 1'b0;
    assign ts_i[1] = 1'b0;
    assign ts_i[0] = 1'b0;
    assign adr_i[28] = tc_a_60;
    assign adr_i[26] = tc_a_58;
    assign dat_i[31] = tc_wd_63;
    assign dat_i[30] = tc_wd_62;
    assign dat_i[29] = tc_wd_61;
    assign dat_i[28] = tc_wd_60;
    assign dat_i[27] = tc_wd_59;
    assign dat_i[26] = tc_wd_58;
    assign dat_i[24] = tc_wd_56;
    assign dat_i[23] = tc_wd_55;
    assign dat_i[22] = tc_wd_54;
    assign dat_i[21] = tc_wd_53;
    assign dat_i[20] = tc_wd_52;
    assign dat_i[19] = tc_wd_51;
    assign dat_i[18] = tc_wd_50;
    assign dat_i[17] = tc_wd_49;
    assign dat_i[16] = tc_wd_48;
    assign dat_i[15] = tc_wd_47;
    assign dat_i[14] = tc_wd_46;
    assign dat_i[13] = tc_wd_45;
    assign dat_i[12] = tc_wd_44;
    assign dat_i[11] = tc_wd_43;
    assign dat_i[8] = tc_wd_40;
    assign dat_i[7] = tc_wd_39;
    assign dat_i[6] = tc_wd_38;
    assign dat_i[4] = tc_wd_36;
    assign dat_i[0] = tc_wd_32;
    assign prd_i = 1'b0;
    assign sel_i[3] = sel_i_3;
    assign sel_i[2] = sel_i_3;
    assign sel_i[0] = 1'b1;
    assign tc_ack = ack_in;
    assign ack_out = tr_ack;
    sr2dr_word_6 Urd ( .i(dat_o), .req(n1), .h(tr_rd[63:32]), .l(tr_rd[31:0])
         );
    inv_1 U3 ( .x(n334), .a(tc_a[7]) );
    inv_1 U5 ( .x(n311), .a(tc_a[21]) );
    and2_1 U6 ( .x(n129), .a(n309), .b(n310) );
    inv_1 U7 ( .x(n309), .a(tc_a[6]) );
    inv_1 U9 ( .x(n315), .a(tc_itag[4]) );
    nand2_1 U10 ( .x(n348), .a(n349), .b(n350) );
    inv_1 U11 ( .x(n349), .a(tc_a[12]) );
    inv_1 U12 ( .x(n456), .a(n348) );
    inv_1 U13 ( .x(n336), .a(tc_a[30]) );
    inv_1 U14 ( .x(n457), .a(n345) );
    inv_1 U15 ( .x(n303), .a(tc_a[8]) );
    nand3_1 U16 ( .x(n505), .a(n193), .b(n476), .c(n479) );
    inv_1 U17 ( .x(n229), .a(tc_wd[5]) );
    inv_1 U18 ( .x(n226), .a(tc_wd[3]) );
    inv_1 U19 ( .x(n257), .a(tc_wd[16]) );
    inv_1 U20 ( .x(n263), .a(tc_wd[21]) );
    inv_1 U21 ( .x(n260), .a(tc_wd[19]) );
    nand2_1 U22 ( .x(n268), .a(n269), .b(n270) );
    inv_1 U23 ( .x(n269), .a(tc_wd[23]) );
    inv_1 U24 ( .x(n270), .a(tc_wd_55) );
    nand2_1 U25 ( .x(n265), .a(n266), .b(n267) );
    inv_1 U26 ( .x(n266), .a(tc_wd[20]) );
    inv_1 U27 ( .x(n277), .a(tc_wd[27]) );
    inv_1 U28 ( .x(n252), .a(tc_wd_47) );
    nand2_1 U29 ( .x(n248), .a(n249), .b(n250) );
    inv_1 U30 ( .x(n249), .a(tc_wd[12]) );
    nand2_1 U31 ( .x(n245), .a(n246), .b(n247) );
    inv_1 U32 ( .x(n246), .a(tc_wd[13]) );
    inv_1 U33 ( .x(n247), .a(tc_wd_45) );
    nand2_1 U34 ( .x(n242), .a(n243), .b(n244) );
    inv_1 U35 ( .x(n243), .a(tc_wd[11]) );
    nand2_1 U36 ( .x(n222), .a(n223), .b(n224) );
    inv_1 U37 ( .x(n223), .a(tc_wd[0]) );
    inv_1 U38 ( .x(n220), .a(tc_wd[1]) );
    nand2_1 U39 ( .x(n234), .a(n235), .b(n236) );
    inv_1 U40 ( .x(n235), .a(tc_wd[7]) );
    nand2_1 U41 ( .x(n231), .a(n232), .b(n233) );
    inv_1 U42 ( .x(n232), .a(tc_wd[4]) );
    nand2_1 U43 ( .x(n205), .a(n206), .b(n207) );
    inv_1 U44 ( .x(n206), .a(tc_wd[18]) );
    inv_1 U45 ( .x(n203), .a(tc_wd[10]) );
    nand2_1 U46 ( .x(n199), .a(n200), .b(n201) );
    inv_1 U47 ( .x(n200), .a(tc_wd[6]) );
    inv_1 U48 ( .x(n197), .a(tc_wd[2]) );
    inv_1 U49 ( .x(n218), .a(tc_wd_46) );
    nand2_1 U50 ( .x(n214), .a(n215), .b(n216) );
    inv_1 U51 ( .x(n215), .a(tc_wd[30]) );
    nand2_1 U52 ( .x(n211), .a(n212), .b(n213) );
    inv_1 U53 ( .x(n213), .a(tc_wd_58) );
    nand2_1 U54 ( .x(n208), .a(n209), .b(n210) );
    inv_1 U55 ( .x(n209), .a(tc_wd[22]) );
    inv_1 U56 ( .x(n374), .a(tc_rnw[0]) );
    inv_1 U57 ( .x(n375), .a(tc_rnw[1]) );
    inv_1 U58 ( .x(n368), .a(tc_a[18]) );
    inv_1 U59 ( .x(n244), .a(tc_wd_43) );
    inv_1 U60 ( .x(n251), .a(tc_wd[15]) );
    inv_1 U61 ( .x(n250), .a(tc_wd_44) );
    inv_1 U62 ( .x(n280), .a(tc_wd[29]) );
    inv_1 U63 ( .x(n267), .a(tc_wd_52) );
    inv_1 U64 ( .x(n274), .a(tc_wd[24]) );
    inv_1 U65 ( .x(n271), .a(tc_wd[25]) );
    inv_1 U66 ( .x(n212), .a(tc_wd[26]) );
    inv_1 U67 ( .x(n210), .a(tc_wd_54) );
    inv_1 U68 ( .x(n216), .a(tc_wd_62) );
    inv_1 U69 ( .x(n201), .a(tc_wd_38) );
    inv_1 U70 ( .x(n427), .a(n196) );
    inv_1 U71 ( .x(n207), .a(tc_wd_50) );
    inv_1 U72 ( .x(n424), .a(n202) );
    inv_1 U73 ( .x(n236), .a(tc_wd_39) );
    inv_1 U74 ( .x(n233), .a(tc_wd_36) );
    inv_1 U75 ( .x(n240), .a(tc_wd[8]) );
    inv_1 U76 ( .x(n237), .a(tc_wd[9]) );
    inv_1 U77 ( .x(n224), .a(tc_wd_32) );
    inv_1 U78 ( .x(n413), .a(n219) );
    nand2_1 U79 ( .x(n421), .a(n418), .b(n416) );
    nand2_1 U80 ( .x(n428), .a(n425), .b(n422) );
    nand2_1 U81 ( .x(n414), .a(n411), .b(n408) );
    inv_1 U82 ( .x(n238), .a(tc_wd[41]) );
    inv_1 U83 ( .x(n272), .a(tc_wd[57]) );
    inv_1 U84 ( .x(n350), .a(tc_a[44]) );
    inv_1 U85 ( .x(n351), .a(tc_a[43]) );
    inv_1 U86 ( .x(n366), .a(tc_a[41]) );
    inv_1 U87 ( .x(n335), .a(tc_a[39]) );
    inv_1 U88 ( .x(n310), .a(tc_a[38]) );
    inv_1 U89 ( .x(n355), .a(tc_a[52]) );
    and3_1 U90 ( .x(tc_ok), .a(n531), .b(n532), .c(respond) );
    and2_1 U91 ( .x(tc_slow), .a(respond), .b(acc_o) );
    inv_1 U94 ( .x(n313), .a(tc_itag[5]) );
    and2_1 U95 ( .x(n121), .a(n334), .b(n335) );
    and2_1 U96 ( .x(n122), .a(n359), .b(n360) );
    and2_1 U97 ( .x(n123), .a(n336), .b(n337) );
    and2_1 U98 ( .x(n124), .a(n237), .b(n238) );
    and2_1 U99 ( .x(n125), .a(n251), .b(n252) );
    and2_1 U100 ( .x(n126), .a(n271), .b(n272) );
    and2_1 U101 ( .x(n127), .a(n217), .b(n218) );
    and2_1 U102 ( .x(n128), .a(n311), .b(n312) );
    nor2_1 U103 ( .x(n130), .a(tc_size[3]), .b(tc_size[2]) );
    nand2i_1 U105 ( .x(n284), .a(tc_wd[31]), .b(n285) );
    oa22_1 U106 ( .x(n449), .a(tc_a[27]), .b(tc_a[59]), .c(tc_a[54]), .d(tc_a
        [22]) );
    inv_1 U107 ( .x(n359), .a(tc_a[27]) );
    inv_1 U108 ( .x(n360), .a(tc_a[59]) );
    nand2i_1 U109 ( .x(n282), .a(tc_wd[28]), .b(n283) );
    nor2_1 U110 ( .x(n479), .a(tc_itag[0]), .b(tc_itag[5]) );
    nand4_1 U112 ( .x(n380), .a(n279), .b(n276), .c(n284), .d(n282) );
    aoi21_1 U113 ( .x(n425), .a(n200), .b(n201), .c(n427) );
    oa22_1 U114 ( .x(n397), .a(tc_wd[13]), .b(tc_wd_45), .c(tc_wd[11]), .d(
        tc_wd_43) );
    nor2_1 U115 ( .x(n454), .a(tc_a[20]), .b(tc_a[52]) );
    aoi21_1 U116 ( .x(n422), .a(n206), .b(n207), .c(n424) );
    oa22_1 U117 ( .x(n418), .a(tc_wd[26]), .b(tc_wd_58), .c(tc_wd[22]), .d(
        tc_wd_54) );
    oa22_1 U118 ( .x(n416), .a(tc_wd[14]), .b(tc_wd_46), .c(tc_wd[30]), .d(
        tc_wd_62) );
    inv_1 U119 ( .x(n217), .a(tc_wd[14]) );
    aoi22_1 U120 ( .x(n463), .a(n336), .b(n337), .c(n334), .d(n335) );
    nor2_1 U121 ( .x(n453), .a(tc_a[11]), .b(tc_a[43]) );
    oa22_1 U122 ( .x(n395), .a(tc_wd[15]), .b(tc_wd_47), .c(tc_wd[12]), .d(
        tc_wd_44) );
    oa22_1 U123 ( .x(n404), .a(tc_wd[7]), .b(tc_wd_39), .c(tc_wd[4]), .d(
        tc_wd_36) );
    oa22_1 U124 ( .x(n383), .a(tc_wd[23]), .b(tc_wd_55), .c(tc_wd[20]), .d(
        tc_wd_52) );
    aoi21_1 U125 ( .x(n411), .a(n223), .b(n224), .c(n413) );
    nor2_1 U126 ( .x(n443), .a(tc_a[49]), .b(tc_a[17]) );
    aoi22_1 U127 ( .x(n477), .a(n311), .b(n312), .c(n309), .d(n310) );
    oa21_1 U128 ( .x(n455), .a(tc_a[12]), .b(tc_a[44]), .c(n345) );
    inv_1 U129 ( .x(dat_i[5]), .a(n230) );
    inv_1 U130 ( .x(dat_i[9]), .a(n238) );
    inv_1 U131 ( .x(dat_i[25]), .a(n272) );
    buf_1 U132 ( .x(sel_i_3), .a(tc_size[3]) );
    buf_1 U133 ( .x(adr_i[16]), .a(tc_a[48]) );
    nor2_1 U134 ( .x(n135), .a(tc_a[14]), .b(tc_a[46]) );
    inv_1 U135 ( .x(n305), .a(tc_a[46]) );
    inv_1 U136 ( .x(n487), .a(n302) );
    nand2i_1 U137 ( .x(n445), .a(n446), .b(n442) );
    nor2_1 U138 ( .x(n136), .a(tc_a[29]), .b(tc_a[61]) );
    inv_1 U139 ( .x(n320), .a(tc_a[61]) );
    nand2_1 U140 ( .x(n400), .a(n397), .b(n395) );
    inv_1 U141 ( .x(n137), .a(n340) );
    inv_1 U142 ( .x(dat_i[2]), .a(n198) );
    nand2_1 U143 ( .x(n386), .a(n383), .b(n381) );
    nand3i_1 U144 ( .x(n478), .a(n479), .b(n477), .c(n475) );
    nand2_1 U145 ( .x(n407), .a(n404), .b(n402) );
    inv_1 U146 ( .x(dat_i[10]), .a(n204) );
    inv_1 U147 ( .x(dat_i[1]), .a(n221) );
    nor2_1 U148 ( .x(n141), .a(tc_a[3]), .b(tc_a[35]) );
    inv_1 U149 ( .x(n321), .a(tc_a[35]) );
    nor2_1 U151 ( .x(n483), .a(n484), .b(n485) );
    nor2_1 U152 ( .x(n480), .a(n474), .b(n478) );
    inv_1 U153 ( .x(dat_i[3]), .a(n227) );
    nor2_1 U154 ( .x(n188), .a(n517), .b(n525) );
    nand2_1 U155 ( .x(n180), .a(n401), .b(n387) );
    nor2_1 U156 ( .x(n401), .a(n394), .b(n400) );
    nor2_1 U157 ( .x(n387), .a(n380), .b(n386) );
    nor2_1 U158 ( .x(n481), .a(n482), .b(n135) );
    nor2_1 U159 ( .x(n491), .a(n195), .b(n492) );
    nor2_1 U160 ( .x(n195), .a(tc_size[1]), .b(tc_size[3]) );
    inv_1 U161 ( .x(adr_i[18]), .a(n369) );
    nand2_1 U162 ( .x(n181), .a(n429), .b(n415) );
    nor2_1 U163 ( .x(n429), .a(n421), .b(n428) );
    nor2_1 U164 ( .x(n415), .a(n407), .b(n414) );
    inv_1 U165 ( .x(adr_i[0]), .a(n324) );
    inv_1 U166 ( .x(n324), .a(tc_a[32]) );
    inv_1 U167 ( .x(sel_i[1]), .a(n130) );
    inv_1 U168 ( .x(st_i[2]), .a(n343) );
    inv_1 U169 ( .x(adr_i[9]), .a(n366) );
    inv_1 U170 ( .x(adr_i[24]), .a(n363) );
    inv_1 U171 ( .x(adr_i[19]), .a(n319) );
    inv_1 U172 ( .x(n319), .a(tc_a[51]) );
    inv_1 U173 ( .x(n369), .a(tc_a[50]) );
    inv_1 U174 ( .x(st_i[3]), .a(n344) );
    inv_1 U175 ( .x(adr_i[13]), .a(n354) );
    inv_1 U176 ( .x(adr_i[12]), .a(n350) );
    inv_1 U177 ( .x(adr_i[8]), .a(n304) );
    inv_1 U178 ( .x(n304), .a(tc_a[40]) );
    inv_1 U179 ( .x(adr_i[2]), .a(n330) );
    buf_1 U180 ( .x(adr_i[17]), .a(tc_a[49]) );
    nand2_1 U181 ( .x(n497), .a(n496), .b(n130) );
    inv_1 U182 ( .x(adr_i[10]), .a(n291) );
    and2_1 U183 ( .x(n438), .a(n373), .b(n367) );
    inv_1 U184 ( .x(n439), .a(n373) );
    inv_1 U185 ( .x(n440), .a(n367) );
    inv_1 U186 ( .x(adr_i[20]), .a(n355) );
    inv_1 U187 ( .x(adr_i[27]), .a(n360) );
    inv_1 U188 ( .x(adr_i[4]), .a(n333) );
    inv_1 U189 ( .x(adr_i[25]), .a(n308) );
    inv_1 U190 ( .x(adr_i[30]), .a(n337) );
    inv_1 U191 ( .x(adr_i[31]), .a(n297) );
    inv_1 U192 ( .x(n297), .a(tc_a[63]) );
    inv_1 U193 ( .x(adr_i[15]), .a(n347) );
    inv_1 U194 ( .x(adr_i[11]), .a(n351) );
    inv_1 U195 ( .x(adr_i[1]), .a(n301) );
    inv_1 U196 ( .x(n301), .a(tc_a[33]) );
    nand2_1 U197 ( .x(n503), .a(n499), .b(n502) );
    nor2_1 U198 ( .x(n499), .a(n497), .b(n498) );
    inv_1 U199 ( .x(adr_i[21]), .a(n312) );
    inv_1 U200 ( .x(n312), .a(tc_a[53]) );
    inv_1 U201 ( .x(seq_i), .a(n288) );
    inv_1 U202 ( .x(adr_i[5]), .a(n327) );
    inv_1 U203 ( .x(st_i[4]), .a(n316) );
    inv_1 U204 ( .x(n316), .a(tc_itag[9]) );
    inv_1 U205 ( .x(st_i[1]), .a(n298) );
    inv_1 U206 ( .x(adr_i[23]), .a(n294) );
    inv_1 U207 ( .x(adr_i[22]), .a(n358) );
    nand2_1 U208 ( .x(complb0), .a(n188), .b(n189) );
    nor2_1 U209 ( .x(n189), .a(n503), .b(n510) );
    inv_1 U210 ( .x(adr_i[29]), .a(n320) );
    inv_1 U211 ( .x(adr_i[7]), .a(n335) );
    inv_1 U212 ( .x(adr_i[14]), .a(n305) );
    inv_1 U213 ( .x(adr_i[6]), .a(n310) );
    inv_1 U214 ( .x(st_i[0]), .a(n313) );
    inv_1 U215 ( .x(adr_i[3]), .a(n321) );
    nand3_1 U218 ( .x(n507), .a(n192), .b(n136), .c(n473) );
    nand2_1 U219 ( .x(n508), .a(n471), .b(n141) );
    nor2_1 U220 ( .x(n488), .a(n489), .b(n490) );
    nand4_1 U222 ( .x(complw0), .a(n182), .b(n183), .c(n184), .d(n185) );
    nor2_1 U223 ( .x(n192), .a(tc_a_58), .b(tc_a[26]) );
    nor2_1 U224 ( .x(n193), .a(tc_a[48]), .b(tc_a[16]) );
    nand2_1 U225 ( .x(n364), .a(n365), .b(n366) );
    nand2_1 U226 ( .x(n394), .a(n391), .b(n388) );
    nand4_1 U227 ( .x(n430), .a(n423), .b(n424), .c(n426), .d(n427) );
    nand4_1 U228 ( .x(n431), .a(n127), .b(n417), .c(n419), .d(n420) );
    nor2_1 U229 ( .x(n185), .a(n430), .b(n431) );
    nand4_1 U230 ( .x(n432), .a(n409), .b(n410), .c(n412), .d(n413) );
    nand4_1 U231 ( .x(n433), .a(n403), .b(n124), .c(n405), .d(n406) );
    nor2_1 U232 ( .x(n184), .a(n432), .b(n433) );
    nand4_1 U233 ( .x(n434), .a(n125), .b(n396), .c(n398), .d(n399) );
    nand4_1 U234 ( .x(n435), .a(n389), .b(n390), .c(n392), .d(n393) );
    nor2_1 U235 ( .x(n183), .a(n434), .b(n435) );
    nand4_1 U236 ( .x(n436), .a(n382), .b(n126), .c(n384), .d(n385) );
    nand4_1 U237 ( .x(n437), .a(n376), .b(n377), .c(n378), .d(n379) );
    nor2_1 U238 ( .x(n182), .a(n436), .b(n437) );
    nand2_1 U239 ( .x(n441), .a(n438), .b(n370) );
    nor2_1 U240 ( .x(n442), .a(n443), .b(n444) );
    nor3_1 U241 ( .x(n470), .a(n471), .b(n136), .c(n141) );
    nor3_1 U242 ( .x(n472), .a(n473), .b(n192), .c(n193) );
    nand2_1 U243 ( .x(n474), .a(n472), .b(n470) );
    nor2_1 U244 ( .x(n475), .a(n476), .b(n194) );
    nand3i_1 U245 ( .x(n486), .a(n487), .b(n481), .c(n483) );
    nand3i_1 U246 ( .x(n493), .a(n494), .b(n488), .c(n491) );
    nor2_1 U247 ( .x(n495), .a(n493), .b(n486) );
    nand2_1 U248 ( .x(n191), .a(n495), .b(n480) );
    nand3_1 U249 ( .x(n498), .a(n489), .b(n492), .c(n490) );
    nand3_1 U250 ( .x(n500), .a(n485), .b(n494), .c(n484) );
    nand2_1 U251 ( .x(n501), .a(n135), .b(n487) );
    nor2_1 U252 ( .x(n502), .a(n500), .b(n501) );
    nand3_1 U253 ( .x(n504), .a(n128), .b(n482), .c(n129) );
    nor2_1 U254 ( .x(n506), .a(n504), .b(n505) );
    nor2_1 U255 ( .x(n509), .a(n507), .b(n508) );
    nand2_1 U256 ( .x(n510), .a(n509), .b(n506) );
    nand3_1 U257 ( .x(n511), .a(n465), .b(n466), .c(n468) );
    nand3_1 U258 ( .x(n512), .a(n123), .b(n121), .c(n460) );
    nor2_1 U259 ( .x(n513), .a(n511), .b(n512) );
    nand3_1 U260 ( .x(n514), .a(n462), .b(n459), .c(n457) );
    nand2_1 U261 ( .x(n515), .a(n453), .b(n456) );
    nor2_1 U262 ( .x(n516), .a(n514), .b(n515) );
    nand2_1 U263 ( .x(n517), .a(n516), .b(n513) );
    nand2_1 U264 ( .x(n518), .a(n454), .b(n452) );
    nor2i_1 U265 ( .x(n519), .a(n450), .b(n518) );
    nand2_1 U266 ( .x(n520), .a(n444), .b(n122) );
    nor2i_1 U267 ( .x(n522), .a(n446), .b(n521) );
    nand2_1 U268 ( .x(n523), .a(n439), .b(n524) );
    inv_1 U270 ( .x(n365), .a(tc_a[9]) );
    inv_1 U271 ( .x(n371), .a(tc_a_60) );
    inv_1 U272 ( .x(n446), .a(n364) );
    nor2_1 U273 ( .x(complb1), .a(n190), .b(n191) );
    nor2_1 U274 ( .x(complw1), .a(n180), .b(n181) );
    nand3i_1 U276 ( .x(n190), .a(n441), .b(n447), .c(n469) );
    and4_1 U277 ( .x(n5), .a(n3), .b(n4), .c(n519), .d(n522) );
    inv_1 U216 ( .x(n3), .a(n520) );
    inv_1 U217 ( .x(n4), .a(n523) );
    inv_1 U428 ( .x(n525), .a(n5) );
    nor2_1 U278 ( .x(n447), .a(n448), .b(n445) );
    nor2_1 U279 ( .x(n469), .a(n467), .b(n461) );
    nand2_1 U280 ( .x(n370), .a(n371), .b(n372) );
    nand3i_1 U281 ( .x(n448), .a(n454), .b(n449), .c(n451) );
    nand3i_1 U282 ( .x(n461), .a(n462), .b(n455), .c(n458) );
    nand3i_1 U283 ( .x(n467), .a(n468), .b(n463), .c(n464) );
    inv_1 U284 ( .x(n382), .a(n273) );
    inv_1 U285 ( .x(n384), .a(n268) );
    inv_1 U286 ( .x(n385), .a(n265) );
    inv_1 U287 ( .x(n376), .a(n284) );
    inv_1 U288 ( .x(n377), .a(n282) );
    inv_1 U289 ( .x(n378), .a(n279) );
    inv_1 U290 ( .x(n379), .a(n276) );
    inv_1 U291 ( .x(n396), .a(n248) );
    inv_1 U292 ( .x(n398), .a(n245) );
    inv_1 U293 ( .x(n399), .a(n242) );
    inv_1 U294 ( .x(n389), .a(n262) );
    inv_1 U295 ( .x(n390), .a(n259) );
    inv_1 U296 ( .x(n392), .a(n256) );
    inv_1 U297 ( .x(n393), .a(n253) );
    inv_1 U298 ( .x(n409), .a(n228) );
    inv_1 U299 ( .x(n410), .a(n225) );
    inv_1 U300 ( .x(n412), .a(n222) );
    inv_1 U301 ( .x(n403), .a(n239) );
    inv_1 U302 ( .x(n405), .a(n234) );
    inv_1 U303 ( .x(n406), .a(n231) );
    inv_1 U304 ( .x(n423), .a(n205) );
    inv_1 U305 ( .x(n426), .a(n199) );
    inv_1 U306 ( .x(n417), .a(n214) );
    inv_1 U307 ( .x(n419), .a(n211) );
    inv_1 U308 ( .x(n420), .a(n208) );
    inv_1 U309 ( .x(n444), .a(n361) );
    inv_1 U310 ( .x(n524), .a(n370) );
    inv_1 U311 ( .x(n450), .a(n356) );
    nand2_1 U312 ( .x(n521), .a(n443), .b(n440) );
    inv_1 U313 ( .x(n372), .a(tc_a[28]) );
    nor2_1 U314 ( .x(n451), .a(n452), .b(n453) );
    nor2_1 U315 ( .x(n458), .a(n459), .b(n460) );
    inv_1 U316 ( .x(n468), .a(n331) );
    nor2_1 U317 ( .x(n464), .a(n465), .b(n466) );
    inv_1 U318 ( .x(n494), .a(n295) );
    nand2_1 U319 ( .x(n273), .a(n274), .b(n275) );
    nand2_1 U320 ( .x(n279), .a(n280), .b(n281) );
    nand2_1 U321 ( .x(n276), .a(n277), .b(n278) );
    nand2_1 U322 ( .x(n262), .a(n263), .b(n264) );
    nand2_1 U323 ( .x(n259), .a(n260), .b(n261) );
    nand2_1 U324 ( .x(n256), .a(n257), .b(n258) );
    nand2_1 U325 ( .x(n253), .a(n254), .b(n255) );
    nand2_1 U326 ( .x(n228), .a(n229), .b(n230) );
    nand2_1 U327 ( .x(n225), .a(n226), .b(n227) );
    nand2_1 U328 ( .x(n219), .a(n220), .b(n221) );
    nand2_1 U329 ( .x(n239), .a(n240), .b(n241) );
    nand2_1 U330 ( .x(n202), .a(n203), .b(n204) );
    nand2_1 U331 ( .x(n196), .a(n197), .b(n198) );
    nor2_1 U332 ( .x(n391), .a(n392), .b(n393) );
    nor2_1 U333 ( .x(n388), .a(n389), .b(n390) );
    nor2_1 U334 ( .x(n381), .a(n382), .b(n126) );
    nor2_1 U335 ( .x(n402), .a(n403), .b(n124) );
    nor2_1 U336 ( .x(n408), .a(n409), .b(n410) );
    inv_1 U337 ( .x(n459), .a(n341) );
    inv_1 U338 ( .x(n465), .a(n328) );
    inv_1 U339 ( .x(n466), .a(n325) );
    inv_1 U340 ( .x(n460), .a(n338) );
    nand2_1 U341 ( .x(n361), .a(n362), .b(n363) );
    nand2_1 U342 ( .x(n373), .a(n374), .b(n375) );
    nand2_1 U343 ( .x(n356), .a(n358), .b(n357) );
    inv_1 U344 ( .x(n452), .a(n352) );
    inv_1 U345 ( .x(n484), .a(n299) );
    inv_1 U346 ( .x(n489), .a(n289) );
    inv_1 U347 ( .x(n492), .a(n286) );
    inv_1 U348 ( .x(n490), .a(n292) );
    inv_1 U349 ( .x(n473), .a(n317) );
    inv_1 U350 ( .x(n471), .a(n322) );
    inv_1 U351 ( .x(n482), .a(n306) );
    inv_1 U352 ( .x(n476), .a(n314) );
    nand2_1 U353 ( .x(n367), .a(n368), .b(n369) );
    nand2_1 U354 ( .x(n331), .a(n332), .b(n333) );
    nand2_1 U355 ( .x(n302), .a(n303), .b(n304) );
    nand2_1 U356 ( .x(n295), .a(n296), .b(n297) );
    inv_1 U357 ( .x(n275), .a(tc_wd_56) );
    inv_1 U358 ( .x(n285), .a(tc_wd_63) );
    inv_1 U359 ( .x(n283), .a(tc_wd_60) );
    inv_1 U360 ( .x(n281), .a(tc_wd_61) );
    inv_1 U361 ( .x(n278), .a(tc_wd_59) );
    inv_1 U362 ( .x(n264), .a(tc_wd_53) );
    inv_1 U363 ( .x(n261), .a(tc_wd_51) );
    inv_1 U364 ( .x(n258), .a(tc_wd_48) );
    inv_1 U365 ( .x(n254), .a(tc_wd[17]) );
    inv_1 U366 ( .x(n255), .a(tc_wd_49) );
    inv_1 U367 ( .x(n230), .a(tc_wd[37]) );
    inv_1 U368 ( .x(n227), .a(tc_wd[35]) );
    inv_1 U369 ( .x(n221), .a(tc_wd[33]) );
    inv_1 U370 ( .x(n241), .a(tc_wd_40) );
    inv_1 U371 ( .x(n204), .a(tc_wd[42]) );
    inv_1 U372 ( .x(n198), .a(tc_wd[34]) );
    nand2_1 U373 ( .x(n341), .a(n342), .b(n343) );
    nand2_1 U374 ( .x(n345), .a(n347), .b(n346) );
    nand2_1 U375 ( .x(n328), .a(n329), .b(n330) );
    nand2_1 U376 ( .x(n325), .a(n326), .b(n327) );
    nand2_1 U377 ( .x(n338), .a(n340), .b(n339) );
    inv_1 U378 ( .x(n362), .a(tc_a[24]) );
    inv_1 U379 ( .x(n363), .a(tc_a[56]) );
    inv_1 U380 ( .x(n357), .a(tc_a[22]) );
    inv_1 U381 ( .x(n358), .a(tc_a[54]) );
    nand2_1 U382 ( .x(n352), .a(n353), .b(n354) );
    nand2_1 U383 ( .x(n299), .a(n300), .b(n301) );
    nand2_1 U384 ( .x(n289), .a(n290), .b(n291) );
    nand2_1 U385 ( .x(n286), .a(n287), .b(n288) );
    nand2_1 U386 ( .x(n292), .a(n293), .b(n294) );
    nand2_1 U387 ( .x(n317), .a(n318), .b(n319) );
    nand2_1 U388 ( .x(n322), .a(n323), .b(n324) );
    nand2_1 U389 ( .x(n306), .a(n307), .b(n308) );
    nand2_1 U390 ( .x(n314), .a(n315), .b(n316) );
    inv_1 U391 ( .x(n332), .a(tc_a[4]) );
    inv_1 U392 ( .x(n333), .a(tc_a[36]) );
    inv_1 U393 ( .x(n296), .a(tc_a[31]) );
    inv_1 U394 ( .x(n342), .a(tc_itag[2]) );
    inv_1 U395 ( .x(n343), .a(tc_itag[7]) );
    inv_1 U396 ( .x(n346), .a(tc_a[15]) );
    inv_1 U397 ( .x(n347), .a(tc_a[47]) );
    inv_1 U398 ( .x(n329), .a(tc_a[2]) );
    inv_1 U399 ( .x(n330), .a(tc_a[34]) );
    inv_1 U400 ( .x(n326), .a(tc_a[5]) );
    inv_1 U401 ( .x(n327), .a(tc_a[37]) );
    inv_1 U402 ( .x(n337), .a(tc_a[62]) );
    inv_1 U403 ( .x(n339), .a(tc_lock[0]) );
    inv_1 U404 ( .x(n340), .a(tc_lock[1]) );
    inv_1 U405 ( .x(n353), .a(tc_a[13]) );
    inv_1 U406 ( .x(n354), .a(tc_a[45]) );
    inv_1 U407 ( .x(n300), .a(tc_a[1]) );
    inv_1 U408 ( .x(n290), .a(tc_a[10]) );
    inv_1 U409 ( .x(n291), .a(tc_a[42]) );
    inv_1 U410 ( .x(n287), .a(tc_seq[0]) );
    inv_1 U411 ( .x(n288), .a(tc_seq[1]) );
    inv_1 U412 ( .x(n293), .a(tc_a[23]) );
    inv_1 U413 ( .x(n294), .a(tc_a[55]) );
    inv_1 U414 ( .x(n318), .a(tc_a[19]) );
    inv_1 U415 ( .x(n323), .a(tc_a[0]) );
    inv_1 U416 ( .x(n307), .a(tc_a[25]) );
    inv_1 U417 ( .x(n308), .a(tc_a[57]) );
    buf_1 U418 ( .x(we_i), .a(tc_rnw[0]) );
    matched_delay_cp2slave_resp_wb U419 ( .x(req_out_delayed), .a(req_out) );
    and4_1 U420 ( .x(_25_net_), .a(sel_o[0]), .b(sel_o[1]), .c(n529), .d(n530)
         );
    inv_1 U421 ( .x(_24_net_), .a(we_i) );
    and2_1 U422 ( .x(tc_defer), .a(rty_o), .b(respond) );
    and4_1 U423 ( .x(_26_net_), .a(sel_o[0]), .b(sel_o[1]), .c(sel_o[3]), .d(
        sel_o[2]) );
    inv_1 U424 ( .x(n532), .a(acc_o) );
    inv_1 U425 ( .x(n531), .a(rty_o) );
    inv_1 U426 ( .x(n529), .a(sel_o[2]) );
    inv_1 U427 ( .x(n530), .a(sel_o[3]) );
    buf_1 U150 ( .x(n142), .a(req_in_i) );
    matched_delay_cp2slave_com_wb matchDelCom ( .x(req_in), .a(req_in_i) );
    nand2_1 U275 ( .x(req_in_i), .a(n186), .b(n187) );
    inv_1 U221 ( .x(n186), .a(all_w) );
    inv_1 U269 ( .x(n187), .a(all_r) );
    dffp_1 mult_i_reg ( .q(mult_i), .d(n137), .ck(n142) );
    ao222_1 \cg_respond/__tmp99/U1  ( .x(respond), .a(req_out), .b(tc_ack), 
        .c(req_out), .d(respond), .e(tc_ack), .f(respond) );
    oa21_1 \cg_all_r/__tmp99/U1  ( .x(all_r), .a(tc_rnw[1]), .b(all_r), .c(
        comp_basic) );
    ao31_1 \cg_all_w/__tmp99/aoi  ( .x(\cg_all_w/__tmp99/loop ), .a(comp_basic
        ), .b(comp_wd), .c(we_i), .d(all_w) );
    oa21_1 \cg_all_w/__tmp99/outGate  ( .x(all_w), .a(comp_basic), .b(comp_wd), 
        .c(\cg_all_w/__tmp99/loop ) );
    ao222_1 \cg_wd/__tmp99/U1  ( .x(comp_wd), .a(complw0), .b(complw1), .c(
        complw0), .d(comp_wd), .e(complw1), .f(comp_wd) );
    ao222_1 \cg_basic/__tmp99/U1  ( .x(comp_basic), .a(complb0), .b(complb1), 
        .c(complb0), .d(comp_basic), .e(complb1), .f(comp_basic) );
    inv_1 \Usze1/Uii  ( .x(\Usze1/ni ), .a(_26_net_) );
    inv_1 \Usze1/Uih  ( .x(\Usze1/nh ), .a(tr_size[3]) );
    inv_1 \Usze1/Uil  ( .x(\Usze1/nl ), .a(tr_size[1]) );
    ao23_1 \Usze1/Ucl/U1/U1  ( .x(tr_size[1]), .a(n2), .b(tr_size[1]), .c(n1), 
        .d(\Usze1/ni ), .e(\Usze1/nh ) );
    ao23_1 \Usze1/Uch/U1/U1  ( .x(tr_size[3]), .a(n1), .b(tr_size[3]), .c(n1), 
        .d(_26_net_), .e(\Usze1/nl ) );
    inv_1 \Usze0/Uii  ( .x(\Usze0/ni ), .a(_25_net_) );
    inv_1 \Usze0/Uih  ( .x(\Usze0/nh ), .a(tr_size[2]) );
    inv_1 \Usze0/Uil  ( .x(\Usze0/nl ), .a(tr_size[0]) );
    ao23_1 \Usze0/Ucl/U1/U1  ( .x(tr_size[0]), .a(n2), .b(tr_size[0]), .c(n1), 
        .d(\Usze0/ni ), .e(\Usze0/nh ) );
    ao23_1 \Usze0/Uch/U1/U1  ( .x(tr_size[2]), .a(n2), .b(tr_size[2]), .c(n1), 
        .d(_25_net_), .e(\Usze0/nl ) );
    inv_1 \Urnw/Uii  ( .x(\Urnw/ni ), .a(_24_net_) );
    inv_1 \Urnw/Uih  ( .x(\Urnw/nh ), .a(tr_rnw[1]) );
    inv_1 \Urnw/Uil  ( .x(\Urnw/nl ), .a(tr_rnw[0]) );
    ao23_1 \Urnw/Ucl/U1/U1  ( .x(tr_rnw[0]), .a(n1), .b(tr_rnw[0]), .c(n1), 
        .d(\Urnw/ni ), .e(\Urnw/nh ) );
    ao23_1 \Urnw/Uch/U1/U1  ( .x(tr_rnw[1]), .a(n1), .b(tr_rnw[1]), .c(n1), 
        .d(_24_net_), .e(\Urnw/nl ) );
    inv_1 \Uerr/Uii  ( .x(\Uerr/ni ), .a(err_o) );
    inv_1 \Uerr/Uih  ( .x(\Uerr/nh ), .a(tr_err[1]) );
    inv_1 \Uerr/Uil  ( .x(\Uerr/nl ), .a(tr_err[0]) );
    ao23_1 \Uerr/Ucl/U1/U1  ( .x(tr_err[0]), .a(n1), .b(tr_err[0]), .c(n1), 
        .d(\Uerr/ni ), .e(\Uerr/nh ) );
    ao23_1 \Uerr/Uch/U1/U1  ( .x(tr_err[1]), .a(n1), .b(tr_err[1]), .c(n1), 
        .d(err_o), .e(\Uerr/nl ) );
    inv_0 U1 ( .x(n298), .a(tc_itag[6]) );
    nor2_0 U2 ( .x(n485), .a(tc_itag[1]), .b(tc_itag[6]) );
    inv_0 U4 ( .x(n344), .a(tc_itag[8]) );
    nor2_0 U8 ( .x(n462), .a(tc_itag[3]), .b(tc_itag[8]) );
    nor2_0 U92 ( .x(n496), .a(tc_size[0]), .b(tc_size[1]) );
    nor2_0 U93 ( .x(n194), .a(tc_size[0]), .b(tc_size[2]) );
    buf_16 U104 ( .x(n1), .a(req_out_delayed) );
    buf_16 U111 ( .x(n2), .a(req_out_delayed) );
endmodule


module slave_if_wb ( nReset, sc_req, sc_we, sc_mult, sc_seq, sc_prd, sc_ts, 
    sc_st, sc_sel, sc_adr, sc_dat, sc_ack, sr_req, sr_err, sr_rty, sr_acc, 
    sr_mult, sr_ts, sr_rt, sr_sel, sr_dat, sr_ack, chaincommand, 
    nchaincommandack, chainresponse, nchainresponseack, e_dp, e_ip, e_tic, 
    r_dp, r_ip, r_tic );
output [2:0] sc_ts;
output [4:0] sc_st;
output [3:0] sc_sel;
output [31:0] sc_adr;
output [31:0] sc_dat;
input  [2:0] sr_ts;
input  [4:0] sr_rt;
input  [3:0] sr_sel;
input  [31:0] sr_dat;
input  [4:0] chaincommand;
output [4:0] chainresponse;
input  [2:0] e_dp;
input  [2:0] e_ip;
input  [2:0] e_tic;
input  [2:0] r_dp;
input  [2:0] r_ip;
input  [2:0] r_tic;
input  nReset, sc_ack, sr_req, sr_err, sr_rty, sr_acc, sr_mult, 
    nchainresponseack;
output sc_req, sc_we, sc_mult, sc_seq, sc_prd, sr_ack, nchaincommandack;
    wire nroute_ack, rt_ack, routetx_req, ct_ack, ct_defer, ct_slow, ct_ok, 
        routetx_ack, \route[4] , \route[1] , \route[0] , \rt_rd[63] , 
        \rt_rd[62] , \rt_rd[61] , \rt_rd[60] , \rt_rd[59] , \rt_rd[58] , 
        \rt_rd[57] , \rt_rd[56] , \rt_rd[55] , \rt_rd[54] , \rt_rd[53] , 
        \rt_rd[52] , \rt_rd[51] , \rt_rd[50] , \rt_rd[49] , \rt_rd[48] , 
        \rt_rd[47] , \rt_rd[46] , \rt_rd[45] , \rt_rd[44] , \rt_rd[43] , 
        \rt_rd[42] , \rt_rd[41] , \rt_rd[40] , \rt_rd[39] , \rt_rd[38] , 
        \rt_rd[37] , \rt_rd[36] , \rt_rd[35] , \rt_rd[34] , \rt_rd[33] , 
        \rt_rd[32] , \rt_rd[31] , \rt_rd[30] , \rt_rd[29] , \rt_rd[28] , 
        \rt_rd[27] , \rt_rd[26] , \rt_rd[25] , \rt_rd[24] , \rt_rd[23] , 
        \rt_rd[22] , \rt_rd[21] , \rt_rd[20] , \rt_rd[19] , \rt_rd[18] , 
        \rt_rd[17] , \rt_rd[16] , \rt_rd[15] , \rt_rd[14] , \rt_rd[13] , 
        \rt_rd[12] , \rt_rd[11] , \rt_rd[10] , \rt_rd[9] , \rt_rd[8] , 
        \rt_rd[7] , \rt_rd[6] , \rt_rd[5] , \rt_rd[4] , \rt_rd[3] , \rt_rd[2] , 
        \rt_rd[1] , \rt_rd[0] , \rt_err[1] , \rt_err[0] , \ct_wd[63] , 
        \ct_wd[62] , \ct_wd[61] , \ct_wd[60] , \ct_wd[59] , \ct_wd[58] , 
        \ct_wd[57] , \ct_wd[56] , \ct_wd[55] , \ct_wd[54] , \ct_wd[53] , 
        \ct_wd[52] , \ct_wd[51] , \ct_wd[50] , \ct_wd[49] , \ct_wd[48] , 
        \ct_wd[47] , \ct_wd[46] , \ct_wd[45] , \ct_wd[44] , \ct_wd[43] , 
        \ct_wd[42] , \ct_wd[41] , \ct_wd[40] , \ct_wd[39] , \ct_wd[38] , 
        \ct_wd[37] , \ct_wd[36] , \ct_wd[35] , \ct_wd[34] , \ct_wd[33] , 
        \ct_wd[32] , \ct_wd[31] , \ct_wd[30] , \ct_wd[29] , \ct_wd[28] , 
        \ct_wd[27] , \ct_wd[26] , \ct_wd[25] , \ct_wd[24] , \ct_wd[23] , 
        \ct_wd[22] , \ct_wd[21] , \ct_wd[20] , \ct_wd[19] , \ct_wd[18] , 
        \ct_wd[17] , \ct_wd[16] , \ct_wd[15] , \ct_wd[14] , \ct_wd[13] , 
        \ct_wd[12] , \ct_wd[11] , \ct_wd[10] , \ct_wd[9] , \ct_wd[8] , 
        \ct_wd[7] , \ct_wd[6] , \ct_wd[5] , \ct_wd[4] , \ct_wd[3] , \ct_wd[2] , 
        \ct_wd[1] , \ct_wd[0] , \tag_l[4] , \tag_l[3] , \tag_l[2] , \tag_l[1] , 
        \tag_l[0] , \tag_h[4] , \tag_h[3] , \tag_h[2] , \tag_h[1] , \tag_h[0] , 
        \ct_seq[1] , \ct_seq[0] , \ct_lock[1] , \ct_lock[0] , \ct_itag[9] , 
        \ct_itag[8] , \ct_itag[7] , \ct_itag[6] , \ct_itag[5] , \ct_itag[4] , 
        \ct_itag[3] , \ct_itag[2] , \ct_itag[1] , \ct_itag[0] , \ct_size[3] , 
        \ct_size[2] , \ct_size[1] , \ct_size[0] , \ct_rnw[1] , \ct_rnw[0] , 
        \ct_a[63] , \ct_a[62] , \ct_a[61] , \ct_a[60] , \ct_a[59] , \ct_a[58] , 
        \ct_a[57] , \ct_a[56] , \ct_a[55] , \ct_a[54] , \ct_a[53] , \ct_a[52] , 
        \ct_a[51] , \ct_a[50] , \ct_a[49] , \ct_a[48] , \ct_a[47] , \ct_a[46] , 
        \ct_a[45] , \ct_a[44] , \ct_a[43] , \ct_a[42] , \ct_a[41] , \ct_a[40] , 
        \ct_a[39] , \ct_a[38] , \ct_a[37] , \ct_a[36] , \ct_a[35] , \ct_a[34] , 
        \ct_a[33] , \ct_a[32] , \ct_a[31] , \ct_a[30] , \ct_a[29] , \ct_a[28] , 
        \ct_a[27] , \ct_a[26] , \ct_a[25] , \ct_a[24] , \ct_a[23] , \ct_a[22] , 
        \ct_a[21] , \ct_a[20] , \ct_a[19] , \ct_a[18] , \ct_a[17] , \ct_a[16] , 
        \ct_a[15] , \ct_a[14] , \ct_a[13] , \ct_a[12] , \ct_a[11] , \ct_a[10] , 
        \ct_a[9] , \ct_a[8] , \ct_a[7] , \ct_a[6] , \ct_a[5] , \ct_a[4] , 
        \ct_a[3] , \ct_a[2] , \ct_a[1] , \ct_a[0] , \rl[2] , \rl[1] , \rl[0] , 
        \rh[2] , \rh[1] , SYNOPSYS_UNCONNECTED_2, \el[2] , \el[1] , \el[0] , 
        SYNOPSYS_UNCONNECTED_1, \eh[1] , \eh[0] , SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4, reset, SYNOPSYS_UNCONNECTED_5;
    assign sc_prd = 1'b0;
    assign sc_ts[2] = 1'b0;
    assign sc_ts[1] = 1'b0;
    assign sc_ts[0] = 1'b0;
    assign sc_sel[0] = 1'b1;
    target_wb tg ( .addr({\ct_a[63] , \ct_a[62] , \ct_a[61] , \ct_a[60] , 
        \ct_a[59] , \ct_a[58] , \ct_a[57] , \ct_a[56] , \ct_a[55] , \ct_a[54] , 
        \ct_a[53] , \ct_a[52] , \ct_a[51] , \ct_a[50] , \ct_a[49] , \ct_a[48] , 
        \ct_a[47] , \ct_a[46] , \ct_a[45] , \ct_a[44] , \ct_a[43] , \ct_a[42] , 
        \ct_a[41] , \ct_a[40] , \ct_a[39] , \ct_a[38] , \ct_a[37] , \ct_a[36] , 
        \ct_a[35] , \ct_a[34] , \ct_a[33] , \ct_a[32] , \ct_a[31] , \ct_a[30] , 
        \ct_a[29] , \ct_a[28] , \ct_a[27] , \ct_a[26] , \ct_a[25] , \ct_a[24] , 
        \ct_a[23] , \ct_a[22] , \ct_a[21] , \ct_a[20] , \ct_a[19] , \ct_a[18] , 
        \ct_a[17] , \ct_a[16] , \ct_a[15] , \ct_a[14] , \ct_a[13] , \ct_a[12] , 
        \ct_a[11] , \ct_a[10] , \ct_a[9] , \ct_a[8] , \ct_a[7] , \ct_a[6] , 
        \ct_a[5] , \ct_a[4] , \ct_a[3] , \ct_a[2] , \ct_a[1] , \ct_a[0] }), 
        .chainresponse(chainresponse), .crnw({\ct_rnw[1] , \ct_rnw[0] }), 
        .csize({\ct_size[3] , \ct_size[2] , \ct_size[1] , \ct_size[0] }), 
        .ctag({\ct_itag[9] , \ct_itag[8] , \ct_itag[7] , \ct_itag[6] , 
        \ct_itag[5] , \ct_itag[4] , \ct_itag[3] , \ct_itag[2] , \ct_itag[1] , 
        \ct_itag[0] }), .lock({\ct_lock[1] , \ct_lock[0] }), 
        .nchaincommandack(nchaincommandack), .nrouteack(nroute_ack), .rack(
        rt_ack), .routetxreq(routetx_req), .seq({\ct_seq[1] , \ct_seq[0] }), 
        .tag_h({\tag_h[4] , \tag_h[3] , \tag_h[2] , \tag_h[1] , \tag_h[0] }), 
        .tag_l({\tag_l[4] , \tag_l[3] , \tag_l[2] , \tag_l[1] , \tag_l[0] }), 
        .wd({\ct_wd[63] , \ct_wd[62] , \ct_wd[61] , \ct_wd[60] , \ct_wd[59] , 
        \ct_wd[58] , \ct_wd[57] , \ct_wd[56] , \ct_wd[55] , \ct_wd[54] , 
        \ct_wd[53] , \ct_wd[52] , \ct_wd[51] , \ct_wd[50] , \ct_wd[49] , 
        \ct_wd[48] , \ct_wd[47] , \ct_wd[46] , \ct_wd[45] , \ct_wd[44] , 
        \ct_wd[43] , \ct_wd[42] , \ct_wd[41] , \ct_wd[40] , \ct_wd[39] , 
        \ct_wd[38] , \ct_wd[37] , \ct_wd[36] , \ct_wd[35] , \ct_wd[34] , 
        \ct_wd[33] , \ct_wd[32] , \ct_wd[31] , \ct_wd[30] , \ct_wd[29] , 
        \ct_wd[28] , \ct_wd[27] , \ct_wd[26] , \ct_wd[25] , \ct_wd[24] , 
        \ct_wd[23] , \ct_wd[22] , \ct_wd[21] , \ct_wd[20] , \ct_wd[19] , 
        \ct_wd[18] , \ct_wd[17] , \ct_wd[16] , \ct_wd[15] , \ct_wd[14] , 
        \ct_wd[13] , \ct_wd[12] , \ct_wd[11] , \ct_wd[10] , \ct_wd[9] , 
        \ct_wd[8] , \ct_wd[7] , \ct_wd[6] , \ct_wd[5] , \ct_wd[4] , \ct_wd[3] , 
        \ct_wd[2] , \ct_wd[1] , \ct_wd[0] }), .cack(ct_ack), .cdefer(ct_defer), 
        .chaincommand(chaincommand), .cndefer(ct_slow), .cok(ct_ok), .err({
        \rt_err[1] , \rt_err[0] }), .nReset(nReset), .nchainresponseack(
        nchainresponseack), .rd({\rt_rd[63] , \rt_rd[62] , \rt_rd[61] , 
        \rt_rd[60] , \rt_rd[59] , \rt_rd[58] , \rt_rd[57] , \rt_rd[56] , 
        \rt_rd[55] , \rt_rd[54] , \rt_rd[53] , \rt_rd[52] , \rt_rd[51] , 
        \rt_rd[50] , \rt_rd[49] , \rt_rd[48] , \rt_rd[47] , \rt_rd[46] , 
        \rt_rd[45] , \rt_rd[44] , \rt_rd[43] , \rt_rd[42] , \rt_rd[41] , 
        \rt_rd[40] , \rt_rd[39] , \rt_rd[38] , \rt_rd[37] , \rt_rd[36] , 
        \rt_rd[35] , \rt_rd[34] , \rt_rd[33] , \rt_rd[32] , \rt_rd[31] , 
        \rt_rd[30] , \rt_rd[29] , \rt_rd[28] , \rt_rd[27] , \rt_rd[26] , 
        \rt_rd[25] , \rt_rd[24] , \rt_rd[23] , \rt_rd[22] , \rt_rd[21] , 
        \rt_rd[20] , \rt_rd[19] , \rt_rd[18] , \rt_rd[17] , \rt_rd[16] , 
        \rt_rd[15] , \rt_rd[14] , \rt_rd[13] , \rt_rd[12] , \rt_rd[11] , 
        \rt_rd[10] , \rt_rd[9] , \rt_rd[8] , \rt_rd[7] , \rt_rd[6] , 
        \rt_rd[5] , \rt_rd[4] , \rt_rd[3] , \rt_rd[2] , \rt_rd[1] , \rt_rd[0] 
        }), .route({\route[4] , 1'b0, 1'b0, \route[1] , \route[0] }), 
        .routetxack(routetx_ack) );
    t_adec_wb dec ( .e_h({SYNOPSYS_UNCONNECTED_1, \eh[1] , \eh[0] }), .e_l({
        \el[2] , \el[1] , \el[0] }), .r_h({\rh[2] , \rh[1] , 
        SYNOPSYS_UNCONNECTED_2}), .r_l({\rl[2] , \rl[1] , \rl[0] }), .e_dp(
        e_dp), .e_ip(e_ip), .e_tic(e_tic), .r_dp(r_dp), .r_ip(r_ip), .r_tic(
        r_tic), .tag_h({\tag_h[4] , \tag_h[3] , \tag_h[2] , \tag_h[1] , 
        \tag_h[0] }), .tag_l({\tag_l[4] , \tag_l[3] , \tag_l[2] , \tag_l[1] , 
        \tag_l[0] }) );
    resp_route_tx_wb rt ( .o({\route[4] , SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4, \route[1] , \route[0] }), .rtxack(routetx_ack), 
        .e_h({1'b0, \eh[1] , \eh[0] }), .e_l({\el[2] , \el[1] , \el[0] }), 
        .noa(nroute_ack), .r_h({\rh[2] , \rh[1] , 1'b0}), .r_l({\rl[2] , 
        \rl[1] , \rl[0] }), .rtxreq(routetx_req) );
    inv_2 U1 ( .x(reset), .a(nReset) );
    cp2slave_wb chainif2slave ( .tc_seq({\ct_seq[1] , \ct_seq[0] }), .tc_size(
        {\ct_size[3] , \ct_size[2] , \ct_size[1] , \ct_size[0] }), .tc_itag({
        \ct_itag[9] , \ct_itag[8] , \ct_itag[7] , \ct_itag[6] , \ct_itag[5] , 
        \ct_itag[4] , \ct_itag[3] , \ct_itag[2] , \ct_itag[1] , \ct_itag[0] }), 
        .tc_wd({\ct_wd[63] , \ct_wd[62] , \ct_wd[61] , \ct_wd[60] , 
        \ct_wd[59] , \ct_wd[58] , \ct_wd[57] , \ct_wd[56] , \ct_wd[55] , 
        \ct_wd[54] , \ct_wd[53] , \ct_wd[52] , \ct_wd[51] , \ct_wd[50] , 
        \ct_wd[49] , \ct_wd[48] , \ct_wd[47] , \ct_wd[46] , \ct_wd[45] , 
        \ct_wd[44] , \ct_wd[43] , \ct_wd[42] , \ct_wd[41] , \ct_wd[40] , 
        \ct_wd[39] , \ct_wd[38] , \ct_wd[37] , \ct_wd[36] , \ct_wd[35] , 
        \ct_wd[34] , \ct_wd[33] , \ct_wd[32] , \ct_wd[31] , \ct_wd[30] , 
        \ct_wd[29] , \ct_wd[28] , \ct_wd[27] , \ct_wd[26] , \ct_wd[25] , 
        \ct_wd[24] , \ct_wd[23] , \ct_wd[22] , \ct_wd[21] , \ct_wd[20] , 
        \ct_wd[19] , \ct_wd[18] , \ct_wd[17] , \ct_wd[16] , \ct_wd[15] , 
        \ct_wd[14] , \ct_wd[13] , \ct_wd[12] , \ct_wd[11] , \ct_wd[10] , 
        \ct_wd[9] , \ct_wd[8] , \ct_wd[7] , \ct_wd[6] , \ct_wd[5] , \ct_wd[4] , 
        \ct_wd[3] , \ct_wd[2] , \ct_wd[1] , \ct_wd[0] }), .tc_lock({
        \ct_lock[1] , \ct_lock[0] }), .tc_a({\ct_a[63] , \ct_a[62] , 
        \ct_a[61] , \ct_a[60] , \ct_a[59] , \ct_a[58] , \ct_a[57] , \ct_a[56] , 
        \ct_a[55] , \ct_a[54] , \ct_a[53] , \ct_a[52] , \ct_a[51] , \ct_a[50] , 
        \ct_a[49] , \ct_a[48] , \ct_a[47] , \ct_a[46] , \ct_a[45] , \ct_a[44] , 
        \ct_a[43] , \ct_a[42] , \ct_a[41] , \ct_a[40] , \ct_a[39] , \ct_a[38] , 
        \ct_a[37] , \ct_a[36] , \ct_a[35] , \ct_a[34] , \ct_a[33] , \ct_a[32] , 
        \ct_a[31] , \ct_a[30] , \ct_a[29] , \ct_a[28] , \ct_a[27] , \ct_a[26] , 
        \ct_a[25] , \ct_a[24] , \ct_a[23] , \ct_a[22] , \ct_a[21] , \ct_a[20] , 
        \ct_a[19] , \ct_a[18] , \ct_a[17] , \ct_a[16] , \ct_a[15] , \ct_a[14] , 
        \ct_a[13] , \ct_a[12] , \ct_a[11] , \ct_a[10] , \ct_a[9] , \ct_a[8] , 
        \ct_a[7] , \ct_a[6] , \ct_a[5] , \ct_a[4] , \ct_a[3] , \ct_a[2] , 
        \ct_a[1] , \ct_a[0] }), .tc_rnw({\ct_rnw[1] , \ct_rnw[0] }), .tc_ok(
        ct_ok), .tc_defer(ct_defer), .tc_slow(ct_slow), .tc_ack(ct_ack), 
        .req_in(sc_req), .st_i(sc_st), .we_i(sc_we), .mult_i(sc_mult), .adr_i(
        sc_adr), .dat_i(sc_dat), .seq_i(sc_seq), .sel_i({sc_sel[3], sc_sel[2], 
        sc_sel[1], SYNOPSYS_UNCONNECTED_5}), .ack_in(sc_ack), .tr_rd({
        \rt_rd[63] , \rt_rd[62] , \rt_rd[61] , \rt_rd[60] , \rt_rd[59] , 
        \rt_rd[58] , \rt_rd[57] , \rt_rd[56] , \rt_rd[55] , \rt_rd[54] , 
        \rt_rd[53] , \rt_rd[52] , \rt_rd[51] , \rt_rd[50] , \rt_rd[49] , 
        \rt_rd[48] , \rt_rd[47] , \rt_rd[46] , \rt_rd[45] , \rt_rd[44] , 
        \rt_rd[43] , \rt_rd[42] , \rt_rd[41] , \rt_rd[40] , \rt_rd[39] , 
        \rt_rd[38] , \rt_rd[37] , \rt_rd[36] , \rt_rd[35] , \rt_rd[34] , 
        \rt_rd[33] , \rt_rd[32] , \rt_rd[31] , \rt_rd[30] , \rt_rd[29] , 
        \rt_rd[28] , \rt_rd[27] , \rt_rd[26] , \rt_rd[25] , \rt_rd[24] , 
        \rt_rd[23] , \rt_rd[22] , \rt_rd[21] , \rt_rd[20] , \rt_rd[19] , 
        \rt_rd[18] , \rt_rd[17] , \rt_rd[16] , \rt_rd[15] , \rt_rd[14] , 
        \rt_rd[13] , \rt_rd[12] , \rt_rd[11] , \rt_rd[10] , \rt_rd[9] , 
        \rt_rd[8] , \rt_rd[7] , \rt_rd[6] , \rt_rd[5] , \rt_rd[4] , \rt_rd[3] , 
        \rt_rd[2] , \rt_rd[1] , \rt_rd[0] }), .tr_err({\rt_err[1] , 
        \rt_err[0] }), .tr_ack(rt_ack), .req_out(sr_req), .dat_o(sr_dat), 
        .err_o(sr_err), .rty_o(sr_rty), .acc_o(sr_acc), .sel_o(sr_sel), 
        .mult_o(sr_mult), .rt_o(sr_rt), .ack_out(sr_ack), .reset(reset) );
endmodule


module wishbone ( reset_b, clk, ch_we_i, ch_dat_i, ch_adr_i, ch_req_i, 
    ch_ack_i, ch_req_o, ch_dat_o, ch_ack_o, wb_we_o, wb_stb_cyc_o, wb_dat_o, 
    wb_adr_o, wb_dat_i, wb_ack_i );
input  [31:0] ch_dat_i;
input  [11:0] ch_adr_i;
output [31:0] ch_dat_o;
output [31:0] wb_dat_o;
output [11:0] wb_adr_o;
input  [31:0] wb_dat_i;
input  reset_b, clk, ch_we_i, ch_req_i, ch_ack_o, wb_ack_i;
output ch_ack_i, ch_req_o, wb_we_o, wb_stb_cyc_o;
    wire ch_dat_i_31, ch_dat_i_30, ch_dat_i_29, ch_dat_i_28, ch_dat_i_27, 
        ch_dat_i_26, ch_dat_i_25, ch_dat_i_24, ch_dat_i_23, ch_dat_i_22, 
        ch_dat_i_21, ch_dat_i_20, ch_dat_i_19, ch_dat_i_18, ch_dat_i_17, 
        ch_dat_i_16, ch_dat_i_15, ch_dat_i_14, ch_dat_i_13, ch_dat_i_12, 
        ch_dat_i_11, ch_dat_i_10, ch_dat_i_9, ch_dat_i_8, ch_dat_i_7, 
        ch_dat_i_6, ch_dat_i_5, ch_dat_i_4, ch_dat_i_3, ch_dat_i_2, ch_dat_i_1, 
        ch_dat_i_0, ch_adr_i_11, ch_adr_i_10, ch_adr_i_9, ch_adr_i_8, 
        ch_adr_i_7, ch_adr_i_6, ch_adr_i_5, ch_adr_i_4, ch_adr_i_3, ch_adr_i_2, 
        ch_adr_i_1, ch_adr_i_0, n7, n4, n3, \reqoGate/n2 , \reqoGate/nr , 
        \reqoGate/nd , sync_ack_inv, rsync, ch_idle, n5, n2, n6, rin1, 
        sync_ack_l, n1, ch_req_o_wire;
    assign wb_we_o = ch_we_i;
    assign ch_dat_i_31 = ch_dat_i[31];
    assign ch_dat_i_30 = ch_dat_i[30];
    assign ch_dat_i_29 = ch_dat_i[29];
    assign ch_dat_i_28 = ch_dat_i[28];
    assign ch_dat_i_27 = ch_dat_i[27];
    assign ch_dat_i_26 = ch_dat_i[26];
    assign ch_dat_i_25 = ch_dat_i[25];
    assign ch_dat_i_24 = ch_dat_i[24];
    assign ch_dat_i_23 = ch_dat_i[23];
    assign ch_dat_i_22 = ch_dat_i[22];
    assign ch_dat_i_21 = ch_dat_i[21];
    assign ch_dat_i_20 = ch_dat_i[20];
    assign ch_dat_i_19 = ch_dat_i[19];
    assign ch_dat_i_18 = ch_dat_i[18];
    assign ch_dat_i_17 = ch_dat_i[17];
    assign ch_dat_i_16 = ch_dat_i[16];
    assign ch_dat_i_15 = ch_dat_i[15];
    assign ch_dat_i_14 = ch_dat_i[14];
    assign ch_dat_i_13 = ch_dat_i[13];
    assign ch_dat_i_12 = ch_dat_i[12];
    assign ch_dat_i_11 = ch_dat_i[11];
    assign ch_dat_i_10 = ch_dat_i[10];
    assign ch_dat_i_9 = ch_dat_i[9];
    assign ch_dat_i_8 = ch_dat_i[8];
    assign ch_dat_i_7 = ch_dat_i[7];
    assign ch_dat_i_6 = ch_dat_i[6];
    assign ch_dat_i_5 = ch_dat_i[5];
    assign ch_dat_i_4 = ch_dat_i[4];
    assign ch_dat_i_3 = ch_dat_i[3];
    assign ch_dat_i_2 = ch_dat_i[2];
    assign ch_dat_i_1 = ch_dat_i[1];
    assign ch_dat_i_0 = ch_dat_i[0];
    assign ch_adr_i_11 = ch_adr_i[11];
    assign ch_adr_i_10 = ch_adr_i[10];
    assign ch_adr_i_9 = ch_adr_i[9];
    assign ch_adr_i_8 = ch_adr_i[8];
    assign ch_adr_i_7 = ch_adr_i[7];
    assign ch_adr_i_6 = ch_adr_i[6];
    assign ch_adr_i_5 = ch_adr_i[5];
    assign ch_adr_i_4 = ch_adr_i[4];
    assign ch_adr_i_3 = ch_adr_i[3];
    assign ch_adr_i_2 = ch_adr_i[2];
    assign ch_adr_i_1 = ch_adr_i[1];
    assign ch_adr_i_0 = ch_adr_i[0];
    assign ch_req_o = ch_ack_i;
    assign wb_dat_o[31] = ch_dat_i_31;
    assign wb_dat_o[30] = ch_dat_i_30;
    assign wb_dat_o[29] = ch_dat_i_29;
    assign wb_dat_o[28] = ch_dat_i_28;
    assign wb_dat_o[27] = ch_dat_i_27;
    assign wb_dat_o[26] = ch_dat_i_26;
    assign wb_dat_o[25] = ch_dat_i_25;
    assign wb_dat_o[24] = ch_dat_i_24;
    assign wb_dat_o[23] = ch_dat_i_23;
    assign wb_dat_o[22] = ch_dat_i_22;
    assign wb_dat_o[21] = ch_dat_i_21;
    assign wb_dat_o[20] = ch_dat_i_20;
    assign wb_dat_o[19] = ch_dat_i_19;
    assign wb_dat_o[18] = ch_dat_i_18;
    assign wb_dat_o[17] = ch_dat_i_17;
    assign wb_dat_o[16] = ch_dat_i_16;
    assign wb_dat_o[15] = ch_dat_i_15;
    assign wb_dat_o[14] = ch_dat_i_14;
    assign wb_dat_o[13] = ch_dat_i_13;
    assign wb_dat_o[12] = ch_dat_i_12;
    assign wb_dat_o[11] = ch_dat_i_11;
    assign wb_dat_o[10] = ch_dat_i_10;
    assign wb_dat_o[9] = ch_dat_i_9;
    assign wb_dat_o[8] = ch_dat_i_8;
    assign wb_dat_o[7] = ch_dat_i_7;
    assign wb_dat_o[6] = ch_dat_i_6;
    assign wb_dat_o[5] = ch_dat_i_5;
    assign wb_dat_o[4] = ch_dat_i_4;
    assign wb_dat_o[3] = ch_dat_i_3;
    assign wb_dat_o[2] = ch_dat_i_2;
    assign wb_dat_o[1] = ch_dat_i_1;
    assign wb_dat_o[0] = ch_dat_i_0;
    assign wb_adr_o[11] = ch_adr_i_11;
    assign wb_adr_o[10] = ch_adr_i_10;
    assign wb_adr_o[9] = ch_adr_i_9;
    assign wb_adr_o[8] = ch_adr_i_8;
    assign wb_adr_o[7] = ch_adr_i_7;
    assign wb_adr_o[6] = ch_adr_i_6;
    assign wb_adr_o[5] = ch_adr_i_5;
    assign wb_adr_o[4] = ch_adr_i_4;
    assign wb_adr_o[3] = ch_adr_i_3;
    assign wb_adr_o[2] = ch_adr_i_2;
    assign wb_adr_o[1] = ch_adr_i_1;
    assign wb_adr_o[0] = ch_adr_i_0;
    dffph_2 \ch_dat_o_reg[4]  ( .q(ch_dat_o[4]), .d(wb_dat_i[4]), .ck(n7), .g(
        n4) );
    dffph_2 \ch_dat_o_reg[3]  ( .q(ch_dat_o[3]), .d(wb_dat_i[3]), .ck(n7), .g(
        n4) );
    dffph_2 \ch_dat_o_reg[2]  ( .q(ch_dat_o[2]), .d(wb_dat_i[2]), .ck(n7), .g(
        n4) );
    dffph_2 \ch_dat_o_reg[1]  ( .q(ch_dat_o[1]), .d(wb_dat_i[1]), .ck(n7), .g(
        n4) );
    dffph_2 \ch_dat_o_reg[0]  ( .q(ch_dat_o[0]), .d(wb_dat_i[0]), .ck(n7), .g(
        n3) );
    oa21_2 \reqoGate/U1  ( .x(\reqoGate/n2 ), .a(\reqoGate/n2 ), .b(
        \reqoGate/nr ), .c(\reqoGate/nd ) );
    ao33_1 \cycGate/U1/U1  ( .x(wb_stb_cyc_o), .a(sync_ack_inv), .b(
        wb_stb_cyc_o), .c(reset_b), .d(sync_ack_inv), .e(rsync), .f(ch_idle)
         );
    dffph_2 \ch_dat_o_reg[19]  ( .q(ch_dat_o[19]), .d(wb_dat_i[19]), .ck(n5), 
        .g(n2) );
    dffph_2 \ch_dat_o_reg[18]  ( .q(ch_dat_o[18]), .d(wb_dat_i[18]), .ck(n5), 
        .g(n2) );
    dffph_2 \ch_dat_o_reg[17]  ( .q(ch_dat_o[17]), .d(wb_dat_i[17]), .ck(n6), 
        .g(n2) );
    dffph_2 \ch_dat_o_reg[16]  ( .q(ch_dat_o[16]), .d(wb_dat_i[16]), .ck(n5), 
        .g(n3) );
    dffph_2 \ch_dat_o_reg[15]  ( .q(ch_dat_o[15]), .d(wb_dat_i[15]), .ck(n6), 
        .g(n3) );
    dffph_2 \ch_dat_o_reg[14]  ( .q(ch_dat_o[14]), .d(wb_dat_i[14]), .ck(n6), 
        .g(n3) );
    dffph_2 \ch_dat_o_reg[13]  ( .q(ch_dat_o[13]), .d(wb_dat_i[13]), .ck(n6), 
        .g(n3) );
    dffph_2 \ch_dat_o_reg[12]  ( .q(ch_dat_o[12]), .d(wb_dat_i[12]), .ck(n6), 
        .g(n3) );
    dffph_2 \ch_dat_o_reg[11]  ( .q(ch_dat_o[11]), .d(wb_dat_i[11]), .ck(n7), 
        .g(n4) );
    dffph_2 \ch_dat_o_reg[10]  ( .q(ch_dat_o[10]), .d(wb_dat_i[10]), .ck(n7), 
        .g(n4) );
    dffph_2 \ch_dat_o_reg[9]  ( .q(ch_dat_o[9]), .d(wb_dat_i[9]), .ck(n7), .g(
        n4) );
    dffph_2 \ch_dat_o_reg[8]  ( .q(ch_dat_o[8]), .d(wb_dat_i[8]), .ck(n7), .g(
        n4) );
    dffph_2 \ch_dat_o_reg[7]  ( .q(ch_dat_o[7]), .d(wb_dat_i[7]), .ck(n7), .g(
        n4) );
    dffph_2 \ch_dat_o_reg[6]  ( .q(ch_dat_o[6]), .d(wb_dat_i[6]), .ck(n7), .g(
        n4) );
    dffph_2 \ch_dat_o_reg[5]  ( .q(ch_dat_o[5]), .d(wb_dat_i[5]), .ck(n7), .g(
        n4) );
    dffpr_2 rsync_reg ( .q(rsync), .rb(reset_b), .d(rin1), .ck(n6) );
    dffpr_2 rin1_reg ( .q(rin1), .rb(reset_b), .d(ch_req_i), .ck(n6) );
    dffpr_2 sync_ack_l_reg ( .q(sync_ack_l), .qb(sync_ack_inv), .rb(reset_b), 
        .d(n2), .ck(n6) );
    dffph_2 \ch_dat_o_reg[31]  ( .q(ch_dat_o[31]), .d(wb_dat_i[31]), .ck(n5), 
        .g(n3) );
    dffph_2 \ch_dat_o_reg[30]  ( .q(ch_dat_o[30]), .d(wb_dat_i[30]), .ck(n6), 
        .g(n2) );
    dffph_2 \ch_dat_o_reg[29]  ( .q(ch_dat_o[29]), .d(wb_dat_i[29]), .ck(n5), 
        .g(n3) );
    dffph_2 \ch_dat_o_reg[28]  ( .q(ch_dat_o[28]), .d(wb_dat_i[28]), .ck(n6), 
        .g(n2) );
    dffph_2 \ch_dat_o_reg[27]  ( .q(ch_dat_o[27]), .d(wb_dat_i[27]), .ck(n5), 
        .g(n3) );
    dffph_2 \ch_dat_o_reg[26]  ( .q(ch_dat_o[26]), .d(wb_dat_i[26]), .ck(n6), 
        .g(n2) );
    dffph_2 \ch_dat_o_reg[25]  ( .q(ch_dat_o[25]), .d(wb_dat_i[25]), .ck(n5), 
        .g(n3) );
    dffph_2 \ch_dat_o_reg[24]  ( .q(ch_dat_o[24]), .d(wb_dat_i[24]), .ck(n5), 
        .g(n2) );
    dffph_2 \ch_dat_o_reg[23]  ( .q(ch_dat_o[23]), .d(wb_dat_i[23]), .ck(n5), 
        .g(n3) );
    dffph_2 \ch_dat_o_reg[22]  ( .q(ch_dat_o[22]), .d(wb_dat_i[22]), .ck(n5), 
        .g(n2) );
    dffph_2 \ch_dat_o_reg[21]  ( .q(ch_dat_o[21]), .d(wb_dat_i[21]), .ck(n5), 
        .g(n2) );
    dffph_2 \ch_dat_o_reg[20]  ( .q(ch_dat_o[20]), .d(wb_dat_i[20]), .ck(n5), 
        .g(n2) );
    nor3_0 U3 ( .x(\reqoGate/nr ), .a(n1), .b(sync_ack_l), .c(rsync) );
    nand3_0 U4 ( .x(\reqoGate/nd ), .a(rsync), .b(n1), .c(sync_ack_l) );
    inv_0 U5 ( .x(ch_req_o_wire), .a(\reqoGate/n2 ) );
    nor2_0 U6 ( .x(ch_idle), .a(ch_ack_i), .b(ch_ack_o) );
    nor2i_0 U7 ( .x(n1), .a(reset_b), .b(ch_ack_o) );
    buf_3 U8 ( .x(n2), .a(wb_ack_i) );
    buf_3 U9 ( .x(n4), .a(wb_ack_i) );
    buf_3 U10 ( .x(n3), .a(wb_ack_i) );
    buf_3 U11 ( .x(n5), .a(clk) );
    buf_3 U12 ( .x(n7), .a(clk) );
    buf_3 U13 ( .x(n6), .a(clk) );
    buf_3 U14 ( .x(ch_ack_i), .a(ch_req_o_wire) );
endmodule


module wb_block ( nReset, clk, chaincommand, nchaincommandack, chainresponse, 
    nchainresponseack, e_dp, e_ip, e_tic, r_dp, r_ip, r_tic, wb_we_o, 
    wb_stb_cyc_o, wb_ack_i, wb_adr_o, wb_dat_i, wb_dat_o );
input  [4:0] chaincommand;
output [4:0] chainresponse;
input  [2:0] e_dp;
input  [2:0] e_ip;
input  [2:0] e_tic;
input  [2:0] r_dp;
input  [2:0] r_ip;
input  [2:0] r_tic;
output [11:0] wb_adr_o;
input  [31:0] wb_dat_i;
output [31:0] wb_dat_o;
input  nReset, clk, nchainresponseack, wb_ack_i;
output nchaincommandack, wb_we_o, wb_stb_cyc_o;
    wire sc_req, sc_we, sc_ack, sr_req, sr_ack, \sr_dat[31] , \sr_dat[30] , 
        \sr_dat[29] , \sr_dat[28] , \sr_dat[27] , \sr_dat[26] , \sr_dat[25] , 
        \sr_dat[24] , \sr_dat[23] , \sr_dat[22] , \sr_dat[21] , \sr_dat[20] , 
        \sr_dat[19] , \sr_dat[18] , \sr_dat[17] , \sr_dat[16] , \sr_dat[15] , 
        \sr_dat[14] , \sr_dat[13] , \sr_dat[12] , \sr_dat[11] , \sr_dat[10] , 
        \sr_dat[9] , \sr_dat[8] , \sr_dat[7] , \sr_dat[6] , \sr_dat[5] , 
        \sr_dat[4] , \sr_dat[3] , \sr_dat[2] , \sr_dat[1] , \sr_dat[0] , 
        \sc_st[4] , \sc_st[3] , \sc_st[2] , \sc_st[1] , \sc_st[0] , 
        \sc_dat[31] , \sc_dat[30] , \sc_dat[29] , \sc_dat[28] , \sc_dat[27] , 
        \sc_dat[26] , \sc_dat[25] , \sc_dat[24] , \sc_dat[23] , \sc_dat[22] , 
        \sc_dat[21] , \sc_dat[20] , \sc_dat[19] , \sc_dat[18] , \sc_dat[17] , 
        \sc_dat[16] , \sc_dat[15] , \sc_dat[14] , \sc_dat[13] , \sc_dat[12] , 
        \sc_dat[11] , \sc_dat[10] , \sc_dat[9] , \sc_dat[8] , \sc_dat[7] , 
        \sc_dat[6] , \sc_dat[5] , \sc_dat[4] , \sc_dat[3] , \sc_dat[2] , 
        \sc_dat[1] , \sc_dat[0] , SYNOPSYS_UNCONNECTED_1, 
        SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, 
        SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, 
        SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, \sc_adr[13] , \sc_adr[12] , \sc_adr[11] , 
        \sc_adr[10] , \sc_adr[9] , \sc_adr[8] , \sc_adr[7] , \sc_adr[6] , 
        \sc_adr[5] , \sc_adr[4] , \sc_adr[3] , \sc_adr[2] , 
        SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20;
    slave_if_wb wbIf ( .nReset(nReset), .sc_req(sc_req), .sc_we(sc_we), 
        .sc_st({\sc_st[4] , \sc_st[3] , \sc_st[2] , \sc_st[1] , \sc_st[0] }), 
        .sc_adr({SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, 
        SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, 
        SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, 
        SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10, 
        SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12, 
        SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14, 
        SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16, 
        SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18, \sc_adr[13] , 
        \sc_adr[12] , \sc_adr[11] , \sc_adr[10] , \sc_adr[9] , \sc_adr[8] , 
        \sc_adr[7] , \sc_adr[6] , \sc_adr[5] , \sc_adr[4] , \sc_adr[3] , 
        \sc_adr[2] , SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20}), 
        .sc_dat({\sc_dat[31] , \sc_dat[30] , \sc_dat[29] , \sc_dat[28] , 
        \sc_dat[27] , \sc_dat[26] , \sc_dat[25] , \sc_dat[24] , \sc_dat[23] , 
        \sc_dat[22] , \sc_dat[21] , \sc_dat[20] , \sc_dat[19] , \sc_dat[18] , 
        \sc_dat[17] , \sc_dat[16] , \sc_dat[15] , \sc_dat[14] , \sc_dat[13] , 
        \sc_dat[12] , \sc_dat[11] , \sc_dat[10] , \sc_dat[9] , \sc_dat[8] , 
        \sc_dat[7] , \sc_dat[6] , \sc_dat[5] , \sc_dat[4] , \sc_dat[3] , 
        \sc_dat[2] , \sc_dat[1] , \sc_dat[0] }), .sc_ack(sc_ack), .sr_req(
        sr_req), .sr_err(1'b0), .sr_rty(1'b0), .sr_acc(1'b0), .sr_mult(1'b0), 
        .sr_ts({1'b0, 1'b0, 1'b0}), .sr_rt({\sc_st[4] , \sc_st[3] , \sc_st[2] , 
        \sc_st[1] , \sc_st[0] }), .sr_sel({1'b1, 1'b1, 1'b1, 1'b1}), .sr_dat({
        \sr_dat[31] , \sr_dat[30] , \sr_dat[29] , \sr_dat[28] , \sr_dat[27] , 
        \sr_dat[26] , \sr_dat[25] , \sr_dat[24] , \sr_dat[23] , \sr_dat[22] , 
        \sr_dat[21] , \sr_dat[20] , \sr_dat[19] , \sr_dat[18] , \sr_dat[17] , 
        \sr_dat[16] , \sr_dat[15] , \sr_dat[14] , \sr_dat[13] , \sr_dat[12] , 
        \sr_dat[11] , \sr_dat[10] , \sr_dat[9] , \sr_dat[8] , \sr_dat[7] , 
        \sr_dat[6] , \sr_dat[5] , \sr_dat[4] , \sr_dat[3] , \sr_dat[2] , 
        \sr_dat[1] , \sr_dat[0] }), .sr_ack(sr_ack), .chaincommand(
        chaincommand), .nchaincommandack(nchaincommandack), .chainresponse(
        chainresponse), .nchainresponseack(nchainresponseack), .e_dp(e_dp), 
        .e_ip(e_ip), .e_tic(e_tic), .r_dp(r_dp), .r_ip(r_ip), .r_tic(r_tic) );
    wishbone wbconv ( .reset_b(nReset), .clk(clk), .ch_we_i(sc_we), .ch_dat_i(
        {\sc_dat[31] , \sc_dat[30] , \sc_dat[29] , \sc_dat[28] , \sc_dat[27] , 
        \sc_dat[26] , \sc_dat[25] , \sc_dat[24] , \sc_dat[23] , \sc_dat[22] , 
        \sc_dat[21] , \sc_dat[20] , \sc_dat[19] , \sc_dat[18] , \sc_dat[17] , 
        \sc_dat[16] , \sc_dat[15] , \sc_dat[14] , \sc_dat[13] , \sc_dat[12] , 
        \sc_dat[11] , \sc_dat[10] , \sc_dat[9] , \sc_dat[8] , \sc_dat[7] , 
        \sc_dat[6] , \sc_dat[5] , \sc_dat[4] , \sc_dat[3] , \sc_dat[2] , 
        \sc_dat[1] , \sc_dat[0] }), .ch_adr_i({\sc_adr[13] , \sc_adr[12] , 
        \sc_adr[11] , \sc_adr[10] , \sc_adr[9] , \sc_adr[8] , \sc_adr[7] , 
        \sc_adr[6] , \sc_adr[5] , \sc_adr[4] , \sc_adr[3] , \sc_adr[2] }), 
        .ch_req_i(sc_req), .ch_ack_i(sc_ack), .ch_req_o(sr_req), .ch_dat_o({
        \sr_dat[31] , \sr_dat[30] , \sr_dat[29] , \sr_dat[28] , \sr_dat[27] , 
        \sr_dat[26] , \sr_dat[25] , \sr_dat[24] , \sr_dat[23] , \sr_dat[22] , 
        \sr_dat[21] , \sr_dat[20] , \sr_dat[19] , \sr_dat[18] , \sr_dat[17] , 
        \sr_dat[16] , \sr_dat[15] , \sr_dat[14] , \sr_dat[13] , \sr_dat[12] , 
        \sr_dat[11] , \sr_dat[10] , \sr_dat[9] , \sr_dat[8] , \sr_dat[7] , 
        \sr_dat[6] , \sr_dat[5] , \sr_dat[4] , \sr_dat[3] , \sr_dat[2] , 
        \sr_dat[1] , \sr_dat[0] }), .ch_ack_o(sr_ack), .wb_we_o(wb_we_o), 
        .wb_stb_cyc_o(wb_stb_cyc_o), .wb_dat_o(wb_dat_o), .wb_adr_o(wb_adr_o), 
        .wb_dat_i(wb_dat_i), .wb_ack_i(wb_ack_i) );
endmodule


module chain_sendmux8_14 ( ctrlack, oh, ol, i_h, i_l, ctrlreq, oa );
output [7:0] oh;
output [7:0] ol;
input  [7:0] i_h;
input  [7:0] i_l;
input  ctrlreq, oa;
output ctrlack;
    wire \drive[1] , \drive[0] , \U1693/drivemonitor , \U1693/naa , 
        \U1693/net2 , \U1693/net3 , \U1693/bdone , \U1693/U1702/Z ;
    and2_1 \U33_0_/U8  ( .x(oh[0]), .a(i_h[0]), .b(\drive[1] ) );
    and2_1 \U33_1_/U8  ( .x(oh[1]), .a(i_h[1]), .b(\drive[1] ) );
    and2_1 \U33_2_/U8  ( .x(oh[2]), .a(i_h[2]), .b(\drive[1] ) );
    and2_1 \U33_3_/U8  ( .x(oh[3]), .a(i_h[3]), .b(\drive[1] ) );
    and2_1 \U33_4_/U8  ( .x(oh[4]), .a(i_h[4]), .b(\drive[1] ) );
    and2_1 \U33_5_/U8  ( .x(oh[5]), .a(i_h[5]), .b(\drive[1] ) );
    and2_1 \U33_6_/U8  ( .x(oh[6]), .a(i_h[6]), .b(\drive[1] ) );
    and2_1 \U33_7_/U8  ( .x(oh[7]), .a(i_h[7]), .b(\drive[1] ) );
    and2_1 \U1670_0_/U8  ( .x(ol[0]), .a(\drive[0] ), .b(i_l[0]) );
    and2_1 \U1670_1_/U8  ( .x(ol[1]), .a(\drive[0] ), .b(i_l[1]) );
    and2_1 \U1670_2_/U8  ( .x(ol[2]), .a(\drive[0] ), .b(i_l[2]) );
    and2_1 \U1670_3_/U8  ( .x(ol[3]), .a(\drive[0] ), .b(i_l[3]) );
    and2_1 \U1670_4_/U8  ( .x(ol[4]), .a(\drive[0] ), .b(i_l[4]) );
    and2_1 \U1670_5_/U8  ( .x(ol[5]), .a(\drive[0] ), .b(i_l[5]) );
    and2_1 \U1670_6_/U8  ( .x(ol[6]), .a(\drive[0] ), .b(i_l[6]) );
    and2_1 \U1670_7_/U8  ( .x(ol[7]), .a(\drive[0] ), .b(i_l[7]) );
    nor2_2 \U1693/U1703/U6  ( .x(ctrlack), .a(\U1693/drivemonitor ), .b(
        \U1693/naa ) );
    inv_2 \U1693/U1699/U3  ( .x(\U1693/net2 ), .a(\U1693/net3 ) );
    and2_4 \U1693/U2_0_/U8  ( .x(\drive[0] ), .a(ctrlreq), .b(\U1693/net2 ) );
    and2_4 \U1693/U2_1_/U8  ( .x(\drive[1] ), .a(ctrlreq), .b(\U1693/net2 ) );
    inv_1 \U1693/U1701/U3  ( .x(\U1693/naa ), .a(\U1693/bdone ) );
    ao222_1 \U1693/U13/U18/U1/U1  ( .x(\U1693/drivemonitor ), .a(\drive[1] ), 
        .b(\drive[0] ), .c(\drive[1] ), .d(\U1693/drivemonitor ), .e(
        \drive[0] ), .f(\U1693/drivemonitor ) );
    aoi21_1 \U1693/U1702/U30/U1/U1  ( .x(\U1693/bdone ), .a(\U1693/U1702/Z ), 
        .b(oa), .c(\U1693/net2 ) );
    inv_1 \U1693/U1702/U30/U1/U2  ( .x(\U1693/U1702/Z ), .a(\U1693/bdone ) );
    ao23_1 \U1693/U1693/U21/U1/U1  ( .x(\U1693/net3 ), .a(ctrlreq), .b(
        \U1693/net3 ), .c(ctrlreq), .d(\U1693/drivemonitor ), .e(oa) );
endmodule


module chain_sendmux8_13 ( ctrlack, oh, ol, i_h, i_l, ctrlreq, oa );
output [7:0] oh;
output [7:0] ol;
input  [7:0] i_h;
input  [7:0] i_l;
input  ctrlreq, oa;
output ctrlack;
    wire \drive[1] , \drive[0] , \U1693/drivemonitor , \U1693/naa , 
        \U1693/net2 , \U1693/net3 , \U1693/bdone , \U1693/U1702/Z ;
    and2_1 \U33_0_/U8  ( .x(oh[0]), .a(i_h[0]), .b(\drive[1] ) );
    and2_1 \U33_1_/U8  ( .x(oh[1]), .a(i_h[1]), .b(\drive[1] ) );
    and2_1 \U33_2_/U8  ( .x(oh[2]), .a(i_h[2]), .b(\drive[1] ) );
    and2_1 \U33_3_/U8  ( .x(oh[3]), .a(i_h[3]), .b(\drive[1] ) );
    and2_1 \U33_4_/U8  ( .x(oh[4]), .a(i_h[4]), .b(\drive[1] ) );
    and2_1 \U33_5_/U8  ( .x(oh[5]), .a(i_h[5]), .b(\drive[1] ) );
    and2_1 \U33_6_/U8  ( .x(oh[6]), .a(i_h[6]), .b(\drive[1] ) );
    and2_1 \U33_7_/U8  ( .x(oh[7]), .a(i_h[7]), .b(\drive[1] ) );
    and2_1 \U1670_0_/U8  ( .x(ol[0]), .a(\drive[0] ), .b(i_l[0]) );
    and2_1 \U1670_1_/U8  ( .x(ol[1]), .a(\drive[0] ), .b(i_l[1]) );
    and2_1 \U1670_2_/U8  ( .x(ol[2]), .a(\drive[0] ), .b(i_l[2]) );
    and2_1 \U1670_3_/U8  ( .x(ol[3]), .a(\drive[0] ), .b(i_l[3]) );
    and2_1 \U1670_4_/U8  ( .x(ol[4]), .a(\drive[0] ), .b(i_l[4]) );
    and2_1 \U1670_5_/U8  ( .x(ol[5]), .a(\drive[0] ), .b(i_l[5]) );
    and2_1 \U1670_6_/U8  ( .x(ol[6]), .a(\drive[0] ), .b(i_l[6]) );
    and2_1 \U1670_7_/U8  ( .x(ol[7]), .a(\drive[0] ), .b(i_l[7]) );
    nor2_2 \U1693/U1703/U6  ( .x(ctrlack), .a(\U1693/drivemonitor ), .b(
        \U1693/naa ) );
    inv_2 \U1693/U1699/U3  ( .x(\U1693/net2 ), .a(\U1693/net3 ) );
    and2_4 \U1693/U2_0_/U8  ( .x(\drive[0] ), .a(ctrlreq), .b(\U1693/net2 ) );
    and2_4 \U1693/U2_1_/U8  ( .x(\drive[1] ), .a(ctrlreq), .b(\U1693/net2 ) );
    inv_1 \U1693/U1701/U3  ( .x(\U1693/naa ), .a(\U1693/bdone ) );
    ao222_1 \U1693/U13/U18/U1/U1  ( .x(\U1693/drivemonitor ), .a(\drive[1] ), 
        .b(\drive[0] ), .c(\drive[1] ), .d(\U1693/drivemonitor ), .e(
        \drive[0] ), .f(\U1693/drivemonitor ) );
    aoi21_1 \U1693/U1702/U30/U1/U1  ( .x(\U1693/bdone ), .a(\U1693/U1702/Z ), 
        .b(oa), .c(\U1693/net2 ) );
    inv_1 \U1693/U1702/U30/U1/U2  ( .x(\U1693/U1702/Z ), .a(\U1693/bdone ) );
    ao23_1 \U1693/U1693/U21/U1/U1  ( .x(\U1693/net3 ), .a(ctrlreq), .b(
        \U1693/net3 ), .c(ctrlreq), .d(\U1693/drivemonitor ), .e(oa) );
endmodule


module chain_sendmux8_12 ( ctrlack, oh, ol, i_h, i_l, ctrlreq, oa );
output [7:0] oh;
output [7:0] ol;
input  [7:0] i_h;
input  [7:0] i_l;
input  ctrlreq, oa;
output ctrlack;
    wire \drive[1] , \drive[0] , \U1693/drivemonitor , \U1693/naa , 
        \U1693/net2 , \U1693/net3 , \U1693/bdone , \U1693/U1702/Z ;
    and2_1 \U33_0_/U8  ( .x(oh[0]), .a(i_h[0]), .b(\drive[1] ) );
    and2_1 \U33_1_/U8  ( .x(oh[1]), .a(i_h[1]), .b(\drive[1] ) );
    and2_1 \U33_2_/U8  ( .x(oh[2]), .a(i_h[2]), .b(\drive[1] ) );
    and2_1 \U33_3_/U8  ( .x(oh[3]), .a(i_h[3]), .b(\drive[1] ) );
    and2_1 \U33_4_/U8  ( .x(oh[4]), .a(i_h[4]), .b(\drive[1] ) );
    and2_1 \U33_5_/U8  ( .x(oh[5]), .a(i_h[5]), .b(\drive[1] ) );
    and2_1 \U33_6_/U8  ( .x(oh[6]), .a(i_h[6]), .b(\drive[1] ) );
    and2_1 \U33_7_/U8  ( .x(oh[7]), .a(i_h[7]), .b(\drive[1] ) );
    and2_1 \U1670_0_/U8  ( .x(ol[0]), .a(\drive[0] ), .b(i_l[0]) );
    and2_1 \U1670_1_/U8  ( .x(ol[1]), .a(\drive[0] ), .b(i_l[1]) );
    and2_1 \U1670_2_/U8  ( .x(ol[2]), .a(\drive[0] ), .b(i_l[2]) );
    and2_1 \U1670_3_/U8  ( .x(ol[3]), .a(\drive[0] ), .b(i_l[3]) );
    and2_1 \U1670_4_/U8  ( .x(ol[4]), .a(\drive[0] ), .b(i_l[4]) );
    and2_1 \U1670_5_/U8  ( .x(ol[5]), .a(\drive[0] ), .b(i_l[5]) );
    and2_1 \U1670_6_/U8  ( .x(ol[6]), .a(\drive[0] ), .b(i_l[6]) );
    and2_1 \U1670_7_/U8  ( .x(ol[7]), .a(\drive[0] ), .b(i_l[7]) );
    nor2_2 \U1693/U1703/U6  ( .x(ctrlack), .a(\U1693/drivemonitor ), .b(
        \U1693/naa ) );
    inv_2 \U1693/U1699/U3  ( .x(\U1693/net2 ), .a(\U1693/net3 ) );
    and2_4 \U1693/U2_0_/U8  ( .x(\drive[0] ), .a(ctrlreq), .b(\U1693/net2 ) );
    and2_4 \U1693/U2_1_/U8  ( .x(\drive[1] ), .a(ctrlreq), .b(\U1693/net2 ) );
    inv_1 \U1693/U1701/U3  ( .x(\U1693/naa ), .a(\U1693/bdone ) );
    ao222_1 \U1693/U13/U18/U1/U1  ( .x(\U1693/drivemonitor ), .a(\drive[1] ), 
        .b(\drive[0] ), .c(\drive[1] ), .d(\U1693/drivemonitor ), .e(
        \drive[0] ), .f(\U1693/drivemonitor ) );
    aoi21_1 \U1693/U1702/U30/U1/U1  ( .x(\U1693/bdone ), .a(\U1693/U1702/Z ), 
        .b(oa), .c(\U1693/net2 ) );
    inv_1 \U1693/U1702/U30/U1/U2  ( .x(\U1693/U1702/Z ), .a(\U1693/bdone ) );
    ao23_1 \U1693/U1693/U21/U1/U1  ( .x(\U1693/net3 ), .a(ctrlreq), .b(
        \U1693/net3 ), .c(ctrlreq), .d(\U1693/drivemonitor ), .e(oa) );
endmodule


module chain_sendmux8_15 ( ctrlack, oh, ol, i_h, i_l, ctrlreq, oa );
output [7:0] oh;
output [7:0] ol;
input  [7:0] i_h;
input  [7:0] i_l;
input  ctrlreq, oa;
output ctrlack;
    wire \drive[1] , \drive[0] , \U1693/drivemonitor , \U1693/naa , 
        \U1693/net2 , \U1693/net3 , \U1693/bdone , \U1693/U1702/Z ;
    and2_1 \U33_0_/U8  ( .x(oh[0]), .a(i_h[0]), .b(\drive[1] ) );
    and2_1 \U33_1_/U8  ( .x(oh[1]), .a(i_h[1]), .b(\drive[1] ) );
    and2_1 \U33_2_/U8  ( .x(oh[2]), .a(i_h[2]), .b(\drive[1] ) );
    and2_1 \U33_3_/U8  ( .x(oh[3]), .a(i_h[3]), .b(\drive[1] ) );
    and2_1 \U33_4_/U8  ( .x(oh[4]), .a(i_h[4]), .b(\drive[1] ) );
    and2_1 \U33_5_/U8  ( .x(oh[5]), .a(i_h[5]), .b(\drive[1] ) );
    and2_1 \U33_6_/U8  ( .x(oh[6]), .a(i_h[6]), .b(\drive[1] ) );
    and2_1 \U33_7_/U8  ( .x(oh[7]), .a(i_h[7]), .b(\drive[1] ) );
    and2_1 \U1670_0_/U8  ( .x(ol[0]), .a(\drive[0] ), .b(i_l[0]) );
    and2_1 \U1670_1_/U8  ( .x(ol[1]), .a(\drive[0] ), .b(i_l[1]) );
    and2_1 \U1670_2_/U8  ( .x(ol[2]), .a(\drive[0] ), .b(i_l[2]) );
    and2_1 \U1670_3_/U8  ( .x(ol[3]), .a(\drive[0] ), .b(i_l[3]) );
    and2_1 \U1670_4_/U8  ( .x(ol[4]), .a(\drive[0] ), .b(i_l[4]) );
    and2_1 \U1670_5_/U8  ( .x(ol[5]), .a(\drive[0] ), .b(i_l[5]) );
    and2_1 \U1670_6_/U8  ( .x(ol[6]), .a(\drive[0] ), .b(i_l[6]) );
    and2_1 \U1670_7_/U8  ( .x(ol[7]), .a(\drive[0] ), .b(i_l[7]) );
    nor2_2 \U1693/U1703/U6  ( .x(ctrlack), .a(\U1693/drivemonitor ), .b(
        \U1693/naa ) );
    inv_2 \U1693/U1699/U3  ( .x(\U1693/net2 ), .a(\U1693/net3 ) );
    and2_4 \U1693/U2_0_/U8  ( .x(\drive[0] ), .a(ctrlreq), .b(\U1693/net2 ) );
    and2_4 \U1693/U2_1_/U8  ( .x(\drive[1] ), .a(ctrlreq), .b(\U1693/net2 ) );
    inv_1 \U1693/U1701/U3  ( .x(\U1693/naa ), .a(\U1693/bdone ) );
    ao222_1 \U1693/U13/U18/U1/U1  ( .x(\U1693/drivemonitor ), .a(\drive[1] ), 
        .b(\drive[0] ), .c(\drive[1] ), .d(\U1693/drivemonitor ), .e(
        \drive[0] ), .f(\U1693/drivemonitor ) );
    aoi21_1 \U1693/U1702/U30/U1/U1  ( .x(\U1693/bdone ), .a(\U1693/U1702/Z ), 
        .b(oa), .c(\U1693/net2 ) );
    inv_1 \U1693/U1702/U30/U1/U2  ( .x(\U1693/U1702/Z ), .a(\U1693/bdone ) );
    ao23_1 \U1693/U1693/U21/U1/U1  ( .x(\U1693/net3 ), .a(ctrlreq), .b(
        \U1693/net3 ), .c(ctrlreq), .d(\U1693/drivemonitor ), .e(oa) );
endmodule


module chain_sendword_2 ( ctrlack, oh, ol, chainackff, ctrlreq, ih, il );
output [7:0] oh;
output [7:0] ol;
input  [31:0] ih;
input  [31:0] il;
input  chainackff, ctrlreq;
output ctrlack;
    wire net44, \fourth_ol[7] , \fourth_ol[6] , \fourth_ol[5] , \fourth_ol[4] , 
        \fourth_ol[3] , \fourth_ol[2] , \fourth_ol[1] , \fourth_ol[0] , 
        \fourth_oh[7] , \fourth_oh[6] , \fourth_oh[5] , \fourth_oh[4] , 
        \fourth_oh[3] , \fourth_oh[2] , \fourth_oh[1] , \fourth_oh[0] , net51, 
        \third_ol[7] , \third_ol[6] , \third_ol[5] , \third_ol[4] , 
        \third_ol[3] , \third_ol[2] , \third_ol[1] , \third_ol[0] , 
        \third_oh[7] , \third_oh[6] , \third_oh[5] , \third_oh[4] , 
        \third_oh[3] , \third_oh[2] , \third_oh[1] , \third_oh[0] , net58, 
        \second_ol[7] , \second_ol[6] , \second_ol[5] , \second_ol[4] , 
        \second_ol[3] , \second_ol[2] , \second_ol[1] , \second_ol[0] , 
        \second_oh[7] , \second_oh[6] , \second_oh[5] , \second_oh[4] , 
        \second_oh[3] , \second_oh[2] , \second_oh[1] , \second_oh[0] , 
        bctrlreq, \first_ol[7] , \first_ol[6] , \first_ol[5] , \first_ol[4] , 
        \first_ol[3] , \first_ol[2] , \first_ol[1] , \first_ol[0] , 
        \first_oh[7] , \first_oh[6] , \first_oh[5] , \first_oh[4] , 
        \first_oh[3] , \first_oh[2] , \first_oh[1] , \first_oh[0] , 
        \U309_0_/n5 , \U309_0_/n1 , \U309_0_/n2 , \U309_0_/n3 , \U309_0_/n4 , 
        \U309_1_/n5 , \U309_1_/n1 , \U309_1_/n2 , \U309_1_/n3 , \U309_1_/n4 , 
        \U309_2_/n5 , \U309_2_/n1 , \U309_2_/n2 , \U309_2_/n3 , \U309_2_/n4 , 
        \U309_3_/n5 , \U309_3_/n1 , \U309_3_/n2 , \U309_3_/n3 , \U309_3_/n4 , 
        \U309_4_/n5 , \U309_4_/n1 , \U309_4_/n2 , \U309_4_/n3 , \U309_4_/n4 , 
        \U309_5_/n5 , \U309_5_/n1 , \U309_5_/n2 , \U309_5_/n3 , \U309_5_/n4 , 
        \U309_6_/n5 , \U309_6_/n1 , \U309_6_/n2 , \U309_6_/n3 , \U309_6_/n4 , 
        \U309_7_/n5 , \U309_7_/n1 , \U309_7_/n2 , \U309_7_/n3 , \U309_7_/n4 , 
        \U310_0_/n5 , \U310_0_/n1 , \U310_0_/n2 , \U310_0_/n3 , \U310_0_/n4 , 
        \U310_1_/n5 , \U310_1_/n1 , \U310_1_/n2 , \U310_1_/n3 , \U310_1_/n4 , 
        \U310_2_/n5 , \U310_2_/n1 , \U310_2_/n2 , \U310_2_/n3 , \U310_2_/n4 , 
        \U310_3_/n5 , \U310_3_/n1 , \U310_3_/n2 , \U310_3_/n3 , \U310_3_/n4 , 
        \U310_4_/n5 , \U310_4_/n1 , \U310_4_/n2 , \U310_4_/n3 , \U310_4_/n4 , 
        \U310_5_/n5 , \U310_5_/n1 , \U310_5_/n2 , \U310_5_/n3 , \U310_5_/n4 , 
        \U310_6_/n5 , \U310_6_/n1 , \U310_6_/n2 , \U310_6_/n3 , \U310_6_/n4 , 
        \U310_7_/n5 , \U310_7_/n1 , \U310_7_/n2 , \U310_7_/n3 , \U310_7_/n4 ;
    chain_sendmux8_14 I4 ( .ctrlack(ctrlack), .oh({\fourth_oh[7] , 
        \fourth_oh[6] , \fourth_oh[5] , \fourth_oh[4] , \fourth_oh[3] , 
        \fourth_oh[2] , \fourth_oh[1] , \fourth_oh[0] }), .ol({\fourth_ol[7] , 
        \fourth_ol[6] , \fourth_ol[5] , \fourth_ol[4] , \fourth_ol[3] , 
        \fourth_ol[2] , \fourth_ol[1] , \fourth_ol[0] }), .i_h(ih[7:0]), .i_l(
        il[7:0]), .ctrlreq(net44), .oa(chainackff) );
    chain_sendmux8_13 I3 ( .ctrlack(net44), .oh({\third_oh[7] , \third_oh[6] , 
        \third_oh[5] , \third_oh[4] , \third_oh[3] , \third_oh[2] , 
        \third_oh[1] , \third_oh[0] }), .ol({\third_ol[7] , \third_ol[6] , 
        \third_ol[5] , \third_ol[4] , \third_ol[3] , \third_ol[2] , 
        \third_ol[1] , \third_ol[0] }), .i_h(ih[15:8]), .i_l(il[15:8]), 
        .ctrlreq(net51), .oa(chainackff) );
    chain_sendmux8_12 I2 ( .ctrlack(net51), .oh({\second_oh[7] , 
        \second_oh[6] , \second_oh[5] , \second_oh[4] , \second_oh[3] , 
        \second_oh[2] , \second_oh[1] , \second_oh[0] }), .ol({\second_ol[7] , 
        \second_ol[6] , \second_ol[5] , \second_ol[4] , \second_ol[3] , 
        \second_ol[2] , \second_ol[1] , \second_ol[0] }), .i_h(ih[23:16]), 
        .i_l(il[23:16]), .ctrlreq(net58), .oa(chainackff) );
    chain_sendmux8_15 U320 ( .ctrlack(net58), .oh({\first_oh[7] , 
        \first_oh[6] , \first_oh[5] , \first_oh[4] , \first_oh[3] , 
        \first_oh[2] , \first_oh[1] , \first_oh[0] }), .ol({\first_ol[7] , 
        \first_ol[6] , \first_ol[5] , \first_ol[4] , \first_ol[3] , 
        \first_ol[2] , \first_ol[1] , \first_ol[0] }), .i_h(ih[31:24]), .i_l(
        il[31:24]), .ctrlreq(bctrlreq), .oa(chainackff) );
    buf_2 \U328/U7  ( .x(bctrlreq), .a(ctrlreq) );
    and4_2 \U309_0_/U24  ( .x(\U309_0_/n5 ), .a(\U309_0_/n1 ), .b(\U309_0_/n2 
        ), .c(\U309_0_/n3 ), .d(\U309_0_/n4 ) );
    inv_1 \U309_0_/U1  ( .x(\U309_0_/n1 ), .a(\fourth_oh[0] ) );
    inv_1 \U309_0_/U2  ( .x(\U309_0_/n2 ), .a(\third_oh[0] ) );
    inv_1 \U309_0_/U3  ( .x(\U309_0_/n3 ), .a(\second_oh[0] ) );
    inv_1 \U309_0_/U4  ( .x(\U309_0_/n4 ), .a(\first_oh[0] ) );
    inv_4 \U309_0_/U5  ( .x(oh[0]), .a(\U309_0_/n5 ) );
    and4_2 \U309_1_/U24  ( .x(\U309_1_/n5 ), .a(\U309_1_/n1 ), .b(\U309_1_/n2 
        ), .c(\U309_1_/n3 ), .d(\U309_1_/n4 ) );
    inv_1 \U309_1_/U1  ( .x(\U309_1_/n1 ), .a(\fourth_oh[1] ) );
    inv_1 \U309_1_/U2  ( .x(\U309_1_/n2 ), .a(\third_oh[1] ) );
    inv_1 \U309_1_/U3  ( .x(\U309_1_/n3 ), .a(\second_oh[1] ) );
    inv_1 \U309_1_/U4  ( .x(\U309_1_/n4 ), .a(\first_oh[1] ) );
    inv_4 \U309_1_/U5  ( .x(oh[1]), .a(\U309_1_/n5 ) );
    and4_2 \U309_2_/U24  ( .x(\U309_2_/n5 ), .a(\U309_2_/n1 ), .b(\U309_2_/n2 
        ), .c(\U309_2_/n3 ), .d(\U309_2_/n4 ) );
    inv_1 \U309_2_/U1  ( .x(\U309_2_/n1 ), .a(\fourth_oh[2] ) );
    inv_1 \U309_2_/U2  ( .x(\U309_2_/n2 ), .a(\third_oh[2] ) );
    inv_1 \U309_2_/U3  ( .x(\U309_2_/n3 ), .a(\second_oh[2] ) );
    inv_1 \U309_2_/U4  ( .x(\U309_2_/n4 ), .a(\first_oh[2] ) );
    inv_4 \U309_2_/U5  ( .x(oh[2]), .a(\U309_2_/n5 ) );
    and4_2 \U309_3_/U24  ( .x(\U309_3_/n5 ), .a(\U309_3_/n1 ), .b(\U309_3_/n2 
        ), .c(\U309_3_/n3 ), .d(\U309_3_/n4 ) );
    inv_1 \U309_3_/U1  ( .x(\U309_3_/n1 ), .a(\fourth_oh[3] ) );
    inv_1 \U309_3_/U2  ( .x(\U309_3_/n2 ), .a(\third_oh[3] ) );
    inv_1 \U309_3_/U3  ( .x(\U309_3_/n3 ), .a(\second_oh[3] ) );
    inv_1 \U309_3_/U4  ( .x(\U309_3_/n4 ), .a(\first_oh[3] ) );
    inv_4 \U309_3_/U5  ( .x(oh[3]), .a(\U309_3_/n5 ) );
    and4_2 \U309_4_/U24  ( .x(\U309_4_/n5 ), .a(\U309_4_/n1 ), .b(\U309_4_/n2 
        ), .c(\U309_4_/n3 ), .d(\U309_4_/n4 ) );
    inv_1 \U309_4_/U1  ( .x(\U309_4_/n1 ), .a(\fourth_oh[4] ) );
    inv_1 \U309_4_/U2  ( .x(\U309_4_/n2 ), .a(\third_oh[4] ) );
    inv_1 \U309_4_/U3  ( .x(\U309_4_/n3 ), .a(\second_oh[4] ) );
    inv_1 \U309_4_/U4  ( .x(\U309_4_/n4 ), .a(\first_oh[4] ) );
    inv_4 \U309_4_/U5  ( .x(oh[4]), .a(\U309_4_/n5 ) );
    and4_2 \U309_5_/U24  ( .x(\U309_5_/n5 ), .a(\U309_5_/n1 ), .b(\U309_5_/n2 
        ), .c(\U309_5_/n3 ), .d(\U309_5_/n4 ) );
    inv_1 \U309_5_/U1  ( .x(\U309_5_/n1 ), .a(\fourth_oh[5] ) );
    inv_1 \U309_5_/U2  ( .x(\U309_5_/n2 ), .a(\third_oh[5] ) );
    inv_1 \U309_5_/U3  ( .x(\U309_5_/n3 ), .a(\second_oh[5] ) );
    inv_1 \U309_5_/U4  ( .x(\U309_5_/n4 ), .a(\first_oh[5] ) );
    inv_4 \U309_5_/U5  ( .x(oh[5]), .a(\U309_5_/n5 ) );
    and4_2 \U309_6_/U24  ( .x(\U309_6_/n5 ), .a(\U309_6_/n1 ), .b(\U309_6_/n2 
        ), .c(\U309_6_/n3 ), .d(\U309_6_/n4 ) );
    inv_1 \U309_6_/U1  ( .x(\U309_6_/n1 ), .a(\fourth_oh[6] ) );
    inv_1 \U309_6_/U2  ( .x(\U309_6_/n2 ), .a(\third_oh[6] ) );
    inv_1 \U309_6_/U3  ( .x(\U309_6_/n3 ), .a(\second_oh[6] ) );
    inv_1 \U309_6_/U4  ( .x(\U309_6_/n4 ), .a(\first_oh[6] ) );
    inv_4 \U309_6_/U5  ( .x(oh[6]), .a(\U309_6_/n5 ) );
    and4_2 \U309_7_/U24  ( .x(\U309_7_/n5 ), .a(\U309_7_/n1 ), .b(\U309_7_/n2 
        ), .c(\U309_7_/n3 ), .d(\U309_7_/n4 ) );
    inv_1 \U309_7_/U1  ( .x(\U309_7_/n1 ), .a(\fourth_oh[7] ) );
    inv_1 \U309_7_/U2  ( .x(\U309_7_/n2 ), .a(\third_oh[7] ) );
    inv_1 \U309_7_/U3  ( .x(\U309_7_/n3 ), .a(\second_oh[7] ) );
    inv_1 \U309_7_/U4  ( .x(\U309_7_/n4 ), .a(\first_oh[7] ) );
    inv_4 \U309_7_/U5  ( .x(oh[7]), .a(\U309_7_/n5 ) );
    and4_2 \U310_0_/U24  ( .x(\U310_0_/n5 ), .a(\U310_0_/n1 ), .b(\U310_0_/n2 
        ), .c(\U310_0_/n3 ), .d(\U310_0_/n4 ) );
    inv_1 \U310_0_/U1  ( .x(\U310_0_/n1 ), .a(\fourth_ol[0] ) );
    inv_1 \U310_0_/U2  ( .x(\U310_0_/n2 ), .a(\third_ol[0] ) );
    inv_1 \U310_0_/U3  ( .x(\U310_0_/n3 ), .a(\second_ol[0] ) );
    inv_1 \U310_0_/U4  ( .x(\U310_0_/n4 ), .a(\first_ol[0] ) );
    inv_4 \U310_0_/U5  ( .x(ol[0]), .a(\U310_0_/n5 ) );
    and4_2 \U310_1_/U24  ( .x(\U310_1_/n5 ), .a(\U310_1_/n1 ), .b(\U310_1_/n2 
        ), .c(\U310_1_/n3 ), .d(\U310_1_/n4 ) );
    inv_1 \U310_1_/U1  ( .x(\U310_1_/n1 ), .a(\fourth_ol[1] ) );
    inv_1 \U310_1_/U2  ( .x(\U310_1_/n2 ), .a(\third_ol[1] ) );
    inv_1 \U310_1_/U3  ( .x(\U310_1_/n3 ), .a(\second_ol[1] ) );
    inv_1 \U310_1_/U4  ( .x(\U310_1_/n4 ), .a(\first_ol[1] ) );
    inv_4 \U310_1_/U5  ( .x(ol[1]), .a(\U310_1_/n5 ) );
    and4_2 \U310_2_/U24  ( .x(\U310_2_/n5 ), .a(\U310_2_/n1 ), .b(\U310_2_/n2 
        ), .c(\U310_2_/n3 ), .d(\U310_2_/n4 ) );
    inv_1 \U310_2_/U1  ( .x(\U310_2_/n1 ), .a(\fourth_ol[2] ) );
    inv_1 \U310_2_/U2  ( .x(\U310_2_/n2 ), .a(\third_ol[2] ) );
    inv_1 \U310_2_/U3  ( .x(\U310_2_/n3 ), .a(\second_ol[2] ) );
    inv_1 \U310_2_/U4  ( .x(\U310_2_/n4 ), .a(\first_ol[2] ) );
    inv_4 \U310_2_/U5  ( .x(ol[2]), .a(\U310_2_/n5 ) );
    and4_2 \U310_3_/U24  ( .x(\U310_3_/n5 ), .a(\U310_3_/n1 ), .b(\U310_3_/n2 
        ), .c(\U310_3_/n3 ), .d(\U310_3_/n4 ) );
    inv_1 \U310_3_/U1  ( .x(\U310_3_/n1 ), .a(\fourth_ol[3] ) );
    inv_1 \U310_3_/U2  ( .x(\U310_3_/n2 ), .a(\third_ol[3] ) );
    inv_1 \U310_3_/U3  ( .x(\U310_3_/n3 ), .a(\second_ol[3] ) );
    inv_1 \U310_3_/U4  ( .x(\U310_3_/n4 ), .a(\first_ol[3] ) );
    inv_4 \U310_3_/U5  ( .x(ol[3]), .a(\U310_3_/n5 ) );
    and4_2 \U310_4_/U24  ( .x(\U310_4_/n5 ), .a(\U310_4_/n1 ), .b(\U310_4_/n2 
        ), .c(\U310_4_/n3 ), .d(\U310_4_/n4 ) );
    inv_1 \U310_4_/U1  ( .x(\U310_4_/n1 ), .a(\fourth_ol[4] ) );
    inv_1 \U310_4_/U2  ( .x(\U310_4_/n2 ), .a(\third_ol[4] ) );
    inv_1 \U310_4_/U3  ( .x(\U310_4_/n3 ), .a(\second_ol[4] ) );
    inv_1 \U310_4_/U4  ( .x(\U310_4_/n4 ), .a(\first_ol[4] ) );
    inv_4 \U310_4_/U5  ( .x(ol[4]), .a(\U310_4_/n5 ) );
    and4_2 \U310_5_/U24  ( .x(\U310_5_/n5 ), .a(\U310_5_/n1 ), .b(\U310_5_/n2 
        ), .c(\U310_5_/n3 ), .d(\U310_5_/n4 ) );
    inv_1 \U310_5_/U1  ( .x(\U310_5_/n1 ), .a(\fourth_ol[5] ) );
    inv_1 \U310_5_/U2  ( .x(\U310_5_/n2 ), .a(\third_ol[5] ) );
    inv_1 \U310_5_/U3  ( .x(\U310_5_/n3 ), .a(\second_ol[5] ) );
    inv_1 \U310_5_/U4  ( .x(\U310_5_/n4 ), .a(\first_ol[5] ) );
    inv_4 \U310_5_/U5  ( .x(ol[5]), .a(\U310_5_/n5 ) );
    and4_2 \U310_6_/U24  ( .x(\U310_6_/n5 ), .a(\U310_6_/n1 ), .b(\U310_6_/n2 
        ), .c(\U310_6_/n3 ), .d(\U310_6_/n4 ) );
    inv_1 \U310_6_/U1  ( .x(\U310_6_/n1 ), .a(\fourth_ol[6] ) );
    inv_1 \U310_6_/U2  ( .x(\U310_6_/n2 ), .a(\third_ol[6] ) );
    inv_1 \U310_6_/U3  ( .x(\U310_6_/n3 ), .a(\second_ol[6] ) );
    inv_1 \U310_6_/U4  ( .x(\U310_6_/n4 ), .a(\first_ol[6] ) );
    inv_4 \U310_6_/U5  ( .x(ol[6]), .a(\U310_6_/n5 ) );
    and4_2 \U310_7_/U24  ( .x(\U310_7_/n5 ), .a(\U310_7_/n1 ), .b(\U310_7_/n2 
        ), .c(\U310_7_/n3 ), .d(\U310_7_/n4 ) );
    inv_1 \U310_7_/U1  ( .x(\U310_7_/n1 ), .a(\fourth_ol[7] ) );
    inv_1 \U310_7_/U2  ( .x(\U310_7_/n2 ), .a(\third_ol[7] ) );
    inv_1 \U310_7_/U3  ( .x(\U310_7_/n3 ), .a(\second_ol[7] ) );
    inv_1 \U310_7_/U4  ( .x(\U310_7_/n4 ), .a(\first_ol[7] ) );
    inv_4 \U310_7_/U5  ( .x(ol[7]), .a(\U310_7_/n5 ) );
endmodule


module chain_dr8bit_completion_44 ( o, i );
input  [15:0] i;
output o;
    wire \nx[0] , \nx[1] , \nx[2] , \nx[3] , \ny[0] , \ny[1] , \ny[2] , 
        \ny[3] , y, x, \U6/Z , \U3/net3 , \U3/U20/Z , \U3/net2 , \U3/U21/Z , 
        \U3/U19/Z , \U5/net3 , \U5/U20/Z , \U5/net2 , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_47 ( o, i );
input  [15:0] i;
output o;
    wire \nx[0] , \nx[1] , \nx[2] , \nx[3] , \ny[0] , \ny[1] , \ny[2] , 
        \ny[3] , y, x, \U6/Z , \U3/net3 , \U3/U20/Z , \U3/net2 , \U3/U21/Z , 
        \U3/U19/Z , \U5/net3 , \U5/U20/Z , \U5/net2 , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_46 ( o, i );
input  [15:0] i;
output o;
    wire \nx[0] , \nx[1] , \nx[2] , \nx[3] , \ny[0] , \ny[1] , \ny[2] , 
        \ny[3] , y, x, \U6/Z , \U3/net3 , \U3/U20/Z , \U3/net2 , \U3/U21/Z , 
        \U3/U19/Z , \U5/net3 , \U5/U20/Z , \U5/net2 , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_45 ( o, i );
input  [15:0] i;
output o;
    wire \nx[0] , \nx[1] , \nx[2] , \nx[3] , \ny[0] , \ny[1] , \ny[2] , 
        \ny[3] , y, x, \U6/Z , \U3/net3 , \U3/U20/Z , \U3/net2 , \U3/U21/Z , 
        \U3/U19/Z , \U5/net3 , \U5/U20/Z , \U5/net2 , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr32bit_completion_10 ( o, i );
input  [63:0] i;
output o;
    wire \cd[3] , \cd[2] , \cd[1] , \cd[0] , ny, \U16/Z , nx, \U6/Z , \U15/Z ;
    chain_dr8bit_completion_44 U11 ( .o(\cd[3] ), .i({i[63], i[62], i[61], 
        i[60], i[59], i[58], i[57], i[56], i[31], i[30], i[29], i[28], i[27], 
        i[26], i[25], i[24]}) );
    chain_dr8bit_completion_47 U14 ( .o(\cd[2] ), .i({i[55], i[54], i[53], 
        i[52], i[51], i[50], i[49], i[48], i[23], i[22], i[21], i[20], i[19], 
        i[18], i[17], i[16]}) );
    chain_dr8bit_completion_46 U13 ( .o(\cd[1] ), .i({i[47], i[46], i[45], 
        i[44], i[43], i[42], i[41], i[40], i[15], i[14], i[13], i[12], i[11], 
        i[10], i[9], i[8]}) );
    chain_dr8bit_completion_45 U12 ( .o(\cd[0] ), .i({i[39], i[38], i[37], 
        i[36], i[35], i[34], i[33], i[32], i[7], i[6], i[5], i[4], i[3], i[2], 
        i[1], i[0]}) );
    aoi222_1 \U16/U30/U1  ( .x(ny), .a(\cd[0] ), .b(\cd[1] ), .c(\cd[0] ), .d(
        \U16/Z ), .e(\cd[1] ), .f(\U16/Z ) );
    inv_1 \U16/U30/Uinv  ( .x(\U16/Z ), .a(ny) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(ny), .b(nx), .c(ny), .d(\U6/Z ), .e(nx), 
        .f(\U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U15/U30/U1  ( .x(nx), .a(\cd[3] ), .b(\cd[2] ), .c(\cd[3] ), .d(
        \U15/Z ), .e(\cd[2] ), .f(\U15/Z ) );
    inv_1 \U15/U30/Uinv  ( .x(\U15/Z ), .a(nx) );
endmodule


module chain_selement_ga_65 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_trhdr_2 ( chainff_ack, chainh, chainl, eop, hdrack, normal_ack, 
    notify_ack, read_req, routereq, chain_ff_h, chainack, chainff_l, eopack, 
    err, nReset, normal_response, notify_accept, notify_defer, rcol_h, rcol_l, 
    read_ack, rnw_h, rnw_l, routeack, rsize_h, rsize_l, rtag_h, rtag_l );
output [7:0] chainh;
output [7:0] chainl;
input  [7:0] chain_ff_h;
input  [7:0] chainff_l;
input  [1:0] err;
input  [2:0] rcol_h;
input  [2:0] rcol_l;
input  [1:0] rsize_h;
input  [1:0] rsize_l;
input  [4:0] rtag_h;
input  [4:0] rtag_l;
input  chainack, eopack, nReset, normal_response, notify_accept, notify_defer, 
    read_ack, rnw_h, rnw_l, routeack;
output chainff_ack, eop, hdrack, normal_ack, notify_ack, read_req, routereq;
    wire done_eop, done_pl, \net413[15] , \hdr[16] , \hdr[0] , \net413[14] , 
        \hdr[17] , \hdr[1] , \net413[13] , \net413[12] , \net413[11] , 
        \net413[10] , \net413[9] , \net413[8] , \net413[7] , \net413[6] , 
        \net413[5] , \net413[4] , \net413[3] , \net413[2] , \net413[1] , 
        \net413[0] , net364, donotify, dowrite, net383, done_defer, done_write, 
        done_read, \net343[7] , \drive_l[0] , \net343[6] , \net343[5] , 
        \net343[3] , \net343[2] , \net343[1] , \net343[0] , net340, net337, 
        \net334[7] , \drive_l[1] , \net334[6] , \net334[4] , \net334[2] , 
        \net334[1] , \net334[0] , \net284[7] , \drive_h[1] , \net284[6] , 
        \net284[5] , \net284[4] , \net284[3] , \net284[2] , \net284[1] , 
        \net284[0] , \net288[7] , \drive_h[0] , \net288[6] , \net288[5] , 
        \net288[4] , \net288[3] , \net288[2] , \net288[1] , \net288[0] , 
        net332, done_accept, net321, net359, net362, ctrl_cd, \U311/nz[0] , 
        \U311/nz[1] , \U311/x[3] , \U311/U28/Z , \U311/x[0] , \U311/U32/Z , 
        \U311/x[5] , \U311/U20/Z , \U311/x[2] , \U311/U29/Z , \U311/x[7] , 
        \U311/U25/Z , \U311/y[0] , \U311/x[1] , \U311/U33/Z , \U311/y[2] , 
        \U311/x[4] , \U311/U21/Z , \U311/x[6] , \U311/U26/Z , \U311/y[1] , 
        \U311/U34/Z , \U311/U30/Z , \U311/U19/Z , \U311/y[3] , \U311/U27/Z , 
        \U311/U35/Z , \U311/U31/Z , net407, \U151/Z , done_hdr, 
        \U319/U21/U1/loop , \U323/U21/U1/loop , \U320/U21/U1/loop , 
        \U321/U21/U1/loop , \U322/U21/U1/loop , \U210/drivemonitor , 
        \U210/naa , \U210/net2 , \U210/net3 , net0230, \U210/bdone , 
        \U210/U1702/Z , \I0/drivemonitor , \I0/naa , \I0/net2 , \I0/net3 , 
        \I0/bdone , \I0/U1702/Z ;
    chain_selement_ga_65 U215 ( .Aa(done_eop), .Br(eop), .Ar(done_pl), .Ba(
        eopack) );
    nor2_1 \U308_0_/U5  ( .x(\net413[15] ), .a(\hdr[16] ), .b(\hdr[0] ) );
    nor2_1 \U308_1_/U5  ( .x(\net413[14] ), .a(\hdr[17] ), .b(\hdr[1] ) );
    nor2_1 \U308_2_/U5  ( .x(\net413[13] ), .a(1'b0), .b(routereq) );
    nor2_1 \U308_3_/U5  ( .x(\net413[12] ), .a(routereq), .b(1'b0) );
    nor2_1 \U308_4_/U5  ( .x(\net413[11] ), .a(1'b0), .b(routereq) );
    nor2_1 \U308_5_/U5  ( .x(\net413[10] ), .a(rnw_h), .b(rnw_l) );
    nor2_1 \U308_6_/U5  ( .x(\net413[9] ), .a(rsize_h[0]), .b(rsize_l[0]) );
    nor2_1 \U308_7_/U5  ( .x(\net413[8] ), .a(rsize_h[1]), .b(rsize_l[1]) );
    nor2_1 \U308_8_/U5  ( .x(\net413[7] ), .a(rtag_h[0]), .b(rtag_l[0]) );
    nor2_1 \U308_9_/U5  ( .x(\net413[6] ), .a(rtag_h[1]), .b(rtag_l[1]) );
    nor2_1 \U308_10_/U5  ( .x(\net413[5] ), .a(rtag_h[2]), .b(rtag_l[2]) );
    nor2_1 \U308_11_/U5  ( .x(\net413[4] ), .a(rtag_h[3]), .b(rtag_l[3]) );
    nor2_1 \U308_12_/U5  ( .x(\net413[3] ), .a(rtag_h[4]), .b(rtag_l[4]) );
    nor2_1 \U308_13_/U5  ( .x(\net413[2] ), .a(rcol_h[0]), .b(rcol_l[0]) );
    nor2_1 \U308_14_/U5  ( .x(\net413[1] ), .a(rcol_h[1]), .b(rcol_l[1]) );
    nor2_1 \U308_15_/U5  ( .x(\net413[0] ), .a(rcol_h[2]), .b(rcol_l[2]) );
    or3_1 \U257/U12  ( .x(net364), .a(donotify), .b(dowrite), .c(read_ack) );
    or3_1 \U297/U12  ( .x(net383), .a(done_defer), .b(done_write), .c(
        done_read) );
    and2_2 \U237/U8  ( .x(\hdr[1] ), .a(nReset), .b(normal_response) );
    and2_1 \U307_0_/U8  ( .x(\net343[7] ), .a(\drive_l[0] ), .b(\hdr[0] ) );
    and2_1 \U307_1_/U8  ( .x(\net343[6] ), .a(\drive_l[0] ), .b(\hdr[1] ) );
    and2_1 \U307_2_/U8  ( .x(\net343[5] ), .a(\drive_l[0] ), .b(routereq) );
    and2_1 \U307_4_/U8  ( .x(\net343[3] ), .a(\drive_l[0] ), .b(routereq) );
    and2_1 \U307_5_/U8  ( .x(\net343[2] ), .a(\drive_l[0] ), .b(rnw_l) );
    and2_1 \U307_6_/U8  ( .x(\net343[1] ), .a(\drive_l[0] ), .b(rsize_l[0]) );
    and2_1 \U307_7_/U8  ( .x(\net343[0] ), .a(\drive_l[0] ), .b(rsize_l[1]) );
    and2_1 \U235/U8  ( .x(net340), .a(err[1]), .b(nReset) );
    and2_1 \U236/U8  ( .x(net337), .a(nReset), .b(err[0]) );
    and2_1 \U306_0_/U8  ( .x(\net334[7] ), .a(\hdr[16] ), .b(\drive_l[1] ) );
    and2_1 \U306_1_/U8  ( .x(\net334[6] ), .a(\hdr[17] ), .b(\drive_l[1] ) );
    and2_1 \U306_3_/U8  ( .x(\net334[4] ), .a(routereq), .b(\drive_l[1] ) );
    and2_1 \U306_5_/U8  ( .x(\net334[2] ), .a(rnw_h), .b(\drive_l[1] ) );
    and2_1 \U306_6_/U8  ( .x(\net334[1] ), .a(rsize_h[0]), .b(\drive_l[1] ) );
    and2_1 \U306_7_/U8  ( .x(\net334[0] ), .a(rsize_h[1]), .b(\drive_l[1] ) );
    and2_1 \I1_0_/U8  ( .x(\net284[7] ), .a(rtag_h[0]), .b(\drive_h[1] ) );
    and2_1 \I1_1_/U8  ( .x(\net284[6] ), .a(rtag_h[1]), .b(\drive_h[1] ) );
    and2_1 \I1_2_/U8  ( .x(\net284[5] ), .a(rtag_h[2]), .b(\drive_h[1] ) );
    and2_1 \I1_3_/U8  ( .x(\net284[4] ), .a(rtag_h[3]), .b(\drive_h[1] ) );
    and2_1 \I1_4_/U8  ( .x(\net284[3] ), .a(rtag_h[4]), .b(\drive_h[1] ) );
    and2_1 \I1_5_/U8  ( .x(\net284[2] ), .a(rcol_h[0]), .b(\drive_h[1] ) );
    and2_1 \I1_6_/U8  ( .x(\net284[1] ), .a(rcol_h[1]), .b(\drive_h[1] ) );
    and2_1 \I1_7_/U8  ( .x(\net284[0] ), .a(rcol_h[2]), .b(\drive_h[1] ) );
    and2_1 \I2_0_/U8  ( .x(\net288[7] ), .a(\drive_h[0] ), .b(rtag_l[0]) );
    and2_1 \I2_1_/U8  ( .x(\net288[6] ), .a(\drive_h[0] ), .b(rtag_l[1]) );
    and2_1 \I2_2_/U8  ( .x(\net288[5] ), .a(\drive_h[0] ), .b(rtag_l[2]) );
    and2_1 \I2_3_/U8  ( .x(\net288[4] ), .a(\drive_h[0] ), .b(rtag_l[3]) );
    and2_1 \I2_4_/U8  ( .x(\net288[3] ), .a(\drive_h[0] ), .b(rtag_l[4]) );
    and2_1 \I2_5_/U8  ( .x(\net288[2] ), .a(\drive_h[0] ), .b(rcol_l[0]) );
    and2_1 \I2_6_/U8  ( .x(\net288[1] ), .a(\drive_h[0] ), .b(rcol_l[1]) );
    and2_1 \I2_7_/U8  ( .x(\net288[0] ), .a(\drive_h[0] ), .b(rcol_l[2]) );
    inv_1 \U318/U3  ( .x(net332), .a(routereq) );
    or2_4 \U255/U12  ( .x(notify_ack), .a(done_accept), .b(done_defer) );
    or2_4 \U228/U12  ( .x(\hdr[17] ), .a(notify_defer), .b(notify_accept) );
    or2_4 \U204/U12  ( .x(net321), .a(net359), .b(net362) );
    or2_4 \U221/U12  ( .x(\hdr[16] ), .a(net359), .b(notify_defer) );
    or2_4 \U252/U12  ( .x(normal_ack), .a(done_write), .b(done_read) );
    or2_4 \U280/U12  ( .x(\hdr[0] ), .a(net362), .b(notify_accept) );
    or2_4 \U317/U12  ( .x(routereq), .a(\hdr[17] ), .b(net321) );
    or3_4 \U309_0_/U12  ( .x(chainh[0]), .a(\net334[7] ), .b(\net284[7] ), .c(
        chain_ff_h[0]) );
    or3_4 \U309_1_/U12  ( .x(chainh[1]), .a(\net334[6] ), .b(\net284[6] ), .c(
        chain_ff_h[1]) );
    or3_4 \U309_3_/U12  ( .x(chainh[3]), .a(\net334[4] ), .b(\net284[4] ), .c(
        chain_ff_h[3]) );
    or3_4 \U309_5_/U12  ( .x(chainh[5]), .a(\net334[2] ), .b(\net284[2] ), .c(
        chain_ff_h[5]) );
    or3_4 \U309_6_/U12  ( .x(chainh[6]), .a(\net334[1] ), .b(\net284[1] ), .c(
        chain_ff_h[6]) );
    or3_4 \U309_7_/U12  ( .x(chainh[7]), .a(\net334[0] ), .b(\net284[0] ), .c(
        chain_ff_h[7]) );
    or3_4 \U310_0_/U12  ( .x(chainl[0]), .a(\net343[7] ), .b(\net288[7] ), .c(
        chainff_l[0]) );
    or3_4 \U310_1_/U12  ( .x(chainl[1]), .a(\net343[6] ), .b(\net288[6] ), .c(
        chainff_l[1]) );
    or3_4 \U310_2_/U12  ( .x(chainl[2]), .a(\net343[5] ), .b(\net288[5] ), .c(
        chainff_l[2]) );
    or3_4 \U310_4_/U12  ( .x(chainl[4]), .a(\net343[3] ), .b(\net288[3] ), .c(
        chainff_l[4]) );
    or3_4 \U310_5_/U12  ( .x(chainl[5]), .a(\net343[2] ), .b(\net288[2] ), .c(
        chainff_l[5]) );
    or3_4 \U310_6_/U12  ( .x(chainl[6]), .a(\net343[1] ), .b(\net288[1] ), .c(
        chainff_l[6]) );
    or3_4 \U310_7_/U12  ( .x(chainl[7]), .a(\net343[0] ), .b(\net288[0] ), .c(
        chainff_l[7]) );
    ao222_1 \U311/U37/U18/U1/U1  ( .x(ctrl_cd), .a(\U311/nz[0] ), .b(
        \U311/nz[1] ), .c(\U311/nz[0] ), .d(ctrl_cd), .e(\U311/nz[1] ), .f(
        ctrl_cd) );
    aoi222_1 \U311/U28/U30/U1  ( .x(\U311/x[3] ), .a(\net413[8] ), .b(
        \net413[9] ), .c(\net413[8] ), .d(\U311/U28/Z ), .e(\net413[9] ), .f(
        \U311/U28/Z ) );
    inv_1 \U311/U28/U30/Uinv  ( .x(\U311/U28/Z ), .a(\U311/x[3] ) );
    aoi222_1 \U311/U32/U30/U1  ( .x(\U311/x[0] ), .a(\net413[14] ), .b(
        \net413[15] ), .c(\net413[14] ), .d(\U311/U32/Z ), .e(\net413[15] ), 
        .f(\U311/U32/Z ) );
    inv_1 \U311/U32/U30/Uinv  ( .x(\U311/U32/Z ), .a(\U311/x[0] ) );
    aoi222_1 \U311/U20/U30/U1  ( .x(\U311/x[5] ), .a(\net413[4] ), .b(
        \net413[5] ), .c(\net413[4] ), .d(\U311/U20/Z ), .e(\net413[5] ), .f(
        \U311/U20/Z ) );
    inv_1 \U311/U20/U30/Uinv  ( .x(\U311/U20/Z ), .a(\U311/x[5] ) );
    aoi222_1 \U311/U29/U30/U1  ( .x(\U311/x[2] ), .a(\net413[10] ), .b(
        \net413[11] ), .c(\net413[10] ), .d(\U311/U29/Z ), .e(\net413[11] ), 
        .f(\U311/U29/Z ) );
    inv_1 \U311/U29/U30/Uinv  ( .x(\U311/U29/Z ), .a(\U311/x[2] ) );
    aoi222_1 \U311/U25/U30/U1  ( .x(\U311/x[7] ), .a(\net413[0] ), .b(
        \net413[1] ), .c(\net413[0] ), .d(\U311/U25/Z ), .e(\net413[1] ), .f(
        \U311/U25/Z ) );
    inv_1 \U311/U25/U30/Uinv  ( .x(\U311/U25/Z ), .a(\U311/x[7] ) );
    aoi222_1 \U311/U33/U30/U1  ( .x(\U311/y[0] ), .a(\U311/x[1] ), .b(
        \U311/x[0] ), .c(\U311/x[1] ), .d(\U311/U33/Z ), .e(\U311/x[0] ), .f(
        \U311/U33/Z ) );
    inv_1 \U311/U33/U30/Uinv  ( .x(\U311/U33/Z ), .a(\U311/y[0] ) );
    aoi222_1 \U311/U21/U30/U1  ( .x(\U311/y[2] ), .a(\U311/x[5] ), .b(
        \U311/x[4] ), .c(\U311/x[5] ), .d(\U311/U21/Z ), .e(\U311/x[4] ), .f(
        \U311/U21/Z ) );
    inv_1 \U311/U21/U30/Uinv  ( .x(\U311/U21/Z ), .a(\U311/y[2] ) );
    aoi222_1 \U311/U26/U30/U1  ( .x(\U311/x[6] ), .a(\net413[2] ), .b(
        \net413[3] ), .c(\net413[2] ), .d(\U311/U26/Z ), .e(\net413[3] ), .f(
        \U311/U26/Z ) );
    inv_1 \U311/U26/U30/Uinv  ( .x(\U311/U26/Z ), .a(\U311/x[6] ) );
    aoi222_1 \U311/U34/U30/U1  ( .x(\U311/nz[0] ), .a(\U311/y[1] ), .b(
        \U311/y[0] ), .c(\U311/y[1] ), .d(\U311/U34/Z ), .e(\U311/y[0] ), .f(
        \U311/U34/Z ) );
    inv_1 \U311/U34/U30/Uinv  ( .x(\U311/U34/Z ), .a(\U311/nz[0] ) );
    aoi222_1 \U311/U30/U30/U1  ( .x(\U311/y[1] ), .a(\U311/x[3] ), .b(
        \U311/x[2] ), .c(\U311/x[3] ), .d(\U311/U30/Z ), .e(\U311/x[2] ), .f(
        \U311/U30/Z ) );
    inv_1 \U311/U30/U30/Uinv  ( .x(\U311/U30/Z ), .a(\U311/y[1] ) );
    aoi222_1 \U311/U19/U30/U1  ( .x(\U311/x[4] ), .a(\net413[6] ), .b(
        \net413[7] ), .c(\net413[6] ), .d(\U311/U19/Z ), .e(\net413[7] ), .f(
        \U311/U19/Z ) );
    inv_1 \U311/U19/U30/Uinv  ( .x(\U311/U19/Z ), .a(\U311/x[4] ) );
    aoi222_1 \U311/U27/U30/U1  ( .x(\U311/y[3] ), .a(\U311/x[7] ), .b(
        \U311/x[6] ), .c(\U311/x[7] ), .d(\U311/U27/Z ), .e(\U311/x[6] ), .f(
        \U311/U27/Z ) );
    inv_1 \U311/U27/U30/Uinv  ( .x(\U311/U27/Z ), .a(\U311/y[3] ) );
    aoi222_1 \U311/U35/U30/U1  ( .x(\U311/nz[1] ), .a(\U311/y[3] ), .b(
        \U311/y[2] ), .c(\U311/y[3] ), .d(\U311/U35/Z ), .e(\U311/y[2] ), .f(
        \U311/U35/Z ) );
    inv_1 \U311/U35/U30/Uinv  ( .x(\U311/U35/Z ), .a(\U311/nz[1] ) );
    aoi222_1 \U311/U31/U30/U1  ( .x(\U311/x[1] ), .a(\net413[12] ), .b(
        \net413[13] ), .c(\net413[12] ), .d(\U311/U31/Z ), .e(\net413[13] ), 
        .f(\U311/U31/Z ) );
    inv_1 \U311/U31/U30/Uinv  ( .x(\U311/U31/Z ), .a(\U311/x[1] ) );
    aoi21_1 \U151/U30/U1/U1  ( .x(net407), .a(\U151/Z ), .b(chainff_ack), .c(
        net332) );
    inv_1 \U151/U30/U1/U2  ( .x(\U151/Z ), .a(net407) );
    ao222_1 \U324/U18/U1/U1  ( .x(hdrack), .a(ctrl_cd), .b(net383), .c(ctrl_cd
        ), .d(hdrack), .e(net383), .f(hdrack) );
    ao222_1 \U244/U18/U1/U1  ( .x(donotify), .a(done_hdr), .b(\hdr[17] ), .c(
        done_hdr), .d(donotify), .e(\hdr[17] ), .f(donotify) );
    ao222_1 \U260/U18/U1/U1  ( .x(net362), .a(net337), .b(\hdr[1] ), .c(net337
        ), .d(net362), .e(\hdr[1] ), .f(net362) );
    ao222_1 \U296/U18/U1/U1  ( .x(done_accept), .a(done_eop), .b(notify_accept
        ), .c(done_eop), .d(done_accept), .e(notify_accept), .f(done_accept)
         );
    ao222_1 \U261/U18/U1/U1  ( .x(net359), .a(net340), .b(\hdr[1] ), .c(net340
        ), .d(net359), .e(\hdr[1] ), .f(net359) );
    ao222_1 \U316/U18/U1/U1  ( .x(done_pl), .a(net364), .b(routeack), .c(
        net364), .d(done_pl), .e(routeack), .f(done_pl) );
    ao31_1 \U319/U21/U1/aoi  ( .x(\U319/U21/U1/loop ), .a(\hdr[1] ), .b(
        done_hdr), .c(rnw_h), .d(read_req) );
    oa21_1 \U319/U21/U1/outGate  ( .x(read_req), .a(\hdr[1] ), .b(done_hdr), 
        .c(\U319/U21/U1/loop ) );
    ao31_1 \U323/U21/U1/aoi  ( .x(\U323/U21/U1/loop ), .a(done_eop), .b(
        notify_defer), .c(ctrl_cd), .d(done_defer) );
    oa21_1 \U323/U21/U1/outGate  ( .x(done_defer), .a(done_eop), .b(
        notify_defer), .c(\U323/U21/U1/loop ) );
    ao31_1 \U320/U21/U1/aoi  ( .x(\U320/U21/U1/loop ), .a(\hdr[1] ), .b(
        done_hdr), .c(rnw_l), .d(dowrite) );
    oa21_1 \U320/U21/U1/outGate  ( .x(dowrite), .a(\hdr[1] ), .b(done_hdr), 
        .c(\U320/U21/U1/loop ) );
    ao31_1 \U321/U21/U1/aoi  ( .x(\U321/U21/U1/loop ), .a(read_req), .b(
        done_eop), .c(ctrl_cd), .d(done_read) );
    oa21_1 \U321/U21/U1/outGate  ( .x(done_read), .a(read_req), .b(done_eop), 
        .c(\U321/U21/U1/loop ) );
    ao31_1 \U322/U21/U1/aoi  ( .x(\U322/U21/U1/loop ), .a(dowrite), .b(
        done_eop), .c(ctrl_cd), .d(done_write) );
    oa21_1 \U322/U21/U1/outGate  ( .x(done_write), .a(dowrite), .b(done_eop), 
        .c(\U322/U21/U1/loop ) );
    nor2_2 \U210/U1703/U6  ( .x(done_hdr), .a(\U210/drivemonitor ), .b(
        \U210/naa ) );
    inv_2 \U210/U1699/U3  ( .x(\U210/net2 ), .a(\U210/net3 ) );
    and2_4 \U210/U2_0_/U8  ( .x(\drive_l[0] ), .a(net0230), .b(\U210/net2 ) );
    and2_4 \U210/U2_1_/U8  ( .x(\drive_l[1] ), .a(net0230), .b(\U210/net2 ) );
    inv_1 \U210/U1701/U3  ( .x(\U210/naa ), .a(\U210/bdone ) );
    ao222_1 \U210/U13/U18/U1/U1  ( .x(\U210/drivemonitor ), .a(\drive_l[1] ), 
        .b(\drive_l[0] ), .c(\drive_l[1] ), .d(\U210/drivemonitor ), .e(
        \drive_l[0] ), .f(\U210/drivemonitor ) );
    aoi21_1 \U210/U1702/U30/U1/U1  ( .x(\U210/bdone ), .a(\U210/U1702/Z ), .b(
        chainff_ack), .c(\U210/net2 ) );
    inv_1 \U210/U1702/U30/U1/U2  ( .x(\U210/U1702/Z ), .a(\U210/bdone ) );
    ao23_1 \U210/U1693/U21/U1/U1  ( .x(\U210/net3 ), .a(net0230), .b(
        \U210/net3 ), .c(net0230), .d(\U210/drivemonitor ), .e(chainff_ack) );
    nor2_2 \I0/U1703/U6  ( .x(net0230), .a(\I0/drivemonitor ), .b(\I0/naa ) );
    inv_2 \I0/U1699/U3  ( .x(\I0/net2 ), .a(\I0/net3 ) );
    and2_4 \I0/U2_0_/U8  ( .x(\drive_h[0] ), .a(net407), .b(\I0/net2 ) );
    and2_4 \I0/U2_1_/U8  ( .x(\drive_h[1] ), .a(net407), .b(\I0/net2 ) );
    inv_1 \I0/U1701/U3  ( .x(\I0/naa ), .a(\I0/bdone ) );
    ao222_1 \I0/U13/U18/U1/U1  ( .x(\I0/drivemonitor ), .a(\drive_h[1] ), .b(
        \drive_h[0] ), .c(\drive_h[1] ), .d(\I0/drivemonitor ), .e(
        \drive_h[0] ), .f(\I0/drivemonitor ) );
    aoi21_1 \I0/U1702/U30/U1/U1  ( .x(\I0/bdone ), .a(\I0/U1702/Z ), .b(
        chainff_ack), .c(\I0/net2 ) );
    inv_1 \I0/U1702/U30/U1/U2  ( .x(\I0/U1702/Z ), .a(\I0/bdone ) );
    ao23_1 \I0/U1693/U21/U1/U1  ( .x(\I0/net3 ), .a(net407), .b(\I0/net3 ), 
        .c(net407), .d(\I0/drivemonitor ), .e(chainff_ack) );
    buf_3 U1 ( .x(chainff_ack), .a(chainack) );
    or2_1 U2 ( .x(chainh[4]), .a(chain_ff_h[4]), .b(\net284[3] ) );
    or2_1 U3 ( .x(chainh[2]), .a(chain_ff_h[2]), .b(\net284[5] ) );
    or2_1 U4 ( .x(chainl[3]), .a(chainff_l[3]), .b(\net288[4] ) );
endmodule


module chain_dr2fr_byte_5 ( eop_ack, ia, o, eop, ih, il, nReset, noa );
output [4:0] o;
input  [7:0] ih;
input  [7:0] il;
input  eop, nReset, noa;
output eop_ack, ia;
    wire eop_ack_wire, nbReset, eop_pass, nxa, naa, nlowack, \twobitack[0] , 
        \twobitack[1] , nhighack, \twobitack[2] , \twobitack[3] , \U1018/Z , 
        \U1270/net189 , \U1270/net192 , \U1270/net191 , net199, \U1270/net190 , 
        \U1270/U1141/Z , \U1268/net189 , \U1268/net192 , \U1268/net191 , 
        net194, \U1268/net190 , \U1268/U1141/Z , \U1224/nack[0] , \x[3] , 
        \x[2] , \U1224/nack[1] , \x[1] , \U1224/net4 , \x[0] , 
        \U1224/U1125/U28/U1/clr , asel, \U1224/U1125/U28/U1/set , 
        \U1224/U1122/U28/U1/clr , csel, nca, \U1224/U1122/U28/U1/set , 
        \U1224/U916_0_/U25/U1/clr , \a[0] , \c[0] , \U1224/U916_0_/U25/U1/ob , 
        \U1224/U916_1_/U25/U1/clr , \a[1] , \c[1] , \U1224/U916_1_/U25/U1/ob , 
        \U1224/U916_2_/U25/U1/clr , \a[2] , \c[2] , \U1224/U916_2_/U25/U1/ob , 
        \U1224/U916_3_/U25/U1/clr , \a[3] , \c[3] , \U1224/U916_3_/U25/U1/ob , 
        \U1209/nack[0] , \U1209/nack[1] , \U1209/net4 , 
        \U1209/U1125/U28/U1/clr , xsel, \U1209/U1125/U28/U1/set , 
        \U1209/U1122/U28/U1/clr , ysel, nyla, \U1209/U1122/U28/U1/set , 
        \U1209/U916_0_/U25/U1/clr , \yl[0] , \U1209/U916_0_/U25/U1/ob , 
        \U1209/U916_1_/U25/U1/clr , \yl[1] , \U1209/U916_1_/U25/U1/ob , 
        \U1209/U916_2_/U25/U1/clr , \yl[2] , \U1209/U916_2_/U25/U1/ob , 
        \U1209/U916_3_/U25/U1/clr , \yl[3] , \U1209/U916_3_/U25/U1/ob , 
        \U1213/nack[0] , \y[3] , \y[2] , \U1213/nack[1] , \y[1] , \U1213/net4 , 
        \y[0] , \U1213/U1125/U28/U1/clr , bsel, nba, \U1213/U1125/U28/U1/set , 
        \U1213/U1122/U28/U1/clr , dsel, nda, \U1213/U1122/U28/U1/set , 
        \U1213/U916_0_/U25/U1/clr , nya, \b[0] , \d[0] , 
        \U1213/U916_0_/U25/U1/ob , \U1213/U916_1_/U25/U1/clr , \b[1] , \d[1] , 
        \U1213/U916_1_/U25/U1/ob , \U1213/U916_2_/U25/U1/clr , \b[2] , \d[2] , 
        \U1213/U916_2_/U25/U1/ob , \U1213/U916_3_/U25/U1/clr , \b[3] , \d[3] , 
        \U1213/U916_3_/U25/U1/ob , \cdh[0] , \cdh[1] , \cdl[0] , \cdl[1] , 
        \cdh[2] , \cdh[3] , \cdl[2] , \cdl[3] , cg, \U1296/ng , net195, 
        \U1296/U1384/Z , \U1296/U1386/U25/U1/clr , \U1296/U1386/U25/U1/ob , dg, 
        \U1298/ng , net193, \U1298/U1384/Z , \U1298/U1386/U25/U1/clr , 
        \U1298/U1386/U25/U1/ob , bg, \U1306/ng , \U1306/U1384/Z , 
        \U1306/U1386/U25/U1/clr , \U1306/U1386/U25/U1/ob , ag, \U1295/ng , 
        \U1295/U1384/Z , \U1295/U1386/U25/U1/clr , \U1295/U1386/U25/U1/ob , 
        \U1297/s , \U1297/r , \U1297/nback , \U1297/naack , \U1297/reset , 
        \U1297/U1128/U28/U1/clr , \U1297/U1128/U28/U1/set , 
        \U1297/U1127/U28/U1/clr , \U1297/U1127/U28/U1/set , \U1300/s , 
        \U1300/r , \U1300/nback , \U1300/naack , \U1300/reset , 
        \U1300/U1128/U28/U1/clr , \U1300/U1128/U28/U1/set , 
        \U1300/U1127/U28/U1/clr , \U1300/U1127/U28/U1/set , 
        \U1289/U1150/U28/U1/clr , \U1289/bnreset , \U1289/U1150/U28/U1/set , 
        \U1289/U1152/U28/U1/clr , \U1289/U1152/U28/U1/set , 
        \U1289/U1149/U28/U1/clr , \U1289/U1149/U28/U1/set , 
        \U1289/U1151/U28/U1/clr , \U1289/U1151/U28/U1/set , 
        \U1289/U1148/net189 , \U1289/U1148/net192 , \U1289/U1148/net191 , 
        \U1289/U1148/net190 , \U1289/U1148/U1141/Z , \U1271/U1150/U28/U1/clr , 
        \U1271/bnreset , \U1271/U1150/U28/U1/set , \U1271/U1152/U28/U1/clr , 
        \U1271/U1152/U28/U1/set , \U1271/U1149/U28/U1/clr , 
        \U1271/U1149/U28/U1/set , \U1271/U1151/U28/U1/clr , 
        \U1271/U1151/U28/U1/set , \U1271/U1148/net189 , \U1271/U1148/net192 , 
        \U1271/U1148/net191 , \U1271/U1148/net190 , \U1271/U1148/U1141/Z , 
        \U1225/s , \U1225/r , \U1225/nback , \U1225/naack , \U1225/reset , 
        \U1308/nack[1] , \U1308/nack[0] ;
    assign eop_ack = eop_ack_wire;
    assign o[4] = eop_ack_wire;
    buf_2 U1231 ( .x(nbReset), .a(nReset) );
    and3_1 \U1194/U9  ( .x(eop_pass), .a(nxa), .b(naa), .c(eop) );
    ao222_1 \U1301/U18/U1/U1  ( .x(nlowack), .a(\twobitack[0] ), .b(
        \twobitack[1] ), .c(\twobitack[0] ), .d(nlowack), .e(\twobitack[1] ), 
        .f(nlowack) );
    ao222_1 \U1302/U18/U1/U1  ( .x(nhighack), .a(\twobitack[2] ), .b(
        \twobitack[3] ), .c(\twobitack[2] ), .d(nhighack), .e(\twobitack[3] ), 
        .f(nhighack) );
    aoi222_1 \U1018/U30/U1  ( .x(ia), .a(nhighack), .b(nlowack), .c(nhighack), 
        .d(\U1018/Z ), .e(nlowack), .f(\U1018/Z ) );
    inv_1 \U1018/U30/Uinv  ( .x(\U1018/Z ), .a(ia) );
    ao222_2 \U1038/U19/U1/U1  ( .x(eop_ack_wire), .a(eop_pass), .b(noa), .c(
        eop_pass), .d(eop_ack_wire), .e(noa), .f(eop_ack_wire) );
    inv_1 \U1270/U1147/U3  ( .x(\U1270/net189 ), .a(nbReset) );
    nor2_1 \U1270/U582/U5  ( .x(\U1270/net192 ), .a(il[4]), .b(ih[4]) );
    nor2_1 \U1270/U580/U5  ( .x(\U1270/net191 ), .a(il[5]), .b(ih[5]) );
    nor2_2 \U1270/U1146/U6  ( .x(net199), .a(\U1270/net190 ), .b(
        \U1270/net189 ) );
    aoi222_1 \U1270/U1141/U30/U1  ( .x(\U1270/net190 ), .a(\U1270/net191 ), 
        .b(\U1270/net192 ), .c(\U1270/net191 ), .d(\U1270/U1141/Z ), .e(
        \U1270/net192 ), .f(\U1270/U1141/Z ) );
    inv_1 \U1270/U1141/U30/Uinv  ( .x(\U1270/U1141/Z ), .a(\U1270/net190 ) );
    inv_1 \U1268/U1147/U3  ( .x(\U1268/net189 ), .a(nbReset) );
    nor2_1 \U1268/U582/U5  ( .x(\U1268/net192 ), .a(il[6]), .b(ih[6]) );
    nor2_1 \U1268/U580/U5  ( .x(\U1268/net191 ), .a(il[7]), .b(ih[7]) );
    nor2_2 \U1268/U1146/U6  ( .x(net194), .a(\U1268/net190 ), .b(
        \U1268/net189 ) );
    aoi222_1 \U1268/U1141/U30/U1  ( .x(\U1268/net190 ), .a(\U1268/net191 ), 
        .b(\U1268/net192 ), .c(\U1268/net191 ), .d(\U1268/U1141/Z ), .e(
        \U1268/net192 ), .f(\U1268/U1141/Z ) );
    inv_1 \U1268/U1141/U30/Uinv  ( .x(\U1268/U1141/Z ), .a(\U1268/net190 ) );
    nor2_1 \U1224/U1128/U5  ( .x(\U1224/nack[0] ), .a(\x[3] ), .b(\x[2] ) );
    nor3_1 \U1224/U1127/U7  ( .x(\U1224/nack[1] ), .a(\x[1] ), .b(\U1224/net4 
        ), .c(\x[0] ) );
    inv_1 \U1224/U907/U3  ( .x(\U1224/net4 ), .a(nbReset) );
    aoai211_1 \U1224/U1125/U28/U1/U1  ( .x(\U1224/U1125/U28/U1/clr ), .a(
        \U1224/nack[1] ), .b(\U1224/nack[0] ), .c(asel), .d(naa) );
    nand3_1 \U1224/U1125/U28/U1/U2  ( .x(\U1224/U1125/U28/U1/set ), .a(asel), 
        .b(\U1224/nack[1] ), .c(\U1224/nack[0] ) );
    nand2_2 \U1224/U1125/U28/U1/U3  ( .x(naa), .a(\U1224/U1125/U28/U1/clr ), 
        .b(\U1224/U1125/U28/U1/set ) );
    aoai211_1 \U1224/U1122/U28/U1/U1  ( .x(\U1224/U1122/U28/U1/clr ), .a(
        \U1224/nack[0] ), .b(\U1224/nack[1] ), .c(csel), .d(nca) );
    nand3_1 \U1224/U1122/U28/U1/U2  ( .x(\U1224/U1122/U28/U1/set ), .a(csel), 
        .b(\U1224/nack[0] ), .c(\U1224/nack[1] ) );
    nand2_2 \U1224/U1122/U28/U1/U3  ( .x(nca), .a(\U1224/U1122/U28/U1/clr ), 
        .b(\U1224/U1122/U28/U1/set ) );
    oa31_1 \U1224/U916_0_/U25/U1/Uclr  ( .x(\U1224/U916_0_/U25/U1/clr ), .a(
        nxa), .b(\a[0] ), .c(\c[0] ), .d(\x[0] ) );
    oaoi211_1 \U1224/U916_0_/U25/U1/Uaoi  ( .x(\U1224/U916_0_/U25/U1/ob ), .a(
        \a[0] ), .b(\c[0] ), .c(nxa), .d(\U1224/U916_0_/U25/U1/clr ) );
    inv_2 \U1224/U916_0_/U25/U1/Ui  ( .x(\x[0] ), .a(\U1224/U916_0_/U25/U1/ob 
        ) );
    oa31_1 \U1224/U916_1_/U25/U1/Uclr  ( .x(\U1224/U916_1_/U25/U1/clr ), .a(
        nxa), .b(\a[1] ), .c(\c[1] ), .d(\x[1] ) );
    oaoi211_1 \U1224/U916_1_/U25/U1/Uaoi  ( .x(\U1224/U916_1_/U25/U1/ob ), .a(
        \a[1] ), .b(\c[1] ), .c(nxa), .d(\U1224/U916_1_/U25/U1/clr ) );
    inv_2 \U1224/U916_1_/U25/U1/Ui  ( .x(\x[1] ), .a(\U1224/U916_1_/U25/U1/ob 
        ) );
    oa31_1 \U1224/U916_2_/U25/U1/Uclr  ( .x(\U1224/U916_2_/U25/U1/clr ), .a(
        nxa), .b(\a[2] ), .c(\c[2] ), .d(\x[2] ) );
    oaoi211_1 \U1224/U916_2_/U25/U1/Uaoi  ( .x(\U1224/U916_2_/U25/U1/ob ), .a(
        \a[2] ), .b(\c[2] ), .c(nxa), .d(\U1224/U916_2_/U25/U1/clr ) );
    inv_2 \U1224/U916_2_/U25/U1/Ui  ( .x(\x[2] ), .a(\U1224/U916_2_/U25/U1/ob 
        ) );
    oa31_1 \U1224/U916_3_/U25/U1/Uclr  ( .x(\U1224/U916_3_/U25/U1/clr ), .a(
        nxa), .b(\a[3] ), .c(\c[3] ), .d(\x[3] ) );
    oaoi211_1 \U1224/U916_3_/U25/U1/Uaoi  ( .x(\U1224/U916_3_/U25/U1/ob ), .a(
        \a[3] ), .b(\c[3] ), .c(nxa), .d(\U1224/U916_3_/U25/U1/clr ) );
    inv_2 \U1224/U916_3_/U25/U1/Ui  ( .x(\x[3] ), .a(\U1224/U916_3_/U25/U1/ob 
        ) );
    nor2_1 \U1209/U1128/U5  ( .x(\U1209/nack[0] ), .a(o[3]), .b(o[2]) );
    nor3_1 \U1209/U1127/U7  ( .x(\U1209/nack[1] ), .a(o[1]), .b(\U1209/net4 ), 
        .c(o[0]) );
    inv_1 \U1209/U907/U3  ( .x(\U1209/net4 ), .a(nbReset) );
    aoai211_1 \U1209/U1125/U28/U1/U1  ( .x(\U1209/U1125/U28/U1/clr ), .a(
        \U1209/nack[1] ), .b(\U1209/nack[0] ), .c(xsel), .d(nxa) );
    nand3_1 \U1209/U1125/U28/U1/U2  ( .x(\U1209/U1125/U28/U1/set ), .a(xsel), 
        .b(\U1209/nack[1] ), .c(\U1209/nack[0] ) );
    nand2_2 \U1209/U1125/U28/U1/U3  ( .x(nxa), .a(\U1209/U1125/U28/U1/clr ), 
        .b(\U1209/U1125/U28/U1/set ) );
    aoai211_1 \U1209/U1122/U28/U1/U1  ( .x(\U1209/U1122/U28/U1/clr ), .a(
        \U1209/nack[0] ), .b(\U1209/nack[1] ), .c(ysel), .d(nyla) );
    nand3_1 \U1209/U1122/U28/U1/U2  ( .x(\U1209/U1122/U28/U1/set ), .a(ysel), 
        .b(\U1209/nack[0] ), .c(\U1209/nack[1] ) );
    nand2_2 \U1209/U1122/U28/U1/U3  ( .x(nyla), .a(\U1209/U1122/U28/U1/clr ), 
        .b(\U1209/U1122/U28/U1/set ) );
    oa31_1 \U1209/U916_0_/U25/U1/Uclr  ( .x(\U1209/U916_0_/U25/U1/clr ), .a(
        noa), .b(\x[0] ), .c(\yl[0] ), .d(o[0]) );
    oaoi211_1 \U1209/U916_0_/U25/U1/Uaoi  ( .x(\U1209/U916_0_/U25/U1/ob ), .a(
        \x[0] ), .b(\yl[0] ), .c(noa), .d(\U1209/U916_0_/U25/U1/clr ) );
    inv_2 \U1209/U916_0_/U25/U1/Ui  ( .x(o[0]), .a(\U1209/U916_0_/U25/U1/ob )
         );
    oa31_1 \U1209/U916_1_/U25/U1/Uclr  ( .x(\U1209/U916_1_/U25/U1/clr ), .a(
        noa), .b(\x[1] ), .c(\yl[1] ), .d(o[1]) );
    oaoi211_1 \U1209/U916_1_/U25/U1/Uaoi  ( .x(\U1209/U916_1_/U25/U1/ob ), .a(
        \x[1] ), .b(\yl[1] ), .c(noa), .d(\U1209/U916_1_/U25/U1/clr ) );
    inv_2 \U1209/U916_1_/U25/U1/Ui  ( .x(o[1]), .a(\U1209/U916_1_/U25/U1/ob )
         );
    oa31_1 \U1209/U916_2_/U25/U1/Uclr  ( .x(\U1209/U916_2_/U25/U1/clr ), .a(
        noa), .b(\x[2] ), .c(\yl[2] ), .d(o[2]) );
    oaoi211_1 \U1209/U916_2_/U25/U1/Uaoi  ( .x(\U1209/U916_2_/U25/U1/ob ), .a(
        \x[2] ), .b(\yl[2] ), .c(noa), .d(\U1209/U916_2_/U25/U1/clr ) );
    inv_2 \U1209/U916_2_/U25/U1/Ui  ( .x(o[2]), .a(\U1209/U916_2_/U25/U1/ob )
         );
    oa31_1 \U1209/U916_3_/U25/U1/Uclr  ( .x(\U1209/U916_3_/U25/U1/clr ), .a(
        noa), .b(\x[3] ), .c(\yl[3] ), .d(o[3]) );
    oaoi211_1 \U1209/U916_3_/U25/U1/Uaoi  ( .x(\U1209/U916_3_/U25/U1/ob ), .a(
        \x[3] ), .b(\yl[3] ), .c(noa), .d(\U1209/U916_3_/U25/U1/clr ) );
    inv_2 \U1209/U916_3_/U25/U1/Ui  ( .x(o[3]), .a(\U1209/U916_3_/U25/U1/ob )
         );
    nor2_1 \U1213/U1128/U5  ( .x(\U1213/nack[0] ), .a(\y[3] ), .b(\y[2] ) );
    nor3_1 \U1213/U1127/U7  ( .x(\U1213/nack[1] ), .a(\y[1] ), .b(\U1213/net4 
        ), .c(\y[0] ) );
    inv_1 \U1213/U907/U3  ( .x(\U1213/net4 ), .a(nbReset) );
    aoai211_1 \U1213/U1125/U28/U1/U1  ( .x(\U1213/U1125/U28/U1/clr ), .a(
        \U1213/nack[1] ), .b(\U1213/nack[0] ), .c(bsel), .d(nba) );
    nand3_1 \U1213/U1125/U28/U1/U2  ( .x(\U1213/U1125/U28/U1/set ), .a(bsel), 
        .b(\U1213/nack[1] ), .c(\U1213/nack[0] ) );
    nand2_2 \U1213/U1125/U28/U1/U3  ( .x(nba), .a(\U1213/U1125/U28/U1/clr ), 
        .b(\U1213/U1125/U28/U1/set ) );
    aoai211_1 \U1213/U1122/U28/U1/U1  ( .x(\U1213/U1122/U28/U1/clr ), .a(
        \U1213/nack[0] ), .b(\U1213/nack[1] ), .c(dsel), .d(nda) );
    nand3_1 \U1213/U1122/U28/U1/U2  ( .x(\U1213/U1122/U28/U1/set ), .a(dsel), 
        .b(\U1213/nack[0] ), .c(\U1213/nack[1] ) );
    nand2_2 \U1213/U1122/U28/U1/U3  ( .x(nda), .a(\U1213/U1122/U28/U1/clr ), 
        .b(\U1213/U1122/U28/U1/set ) );
    oa31_1 \U1213/U916_0_/U25/U1/Uclr  ( .x(\U1213/U916_0_/U25/U1/clr ), .a(
        nya), .b(\b[0] ), .c(\d[0] ), .d(\y[0] ) );
    oaoi211_1 \U1213/U916_0_/U25/U1/Uaoi  ( .x(\U1213/U916_0_/U25/U1/ob ), .a(
        \b[0] ), .b(\d[0] ), .c(nya), .d(\U1213/U916_0_/U25/U1/clr ) );
    inv_2 \U1213/U916_0_/U25/U1/Ui  ( .x(\y[0] ), .a(\U1213/U916_0_/U25/U1/ob 
        ) );
    oa31_1 \U1213/U916_1_/U25/U1/Uclr  ( .x(\U1213/U916_1_/U25/U1/clr ), .a(
        nya), .b(\b[1] ), .c(\d[1] ), .d(\y[1] ) );
    oaoi211_1 \U1213/U916_1_/U25/U1/Uaoi  ( .x(\U1213/U916_1_/U25/U1/ob ), .a(
        \b[1] ), .b(\d[1] ), .c(nya), .d(\U1213/U916_1_/U25/U1/clr ) );
    inv_2 \U1213/U916_1_/U25/U1/Ui  ( .x(\y[1] ), .a(\U1213/U916_1_/U25/U1/ob 
        ) );
    oa31_1 \U1213/U916_2_/U25/U1/Uclr  ( .x(\U1213/U916_2_/U25/U1/clr ), .a(
        nya), .b(\b[2] ), .c(\d[2] ), .d(\y[2] ) );
    oaoi211_1 \U1213/U916_2_/U25/U1/Uaoi  ( .x(\U1213/U916_2_/U25/U1/ob ), .a(
        \b[2] ), .b(\d[2] ), .c(nya), .d(\U1213/U916_2_/U25/U1/clr ) );
    inv_2 \U1213/U916_2_/U25/U1/Ui  ( .x(\y[2] ), .a(\U1213/U916_2_/U25/U1/ob 
        ) );
    oa31_1 \U1213/U916_3_/U25/U1/Uclr  ( .x(\U1213/U916_3_/U25/U1/clr ), .a(
        nya), .b(\b[3] ), .c(\d[3] ), .d(\y[3] ) );
    oaoi211_1 \U1213/U916_3_/U25/U1/Uaoi  ( .x(\U1213/U916_3_/U25/U1/ob ), .a(
        \b[3] ), .b(\d[3] ), .c(nya), .d(\U1213/U916_3_/U25/U1/clr ) );
    inv_2 \U1213/U916_3_/U25/U1/Ui  ( .x(\y[3] ), .a(\U1213/U916_3_/U25/U1/ob 
        ) );
    and3_2 \U1210/U1138/U9  ( .x(\d[3] ), .a(\cdh[0] ), .b(nda), .c(\cdh[1] )
         );
    and3_2 \U1210/U1137/U9  ( .x(\d[2] ), .a(\cdl[0] ), .b(nda), .c(\cdh[1] )
         );
    and3_2 \U1210/U1139/U9  ( .x(\d[1] ), .a(\cdh[0] ), .b(nda), .c(\cdl[1] )
         );
    and3_2 \U1210/U1136/U9  ( .x(\d[0] ), .a(\cdl[0] ), .b(nda), .c(\cdl[1] )
         );
    and3_2 \U1162/U1138/U9  ( .x(\a[3] ), .a(ih[6]), .b(naa), .c(ih[7]) );
    and3_2 \U1162/U1137/U9  ( .x(\a[2] ), .a(il[6]), .b(naa), .c(ih[7]) );
    and3_2 \U1162/U1139/U9  ( .x(\a[1] ), .a(ih[6]), .b(naa), .c(il[7]) );
    and3_2 \U1162/U1136/U9  ( .x(\a[0] ), .a(il[6]), .b(naa), .c(il[7]) );
    and3_2 \U1211/U1138/U9  ( .x(\b[3] ), .a(ih[4]), .b(nba), .c(ih[5]) );
    and3_2 \U1211/U1137/U9  ( .x(\b[2] ), .a(il[4]), .b(nba), .c(ih[5]) );
    and3_2 \U1211/U1139/U9  ( .x(\b[1] ), .a(ih[4]), .b(nba), .c(il[5]) );
    and3_2 \U1211/U1136/U9  ( .x(\b[0] ), .a(il[4]), .b(nba), .c(il[5]) );
    and3_2 \U1163/U1138/U9  ( .x(\c[3] ), .a(\cdh[2] ), .b(nca), .c(\cdh[3] )
         );
    and3_2 \U1163/U1137/U9  ( .x(\c[2] ), .a(\cdl[2] ), .b(nca), .c(\cdh[3] )
         );
    and3_2 \U1163/U1139/U9  ( .x(\c[1] ), .a(\cdh[2] ), .b(nca), .c(\cdl[3] )
         );
    and3_2 \U1163/U1136/U9  ( .x(\c[0] ), .a(\cdl[2] ), .b(nca), .c(\cdl[3] )
         );
    and2_1 \U1296/U1385/U8  ( .x(cg), .a(nbReset), .b(\U1296/ng ) );
    aoi222_1 \U1296/U1384/U30/U1  ( .x(\U1296/ng ), .a(nca), .b(net195), .c(
        nca), .d(\U1296/U1384/Z ), .e(net195), .f(\U1296/U1384/Z ) );
    inv_1 \U1296/U1384/U30/Uinv  ( .x(\U1296/U1384/Z ), .a(\U1296/ng ) );
    oa31_1 \U1296/U1386/U25/U1/Uclr  ( .x(\U1296/U1386/U25/U1/clr ), .a(
        \twobitack[2] ), .b(cg), .c(nca), .d(net195) );
    oaoi211_1 \U1296/U1386/U25/U1/Uaoi  ( .x(\U1296/U1386/U25/U1/ob ), .a(cg), 
        .b(nca), .c(\twobitack[2] ), .d(\U1296/U1386/U25/U1/clr ) );
    inv_2 \U1296/U1386/U25/U1/Ui  ( .x(net195), .a(\U1296/U1386/U25/U1/ob ) );
    and2_1 \U1298/U1385/U8  ( .x(dg), .a(nbReset), .b(\U1298/ng ) );
    aoi222_1 \U1298/U1384/U30/U1  ( .x(\U1298/ng ), .a(nda), .b(net193), .c(
        nda), .d(\U1298/U1384/Z ), .e(net193), .f(\U1298/U1384/Z ) );
    inv_1 \U1298/U1384/U30/Uinv  ( .x(\U1298/U1384/Z ), .a(\U1298/ng ) );
    oa31_1 \U1298/U1386/U25/U1/Uclr  ( .x(\U1298/U1386/U25/U1/clr ), .a(
        \twobitack[0] ), .b(dg), .c(nda), .d(net193) );
    oaoi211_1 \U1298/U1386/U25/U1/Uaoi  ( .x(\U1298/U1386/U25/U1/ob ), .a(dg), 
        .b(nda), .c(\twobitack[0] ), .d(\U1298/U1386/U25/U1/clr ) );
    inv_2 \U1298/U1386/U25/U1/Ui  ( .x(net193), .a(\U1298/U1386/U25/U1/ob ) );
    and2_1 \U1306/U1385/U8  ( .x(bg), .a(nbReset), .b(\U1306/ng ) );
    aoi222_1 \U1306/U1384/U30/U1  ( .x(\U1306/ng ), .a(nba), .b(\twobitack[1] 
        ), .c(nba), .d(\U1306/U1384/Z ), .e(\twobitack[1] ), .f(
        \U1306/U1384/Z ) );
    inv_1 \U1306/U1384/U30/Uinv  ( .x(\U1306/U1384/Z ), .a(\U1306/ng ) );
    oa31_1 \U1306/U1386/U25/U1/Uclr  ( .x(\U1306/U1386/U25/U1/clr ), .a(net199
        ), .b(bg), .c(nba), .d(\twobitack[1] ) );
    oaoi211_1 \U1306/U1386/U25/U1/Uaoi  ( .x(\U1306/U1386/U25/U1/ob ), .a(bg), 
        .b(nba), .c(net199), .d(\U1306/U1386/U25/U1/clr ) );
    inv_2 \U1306/U1386/U25/U1/Ui  ( .x(\twobitack[1] ), .a(
        \U1306/U1386/U25/U1/ob ) );
    and2_1 \U1295/U1385/U8  ( .x(ag), .a(nbReset), .b(\U1295/ng ) );
    aoi222_1 \U1295/U1384/U30/U1  ( .x(\U1295/ng ), .a(naa), .b(\twobitack[3] 
        ), .c(naa), .d(\U1295/U1384/Z ), .e(\twobitack[3] ), .f(
        \U1295/U1384/Z ) );
    inv_1 \U1295/U1384/U30/Uinv  ( .x(\U1295/U1384/Z ), .a(\U1295/ng ) );
    oa31_1 \U1295/U1386/U25/U1/Uclr  ( .x(\U1295/U1386/U25/U1/clr ), .a(net194
        ), .b(ag), .c(naa), .d(\twobitack[3] ) );
    oaoi211_1 \U1295/U1386/U25/U1/Uaoi  ( .x(\U1295/U1386/U25/U1/ob ), .a(ag), 
        .b(naa), .c(net194), .d(\U1295/U1386/U25/U1/clr ) );
    inv_2 \U1295/U1386/U25/U1/Ui  ( .x(\twobitack[3] ), .a(
        \U1295/U1386/U25/U1/ob ) );
    nand2_1 \U1297/U1131/U5  ( .x(\U1297/s ), .a(\U1297/r ), .b(\U1297/nback )
         );
    nand2_1 \U1297/U1103/U5  ( .x(\U1297/r ), .a(\U1297/naack ), .b(\U1297/s )
         );
    inv_1 \U1297/U1111/U3  ( .x(\U1297/reset ), .a(nbReset) );
    inv_1 \U1297/U1112/U3  ( .x(\U1297/naack ), .a(naa) );
    nor2_1 \U1297/U1130/U5  ( .x(\U1297/nback ), .a(nca), .b(\U1297/reset ) );
    aoai211_1 \U1297/U1128/U28/U1/U1  ( .x(\U1297/U1128/U28/U1/clr ), .a(
        \U1297/r ), .b(\U1297/naack ), .c(cg), .d(csel) );
    nand3_1 \U1297/U1128/U28/U1/U2  ( .x(\U1297/U1128/U28/U1/set ), .a(cg), 
        .b(\U1297/r ), .c(\U1297/naack ) );
    nand2_2 \U1297/U1128/U28/U1/U3  ( .x(csel), .a(\U1297/U1128/U28/U1/clr ), 
        .b(\U1297/U1128/U28/U1/set ) );
    aoai211_1 \U1297/U1127/U28/U1/U1  ( .x(\U1297/U1127/U28/U1/clr ), .a(
        \U1297/s ), .b(\U1297/nback ), .c(ag), .d(asel) );
    nand3_1 \U1297/U1127/U28/U1/U2  ( .x(\U1297/U1127/U28/U1/set ), .a(ag), 
        .b(\U1297/s ), .c(\U1297/nback ) );
    nand2_2 \U1297/U1127/U28/U1/U3  ( .x(asel), .a(\U1297/U1127/U28/U1/clr ), 
        .b(\U1297/U1127/U28/U1/set ) );
    nand2_1 \U1300/U1131/U5  ( .x(\U1300/s ), .a(\U1300/r ), .b(\U1300/nback )
         );
    nand2_1 \U1300/U1103/U5  ( .x(\U1300/r ), .a(\U1300/naack ), .b(\U1300/s )
         );
    inv_1 \U1300/U1111/U3  ( .x(\U1300/reset ), .a(nbReset) );
    inv_1 \U1300/U1112/U3  ( .x(\U1300/naack ), .a(nba) );
    nor2_1 \U1300/U1130/U5  ( .x(\U1300/nback ), .a(nda), .b(\U1300/reset ) );
    aoai211_1 \U1300/U1128/U28/U1/U1  ( .x(\U1300/U1128/U28/U1/clr ), .a(
        \U1300/r ), .b(\U1300/naack ), .c(dg), .d(dsel) );
    nand3_1 \U1300/U1128/U28/U1/U2  ( .x(\U1300/U1128/U28/U1/set ), .a(dg), 
        .b(\U1300/r ), .c(\U1300/naack ) );
    nand2_2 \U1300/U1128/U28/U1/U3  ( .x(dsel), .a(\U1300/U1128/U28/U1/clr ), 
        .b(\U1300/U1128/U28/U1/set ) );
    aoai211_1 \U1300/U1127/U28/U1/U1  ( .x(\U1300/U1127/U28/U1/clr ), .a(
        \U1300/s ), .b(\U1300/nback ), .c(bg), .d(bsel) );
    nand3_1 \U1300/U1127/U28/U1/U2  ( .x(\U1300/U1127/U28/U1/set ), .a(bg), 
        .b(\U1300/s ), .c(\U1300/nback ) );
    nand2_2 \U1300/U1127/U28/U1/U3  ( .x(bsel), .a(\U1300/U1127/U28/U1/clr ), 
        .b(\U1300/U1127/U28/U1/set ) );
    aoai211_1 \U1289/U1150/U28/U1/U1  ( .x(\U1289/U1150/U28/U1/clr ), .a(il[2]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdl[2] ) );
    nand3_1 \U1289/U1150/U28/U1/U2  ( .x(\U1289/U1150/U28/U1/set ), .a(net195), 
        .b(il[2]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1150/U28/U1/U3  ( .x(\cdl[2] ), .a(
        \U1289/U1150/U28/U1/clr ), .b(\U1289/U1150/U28/U1/set ) );
    aoai211_1 \U1289/U1152/U28/U1/U1  ( .x(\U1289/U1152/U28/U1/clr ), .a(il[3]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdl[3] ) );
    nand3_1 \U1289/U1152/U28/U1/U2  ( .x(\U1289/U1152/U28/U1/set ), .a(net195), 
        .b(il[3]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1152/U28/U1/U3  ( .x(\cdl[3] ), .a(
        \U1289/U1152/U28/U1/clr ), .b(\U1289/U1152/U28/U1/set ) );
    aoai211_1 \U1289/U1149/U28/U1/U1  ( .x(\U1289/U1149/U28/U1/clr ), .a(ih[2]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdh[2] ) );
    nand3_1 \U1289/U1149/U28/U1/U2  ( .x(\U1289/U1149/U28/U1/set ), .a(net195), 
        .b(ih[2]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1149/U28/U1/U3  ( .x(\cdh[2] ), .a(
        \U1289/U1149/U28/U1/clr ), .b(\U1289/U1149/U28/U1/set ) );
    aoai211_1 \U1289/U1151/U28/U1/U1  ( .x(\U1289/U1151/U28/U1/clr ), .a(ih[3]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdh[3] ) );
    nand3_1 \U1289/U1151/U28/U1/U2  ( .x(\U1289/U1151/U28/U1/set ), .a(net195), 
        .b(ih[3]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1151/U28/U1/U3  ( .x(\cdh[3] ), .a(
        \U1289/U1151/U28/U1/clr ), .b(\U1289/U1151/U28/U1/set ) );
    inv_1 \U1289/U1148/U1147/U3  ( .x(\U1289/U1148/net189 ), .a(
        \U1289/bnreset ) );
    nor2_1 \U1289/U1148/U582/U5  ( .x(\U1289/U1148/net192 ), .a(\cdl[3] ), .b(
        \cdh[3] ) );
    nor2_1 \U1289/U1148/U580/U5  ( .x(\U1289/U1148/net191 ), .a(\cdl[2] ), .b(
        \cdh[2] ) );
    nor2_2 \U1289/U1148/U1146/U6  ( .x(\twobitack[2] ), .a(
        \U1289/U1148/net190 ), .b(\U1289/U1148/net189 ) );
    aoi222_1 \U1289/U1148/U1141/U30/U1  ( .x(\U1289/U1148/net190 ), .a(
        \U1289/U1148/net191 ), .b(\U1289/U1148/net192 ), .c(
        \U1289/U1148/net191 ), .d(\U1289/U1148/U1141/Z ), .e(
        \U1289/U1148/net192 ), .f(\U1289/U1148/U1141/Z ) );
    inv_1 \U1289/U1148/U1141/U30/Uinv  ( .x(\U1289/U1148/U1141/Z ), .a(
        \U1289/U1148/net190 ) );
    aoai211_1 \U1271/U1150/U28/U1/U1  ( .x(\U1271/U1150/U28/U1/clr ), .a(il[0]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdl[0] ) );
    nand3_1 \U1271/U1150/U28/U1/U2  ( .x(\U1271/U1150/U28/U1/set ), .a(net193), 
        .b(il[0]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1150/U28/U1/U3  ( .x(\cdl[0] ), .a(
        \U1271/U1150/U28/U1/clr ), .b(\U1271/U1150/U28/U1/set ) );
    aoai211_1 \U1271/U1152/U28/U1/U1  ( .x(\U1271/U1152/U28/U1/clr ), .a(il[1]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdl[1] ) );
    nand3_1 \U1271/U1152/U28/U1/U2  ( .x(\U1271/U1152/U28/U1/set ), .a(net193), 
        .b(il[1]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1152/U28/U1/U3  ( .x(\cdl[1] ), .a(
        \U1271/U1152/U28/U1/clr ), .b(\U1271/U1152/U28/U1/set ) );
    aoai211_1 \U1271/U1149/U28/U1/U1  ( .x(\U1271/U1149/U28/U1/clr ), .a(ih[0]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdh[0] ) );
    nand3_1 \U1271/U1149/U28/U1/U2  ( .x(\U1271/U1149/U28/U1/set ), .a(net193), 
        .b(ih[0]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1149/U28/U1/U3  ( .x(\cdh[0] ), .a(
        \U1271/U1149/U28/U1/clr ), .b(\U1271/U1149/U28/U1/set ) );
    aoai211_1 \U1271/U1151/U28/U1/U1  ( .x(\U1271/U1151/U28/U1/clr ), .a(ih[1]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdh[1] ) );
    nand3_1 \U1271/U1151/U28/U1/U2  ( .x(\U1271/U1151/U28/U1/set ), .a(net193), 
        .b(ih[1]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1151/U28/U1/U3  ( .x(\cdh[1] ), .a(
        \U1271/U1151/U28/U1/clr ), .b(\U1271/U1151/U28/U1/set ) );
    inv_1 \U1271/U1148/U1147/U3  ( .x(\U1271/U1148/net189 ), .a(
        \U1271/bnreset ) );
    nor2_1 \U1271/U1148/U582/U5  ( .x(\U1271/U1148/net192 ), .a(\cdl[1] ), .b(
        \cdh[1] ) );
    nor2_1 \U1271/U1148/U580/U5  ( .x(\U1271/U1148/net191 ), .a(\cdl[0] ), .b(
        \cdh[0] ) );
    nor2_2 \U1271/U1148/U1146/U6  ( .x(\twobitack[0] ), .a(
        \U1271/U1148/net190 ), .b(\U1271/U1148/net189 ) );
    aoi222_1 \U1271/U1148/U1141/U30/U1  ( .x(\U1271/U1148/net190 ), .a(
        \U1271/U1148/net191 ), .b(\U1271/U1148/net192 ), .c(
        \U1271/U1148/net191 ), .d(\U1271/U1148/U1141/Z ), .e(
        \U1271/U1148/net192 ), .f(\U1271/U1148/U1141/Z ) );
    inv_1 \U1271/U1148/U1141/U30/Uinv  ( .x(\U1271/U1148/U1141/Z ), .a(
        \U1271/U1148/net190 ) );
    nand2_1 \U1225/U1128/U5  ( .x(\U1225/s ), .a(\U1225/r ), .b(\U1225/nback )
         );
    nand2_1 \U1225/U1103/U5  ( .x(\U1225/r ), .a(\U1225/naack ), .b(\U1225/s )
         );
    inv_1 \U1225/U1111/U3  ( .x(\U1225/reset ), .a(nbReset) );
    inv_1 \U1225/U1112/U3  ( .x(\U1225/naack ), .a(nxa) );
    nor2_1 \U1225/U1127/U5  ( .x(\U1225/nback ), .a(nyla), .b(\U1225/reset )
         );
    and2_2 \U1225/U1129/U8  ( .x(xsel), .a(\U1225/nback ), .b(\U1225/s ) );
    and2_2 \U1225/U1124/U8  ( .x(ysel), .a(\U1225/r ), .b(\U1225/naack ) );
    and3_4 \U1308/U20/U9  ( .x(nya), .a(\U1308/nack[1] ), .b(\U1308/nack[0] ), 
        .c(nbReset) );
    nor2_1 \U1308/U18/U5  ( .x(\U1308/nack[0] ), .a(\yl[3] ), .b(\yl[0] ) );
    nor2_1 \U1308/U19/U5  ( .x(\U1308/nack[1] ), .a(\yl[1] ), .b(\yl[2] ) );
    ao222_2 \U1308/U15_0_/U19/U1/U1  ( .x(\yl[0] ), .a(\y[0] ), .b(nyla), .c(
        \y[0] ), .d(\yl[0] ), .e(nyla), .f(\yl[0] ) );
    ao222_2 \U1308/U15_1_/U19/U1/U1  ( .x(\yl[1] ), .a(\y[1] ), .b(nyla), .c(
        \y[1] ), .d(\yl[1] ), .e(nyla), .f(\yl[1] ) );
    ao222_2 \U1308/U15_2_/U19/U1/U1  ( .x(\yl[2] ), .a(\y[2] ), .b(nyla), .c(
        \y[2] ), .d(\yl[2] ), .e(nyla), .f(\yl[2] ) );
    ao222_2 \U1308/U15_3_/U19/U1/U1  ( .x(\yl[3] ), .a(\y[3] ), .b(nyla), .c(
        \y[3] ), .d(\yl[3] ), .e(nyla), .f(\yl[3] ) );
    buf_3 U1 ( .x(\U1271/bnreset ), .a(nbReset) );
    buf_3 U2 ( .x(\U1289/bnreset ), .a(nbReset) );
endmodule


module chain_mergepackets_5 ( naa, nba, o, a, b, nReset, noa );
output [4:0] o;
input  [4:0] a;
input  [4:0] b;
input  nReset, noa;
output naa, nba;
    wire as, seta, asel, bsel, setb, reset, \noack[1] , \noack[0] , 
        \U916_0_/U25/U1/clr , \U916_0_/U25/U1/ob , \U916_1_/U25/U1/clr , 
        \U916_1_/U25/U1/ob , \U916_2_/U25/U1/clr , \U916_2_/U25/U1/ob , 
        \U916_3_/U25/U1/clr , \U916_3_/U25/U1/ob ;
    and2_1 \U1155/U8  ( .x(as), .a(seta), .b(asel) );
    nand2_1 \U1145/U5  ( .x(asel), .a(bsel), .b(seta) );
    nand2_1 \U1103/U5  ( .x(bsel), .a(setb), .b(asel) );
    inv_1 \U1135/U3  ( .x(reset), .a(nReset) );
    inv_1 \U1134/U3  ( .x(setb), .a(a[4]) );
    and3_2 \U1154/U9  ( .x(naa), .a(\noack[1] ), .b(\noack[0] ), .c(as) );
    nor3_1 \U1127/U7  ( .x(\noack[0] ), .a(o[1]), .b(reset), .c(o[0]) );
    nor2_1 \U1132/U5  ( .x(\noack[1] ), .a(o[3]), .b(o[2]) );
    oa31_1 \U916_0_/U25/U1/Uclr  ( .x(\U916_0_/U25/U1/clr ), .a(noa), .b(a[0]), 
        .c(b[0]), .d(o[0]) );
    oaoi211_1 \U916_0_/U25/U1/Uaoi  ( .x(\U916_0_/U25/U1/ob ), .a(a[0]), .b(b
        [0]), .c(noa), .d(\U916_0_/U25/U1/clr ) );
    inv_2 \U916_0_/U25/U1/Ui  ( .x(o[0]), .a(\U916_0_/U25/U1/ob ) );
    oa31_1 \U916_1_/U25/U1/Uclr  ( .x(\U916_1_/U25/U1/clr ), .a(noa), .b(a[1]), 
        .c(b[1]), .d(o[1]) );
    oaoi211_1 \U916_1_/U25/U1/Uaoi  ( .x(\U916_1_/U25/U1/ob ), .a(a[1]), .b(b
        [1]), .c(noa), .d(\U916_1_/U25/U1/clr ) );
    inv_2 \U916_1_/U25/U1/Ui  ( .x(o[1]), .a(\U916_1_/U25/U1/ob ) );
    oa31_1 \U916_2_/U25/U1/Uclr  ( .x(\U916_2_/U25/U1/clr ), .a(noa), .b(a[2]), 
        .c(b[2]), .d(o[2]) );
    oaoi211_1 \U916_2_/U25/U1/Uaoi  ( .x(\U916_2_/U25/U1/ob ), .a(a[2]), .b(b
        [2]), .c(noa), .d(\U916_2_/U25/U1/clr ) );
    inv_2 \U916_2_/U25/U1/Ui  ( .x(o[2]), .a(\U916_2_/U25/U1/ob ) );
    oa31_1 \U916_3_/U25/U1/Uclr  ( .x(\U916_3_/U25/U1/clr ), .a(noa), .b(a[3]), 
        .c(b[3]), .d(o[3]) );
    oaoi211_1 \U916_3_/U25/U1/Uaoi  ( .x(\U916_3_/U25/U1/ob ), .a(a[3]), .b(b
        [3]), .c(noa), .d(\U916_3_/U25/U1/clr ) );
    inv_2 \U916_3_/U25/U1/Ui  ( .x(o[3]), .a(\U916_3_/U25/U1/ob ) );
    ao222_2 \U1148/U19/U1/U1  ( .x(o[4]), .a(noa), .b(b[4]), .c(noa), .d(o[4]), 
        .e(b[4]), .f(o[4]) );
    aoi21_1 \U1153/U11  ( .x(seta), .a(o[4]), .b(setb), .c(reset) );
    and3_3 U1 ( .x(nba), .a(bsel), .b(\noack[0] ), .c(\noack[1] ) );
endmodule


module chain_tchdr_2 ( addr_req, col_h, col_l, itag_h, itag_l, lock, ncback, 
    neop, pred, pullcd, reset, rnw_h, rnw_l, seq, size_h, size_l, write_req, 
    chwh, chwl, addr_ack, addr_pull, nReset, nack, write_ack, write_pull );
output [2:0] col_h;
output [2:0] col_l;
output [4:0] itag_h;
output [4:0] itag_l;
output [1:0] lock;
output [1:0] pred;
output [1:0] seq;
output [1:0] size_h;
output [1:0] size_l;
input  [7:0] chwh;
input  [7:0] chwl;
input  addr_ack, addr_pull, nReset, nack, write_ack, write_pull;
output addr_req, ncback, neop, pullcd, reset, rnw_h, rnw_l, write_req;
    wire n9, pullcdwk, net94, net88, \ncd[0] , \ncd[1] , \ncd[2] , \ncd[3] , 
        \ncd[4] , \ncd[5] , \ncd[6] , \ncd[7] , read, ack, net83, \U1664/x[3] , 
        \U1664/U28/Z , \U1664/x[0] , \U1664/U32/Z , \U1664/x[2] , 
        \U1664/U29/Z , \U1664/y[0] , \U1664/x[1] , \U1664/U33/Z , \U1664/y[1] , 
        \U1664/U30/Z , \U1664/U31/Z , \U1664/U37/Z , receive, \U473/Z , 
        \hdr_hld/net32 , \hdr_hld/net33 , \hdr_hld/low/latch , 
        \hdr_hld/low/nlocalcd , \hdr_hld/low/localcd , \hdr_hld/low/ncd[0] , 
        \hdr_hld/low/ncd[1] , \hdr_hld/low/ncd[2] , \hdr_hld/low/ncd[3] , 
        \hdr_hld/ol[3] , \hdr_hld/oh[3] , \hdr_hld/low/ncd[4] , 
        \hdr_hld/ol[4] , \hdr_hld/oh[4] , \hdr_hld/low/ncd[5] , 
        \hdr_hld/low/ncd[6] , \hdr_hld/low/ncd[7] , 
        \hdr_hld/low/ctrlack_internal , \hdr_hld/low/acb , \hdr_hld/low/ba , 
        \hdr_hld/low/driveh , \hdr_hld/net20 , \hdr_hld/low/drivel , n2, n3, 
        n1, \hdr_hld/low/U4/U28/U1/clr , \hdr_hld/low/U4/U28/U1/set , 
        \hdr_hld/low/U1/Z , \hdr_hld/low/U1664/x[3] , 
        \hdr_hld/low/U1664/U28/Z , \hdr_hld/low/U1664/x[0] , 
        \hdr_hld/low/U1664/U32/Z , \hdr_hld/low/U1664/x[2] , 
        \hdr_hld/low/U1664/U29/Z , \hdr_hld/low/U1664/y[0] , 
        \hdr_hld/low/U1664/x[1] , \hdr_hld/low/U1664/U33/Z , 
        \hdr_hld/low/U1664/y[1] , \hdr_hld/low/U1664/U30/Z , 
        \hdr_hld/low/U1664/U31/Z , \hdr_hld/low/U1664/U37/Z , 
        \hdr_hld/low/U1669/nr , \hdr_hld/low/U1669/nd , \hdr_hld/low/U1669/n2 , 
        \hdr_hld/high/latch , \hdr_hld/high/nlocalcd , \hdr_hld/high/localcd , 
        \hdr_hld/high/ncd[0] , \hdr_hld/high/ncd[1] , \hdr_hld/high/ncd[2] , 
        \hdr_hld/high/ncd[3] , \hdr_hld/high/ncd[4] , \hdr_hld/high/ncd[5] , 
        \hdr_hld/high/ncd[6] , \hdr_hld/high/ncd[7] , 
        \hdr_hld/high/ctrlack_internal , \hdr_hld/high/acb , \hdr_hld/high/ba , 
        \hdr_hld/high/driveh , \hdr_hld/high/drivel , n7, n4, n5, n6, 
        \hdr_hld/high/U4/U28/U1/clr , \hdr_hld/high/U4/U28/U1/set , 
        \hdr_hld/high/U1/Z , \hdr_hld/high/U1664/x[3] , 
        \hdr_hld/high/U1664/U28/Z , \hdr_hld/high/U1664/x[0] , 
        \hdr_hld/high/U1664/U32/Z , \hdr_hld/high/U1664/x[2] , 
        \hdr_hld/high/U1664/U29/Z , \hdr_hld/high/U1664/y[0] , 
        \hdr_hld/high/U1664/x[1] , \hdr_hld/high/U1664/U33/Z , 
        \hdr_hld/high/U1664/y[1] , \hdr_hld/high/U1664/U30/Z , 
        \hdr_hld/high/U1664/U31/Z , \hdr_hld/high/U1664/U37/Z , 
        \hdr_hld/high/U1669/nr , \hdr_hld/high/U1669/nd , 
        \hdr_hld/high/U1669/n2 ;
    buf_1 U262 ( .x(n9), .a(pullcdwk) );
    or3_2 \U1668/U12  ( .x(ncback), .a(net94), .b(addr_pull), .c(write_pull)
         );
    inv_1 \I0/U3  ( .x(net94), .a(net88) );
    nor2_1 \U514_0_/U5  ( .x(\ncd[0] ), .a(chwh[0]), .b(chwl[0]) );
    nor2_1 \U514_1_/U5  ( .x(\ncd[1] ), .a(chwh[1]), .b(chwl[1]) );
    nor2_1 \U514_2_/U5  ( .x(\ncd[2] ), .a(chwh[2]), .b(chwl[2]) );
    nor2_1 \U514_3_/U5  ( .x(\ncd[3] ), .a(chwh[3]), .b(chwl[3]) );
    nor2_1 \U514_4_/U5  ( .x(\ncd[4] ), .a(chwh[4]), .b(chwl[4]) );
    nor2_1 \U514_5_/U5  ( .x(\ncd[5] ), .a(chwh[5]), .b(chwl[5]) );
    nor2_1 \U514_6_/U5  ( .x(\ncd[6] ), .a(chwh[6]), .b(chwl[6]) );
    nor2_1 \U514_7_/U5  ( .x(\ncd[7] ), .a(chwh[7]), .b(chwl[7]) );
    nor2_1 \U1669/U5  ( .x(neop), .a(read), .b(write_ack) );
    nand2_1 \U303/U5  ( .x(ack), .a(nack), .b(nReset) );
    nand2_1 \U1670/U5  ( .x(net83), .a(neop), .b(nReset) );
    ao222_1 \U47/U18/U1/U1  ( .x(read), .a(addr_ack), .b(rnw_h), .c(addr_ack), 
        .d(read), .e(rnw_h), .f(read) );
    ao222_1 \U48/U18/U1/U1  ( .x(write_req), .a(rnw_l), .b(addr_ack), .c(rnw_l
        ), .d(write_req), .e(addr_ack), .f(write_req) );
    aoi222_1 \U1664/U28/U30/U1  ( .x(\U1664/x[3] ), .a(\ncd[7] ), .b(\ncd[6] ), 
        .c(\ncd[7] ), .d(\U1664/U28/Z ), .e(\ncd[6] ), .f(\U1664/U28/Z ) );
    inv_1 \U1664/U28/U30/Uinv  ( .x(\U1664/U28/Z ), .a(\U1664/x[3] ) );
    aoi222_1 \U1664/U32/U30/U1  ( .x(\U1664/x[0] ), .a(\ncd[1] ), .b(\ncd[0] ), 
        .c(\ncd[1] ), .d(\U1664/U32/Z ), .e(\ncd[0] ), .f(\U1664/U32/Z ) );
    inv_1 \U1664/U32/U30/Uinv  ( .x(\U1664/U32/Z ), .a(\U1664/x[0] ) );
    aoi222_1 \U1664/U29/U30/U1  ( .x(\U1664/x[2] ), .a(\ncd[5] ), .b(\ncd[4] ), 
        .c(\ncd[5] ), .d(\U1664/U29/Z ), .e(\ncd[4] ), .f(\U1664/U29/Z ) );
    inv_1 \U1664/U29/U30/Uinv  ( .x(\U1664/U29/Z ), .a(\U1664/x[2] ) );
    aoi222_1 \U1664/U33/U30/U1  ( .x(\U1664/y[0] ), .a(\U1664/x[1] ), .b(
        \U1664/x[0] ), .c(\U1664/x[1] ), .d(\U1664/U33/Z ), .e(\U1664/x[0] ), 
        .f(\U1664/U33/Z ) );
    inv_1 \U1664/U33/U30/Uinv  ( .x(\U1664/U33/Z ), .a(\U1664/y[0] ) );
    aoi222_1 \U1664/U30/U30/U1  ( .x(\U1664/y[1] ), .a(\U1664/x[3] ), .b(
        \U1664/x[2] ), .c(\U1664/x[3] ), .d(\U1664/U30/Z ), .e(\U1664/x[2] ), 
        .f(\U1664/U30/Z ) );
    inv_1 \U1664/U30/U30/Uinv  ( .x(\U1664/U30/Z ), .a(\U1664/y[1] ) );
    aoi222_1 \U1664/U31/U30/U1  ( .x(\U1664/x[1] ), .a(\ncd[3] ), .b(\ncd[2] ), 
        .c(\ncd[3] ), .d(\U1664/U31/Z ), .e(\ncd[2] ), .f(\U1664/U31/Z ) );
    inv_1 \U1664/U31/U30/Uinv  ( .x(\U1664/U31/Z ), .a(\U1664/x[1] ) );
    aoi222_1 \U1664/U37/U30/U1  ( .x(pullcdwk), .a(\U1664/y[0] ), .b(
        \U1664/y[1] ), .c(\U1664/y[0] ), .d(\U1664/U37/Z ), .e(\U1664/y[1] ), 
        .f(\U1664/U37/Z ) );
    inv_1 \U1664/U37/U30/Uinv  ( .x(\U1664/U37/Z ), .a(pullcdwk) );
    aoi222_1 \U473/U30/U1  ( .x(receive), .a(net83), .b(ack), .c(net83), .d(
        \U473/Z ), .e(ack), .f(\U473/Z ) );
    inv_1 \U473/U30/Uinv  ( .x(\U473/Z ), .a(receive) );
    nor2_1 \hdr_hld/U3/U5  ( .x(net88), .a(\hdr_hld/net32 ), .b(
        \hdr_hld/net33 ) );
    buf_2 \hdr_hld/low/U1653  ( .x(\hdr_hld/low/latch ), .a(\hdr_hld/net32 )
         );
    nor2_1 \hdr_hld/low/U264/U5  ( .x(\hdr_hld/low/nlocalcd ), .a(reset), .b(
        \hdr_hld/low/localcd ) );
    nor2_1 \hdr_hld/low/U1659_0_/U5  ( .x(\hdr_hld/low/ncd[0] ), .a(seq[0]), 
        .b(seq[1]) );
    nor2_1 \hdr_hld/low/U1659_1_/U5  ( .x(\hdr_hld/low/ncd[1] ), .a(pred[0]), 
        .b(pred[1]) );
    nor2_1 \hdr_hld/low/U1659_2_/U5  ( .x(\hdr_hld/low/ncd[2] ), .a(lock[0]), 
        .b(lock[1]) );
    nor2_1 \hdr_hld/low/U1659_3_/U5  ( .x(\hdr_hld/low/ncd[3] ), .a(
        \hdr_hld/ol[3] ), .b(\hdr_hld/oh[3] ) );
    nor2_1 \hdr_hld/low/U1659_4_/U5  ( .x(\hdr_hld/low/ncd[4] ), .a(
        \hdr_hld/ol[4] ), .b(\hdr_hld/oh[4] ) );
    nor2_1 \hdr_hld/low/U1659_5_/U5  ( .x(\hdr_hld/low/ncd[5] ), .a(rnw_l), 
        .b(rnw_h) );
    nor2_1 \hdr_hld/low/U1659_6_/U5  ( .x(\hdr_hld/low/ncd[6] ), .a(size_l[0]), 
        .b(size_h[0]) );
    nor2_1 \hdr_hld/low/U1659_7_/U5  ( .x(\hdr_hld/low/ncd[7] ), .a(size_l[1]), 
        .b(size_h[1]) );
    nor2_1 \hdr_hld/low/U3/U5  ( .x(\hdr_hld/low/ctrlack_internal ), .a(
        \hdr_hld/low/acb ), .b(\hdr_hld/low/ba ) );
    buf_2 \hdr_hld/low/U1665/U7  ( .x(\hdr_hld/low/driveh ), .a(
        \hdr_hld/net20 ) );
    buf_2 \hdr_hld/low/U1666/U7  ( .x(\hdr_hld/low/drivel ), .a(
        \hdr_hld/net20 ) );
    ao23_1 \hdr_hld/low/U1658_0_/U21/U1/U1  ( .x(seq[0]), .a(n2), .b(seq[0]), 
        .c(\hdr_hld/low/drivel ), .d(chwl[0]), .e(n3) );
    ao23_1 \hdr_hld/low/U1658_1_/U21/U1/U1  ( .x(pred[0]), .a(n1), .b(pred[0]), 
        .c(\hdr_hld/low/drivel ), .d(chwl[1]), .e(n3) );
    ao23_1 \hdr_hld/low/U1658_2_/U21/U1/U1  ( .x(lock[0]), .a(n1), .b(lock[0]), 
        .c(\hdr_hld/low/driveh ), .d(chwl[2]), .e(n3) );
    ao23_1 \hdr_hld/low/U1658_3_/U21/U1/U1  ( .x(\hdr_hld/ol[3] ), .a(n1), .b(
        \hdr_hld/ol[3] ), .c(\hdr_hld/low/driveh ), .d(chwl[3]), .e(
        \hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1658_4_/U21/U1/U1  ( .x(\hdr_hld/ol[4] ), .a(n2), .b(
        \hdr_hld/ol[4] ), .c(\hdr_hld/low/drivel ), .d(chwl[4]), .e(
        \hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1658_5_/U21/U1/U1  ( .x(rnw_l), .a(
        \hdr_hld/low/driveh ), .b(rnw_l), .c(\hdr_hld/low/driveh ), .d(chwl[5]
        ), .e(\hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1658_6_/U21/U1/U1  ( .x(size_l[0]), .a(
        \hdr_hld/low/drivel ), .b(size_l[0]), .c(n2), .d(chwl[6]), .e(
        \hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1658_7_/U21/U1/U1  ( .x(size_l[1]), .a(
        \hdr_hld/low/drivel ), .b(size_l[1]), .c(\hdr_hld/low/drivel ), .d(
        chwl[7]), .e(\hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1651_0_/U21/U1/U1  ( .x(seq[1]), .a(
        \hdr_hld/low/drivel ), .b(seq[1]), .c(\hdr_hld/low/driveh ), .d(chwh
        [0]), .e(\hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1651_1_/U21/U1/U1  ( .x(pred[1]), .a(
        \hdr_hld/low/driveh ), .b(pred[1]), .c(n1), .d(chwh[1]), .e(
        \hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1651_2_/U21/U1/U1  ( .x(lock[1]), .a(
        \hdr_hld/low/driveh ), .b(lock[1]), .c(n1), .d(chwh[2]), .e(
        \hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1651_3_/U21/U1/U1  ( .x(\hdr_hld/oh[3] ), .a(
        \hdr_hld/low/drivel ), .b(\hdr_hld/oh[3] ), .c(n2), .d(chwh[3]), .e(
        \hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1651_4_/U21/U1/U1  ( .x(\hdr_hld/oh[4] ), .a(n2), .b(
        \hdr_hld/oh[4] ), .c(n1), .d(chwh[4]), .e(\hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1651_5_/U21/U1/U1  ( .x(rnw_h), .a(n2), .b(rnw_h), 
        .c(n1), .d(chwh[5]), .e(\hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1651_6_/U21/U1/U1  ( .x(size_h[0]), .a(n1), .b(size_h
        [0]), .c(n2), .d(chwh[6]), .e(\hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1651_7_/U21/U1/U1  ( .x(size_h[1]), .a(
        \hdr_hld/low/driveh ), .b(size_h[1]), .c(n2), .d(chwh[7]), .e(
        \hdr_hld/low/latch ) );
    aoai211_1 \hdr_hld/low/U4/U28/U1/U1  ( .x(\hdr_hld/low/U4/U28/U1/clr ), 
        .a(\hdr_hld/net20 ), .b(\hdr_hld/low/acb ), .c(\hdr_hld/low/nlocalcd ), 
        .d(\hdr_hld/net32 ) );
    nand3_1 \hdr_hld/low/U4/U28/U1/U2  ( .x(\hdr_hld/low/U4/U28/U1/set ), .a(
        \hdr_hld/low/nlocalcd ), .b(\hdr_hld/net20 ), .c(\hdr_hld/low/acb ) );
    nand2_2 \hdr_hld/low/U4/U28/U1/U3  ( .x(\hdr_hld/net32 ), .a(
        \hdr_hld/low/U4/U28/U1/clr ), .b(\hdr_hld/low/U4/U28/U1/set ) );
    oai21_1 \hdr_hld/low/U1/U30/U1/U1  ( .x(\hdr_hld/low/acb ), .a(
        \hdr_hld/low/U1/Z ), .b(\hdr_hld/low/ba ), .c(\hdr_hld/net20 ) );
    inv_1 \hdr_hld/low/U1/U30/U1/U2  ( .x(\hdr_hld/low/U1/Z ), .a(
        \hdr_hld/low/acb ) );
    ao222_1 \hdr_hld/low/U5/U18/U1/U1  ( .x(\hdr_hld/low/ba ), .a(
        \hdr_hld/low/latch ), .b(n9), .c(\hdr_hld/low/latch ), .d(
        \hdr_hld/low/ba ), .e(n9), .f(\hdr_hld/low/ba ) );
    aoi222_1 \hdr_hld/low/U1664/U28/U30/U1  ( .x(\hdr_hld/low/U1664/x[3] ), 
        .a(\hdr_hld/low/ncd[7] ), .b(\hdr_hld/low/ncd[6] ), .c(
        \hdr_hld/low/ncd[7] ), .d(\hdr_hld/low/U1664/U28/Z ), .e(
        \hdr_hld/low/ncd[6] ), .f(\hdr_hld/low/U1664/U28/Z ) );
    inv_1 \hdr_hld/low/U1664/U28/U30/Uinv  ( .x(\hdr_hld/low/U1664/U28/Z ), 
        .a(\hdr_hld/low/U1664/x[3] ) );
    aoi222_1 \hdr_hld/low/U1664/U32/U30/U1  ( .x(\hdr_hld/low/U1664/x[0] ), 
        .a(\hdr_hld/low/ncd[1] ), .b(\hdr_hld/low/ncd[0] ), .c(
        \hdr_hld/low/ncd[1] ), .d(\hdr_hld/low/U1664/U32/Z ), .e(
        \hdr_hld/low/ncd[0] ), .f(\hdr_hld/low/U1664/U32/Z ) );
    inv_1 \hdr_hld/low/U1664/U32/U30/Uinv  ( .x(\hdr_hld/low/U1664/U32/Z ), 
        .a(\hdr_hld/low/U1664/x[0] ) );
    aoi222_1 \hdr_hld/low/U1664/U29/U30/U1  ( .x(\hdr_hld/low/U1664/x[2] ), 
        .a(\hdr_hld/low/ncd[5] ), .b(\hdr_hld/low/ncd[4] ), .c(
        \hdr_hld/low/ncd[5] ), .d(\hdr_hld/low/U1664/U29/Z ), .e(
        \hdr_hld/low/ncd[4] ), .f(\hdr_hld/low/U1664/U29/Z ) );
    inv_1 \hdr_hld/low/U1664/U29/U30/Uinv  ( .x(\hdr_hld/low/U1664/U29/Z ), 
        .a(\hdr_hld/low/U1664/x[2] ) );
    aoi222_1 \hdr_hld/low/U1664/U33/U30/U1  ( .x(\hdr_hld/low/U1664/y[0] ), 
        .a(\hdr_hld/low/U1664/x[1] ), .b(\hdr_hld/low/U1664/x[0] ), .c(
        \hdr_hld/low/U1664/x[1] ), .d(\hdr_hld/low/U1664/U33/Z ), .e(
        \hdr_hld/low/U1664/x[0] ), .f(\hdr_hld/low/U1664/U33/Z ) );
    inv_1 \hdr_hld/low/U1664/U33/U30/Uinv  ( .x(\hdr_hld/low/U1664/U33/Z ), 
        .a(\hdr_hld/low/U1664/y[0] ) );
    aoi222_1 \hdr_hld/low/U1664/U30/U30/U1  ( .x(\hdr_hld/low/U1664/y[1] ), 
        .a(\hdr_hld/low/U1664/x[3] ), .b(\hdr_hld/low/U1664/x[2] ), .c(
        \hdr_hld/low/U1664/x[3] ), .d(\hdr_hld/low/U1664/U30/Z ), .e(
        \hdr_hld/low/U1664/x[2] ), .f(\hdr_hld/low/U1664/U30/Z ) );
    inv_1 \hdr_hld/low/U1664/U30/U30/Uinv  ( .x(\hdr_hld/low/U1664/U30/Z ), 
        .a(\hdr_hld/low/U1664/y[1] ) );
    aoi222_1 \hdr_hld/low/U1664/U31/U30/U1  ( .x(\hdr_hld/low/U1664/x[1] ), 
        .a(\hdr_hld/low/ncd[3] ), .b(\hdr_hld/low/ncd[2] ), .c(
        \hdr_hld/low/ncd[3] ), .d(\hdr_hld/low/U1664/U31/Z ), .e(
        \hdr_hld/low/ncd[2] ), .f(\hdr_hld/low/U1664/U31/Z ) );
    inv_1 \hdr_hld/low/U1664/U31/U30/Uinv  ( .x(\hdr_hld/low/U1664/U31/Z ), 
        .a(\hdr_hld/low/U1664/x[1] ) );
    aoi222_1 \hdr_hld/low/U1664/U37/U30/U1  ( .x(\hdr_hld/low/localcd ), .a(
        \hdr_hld/low/U1664/y[0] ), .b(\hdr_hld/low/U1664/y[1] ), .c(
        \hdr_hld/low/U1664/y[0] ), .d(\hdr_hld/low/U1664/U37/Z ), .e(
        \hdr_hld/low/U1664/y[1] ), .f(\hdr_hld/low/U1664/U37/Z ) );
    inv_1 \hdr_hld/low/U1664/U37/U30/Uinv  ( .x(\hdr_hld/low/U1664/U37/Z ), 
        .a(\hdr_hld/low/localcd ) );
    nor3_1 \hdr_hld/low/U1669/Unr  ( .x(\hdr_hld/low/U1669/nr ), .a(
        \hdr_hld/low/ctrlack_internal ), .b(\hdr_hld/low/driveh ), .c(n1) );
    nand3_1 \hdr_hld/low/U1669/Und  ( .x(\hdr_hld/low/U1669/nd ), .a(
        \hdr_hld/low/ctrlack_internal ), .b(n2), .c(\hdr_hld/low/drivel ) );
    oa21_1 \hdr_hld/low/U1669/U1  ( .x(\hdr_hld/low/U1669/n2 ), .a(
        \hdr_hld/low/U1669/n2 ), .b(\hdr_hld/low/U1669/nr ), .c(
        \hdr_hld/low/U1669/nd ) );
    inv_2 \hdr_hld/low/U1669/U3  ( .x(addr_req), .a(\hdr_hld/low/U1669/n2 ) );
    buf_2 \hdr_hld/high/U1653  ( .x(\hdr_hld/high/latch ), .a(\hdr_hld/net33 )
         );
    nor2_1 \hdr_hld/high/U264/U5  ( .x(\hdr_hld/high/nlocalcd ), .a(reset), 
        .b(\hdr_hld/high/localcd ) );
    nor2_1 \hdr_hld/high/U1659_0_/U5  ( .x(\hdr_hld/high/ncd[0] ), .a(itag_l
        [0]), .b(itag_h[0]) );
    nor2_1 \hdr_hld/high/U1659_1_/U5  ( .x(\hdr_hld/high/ncd[1] ), .a(itag_l
        [1]), .b(itag_h[1]) );
    nor2_1 \hdr_hld/high/U1659_2_/U5  ( .x(\hdr_hld/high/ncd[2] ), .a(itag_l
        [2]), .b(itag_h[2]) );
    nor2_1 \hdr_hld/high/U1659_3_/U5  ( .x(\hdr_hld/high/ncd[3] ), .a(itag_l
        [3]), .b(itag_h[3]) );
    nor2_1 \hdr_hld/high/U1659_4_/U5  ( .x(\hdr_hld/high/ncd[4] ), .a(itag_l
        [4]), .b(itag_h[4]) );
    nor2_1 \hdr_hld/high/U1659_5_/U5  ( .x(\hdr_hld/high/ncd[5] ), .a(col_l[0]
        ), .b(col_h[0]) );
    nor2_1 \hdr_hld/high/U1659_6_/U5  ( .x(\hdr_hld/high/ncd[6] ), .a(col_l[1]
        ), .b(col_h[1]) );
    nor2_1 \hdr_hld/high/U1659_7_/U5  ( .x(\hdr_hld/high/ncd[7] ), .a(col_l[2]
        ), .b(col_h[2]) );
    nor2_1 \hdr_hld/high/U3/U5  ( .x(\hdr_hld/high/ctrlack_internal ), .a(
        \hdr_hld/high/acb ), .b(\hdr_hld/high/ba ) );
    buf_2 \hdr_hld/high/U1665/U7  ( .x(\hdr_hld/high/driveh ), .a(receive) );
    buf_2 \hdr_hld/high/U1666/U7  ( .x(\hdr_hld/high/drivel ), .a(receive) );
    ao23_1 \hdr_hld/high/U1658_0_/U21/U1/U1  ( .x(itag_l[0]), .a(
        \hdr_hld/high/drivel ), .b(itag_l[0]), .c(\hdr_hld/high/drivel ), .d(
        chwl[0]), .e(n7) );
    ao23_1 \hdr_hld/high/U1658_1_/U21/U1/U1  ( .x(itag_l[1]), .a(
        \hdr_hld/high/drivel ), .b(itag_l[1]), .c(\hdr_hld/high/drivel ), .d(
        chwl[1]), .e(n7) );
    ao23_1 \hdr_hld/high/U1658_2_/U21/U1/U1  ( .x(itag_l[2]), .a(
        \hdr_hld/high/drivel ), .b(itag_l[2]), .c(\hdr_hld/high/drivel ), .d(
        chwl[2]), .e(n7) );
    ao23_1 \hdr_hld/high/U1658_3_/U21/U1/U1  ( .x(itag_l[3]), .a(
        \hdr_hld/high/drivel ), .b(itag_l[3]), .c(\hdr_hld/high/drivel ), .d(
        chwl[3]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1658_4_/U21/U1/U1  ( .x(itag_l[4]), .a(n4), .b(
        itag_l[4]), .c(\hdr_hld/high/drivel ), .d(chwl[4]), .e(
        \hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1658_5_/U21/U1/U1  ( .x(col_l[0]), .a(n4), .b(col_l
        [0]), .c(\hdr_hld/high/drivel ), .d(chwl[5]), .e(\hdr_hld/high/latch )
         );
    ao23_1 \hdr_hld/high/U1658_6_/U21/U1/U1  ( .x(col_l[1]), .a(
        \hdr_hld/high/drivel ), .b(col_l[1]), .c(\hdr_hld/high/drivel ), .d(
        chwl[6]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1658_7_/U21/U1/U1  ( .x(col_l[2]), .a(n4), .b(col_l
        [2]), .c(\hdr_hld/high/drivel ), .d(chwl[7]), .e(\hdr_hld/high/latch )
         );
    ao23_1 \hdr_hld/high/U1651_0_/U21/U1/U1  ( .x(itag_h[0]), .a(n5), .b(
        itag_h[0]), .c(n5), .d(chwh[0]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1651_1_/U21/U1/U1  ( .x(itag_h[1]), .a(n5), .b(
        itag_h[1]), .c(n6), .d(chwh[1]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1651_2_/U21/U1/U1  ( .x(itag_h[2]), .a(n5), .b(
        itag_h[2]), .c(n6), .d(chwh[2]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1651_3_/U21/U1/U1  ( .x(itag_h[3]), .a(n5), .b(
        itag_h[3]), .c(n6), .d(chwh[3]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1651_4_/U21/U1/U1  ( .x(itag_h[4]), .a(n5), .b(
        itag_h[4]), .c(n6), .d(chwh[4]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1651_5_/U21/U1/U1  ( .x(col_h[0]), .a(n5), .b(col_h
        [0]), .c(n6), .d(chwh[5]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1651_6_/U21/U1/U1  ( .x(col_h[1]), .a(n5), .b(col_h
        [1]), .c(n5), .d(chwh[6]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1651_7_/U21/U1/U1  ( .x(col_h[2]), .a(n5), .b(col_h
        [2]), .c(n5), .d(chwh[7]), .e(\hdr_hld/high/latch ) );
    aoai211_1 \hdr_hld/high/U4/U28/U1/U1  ( .x(\hdr_hld/high/U4/U28/U1/clr ), 
        .a(receive), .b(\hdr_hld/high/acb ), .c(\hdr_hld/high/nlocalcd ), .d(
        \hdr_hld/net33 ) );
    nand3_1 \hdr_hld/high/U4/U28/U1/U2  ( .x(\hdr_hld/high/U4/U28/U1/set ), 
        .a(\hdr_hld/high/nlocalcd ), .b(receive), .c(\hdr_hld/high/acb ) );
    nand2_2 \hdr_hld/high/U4/U28/U1/U3  ( .x(\hdr_hld/net33 ), .a(
        \hdr_hld/high/U4/U28/U1/clr ), .b(\hdr_hld/high/U4/U28/U1/set ) );
    oai21_1 \hdr_hld/high/U1/U30/U1/U1  ( .x(\hdr_hld/high/acb ), .a(
        \hdr_hld/high/U1/Z ), .b(\hdr_hld/high/ba ), .c(receive) );
    inv_1 \hdr_hld/high/U1/U30/U1/U2  ( .x(\hdr_hld/high/U1/Z ), .a(
        \hdr_hld/high/acb ) );
    ao222_1 \hdr_hld/high/U5/U18/U1/U1  ( .x(\hdr_hld/high/ba ), .a(
        \hdr_hld/high/latch ), .b(n9), .c(\hdr_hld/high/latch ), .d(
        \hdr_hld/high/ba ), .e(n9), .f(\hdr_hld/high/ba ) );
    aoi222_1 \hdr_hld/high/U1664/U28/U30/U1  ( .x(\hdr_hld/high/U1664/x[3] ), 
        .a(\hdr_hld/high/ncd[7] ), .b(\hdr_hld/high/ncd[6] ), .c(
        \hdr_hld/high/ncd[7] ), .d(\hdr_hld/high/U1664/U28/Z ), .e(
        \hdr_hld/high/ncd[6] ), .f(\hdr_hld/high/U1664/U28/Z ) );
    inv_1 \hdr_hld/high/U1664/U28/U30/Uinv  ( .x(\hdr_hld/high/U1664/U28/Z ), 
        .a(\hdr_hld/high/U1664/x[3] ) );
    aoi222_1 \hdr_hld/high/U1664/U32/U30/U1  ( .x(\hdr_hld/high/U1664/x[0] ), 
        .a(\hdr_hld/high/ncd[1] ), .b(\hdr_hld/high/ncd[0] ), .c(
        \hdr_hld/high/ncd[1] ), .d(\hdr_hld/high/U1664/U32/Z ), .e(
        \hdr_hld/high/ncd[0] ), .f(\hdr_hld/high/U1664/U32/Z ) );
    inv_1 \hdr_hld/high/U1664/U32/U30/Uinv  ( .x(\hdr_hld/high/U1664/U32/Z ), 
        .a(\hdr_hld/high/U1664/x[0] ) );
    aoi222_1 \hdr_hld/high/U1664/U29/U30/U1  ( .x(\hdr_hld/high/U1664/x[2] ), 
        .a(\hdr_hld/high/ncd[5] ), .b(\hdr_hld/high/ncd[4] ), .c(
        \hdr_hld/high/ncd[5] ), .d(\hdr_hld/high/U1664/U29/Z ), .e(
        \hdr_hld/high/ncd[4] ), .f(\hdr_hld/high/U1664/U29/Z ) );
    inv_1 \hdr_hld/high/U1664/U29/U30/Uinv  ( .x(\hdr_hld/high/U1664/U29/Z ), 
        .a(\hdr_hld/high/U1664/x[2] ) );
    aoi222_1 \hdr_hld/high/U1664/U33/U30/U1  ( .x(\hdr_hld/high/U1664/y[0] ), 
        .a(\hdr_hld/high/U1664/x[1] ), .b(\hdr_hld/high/U1664/x[0] ), .c(
        \hdr_hld/high/U1664/x[1] ), .d(\hdr_hld/high/U1664/U33/Z ), .e(
        \hdr_hld/high/U1664/x[0] ), .f(\hdr_hld/high/U1664/U33/Z ) );
    inv_1 \hdr_hld/high/U1664/U33/U30/Uinv  ( .x(\hdr_hld/high/U1664/U33/Z ), 
        .a(\hdr_hld/high/U1664/y[0] ) );
    aoi222_1 \hdr_hld/high/U1664/U30/U30/U1  ( .x(\hdr_hld/high/U1664/y[1] ), 
        .a(\hdr_hld/high/U1664/x[3] ), .b(\hdr_hld/high/U1664/x[2] ), .c(
        \hdr_hld/high/U1664/x[3] ), .d(\hdr_hld/high/U1664/U30/Z ), .e(
        \hdr_hld/high/U1664/x[2] ), .f(\hdr_hld/high/U1664/U30/Z ) );
    inv_1 \hdr_hld/high/U1664/U30/U30/Uinv  ( .x(\hdr_hld/high/U1664/U30/Z ), 
        .a(\hdr_hld/high/U1664/y[1] ) );
    aoi222_1 \hdr_hld/high/U1664/U31/U30/U1  ( .x(\hdr_hld/high/U1664/x[1] ), 
        .a(\hdr_hld/high/ncd[3] ), .b(\hdr_hld/high/ncd[2] ), .c(
        \hdr_hld/high/ncd[3] ), .d(\hdr_hld/high/U1664/U31/Z ), .e(
        \hdr_hld/high/ncd[2] ), .f(\hdr_hld/high/U1664/U31/Z ) );
    inv_1 \hdr_hld/high/U1664/U31/U30/Uinv  ( .x(\hdr_hld/high/U1664/U31/Z ), 
        .a(\hdr_hld/high/U1664/x[1] ) );
    aoi222_1 \hdr_hld/high/U1664/U37/U30/U1  ( .x(\hdr_hld/high/localcd ), .a(
        \hdr_hld/high/U1664/y[0] ), .b(\hdr_hld/high/U1664/y[1] ), .c(
        \hdr_hld/high/U1664/y[0] ), .d(\hdr_hld/high/U1664/U37/Z ), .e(
        \hdr_hld/high/U1664/y[1] ), .f(\hdr_hld/high/U1664/U37/Z ) );
    inv_1 \hdr_hld/high/U1664/U37/U30/Uinv  ( .x(\hdr_hld/high/U1664/U37/Z ), 
        .a(\hdr_hld/high/localcd ) );
    nor3_1 \hdr_hld/high/U1669/Unr  ( .x(\hdr_hld/high/U1669/nr ), .a(
        \hdr_hld/high/ctrlack_internal ), .b(\hdr_hld/high/drivel ), .c(n6) );
    nand3_1 \hdr_hld/high/U1669/Und  ( .x(\hdr_hld/high/U1669/nd ), .a(
        \hdr_hld/high/ctrlack_internal ), .b(\hdr_hld/high/drivel ), .c(n6) );
    oa21_1 \hdr_hld/high/U1669/U1  ( .x(\hdr_hld/high/U1669/n2 ), .a(
        \hdr_hld/high/U1669/n2 ), .b(\hdr_hld/high/U1669/nr ), .c(
        \hdr_hld/high/U1669/nd ) );
    inv_2 \hdr_hld/high/U1669/U3  ( .x(\hdr_hld/net20 ), .a(
        \hdr_hld/high/U1669/n2 ) );
    buf_2 U1 ( .x(n2), .a(\hdr_hld/net20 ) );
    buf_2 U2 ( .x(n1), .a(\hdr_hld/net20 ) );
    buf_1 U3 ( .x(n3), .a(\hdr_hld/low/latch ) );
    buf_1 U4 ( .x(n4), .a(\hdr_hld/high/drivel ) );
    buf_3 U5 ( .x(n5), .a(\hdr_hld/high/driveh ) );
    buf_3 U6 ( .x(n6), .a(\hdr_hld/high/driveh ) );
    buf_1 U7 ( .x(n7), .a(\hdr_hld/high/latch ) );
    inv_2 U8 ( .x(reset), .a(nReset) );
    buf_3 U9 ( .x(pullcd), .a(n9) );
endmodule


module chain_irdemux_32new_5 ( ctrlack, oh, ol, pullreq, pull_h, pull_l, 
    pullcd, reset, ctrlreq );
output [31:0] oh;
output [31:0] ol;
input  [7:0] pull_h;
input  [7:0] pull_l;
input  pullcd, reset, ctrlreq;
output ctrlack, pullreq;
    wire net30, net31, \I0/net32 , \I0/net33 , \I0/low/latch , 
        \I0/low/nlocalcd , \I0/low/localcd , \I0/low/ncd[0] , \I0/low/ncd[1] , 
        \I0/low/ncd[2] , \I0/low/ncd[3] , \I0/low/ncd[4] , \I0/low/ncd[5] , 
        \I0/low/ncd[6] , \I0/low/ncd[7] , \I0/low/ctrlack_internal , 
        \I0/low/acb , \I0/low/ba , \I0/low/driveh , \I0/net20 , 
        \I0/low/drivel , n1, n2, \I0/low/U4/U28/U1/clr , 
        \I0/low/U4/U28/U1/set , \I0/low/U1/Z , \I0/low/U1664/x[3] , 
        \I0/low/U1664/U28/Z , \I0/low/U1664/x[0] , \I0/low/U1664/U32/Z , 
        \I0/low/U1664/x[2] , \I0/low/U1664/U29/Z , \I0/low/U1664/y[0] , 
        \I0/low/U1664/x[1] , \I0/low/U1664/U33/Z , \I0/low/U1664/y[1] , 
        \I0/low/U1664/U30/Z , \I0/low/U1664/U31/Z , \I0/low/U1664/U37/Z , 
        \I0/low/U1669/nr , \I0/low/U1669/nd , \I0/low/U1669/n2 , 
        \I0/high/latch , \I0/high/nlocalcd , \I0/high/localcd , 
        \I0/high/ncd[0] , \I0/high/ncd[1] , \I0/high/ncd[2] , \I0/high/ncd[3] , 
        \I0/high/ncd[4] , \I0/high/ncd[5] , \I0/high/ncd[6] , \I0/high/ncd[7] , 
        \I0/high/ctrlack_internal , \I0/high/acb , \I0/high/ba , 
        \I0/high/driveh , net17, \I0/high/drivel , n3, n4, 
        \I0/high/U4/U28/U1/clr , \I0/high/U4/U28/U1/set , \I0/high/U1/Z , 
        \I0/high/U1664/x[3] , \I0/high/U1664/U28/Z , \I0/high/U1664/x[0] , 
        \I0/high/U1664/U32/Z , \I0/high/U1664/x[2] , \I0/high/U1664/U29/Z , 
        \I0/high/U1664/y[0] , \I0/high/U1664/x[1] , \I0/high/U1664/U33/Z , 
        \I0/high/U1664/y[1] , \I0/high/U1664/U30/Z , \I0/high/U1664/U31/Z , 
        \I0/high/U1664/U37/Z , \I0/high/U1669/nr , \I0/high/U1669/nd , 
        \I0/high/U1669/n2 , \I1/net32 , \I1/net33 , \I1/low/latch , 
        \I1/low/nlocalcd , \I1/low/localcd , \I1/low/ncd[0] , \I1/low/ncd[1] , 
        \I1/low/ncd[2] , \I1/low/ncd[3] , \I1/low/ncd[4] , \I1/low/ncd[5] , 
        \I1/low/ncd[6] , \I1/low/ncd[7] , \I1/low/ctrlack_internal , 
        \I1/low/acb , \I1/low/ba , \I1/low/driveh , \I1/net20 , 
        \I1/low/drivel , n5, n6, \I1/low/U4/U28/U1/clr , 
        \I1/low/U4/U28/U1/set , \I1/low/U1/Z , \I1/low/U1664/x[3] , 
        \I1/low/U1664/U28/Z , \I1/low/U1664/x[0] , \I1/low/U1664/U32/Z , 
        \I1/low/U1664/x[2] , \I1/low/U1664/U29/Z , \I1/low/U1664/y[0] , 
        \I1/low/U1664/x[1] , \I1/low/U1664/U33/Z , \I1/low/U1664/y[1] , 
        \I1/low/U1664/U30/Z , \I1/low/U1664/U31/Z , \I1/low/U1664/U37/Z , 
        \I1/low/U1669/nr , \I1/low/U1669/nd , \I1/low/U1669/n2 , 
        \I1/high/latch , \I1/high/nlocalcd , \I1/high/localcd , 
        \I1/high/ncd[0] , \I1/high/ncd[1] , \I1/high/ncd[2] , \I1/high/ncd[3] , 
        \I1/high/ncd[4] , \I1/high/ncd[5] , \I1/high/ncd[6] , \I1/high/ncd[7] , 
        \I1/high/ctrlack_internal , \I1/high/acb , \I1/high/ba , n7, n8, n12, 
        n10, n11, \I1/high/U4/U28/U1/clr , \I1/high/U4/U28/U1/set , 
        \I1/high/U1/Z , \I1/high/U1664/x[3] , \I1/high/U1664/U28/Z , 
        \I1/high/U1664/x[0] , \I1/high/U1664/U32/Z , \I1/high/U1664/x[2] , 
        \I1/high/U1664/U29/Z , \I1/high/U1664/y[0] , \I1/high/U1664/x[1] , 
        \I1/high/U1664/U33/Z , \I1/high/U1664/y[1] , \I1/high/U1664/U30/Z , 
        \I1/high/U1664/U31/Z , \I1/high/U1664/U37/Z , \I1/high/U1669/nr , 
        \I1/high/U1669/nd , \I1/high/U1669/n2 , n9;
    nand2_1 \U3/U5  ( .x(pullreq), .a(net30), .b(net31) );
    nor2_1 \I0/U3/U5  ( .x(net30), .a(\I0/net32 ), .b(\I0/net33 ) );
    buf_2 \I0/low/U1653  ( .x(\I0/low/latch ), .a(\I0/net32 ) );
    nor2_1 \I0/low/U264/U5  ( .x(\I0/low/nlocalcd ), .a(reset), .b(
        \I0/low/localcd ) );
    nor2_1 \I0/low/U1659_0_/U5  ( .x(\I0/low/ncd[0] ), .a(ol[0]), .b(oh[0]) );
    nor2_1 \I0/low/U1659_1_/U5  ( .x(\I0/low/ncd[1] ), .a(ol[1]), .b(oh[1]) );
    nor2_1 \I0/low/U1659_2_/U5  ( .x(\I0/low/ncd[2] ), .a(ol[2]), .b(oh[2]) );
    nor2_1 \I0/low/U1659_3_/U5  ( .x(\I0/low/ncd[3] ), .a(ol[3]), .b(oh[3]) );
    nor2_1 \I0/low/U1659_4_/U5  ( .x(\I0/low/ncd[4] ), .a(ol[4]), .b(oh[4]) );
    nor2_1 \I0/low/U1659_5_/U5  ( .x(\I0/low/ncd[5] ), .a(ol[5]), .b(oh[5]) );
    nor2_1 \I0/low/U1659_6_/U5  ( .x(\I0/low/ncd[6] ), .a(ol[6]), .b(oh[6]) );
    nor2_1 \I0/low/U1659_7_/U5  ( .x(\I0/low/ncd[7] ), .a(ol[7]), .b(oh[7]) );
    nor2_1 \I0/low/U3/U5  ( .x(\I0/low/ctrlack_internal ), .a(\I0/low/acb ), 
        .b(\I0/low/ba ) );
    buf_2 \I0/low/U1665/U7  ( .x(\I0/low/driveh ), .a(\I0/net20 ) );
    buf_2 \I0/low/U1666/U7  ( .x(\I0/low/drivel ), .a(\I0/net20 ) );
    ao23_1 \I0/low/U1658_0_/U21/U1/U1  ( .x(ol[0]), .a(\I0/low/driveh ), .b(ol
        [0]), .c(n1), .d(pull_l[0]), .e(n2) );
    ao23_1 \I0/low/U1658_1_/U21/U1/U1  ( .x(ol[1]), .a(\I0/low/drivel ), .b(ol
        [1]), .c(\I0/low/driveh ), .d(pull_l[1]), .e(n2) );
    ao23_1 \I0/low/U1658_2_/U21/U1/U1  ( .x(ol[2]), .a(\I0/low/drivel ), .b(ol
        [2]), .c(\I0/low/driveh ), .d(pull_l[2]), .e(n2) );
    ao23_1 \I0/low/U1658_3_/U21/U1/U1  ( .x(ol[3]), .a(\I0/low/driveh ), .b(ol
        [3]), .c(\I0/low/drivel ), .d(pull_l[3]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_4_/U21/U1/U1  ( .x(ol[4]), .a(n1), .b(ol[4]), .c(
        \I0/low/drivel ), .d(pull_l[4]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_5_/U21/U1/U1  ( .x(ol[5]), .a(\I0/low/driveh ), .b(ol
        [5]), .c(n1), .d(pull_l[5]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_6_/U21/U1/U1  ( .x(ol[6]), .a(\I0/low/drivel ), .b(ol
        [6]), .c(\I0/low/driveh ), .d(pull_l[6]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_7_/U21/U1/U1  ( .x(ol[7]), .a(n1), .b(ol[7]), .c(n1), 
        .d(pull_l[7]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_0_/U21/U1/U1  ( .x(oh[0]), .a(\I0/low/driveh ), .b(oh
        [0]), .c(n1), .d(pull_h[0]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_1_/U21/U1/U1  ( .x(oh[1]), .a(n1), .b(oh[1]), .c(
        \I0/low/drivel ), .d(pull_h[1]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_2_/U21/U1/U1  ( .x(oh[2]), .a(\I0/low/drivel ), .b(oh
        [2]), .c(\I0/low/drivel ), .d(pull_h[2]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_3_/U21/U1/U1  ( .x(oh[3]), .a(n1), .b(oh[3]), .c(
        \I0/low/driveh ), .d(pull_h[3]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_4_/U21/U1/U1  ( .x(oh[4]), .a(n1), .b(oh[4]), .c(n1), 
        .d(pull_h[4]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_5_/U21/U1/U1  ( .x(oh[5]), .a(\I0/low/drivel ), .b(oh
        [5]), .c(n1), .d(pull_h[5]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_6_/U21/U1/U1  ( .x(oh[6]), .a(\I0/low/drivel ), .b(oh
        [6]), .c(\I0/low/driveh ), .d(pull_h[6]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_7_/U21/U1/U1  ( .x(oh[7]), .a(\I0/low/driveh ), .b(oh
        [7]), .c(\I0/low/drivel ), .d(pull_h[7]), .e(\I0/low/latch ) );
    aoai211_1 \I0/low/U4/U28/U1/U1  ( .x(\I0/low/U4/U28/U1/clr ), .a(
        \I0/net20 ), .b(\I0/low/acb ), .c(\I0/low/nlocalcd ), .d(\I0/net32 )
         );
    nand3_1 \I0/low/U4/U28/U1/U2  ( .x(\I0/low/U4/U28/U1/set ), .a(
        \I0/low/nlocalcd ), .b(\I0/net20 ), .c(\I0/low/acb ) );
    nand2_2 \I0/low/U4/U28/U1/U3  ( .x(\I0/net32 ), .a(\I0/low/U4/U28/U1/clr ), 
        .b(\I0/low/U4/U28/U1/set ) );
    oai21_1 \I0/low/U1/U30/U1/U1  ( .x(\I0/low/acb ), .a(\I0/low/U1/Z ), .b(
        \I0/low/ba ), .c(\I0/net20 ) );
    inv_1 \I0/low/U1/U30/U1/U2  ( .x(\I0/low/U1/Z ), .a(\I0/low/acb ) );
    ao222_1 \I0/low/U5/U18/U1/U1  ( .x(\I0/low/ba ), .a(\I0/low/latch ), .b(
        pullcd), .c(\I0/low/latch ), .d(\I0/low/ba ), .e(pullcd), .f(
        \I0/low/ba ) );
    aoi222_1 \I0/low/U1664/U28/U30/U1  ( .x(\I0/low/U1664/x[3] ), .a(
        \I0/low/ncd[7] ), .b(\I0/low/ncd[6] ), .c(\I0/low/ncd[7] ), .d(
        \I0/low/U1664/U28/Z ), .e(\I0/low/ncd[6] ), .f(\I0/low/U1664/U28/Z )
         );
    inv_1 \I0/low/U1664/U28/U30/Uinv  ( .x(\I0/low/U1664/U28/Z ), .a(
        \I0/low/U1664/x[3] ) );
    aoi222_1 \I0/low/U1664/U32/U30/U1  ( .x(\I0/low/U1664/x[0] ), .a(
        \I0/low/ncd[1] ), .b(\I0/low/ncd[0] ), .c(\I0/low/ncd[1] ), .d(
        \I0/low/U1664/U32/Z ), .e(\I0/low/ncd[0] ), .f(\I0/low/U1664/U32/Z )
         );
    inv_1 \I0/low/U1664/U32/U30/Uinv  ( .x(\I0/low/U1664/U32/Z ), .a(
        \I0/low/U1664/x[0] ) );
    aoi222_1 \I0/low/U1664/U29/U30/U1  ( .x(\I0/low/U1664/x[2] ), .a(
        \I0/low/ncd[5] ), .b(\I0/low/ncd[4] ), .c(\I0/low/ncd[5] ), .d(
        \I0/low/U1664/U29/Z ), .e(\I0/low/ncd[4] ), .f(\I0/low/U1664/U29/Z )
         );
    inv_1 \I0/low/U1664/U29/U30/Uinv  ( .x(\I0/low/U1664/U29/Z ), .a(
        \I0/low/U1664/x[2] ) );
    aoi222_1 \I0/low/U1664/U33/U30/U1  ( .x(\I0/low/U1664/y[0] ), .a(
        \I0/low/U1664/x[1] ), .b(\I0/low/U1664/x[0] ), .c(\I0/low/U1664/x[1] ), 
        .d(\I0/low/U1664/U33/Z ), .e(\I0/low/U1664/x[0] ), .f(
        \I0/low/U1664/U33/Z ) );
    inv_1 \I0/low/U1664/U33/U30/Uinv  ( .x(\I0/low/U1664/U33/Z ), .a(
        \I0/low/U1664/y[0] ) );
    aoi222_1 \I0/low/U1664/U30/U30/U1  ( .x(\I0/low/U1664/y[1] ), .a(
        \I0/low/U1664/x[3] ), .b(\I0/low/U1664/x[2] ), .c(\I0/low/U1664/x[3] ), 
        .d(\I0/low/U1664/U30/Z ), .e(\I0/low/U1664/x[2] ), .f(
        \I0/low/U1664/U30/Z ) );
    inv_1 \I0/low/U1664/U30/U30/Uinv  ( .x(\I0/low/U1664/U30/Z ), .a(
        \I0/low/U1664/y[1] ) );
    aoi222_1 \I0/low/U1664/U31/U30/U1  ( .x(\I0/low/U1664/x[1] ), .a(
        \I0/low/ncd[3] ), .b(\I0/low/ncd[2] ), .c(\I0/low/ncd[3] ), .d(
        \I0/low/U1664/U31/Z ), .e(\I0/low/ncd[2] ), .f(\I0/low/U1664/U31/Z )
         );
    inv_1 \I0/low/U1664/U31/U30/Uinv  ( .x(\I0/low/U1664/U31/Z ), .a(
        \I0/low/U1664/x[1] ) );
    aoi222_1 \I0/low/U1664/U37/U30/U1  ( .x(\I0/low/localcd ), .a(
        \I0/low/U1664/y[0] ), .b(\I0/low/U1664/y[1] ), .c(\I0/low/U1664/y[0] ), 
        .d(\I0/low/U1664/U37/Z ), .e(\I0/low/U1664/y[1] ), .f(
        \I0/low/U1664/U37/Z ) );
    inv_1 \I0/low/U1664/U37/U30/Uinv  ( .x(\I0/low/U1664/U37/Z ), .a(
        \I0/low/localcd ) );
    nor3_1 \I0/low/U1669/Unr  ( .x(\I0/low/U1669/nr ), .a(
        \I0/low/ctrlack_internal ), .b(n1), .c(\I0/low/driveh ) );
    nand3_1 \I0/low/U1669/Und  ( .x(\I0/low/U1669/nd ), .a(
        \I0/low/ctrlack_internal ), .b(\I0/low/drivel ), .c(\I0/low/driveh )
         );
    oa21_1 \I0/low/U1669/U1  ( .x(\I0/low/U1669/n2 ), .a(\I0/low/U1669/n2 ), 
        .b(\I0/low/U1669/nr ), .c(\I0/low/U1669/nd ) );
    inv_2 \I0/low/U1669/U3  ( .x(ctrlack), .a(\I0/low/U1669/n2 ) );
    buf_2 \I0/high/U1653  ( .x(\I0/high/latch ), .a(\I0/net33 ) );
    nor2_1 \I0/high/U264/U5  ( .x(\I0/high/nlocalcd ), .a(reset), .b(
        \I0/high/localcd ) );
    nor2_1 \I0/high/U1659_0_/U5  ( .x(\I0/high/ncd[0] ), .a(ol[8]), .b(oh[8])
         );
    nor2_1 \I0/high/U1659_1_/U5  ( .x(\I0/high/ncd[1] ), .a(ol[9]), .b(oh[9])
         );
    nor2_1 \I0/high/U1659_2_/U5  ( .x(\I0/high/ncd[2] ), .a(ol[10]), .b(oh[10]
        ) );
    nor2_1 \I0/high/U1659_3_/U5  ( .x(\I0/high/ncd[3] ), .a(ol[11]), .b(oh[11]
        ) );
    nor2_1 \I0/high/U1659_4_/U5  ( .x(\I0/high/ncd[4] ), .a(ol[12]), .b(oh[12]
        ) );
    nor2_1 \I0/high/U1659_5_/U5  ( .x(\I0/high/ncd[5] ), .a(ol[13]), .b(oh[13]
        ) );
    nor2_1 \I0/high/U1659_6_/U5  ( .x(\I0/high/ncd[6] ), .a(ol[14]), .b(oh[14]
        ) );
    nor2_1 \I0/high/U1659_7_/U5  ( .x(\I0/high/ncd[7] ), .a(ol[15]), .b(oh[15]
        ) );
    nor2_1 \I0/high/U3/U5  ( .x(\I0/high/ctrlack_internal ), .a(\I0/high/acb ), 
        .b(\I0/high/ba ) );
    buf_2 \I0/high/U1665/U7  ( .x(\I0/high/driveh ), .a(net17) );
    buf_2 \I0/high/U1666/U7  ( .x(\I0/high/drivel ), .a(net17) );
    ao23_1 \I0/high/U1658_0_/U21/U1/U1  ( .x(ol[8]), .a(\I0/high/driveh ), .b(
        ol[8]), .c(n3), .d(pull_l[0]), .e(n4) );
    ao23_1 \I0/high/U1658_1_/U21/U1/U1  ( .x(ol[9]), .a(\I0/high/drivel ), .b(
        ol[9]), .c(\I0/high/driveh ), .d(pull_l[1]), .e(n4) );
    ao23_1 \I0/high/U1658_2_/U21/U1/U1  ( .x(ol[10]), .a(\I0/high/drivel ), 
        .b(ol[10]), .c(\I0/high/driveh ), .d(pull_l[2]), .e(n4) );
    ao23_1 \I0/high/U1658_3_/U21/U1/U1  ( .x(ol[11]), .a(\I0/high/driveh ), 
        .b(ol[11]), .c(\I0/high/drivel ), .d(pull_l[3]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1658_4_/U21/U1/U1  ( .x(ol[12]), .a(n3), .b(ol[12]), .c(
        \I0/high/drivel ), .d(pull_l[4]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1658_5_/U21/U1/U1  ( .x(ol[13]), .a(\I0/high/driveh ), 
        .b(ol[13]), .c(n3), .d(pull_l[5]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1658_6_/U21/U1/U1  ( .x(ol[14]), .a(\I0/high/drivel ), 
        .b(ol[14]), .c(\I0/high/driveh ), .d(pull_l[6]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1658_7_/U21/U1/U1  ( .x(ol[15]), .a(n3), .b(ol[15]), .c(
        n3), .d(pull_l[7]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_0_/U21/U1/U1  ( .x(oh[8]), .a(\I0/high/driveh ), .b(
        oh[8]), .c(n3), .d(pull_h[0]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_1_/U21/U1/U1  ( .x(oh[9]), .a(n3), .b(oh[9]), .c(
        \I0/high/drivel ), .d(pull_h[1]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_2_/U21/U1/U1  ( .x(oh[10]), .a(\I0/high/drivel ), 
        .b(oh[10]), .c(\I0/high/drivel ), .d(pull_h[2]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1651_3_/U21/U1/U1  ( .x(oh[11]), .a(n3), .b(oh[11]), .c(
        \I0/high/driveh ), .d(pull_h[3]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_4_/U21/U1/U1  ( .x(oh[12]), .a(n3), .b(oh[12]), .c(
        n3), .d(pull_h[4]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_5_/U21/U1/U1  ( .x(oh[13]), .a(\I0/high/drivel ), 
        .b(oh[13]), .c(n3), .d(pull_h[5]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_6_/U21/U1/U1  ( .x(oh[14]), .a(\I0/high/drivel ), 
        .b(oh[14]), .c(\I0/high/driveh ), .d(pull_h[6]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1651_7_/U21/U1/U1  ( .x(oh[15]), .a(\I0/high/driveh ), 
        .b(oh[15]), .c(\I0/high/drivel ), .d(pull_h[7]), .e(\I0/high/latch )
         );
    aoai211_1 \I0/high/U4/U28/U1/U1  ( .x(\I0/high/U4/U28/U1/clr ), .a(net17), 
        .b(\I0/high/acb ), .c(\I0/high/nlocalcd ), .d(\I0/net33 ) );
    nand3_1 \I0/high/U4/U28/U1/U2  ( .x(\I0/high/U4/U28/U1/set ), .a(
        \I0/high/nlocalcd ), .b(net17), .c(\I0/high/acb ) );
    nand2_2 \I0/high/U4/U28/U1/U3  ( .x(\I0/net33 ), .a(
        \I0/high/U4/U28/U1/clr ), .b(\I0/high/U4/U28/U1/set ) );
    oai21_1 \I0/high/U1/U30/U1/U1  ( .x(\I0/high/acb ), .a(\I0/high/U1/Z ), 
        .b(\I0/high/ba ), .c(net17) );
    inv_1 \I0/high/U1/U30/U1/U2  ( .x(\I0/high/U1/Z ), .a(\I0/high/acb ) );
    ao222_1 \I0/high/U5/U18/U1/U1  ( .x(\I0/high/ba ), .a(\I0/high/latch ), 
        .b(pullcd), .c(\I0/high/latch ), .d(\I0/high/ba ), .e(pullcd), .f(
        \I0/high/ba ) );
    aoi222_1 \I0/high/U1664/U28/U30/U1  ( .x(\I0/high/U1664/x[3] ), .a(
        \I0/high/ncd[7] ), .b(\I0/high/ncd[6] ), .c(\I0/high/ncd[7] ), .d(
        \I0/high/U1664/U28/Z ), .e(\I0/high/ncd[6] ), .f(\I0/high/U1664/U28/Z 
        ) );
    inv_1 \I0/high/U1664/U28/U30/Uinv  ( .x(\I0/high/U1664/U28/Z ), .a(
        \I0/high/U1664/x[3] ) );
    aoi222_1 \I0/high/U1664/U32/U30/U1  ( .x(\I0/high/U1664/x[0] ), .a(
        \I0/high/ncd[1] ), .b(\I0/high/ncd[0] ), .c(\I0/high/ncd[1] ), .d(
        \I0/high/U1664/U32/Z ), .e(\I0/high/ncd[0] ), .f(\I0/high/U1664/U32/Z 
        ) );
    inv_1 \I0/high/U1664/U32/U30/Uinv  ( .x(\I0/high/U1664/U32/Z ), .a(
        \I0/high/U1664/x[0] ) );
    aoi222_1 \I0/high/U1664/U29/U30/U1  ( .x(\I0/high/U1664/x[2] ), .a(
        \I0/high/ncd[5] ), .b(\I0/high/ncd[4] ), .c(\I0/high/ncd[5] ), .d(
        \I0/high/U1664/U29/Z ), .e(\I0/high/ncd[4] ), .f(\I0/high/U1664/U29/Z 
        ) );
    inv_1 \I0/high/U1664/U29/U30/Uinv  ( .x(\I0/high/U1664/U29/Z ), .a(
        \I0/high/U1664/x[2] ) );
    aoi222_1 \I0/high/U1664/U33/U30/U1  ( .x(\I0/high/U1664/y[0] ), .a(
        \I0/high/U1664/x[1] ), .b(\I0/high/U1664/x[0] ), .c(
        \I0/high/U1664/x[1] ), .d(\I0/high/U1664/U33/Z ), .e(
        \I0/high/U1664/x[0] ), .f(\I0/high/U1664/U33/Z ) );
    inv_1 \I0/high/U1664/U33/U30/Uinv  ( .x(\I0/high/U1664/U33/Z ), .a(
        \I0/high/U1664/y[0] ) );
    aoi222_1 \I0/high/U1664/U30/U30/U1  ( .x(\I0/high/U1664/y[1] ), .a(
        \I0/high/U1664/x[3] ), .b(\I0/high/U1664/x[2] ), .c(
        \I0/high/U1664/x[3] ), .d(\I0/high/U1664/U30/Z ), .e(
        \I0/high/U1664/x[2] ), .f(\I0/high/U1664/U30/Z ) );
    inv_1 \I0/high/U1664/U30/U30/Uinv  ( .x(\I0/high/U1664/U30/Z ), .a(
        \I0/high/U1664/y[1] ) );
    aoi222_1 \I0/high/U1664/U31/U30/U1  ( .x(\I0/high/U1664/x[1] ), .a(
        \I0/high/ncd[3] ), .b(\I0/high/ncd[2] ), .c(\I0/high/ncd[3] ), .d(
        \I0/high/U1664/U31/Z ), .e(\I0/high/ncd[2] ), .f(\I0/high/U1664/U31/Z 
        ) );
    inv_1 \I0/high/U1664/U31/U30/Uinv  ( .x(\I0/high/U1664/U31/Z ), .a(
        \I0/high/U1664/x[1] ) );
    aoi222_1 \I0/high/U1664/U37/U30/U1  ( .x(\I0/high/localcd ), .a(
        \I0/high/U1664/y[0] ), .b(\I0/high/U1664/y[1] ), .c(
        \I0/high/U1664/y[0] ), .d(\I0/high/U1664/U37/Z ), .e(
        \I0/high/U1664/y[1] ), .f(\I0/high/U1664/U37/Z ) );
    inv_1 \I0/high/U1664/U37/U30/Uinv  ( .x(\I0/high/U1664/U37/Z ), .a(
        \I0/high/localcd ) );
    nor3_1 \I0/high/U1669/Unr  ( .x(\I0/high/U1669/nr ), .a(
        \I0/high/ctrlack_internal ), .b(n3), .c(\I0/high/driveh ) );
    nand3_1 \I0/high/U1669/Und  ( .x(\I0/high/U1669/nd ), .a(
        \I0/high/ctrlack_internal ), .b(\I0/high/drivel ), .c(\I0/high/driveh 
        ) );
    oa21_1 \I0/high/U1669/U1  ( .x(\I0/high/U1669/n2 ), .a(\I0/high/U1669/n2 ), 
        .b(\I0/high/U1669/nr ), .c(\I0/high/U1669/nd ) );
    inv_2 \I0/high/U1669/U3  ( .x(\I0/net20 ), .a(\I0/high/U1669/n2 ) );
    nor2_1 \I1/U3/U5  ( .x(net31), .a(\I1/net32 ), .b(\I1/net33 ) );
    buf_2 \I1/low/U1653  ( .x(\I1/low/latch ), .a(\I1/net32 ) );
    nor2_1 \I1/low/U264/U5  ( .x(\I1/low/nlocalcd ), .a(reset), .b(
        \I1/low/localcd ) );
    nor2_1 \I1/low/U1659_0_/U5  ( .x(\I1/low/ncd[0] ), .a(ol[16]), .b(oh[16])
         );
    nor2_1 \I1/low/U1659_1_/U5  ( .x(\I1/low/ncd[1] ), .a(ol[17]), .b(oh[17])
         );
    nor2_1 \I1/low/U1659_2_/U5  ( .x(\I1/low/ncd[2] ), .a(ol[18]), .b(oh[18])
         );
    nor2_1 \I1/low/U1659_3_/U5  ( .x(\I1/low/ncd[3] ), .a(ol[19]), .b(oh[19])
         );
    nor2_1 \I1/low/U1659_4_/U5  ( .x(\I1/low/ncd[4] ), .a(ol[20]), .b(oh[20])
         );
    nor2_1 \I1/low/U1659_5_/U5  ( .x(\I1/low/ncd[5] ), .a(ol[21]), .b(oh[21])
         );
    nor2_1 \I1/low/U1659_6_/U5  ( .x(\I1/low/ncd[6] ), .a(ol[22]), .b(oh[22])
         );
    nor2_1 \I1/low/U1659_7_/U5  ( .x(\I1/low/ncd[7] ), .a(ol[23]), .b(oh[23])
         );
    nor2_1 \I1/low/U3/U5  ( .x(\I1/low/ctrlack_internal ), .a(\I1/low/acb ), 
        .b(\I1/low/ba ) );
    buf_2 \I1/low/U1665/U7  ( .x(\I1/low/driveh ), .a(\I1/net20 ) );
    buf_2 \I1/low/U1666/U7  ( .x(\I1/low/drivel ), .a(\I1/net20 ) );
    ao23_1 \I1/low/U1658_0_/U21/U1/U1  ( .x(ol[16]), .a(\I1/low/drivel ), .b(
        ol[16]), .c(n5), .d(pull_l[0]), .e(n6) );
    ao23_1 \I1/low/U1658_1_/U21/U1/U1  ( .x(ol[17]), .a(\I1/low/driveh ), .b(
        ol[17]), .c(n5), .d(pull_l[1]), .e(n6) );
    ao23_1 \I1/low/U1658_2_/U21/U1/U1  ( .x(ol[18]), .a(\I1/low/drivel ), .b(
        ol[18]), .c(\I1/low/driveh ), .d(pull_l[2]), .e(n6) );
    ao23_1 \I1/low/U1658_3_/U21/U1/U1  ( .x(ol[19]), .a(n5), .b(ol[19]), .c(
        \I1/low/driveh ), .d(pull_l[3]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_4_/U21/U1/U1  ( .x(ol[20]), .a(\I1/low/driveh ), .b(
        ol[20]), .c(\I1/low/drivel ), .d(pull_l[4]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_5_/U21/U1/U1  ( .x(ol[21]), .a(n5), .b(ol[21]), .c(
        \I1/low/drivel ), .d(pull_l[5]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_6_/U21/U1/U1  ( .x(ol[22]), .a(\I1/low/driveh ), .b(
        ol[22]), .c(n5), .d(pull_l[6]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_7_/U21/U1/U1  ( .x(ol[23]), .a(\I1/low/drivel ), .b(
        ol[23]), .c(\I1/low/driveh ), .d(pull_l[7]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_0_/U21/U1/U1  ( .x(oh[16]), .a(\I1/low/driveh ), .b(
        oh[16]), .c(\I1/low/drivel ), .d(pull_h[0]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_1_/U21/U1/U1  ( .x(oh[17]), .a(\I1/low/drivel ), .b(
        oh[17]), .c(n5), .d(pull_h[1]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_2_/U21/U1/U1  ( .x(oh[18]), .a(\I1/low/drivel ), .b(
        oh[18]), .c(\I1/low/driveh ), .d(pull_h[2]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_3_/U21/U1/U1  ( .x(oh[19]), .a(n5), .b(oh[19]), .c(n5
        ), .d(pull_h[3]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_4_/U21/U1/U1  ( .x(oh[20]), .a(n5), .b(oh[20]), .c(n5
        ), .d(pull_h[4]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_5_/U21/U1/U1  ( .x(oh[21]), .a(\I1/low/drivel ), .b(
        oh[21]), .c(\I1/low/driveh ), .d(pull_h[5]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_6_/U21/U1/U1  ( .x(oh[22]), .a(n5), .b(oh[22]), .c(
        \I1/low/drivel ), .d(pull_h[6]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_7_/U21/U1/U1  ( .x(oh[23]), .a(\I1/low/driveh ), .b(
        oh[23]), .c(\I1/low/drivel ), .d(pull_h[7]), .e(\I1/low/latch ) );
    aoai211_1 \I1/low/U4/U28/U1/U1  ( .x(\I1/low/U4/U28/U1/clr ), .a(
        \I1/net20 ), .b(\I1/low/acb ), .c(\I1/low/nlocalcd ), .d(\I1/net32 )
         );
    nand3_1 \I1/low/U4/U28/U1/U2  ( .x(\I1/low/U4/U28/U1/set ), .a(
        \I1/low/nlocalcd ), .b(\I1/net20 ), .c(\I1/low/acb ) );
    nand2_2 \I1/low/U4/U28/U1/U3  ( .x(\I1/net32 ), .a(\I1/low/U4/U28/U1/clr ), 
        .b(\I1/low/U4/U28/U1/set ) );
    oai21_1 \I1/low/U1/U30/U1/U1  ( .x(\I1/low/acb ), .a(\I1/low/U1/Z ), .b(
        \I1/low/ba ), .c(\I1/net20 ) );
    inv_1 \I1/low/U1/U30/U1/U2  ( .x(\I1/low/U1/Z ), .a(\I1/low/acb ) );
    ao222_1 \I1/low/U5/U18/U1/U1  ( .x(\I1/low/ba ), .a(\I1/low/latch ), .b(
        pullcd), .c(\I1/low/latch ), .d(\I1/low/ba ), .e(pullcd), .f(
        \I1/low/ba ) );
    aoi222_1 \I1/low/U1664/U28/U30/U1  ( .x(\I1/low/U1664/x[3] ), .a(
        \I1/low/ncd[7] ), .b(\I1/low/ncd[6] ), .c(\I1/low/ncd[7] ), .d(
        \I1/low/U1664/U28/Z ), .e(\I1/low/ncd[6] ), .f(\I1/low/U1664/U28/Z )
         );
    inv_1 \I1/low/U1664/U28/U30/Uinv  ( .x(\I1/low/U1664/U28/Z ), .a(
        \I1/low/U1664/x[3] ) );
    aoi222_1 \I1/low/U1664/U32/U30/U1  ( .x(\I1/low/U1664/x[0] ), .a(
        \I1/low/ncd[1] ), .b(\I1/low/ncd[0] ), .c(\I1/low/ncd[1] ), .d(
        \I1/low/U1664/U32/Z ), .e(\I1/low/ncd[0] ), .f(\I1/low/U1664/U32/Z )
         );
    inv_1 \I1/low/U1664/U32/U30/Uinv  ( .x(\I1/low/U1664/U32/Z ), .a(
        \I1/low/U1664/x[0] ) );
    aoi222_1 \I1/low/U1664/U29/U30/U1  ( .x(\I1/low/U1664/x[2] ), .a(
        \I1/low/ncd[5] ), .b(\I1/low/ncd[4] ), .c(\I1/low/ncd[5] ), .d(
        \I1/low/U1664/U29/Z ), .e(\I1/low/ncd[4] ), .f(\I1/low/U1664/U29/Z )
         );
    inv_1 \I1/low/U1664/U29/U30/Uinv  ( .x(\I1/low/U1664/U29/Z ), .a(
        \I1/low/U1664/x[2] ) );
    aoi222_1 \I1/low/U1664/U33/U30/U1  ( .x(\I1/low/U1664/y[0] ), .a(
        \I1/low/U1664/x[1] ), .b(\I1/low/U1664/x[0] ), .c(\I1/low/U1664/x[1] ), 
        .d(\I1/low/U1664/U33/Z ), .e(\I1/low/U1664/x[0] ), .f(
        \I1/low/U1664/U33/Z ) );
    inv_1 \I1/low/U1664/U33/U30/Uinv  ( .x(\I1/low/U1664/U33/Z ), .a(
        \I1/low/U1664/y[0] ) );
    aoi222_1 \I1/low/U1664/U30/U30/U1  ( .x(\I1/low/U1664/y[1] ), .a(
        \I1/low/U1664/x[3] ), .b(\I1/low/U1664/x[2] ), .c(\I1/low/U1664/x[3] ), 
        .d(\I1/low/U1664/U30/Z ), .e(\I1/low/U1664/x[2] ), .f(
        \I1/low/U1664/U30/Z ) );
    inv_1 \I1/low/U1664/U30/U30/Uinv  ( .x(\I1/low/U1664/U30/Z ), .a(
        \I1/low/U1664/y[1] ) );
    aoi222_1 \I1/low/U1664/U31/U30/U1  ( .x(\I1/low/U1664/x[1] ), .a(
        \I1/low/ncd[3] ), .b(\I1/low/ncd[2] ), .c(\I1/low/ncd[3] ), .d(
        \I1/low/U1664/U31/Z ), .e(\I1/low/ncd[2] ), .f(\I1/low/U1664/U31/Z )
         );
    inv_1 \I1/low/U1664/U31/U30/Uinv  ( .x(\I1/low/U1664/U31/Z ), .a(
        \I1/low/U1664/x[1] ) );
    aoi222_1 \I1/low/U1664/U37/U30/U1  ( .x(\I1/low/localcd ), .a(
        \I1/low/U1664/y[0] ), .b(\I1/low/U1664/y[1] ), .c(\I1/low/U1664/y[0] ), 
        .d(\I1/low/U1664/U37/Z ), .e(\I1/low/U1664/y[1] ), .f(
        \I1/low/U1664/U37/Z ) );
    inv_1 \I1/low/U1664/U37/U30/Uinv  ( .x(\I1/low/U1664/U37/Z ), .a(
        \I1/low/localcd ) );
    nor3_1 \I1/low/U1669/Unr  ( .x(\I1/low/U1669/nr ), .a(
        \I1/low/ctrlack_internal ), .b(n5), .c(\I1/low/driveh ) );
    nand3_1 \I1/low/U1669/Und  ( .x(\I1/low/U1669/nd ), .a(
        \I1/low/ctrlack_internal ), .b(\I1/low/drivel ), .c(\I1/low/driveh )
         );
    oa21_1 \I1/low/U1669/U1  ( .x(\I1/low/U1669/n2 ), .a(\I1/low/U1669/n2 ), 
        .b(\I1/low/U1669/nr ), .c(\I1/low/U1669/nd ) );
    inv_2 \I1/low/U1669/U3  ( .x(net17), .a(\I1/low/U1669/n2 ) );
    buf_2 \I1/high/U1653  ( .x(\I1/high/latch ), .a(\I1/net33 ) );
    nor2_1 \I1/high/U264/U5  ( .x(\I1/high/nlocalcd ), .a(reset), .b(
        \I1/high/localcd ) );
    nor2_1 \I1/high/U1659_0_/U5  ( .x(\I1/high/ncd[0] ), .a(ol[24]), .b(oh[24]
        ) );
    nor2_1 \I1/high/U1659_1_/U5  ( .x(\I1/high/ncd[1] ), .a(ol[25]), .b(oh[25]
        ) );
    nor2_1 \I1/high/U1659_2_/U5  ( .x(\I1/high/ncd[2] ), .a(ol[26]), .b(oh[26]
        ) );
    nor2_1 \I1/high/U1659_3_/U5  ( .x(\I1/high/ncd[3] ), .a(ol[27]), .b(oh[27]
        ) );
    nor2_1 \I1/high/U1659_4_/U5  ( .x(\I1/high/ncd[4] ), .a(ol[28]), .b(oh[28]
        ) );
    nor2_1 \I1/high/U1659_5_/U5  ( .x(\I1/high/ncd[5] ), .a(ol[29]), .b(oh[29]
        ) );
    nor2_1 \I1/high/U1659_6_/U5  ( .x(\I1/high/ncd[6] ), .a(ol[30]), .b(oh[30]
        ) );
    nor2_1 \I1/high/U1659_7_/U5  ( .x(\I1/high/ncd[7] ), .a(ol[31]), .b(oh[31]
        ) );
    nor2_1 \I1/high/U3/U5  ( .x(\I1/high/ctrlack_internal ), .a(\I1/high/acb ), 
        .b(\I1/high/ba ) );
    ao23_1 \I1/high/U1658_0_/U21/U1/U1  ( .x(ol[24]), .a(n7), .b(ol[24]), .c(
        n8), .d(pull_l[0]), .e(n12) );
    ao23_1 \I1/high/U1658_1_/U21/U1/U1  ( .x(ol[25]), .a(n7), .b(ol[25]), .c(
        n8), .d(pull_l[1]), .e(n12) );
    ao23_1 \I1/high/U1658_2_/U21/U1/U1  ( .x(ol[26]), .a(n7), .b(ol[26]), .c(
        n7), .d(pull_l[2]), .e(n12) );
    ao23_1 \I1/high/U1658_3_/U21/U1/U1  ( .x(ol[27]), .a(n7), .b(ol[27]), .c(
        n7), .d(pull_l[3]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1658_4_/U21/U1/U1  ( .x(ol[28]), .a(n7), .b(ol[28]), .c(
        n7), .d(pull_l[4]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1658_5_/U21/U1/U1  ( .x(ol[29]), .a(n7), .b(ol[29]), .c(
        n8), .d(pull_l[5]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1658_6_/U21/U1/U1  ( .x(ol[30]), .a(n7), .b(ol[30]), .c(
        n8), .d(pull_l[6]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1658_7_/U21/U1/U1  ( .x(ol[31]), .a(n7), .b(ol[31]), .c(
        n8), .d(pull_l[7]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_0_/U21/U1/U1  ( .x(oh[24]), .a(n10), .b(oh[24]), .c(
        n10), .d(pull_h[0]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_1_/U21/U1/U1  ( .x(oh[25]), .a(n10), .b(oh[25]), .c(
        n11), .d(pull_h[1]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_2_/U21/U1/U1  ( .x(oh[26]), .a(n10), .b(oh[26]), .c(
        n11), .d(pull_h[2]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_3_/U21/U1/U1  ( .x(oh[27]), .a(n10), .b(oh[27]), .c(
        n10), .d(pull_h[3]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_4_/U21/U1/U1  ( .x(oh[28]), .a(n10), .b(oh[28]), .c(
        n11), .d(pull_h[4]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_5_/U21/U1/U1  ( .x(oh[29]), .a(n10), .b(oh[29]), .c(
        n11), .d(pull_h[5]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_6_/U21/U1/U1  ( .x(oh[30]), .a(n10), .b(oh[30]), .c(
        n11), .d(pull_h[6]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_7_/U21/U1/U1  ( .x(oh[31]), .a(n10), .b(oh[31]), .c(
        n10), .d(pull_h[7]), .e(\I1/high/latch ) );
    aoai211_1 \I1/high/U4/U28/U1/U1  ( .x(\I1/high/U4/U28/U1/clr ), .a(ctrlreq
        ), .b(\I1/high/acb ), .c(\I1/high/nlocalcd ), .d(\I1/net33 ) );
    nand3_1 \I1/high/U4/U28/U1/U2  ( .x(\I1/high/U4/U28/U1/set ), .a(
        \I1/high/nlocalcd ), .b(ctrlreq), .c(\I1/high/acb ) );
    nand2_2 \I1/high/U4/U28/U1/U3  ( .x(\I1/net33 ), .a(
        \I1/high/U4/U28/U1/clr ), .b(\I1/high/U4/U28/U1/set ) );
    oai21_1 \I1/high/U1/U30/U1/U1  ( .x(\I1/high/acb ), .a(\I1/high/U1/Z ), 
        .b(\I1/high/ba ), .c(ctrlreq) );
    inv_1 \I1/high/U1/U30/U1/U2  ( .x(\I1/high/U1/Z ), .a(\I1/high/acb ) );
    ao222_1 \I1/high/U5/U18/U1/U1  ( .x(\I1/high/ba ), .a(\I1/high/latch ), 
        .b(pullcd), .c(\I1/high/latch ), .d(\I1/high/ba ), .e(pullcd), .f(
        \I1/high/ba ) );
    aoi222_1 \I1/high/U1664/U28/U30/U1  ( .x(\I1/high/U1664/x[3] ), .a(
        \I1/high/ncd[7] ), .b(\I1/high/ncd[6] ), .c(\I1/high/ncd[7] ), .d(
        \I1/high/U1664/U28/Z ), .e(\I1/high/ncd[6] ), .f(\I1/high/U1664/U28/Z 
        ) );
    inv_1 \I1/high/U1664/U28/U30/Uinv  ( .x(\I1/high/U1664/U28/Z ), .a(
        \I1/high/U1664/x[3] ) );
    aoi222_1 \I1/high/U1664/U32/U30/U1  ( .x(\I1/high/U1664/x[0] ), .a(
        \I1/high/ncd[1] ), .b(\I1/high/ncd[0] ), .c(\I1/high/ncd[1] ), .d(
        \I1/high/U1664/U32/Z ), .e(\I1/high/ncd[0] ), .f(\I1/high/U1664/U32/Z 
        ) );
    inv_1 \I1/high/U1664/U32/U30/Uinv  ( .x(\I1/high/U1664/U32/Z ), .a(
        \I1/high/U1664/x[0] ) );
    aoi222_1 \I1/high/U1664/U29/U30/U1  ( .x(\I1/high/U1664/x[2] ), .a(
        \I1/high/ncd[5] ), .b(\I1/high/ncd[4] ), .c(\I1/high/ncd[5] ), .d(
        \I1/high/U1664/U29/Z ), .e(\I1/high/ncd[4] ), .f(\I1/high/U1664/U29/Z 
        ) );
    inv_1 \I1/high/U1664/U29/U30/Uinv  ( .x(\I1/high/U1664/U29/Z ), .a(
        \I1/high/U1664/x[2] ) );
    aoi222_1 \I1/high/U1664/U33/U30/U1  ( .x(\I1/high/U1664/y[0] ), .a(
        \I1/high/U1664/x[1] ), .b(\I1/high/U1664/x[0] ), .c(
        \I1/high/U1664/x[1] ), .d(\I1/high/U1664/U33/Z ), .e(
        \I1/high/U1664/x[0] ), .f(\I1/high/U1664/U33/Z ) );
    inv_1 \I1/high/U1664/U33/U30/Uinv  ( .x(\I1/high/U1664/U33/Z ), .a(
        \I1/high/U1664/y[0] ) );
    aoi222_1 \I1/high/U1664/U30/U30/U1  ( .x(\I1/high/U1664/y[1] ), .a(
        \I1/high/U1664/x[3] ), .b(\I1/high/U1664/x[2] ), .c(
        \I1/high/U1664/x[3] ), .d(\I1/high/U1664/U30/Z ), .e(
        \I1/high/U1664/x[2] ), .f(\I1/high/U1664/U30/Z ) );
    inv_1 \I1/high/U1664/U30/U30/Uinv  ( .x(\I1/high/U1664/U30/Z ), .a(
        \I1/high/U1664/y[1] ) );
    aoi222_1 \I1/high/U1664/U31/U30/U1  ( .x(\I1/high/U1664/x[1] ), .a(
        \I1/high/ncd[3] ), .b(\I1/high/ncd[2] ), .c(\I1/high/ncd[3] ), .d(
        \I1/high/U1664/U31/Z ), .e(\I1/high/ncd[2] ), .f(\I1/high/U1664/U31/Z 
        ) );
    inv_1 \I1/high/U1664/U31/U30/Uinv  ( .x(\I1/high/U1664/U31/Z ), .a(
        \I1/high/U1664/x[1] ) );
    aoi222_1 \I1/high/U1664/U37/U30/U1  ( .x(\I1/high/localcd ), .a(
        \I1/high/U1664/y[0] ), .b(\I1/high/U1664/y[1] ), .c(
        \I1/high/U1664/y[0] ), .d(\I1/high/U1664/U37/Z ), .e(
        \I1/high/U1664/y[1] ), .f(\I1/high/U1664/U37/Z ) );
    inv_1 \I1/high/U1664/U37/U30/Uinv  ( .x(\I1/high/U1664/U37/Z ), .a(
        \I1/high/localcd ) );
    nor3_1 \I1/high/U1669/Unr  ( .x(\I1/high/U1669/nr ), .a(
        \I1/high/ctrlack_internal ), .b(n8), .c(n11) );
    nand3_1 \I1/high/U1669/Und  ( .x(\I1/high/U1669/nd ), .a(
        \I1/high/ctrlack_internal ), .b(n8), .c(n11) );
    oa21_1 \I1/high/U1669/U1  ( .x(\I1/high/U1669/n2 ), .a(\I1/high/U1669/n2 ), 
        .b(\I1/high/U1669/nr ), .c(\I1/high/U1669/nd ) );
    inv_2 \I1/high/U1669/U3  ( .x(\I1/net20 ), .a(\I1/high/U1669/n2 ) );
    buf_2 U1 ( .x(n1), .a(\I0/net20 ) );
    buf_1 U2 ( .x(n2), .a(\I0/low/latch ) );
    buf_2 U3 ( .x(n3), .a(net17) );
    buf_1 U4 ( .x(n4), .a(\I0/high/latch ) );
    buf_2 U5 ( .x(n5), .a(\I1/net20 ) );
    buf_1 U6 ( .x(n6), .a(\I1/low/latch ) );
    inv_2 U7 ( .x(n7), .a(n9) );
    inv_1 U8 ( .x(n8), .a(n9) );
    inv_0 U9 ( .x(n9), .a(ctrlreq) );
    inv_2 U10 ( .x(n10), .a(n9) );
    inv_1 U11 ( .x(n11), .a(n9) );
    buf_1 U12 ( .x(n12), .a(\I1/high/latch ) );
endmodule


module chain_irdemux_32new_4 ( ctrlack, oh, ol, pullreq, pull_h, pull_l, 
    pullcd, reset, ctrlreq );
output [31:0] oh;
output [31:0] ol;
input  [7:0] pull_h;
input  [7:0] pull_l;
input  pullcd, reset, ctrlreq;
output ctrlack, pullreq;
    wire net30, net31, \I0/net32 , \I0/net33 , \I0/low/latch , 
        \I0/low/nlocalcd , \I0/low/localcd , \I0/low/ncd[0] , \I0/low/ncd[1] , 
        \I0/low/ncd[2] , \I0/low/ncd[3] , \I0/low/ncd[4] , \I0/low/ncd[5] , 
        \I0/low/ncd[6] , \I0/low/ncd[7] , \I0/low/ctrlack_internal , 
        \I0/low/acb , \I0/low/ba , \I0/low/driveh , \I0/net20 , 
        \I0/low/drivel , n1, n2, \I0/low/U4/U28/U1/clr , 
        \I0/low/U4/U28/U1/set , \I0/low/U1/Z , \I0/low/U1664/x[3] , 
        \I0/low/U1664/U28/Z , \I0/low/U1664/x[0] , \I0/low/U1664/U32/Z , 
        \I0/low/U1664/x[2] , \I0/low/U1664/U29/Z , \I0/low/U1664/y[0] , 
        \I0/low/U1664/x[1] , \I0/low/U1664/U33/Z , \I0/low/U1664/y[1] , 
        \I0/low/U1664/U30/Z , \I0/low/U1664/U31/Z , \I0/low/U1664/U37/Z , 
        \I0/low/U1669/nr , \I0/low/U1669/nd , \I0/low/U1669/n2 , 
        \I0/high/latch , \I0/high/nlocalcd , \I0/high/localcd , 
        \I0/high/ncd[0] , \I0/high/ncd[1] , \I0/high/ncd[2] , \I0/high/ncd[3] , 
        \I0/high/ncd[4] , \I0/high/ncd[5] , \I0/high/ncd[6] , \I0/high/ncd[7] , 
        \I0/high/ctrlack_internal , \I0/high/acb , \I0/high/ba , 
        \I0/high/driveh , net17, \I0/high/drivel , n3, n4, 
        \I0/high/U4/U28/U1/clr , \I0/high/U4/U28/U1/set , \I0/high/U1/Z , 
        \I0/high/U1664/x[3] , \I0/high/U1664/U28/Z , \I0/high/U1664/x[0] , 
        \I0/high/U1664/U32/Z , \I0/high/U1664/x[2] , \I0/high/U1664/U29/Z , 
        \I0/high/U1664/y[0] , \I0/high/U1664/x[1] , \I0/high/U1664/U33/Z , 
        \I0/high/U1664/y[1] , \I0/high/U1664/U30/Z , \I0/high/U1664/U31/Z , 
        \I0/high/U1664/U37/Z , \I0/high/U1669/nr , \I0/high/U1669/nd , 
        \I0/high/U1669/n2 , \I1/net32 , \I1/net33 , \I1/low/latch , 
        \I1/low/nlocalcd , \I1/low/localcd , \I1/low/ncd[0] , \I1/low/ncd[1] , 
        \I1/low/ncd[2] , \I1/low/ncd[3] , \I1/low/ncd[4] , \I1/low/ncd[5] , 
        \I1/low/ncd[6] , \I1/low/ncd[7] , \I1/low/ctrlack_internal , 
        \I1/low/acb , \I1/low/ba , \I1/low/driveh , \I1/net20 , 
        \I1/low/drivel , n5, n6, \I1/low/U4/U28/U1/clr , 
        \I1/low/U4/U28/U1/set , \I1/low/U1/Z , \I1/low/U1664/x[3] , 
        \I1/low/U1664/U28/Z , \I1/low/U1664/x[0] , \I1/low/U1664/U32/Z , 
        \I1/low/U1664/x[2] , \I1/low/U1664/U29/Z , \I1/low/U1664/y[0] , 
        \I1/low/U1664/x[1] , \I1/low/U1664/U33/Z , \I1/low/U1664/y[1] , 
        \I1/low/U1664/U30/Z , \I1/low/U1664/U31/Z , \I1/low/U1664/U37/Z , 
        \I1/low/U1669/nr , \I1/low/U1669/nd , \I1/low/U1669/n2 , 
        \I1/high/latch , \I1/high/nlocalcd , \I1/high/localcd , 
        \I1/high/ncd[0] , \I1/high/ncd[1] , \I1/high/ncd[2] , \I1/high/ncd[3] , 
        \I1/high/ncd[4] , \I1/high/ncd[5] , \I1/high/ncd[6] , \I1/high/ncd[7] , 
        \I1/high/ctrlack_internal , \I1/high/acb , \I1/high/ba , 
        \I1/high/driveh , \I1/high/drivel , n7, n8, \I1/high/U4/U28/U1/clr , 
        \I1/high/U4/U28/U1/set , \I1/high/U1/Z , \I1/high/U1664/x[3] , 
        \I1/high/U1664/U28/Z , \I1/high/U1664/x[0] , \I1/high/U1664/U32/Z , 
        \I1/high/U1664/x[2] , \I1/high/U1664/U29/Z , \I1/high/U1664/y[0] , 
        \I1/high/U1664/x[1] , \I1/high/U1664/U33/Z , \I1/high/U1664/y[1] , 
        \I1/high/U1664/U30/Z , \I1/high/U1664/U31/Z , \I1/high/U1664/U37/Z , 
        \I1/high/U1669/nr , \I1/high/U1669/nd , \I1/high/U1669/n2 ;
    nand2_1 \U3/U5  ( .x(pullreq), .a(net30), .b(net31) );
    nor2_1 \I0/U3/U5  ( .x(net30), .a(\I0/net32 ), .b(\I0/net33 ) );
    buf_2 \I0/low/U1653  ( .x(\I0/low/latch ), .a(\I0/net32 ) );
    nor2_1 \I0/low/U264/U5  ( .x(\I0/low/nlocalcd ), .a(reset), .b(
        \I0/low/localcd ) );
    nor2_1 \I0/low/U1659_0_/U5  ( .x(\I0/low/ncd[0] ), .a(ol[0]), .b(oh[0]) );
    nor2_1 \I0/low/U1659_1_/U5  ( .x(\I0/low/ncd[1] ), .a(ol[1]), .b(oh[1]) );
    nor2_1 \I0/low/U1659_2_/U5  ( .x(\I0/low/ncd[2] ), .a(ol[2]), .b(oh[2]) );
    nor2_1 \I0/low/U1659_3_/U5  ( .x(\I0/low/ncd[3] ), .a(ol[3]), .b(oh[3]) );
    nor2_1 \I0/low/U1659_4_/U5  ( .x(\I0/low/ncd[4] ), .a(ol[4]), .b(oh[4]) );
    nor2_1 \I0/low/U1659_5_/U5  ( .x(\I0/low/ncd[5] ), .a(ol[5]), .b(oh[5]) );
    nor2_1 \I0/low/U1659_6_/U5  ( .x(\I0/low/ncd[6] ), .a(ol[6]), .b(oh[6]) );
    nor2_1 \I0/low/U1659_7_/U5  ( .x(\I0/low/ncd[7] ), .a(ol[7]), .b(oh[7]) );
    nor2_1 \I0/low/U3/U5  ( .x(\I0/low/ctrlack_internal ), .a(\I0/low/acb ), 
        .b(\I0/low/ba ) );
    buf_2 \I0/low/U1665/U7  ( .x(\I0/low/driveh ), .a(\I0/net20 ) );
    buf_2 \I0/low/U1666/U7  ( .x(\I0/low/drivel ), .a(\I0/net20 ) );
    ao23_1 \I0/low/U1658_0_/U21/U1/U1  ( .x(ol[0]), .a(\I0/low/driveh ), .b(ol
        [0]), .c(n1), .d(pull_l[0]), .e(n2) );
    ao23_1 \I0/low/U1658_1_/U21/U1/U1  ( .x(ol[1]), .a(\I0/low/drivel ), .b(ol
        [1]), .c(\I0/low/driveh ), .d(pull_l[1]), .e(n2) );
    ao23_1 \I0/low/U1658_2_/U21/U1/U1  ( .x(ol[2]), .a(\I0/low/drivel ), .b(ol
        [2]), .c(\I0/low/driveh ), .d(pull_l[2]), .e(n2) );
    ao23_1 \I0/low/U1658_3_/U21/U1/U1  ( .x(ol[3]), .a(\I0/low/driveh ), .b(ol
        [3]), .c(\I0/low/drivel ), .d(pull_l[3]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_4_/U21/U1/U1  ( .x(ol[4]), .a(n1), .b(ol[4]), .c(
        \I0/low/drivel ), .d(pull_l[4]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_5_/U21/U1/U1  ( .x(ol[5]), .a(\I0/low/driveh ), .b(ol
        [5]), .c(n1), .d(pull_l[5]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_6_/U21/U1/U1  ( .x(ol[6]), .a(\I0/low/drivel ), .b(ol
        [6]), .c(\I0/low/driveh ), .d(pull_l[6]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_7_/U21/U1/U1  ( .x(ol[7]), .a(n1), .b(ol[7]), .c(n1), 
        .d(pull_l[7]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_0_/U21/U1/U1  ( .x(oh[0]), .a(\I0/low/driveh ), .b(oh
        [0]), .c(n1), .d(pull_h[0]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_1_/U21/U1/U1  ( .x(oh[1]), .a(n1), .b(oh[1]), .c(
        \I0/low/drivel ), .d(pull_h[1]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_2_/U21/U1/U1  ( .x(oh[2]), .a(\I0/low/drivel ), .b(oh
        [2]), .c(\I0/low/drivel ), .d(pull_h[2]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_3_/U21/U1/U1  ( .x(oh[3]), .a(n1), .b(oh[3]), .c(
        \I0/low/driveh ), .d(pull_h[3]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_4_/U21/U1/U1  ( .x(oh[4]), .a(n1), .b(oh[4]), .c(n1), 
        .d(pull_h[4]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_5_/U21/U1/U1  ( .x(oh[5]), .a(\I0/low/drivel ), .b(oh
        [5]), .c(n1), .d(pull_h[5]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_6_/U21/U1/U1  ( .x(oh[6]), .a(\I0/low/drivel ), .b(oh
        [6]), .c(\I0/low/driveh ), .d(pull_h[6]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_7_/U21/U1/U1  ( .x(oh[7]), .a(\I0/low/driveh ), .b(oh
        [7]), .c(\I0/low/drivel ), .d(pull_h[7]), .e(\I0/low/latch ) );
    aoai211_1 \I0/low/U4/U28/U1/U1  ( .x(\I0/low/U4/U28/U1/clr ), .a(
        \I0/net20 ), .b(\I0/low/acb ), .c(\I0/low/nlocalcd ), .d(\I0/net32 )
         );
    nand3_1 \I0/low/U4/U28/U1/U2  ( .x(\I0/low/U4/U28/U1/set ), .a(
        \I0/low/nlocalcd ), .b(\I0/net20 ), .c(\I0/low/acb ) );
    nand2_2 \I0/low/U4/U28/U1/U3  ( .x(\I0/net32 ), .a(\I0/low/U4/U28/U1/clr ), 
        .b(\I0/low/U4/U28/U1/set ) );
    oai21_1 \I0/low/U1/U30/U1/U1  ( .x(\I0/low/acb ), .a(\I0/low/U1/Z ), .b(
        \I0/low/ba ), .c(\I0/net20 ) );
    inv_1 \I0/low/U1/U30/U1/U2  ( .x(\I0/low/U1/Z ), .a(\I0/low/acb ) );
    ao222_1 \I0/low/U5/U18/U1/U1  ( .x(\I0/low/ba ), .a(\I0/low/latch ), .b(
        pullcd), .c(\I0/low/latch ), .d(\I0/low/ba ), .e(pullcd), .f(
        \I0/low/ba ) );
    aoi222_1 \I0/low/U1664/U28/U30/U1  ( .x(\I0/low/U1664/x[3] ), .a(
        \I0/low/ncd[7] ), .b(\I0/low/ncd[6] ), .c(\I0/low/ncd[7] ), .d(
        \I0/low/U1664/U28/Z ), .e(\I0/low/ncd[6] ), .f(\I0/low/U1664/U28/Z )
         );
    inv_1 \I0/low/U1664/U28/U30/Uinv  ( .x(\I0/low/U1664/U28/Z ), .a(
        \I0/low/U1664/x[3] ) );
    aoi222_1 \I0/low/U1664/U32/U30/U1  ( .x(\I0/low/U1664/x[0] ), .a(
        \I0/low/ncd[1] ), .b(\I0/low/ncd[0] ), .c(\I0/low/ncd[1] ), .d(
        \I0/low/U1664/U32/Z ), .e(\I0/low/ncd[0] ), .f(\I0/low/U1664/U32/Z )
         );
    inv_1 \I0/low/U1664/U32/U30/Uinv  ( .x(\I0/low/U1664/U32/Z ), .a(
        \I0/low/U1664/x[0] ) );
    aoi222_1 \I0/low/U1664/U29/U30/U1  ( .x(\I0/low/U1664/x[2] ), .a(
        \I0/low/ncd[5] ), .b(\I0/low/ncd[4] ), .c(\I0/low/ncd[5] ), .d(
        \I0/low/U1664/U29/Z ), .e(\I0/low/ncd[4] ), .f(\I0/low/U1664/U29/Z )
         );
    inv_1 \I0/low/U1664/U29/U30/Uinv  ( .x(\I0/low/U1664/U29/Z ), .a(
        \I0/low/U1664/x[2] ) );
    aoi222_1 \I0/low/U1664/U33/U30/U1  ( .x(\I0/low/U1664/y[0] ), .a(
        \I0/low/U1664/x[1] ), .b(\I0/low/U1664/x[0] ), .c(\I0/low/U1664/x[1] ), 
        .d(\I0/low/U1664/U33/Z ), .e(\I0/low/U1664/x[0] ), .f(
        \I0/low/U1664/U33/Z ) );
    inv_1 \I0/low/U1664/U33/U30/Uinv  ( .x(\I0/low/U1664/U33/Z ), .a(
        \I0/low/U1664/y[0] ) );
    aoi222_1 \I0/low/U1664/U30/U30/U1  ( .x(\I0/low/U1664/y[1] ), .a(
        \I0/low/U1664/x[3] ), .b(\I0/low/U1664/x[2] ), .c(\I0/low/U1664/x[3] ), 
        .d(\I0/low/U1664/U30/Z ), .e(\I0/low/U1664/x[2] ), .f(
        \I0/low/U1664/U30/Z ) );
    inv_1 \I0/low/U1664/U30/U30/Uinv  ( .x(\I0/low/U1664/U30/Z ), .a(
        \I0/low/U1664/y[1] ) );
    aoi222_1 \I0/low/U1664/U31/U30/U1  ( .x(\I0/low/U1664/x[1] ), .a(
        \I0/low/ncd[3] ), .b(\I0/low/ncd[2] ), .c(\I0/low/ncd[3] ), .d(
        \I0/low/U1664/U31/Z ), .e(\I0/low/ncd[2] ), .f(\I0/low/U1664/U31/Z )
         );
    inv_1 \I0/low/U1664/U31/U30/Uinv  ( .x(\I0/low/U1664/U31/Z ), .a(
        \I0/low/U1664/x[1] ) );
    aoi222_1 \I0/low/U1664/U37/U30/U1  ( .x(\I0/low/localcd ), .a(
        \I0/low/U1664/y[0] ), .b(\I0/low/U1664/y[1] ), .c(\I0/low/U1664/y[0] ), 
        .d(\I0/low/U1664/U37/Z ), .e(\I0/low/U1664/y[1] ), .f(
        \I0/low/U1664/U37/Z ) );
    inv_1 \I0/low/U1664/U37/U30/Uinv  ( .x(\I0/low/U1664/U37/Z ), .a(
        \I0/low/localcd ) );
    nor3_1 \I0/low/U1669/Unr  ( .x(\I0/low/U1669/nr ), .a(
        \I0/low/ctrlack_internal ), .b(n1), .c(\I0/low/driveh ) );
    nand3_1 \I0/low/U1669/Und  ( .x(\I0/low/U1669/nd ), .a(
        \I0/low/ctrlack_internal ), .b(\I0/low/drivel ), .c(\I0/low/driveh )
         );
    oa21_1 \I0/low/U1669/U1  ( .x(\I0/low/U1669/n2 ), .a(\I0/low/U1669/n2 ), 
        .b(\I0/low/U1669/nr ), .c(\I0/low/U1669/nd ) );
    inv_2 \I0/low/U1669/U3  ( .x(ctrlack), .a(\I0/low/U1669/n2 ) );
    buf_2 \I0/high/U1653  ( .x(\I0/high/latch ), .a(\I0/net33 ) );
    nor2_1 \I0/high/U264/U5  ( .x(\I0/high/nlocalcd ), .a(reset), .b(
        \I0/high/localcd ) );
    nor2_1 \I0/high/U1659_0_/U5  ( .x(\I0/high/ncd[0] ), .a(ol[8]), .b(oh[8])
         );
    nor2_1 \I0/high/U1659_1_/U5  ( .x(\I0/high/ncd[1] ), .a(ol[9]), .b(oh[9])
         );
    nor2_1 \I0/high/U1659_2_/U5  ( .x(\I0/high/ncd[2] ), .a(ol[10]), .b(oh[10]
        ) );
    nor2_1 \I0/high/U1659_3_/U5  ( .x(\I0/high/ncd[3] ), .a(ol[11]), .b(oh[11]
        ) );
    nor2_1 \I0/high/U1659_4_/U5  ( .x(\I0/high/ncd[4] ), .a(ol[12]), .b(oh[12]
        ) );
    nor2_1 \I0/high/U1659_5_/U5  ( .x(\I0/high/ncd[5] ), .a(ol[13]), .b(oh[13]
        ) );
    nor2_1 \I0/high/U1659_6_/U5  ( .x(\I0/high/ncd[6] ), .a(ol[14]), .b(oh[14]
        ) );
    nor2_1 \I0/high/U1659_7_/U5  ( .x(\I0/high/ncd[7] ), .a(ol[15]), .b(oh[15]
        ) );
    nor2_1 \I0/high/U3/U5  ( .x(\I0/high/ctrlack_internal ), .a(\I0/high/acb ), 
        .b(\I0/high/ba ) );
    buf_2 \I0/high/U1665/U7  ( .x(\I0/high/driveh ), .a(net17) );
    buf_2 \I0/high/U1666/U7  ( .x(\I0/high/drivel ), .a(net17) );
    ao23_1 \I0/high/U1658_0_/U21/U1/U1  ( .x(ol[8]), .a(\I0/high/driveh ), .b(
        ol[8]), .c(n3), .d(pull_l[0]), .e(n4) );
    ao23_1 \I0/high/U1658_1_/U21/U1/U1  ( .x(ol[9]), .a(\I0/high/drivel ), .b(
        ol[9]), .c(\I0/high/driveh ), .d(pull_l[1]), .e(n4) );
    ao23_1 \I0/high/U1658_2_/U21/U1/U1  ( .x(ol[10]), .a(\I0/high/drivel ), 
        .b(ol[10]), .c(\I0/high/driveh ), .d(pull_l[2]), .e(n4) );
    ao23_1 \I0/high/U1658_3_/U21/U1/U1  ( .x(ol[11]), .a(\I0/high/driveh ), 
        .b(ol[11]), .c(\I0/high/drivel ), .d(pull_l[3]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1658_4_/U21/U1/U1  ( .x(ol[12]), .a(n3), .b(ol[12]), .c(
        \I0/high/drivel ), .d(pull_l[4]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1658_5_/U21/U1/U1  ( .x(ol[13]), .a(\I0/high/driveh ), 
        .b(ol[13]), .c(n3), .d(pull_l[5]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1658_6_/U21/U1/U1  ( .x(ol[14]), .a(\I0/high/drivel ), 
        .b(ol[14]), .c(\I0/high/driveh ), .d(pull_l[6]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1658_7_/U21/U1/U1  ( .x(ol[15]), .a(n3), .b(ol[15]), .c(
        n3), .d(pull_l[7]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_0_/U21/U1/U1  ( .x(oh[8]), .a(\I0/high/driveh ), .b(
        oh[8]), .c(n3), .d(pull_h[0]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_1_/U21/U1/U1  ( .x(oh[9]), .a(n3), .b(oh[9]), .c(
        \I0/high/drivel ), .d(pull_h[1]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_2_/U21/U1/U1  ( .x(oh[10]), .a(\I0/high/drivel ), 
        .b(oh[10]), .c(\I0/high/drivel ), .d(pull_h[2]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1651_3_/U21/U1/U1  ( .x(oh[11]), .a(n3), .b(oh[11]), .c(
        \I0/high/driveh ), .d(pull_h[3]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_4_/U21/U1/U1  ( .x(oh[12]), .a(n3), .b(oh[12]), .c(
        n3), .d(pull_h[4]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_5_/U21/U1/U1  ( .x(oh[13]), .a(\I0/high/drivel ), 
        .b(oh[13]), .c(n3), .d(pull_h[5]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_6_/U21/U1/U1  ( .x(oh[14]), .a(\I0/high/drivel ), 
        .b(oh[14]), .c(\I0/high/driveh ), .d(pull_h[6]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1651_7_/U21/U1/U1  ( .x(oh[15]), .a(\I0/high/driveh ), 
        .b(oh[15]), .c(\I0/high/drivel ), .d(pull_h[7]), .e(\I0/high/latch )
         );
    aoai211_1 \I0/high/U4/U28/U1/U1  ( .x(\I0/high/U4/U28/U1/clr ), .a(net17), 
        .b(\I0/high/acb ), .c(\I0/high/nlocalcd ), .d(\I0/net33 ) );
    nand3_1 \I0/high/U4/U28/U1/U2  ( .x(\I0/high/U4/U28/U1/set ), .a(
        \I0/high/nlocalcd ), .b(net17), .c(\I0/high/acb ) );
    nand2_2 \I0/high/U4/U28/U1/U3  ( .x(\I0/net33 ), .a(
        \I0/high/U4/U28/U1/clr ), .b(\I0/high/U4/U28/U1/set ) );
    oai21_1 \I0/high/U1/U30/U1/U1  ( .x(\I0/high/acb ), .a(\I0/high/U1/Z ), 
        .b(\I0/high/ba ), .c(net17) );
    inv_1 \I0/high/U1/U30/U1/U2  ( .x(\I0/high/U1/Z ), .a(\I0/high/acb ) );
    ao222_1 \I0/high/U5/U18/U1/U1  ( .x(\I0/high/ba ), .a(\I0/high/latch ), 
        .b(pullcd), .c(\I0/high/latch ), .d(\I0/high/ba ), .e(pullcd), .f(
        \I0/high/ba ) );
    aoi222_1 \I0/high/U1664/U28/U30/U1  ( .x(\I0/high/U1664/x[3] ), .a(
        \I0/high/ncd[7] ), .b(\I0/high/ncd[6] ), .c(\I0/high/ncd[7] ), .d(
        \I0/high/U1664/U28/Z ), .e(\I0/high/ncd[6] ), .f(\I0/high/U1664/U28/Z 
        ) );
    inv_1 \I0/high/U1664/U28/U30/Uinv  ( .x(\I0/high/U1664/U28/Z ), .a(
        \I0/high/U1664/x[3] ) );
    aoi222_1 \I0/high/U1664/U32/U30/U1  ( .x(\I0/high/U1664/x[0] ), .a(
        \I0/high/ncd[1] ), .b(\I0/high/ncd[0] ), .c(\I0/high/ncd[1] ), .d(
        \I0/high/U1664/U32/Z ), .e(\I0/high/ncd[0] ), .f(\I0/high/U1664/U32/Z 
        ) );
    inv_1 \I0/high/U1664/U32/U30/Uinv  ( .x(\I0/high/U1664/U32/Z ), .a(
        \I0/high/U1664/x[0] ) );
    aoi222_1 \I0/high/U1664/U29/U30/U1  ( .x(\I0/high/U1664/x[2] ), .a(
        \I0/high/ncd[5] ), .b(\I0/high/ncd[4] ), .c(\I0/high/ncd[5] ), .d(
        \I0/high/U1664/U29/Z ), .e(\I0/high/ncd[4] ), .f(\I0/high/U1664/U29/Z 
        ) );
    inv_1 \I0/high/U1664/U29/U30/Uinv  ( .x(\I0/high/U1664/U29/Z ), .a(
        \I0/high/U1664/x[2] ) );
    aoi222_1 \I0/high/U1664/U33/U30/U1  ( .x(\I0/high/U1664/y[0] ), .a(
        \I0/high/U1664/x[1] ), .b(\I0/high/U1664/x[0] ), .c(
        \I0/high/U1664/x[1] ), .d(\I0/high/U1664/U33/Z ), .e(
        \I0/high/U1664/x[0] ), .f(\I0/high/U1664/U33/Z ) );
    inv_1 \I0/high/U1664/U33/U30/Uinv  ( .x(\I0/high/U1664/U33/Z ), .a(
        \I0/high/U1664/y[0] ) );
    aoi222_1 \I0/high/U1664/U30/U30/U1  ( .x(\I0/high/U1664/y[1] ), .a(
        \I0/high/U1664/x[3] ), .b(\I0/high/U1664/x[2] ), .c(
        \I0/high/U1664/x[3] ), .d(\I0/high/U1664/U30/Z ), .e(
        \I0/high/U1664/x[2] ), .f(\I0/high/U1664/U30/Z ) );
    inv_1 \I0/high/U1664/U30/U30/Uinv  ( .x(\I0/high/U1664/U30/Z ), .a(
        \I0/high/U1664/y[1] ) );
    aoi222_1 \I0/high/U1664/U31/U30/U1  ( .x(\I0/high/U1664/x[1] ), .a(
        \I0/high/ncd[3] ), .b(\I0/high/ncd[2] ), .c(\I0/high/ncd[3] ), .d(
        \I0/high/U1664/U31/Z ), .e(\I0/high/ncd[2] ), .f(\I0/high/U1664/U31/Z 
        ) );
    inv_1 \I0/high/U1664/U31/U30/Uinv  ( .x(\I0/high/U1664/U31/Z ), .a(
        \I0/high/U1664/x[1] ) );
    aoi222_1 \I0/high/U1664/U37/U30/U1  ( .x(\I0/high/localcd ), .a(
        \I0/high/U1664/y[0] ), .b(\I0/high/U1664/y[1] ), .c(
        \I0/high/U1664/y[0] ), .d(\I0/high/U1664/U37/Z ), .e(
        \I0/high/U1664/y[1] ), .f(\I0/high/U1664/U37/Z ) );
    inv_1 \I0/high/U1664/U37/U30/Uinv  ( .x(\I0/high/U1664/U37/Z ), .a(
        \I0/high/localcd ) );
    nor3_1 \I0/high/U1669/Unr  ( .x(\I0/high/U1669/nr ), .a(
        \I0/high/ctrlack_internal ), .b(n3), .c(\I0/high/driveh ) );
    nand3_1 \I0/high/U1669/Und  ( .x(\I0/high/U1669/nd ), .a(
        \I0/high/ctrlack_internal ), .b(\I0/high/drivel ), .c(\I0/high/driveh 
        ) );
    oa21_1 \I0/high/U1669/U1  ( .x(\I0/high/U1669/n2 ), .a(\I0/high/U1669/n2 ), 
        .b(\I0/high/U1669/nr ), .c(\I0/high/U1669/nd ) );
    inv_2 \I0/high/U1669/U3  ( .x(\I0/net20 ), .a(\I0/high/U1669/n2 ) );
    nor2_1 \I1/U3/U5  ( .x(net31), .a(\I1/net32 ), .b(\I1/net33 ) );
    buf_2 \I1/low/U1653  ( .x(\I1/low/latch ), .a(\I1/net32 ) );
    nor2_1 \I1/low/U264/U5  ( .x(\I1/low/nlocalcd ), .a(reset), .b(
        \I1/low/localcd ) );
    nor2_1 \I1/low/U1659_0_/U5  ( .x(\I1/low/ncd[0] ), .a(ol[16]), .b(oh[16])
         );
    nor2_1 \I1/low/U1659_1_/U5  ( .x(\I1/low/ncd[1] ), .a(ol[17]), .b(oh[17])
         );
    nor2_1 \I1/low/U1659_2_/U5  ( .x(\I1/low/ncd[2] ), .a(ol[18]), .b(oh[18])
         );
    nor2_1 \I1/low/U1659_3_/U5  ( .x(\I1/low/ncd[3] ), .a(ol[19]), .b(oh[19])
         );
    nor2_1 \I1/low/U1659_4_/U5  ( .x(\I1/low/ncd[4] ), .a(ol[20]), .b(oh[20])
         );
    nor2_1 \I1/low/U1659_5_/U5  ( .x(\I1/low/ncd[5] ), .a(ol[21]), .b(oh[21])
         );
    nor2_1 \I1/low/U1659_6_/U5  ( .x(\I1/low/ncd[6] ), .a(ol[22]), .b(oh[22])
         );
    nor2_1 \I1/low/U1659_7_/U5  ( .x(\I1/low/ncd[7] ), .a(ol[23]), .b(oh[23])
         );
    nor2_1 \I1/low/U3/U5  ( .x(\I1/low/ctrlack_internal ), .a(\I1/low/acb ), 
        .b(\I1/low/ba ) );
    buf_2 \I1/low/U1665/U7  ( .x(\I1/low/driveh ), .a(\I1/net20 ) );
    buf_2 \I1/low/U1666/U7  ( .x(\I1/low/drivel ), .a(\I1/net20 ) );
    ao23_1 \I1/low/U1658_0_/U21/U1/U1  ( .x(ol[16]), .a(\I1/low/driveh ), .b(
        ol[16]), .c(n5), .d(pull_l[0]), .e(n6) );
    ao23_1 \I1/low/U1658_1_/U21/U1/U1  ( .x(ol[17]), .a(\I1/low/drivel ), .b(
        ol[17]), .c(\I1/low/driveh ), .d(pull_l[1]), .e(n6) );
    ao23_1 \I1/low/U1658_2_/U21/U1/U1  ( .x(ol[18]), .a(\I1/low/drivel ), .b(
        ol[18]), .c(\I1/low/driveh ), .d(pull_l[2]), .e(n6) );
    ao23_1 \I1/low/U1658_3_/U21/U1/U1  ( .x(ol[19]), .a(\I1/low/driveh ), .b(
        ol[19]), .c(\I1/low/drivel ), .d(pull_l[3]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_4_/U21/U1/U1  ( .x(ol[20]), .a(n5), .b(ol[20]), .c(
        \I1/low/drivel ), .d(pull_l[4]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_5_/U21/U1/U1  ( .x(ol[21]), .a(\I1/low/driveh ), .b(
        ol[21]), .c(n5), .d(pull_l[5]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_6_/U21/U1/U1  ( .x(ol[22]), .a(\I1/low/drivel ), .b(
        ol[22]), .c(\I1/low/driveh ), .d(pull_l[6]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_7_/U21/U1/U1  ( .x(ol[23]), .a(n5), .b(ol[23]), .c(n5
        ), .d(pull_l[7]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_0_/U21/U1/U1  ( .x(oh[16]), .a(\I1/low/driveh ), .b(
        oh[16]), .c(n5), .d(pull_h[0]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_1_/U21/U1/U1  ( .x(oh[17]), .a(n5), .b(oh[17]), .c(
        \I1/low/drivel ), .d(pull_h[1]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_2_/U21/U1/U1  ( .x(oh[18]), .a(\I1/low/drivel ), .b(
        oh[18]), .c(\I1/low/drivel ), .d(pull_h[2]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_3_/U21/U1/U1  ( .x(oh[19]), .a(n5), .b(oh[19]), .c(
        \I1/low/driveh ), .d(pull_h[3]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_4_/U21/U1/U1  ( .x(oh[20]), .a(n5), .b(oh[20]), .c(n5
        ), .d(pull_h[4]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_5_/U21/U1/U1  ( .x(oh[21]), .a(\I1/low/drivel ), .b(
        oh[21]), .c(n5), .d(pull_h[5]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_6_/U21/U1/U1  ( .x(oh[22]), .a(\I1/low/drivel ), .b(
        oh[22]), .c(\I1/low/driveh ), .d(pull_h[6]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_7_/U21/U1/U1  ( .x(oh[23]), .a(\I1/low/driveh ), .b(
        oh[23]), .c(\I1/low/drivel ), .d(pull_h[7]), .e(\I1/low/latch ) );
    aoai211_1 \I1/low/U4/U28/U1/U1  ( .x(\I1/low/U4/U28/U1/clr ), .a(
        \I1/net20 ), .b(\I1/low/acb ), .c(\I1/low/nlocalcd ), .d(\I1/net32 )
         );
    nand3_1 \I1/low/U4/U28/U1/U2  ( .x(\I1/low/U4/U28/U1/set ), .a(
        \I1/low/nlocalcd ), .b(\I1/net20 ), .c(\I1/low/acb ) );
    nand2_2 \I1/low/U4/U28/U1/U3  ( .x(\I1/net32 ), .a(\I1/low/U4/U28/U1/clr ), 
        .b(\I1/low/U4/U28/U1/set ) );
    oai21_1 \I1/low/U1/U30/U1/U1  ( .x(\I1/low/acb ), .a(\I1/low/U1/Z ), .b(
        \I1/low/ba ), .c(\I1/net20 ) );
    inv_1 \I1/low/U1/U30/U1/U2  ( .x(\I1/low/U1/Z ), .a(\I1/low/acb ) );
    ao222_1 \I1/low/U5/U18/U1/U1  ( .x(\I1/low/ba ), .a(\I1/low/latch ), .b(
        pullcd), .c(\I1/low/latch ), .d(\I1/low/ba ), .e(pullcd), .f(
        \I1/low/ba ) );
    aoi222_1 \I1/low/U1664/U28/U30/U1  ( .x(\I1/low/U1664/x[3] ), .a(
        \I1/low/ncd[7] ), .b(\I1/low/ncd[6] ), .c(\I1/low/ncd[7] ), .d(
        \I1/low/U1664/U28/Z ), .e(\I1/low/ncd[6] ), .f(\I1/low/U1664/U28/Z )
         );
    inv_1 \I1/low/U1664/U28/U30/Uinv  ( .x(\I1/low/U1664/U28/Z ), .a(
        \I1/low/U1664/x[3] ) );
    aoi222_1 \I1/low/U1664/U32/U30/U1  ( .x(\I1/low/U1664/x[0] ), .a(
        \I1/low/ncd[1] ), .b(\I1/low/ncd[0] ), .c(\I1/low/ncd[1] ), .d(
        \I1/low/U1664/U32/Z ), .e(\I1/low/ncd[0] ), .f(\I1/low/U1664/U32/Z )
         );
    inv_1 \I1/low/U1664/U32/U30/Uinv  ( .x(\I1/low/U1664/U32/Z ), .a(
        \I1/low/U1664/x[0] ) );
    aoi222_1 \I1/low/U1664/U29/U30/U1  ( .x(\I1/low/U1664/x[2] ), .a(
        \I1/low/ncd[5] ), .b(\I1/low/ncd[4] ), .c(\I1/low/ncd[5] ), .d(
        \I1/low/U1664/U29/Z ), .e(\I1/low/ncd[4] ), .f(\I1/low/U1664/U29/Z )
         );
    inv_1 \I1/low/U1664/U29/U30/Uinv  ( .x(\I1/low/U1664/U29/Z ), .a(
        \I1/low/U1664/x[2] ) );
    aoi222_1 \I1/low/U1664/U33/U30/U1  ( .x(\I1/low/U1664/y[0] ), .a(
        \I1/low/U1664/x[1] ), .b(\I1/low/U1664/x[0] ), .c(\I1/low/U1664/x[1] ), 
        .d(\I1/low/U1664/U33/Z ), .e(\I1/low/U1664/x[0] ), .f(
        \I1/low/U1664/U33/Z ) );
    inv_1 \I1/low/U1664/U33/U30/Uinv  ( .x(\I1/low/U1664/U33/Z ), .a(
        \I1/low/U1664/y[0] ) );
    aoi222_1 \I1/low/U1664/U30/U30/U1  ( .x(\I1/low/U1664/y[1] ), .a(
        \I1/low/U1664/x[3] ), .b(\I1/low/U1664/x[2] ), .c(\I1/low/U1664/x[3] ), 
        .d(\I1/low/U1664/U30/Z ), .e(\I1/low/U1664/x[2] ), .f(
        \I1/low/U1664/U30/Z ) );
    inv_1 \I1/low/U1664/U30/U30/Uinv  ( .x(\I1/low/U1664/U30/Z ), .a(
        \I1/low/U1664/y[1] ) );
    aoi222_1 \I1/low/U1664/U31/U30/U1  ( .x(\I1/low/U1664/x[1] ), .a(
        \I1/low/ncd[3] ), .b(\I1/low/ncd[2] ), .c(\I1/low/ncd[3] ), .d(
        \I1/low/U1664/U31/Z ), .e(\I1/low/ncd[2] ), .f(\I1/low/U1664/U31/Z )
         );
    inv_1 \I1/low/U1664/U31/U30/Uinv  ( .x(\I1/low/U1664/U31/Z ), .a(
        \I1/low/U1664/x[1] ) );
    aoi222_1 \I1/low/U1664/U37/U30/U1  ( .x(\I1/low/localcd ), .a(
        \I1/low/U1664/y[0] ), .b(\I1/low/U1664/y[1] ), .c(\I1/low/U1664/y[0] ), 
        .d(\I1/low/U1664/U37/Z ), .e(\I1/low/U1664/y[1] ), .f(
        \I1/low/U1664/U37/Z ) );
    inv_1 \I1/low/U1664/U37/U30/Uinv  ( .x(\I1/low/U1664/U37/Z ), .a(
        \I1/low/localcd ) );
    nor3_1 \I1/low/U1669/Unr  ( .x(\I1/low/U1669/nr ), .a(
        \I1/low/ctrlack_internal ), .b(n5), .c(\I1/low/driveh ) );
    nand3_1 \I1/low/U1669/Und  ( .x(\I1/low/U1669/nd ), .a(
        \I1/low/ctrlack_internal ), .b(\I1/low/drivel ), .c(\I1/low/driveh )
         );
    oa21_1 \I1/low/U1669/U1  ( .x(\I1/low/U1669/n2 ), .a(\I1/low/U1669/n2 ), 
        .b(\I1/low/U1669/nr ), .c(\I1/low/U1669/nd ) );
    inv_2 \I1/low/U1669/U3  ( .x(net17), .a(\I1/low/U1669/n2 ) );
    buf_2 \I1/high/U1653  ( .x(\I1/high/latch ), .a(\I1/net33 ) );
    nor2_1 \I1/high/U264/U5  ( .x(\I1/high/nlocalcd ), .a(reset), .b(
        \I1/high/localcd ) );
    nor2_1 \I1/high/U1659_0_/U5  ( .x(\I1/high/ncd[0] ), .a(ol[24]), .b(oh[24]
        ) );
    nor2_1 \I1/high/U1659_1_/U5  ( .x(\I1/high/ncd[1] ), .a(ol[25]), .b(oh[25]
        ) );
    nor2_1 \I1/high/U1659_2_/U5  ( .x(\I1/high/ncd[2] ), .a(ol[26]), .b(oh[26]
        ) );
    nor2_1 \I1/high/U1659_3_/U5  ( .x(\I1/high/ncd[3] ), .a(ol[27]), .b(oh[27]
        ) );
    nor2_1 \I1/high/U1659_4_/U5  ( .x(\I1/high/ncd[4] ), .a(ol[28]), .b(oh[28]
        ) );
    nor2_1 \I1/high/U1659_5_/U5  ( .x(\I1/high/ncd[5] ), .a(ol[29]), .b(oh[29]
        ) );
    nor2_1 \I1/high/U1659_6_/U5  ( .x(\I1/high/ncd[6] ), .a(ol[30]), .b(oh[30]
        ) );
    nor2_1 \I1/high/U1659_7_/U5  ( .x(\I1/high/ncd[7] ), .a(ol[31]), .b(oh[31]
        ) );
    nor2_1 \I1/high/U3/U5  ( .x(\I1/high/ctrlack_internal ), .a(\I1/high/acb ), 
        .b(\I1/high/ba ) );
    buf_2 \I1/high/U1665/U7  ( .x(\I1/high/driveh ), .a(ctrlreq) );
    buf_2 \I1/high/U1666/U7  ( .x(\I1/high/drivel ), .a(ctrlreq) );
    ao23_1 \I1/high/U1658_0_/U21/U1/U1  ( .x(ol[24]), .a(\I1/high/driveh ), 
        .b(ol[24]), .c(n7), .d(pull_l[0]), .e(n8) );
    ao23_1 \I1/high/U1658_1_/U21/U1/U1  ( .x(ol[25]), .a(\I1/high/drivel ), 
        .b(ol[25]), .c(\I1/high/driveh ), .d(pull_l[1]), .e(n8) );
    ao23_1 \I1/high/U1658_2_/U21/U1/U1  ( .x(ol[26]), .a(\I1/high/drivel ), 
        .b(ol[26]), .c(\I1/high/driveh ), .d(pull_l[2]), .e(n8) );
    ao23_1 \I1/high/U1658_3_/U21/U1/U1  ( .x(ol[27]), .a(\I1/high/driveh ), 
        .b(ol[27]), .c(\I1/high/drivel ), .d(pull_l[3]), .e(\I1/high/latch )
         );
    ao23_1 \I1/high/U1658_4_/U21/U1/U1  ( .x(ol[28]), .a(n7), .b(ol[28]), .c(
        \I1/high/drivel ), .d(pull_l[4]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1658_5_/U21/U1/U1  ( .x(ol[29]), .a(\I1/high/driveh ), 
        .b(ol[29]), .c(n7), .d(pull_l[5]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1658_6_/U21/U1/U1  ( .x(ol[30]), .a(\I1/high/drivel ), 
        .b(ol[30]), .c(\I1/high/driveh ), .d(pull_l[6]), .e(\I1/high/latch )
         );
    ao23_1 \I1/high/U1658_7_/U21/U1/U1  ( .x(ol[31]), .a(n7), .b(ol[31]), .c(
        n7), .d(pull_l[7]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_0_/U21/U1/U1  ( .x(oh[24]), .a(\I1/high/driveh ), 
        .b(oh[24]), .c(n7), .d(pull_h[0]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_1_/U21/U1/U1  ( .x(oh[25]), .a(n7), .b(oh[25]), .c(
        \I1/high/drivel ), .d(pull_h[1]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_2_/U21/U1/U1  ( .x(oh[26]), .a(\I1/high/drivel ), 
        .b(oh[26]), .c(\I1/high/drivel ), .d(pull_h[2]), .e(\I1/high/latch )
         );
    ao23_1 \I1/high/U1651_3_/U21/U1/U1  ( .x(oh[27]), .a(n7), .b(oh[27]), .c(
        \I1/high/driveh ), .d(pull_h[3]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_4_/U21/U1/U1  ( .x(oh[28]), .a(n7), .b(oh[28]), .c(
        n7), .d(pull_h[4]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_5_/U21/U1/U1  ( .x(oh[29]), .a(\I1/high/drivel ), 
        .b(oh[29]), .c(n7), .d(pull_h[5]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_6_/U21/U1/U1  ( .x(oh[30]), .a(\I1/high/drivel ), 
        .b(oh[30]), .c(\I1/high/driveh ), .d(pull_h[6]), .e(\I1/high/latch )
         );
    ao23_1 \I1/high/U1651_7_/U21/U1/U1  ( .x(oh[31]), .a(\I1/high/driveh ), 
        .b(oh[31]), .c(\I1/high/drivel ), .d(pull_h[7]), .e(\I1/high/latch )
         );
    aoai211_1 \I1/high/U4/U28/U1/U1  ( .x(\I1/high/U4/U28/U1/clr ), .a(ctrlreq
        ), .b(\I1/high/acb ), .c(\I1/high/nlocalcd ), .d(\I1/net33 ) );
    nand3_1 \I1/high/U4/U28/U1/U2  ( .x(\I1/high/U4/U28/U1/set ), .a(
        \I1/high/nlocalcd ), .b(ctrlreq), .c(\I1/high/acb ) );
    nand2_2 \I1/high/U4/U28/U1/U3  ( .x(\I1/net33 ), .a(
        \I1/high/U4/U28/U1/clr ), .b(\I1/high/U4/U28/U1/set ) );
    oai21_1 \I1/high/U1/U30/U1/U1  ( .x(\I1/high/acb ), .a(\I1/high/U1/Z ), 
        .b(\I1/high/ba ), .c(ctrlreq) );
    inv_1 \I1/high/U1/U30/U1/U2  ( .x(\I1/high/U1/Z ), .a(\I1/high/acb ) );
    ao222_1 \I1/high/U5/U18/U1/U1  ( .x(\I1/high/ba ), .a(\I1/high/latch ), 
        .b(pullcd), .c(\I1/high/latch ), .d(\I1/high/ba ), .e(pullcd), .f(
        \I1/high/ba ) );
    aoi222_1 \I1/high/U1664/U28/U30/U1  ( .x(\I1/high/U1664/x[3] ), .a(
        \I1/high/ncd[7] ), .b(\I1/high/ncd[6] ), .c(\I1/high/ncd[7] ), .d(
        \I1/high/U1664/U28/Z ), .e(\I1/high/ncd[6] ), .f(\I1/high/U1664/U28/Z 
        ) );
    inv_1 \I1/high/U1664/U28/U30/Uinv  ( .x(\I1/high/U1664/U28/Z ), .a(
        \I1/high/U1664/x[3] ) );
    aoi222_1 \I1/high/U1664/U32/U30/U1  ( .x(\I1/high/U1664/x[0] ), .a(
        \I1/high/ncd[1] ), .b(\I1/high/ncd[0] ), .c(\I1/high/ncd[1] ), .d(
        \I1/high/U1664/U32/Z ), .e(\I1/high/ncd[0] ), .f(\I1/high/U1664/U32/Z 
        ) );
    inv_1 \I1/high/U1664/U32/U30/Uinv  ( .x(\I1/high/U1664/U32/Z ), .a(
        \I1/high/U1664/x[0] ) );
    aoi222_1 \I1/high/U1664/U29/U30/U1  ( .x(\I1/high/U1664/x[2] ), .a(
        \I1/high/ncd[5] ), .b(\I1/high/ncd[4] ), .c(\I1/high/ncd[5] ), .d(
        \I1/high/U1664/U29/Z ), .e(\I1/high/ncd[4] ), .f(\I1/high/U1664/U29/Z 
        ) );
    inv_1 \I1/high/U1664/U29/U30/Uinv  ( .x(\I1/high/U1664/U29/Z ), .a(
        \I1/high/U1664/x[2] ) );
    aoi222_1 \I1/high/U1664/U33/U30/U1  ( .x(\I1/high/U1664/y[0] ), .a(
        \I1/high/U1664/x[1] ), .b(\I1/high/U1664/x[0] ), .c(
        \I1/high/U1664/x[1] ), .d(\I1/high/U1664/U33/Z ), .e(
        \I1/high/U1664/x[0] ), .f(\I1/high/U1664/U33/Z ) );
    inv_1 \I1/high/U1664/U33/U30/Uinv  ( .x(\I1/high/U1664/U33/Z ), .a(
        \I1/high/U1664/y[0] ) );
    aoi222_1 \I1/high/U1664/U30/U30/U1  ( .x(\I1/high/U1664/y[1] ), .a(
        \I1/high/U1664/x[3] ), .b(\I1/high/U1664/x[2] ), .c(
        \I1/high/U1664/x[3] ), .d(\I1/high/U1664/U30/Z ), .e(
        \I1/high/U1664/x[2] ), .f(\I1/high/U1664/U30/Z ) );
    inv_1 \I1/high/U1664/U30/U30/Uinv  ( .x(\I1/high/U1664/U30/Z ), .a(
        \I1/high/U1664/y[1] ) );
    aoi222_1 \I1/high/U1664/U31/U30/U1  ( .x(\I1/high/U1664/x[1] ), .a(
        \I1/high/ncd[3] ), .b(\I1/high/ncd[2] ), .c(\I1/high/ncd[3] ), .d(
        \I1/high/U1664/U31/Z ), .e(\I1/high/ncd[2] ), .f(\I1/high/U1664/U31/Z 
        ) );
    inv_1 \I1/high/U1664/U31/U30/Uinv  ( .x(\I1/high/U1664/U31/Z ), .a(
        \I1/high/U1664/x[1] ) );
    aoi222_1 \I1/high/U1664/U37/U30/U1  ( .x(\I1/high/localcd ), .a(
        \I1/high/U1664/y[0] ), .b(\I1/high/U1664/y[1] ), .c(
        \I1/high/U1664/y[0] ), .d(\I1/high/U1664/U37/Z ), .e(
        \I1/high/U1664/y[1] ), .f(\I1/high/U1664/U37/Z ) );
    inv_1 \I1/high/U1664/U37/U30/Uinv  ( .x(\I1/high/U1664/U37/Z ), .a(
        \I1/high/localcd ) );
    nor3_1 \I1/high/U1669/Unr  ( .x(\I1/high/U1669/nr ), .a(
        \I1/high/ctrlack_internal ), .b(n7), .c(\I1/high/driveh ) );
    nand3_1 \I1/high/U1669/Und  ( .x(\I1/high/U1669/nd ), .a(
        \I1/high/ctrlack_internal ), .b(\I1/high/drivel ), .c(\I1/high/driveh 
        ) );
    oa21_1 \I1/high/U1669/U1  ( .x(\I1/high/U1669/n2 ), .a(\I1/high/U1669/n2 ), 
        .b(\I1/high/U1669/nr ), .c(\I1/high/U1669/nd ) );
    inv_2 \I1/high/U1669/U3  ( .x(\I1/net20 ), .a(\I1/high/U1669/n2 ) );
    buf_2 U1 ( .x(n1), .a(\I0/net20 ) );
    buf_1 U2 ( .x(n2), .a(\I0/low/latch ) );
    buf_2 U3 ( .x(n3), .a(net17) );
    buf_1 U4 ( .x(n4), .a(\I0/high/latch ) );
    buf_2 U5 ( .x(n5), .a(\I1/net20 ) );
    buf_1 U6 ( .x(n6), .a(\I1/low/latch ) );
    buf_2 U7 ( .x(n7), .a(ctrlreq) );
    buf_1 U8 ( .x(n8), .a(\I1/high/latch ) );
endmodule


module chain_fr2dr_byte_2 ( nia, oh, ol, i, nReset, noa );
output [7:0] oh;
output [7:0] ol;
input  [4:0] i;
input  nReset, noa;
output nia;
    wire nbReset, eop, ncla, csela, asela, \U891/reset , \U891/neopack , 
        \U891/iay , \U891/naack[0] , \U891/naack[1] , \U891/U1128/nb , \b[3] , 
        \b[2] , \U891/U1128/na , \b[1] , \b[0] , \U891/ackb , \a[3] , \a[2] , 
        \U891/nack , \U891/acka , \a[1] , \a[0] , bsela, bsel, asel, 
        \U891/U1118_0_/nr , naa, \U891/U1118_0_/nd , \U891/U1118_0_/n2 , 
        \U891/U1118_1_/nr , \U891/U1118_1_/nd , \U891/U1118_1_/n2 , 
        \U891/U1118_2_/nr , \U891/U1118_2_/nd , \U891/U1118_2_/n2 , 
        \U891/U1118_3_/nr , \U891/U1118_3_/nd , \U891/U1118_3_/n2 , 
        \U891/U1117_0_/nr , nba, \U891/U1117_0_/nd , \U891/U1117_0_/n2 , 
        \U891/U1117_1_/nr , \U891/U1117_1_/nd , \U891/U1117_1_/n2 , 
        \U891/U1117_2_/nr , \U891/U1117_2_/nd , \U891/U1117_2_/n2 , 
        \U891/U1117_3_/nr , \U891/U1117_3_/nd , \U891/U1117_3_/n2 , 
        \U886/reset , \U886/U1128/nb , \f[3] , \f[2] , \U886/U1128/na , \f[1] , 
        \f[0] , \U886/ackb , \U886/nack , \U886/acka , \U886/U1127/n5 , 
        \U886/U1127/n1 , \U886/U1127/n2 , \U886/U1127/n3 , \U886/U1127/n4 , 
        \e[3] , \e[2] , \e[1] , \e[0] , fsela, fsel, esela, esel, 
        \U886/U1118_0_/nr , nea, \U886/U1118_0_/nd , \U886/U1118_0_/n2 , 
        \U886/U1118_1_/nr , \U886/U1118_1_/nd , \U886/U1118_1_/n2 , 
        \U886/U1118_2_/nr , \U886/U1118_2_/nd , \U886/U1118_2_/n2 , 
        \U886/U1118_3_/nr , \U886/U1118_3_/nd , \U886/U1118_3_/n2 , 
        \U886/U1117_0_/nr , nfa, \U886/U1117_0_/nd , \U886/U1117_0_/n2 , 
        \U886/U1117_1_/nr , \U886/U1117_1_/nd , \U886/U1117_1_/n2 , 
        \U886/U1117_2_/nr , \U886/U1117_2_/nd , \U886/U1117_2_/n2 , 
        \U886/U1117_3_/nr , \U886/U1117_3_/nd , \U886/U1117_3_/n2 , 
        \U884/reset , \U884/U1128/nb , \d[3] , \d[2] , \U884/U1128/na , \d[1] , 
        \d[0] , \U884/ackb , \U884/nack , \U884/acka , \U884/U1127/n5 , 
        \U884/U1127/n1 , \U884/U1127/n2 , \U884/U1127/n3 , \U884/U1127/n4 , 
        \c[3] , \c[2] , \c[1] , \c[0] , dsela, dsel, csel, \U884/U1118_0_/nr , 
        nca, \U884/U1118_0_/nd , \U884/U1118_0_/n2 , \U884/U1118_1_/nr , 
        \U884/U1118_1_/nd , \U884/U1118_1_/n2 , \U884/U1118_2_/nr , 
        \U884/U1118_2_/nd , \U884/U1118_2_/n2 , \U884/U1118_3_/nr , 
        \U884/U1118_3_/nd , \U884/U1118_3_/n2 , \U884/U1117_0_/nr , nda, 
        \U884/U1117_0_/nd , \U884/U1117_0_/n2 , \U884/U1117_1_/nr , 
        \U884/U1117_1_/nd , \U884/U1117_1_/n2 , \U884/U1117_2_/nr , 
        \U884/U1117_2_/nd , \U884/U1117_2_/n2 , \U884/U1117_3_/nr , 
        \U884/U1117_3_/nd , \U884/U1117_3_/n2 , \U888/s , \U888/r , 
        \U888/nback , \U888/naack , \U888/reset , \U887/s , \U887/r , 
        \U887/nback , \U887/naack , \U887/reset , \U885/s , \U885/r , 
        \U885/nback , \U885/naack , \U885/reset , \U877/x , \U877/reset , 
        \U877/y , \U877/U590/U25/U1/clr , net135, \cl[3] , \cl[1] , 
        \U877/U590/U25/U1/ob , n1, \U877/U589/U25/U1/clr , \cl[0] , 
        \U877/U589/U25/U1/ob , \U877/U588/U25/U1/clr , \cl[2] , 
        \U877/U588/U25/U1/ob , \U877/U591/U25/U1/clr , \U877/U591/U25/U1/ob , 
        \U876/x , \U876/reset , \U876/y , \U876/U590/U25/U1/clr , 
        \U876/U590/U25/U1/ob , \U876/U589/U25/U1/clr , \U876/U589/U25/U1/ob , 
        \U876/U588/U25/U1/clr , \U876/U588/U25/U1/ob , \U876/U591/U25/U1/clr , 
        \U876/U591/U25/U1/ob , \U2/x , \U2/reset , \U2/y , 
        \U2/U590/U25/U1/clr , \U2/U590/U25/U1/ob , \U2/U589/U25/U1/clr , 
        \U2/U589/U25/U1/ob , \U2/U588/U25/U1/clr , \U2/U588/U25/U1/ob , 
        \U2/U591/U25/U1/clr , \U2/U591/U25/U1/ob , \U1/x , \U1/reset , \U1/y , 
        \U1/U590/U25/U1/clr , \U1/U590/U25/U1/ob , \U1/U589/U25/U1/clr , 
        \U1/U589/U25/U1/ob , \U1/U588/U25/U1/clr , \U1/U588/U25/U1/ob , 
        \U1/U591/U25/U1/clr , \U1/U591/U25/U1/ob , \U881/nack[1] , 
        \U881/nack[0] ;
    buf_2 U897 ( .x(nbReset), .a(nReset) );
    and4_1 \U894/U12  ( .x(eop), .a(ncla), .b(csela), .c(asela), .d(i[4]) );
    inv_1 \U891/U1126/U3  ( .x(\U891/reset ), .a(nbReset) );
    inv_1 \U891/U1139/U3  ( .x(\U891/neopack ), .a(eop) );
    nand3_1 \U891/U1131/U9  ( .x(\U891/iay ), .a(\U891/neopack ), .b(
        \U891/naack[0] ), .c(\U891/naack[1] ) );
    nor3_1 \U891/U1128/U27  ( .x(\U891/U1128/nb ), .a(\U891/reset ), .b(\b[3] 
        ), .c(\b[2] ) );
    nor2_1 \U891/U1128/U26  ( .x(\U891/U1128/na ), .a(\b[1] ), .b(\b[0] ) );
    nand2_2 \U891/U1128/U29  ( .x(\U891/ackb ), .a(\U891/U1128/nb ), .b(
        \U891/U1128/na ) );
    nor2_1 \U891/U1133/U5  ( .x(\U891/naack[0] ), .a(\a[3] ), .b(\a[2] ) );
    nor2_1 \U891/U1108/U5  ( .x(\U891/nack ), .a(\U891/acka ), .b(\U891/ackb )
         );
    nor2_1 \U891/U1134/U5  ( .x(\U891/naack[1] ), .a(\a[1] ), .b(\a[0] ) );
    nor2_2 \U891/U914/U6  ( .x(nia), .a(\U891/iay ), .b(\U891/ackb ) );
    nand2_1 \U891/U1130/U5  ( .x(\U891/acka ), .a(\U891/naack[0] ), .b(
        \U891/naack[1] ) );
    ao222_4 \U891/U1121/U1/U1  ( .x(bsela), .a(\U891/nack ), .b(bsel), .c(
        \U891/nack ), .d(bsela), .e(bsel), .f(bsela) );
    ao222_4 \U891/U1120/U1/U1  ( .x(asela), .a(asel), .b(\U891/nack ), .c(asel
        ), .d(asela), .e(\U891/nack ), .f(asela) );
    nor3_1 \U891/U1118_0_/Unr  ( .x(\U891/U1118_0_/nr ), .a(i[0]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_0_/Und  ( .x(\U891/U1118_0_/nd ), .a(i[0]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_0_/U1  ( .x(\U891/U1118_0_/n2 ), .a(\U891/U1118_0_/n2 ), 
        .b(\U891/U1118_0_/nr ), .c(\U891/U1118_0_/nd ) );
    inv_2 \U891/U1118_0_/U3  ( .x(\a[0] ), .a(\U891/U1118_0_/n2 ) );
    nor3_1 \U891/U1118_1_/Unr  ( .x(\U891/U1118_1_/nr ), .a(i[1]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_1_/Und  ( .x(\U891/U1118_1_/nd ), .a(i[1]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_1_/U1  ( .x(\U891/U1118_1_/n2 ), .a(\U891/U1118_1_/n2 ), 
        .b(\U891/U1118_1_/nr ), .c(\U891/U1118_1_/nd ) );
    inv_2 \U891/U1118_1_/U3  ( .x(\a[1] ), .a(\U891/U1118_1_/n2 ) );
    nor3_1 \U891/U1118_2_/Unr  ( .x(\U891/U1118_2_/nr ), .a(i[2]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_2_/Und  ( .x(\U891/U1118_2_/nd ), .a(i[2]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_2_/U1  ( .x(\U891/U1118_2_/n2 ), .a(\U891/U1118_2_/n2 ), 
        .b(\U891/U1118_2_/nr ), .c(\U891/U1118_2_/nd ) );
    inv_2 \U891/U1118_2_/U3  ( .x(\a[2] ), .a(\U891/U1118_2_/n2 ) );
    nor3_1 \U891/U1118_3_/Unr  ( .x(\U891/U1118_3_/nr ), .a(i[3]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_3_/Und  ( .x(\U891/U1118_3_/nd ), .a(i[3]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_3_/U1  ( .x(\U891/U1118_3_/n2 ), .a(\U891/U1118_3_/n2 ), 
        .b(\U891/U1118_3_/nr ), .c(\U891/U1118_3_/nd ) );
    inv_2 \U891/U1118_3_/U3  ( .x(\a[3] ), .a(\U891/U1118_3_/n2 ) );
    nor3_1 \U891/U1117_0_/Unr  ( .x(\U891/U1117_0_/nr ), .a(i[0]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_0_/Und  ( .x(\U891/U1117_0_/nd ), .a(i[0]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_0_/U1  ( .x(\U891/U1117_0_/n2 ), .a(\U891/U1117_0_/n2 ), 
        .b(\U891/U1117_0_/nr ), .c(\U891/U1117_0_/nd ) );
    inv_2 \U891/U1117_0_/U3  ( .x(\b[0] ), .a(\U891/U1117_0_/n2 ) );
    nor3_1 \U891/U1117_1_/Unr  ( .x(\U891/U1117_1_/nr ), .a(i[1]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_1_/Und  ( .x(\U891/U1117_1_/nd ), .a(i[1]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_1_/U1  ( .x(\U891/U1117_1_/n2 ), .a(\U891/U1117_1_/n2 ), 
        .b(\U891/U1117_1_/nr ), .c(\U891/U1117_1_/nd ) );
    inv_2 \U891/U1117_1_/U3  ( .x(\b[1] ), .a(\U891/U1117_1_/n2 ) );
    nor3_1 \U891/U1117_2_/Unr  ( .x(\U891/U1117_2_/nr ), .a(i[2]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_2_/Und  ( .x(\U891/U1117_2_/nd ), .a(i[2]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_2_/U1  ( .x(\U891/U1117_2_/n2 ), .a(\U891/U1117_2_/n2 ), 
        .b(\U891/U1117_2_/nr ), .c(\U891/U1117_2_/nd ) );
    inv_2 \U891/U1117_2_/U3  ( .x(\b[2] ), .a(\U891/U1117_2_/n2 ) );
    nor3_1 \U891/U1117_3_/Unr  ( .x(\U891/U1117_3_/nr ), .a(i[3]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_3_/Und  ( .x(\U891/U1117_3_/nd ), .a(i[3]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_3_/U1  ( .x(\U891/U1117_3_/n2 ), .a(\U891/U1117_3_/n2 ), 
        .b(\U891/U1117_3_/nr ), .c(\U891/U1117_3_/nd ) );
    inv_2 \U891/U1117_3_/U3  ( .x(\b[3] ), .a(\U891/U1117_3_/n2 ) );
    inv_1 \U886/U1126/U3  ( .x(\U886/reset ), .a(nbReset) );
    nor3_1 \U886/U1128/U27  ( .x(\U886/U1128/nb ), .a(\U886/reset ), .b(\f[3] 
        ), .c(\f[2] ) );
    nor2_1 \U886/U1128/U26  ( .x(\U886/U1128/na ), .a(\f[1] ), .b(\f[0] ) );
    nand2_2 \U886/U1128/U29  ( .x(\U886/ackb ), .a(\U886/U1128/nb ), .b(
        \U886/U1128/na ) );
    nor2_1 \U886/U1108/U5  ( .x(\U886/nack ), .a(\U886/acka ), .b(\U886/ackb )
         );
    nor2_2 \U886/U914/U6  ( .x(nba), .a(\U886/acka ), .b(\U886/ackb ) );
    and4_1 \U886/U1127/U25  ( .x(\U886/U1127/n5 ), .a(\U886/U1127/n1 ), .b(
        \U886/U1127/n2 ), .c(\U886/U1127/n3 ), .d(\U886/U1127/n4 ) );
    inv_1 \U886/U1127/U1  ( .x(\U886/U1127/n1 ), .a(\e[3] ) );
    inv_1 \U886/U1127/U2  ( .x(\U886/U1127/n2 ), .a(\e[2] ) );
    inv_1 \U886/U1127/U3  ( .x(\U886/U1127/n3 ), .a(\e[1] ) );
    inv_1 \U886/U1127/U4  ( .x(\U886/U1127/n4 ), .a(\e[0] ) );
    inv_2 \U886/U1127/U5  ( .x(\U886/acka ), .a(\U886/U1127/n5 ) );
    ao222_2 \U886/U1121/U19/U1/U1  ( .x(fsela), .a(\U886/nack ), .b(fsel), .c(
        \U886/nack ), .d(fsela), .e(fsel), .f(fsela) );
    ao222_2 \U886/U1120/U19/U1/U1  ( .x(esela), .a(esel), .b(\U886/nack ), .c(
        esel), .d(esela), .e(\U886/nack ), .f(esela) );
    nor3_1 \U886/U1118_0_/Unr  ( .x(\U886/U1118_0_/nr ), .a(\b[0] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_0_/Und  ( .x(\U886/U1118_0_/nd ), .a(\b[0] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_0_/U1  ( .x(\U886/U1118_0_/n2 ), .a(\U886/U1118_0_/n2 ), 
        .b(\U886/U1118_0_/nr ), .c(\U886/U1118_0_/nd ) );
    inv_2 \U886/U1118_0_/U3  ( .x(\e[0] ), .a(\U886/U1118_0_/n2 ) );
    nor3_1 \U886/U1118_1_/Unr  ( .x(\U886/U1118_1_/nr ), .a(\b[1] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_1_/Und  ( .x(\U886/U1118_1_/nd ), .a(\b[1] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_1_/U1  ( .x(\U886/U1118_1_/n2 ), .a(\U886/U1118_1_/n2 ), 
        .b(\U886/U1118_1_/nr ), .c(\U886/U1118_1_/nd ) );
    inv_2 \U886/U1118_1_/U3  ( .x(\e[1] ), .a(\U886/U1118_1_/n2 ) );
    nor3_1 \U886/U1118_2_/Unr  ( .x(\U886/U1118_2_/nr ), .a(\b[2] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_2_/Und  ( .x(\U886/U1118_2_/nd ), .a(\b[2] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_2_/U1  ( .x(\U886/U1118_2_/n2 ), .a(\U886/U1118_2_/n2 ), 
        .b(\U886/U1118_2_/nr ), .c(\U886/U1118_2_/nd ) );
    inv_2 \U886/U1118_2_/U3  ( .x(\e[2] ), .a(\U886/U1118_2_/n2 ) );
    nor3_1 \U886/U1118_3_/Unr  ( .x(\U886/U1118_3_/nr ), .a(\b[3] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_3_/Und  ( .x(\U886/U1118_3_/nd ), .a(\b[3] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_3_/U1  ( .x(\U886/U1118_3_/n2 ), .a(\U886/U1118_3_/n2 ), 
        .b(\U886/U1118_3_/nr ), .c(\U886/U1118_3_/nd ) );
    inv_2 \U886/U1118_3_/U3  ( .x(\e[3] ), .a(\U886/U1118_3_/n2 ) );
    nor3_1 \U886/U1117_0_/Unr  ( .x(\U886/U1117_0_/nr ), .a(\b[0] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_0_/Und  ( .x(\U886/U1117_0_/nd ), .a(\b[0] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_0_/U1  ( .x(\U886/U1117_0_/n2 ), .a(\U886/U1117_0_/n2 ), 
        .b(\U886/U1117_0_/nr ), .c(\U886/U1117_0_/nd ) );
    inv_2 \U886/U1117_0_/U3  ( .x(\f[0] ), .a(\U886/U1117_0_/n2 ) );
    nor3_1 \U886/U1117_1_/Unr  ( .x(\U886/U1117_1_/nr ), .a(\b[1] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_1_/Und  ( .x(\U886/U1117_1_/nd ), .a(\b[1] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_1_/U1  ( .x(\U886/U1117_1_/n2 ), .a(\U886/U1117_1_/n2 ), 
        .b(\U886/U1117_1_/nr ), .c(\U886/U1117_1_/nd ) );
    inv_2 \U886/U1117_1_/U3  ( .x(\f[1] ), .a(\U886/U1117_1_/n2 ) );
    nor3_1 \U886/U1117_2_/Unr  ( .x(\U886/U1117_2_/nr ), .a(\b[2] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_2_/Und  ( .x(\U886/U1117_2_/nd ), .a(\b[2] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_2_/U1  ( .x(\U886/U1117_2_/n2 ), .a(\U886/U1117_2_/n2 ), 
        .b(\U886/U1117_2_/nr ), .c(\U886/U1117_2_/nd ) );
    inv_2 \U886/U1117_2_/U3  ( .x(\f[2] ), .a(\U886/U1117_2_/n2 ) );
    nor3_1 \U886/U1117_3_/Unr  ( .x(\U886/U1117_3_/nr ), .a(\b[3] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_3_/Und  ( .x(\U886/U1117_3_/nd ), .a(\b[3] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_3_/U1  ( .x(\U886/U1117_3_/n2 ), .a(\U886/U1117_3_/n2 ), 
        .b(\U886/U1117_3_/nr ), .c(\U886/U1117_3_/nd ) );
    inv_2 \U886/U1117_3_/U3  ( .x(\f[3] ), .a(\U886/U1117_3_/n2 ) );
    inv_1 \U884/U1126/U3  ( .x(\U884/reset ), .a(nbReset) );
    nor3_1 \U884/U1128/U27  ( .x(\U884/U1128/nb ), .a(\U884/reset ), .b(\d[3] 
        ), .c(\d[2] ) );
    nor2_1 \U884/U1128/U26  ( .x(\U884/U1128/na ), .a(\d[1] ), .b(\d[0] ) );
    nand2_2 \U884/U1128/U29  ( .x(\U884/ackb ), .a(\U884/U1128/nb ), .b(
        \U884/U1128/na ) );
    nor2_1 \U884/U1108/U5  ( .x(\U884/nack ), .a(\U884/acka ), .b(\U884/ackb )
         );
    nor2_2 \U884/U914/U6  ( .x(naa), .a(\U884/acka ), .b(\U884/ackb ) );
    and4_1 \U884/U1127/U25  ( .x(\U884/U1127/n5 ), .a(\U884/U1127/n1 ), .b(
        \U884/U1127/n2 ), .c(\U884/U1127/n3 ), .d(\U884/U1127/n4 ) );
    inv_1 \U884/U1127/U1  ( .x(\U884/U1127/n1 ), .a(\c[3] ) );
    inv_1 \U884/U1127/U2  ( .x(\U884/U1127/n2 ), .a(\c[2] ) );
    inv_1 \U884/U1127/U3  ( .x(\U884/U1127/n3 ), .a(\c[1] ) );
    inv_1 \U884/U1127/U4  ( .x(\U884/U1127/n4 ), .a(\c[0] ) );
    inv_2 \U884/U1127/U5  ( .x(\U884/acka ), .a(\U884/U1127/n5 ) );
    ao222_2 \U884/U1121/U19/U1/U1  ( .x(dsela), .a(\U884/nack ), .b(dsel), .c(
        \U884/nack ), .d(dsela), .e(dsel), .f(dsela) );
    ao222_2 \U884/U1120/U19/U1/U1  ( .x(csela), .a(csel), .b(\U884/nack ), .c(
        csel), .d(csela), .e(\U884/nack ), .f(csela) );
    nor3_1 \U884/U1118_0_/Unr  ( .x(\U884/U1118_0_/nr ), .a(\a[0] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_0_/Und  ( .x(\U884/U1118_0_/nd ), .a(\a[0] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_0_/U1  ( .x(\U884/U1118_0_/n2 ), .a(\U884/U1118_0_/n2 ), 
        .b(\U884/U1118_0_/nr ), .c(\U884/U1118_0_/nd ) );
    inv_2 \U884/U1118_0_/U3  ( .x(\c[0] ), .a(\U884/U1118_0_/n2 ) );
    nor3_1 \U884/U1118_1_/Unr  ( .x(\U884/U1118_1_/nr ), .a(\a[1] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_1_/Und  ( .x(\U884/U1118_1_/nd ), .a(\a[1] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_1_/U1  ( .x(\U884/U1118_1_/n2 ), .a(\U884/U1118_1_/n2 ), 
        .b(\U884/U1118_1_/nr ), .c(\U884/U1118_1_/nd ) );
    inv_2 \U884/U1118_1_/U3  ( .x(\c[1] ), .a(\U884/U1118_1_/n2 ) );
    nor3_1 \U884/U1118_2_/Unr  ( .x(\U884/U1118_2_/nr ), .a(\a[2] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_2_/Und  ( .x(\U884/U1118_2_/nd ), .a(\a[2] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_2_/U1  ( .x(\U884/U1118_2_/n2 ), .a(\U884/U1118_2_/n2 ), 
        .b(\U884/U1118_2_/nr ), .c(\U884/U1118_2_/nd ) );
    inv_2 \U884/U1118_2_/U3  ( .x(\c[2] ), .a(\U884/U1118_2_/n2 ) );
    nor3_1 \U884/U1118_3_/Unr  ( .x(\U884/U1118_3_/nr ), .a(\a[3] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_3_/Und  ( .x(\U884/U1118_3_/nd ), .a(\a[3] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_3_/U1  ( .x(\U884/U1118_3_/n2 ), .a(\U884/U1118_3_/n2 ), 
        .b(\U884/U1118_3_/nr ), .c(\U884/U1118_3_/nd ) );
    inv_2 \U884/U1118_3_/U3  ( .x(\c[3] ), .a(\U884/U1118_3_/n2 ) );
    nor3_1 \U884/U1117_0_/Unr  ( .x(\U884/U1117_0_/nr ), .a(\a[0] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_0_/Und  ( .x(\U884/U1117_0_/nd ), .a(\a[0] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_0_/U1  ( .x(\U884/U1117_0_/n2 ), .a(\U884/U1117_0_/n2 ), 
        .b(\U884/U1117_0_/nr ), .c(\U884/U1117_0_/nd ) );
    inv_2 \U884/U1117_0_/U3  ( .x(\d[0] ), .a(\U884/U1117_0_/n2 ) );
    nor3_1 \U884/U1117_1_/Unr  ( .x(\U884/U1117_1_/nr ), .a(\a[1] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_1_/Und  ( .x(\U884/U1117_1_/nd ), .a(\a[1] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_1_/U1  ( .x(\U884/U1117_1_/n2 ), .a(\U884/U1117_1_/n2 ), 
        .b(\U884/U1117_1_/nr ), .c(\U884/U1117_1_/nd ) );
    inv_2 \U884/U1117_1_/U3  ( .x(\d[1] ), .a(\U884/U1117_1_/n2 ) );
    nor3_1 \U884/U1117_2_/Unr  ( .x(\U884/U1117_2_/nr ), .a(\a[2] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_2_/Und  ( .x(\U884/U1117_2_/nd ), .a(\a[2] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_2_/U1  ( .x(\U884/U1117_2_/n2 ), .a(\U884/U1117_2_/n2 ), 
        .b(\U884/U1117_2_/nr ), .c(\U884/U1117_2_/nd ) );
    inv_2 \U884/U1117_2_/U3  ( .x(\d[2] ), .a(\U884/U1117_2_/n2 ) );
    nor3_1 \U884/U1117_3_/Unr  ( .x(\U884/U1117_3_/nr ), .a(\a[3] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_3_/Und  ( .x(\U884/U1117_3_/nd ), .a(\a[3] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_3_/U1  ( .x(\U884/U1117_3_/n2 ), .a(\U884/U1117_3_/n2 ), 
        .b(\U884/U1117_3_/nr ), .c(\U884/U1117_3_/nd ) );
    inv_2 \U884/U1117_3_/U3  ( .x(\d[3] ), .a(\U884/U1117_3_/n2 ) );
    nand2_1 \U888/U1128/U5  ( .x(\U888/s ), .a(\U888/r ), .b(\U888/nback ) );
    nand2_1 \U888/U1103/U5  ( .x(\U888/r ), .a(\U888/naack ), .b(\U888/s ) );
    inv_1 \U888/U1111/U3  ( .x(\U888/reset ), .a(nbReset) );
    inv_1 \U888/U1112/U3  ( .x(\U888/naack ), .a(esela) );
    nor2_1 \U888/U1127/U5  ( .x(\U888/nback ), .a(fsela), .b(\U888/reset ) );
    and2_2 \U888/U1129/U8  ( .x(esel), .a(\U888/nback ), .b(\U888/s ) );
    and2_2 \U888/U1124/U8  ( .x(fsel), .a(\U888/r ), .b(\U888/naack ) );
    nand2_1 \U887/U1128/U5  ( .x(\U887/s ), .a(\U887/r ), .b(\U887/nback ) );
    nand2_1 \U887/U1103/U5  ( .x(\U887/r ), .a(\U887/naack ), .b(\U887/s ) );
    inv_1 \U887/U1111/U3  ( .x(\U887/reset ), .a(nbReset) );
    inv_1 \U887/U1112/U3  ( .x(\U887/naack ), .a(csela) );
    nor2_1 \U887/U1127/U5  ( .x(\U887/nback ), .a(dsela), .b(\U887/reset ) );
    and2_2 \U887/U1129/U8  ( .x(csel), .a(\U887/nback ), .b(\U887/s ) );
    and2_2 \U887/U1124/U8  ( .x(dsel), .a(\U887/r ), .b(\U887/naack ) );
    nand2_1 \U885/U1128/U5  ( .x(\U885/s ), .a(\U885/r ), .b(\U885/nback ) );
    nand2_1 \U885/U1103/U5  ( .x(\U885/r ), .a(\U885/naack ), .b(\U885/s ) );
    inv_1 \U885/U1111/U3  ( .x(\U885/reset ), .a(nbReset) );
    inv_1 \U885/U1112/U3  ( .x(\U885/naack ), .a(asela) );
    nor2_1 \U885/U1127/U5  ( .x(\U885/nback ), .a(bsela), .b(\U885/reset ) );
    and2_2 \U885/U1129/U8  ( .x(asel), .a(\U885/nback ), .b(\U885/s ) );
    and2_2 \U885/U1124/U8  ( .x(bsel), .a(\U885/r ), .b(\U885/naack ) );
    nor3_1 \U877/U594/U7  ( .x(\U877/x ), .a(ol[7]), .b(\U877/reset ), .c(oh
        [7]) );
    nor3_1 \U877/U593/U7  ( .x(\U877/y ), .a(ol[6]), .b(\U877/reset ), .c(oh
        [6]) );
    inv_1 \U877/U604/U3  ( .x(\U877/reset ), .a(nbReset) );
    oa31_1 \U877/U590/U25/U1/Uclr  ( .x(\U877/U590/U25/U1/clr ), .a(net135), 
        .b(\cl[3] ), .c(\cl[1] ), .d(oh[6]) );
    oaoi211_1 \U877/U590/U25/U1/Uaoi  ( .x(\U877/U590/U25/U1/ob ), .a(\cl[3] ), 
        .b(\cl[1] ), .c(n1), .d(\U877/U590/U25/U1/clr ) );
    inv_2 \U877/U590/U25/U1/Ui  ( .x(oh[6]), .a(\U877/U590/U25/U1/ob ) );
    oa31_1 \U877/U589/U25/U1/Uclr  ( .x(\U877/U589/U25/U1/clr ), .a(net135), 
        .b(\cl[1] ), .c(\cl[0] ), .d(ol[7]) );
    oaoi211_1 \U877/U589/U25/U1/Uaoi  ( .x(\U877/U589/U25/U1/ob ), .a(\cl[1] ), 
        .b(\cl[0] ), .c(n1), .d(\U877/U589/U25/U1/clr ) );
    inv_2 \U877/U589/U25/U1/Ui  ( .x(ol[7]), .a(\U877/U589/U25/U1/ob ) );
    oa31_1 \U877/U588/U25/U1/Uclr  ( .x(\U877/U588/U25/U1/clr ), .a(net135), 
        .b(\cl[3] ), .c(\cl[2] ), .d(oh[7]) );
    oaoi211_1 \U877/U588/U25/U1/Uaoi  ( .x(\U877/U588/U25/U1/ob ), .a(\cl[3] ), 
        .b(\cl[2] ), .c(n1), .d(\U877/U588/U25/U1/clr ) );
    inv_2 \U877/U588/U25/U1/Ui  ( .x(oh[7]), .a(\U877/U588/U25/U1/ob ) );
    oa31_1 \U877/U591/U25/U1/Uclr  ( .x(\U877/U591/U25/U1/clr ), .a(net135), 
        .b(\cl[2] ), .c(\cl[0] ), .d(ol[6]) );
    oaoi211_1 \U877/U591/U25/U1/Uaoi  ( .x(\U877/U591/U25/U1/ob ), .a(\cl[2] ), 
        .b(\cl[0] ), .c(n1), .d(\U877/U591/U25/U1/clr ) );
    inv_2 \U877/U591/U25/U1/Ui  ( .x(ol[6]), .a(\U877/U591/U25/U1/ob ) );
    ao222_2 \U877/U592/U19/U1/U1  ( .x(ncla), .a(\U877/x ), .b(\U877/y ), .c(
        \U877/x ), .d(ncla), .e(\U877/y ), .f(ncla) );
    nor3_1 \U876/U594/U7  ( .x(\U876/x ), .a(ol[3]), .b(\U876/reset ), .c(oh
        [3]) );
    nor3_1 \U876/U593/U7  ( .x(\U876/y ), .a(ol[2]), .b(\U876/reset ), .c(oh
        [2]) );
    inv_1 \U876/U604/U3  ( .x(\U876/reset ), .a(nbReset) );
    oa31_1 \U876/U590/U25/U1/Uclr  ( .x(\U876/U590/U25/U1/clr ), .a(net135), 
        .b(\d[3] ), .c(\d[1] ), .d(oh[2]) );
    oaoi211_1 \U876/U590/U25/U1/Uaoi  ( .x(\U876/U590/U25/U1/ob ), .a(\d[3] ), 
        .b(\d[1] ), .c(n1), .d(\U876/U590/U25/U1/clr ) );
    inv_2 \U876/U590/U25/U1/Ui  ( .x(oh[2]), .a(\U876/U590/U25/U1/ob ) );
    oa31_1 \U876/U589/U25/U1/Uclr  ( .x(\U876/U589/U25/U1/clr ), .a(net135), 
        .b(\d[1] ), .c(\d[0] ), .d(ol[3]) );
    oaoi211_1 \U876/U589/U25/U1/Uaoi  ( .x(\U876/U589/U25/U1/ob ), .a(\d[1] ), 
        .b(\d[0] ), .c(n1), .d(\U876/U589/U25/U1/clr ) );
    inv_2 \U876/U589/U25/U1/Ui  ( .x(ol[3]), .a(\U876/U589/U25/U1/ob ) );
    oa31_1 \U876/U588/U25/U1/Uclr  ( .x(\U876/U588/U25/U1/clr ), .a(net135), 
        .b(\d[3] ), .c(\d[2] ), .d(oh[3]) );
    oaoi211_1 \U876/U588/U25/U1/Uaoi  ( .x(\U876/U588/U25/U1/ob ), .a(\d[3] ), 
        .b(\d[2] ), .c(n1), .d(\U876/U588/U25/U1/clr ) );
    inv_2 \U876/U588/U25/U1/Ui  ( .x(oh[3]), .a(\U876/U588/U25/U1/ob ) );
    oa31_1 \U876/U591/U25/U1/Uclr  ( .x(\U876/U591/U25/U1/clr ), .a(net135), 
        .b(\d[2] ), .c(\d[0] ), .d(ol[2]) );
    oaoi211_1 \U876/U591/U25/U1/Uaoi  ( .x(\U876/U591/U25/U1/ob ), .a(\d[2] ), 
        .b(\d[0] ), .c(n1), .d(\U876/U591/U25/U1/clr ) );
    inv_2 \U876/U591/U25/U1/Ui  ( .x(ol[2]), .a(\U876/U591/U25/U1/ob ) );
    ao222_2 \U876/U592/U19/U1/U1  ( .x(nda), .a(\U876/x ), .b(\U876/y ), .c(
        \U876/x ), .d(nda), .e(\U876/y ), .f(nda) );
    nor3_1 \U2/U594/U7  ( .x(\U2/x ), .a(ol[1]), .b(\U2/reset ), .c(oh[1]) );
    nor3_1 \U2/U593/U7  ( .x(\U2/y ), .a(ol[0]), .b(\U2/reset ), .c(oh[0]) );
    inv_1 \U2/U604/U3  ( .x(\U2/reset ), .a(nbReset) );
    oa31_1 \U2/U590/U25/U1/Uclr  ( .x(\U2/U590/U25/U1/clr ), .a(net135), .b(
        \f[3] ), .c(\f[1] ), .d(oh[0]) );
    oaoi211_1 \U2/U590/U25/U1/Uaoi  ( .x(\U2/U590/U25/U1/ob ), .a(\f[3] ), .b(
        \f[1] ), .c(n1), .d(\U2/U590/U25/U1/clr ) );
    inv_2 \U2/U590/U25/U1/Ui  ( .x(oh[0]), .a(\U2/U590/U25/U1/ob ) );
    oa31_1 \U2/U589/U25/U1/Uclr  ( .x(\U2/U589/U25/U1/clr ), .a(net135), .b(
        \f[1] ), .c(\f[0] ), .d(ol[1]) );
    oaoi211_1 \U2/U589/U25/U1/Uaoi  ( .x(\U2/U589/U25/U1/ob ), .a(\f[1] ), .b(
        \f[0] ), .c(n1), .d(\U2/U589/U25/U1/clr ) );
    inv_2 \U2/U589/U25/U1/Ui  ( .x(ol[1]), .a(\U2/U589/U25/U1/ob ) );
    oa31_1 \U2/U588/U25/U1/Uclr  ( .x(\U2/U588/U25/U1/clr ), .a(net135), .b(
        \f[3] ), .c(\f[2] ), .d(oh[1]) );
    oaoi211_1 \U2/U588/U25/U1/Uaoi  ( .x(\U2/U588/U25/U1/ob ), .a(\f[3] ), .b(
        \f[2] ), .c(n1), .d(\U2/U588/U25/U1/clr ) );
    inv_2 \U2/U588/U25/U1/Ui  ( .x(oh[1]), .a(\U2/U588/U25/U1/ob ) );
    oa31_1 \U2/U591/U25/U1/Uclr  ( .x(\U2/U591/U25/U1/clr ), .a(net135), .b(
        \f[2] ), .c(\f[0] ), .d(ol[0]) );
    oaoi211_1 \U2/U591/U25/U1/Uaoi  ( .x(\U2/U591/U25/U1/ob ), .a(\f[2] ), .b(
        \f[0] ), .c(n1), .d(\U2/U591/U25/U1/clr ) );
    inv_2 \U2/U591/U25/U1/Ui  ( .x(ol[0]), .a(\U2/U591/U25/U1/ob ) );
    ao222_2 \U2/U592/U19/U1/U1  ( .x(nfa), .a(\U2/x ), .b(\U2/y ), .c(\U2/x ), 
        .d(nfa), .e(\U2/y ), .f(nfa) );
    nor3_1 \U1/U594/U7  ( .x(\U1/x ), .a(ol[5]), .b(\U1/reset ), .c(oh[5]) );
    nor3_1 \U1/U593/U7  ( .x(\U1/y ), .a(ol[4]), .b(\U1/reset ), .c(oh[4]) );
    inv_1 \U1/U604/U3  ( .x(\U1/reset ), .a(nbReset) );
    oa31_1 \U1/U590/U25/U1/Uclr  ( .x(\U1/U590/U25/U1/clr ), .a(net135), .b(
        \e[3] ), .c(\e[1] ), .d(oh[4]) );
    oaoi211_1 \U1/U590/U25/U1/Uaoi  ( .x(\U1/U590/U25/U1/ob ), .a(\e[3] ), .b(
        \e[1] ), .c(n1), .d(\U1/U590/U25/U1/clr ) );
    inv_2 \U1/U590/U25/U1/Ui  ( .x(oh[4]), .a(\U1/U590/U25/U1/ob ) );
    oa31_1 \U1/U589/U25/U1/Uclr  ( .x(\U1/U589/U25/U1/clr ), .a(net135), .b(
        \e[1] ), .c(\e[0] ), .d(ol[5]) );
    oaoi211_1 \U1/U589/U25/U1/Uaoi  ( .x(\U1/U589/U25/U1/ob ), .a(\e[1] ), .b(
        \e[0] ), .c(n1), .d(\U1/U589/U25/U1/clr ) );
    inv_2 \U1/U589/U25/U1/Ui  ( .x(ol[5]), .a(\U1/U589/U25/U1/ob ) );
    oa31_1 \U1/U588/U25/U1/Uclr  ( .x(\U1/U588/U25/U1/clr ), .a(net135), .b(
        \e[3] ), .c(\e[2] ), .d(oh[5]) );
    oaoi211_1 \U1/U588/U25/U1/Uaoi  ( .x(\U1/U588/U25/U1/ob ), .a(\e[3] ), .b(
        \e[2] ), .c(n1), .d(\U1/U588/U25/U1/clr ) );
    inv_2 \U1/U588/U25/U1/Ui  ( .x(oh[5]), .a(\U1/U588/U25/U1/ob ) );
    oa31_1 \U1/U591/U25/U1/Uclr  ( .x(\U1/U591/U25/U1/clr ), .a(net135), .b(
        \e[2] ), .c(\e[0] ), .d(ol[4]) );
    oaoi211_1 \U1/U591/U25/U1/Uaoi  ( .x(\U1/U591/U25/U1/ob ), .a(\e[2] ), .b(
        \e[0] ), .c(n1), .d(\U1/U591/U25/U1/clr ) );
    inv_2 \U1/U591/U25/U1/Ui  ( .x(ol[4]), .a(\U1/U591/U25/U1/ob ) );
    ao222_2 \U1/U592/U19/U1/U1  ( .x(nea), .a(\U1/x ), .b(\U1/y ), .c(\U1/x ), 
        .d(nea), .e(\U1/y ), .f(nea) );
    and3_4 \U881/U20/U9  ( .x(nca), .a(\U881/nack[1] ), .b(\U881/nack[0] ), 
        .c(nbReset) );
    nor2_1 \U881/U18/U5  ( .x(\U881/nack[0] ), .a(\cl[3] ), .b(\cl[0] ) );
    nor2_1 \U881/U19/U5  ( .x(\U881/nack[1] ), .a(\cl[1] ), .b(\cl[2] ) );
    ao222_2 \U881/U15_0_/U19/U1/U1  ( .x(\cl[0] ), .a(\c[0] ), .b(ncla), .c(
        \c[0] ), .d(\cl[0] ), .e(ncla), .f(\cl[0] ) );
    ao222_2 \U881/U15_1_/U19/U1/U1  ( .x(\cl[1] ), .a(\c[1] ), .b(ncla), .c(
        \c[1] ), .d(\cl[1] ), .e(ncla), .f(\cl[1] ) );
    ao222_2 \U881/U15_2_/U19/U1/U1  ( .x(\cl[2] ), .a(\c[2] ), .b(ncla), .c(
        \c[2] ), .d(\cl[2] ), .e(ncla), .f(\cl[2] ) );
    ao222_2 \U881/U15_3_/U19/U1/U1  ( .x(\cl[3] ), .a(\c[3] ), .b(ncla), .c(
        \c[3] ), .d(\cl[3] ), .e(ncla), .f(\cl[3] ) );
    and2_5 U1 ( .x(n1), .a(nbReset), .b(noa) );
    and2_3 U2 ( .x(net135), .a(nbReset), .b(noa) );
endmodule


module chain_selement_ga_73 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_72 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_t_ctrl_2 ( cack, fcdefer, fcslowack, screq, ack, defer, fcack, 
    nReset, scack, slowack );
input  ack, defer, fcack, nReset, scack, slowack;
output cack, fcdefer, fcslowack, screq;
    wire net269, net280, net275, net270, net268, net266, net274, net273, 
        net267, net264, net272, net271, net263, net277, net265, net278, net276, 
        net279, \U49/U28/U1/clr , \U49/U28/U1/set , \U50/U28/U1/clr , 
        \U50/U28/U1/set , \U51/U28/U1/clr , \U51/U28/U1/set , \U57/acb , 
        \U57/U1/Z ;
    chain_selement_ga_73 U55 ( .Aa(net269), .Br(fcdefer), .Ar(net280), .Ba(
        fcack) );
    chain_selement_ga_72 U54 ( .Aa(net275), .Br(fcslowack), .Ar(net270), .Ba(
        fcack) );
    or2_4 \U12/U12  ( .x(net268), .a(net266), .b(net270) );
    or2_4 \U56/U12  ( .x(net274), .a(net275), .b(net269) );
    or2_4 \U14/U12  ( .x(net273), .a(net274), .b(net266) );
    or3_1 \U36/U12  ( .x(cack), .a(net267), .b(net264), .c(net272) );
    nor3_1 \U21/U7  ( .x(net271), .a(net270), .b(net266), .c(net280) );
    and2_1 \U53/U8  ( .x(net263), .a(net271), .b(nReset) );
    and2_1 \U43/U8  ( .x(net277), .a(net265), .b(nReset) );
    nor2_1 \U22/U5  ( .x(net265), .a(net278), .b(net276) );
    ao222_2 \U44/U19/U1/U1  ( .x(net276), .a(net280), .b(net273), .c(net280), 
        .d(net276), .e(net273), .f(net276) );
    ao222_2 \U40/U19/U1/U1  ( .x(net280), .a(net272), .b(net277), .c(net272), 
        .d(net280), .e(net277), .f(net280) );
    ao222_2 \U45/U19/U1/U1  ( .x(net279), .a(net273), .b(net268), .c(net273), 
        .d(net279), .e(net268), .f(net279) );
    ao222_2 \U42/U19/U1/U1  ( .x(net266), .a(net277), .b(net267), .c(net277), 
        .d(net266), .e(net267), .f(net266) );
    ao222_2 \U39/U19/U1/U1  ( .x(net270), .a(net277), .b(net264), .c(net277), 
        .d(net270), .e(net264), .f(net270) );
    aoai211_1 \U49/U28/U1/U1  ( .x(\U49/U28/U1/clr ), .a(ack), .b(nReset), .c(
        net263), .d(net267) );
    nand3_1 \U49/U28/U1/U2  ( .x(\U49/U28/U1/set ), .a(net263), .b(ack), .c(
        nReset) );
    nand2_2 \U49/U28/U1/U3  ( .x(net267), .a(\U49/U28/U1/clr ), .b(
        \U49/U28/U1/set ) );
    aoai211_1 \U50/U28/U1/U1  ( .x(\U50/U28/U1/clr ), .a(slowack), .b(nReset), 
        .c(net263), .d(net264) );
    nand3_1 \U50/U28/U1/U2  ( .x(\U50/U28/U1/set ), .a(net263), .b(slowack), 
        .c(nReset) );
    nand2_2 \U50/U28/U1/U3  ( .x(net264), .a(\U50/U28/U1/clr ), .b(
        \U50/U28/U1/set ) );
    aoai211_1 \U51/U28/U1/U1  ( .x(\U51/U28/U1/clr ), .a(defer), .b(nReset), 
        .c(net263), .d(net272) );
    nand2_2 \U51/U28/U1/U3  ( .x(net272), .a(\U51/U28/U1/clr ), .b(
        \U51/U28/U1/set ) );
    and2_1 \U57/U2/U8  ( .x(screq), .a(net279), .b(\U57/acb ) );
    nor2_1 \U57/U3/U5  ( .x(net278), .a(\U57/acb ), .b(scack) );
    oai21_1 \U57/U1/U30/U1/U1  ( .x(\U57/acb ), .a(\U57/U1/Z ), .b(scack), .c(
        net279) );
    inv_1 \U57/U1/U30/U1/U2  ( .x(\U57/U1/Z ), .a(\U57/acb ) );
    nand3_0 U1 ( .x(\U51/U28/U1/set ), .a(net263), .b(defer), .c(nReset) );
endmodule


module target_dmem ( addr, ccol, chainresponse, crnw, csize, ctag, lock, 
    nchaincommandack, nrouteack, pred, rack, routetxreq, seq, tag_h, tag_l, wd, 
    cack, cdefer, chaincommand, cndefer, cok, err, nReset, nchainresponseack, 
    rd, route, routetxack );
output [63:0] addr;
output [5:0] ccol;
output [4:0] chainresponse;
output [1:0] crnw;
output [3:0] csize;
output [9:0] ctag;
output [1:0] lock;
output [1:0] pred;
output [1:0] seq;
output [4:0] tag_h;
output [4:0] tag_l;
output [63:0] wd;
input  [4:0] chaincommand;
input  [1:0] err;
input  [63:0] rd;
input  [4:0] route;
input  cack, cdefer, cndefer, cok, nReset, nchainresponseack, routetxack;
output nchaincommandack, nrouteack, rack, routetxreq;
    wire read_ctrlack, chainff_ack, read_req, \chainff_l[7] , \chainff_l[6] , 
        \chainff_l[5] , \chainff_l[4] , \chainff_l[3] , \chainff_l[2] , 
        \chainff_l[1] , \chainff_l[0] , \chainff_h[7] , \chainff_h[6] , 
        \chainff_h[5] , \chainff_h[4] , \chainff_h[3] , \chainff_h[2] , 
        \chainff_h[1] , \chainff_h[0] , read_cd, teop, rhdrack, fcack, tcba, 
        net145, n6, screq, fcslowack, fcdefer, read_ack, \rhdr_h[7] , 
        \rhdr_l[7] , \rhdr_l[6] , \rhdr_l[5] , \rhdr_h[6] , \rhdr_h[5] , 
        \rhdr_l[15] , \rhdr_l[14] , \rhdr_l[13] , \rhdr_h[15] , \rhdr_h[14] , 
        \rhdr_h[13] , \tcbl[7] , \tcbl[6] , \tcbl[5] , \tcbl[4] , \tcbl[3] , 
        \tcbl[2] , \tcbl[1] , \tcbl[0] , \tcbh[7] , \tcbh[6] , \tcbh[5] , 
        \tcbh[4] , \tcbh[3] , \tcbh[2] , \tcbh[1] , \tcbh[0] , nbreset, 
        ntresponseack, \tresponse[4] , \tresponse[3] , \tresponse[2] , 
        \tresponse[1] , \tresponse[0] , net200, noba, pullcd, net168, n10, n11, 
        net188, net201, net194, net178, net189, net191, \obl[7] , \obl[6] , 
        \obl[5] , \obl[4] , \obl[3] , \obl[2] , \obl[1] , \obl[0] , \obh[7] , 
        \obh[6] , \obh[5] , \obh[4] , \obh[3] , \obh[2] , \obh[1] , \obh[0] , 
        n13, n14, n12, net284, net265, \chdrack[0] , \U1761/y[0] , 
        \U1761/y[1] , chdrctrlack, hdrcd, \U1761/x[3] , \nchdr_ack[7] , 
        \nchdr_ack[6] , \U1761/U28/Z , \U1761/x[0] , \nchdr_ack[1] , 
        \nchdr_ack[0] , \U1761/U32/Z , \U1761/x[2] , \nchdr_ack[5] , 
        \nchdr_ack[4] , \U1761/U29/Z , \U1761/x[1] , \U1761/U33/Z , 
        \U1761/U30/Z , \nchdr_ack[3] , \nchdr_ack[2] , \U1761/U31/Z , 
        \U1632/Z , \chdrack[1] , \U1676/Z , \U1770/U21/nr , \nchdr_ack[10] , 
        \nchdr_ack[9] , \nchdr_ack[8] , \U1770/U21/nd , \U1770/U21/n2 , 
        \net242[10] , \net244[10] , \net243[10] , \net242[9] , \net244[9] , 
        \net243[9] , \net242[8] , \net244[8] , \net243[8] , \net242[7] , 
        \net244[7] , \net243[7] , \net242[6] , \net244[6] , \net243[6] , 
        \net242[5] , \net244[5] , \net243[5] , \net242[4] , \net244[4] , 
        \net243[4] , \net242[3] , \net244[3] , \net243[3] , \net242[2] , 
        \net244[2] , \net243[2] , \net242[1] , \net244[1] , \net243[1] , 
        \net242[0] , \net244[0] , \net243[0] , \U1574_0_/net231 , n9, n8, 
        \U1574_1_/net231 , n7, \U1574_2_/net231 , \U1574_3_/net231 , 
        \U1574_4_/net231 , \U1574_5_/net231 , \U1574_6_/net231 , 
        \U1574_7_/net231 , \U1574_8_/net231 , \U1574_9_/net231 , 
        \U1574_10_/net231 , net248;
    chain_sendword_2 U1765 ( .ctrlack(read_ctrlack), .oh({\chainff_h[7] , 
        \chainff_h[6] , \chainff_h[5] , \chainff_h[4] , \chainff_h[3] , 
        \chainff_h[2] , \chainff_h[1] , \chainff_h[0] }), .ol({\chainff_l[7] , 
        \chainff_l[6] , \chainff_l[5] , \chainff_l[4] , \chainff_l[3] , 
        \chainff_l[2] , \chainff_l[1] , \chainff_l[0] }), .chainackff(
        chainff_ack), .ctrlreq(read_req), .ih(rd[63:32]), .il(rd[31:0]) );
    chain_dr32bit_completion_10 rd_cd ( .o(read_cd), .i(rd) );
    chain_trhdr_2 xmitHdr ( .chainff_ack(chainff_ack), .chainh({\tcbh[7] , 
        \tcbh[6] , \tcbh[5] , \tcbh[4] , \tcbh[3] , \tcbh[2] , \tcbh[1] , 
        \tcbh[0] }), .chainl({\tcbl[7] , \tcbl[6] , \tcbl[5] , \tcbl[4] , 
        \tcbl[3] , \tcbl[2] , \tcbl[1] , \tcbl[0] }), .eop(teop), .hdrack(
        rhdrack), .normal_ack(rack), .notify_ack(fcack), .read_req(read_req), 
        .routereq(routetxreq), .chain_ff_h({\chainff_h[7] , \chainff_h[6] , 
        \chainff_h[5] , \chainff_h[4] , \chainff_h[3] , \chainff_h[2] , 
        \chainff_h[1] , \chainff_h[0] }), .chainack(tcba), .chainff_l({
        \chainff_l[7] , \chainff_l[6] , \chainff_l[5] , \chainff_l[4] , 
        \chainff_l[3] , \chainff_l[2] , \chainff_l[1] , \chainff_l[0] }), 
        .eopack(net145), .err(err), .nReset(n6), .normal_response(screq), 
        .notify_accept(fcslowack), .notify_defer(fcdefer), .rcol_h({
        \rhdr_h[15] , \rhdr_h[14] , \rhdr_h[13] }), .rcol_l({\rhdr_l[15] , 
        \rhdr_l[14] , \rhdr_l[13] }), .read_ack(read_ack), .rnw_h(\rhdr_h[7] ), 
        .rnw_l(\rhdr_l[7] ), .routeack(routetxack), .rsize_h({\rhdr_h[6] , 
        \rhdr_h[5] }), .rsize_l({\rhdr_l[6] , \rhdr_l[5] }), .rtag_h(tag_h), 
        .rtag_l(tag_l) );
    chain_dr2fr_byte_5 dr2fr ( .eop_ack(net145), .ia(tcba), .o({\tresponse[4] , 
        \tresponse[3] , \tresponse[2] , \tresponse[1] , \tresponse[0] }), 
        .eop(teop), .ih({\tcbh[7] , \tcbh[6] , \tcbh[5] , \tcbh[4] , \tcbh[3] , 
        \tcbh[2] , \tcbh[1] , \tcbh[0] }), .il({\tcbl[7] , \tcbl[6] , 
        \tcbl[5] , \tcbl[4] , \tcbl[3] , \tcbl[2] , \tcbl[1] , \tcbl[0] }), 
        .nReset(nbreset), .noa(ntresponseack) );
    chain_mergepackets_5 merger ( .naa(nrouteack), .nba(ntresponseack), .o(
        chainresponse), .a(route), .b({\tresponse[4] , \tresponse[3] , 
        \tresponse[2] , \tresponse[1] , \tresponse[0] }), .nReset(nbreset), 
        .noa(nchainresponseack) );
    chain_tchdr_2 header ( .addr_req(net200), .col_h(ccol[5:3]), .col_l(ccol
        [2:0]), .itag_h(ctag[9:5]), .itag_l(ctag[4:0]), .lock(lock), .ncback(
        noba), .pred(pred), .pullcd(pullcd), .reset(net168), .rnw_h(n10), 
        .rnw_l(n11), .seq(seq), .size_h({n12, csize[2]}), .size_l({n13, n14}), 
        .write_req(net188), .chwh({\obh[7] , \obh[6] , \obh[5] , \obh[4] , 
        \obh[3] , \obh[2] , \obh[1] , \obh[0] }), .chwl({\obl[7] , \obl[6] , 
        \obl[5] , \obl[4] , \obl[3] , \obl[2] , \obl[1] , \obl[0] }), 
        .addr_ack(net201), .addr_pull(net194), .nReset(n6), .nack(net178), 
        .write_ack(net189), .write_pull(net191) );
    chain_irdemux_32new_5 wd_hld ( .ctrlack(net189), .oh(wd[63:32]), .ol(wd
        [31:0]), .pullreq(net191), .pull_h({\obh[7] , \obh[6] , \obh[5] , 
        \obh[4] , \obh[3] , \obh[2] , \obh[1] , \obh[0] }), .pull_l({\obl[7] , 
        \obl[6] , \obl[5] , \obl[4] , \obl[3] , \obl[2] , \obl[1] , \obl[0] }), 
        .pullcd(pullcd), .reset(net168), .ctrlreq(net188) );
    chain_irdemux_32new_4 adr_hld ( .ctrlack(net201), .oh(addr[63:32]), .ol(
        addr[31:0]), .pullreq(net194), .pull_h({\obh[7] , \obh[6] , \obh[5] , 
        \obh[4] , \obh[3] , \obh[2] , \obh[1] , \obh[0] }), .pull_l({\obl[7] , 
        \obl[6] , \obl[5] , \obl[4] , \obl[3] , \obl[2] , \obl[1] , \obl[0] }), 
        .pullcd(pullcd), .reset(net168), .ctrlreq(net200) );
    chain_fr2dr_byte_2 chain_decoder ( .nia(nchaincommandack), .oh({\obh[7] , 
        \obh[6] , \obh[5] , \obh[4] , \obh[3] , \obh[2] , \obh[1] , \obh[0] }), 
        .ol({\obl[7] , \obl[6] , \obl[5] , \obl[4] , \obl[3] , \obl[2] , 
        \obl[1] , \obl[0] }), .i(chaincommand), .nReset(nbreset), .noa(noba)
         );
    chain_t_ctrl_2 cmd_ctrl ( .cack(net284), .fcdefer(fcdefer), .fcslowack(
        fcslowack), .screq(screq), .ack(cok), .defer(cdefer), .fcack(fcack), 
        .nReset(n6), .scack(rack), .slowack(cndefer) );
    inv_1 \I4/U3  ( .x(net265), .a(nbreset) );
    ao222_1 \U1761/U37/U18/U1/U1  ( .x(\chdrack[0] ), .a(\U1761/y[0] ), .b(
        \U1761/y[1] ), .c(\U1761/y[0] ), .d(\chdrack[0] ), .e(\U1761/y[1] ), 
        .f(\chdrack[0] ) );
    ao222_1 \U1762/U18/U1/U1  ( .x(chdrctrlack), .a(hdrcd), .b(net284), .c(
        hdrcd), .d(chdrctrlack), .e(net284), .f(chdrctrlack) );
    ao222_1 \U1769/U18/U1/U1  ( .x(read_ack), .a(read_ctrlack), .b(read_cd), 
        .c(read_ctrlack), .d(read_ack), .e(read_cd), .f(read_ack) );
    aoi222_1 \U1761/U28/U30/U1  ( .x(\U1761/x[3] ), .a(\nchdr_ack[7] ), .b(
        \nchdr_ack[6] ), .c(\nchdr_ack[7] ), .d(\U1761/U28/Z ), .e(
        \nchdr_ack[6] ), .f(\U1761/U28/Z ) );
    inv_1 \U1761/U28/U30/Uinv  ( .x(\U1761/U28/Z ), .a(\U1761/x[3] ) );
    aoi222_1 \U1761/U32/U30/U1  ( .x(\U1761/x[0] ), .a(\nchdr_ack[1] ), .b(
        \nchdr_ack[0] ), .c(\nchdr_ack[1] ), .d(\U1761/U32/Z ), .e(
        \nchdr_ack[0] ), .f(\U1761/U32/Z ) );
    inv_1 \U1761/U32/U30/Uinv  ( .x(\U1761/U32/Z ), .a(\U1761/x[0] ) );
    aoi222_1 \U1761/U29/U30/U1  ( .x(\U1761/x[2] ), .a(\nchdr_ack[5] ), .b(
        \nchdr_ack[4] ), .c(\nchdr_ack[5] ), .d(\U1761/U29/Z ), .e(
        \nchdr_ack[4] ), .f(\U1761/U29/Z ) );
    inv_1 \U1761/U29/U30/Uinv  ( .x(\U1761/U29/Z ), .a(\U1761/x[2] ) );
    aoi222_1 \U1761/U33/U30/U1  ( .x(\U1761/y[0] ), .a(\U1761/x[1] ), .b(
        \U1761/x[0] ), .c(\U1761/x[1] ), .d(\U1761/U33/Z ), .e(\U1761/x[0] ), 
        .f(\U1761/U33/Z ) );
    inv_1 \U1761/U33/U30/Uinv  ( .x(\U1761/U33/Z ), .a(\U1761/y[0] ) );
    aoi222_1 \U1761/U30/U30/U1  ( .x(\U1761/y[1] ), .a(\U1761/x[3] ), .b(
        \U1761/x[2] ), .c(\U1761/x[3] ), .d(\U1761/U30/Z ), .e(\U1761/x[2] ), 
        .f(\U1761/U30/Z ) );
    inv_1 \U1761/U30/U30/Uinv  ( .x(\U1761/U30/Z ), .a(\U1761/y[1] ) );
    aoi222_1 \U1761/U31/U30/U1  ( .x(\U1761/x[1] ), .a(\nchdr_ack[3] ), .b(
        \nchdr_ack[2] ), .c(\nchdr_ack[3] ), .d(\U1761/U31/Z ), .e(
        \nchdr_ack[2] ), .f(\U1761/U31/Z ) );
    inv_1 \U1761/U31/U30/Uinv  ( .x(\U1761/U31/Z ), .a(\U1761/x[1] ) );
    aoi222_1 \U1632/U30/U1  ( .x(net178), .a(cack), .b(chdrctrlack), .c(cack), 
        .d(\U1632/Z ), .e(chdrctrlack), .f(\U1632/Z ) );
    inv_1 \U1632/U30/Uinv  ( .x(\U1632/Z ), .a(net178) );
    aoi222_1 \U1676/U30/U1  ( .x(hdrcd), .a(\chdrack[0] ), .b(\chdrack[1] ), 
        .c(\chdrack[0] ), .d(\U1676/Z ), .e(\chdrack[1] ), .f(\U1676/Z ) );
    inv_1 \U1676/U30/Uinv  ( .x(\U1676/Z ), .a(hdrcd) );
    nor3_1 \U1770/U21/Unr  ( .x(\U1770/U21/nr ), .a(\nchdr_ack[10] ), .b(
        \nchdr_ack[9] ), .c(\nchdr_ack[8] ) );
    nand3_1 \U1770/U21/Und  ( .x(\U1770/U21/nd ), .a(\nchdr_ack[10] ), .b(
        \nchdr_ack[9] ), .c(\nchdr_ack[8] ) );
    oa21_1 \U1770/U21/U1  ( .x(\U1770/U21/n2 ), .a(\U1770/U21/n2 ), .b(
        \U1770/U21/nr ), .c(\U1770/U21/nd ) );
    inv_1 \U1770/U21/U3  ( .x(\chdrack[1] ), .a(\U1770/U21/n2 ) );
    nor2_1 \U1652_0_/U2/U5  ( .x(\nchdr_ack[0] ), .a(\net242[10] ), .b(
        \net244[10] ) );
    ao222_2 \U1652_0_/U12/U19/U1/U1  ( .x(\net244[10] ), .a(\net243[10] ), .b(
        csize[0]), .c(\net243[10] ), .d(\net244[10] ), .e(csize[0]), .f(
        \net244[10] ) );
    ao222_2 \U1652_0_/U11/U19/U1/U1  ( .x(\net242[10] ), .a(csize[2]), .b(
        \net243[10] ), .c(csize[2]), .d(\net242[10] ), .e(\net243[10] ), .f(
        \net242[10] ) );
    nor2_1 \U1652_1_/U2/U5  ( .x(\nchdr_ack[1] ), .a(\net242[9] ), .b(
        \net244[9] ) );
    ao222_2 \U1652_1_/U12/U19/U1/U1  ( .x(\net244[9] ), .a(\net243[9] ), .b(
        csize[1]), .c(\net243[9] ), .d(\net244[9] ), .e(csize[1]), .f(
        \net244[9] ) );
    ao222_2 \U1652_1_/U11/U19/U1/U1  ( .x(\net242[9] ), .a(csize[3]), .b(
        \net243[9] ), .c(csize[3]), .d(\net242[9] ), .e(\net243[9] ), .f(
        \net242[9] ) );
    nor2_1 \U1652_2_/U2/U5  ( .x(\nchdr_ack[2] ), .a(\net242[8] ), .b(
        \net244[8] ) );
    ao222_2 \U1652_2_/U12/U19/U1/U1  ( .x(\net244[8] ), .a(\net243[8] ), .b(
        crnw[0]), .c(\net243[8] ), .d(\net244[8] ), .e(crnw[0]), .f(
        \net244[8] ) );
    ao222_2 \U1652_2_/U11/U19/U1/U1  ( .x(\net242[8] ), .a(crnw[1]), .b(
        \net243[8] ), .c(crnw[1]), .d(\net242[8] ), .e(\net243[8] ), .f(
        \net242[8] ) );
    nor2_1 \U1652_3_/U2/U5  ( .x(\nchdr_ack[3] ), .a(\net242[7] ), .b(
        \net244[7] ) );
    ao222_2 \U1652_3_/U12/U19/U1/U1  ( .x(\net244[7] ), .a(\net243[7] ), .b(
        ctag[0]), .c(\net243[7] ), .d(\net244[7] ), .e(ctag[0]), .f(
        \net244[7] ) );
    ao222_2 \U1652_3_/U11/U19/U1/U1  ( .x(\net242[7] ), .a(ctag[5]), .b(
        \net243[7] ), .c(ctag[5]), .d(\net242[7] ), .e(\net243[7] ), .f(
        \net242[7] ) );
    nor2_1 \U1652_4_/U2/U5  ( .x(\nchdr_ack[4] ), .a(\net242[6] ), .b(
        \net244[6] ) );
    ao222_2 \U1652_4_/U12/U19/U1/U1  ( .x(\net244[6] ), .a(\net243[6] ), .b(
        ctag[1]), .c(\net243[6] ), .d(\net244[6] ), .e(ctag[1]), .f(
        \net244[6] ) );
    ao222_2 \U1652_4_/U11/U19/U1/U1  ( .x(\net242[6] ), .a(ctag[6]), .b(
        \net243[6] ), .c(ctag[6]), .d(\net242[6] ), .e(\net243[6] ), .f(
        \net242[6] ) );
    nor2_1 \U1652_5_/U2/U5  ( .x(\nchdr_ack[5] ), .a(\net242[5] ), .b(
        \net244[5] ) );
    ao222_2 \U1652_5_/U12/U19/U1/U1  ( .x(\net244[5] ), .a(\net243[5] ), .b(
        ctag[2]), .c(\net243[5] ), .d(\net244[5] ), .e(ctag[2]), .f(
        \net244[5] ) );
    ao222_2 \U1652_5_/U11/U19/U1/U1  ( .x(\net242[5] ), .a(ctag[7]), .b(
        \net243[5] ), .c(ctag[7]), .d(\net242[5] ), .e(\net243[5] ), .f(
        \net242[5] ) );
    nor2_1 \U1652_6_/U2/U5  ( .x(\nchdr_ack[6] ), .a(\net242[4] ), .b(
        \net244[4] ) );
    ao222_2 \U1652_6_/U12/U19/U1/U1  ( .x(\net244[4] ), .a(\net243[4] ), .b(
        ctag[3]), .c(\net243[4] ), .d(\net244[4] ), .e(ctag[3]), .f(
        \net244[4] ) );
    ao222_2 \U1652_6_/U11/U19/U1/U1  ( .x(\net242[4] ), .a(ctag[8]), .b(
        \net243[4] ), .c(ctag[8]), .d(\net242[4] ), .e(\net243[4] ), .f(
        \net242[4] ) );
    nor2_1 \U1652_7_/U2/U5  ( .x(\nchdr_ack[7] ), .a(\net242[3] ), .b(
        \net244[3] ) );
    ao222_2 \U1652_7_/U12/U19/U1/U1  ( .x(\net244[3] ), .a(\net243[3] ), .b(
        ctag[4]), .c(\net243[3] ), .d(\net244[3] ), .e(ctag[4]), .f(
        \net244[3] ) );
    ao222_2 \U1652_7_/U11/U19/U1/U1  ( .x(\net242[3] ), .a(ctag[9]), .b(
        \net243[3] ), .c(ctag[9]), .d(\net242[3] ), .e(\net243[3] ), .f(
        \net242[3] ) );
    nor2_1 \U1652_8_/U2/U5  ( .x(\nchdr_ack[8] ), .a(\net242[2] ), .b(
        \net244[2] ) );
    ao222_2 \U1652_8_/U12/U19/U1/U1  ( .x(\net244[2] ), .a(\net243[2] ), .b(
        ccol[0]), .c(\net243[2] ), .d(\net244[2] ), .e(ccol[0]), .f(
        \net244[2] ) );
    ao222_2 \U1652_8_/U11/U19/U1/U1  ( .x(\net242[2] ), .a(ccol[3]), .b(
        \net243[2] ), .c(ccol[3]), .d(\net242[2] ), .e(\net243[2] ), .f(
        \net242[2] ) );
    nor2_1 \U1652_9_/U2/U5  ( .x(\nchdr_ack[9] ), .a(\net242[1] ), .b(
        \net244[1] ) );
    ao222_2 \U1652_9_/U12/U19/U1/U1  ( .x(\net244[1] ), .a(\net243[1] ), .b(
        ccol[1]), .c(\net243[1] ), .d(\net244[1] ), .e(ccol[1]), .f(
        \net244[1] ) );
    ao222_2 \U1652_9_/U11/U19/U1/U1  ( .x(\net242[1] ), .a(ccol[4]), .b(
        \net243[1] ), .c(ccol[4]), .d(\net242[1] ), .e(\net243[1] ), .f(
        \net242[1] ) );
    nor2_1 \U1652_10_/U2/U5  ( .x(\nchdr_ack[10] ), .a(\net242[0] ), .b(
        \net244[0] ) );
    ao222_2 \U1652_10_/U12/U19/U1/U1  ( .x(\net244[0] ), .a(\net243[0] ), .b(
        ccol[2]), .c(\net243[0] ), .d(\net244[0] ), .e(ccol[2]), .f(
        \net244[0] ) );
    ao222_2 \U1652_10_/U11/U19/U1/U1  ( .x(\net242[0] ), .a(ccol[5]), .b(
        \net243[0] ), .c(ccol[5]), .d(\net242[0] ), .e(\net243[0] ), .f(
        \net242[0] ) );
    nor2_1 \U1574_0_/U2/U5  ( .x(\U1574_0_/net231 ), .a(\rhdr_l[5] ), .b(
        \rhdr_h[5] ) );
    and2_1 \U1574_0_/U13/U8  ( .x(\net243[10] ), .a(\U1574_0_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_0_/U12/U19/U1/U1  ( .x(\rhdr_h[5] ), .a(n9), .b(
        \net242[10] ), .c(n9), .d(\rhdr_h[5] ), .e(\net242[10] ), .f(
        \rhdr_h[5] ) );
    ao222_2 \U1574_0_/U11/U19/U1/U1  ( .x(\rhdr_l[5] ), .a(\net244[10] ), .b(
        n8), .c(\net244[10] ), .d(\rhdr_l[5] ), .e(n9), .f(\rhdr_l[5] ) );
    nor2_1 \U1574_1_/U2/U5  ( .x(\U1574_1_/net231 ), .a(\rhdr_l[6] ), .b(
        \rhdr_h[6] ) );
    and2_1 \U1574_1_/U13/U8  ( .x(\net243[9] ), .a(\U1574_1_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_1_/U12/U19/U1/U1  ( .x(\rhdr_h[6] ), .a(n8), .b(\net242[9] 
        ), .c(n7), .d(\rhdr_h[6] ), .e(\net242[9] ), .f(\rhdr_h[6] ) );
    ao222_2 \U1574_1_/U11/U19/U1/U1  ( .x(\rhdr_l[6] ), .a(\net244[9] ), .b(n8
        ), .c(\net244[9] ), .d(\rhdr_l[6] ), .e(n9), .f(\rhdr_l[6] ) );
    nor2_1 \U1574_2_/U2/U5  ( .x(\U1574_2_/net231 ), .a(\rhdr_l[7] ), .b(
        \rhdr_h[7] ) );
    and2_1 \U1574_2_/U13/U8  ( .x(\net243[8] ), .a(\U1574_2_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_2_/U12/U19/U1/U1  ( .x(\rhdr_h[7] ), .a(n7), .b(\net242[8] 
        ), .c(n7), .d(\rhdr_h[7] ), .e(\net242[8] ), .f(\rhdr_h[7] ) );
    ao222_2 \U1574_2_/U11/U19/U1/U1  ( .x(\rhdr_l[7] ), .a(\net244[8] ), .b(n8
        ), .c(\net244[8] ), .d(\rhdr_l[7] ), .e(n9), .f(\rhdr_l[7] ) );
    nor2_1 \U1574_3_/U2/U5  ( .x(\U1574_3_/net231 ), .a(tag_l[0]), .b(tag_h[0]
        ) );
    and2_1 \U1574_3_/U13/U8  ( .x(\net243[7] ), .a(\U1574_3_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_3_/U12/U19/U1/U1  ( .x(tag_h[0]), .a(n9), .b(\net242[7] ), 
        .c(n7), .d(tag_h[0]), .e(\net242[7] ), .f(tag_h[0]) );
    ao222_2 \U1574_3_/U11/U19/U1/U1  ( .x(tag_l[0]), .a(\net244[7] ), .b(n8), 
        .c(\net244[7] ), .d(tag_l[0]), .e(n7), .f(tag_l[0]) );
    nor2_1 \U1574_4_/U2/U5  ( .x(\U1574_4_/net231 ), .a(tag_l[1]), .b(tag_h[1]
        ) );
    and2_1 \U1574_4_/U13/U8  ( .x(\net243[6] ), .a(\U1574_4_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_4_/U12/U19/U1/U1  ( .x(tag_h[1]), .a(n7), .b(\net242[6] ), 
        .c(n7), .d(tag_h[1]), .e(\net242[6] ), .f(tag_h[1]) );
    ao222_2 \U1574_4_/U11/U19/U1/U1  ( .x(tag_l[1]), .a(\net244[6] ), .b(n8), 
        .c(\net244[6] ), .d(tag_l[1]), .e(n7), .f(tag_l[1]) );
    nor2_1 \U1574_5_/U2/U5  ( .x(\U1574_5_/net231 ), .a(tag_l[2]), .b(tag_h[2]
        ) );
    and2_1 \U1574_5_/U13/U8  ( .x(\net243[5] ), .a(\U1574_5_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_5_/U12/U19/U1/U1  ( .x(tag_h[2]), .a(n8), .b(\net242[5] ), 
        .c(n7), .d(tag_h[2]), .e(\net242[5] ), .f(tag_h[2]) );
    ao222_2 \U1574_5_/U11/U19/U1/U1  ( .x(tag_l[2]), .a(\net244[5] ), .b(n8), 
        .c(\net244[5] ), .d(tag_l[2]), .e(n9), .f(tag_l[2]) );
    nor2_1 \U1574_6_/U2/U5  ( .x(\U1574_6_/net231 ), .a(tag_l[3]), .b(tag_h[3]
        ) );
    and2_1 \U1574_6_/U13/U8  ( .x(\net243[4] ), .a(\U1574_6_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_6_/U12/U19/U1/U1  ( .x(tag_h[3]), .a(n7), .b(\net242[4] ), 
        .c(n9), .d(tag_h[3]), .e(\net242[4] ), .f(tag_h[3]) );
    ao222_2 \U1574_6_/U11/U19/U1/U1  ( .x(tag_l[3]), .a(\net244[4] ), .b(n8), 
        .c(\net244[4] ), .d(tag_l[3]), .e(n7), .f(tag_l[3]) );
    nor2_1 \U1574_7_/U2/U5  ( .x(\U1574_7_/net231 ), .a(tag_l[4]), .b(tag_h[4]
        ) );
    and2_1 \U1574_7_/U13/U8  ( .x(\net243[3] ), .a(\U1574_7_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_7_/U12/U19/U1/U1  ( .x(tag_h[4]), .a(n7), .b(\net242[3] ), 
        .c(n9), .d(tag_h[4]), .e(\net242[3] ), .f(tag_h[4]) );
    ao222_2 \U1574_7_/U11/U19/U1/U1  ( .x(tag_l[4]), .a(\net244[3] ), .b(n8), 
        .c(\net244[3] ), .d(tag_l[4]), .e(n7), .f(tag_l[4]) );
    nor2_1 \U1574_8_/U2/U5  ( .x(\U1574_8_/net231 ), .a(\rhdr_l[13] ), .b(
        \rhdr_h[13] ) );
    and2_1 \U1574_8_/U13/U8  ( .x(\net243[2] ), .a(\U1574_8_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_8_/U12/U19/U1/U1  ( .x(\rhdr_h[13] ), .a(n8), .b(
        \net242[2] ), .c(n9), .d(\rhdr_h[13] ), .e(\net242[2] ), .f(
        \rhdr_h[13] ) );
    ao222_2 \U1574_8_/U11/U19/U1/U1  ( .x(\rhdr_l[13] ), .a(\net244[2] ), .b(
        n8), .c(\net244[2] ), .d(\rhdr_l[13] ), .e(n7), .f(\rhdr_l[13] ) );
    nor2_1 \U1574_9_/U2/U5  ( .x(\U1574_9_/net231 ), .a(\rhdr_l[14] ), .b(
        \rhdr_h[14] ) );
    and2_1 \U1574_9_/U13/U8  ( .x(\net243[1] ), .a(\U1574_9_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_9_/U12/U19/U1/U1  ( .x(\rhdr_h[14] ), .a(n9), .b(
        \net242[1] ), .c(n7), .d(\rhdr_h[14] ), .e(\net242[1] ), .f(
        \rhdr_h[14] ) );
    ao222_2 \U1574_9_/U11/U19/U1/U1  ( .x(\rhdr_l[14] ), .a(\net244[1] ), .b(
        n8), .c(\net244[1] ), .d(\rhdr_l[14] ), .e(n9), .f(\rhdr_l[14] ) );
    nor2_1 \U1574_10_/U2/U5  ( .x(\U1574_10_/net231 ), .a(\rhdr_l[15] ), .b(
        \rhdr_h[15] ) );
    and2_1 \U1574_10_/U13/U8  ( .x(\net243[0] ), .a(\U1574_10_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_10_/U12/U19/U1/U1  ( .x(\rhdr_h[15] ), .a(n9), .b(
        \net242[0] ), .c(n9), .d(\rhdr_h[15] ), .e(\net242[0] ), .f(
        \rhdr_h[15] ) );
    ao222_2 \U1574_10_/U11/U19/U1/U1  ( .x(\rhdr_l[15] ), .a(\net244[0] ), .b(
        n8), .c(\net244[0] ), .d(\rhdr_l[15] ), .e(n9), .f(\rhdr_l[15] ) );
    buf_1 U1 ( .x(csize[0]), .a(n14) );
    buf_1 U2 ( .x(csize[1]), .a(n13) );
    buf_1 U3 ( .x(csize[3]), .a(n12) );
    buf_1 U4 ( .x(crnw[0]), .a(n11) );
    buf_1 U5 ( .x(crnw[1]), .a(n10) );
    inv_5 U6 ( .x(n6), .a(net265) );
    buf_3 U7 ( .x(nbreset), .a(nReset) );
    buf_3 U8 ( .x(n7), .a(net248) );
    buf_3 U9 ( .x(n9), .a(net248) );
    buf_3 U10 ( .x(n8), .a(net248) );
    nor2_1 U11 ( .x(net248), .a(net265), .b(rhdrack) );
endmodule


module t_adec_dmem ( e_h, e_l, r_h, r_l, e_dp, e_ip, e_tic, r_dp, r_ip, r_tic, 
    tag_h, tag_l );
output [2:0] e_h;
output [2:0] e_l;
output [2:0] r_h;
output [2:0] r_l;
input  [2:0] e_dp;
input  [2:0] e_ip;
input  [2:0] e_tic;
input  [2:0] r_dp;
input  [2:0] r_ip;
input  [2:0] r_tic;
input  [4:0] tag_h;
input  [4:0] tag_l;
    wire e_h_1, e_h_0, e_l_2, r_h_1;
    assign e_h[2] = 1'b0;
    assign e_h[1] = e_h_1;
    assign e_h[0] = e_h_0;
    assign e_l[2] = e_l_2;
    assign e_l[1] = e_h_0;
    assign e_l[0] = e_h_1;
    assign r_h[2] = e_h_0;
    assign r_h[1] = r_h_1;
    assign r_h[0] = 1'b0;
    assign r_l[2] = e_h_1;
    assign r_l[0] = e_l_2;
    assign r_h_1 = tag_h[4];
    or2_1 U3 ( .x(r_l[1]), .a(e_h_1), .b(tag_h[3]) );
    buf_3 U6 ( .x(e_h_1), .a(tag_h[2]) );
    or2_2 U7 ( .x(e_h_0), .a(tag_h[3]), .b(r_h_1) );
    or2_2 U8 ( .x(e_l_2), .a(r_h_1), .b(r_l[1]) );
endmodule


module chain_selement_ga_76 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_20 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_symbol_19 ( o, txack, txack_last, e, oa, r, txreq );
output [2:0] o;
input  [1:0] e;
input  [1:0] r;
input  oa, txreq;
output txack, txack_last;
    wire ack, net10, \c[0] , \c[1] ;
    chain_selement_ga_20 U1239 ( .Aa(ack), .Br(net10), .Ar(txreq), .Ba(oa) );
    and2_1 \U1229_0_/U8  ( .x(o[0]), .a(\c[0] ), .b(net10) );
    and2_1 \U1229_1_/U8  ( .x(o[1]), .a(\c[1] ), .b(net10) );
    and2_1 \U1229_2_/U8  ( .x(o[2]), .a(e[1]), .b(net10) );
    ao23_1 \U1251/U19/U21/U1/U1  ( .x(txack_last), .a(ack), .b(txack_last), 
        .c(ack), .d(e[1]), .e(e[1]) );
    ao23_1 \U1250/U19/U21/U1/U1  ( .x(txack), .a(ack), .b(txack), .c(ack), .d(
        e[0]), .e(e[0]) );
    ao222_1 \U1210/U18/U1/U1  ( .x(\c[0] ), .a(e[0]), .b(r[0]), .c(e[0]), .d(
        \c[0] ), .e(r[0]), .f(\c[0] ) );
    ao222_1 \U1209/U18/U1/U1  ( .x(\c[1] ), .a(e[0]), .b(r[1]), .c(e[0]), .d(
        \c[1] ), .e(r[1]), .f(\c[1] ) );
endmodule


module chain_selement_ga_21 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_symbol_20 ( o, txack, txack_last, e, oa, r, txreq );
output [2:0] o;
input  [1:0] e;
input  [1:0] r;
input  oa, txreq;
output txack, txack_last;
    wire ack, net10, \c[0] , \c[1] , n2, n1;
    chain_selement_ga_21 U1239 ( .Aa(ack), .Br(net10), .Ar(txreq), .Ba(oa) );
    and2_1 \U1229_0_/U8  ( .x(o[0]), .a(\c[0] ), .b(net10) );
    and2_1 \U1229_1_/U8  ( .x(o[1]), .a(\c[1] ), .b(net10) );
    and2_1 \U1229_2_/U8  ( .x(o[2]), .a(e[1]), .b(net10) );
    ao23_1 \U1251/U19/U21/U1/U1  ( .x(txack_last), .a(ack), .b(txack_last), 
        .c(ack), .d(e[1]), .e(e[1]) );
    ao23_1 \U1250/U19/U21/U1/U1  ( .x(txack), .a(ack), .b(txack), .c(ack), .d(
        n2), .e(n2) );
    ao222_1 \U1210/U18/U1/U1  ( .x(\c[0] ), .a(n2), .b(r[0]), .c(n2), .d(
        \c[0] ), .e(r[0]), .f(\c[0] ) );
    ao222_1 \U1209/U18/U1/U1  ( .x(\c[1] ), .a(n2), .b(r[1]), .c(n2), .d(
        \c[1] ), .e(r[1]), .f(\c[1] ) );
    inv_0 U1 ( .x(n1), .a(e[0]) );
    inv_2 U2 ( .x(n2), .a(n1) );
endmodule


module chain_selement_ga_19 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_symbol_18 ( o, txack, txack_last, e, oa, r, txreq );
output [2:0] o;
input  [1:0] e;
input  [1:0] r;
input  oa, txreq;
output txack, txack_last;
    wire ack, net10, \c[0] , \c[1] ;
    chain_selement_ga_19 U1239 ( .Aa(ack), .Br(net10), .Ar(txreq), .Ba(oa) );
    and2_1 \U1229_0_/U8  ( .x(o[0]), .a(\c[0] ), .b(net10) );
    and2_1 \U1229_1_/U8  ( .x(o[1]), .a(\c[1] ), .b(net10) );
    and2_1 \U1229_2_/U8  ( .x(o[2]), .a(e[1]), .b(net10) );
    ao23_1 \U1251/U19/U21/U1/U1  ( .x(txack_last), .a(ack), .b(txack_last), 
        .c(ack), .d(e[1]), .e(e[1]) );
    ao23_1 \U1250/U19/U21/U1/U1  ( .x(txack), .a(ack), .b(txack), .c(ack), .d(
        e[0]), .e(e[0]) );
    ao222_1 \U1210/U18/U1/U1  ( .x(\c[0] ), .a(e[0]), .b(r[0]), .c(e[0]), .d(
        \c[0] ), .e(r[0]), .f(\c[0] ) );
    ao222_1 \U1209/U18/U1/U1  ( .x(\c[1] ), .a(e[0]), .b(r[1]), .c(e[0]), .d(
        \c[1] ), .e(r[1]), .f(\c[1] ) );
endmodule


module resp_route_tx_dmem ( o, rtxack, e_h, e_l, noa, r_h, r_l, rtxreq );
output [4:0] o;
input  [2:0] e_h;
input  [2:0] e_l;
input  [2:0] r_h;
input  [2:0] r_l;
input  noa, rtxreq;
output rtxack;
    wire \last[0] , eopsym, net87, net66, net84, \last[2] , net77, \r1[2] , 
        \r1[1] , \r1[0] , \last[1] , \r0[2] , \r0[1] , \r0[0] , \last[3] , 
        \r2[2] , \r2[1] , \r2[0] , net106, net103, \net72[1] , \net72[0] , 
        \I8/nb , \I8/na , \I11/n5 , \I11/n1 , \I11/n2 , \I11/n3 , \I11/n4 , 
        net56, \I7_0_/U25/U1/clr , \I7_0_/U25/U1/ob , \I7_1_/U25/U1/clr , 
        \I7_1_/U25/U1/ob ;
    assign o[3] = 1'b0;
    assign o[2] = 1'b0;
    chain_selement_ga_76 I9 ( .Aa(\last[0] ), .Br(eopsym), .Ar(net87), .Ba(
        net66) );
    route_symbol_19 I2 ( .o({\r1[2] , \r1[1] , \r1[0] }), .txack(net84), 
        .txack_last(\last[2] ), .e({e_h[1], e_l[1]}), .oa(net66), .r({r_h[1], 
        r_l[1]}), .txreq(net77) );
    route_symbol_20 I3 ( .o({\r0[2] , \r0[1] , \r0[0] }), .txack(net87), 
        .txack_last(\last[1] ), .e({e_h[0], e_l[0]}), .oa(net66), .r({r_h[0], 
        r_l[0]}), .txreq(net84) );
    route_symbol_18 I1 ( .o({\r2[2] , \r2[1] , \r2[0] }), .txack(net77), 
        .txack_last(\last[3] ), .e({e_h[2], e_l[2]}), .oa(net66), .r({r_h[2], 
        r_l[2]}), .txreq(rtxreq) );
    nor2_1 \I5/U5  ( .x(net106), .a(eopsym), .b(\r2[2] ) );
    nor2_1 \I16/U5  ( .x(net103), .a(\r1[2] ), .b(\r0[2] ) );
    or2_1 \I14_0_/U12  ( .x(\net72[1] ), .a(\r2[0] ), .b(\r1[0] ) );
    or2_1 \I14_1_/U12  ( .x(\net72[0] ), .a(\r2[1] ), .b(\r1[1] ) );
    nor3_1 \I8/U27  ( .x(\I8/nb ), .a(o[4]), .b(1'b0), .c(1'b0) );
    nor2_1 \I8/U26  ( .x(\I8/na ), .a(o[1]), .b(o[0]) );
    nand2_2 \I8/U29  ( .x(net66), .a(\I8/nb ), .b(\I8/na ) );
    and4_1 \I11/U16  ( .x(\I11/n5 ), .a(\I11/n1 ), .b(\I11/n2 ), .c(\I11/n3 ), 
        .d(\I11/n4 ) );
    inv_1 \I11/U1  ( .x(\I11/n1 ), .a(\last[3] ) );
    inv_1 \I11/U2  ( .x(\I11/n2 ), .a(\last[2] ) );
    inv_1 \I11/U3  ( .x(\I11/n3 ), .a(\last[1] ) );
    inv_1 \I11/U4  ( .x(\I11/n4 ), .a(\last[0] ) );
    inv_1 \I11/U5  ( .x(rtxack), .a(\I11/n5 ) );
    nand2_1 \I17/U5  ( .x(net56), .a(net106), .b(net103) );
    ao222_1 \I15/U18/U1/U1  ( .x(o[4]), .a(noa), .b(net56), .c(noa), .d(o[4]), 
        .e(net56), .f(o[4]) );
    oa31_1 \I7_0_/U25/U1/Uclr  ( .x(\I7_0_/U25/U1/clr ), .a(noa), .b(\r0[0] ), 
        .c(\net72[1] ), .d(o[0]) );
    oaoi211_1 \I7_0_/U25/U1/Uaoi  ( .x(\I7_0_/U25/U1/ob ), .a(\r0[0] ), .b(
        \net72[1] ), .c(noa), .d(\I7_0_/U25/U1/clr ) );
    inv_2 \I7_0_/U25/U1/Ui  ( .x(o[0]), .a(\I7_0_/U25/U1/ob ) );
    oa31_1 \I7_1_/U25/U1/Uclr  ( .x(\I7_1_/U25/U1/clr ), .a(noa), .b(\r0[1] ), 
        .c(\net72[0] ), .d(o[1]) );
    oaoi211_1 \I7_1_/U25/U1/Uaoi  ( .x(\I7_1_/U25/U1/ob ), .a(\r0[1] ), .b(
        \net72[0] ), .c(noa), .d(\I7_1_/U25/U1/clr ) );
    inv_2 \I7_1_/U25/U1/Ui  ( .x(o[1]), .a(\I7_1_/U25/U1/ob ) );
endmodule


module sr2dr_word_8 ( i, req, h, l );
input  [31:0] i;
output [31:0] h;
output [31:0] l;
input  req;
    wire \U31/ni , \U31/nh , \U31/nl , n9, n1, n2, \U30/ni , \U30/nh , 
        \U30/nl , n8, \U29/ni , \U29/nh , \U29/nl , \U28/ni , \U28/nh , 
        \U28/nl , \U27/ni , \U27/nh , \U27/nl , \U26/ni , \U26/nh , \U26/nl , 
        n7, n4, \U25/ni , \U25/nh , \U25/nl , \U24/ni , \U24/nh , \U24/nl , 
        \U23/ni , \U23/nh , \U23/nl , n3, \U22/ni , \U22/nh , \U22/nl , n6, 
        \U21/ni , \U21/nh , \U21/nl , \U20/ni , \U20/nh , \U20/nl , n5, 
        \U19/ni , \U19/nh , \U19/nl , \U18/ni , \U18/nh , \U18/nl , \U17/ni , 
        \U17/nh , \U17/nl , \U16/ni , \U16/nh , \U16/nl , \U15/ni , \U15/nh , 
        \U15/nl , \U14/ni , \U14/nh , \U14/nl , \U13/ni , \U13/nh , \U13/nl , 
        \U12/ni , \U12/nh , \U12/nl , \U11/ni , \U11/nh , \U11/nl , \U10/ni , 
        \U10/nh , \U10/nl , \U9/ni , \U9/nh , \U9/nl , \U8/ni , \U8/nh , 
        \U8/nl , \U7/ni , \U7/nh , \U7/nl , \U6/ni , \U6/nh , \U6/nl , \U5/ni , 
        \U5/nh , \U5/nl , \U4/ni , \U4/nh , \U4/nl , \U3/ni , \U3/nh , \U3/nl , 
        \U2/ni , \U2/nh , \U2/nl , \U1/ni , \U1/nh , \U1/nl , \U0/ni , \U0/nh , 
        \U0/nl , n12, n11, n10;
    inv_1 \U31/Uii  ( .x(\U31/ni ), .a(i[31]) );
    inv_1 \U31/Uih  ( .x(\U31/nh ), .a(h[31]) );
    inv_1 \U31/Uil  ( .x(\U31/nl ), .a(l[31]) );
    ao23_1 \U31/Ucl/U1/U1  ( .x(l[31]), .a(n9), .b(l[31]), .c(n1), .d(\U31/ni 
        ), .e(\U31/nh ) );
    ao23_1 \U31/Uch/U1/U1  ( .x(h[31]), .a(n9), .b(h[31]), .c(n2), .d(i[31]), 
        .e(\U31/nl ) );
    inv_1 \U30/Uii  ( .x(\U30/ni ), .a(i[30]) );
    inv_1 \U30/Uih  ( .x(\U30/nh ), .a(h[30]) );
    inv_1 \U30/Uil  ( .x(\U30/nl ), .a(l[30]) );
    ao23_1 \U30/Ucl/U1/U1  ( .x(l[30]), .a(n8), .b(l[30]), .c(n1), .d(\U30/ni 
        ), .e(\U30/nh ) );
    ao23_1 \U30/Uch/U1/U1  ( .x(h[30]), .a(n8), .b(h[30]), .c(n1), .d(i[30]), 
        .e(\U30/nl ) );
    inv_1 \U29/Uii  ( .x(\U29/ni ), .a(i[29]) );
    inv_1 \U29/Uih  ( .x(\U29/nh ), .a(h[29]) );
    inv_1 \U29/Uil  ( .x(\U29/nl ), .a(l[29]) );
    ao23_1 \U29/Ucl/U1/U1  ( .x(l[29]), .a(n8), .b(l[29]), .c(n1), .d(\U29/ni 
        ), .e(\U29/nh ) );
    ao23_1 \U29/Uch/U1/U1  ( .x(h[29]), .a(n8), .b(h[29]), .c(n2), .d(i[29]), 
        .e(\U29/nl ) );
    inv_1 \U28/Uii  ( .x(\U28/ni ), .a(i[28]) );
    inv_1 \U28/Uih  ( .x(\U28/nh ), .a(h[28]) );
    inv_1 \U28/Uil  ( .x(\U28/nl ), .a(l[28]) );
    ao23_1 \U28/Ucl/U1/U1  ( .x(l[28]), .a(n8), .b(l[28]), .c(n2), .d(\U28/ni 
        ), .e(\U28/nh ) );
    ao23_1 \U28/Uch/U1/U1  ( .x(h[28]), .a(n8), .b(h[28]), .c(n2), .d(i[28]), 
        .e(\U28/nl ) );
    inv_1 \U27/Uii  ( .x(\U27/ni ), .a(i[27]) );
    inv_1 \U27/Uih  ( .x(\U27/nh ), .a(h[27]) );
    inv_1 \U27/Uil  ( .x(\U27/nl ), .a(l[27]) );
    ao23_1 \U27/Ucl/U1/U1  ( .x(l[27]), .a(n8), .b(l[27]), .c(n2), .d(\U27/ni 
        ), .e(\U27/nh ) );
    ao23_1 \U27/Uch/U1/U1  ( .x(h[27]), .a(n8), .b(h[27]), .c(n2), .d(i[27]), 
        .e(\U27/nl ) );
    inv_1 \U26/Uii  ( .x(\U26/ni ), .a(i[26]) );
    inv_1 \U26/Uih  ( .x(\U26/nh ), .a(h[26]) );
    inv_1 \U26/Uil  ( .x(\U26/nl ), .a(l[26]) );
    ao23_1 \U26/Ucl/U1/U1  ( .x(l[26]), .a(n7), .b(l[26]), .c(n2), .d(\U26/ni 
        ), .e(\U26/nh ) );
    ao23_1 \U26/Uch/U1/U1  ( .x(h[26]), .a(n7), .b(h[26]), .c(n4), .d(i[26]), 
        .e(\U26/nl ) );
    inv_1 \U25/Uii  ( .x(\U25/ni ), .a(i[25]) );
    inv_1 \U25/Uih  ( .x(\U25/nh ), .a(h[25]) );
    inv_1 \U25/Uil  ( .x(\U25/nl ), .a(l[25]) );
    ao23_1 \U25/Ucl/U1/U1  ( .x(l[25]), .a(n7), .b(l[25]), .c(n4), .d(\U25/ni 
        ), .e(\U25/nh ) );
    ao23_1 \U25/Uch/U1/U1  ( .x(h[25]), .a(n7), .b(h[25]), .c(n4), .d(i[25]), 
        .e(\U25/nl ) );
    inv_1 \U24/Uii  ( .x(\U24/ni ), .a(i[24]) );
    inv_1 \U24/Uih  ( .x(\U24/nh ), .a(h[24]) );
    inv_1 \U24/Uil  ( .x(\U24/nl ), .a(l[24]) );
    ao23_1 \U24/Ucl/U1/U1  ( .x(l[24]), .a(n7), .b(l[24]), .c(n4), .d(\U24/ni 
        ), .e(\U24/nh ) );
    ao23_1 \U24/Uch/U1/U1  ( .x(h[24]), .a(n7), .b(h[24]), .c(n4), .d(i[24]), 
        .e(\U24/nl ) );
    inv_1 \U23/Uii  ( .x(\U23/ni ), .a(i[23]) );
    inv_1 \U23/Uih  ( .x(\U23/nh ), .a(h[23]) );
    inv_1 \U23/Uil  ( .x(\U23/nl ), .a(l[23]) );
    ao23_1 \U23/Ucl/U1/U1  ( .x(l[23]), .a(n7), .b(l[23]), .c(n3), .d(\U23/ni 
        ), .e(\U23/nh ) );
    ao23_1 \U23/Uch/U1/U1  ( .x(h[23]), .a(n7), .b(h[23]), .c(n3), .d(i[23]), 
        .e(\U23/nl ) );
    inv_1 \U22/Uii  ( .x(\U22/ni ), .a(i[22]) );
    inv_1 \U22/Uih  ( .x(\U22/nh ), .a(h[22]) );
    inv_1 \U22/Uil  ( .x(\U22/nl ), .a(l[22]) );
    ao23_1 \U22/Ucl/U1/U1  ( .x(l[22]), .a(n6), .b(l[22]), .c(n3), .d(\U22/ni 
        ), .e(\U22/nh ) );
    ao23_1 \U22/Uch/U1/U1  ( .x(h[22]), .a(n6), .b(h[22]), .c(n3), .d(i[22]), 
        .e(\U22/nl ) );
    inv_1 \U21/Uii  ( .x(\U21/ni ), .a(i[21]) );
    inv_1 \U21/Uih  ( .x(\U21/nh ), .a(h[21]) );
    inv_1 \U21/Uil  ( .x(\U21/nl ), .a(l[21]) );
    ao23_1 \U21/Ucl/U1/U1  ( .x(l[21]), .a(n6), .b(l[21]), .c(n3), .d(\U21/ni 
        ), .e(\U21/nh ) );
    ao23_1 \U21/Uch/U1/U1  ( .x(h[21]), .a(n6), .b(h[21]), .c(n3), .d(i[21]), 
        .e(\U21/nl ) );
    inv_1 \U20/Uii  ( .x(\U20/ni ), .a(i[20]) );
    inv_1 \U20/Uih  ( .x(\U20/nh ), .a(h[20]) );
    inv_1 \U20/Uil  ( .x(\U20/nl ), .a(l[20]) );
    ao23_1 \U20/Ucl/U1/U1  ( .x(l[20]), .a(n6), .b(l[20]), .c(n5), .d(\U20/ni 
        ), .e(\U20/nh ) );
    ao23_1 \U20/Uch/U1/U1  ( .x(h[20]), .a(n6), .b(h[20]), .c(n4), .d(i[20]), 
        .e(\U20/nl ) );
    inv_1 \U19/Uii  ( .x(\U19/ni ), .a(i[19]) );
    inv_1 \U19/Uih  ( .x(\U19/nh ), .a(h[19]) );
    inv_1 \U19/Uil  ( .x(\U19/nl ), .a(l[19]) );
    ao23_1 \U19/Ucl/U1/U1  ( .x(l[19]), .a(n6), .b(l[19]), .c(n4), .d(\U19/ni 
        ), .e(\U19/nh ) );
    ao23_1 \U19/Uch/U1/U1  ( .x(h[19]), .a(n6), .b(h[19]), .c(n4), .d(i[19]), 
        .e(\U19/nl ) );
    inv_1 \U18/Uii  ( .x(\U18/ni ), .a(i[18]) );
    inv_1 \U18/Uih  ( .x(\U18/nh ), .a(h[18]) );
    inv_1 \U18/Uil  ( .x(\U18/nl ), .a(l[18]) );
    ao23_1 \U18/Ucl/U1/U1  ( .x(l[18]), .a(n5), .b(l[18]), .c(n5), .d(\U18/ni 
        ), .e(\U18/nh ) );
    ao23_1 \U18/Uch/U1/U1  ( .x(h[18]), .a(n5), .b(h[18]), .c(n5), .d(i[18]), 
        .e(\U18/nl ) );
    inv_1 \U17/Uii  ( .x(\U17/ni ), .a(i[17]) );
    inv_1 \U17/Uih  ( .x(\U17/nh ), .a(h[17]) );
    inv_1 \U17/Uil  ( .x(\U17/nl ), .a(l[17]) );
    ao23_1 \U17/Ucl/U1/U1  ( .x(l[17]), .a(n6), .b(l[17]), .c(n5), .d(\U17/ni 
        ), .e(\U17/nh ) );
    ao23_1 \U17/Uch/U1/U1  ( .x(h[17]), .a(n7), .b(h[17]), .c(n4), .d(i[17]), 
        .e(\U17/nl ) );
    inv_1 \U16/Uii  ( .x(\U16/ni ), .a(i[16]) );
    inv_1 \U16/Uih  ( .x(\U16/nh ), .a(h[16]) );
    inv_1 \U16/Uil  ( .x(\U16/nl ), .a(l[16]) );
    ao23_1 \U16/Ucl/U1/U1  ( .x(l[16]), .a(n9), .b(l[16]), .c(n3), .d(\U16/ni 
        ), .e(\U16/nh ) );
    ao23_1 \U16/Uch/U1/U1  ( .x(h[16]), .a(n9), .b(h[16]), .c(n1), .d(i[16]), 
        .e(\U16/nl ) );
    inv_1 \U15/Uii  ( .x(\U15/ni ), .a(i[15]) );
    inv_1 \U15/Uih  ( .x(\U15/nh ), .a(h[15]) );
    inv_1 \U15/Uil  ( .x(\U15/nl ), .a(l[15]) );
    ao23_1 \U15/Ucl/U1/U1  ( .x(l[15]), .a(n8), .b(l[15]), .c(n1), .d(\U15/ni 
        ), .e(\U15/nh ) );
    ao23_1 \U15/Uch/U1/U1  ( .x(h[15]), .a(n7), .b(h[15]), .c(n1), .d(i[15]), 
        .e(\U15/nl ) );
    inv_1 \U14/Uii  ( .x(\U14/ni ), .a(i[14]) );
    inv_1 \U14/Uih  ( .x(\U14/nh ), .a(h[14]) );
    inv_1 \U14/Uil  ( .x(\U14/nl ), .a(l[14]) );
    ao23_1 \U14/Ucl/U1/U1  ( .x(l[14]), .a(n6), .b(l[14]), .c(n1), .d(\U14/ni 
        ), .e(\U14/nh ) );
    ao23_1 \U14/Uch/U1/U1  ( .x(h[14]), .a(n6), .b(h[14]), .c(n3), .d(i[14]), 
        .e(\U14/nl ) );
    inv_1 \U13/Uii  ( .x(\U13/ni ), .a(i[13]) );
    inv_1 \U13/Uih  ( .x(\U13/nh ), .a(h[13]) );
    inv_1 \U13/Uil  ( .x(\U13/nl ), .a(l[13]) );
    ao23_1 \U13/Ucl/U1/U1  ( .x(l[13]), .a(n6), .b(l[13]), .c(n4), .d(\U13/ni 
        ), .e(\U13/nh ) );
    ao23_1 \U13/Uch/U1/U1  ( .x(h[13]), .a(n6), .b(h[13]), .c(n4), .d(i[13]), 
        .e(\U13/nl ) );
    inv_1 \U12/Uii  ( .x(\U12/ni ), .a(i[12]) );
    inv_1 \U12/Uih  ( .x(\U12/nh ), .a(h[12]) );
    inv_1 \U12/Uil  ( .x(\U12/nl ), .a(l[12]) );
    ao23_1 \U12/Ucl/U1/U1  ( .x(l[12]), .a(n5), .b(l[12]), .c(n4), .d(\U12/ni 
        ), .e(\U12/nh ) );
    ao23_1 \U12/Uch/U1/U1  ( .x(h[12]), .a(n5), .b(h[12]), .c(n4), .d(i[12]), 
        .e(\U12/nl ) );
    inv_1 \U11/Uii  ( .x(\U11/ni ), .a(i[11]) );
    inv_1 \U11/Uih  ( .x(\U11/nh ), .a(h[11]) );
    inv_1 \U11/Uil  ( .x(\U11/nl ), .a(l[11]) );
    ao23_1 \U11/Ucl/U1/U1  ( .x(l[11]), .a(n5), .b(l[11]), .c(n4), .d(\U11/ni 
        ), .e(\U11/nh ) );
    ao23_1 \U11/Uch/U1/U1  ( .x(h[11]), .a(n5), .b(h[11]), .c(n4), .d(i[11]), 
        .e(\U11/nl ) );
    inv_1 \U10/Uii  ( .x(\U10/ni ), .a(i[10]) );
    inv_1 \U10/Uih  ( .x(\U10/nh ), .a(h[10]) );
    inv_1 \U10/Uil  ( .x(\U10/nl ), .a(l[10]) );
    ao23_1 \U10/Ucl/U1/U1  ( .x(l[10]), .a(n5), .b(l[10]), .c(n3), .d(\U10/ni 
        ), .e(\U10/nh ) );
    ao23_1 \U10/Uch/U1/U1  ( .x(h[10]), .a(n5), .b(h[10]), .c(n3), .d(i[10]), 
        .e(\U10/nl ) );
    inv_1 \U9/Uii  ( .x(\U9/ni ), .a(i[9]) );
    inv_1 \U9/Uih  ( .x(\U9/nh ), .a(h[9]) );
    inv_1 \U9/Uil  ( .x(\U9/nl ), .a(l[9]) );
    ao23_1 \U9/Ucl/U1/U1  ( .x(l[9]), .a(n5), .b(l[9]), .c(n3), .d(\U9/ni ), 
        .e(\U9/nh ) );
    ao23_1 \U9/Uch/U1/U1  ( .x(h[9]), .a(n5), .b(h[9]), .c(n3), .d(i[9]), .e(
        \U9/nl ) );
    inv_1 \U8/Uii  ( .x(\U8/ni ), .a(i[8]) );
    inv_1 \U8/Uih  ( .x(\U8/nh ), .a(h[8]) );
    inv_1 \U8/Uil  ( .x(\U8/nl ), .a(l[8]) );
    ao23_1 \U8/Ucl/U1/U1  ( .x(l[8]), .a(n5), .b(l[8]), .c(n3), .d(\U8/ni ), 
        .e(\U8/nh ) );
    ao23_1 \U8/Uch/U1/U1  ( .x(h[8]), .a(n5), .b(h[8]), .c(n3), .d(i[8]), .e(
        \U8/nl ) );
    inv_1 \U7/Uii  ( .x(\U7/ni ), .a(i[7]) );
    inv_1 \U7/Uih  ( .x(\U7/nh ), .a(h[7]) );
    inv_1 \U7/Uil  ( .x(\U7/nl ), .a(l[7]) );
    ao23_1 \U7/Ucl/U1/U1  ( .x(l[7]), .a(n7), .b(l[7]), .c(n3), .d(\U7/ni ), 
        .e(\U7/nh ) );
    ao23_1 \U7/Uch/U1/U1  ( .x(h[7]), .a(n7), .b(h[7]), .c(n2), .d(i[7]), .e(
        \U7/nl ) );
    inv_1 \U6/Uii  ( .x(\U6/ni ), .a(i[6]) );
    inv_1 \U6/Uih  ( .x(\U6/nh ), .a(h[6]) );
    inv_1 \U6/Uil  ( .x(\U6/nl ), .a(l[6]) );
    ao23_1 \U6/Ucl/U1/U1  ( .x(l[6]), .a(n7), .b(l[6]), .c(n2), .d(\U6/ni ), 
        .e(\U6/nh ) );
    ao23_1 \U6/Uch/U1/U1  ( .x(h[6]), .a(n7), .b(h[6]), .c(n2), .d(i[6]), .e(
        \U6/nl ) );
    inv_1 \U5/Uii  ( .x(\U5/ni ), .a(i[5]) );
    inv_1 \U5/Uih  ( .x(\U5/nh ), .a(h[5]) );
    inv_1 \U5/Uil  ( .x(\U5/nl ), .a(l[5]) );
    ao23_1 \U5/Ucl/U1/U1  ( .x(l[5]), .a(n7), .b(l[5]), .c(n2), .d(\U5/ni ), 
        .e(\U5/nh ) );
    ao23_1 \U5/Uch/U1/U1  ( .x(h[5]), .a(n7), .b(h[5]), .c(n2), .d(i[5]), .e(
        \U5/nl ) );
    inv_1 \U4/Uii  ( .x(\U4/ni ), .a(i[4]) );
    inv_1 \U4/Uih  ( .x(\U4/nh ), .a(h[4]) );
    inv_1 \U4/Uil  ( .x(\U4/nl ), .a(l[4]) );
    ao23_1 \U4/Ucl/U1/U1  ( .x(l[4]), .a(n6), .b(l[4]), .c(n2), .d(\U4/ni ), 
        .e(\U4/nh ) );
    ao23_1 \U4/Uch/U1/U1  ( .x(h[4]), .a(n6), .b(h[4]), .c(n2), .d(i[4]), .e(
        \U4/nl ) );
    inv_1 \U3/Uii  ( .x(\U3/ni ), .a(i[3]) );
    inv_1 \U3/Uih  ( .x(\U3/nh ), .a(h[3]) );
    inv_1 \U3/Uil  ( .x(\U3/nl ), .a(l[3]) );
    ao23_1 \U3/Ucl/U1/U1  ( .x(l[3]), .a(n6), .b(l[3]), .c(n2), .d(\U3/ni ), 
        .e(\U3/nh ) );
    ao23_1 \U3/Uch/U1/U1  ( .x(h[3]), .a(n8), .b(h[3]), .c(n1), .d(i[3]), .e(
        \U3/nl ) );
    inv_1 \U2/Uii  ( .x(\U2/ni ), .a(i[2]) );
    inv_1 \U2/Uih  ( .x(\U2/nh ), .a(h[2]) );
    inv_1 \U2/Uil  ( .x(\U2/nl ), .a(l[2]) );
    ao23_1 \U2/Ucl/U1/U1  ( .x(l[2]), .a(n8), .b(l[2]), .c(n1), .d(\U2/ni ), 
        .e(\U2/nh ) );
    ao23_1 \U2/Uch/U1/U1  ( .x(h[2]), .a(n8), .b(h[2]), .c(n1), .d(i[2]), .e(
        \U2/nl ) );
    inv_1 \U1/Uii  ( .x(\U1/ni ), .a(i[1]) );
    inv_1 \U1/Uih  ( .x(\U1/nh ), .a(h[1]) );
    inv_1 \U1/Uil  ( .x(\U1/nl ), .a(l[1]) );
    ao23_1 \U1/Ucl/U1/U1  ( .x(l[1]), .a(n8), .b(l[1]), .c(n1), .d(\U1/ni ), 
        .e(\U1/nh ) );
    ao23_1 \U1/Uch/U1/U1  ( .x(h[1]), .a(n8), .b(h[1]), .c(n1), .d(i[1]), .e(
        \U1/nl ) );
    inv_1 \U0/Uii  ( .x(\U0/ni ), .a(i[0]) );
    inv_1 \U0/Uih  ( .x(\U0/nh ), .a(h[0]) );
    inv_1 \U0/Uil  ( .x(\U0/nl ), .a(l[0]) );
    ao23_1 \U0/Ucl/U1/U1  ( .x(l[0]), .a(n8), .b(l[0]), .c(n1), .d(\U0/ni ), 
        .e(\U0/nh ) );
    ao23_1 \U0/Uch/U1/U1  ( .x(h[0]), .a(n8), .b(h[0]), .c(n1), .d(i[0]), .e(
        \U0/nl ) );
    buf_16 U1 ( .x(n1), .a(n12) );
    buf_16 U2 ( .x(n2), .a(n12) );
    buf_16 U3 ( .x(n3), .a(n12) );
    buf_16 U4 ( .x(n4), .a(n11) );
    buf_16 U5 ( .x(n5), .a(n11) );
    buf_16 U6 ( .x(n6), .a(n11) );
    buf_16 U7 ( .x(n7), .a(n10) );
    buf_16 U8 ( .x(n8), .a(n10) );
    buf_16 U9 ( .x(n9), .a(n10) );
    buf_16 U10 ( .x(n10), .a(req) );
    buf_16 U11 ( .x(n11), .a(req) );
    buf_16 U12 ( .x(n12), .a(req) );
endmodule


module matched_delay_cp2slave_resp_dmem ( x, a );
input  a;
output x;
    buf_1 I1 ( .x(x), .a(a) );
endmodule


module matched_delay_cp2slave_comdmem ( x, a );
input  a;
output x;
    buf_1 I1 ( .x(x), .a(a) );
endmodule


module cp2slave_dmem ( tc_seq, tc_size, tc_itag, tc_wd, tc_lock, tc_a, tc_rnw, 
    tc_ok, tc_defer, tc_slow, tc_ack, req_in, ts_i, st_i, we_i, mult_i, adr_i, 
    dat_i, seq_i, prd_i, sel_i, ack_in, tr_rd, tr_err, tr_size, tr_ack, tr_rnw, 
    req_out, dat_o, err_o, rty_o, acc_o, sel_o, mult_o, rt_o, ack_out, reset
     );
input  [1:0] tc_seq;
input  [3:0] tc_size;
input  [9:0] tc_itag;
input  [63:0] tc_wd;
input  [1:0] tc_lock;
input  [63:0] tc_a;
input  [1:0] tc_rnw;
output [2:0] ts_i;
output [4:0] st_i;
output [31:0] adr_i;
output [31:0] dat_i;
output [3:0] sel_i;
output [63:0] tr_rd;
output [1:0] tr_err;
output [3:0] tr_size;
output [1:0] tr_rnw;
input  [31:0] dat_o;
input  [3:0] sel_o;
input  [4:0] rt_o;
input  ack_in, tr_ack, req_out, err_o, rty_o, acc_o, mult_o, reset;
output tc_ok, tc_defer, tc_slow, tc_ack, req_in, we_i, mult_i, seq_i, prd_i, 
    ack_out;
    wire tc_wd_63, tc_wd_62, tc_wd_61, tc_wd_60, tc_wd_59, tc_wd_58, tc_wd_56, 
        tc_wd_55, tc_wd_54, tc_wd_53, tc_wd_52, tc_wd_51, tc_wd_50, tc_wd_49, 
        tc_wd_48, tc_wd_47, tc_wd_46, tc_wd_45, tc_wd_44, tc_wd_43, tc_wd_40, 
        tc_wd_39, tc_wd_38, tc_wd_36, tc_wd_32, tc_a_60, tc_a_58, sel_i_3, n1, 
        n334, n311, n129, n309, n310, n315, n348, n349, n350, n456, n336, n457, 
        n345, n303, n505, n193, n476, n479, n229, n226, n257, n263, n260, n268, 
        n269, n270, n265, n266, n267, n277, n252, n248, n249, n250, n245, n246, 
        n247, n242, n243, n244, n222, n223, n224, n220, n234, n235, n236, n231, 
        n232, n233, n205, n206, n207, n203, n199, n200, n201, n197, n218, n214, 
        n215, n216, n211, n212, n213, n208, n209, n210, n374, n375, n368, n251, 
        n280, n274, n271, n427, n196, n424, n202, n240, n237, n413, n219, n421, 
        n418, n416, n428, n425, n422, n414, n411, n408, n238, n272, n351, n366, 
        n335, n355, n531, n532, respond, n313, n121, n122, n359, n360, n123, 
        n337, n124, n125, n126, n127, n217, n128, n312, n130, n284, n285, n449, 
        n282, n283, n380, n279, n276, n397, n454, n463, n453, n395, n404, n383, 
        n443, n477, n455, n230, n135, n305, n487, n302, n445, n446, n442, n136, 
        n320, n400, n137, n340, n198, n386, n381, n478, n475, n407, n402, n204, 
        n221, n141, n321, n483, n484, n485, n480, n474, n227, n188, n517, n525, 
        n180, n401, n387, n394, n481, n482, n491, n195, n492, n369, n181, n429, 
        n415, n324, n343, n363, n319, n344, n354, n304, n330, n497, n496, n291, 
        n438, n373, n367, n439, n440, n333, n308, n297, n347, n301, n503, n499, 
        n502, n498, n288, n327, n316, n298, n294, n358, complb0, n189, n510, 
        n507, n192, n473, n508, n471, n488, n489, n490, complw0, n182, n183, 
        n184, n185, n364, n365, n391, n388, n430, n423, n426, n431, n417, n419, 
        n420, n432, n409, n410, n412, n433, n403, n405, n406, n434, n396, n398, 
        n399, n435, n389, n390, n392, n393, n436, n382, n384, n385, n437, n376, 
        n377, n378, n379, n441, n370, n444, n470, n472, n194, n486, n493, n494, 
        n495, n191, n500, n501, n504, n506, n509, n511, n465, n466, n468, n512, 
        n460, n513, n514, n462, n459, n515, n516, n518, n452, n519, n450, n520, 
        n522, n521, n523, n524, n371, complb1, n190, complw1, n447, n469, n5, 
        n3, n4, n448, n467, n461, n372, n451, n458, n464, n273, n262, n259, 
        n256, n253, n228, n225, n239, n361, n356, n331, n295, n275, n281, n278, 
        n264, n261, n258, n254, n255, n241, n341, n328, n325, n338, n362, n357, 
        n352, n299, n289, n286, n292, n317, n322, n306, n314, n332, n296, n342, 
        n346, n329, n326, n339, n353, n300, n290, n287, n293, n318, n323, n307, 
        req_out_delayed, _25_net_, n529, n530, _24_net_, _26_net_, n142, 
        req_in_i, n186, n187, all_w, all_r, comp_basic, 
        \cg_all_w/__tmp99/loop , comp_wd, \Usze1/ni , \Usze1/nh , \Usze1/nl , 
        n2, \Usze0/ni , \Usze0/nh , \Usze0/nl , \Urnw/ni , \Urnw/nh , 
        \Urnw/nl , \Uerr/ni , \Uerr/nh , \Uerr/nl ;
    assign tc_wd_63 = tc_wd[63];
    assign tc_wd_62 = tc_wd[62];
    assign tc_wd_61 = tc_wd[61];
    assign tc_wd_60 = tc_wd[60];
    assign tc_wd_59 = tc_wd[59];
    assign tc_wd_58 = tc_wd[58];
    assign tc_wd_56 = tc_wd[56];
    assign tc_wd_55 = tc_wd[55];
    assign tc_wd_54 = tc_wd[54];
    assign tc_wd_53 = tc_wd[53];
    assign tc_wd_52 = tc_wd[52];
    assign tc_wd_51 = tc_wd[51];
    assign tc_wd_50 = tc_wd[50];
    assign tc_wd_49 = tc_wd[49];
    assign tc_wd_48 = tc_wd[48];
    assign tc_wd_47 = tc_wd[47];
    assign tc_wd_46 = tc_wd[46];
    assign tc_wd_45 = tc_wd[45];
    assign tc_wd_44 = tc_wd[44];
    assign tc_wd_43 = tc_wd[43];
    assign tc_wd_40 = tc_wd[40];
    assign tc_wd_39 = tc_wd[39];
    assign tc_wd_38 = tc_wd[38];
    assign tc_wd_36 = tc_wd[36];
    assign tc_wd_32 = tc_wd[32];
    assign tc_a_60 = tc_a[60];
    assign tc_a_58 = tc_a[58];
    assign ts_i[2] = 1'b0;
    assign ts_i[1] = 1'b0;
    assign ts_i[0] = 1'b0;
    assign adr_i[28] = tc_a_60;
    assign adr_i[26] = tc_a_58;
    assign dat_i[31] = tc_wd_63;
    assign dat_i[30] = tc_wd_62;
    assign dat_i[29] = tc_wd_61;
    assign dat_i[28] = tc_wd_60;
    assign dat_i[27] = tc_wd_59;
    assign dat_i[26] = tc_wd_58;
    assign dat_i[24] = tc_wd_56;
    assign dat_i[23] = tc_wd_55;
    assign dat_i[22] = tc_wd_54;
    assign dat_i[21] = tc_wd_53;
    assign dat_i[20] = tc_wd_52;
    assign dat_i[19] = tc_wd_51;
    assign dat_i[18] = tc_wd_50;
    assign dat_i[17] = tc_wd_49;
    assign dat_i[16] = tc_wd_48;
    assign dat_i[15] = tc_wd_47;
    assign dat_i[14] = tc_wd_46;
    assign dat_i[13] = tc_wd_45;
    assign dat_i[12] = tc_wd_44;
    assign dat_i[11] = tc_wd_43;
    assign dat_i[8] = tc_wd_40;
    assign dat_i[7] = tc_wd_39;
    assign dat_i[6] = tc_wd_38;
    assign dat_i[4] = tc_wd_36;
    assign dat_i[0] = tc_wd_32;
    assign prd_i = 1'b0;
    assign sel_i[3] = sel_i_3;
    assign sel_i[2] = sel_i_3;
    assign sel_i[0] = 1'b1;
    assign tc_ack = ack_in;
    assign ack_out = tr_ack;
    sr2dr_word_8 Urd ( .i(dat_o), .req(n1), .h(tr_rd[63:32]), .l(tr_rd[31:0])
         );
    inv_1 U3 ( .x(n334), .a(tc_a[7]) );
    inv_1 U5 ( .x(n311), .a(tc_a[21]) );
    and2_1 U6 ( .x(n129), .a(n309), .b(n310) );
    inv_1 U7 ( .x(n309), .a(tc_a[6]) );
    inv_1 U9 ( .x(n315), .a(tc_itag[4]) );
    nand2_1 U10 ( .x(n348), .a(n349), .b(n350) );
    inv_1 U11 ( .x(n349), .a(tc_a[12]) );
    inv_1 U12 ( .x(n456), .a(n348) );
    inv_1 U13 ( .x(n336), .a(tc_a[30]) );
    inv_1 U14 ( .x(n457), .a(n345) );
    inv_1 U15 ( .x(n303), .a(tc_a[8]) );
    nand3_1 U16 ( .x(n505), .a(n193), .b(n476), .c(n479) );
    inv_1 U17 ( .x(n229), .a(tc_wd[5]) );
    inv_1 U18 ( .x(n226), .a(tc_wd[3]) );
    inv_1 U19 ( .x(n257), .a(tc_wd[16]) );
    inv_1 U20 ( .x(n263), .a(tc_wd[21]) );
    inv_1 U21 ( .x(n260), .a(tc_wd[19]) );
    nand2_1 U22 ( .x(n268), .a(n269), .b(n270) );
    inv_1 U23 ( .x(n269), .a(tc_wd[23]) );
    inv_1 U24 ( .x(n270), .a(tc_wd_55) );
    nand2_1 U25 ( .x(n265), .a(n266), .b(n267) );
    inv_1 U26 ( .x(n266), .a(tc_wd[20]) );
    inv_1 U27 ( .x(n277), .a(tc_wd[27]) );
    inv_1 U28 ( .x(n252), .a(tc_wd_47) );
    nand2_1 U29 ( .x(n248), .a(n249), .b(n250) );
    inv_1 U30 ( .x(n249), .a(tc_wd[12]) );
    nand2_1 U31 ( .x(n245), .a(n246), .b(n247) );
    inv_1 U32 ( .x(n246), .a(tc_wd[13]) );
    inv_1 U33 ( .x(n247), .a(tc_wd_45) );
    nand2_1 U34 ( .x(n242), .a(n243), .b(n244) );
    inv_1 U35 ( .x(n243), .a(tc_wd[11]) );
    nand2_1 U36 ( .x(n222), .a(n223), .b(n224) );
    inv_1 U37 ( .x(n223), .a(tc_wd[0]) );
    inv_1 U38 ( .x(n220), .a(tc_wd[1]) );
    nand2_1 U39 ( .x(n234), .a(n235), .b(n236) );
    inv_1 U40 ( .x(n235), .a(tc_wd[7]) );
    nand2_1 U41 ( .x(n231), .a(n232), .b(n233) );
    inv_1 U42 ( .x(n232), .a(tc_wd[4]) );
    nand2_1 U43 ( .x(n205), .a(n206), .b(n207) );
    inv_1 U44 ( .x(n206), .a(tc_wd[18]) );
    inv_1 U45 ( .x(n203), .a(tc_wd[10]) );
    nand2_1 U46 ( .x(n199), .a(n200), .b(n201) );
    inv_1 U47 ( .x(n200), .a(tc_wd[6]) );
    inv_1 U48 ( .x(n197), .a(tc_wd[2]) );
    inv_1 U49 ( .x(n218), .a(tc_wd_46) );
    nand2_1 U50 ( .x(n214), .a(n215), .b(n216) );
    inv_1 U51 ( .x(n215), .a(tc_wd[30]) );
    nand2_1 U52 ( .x(n211), .a(n212), .b(n213) );
    inv_1 U53 ( .x(n213), .a(tc_wd_58) );
    nand2_1 U54 ( .x(n208), .a(n209), .b(n210) );
    inv_1 U55 ( .x(n209), .a(tc_wd[22]) );
    inv_1 U56 ( .x(n374), .a(tc_rnw[0]) );
    inv_1 U57 ( .x(n375), .a(tc_rnw[1]) );
    inv_1 U58 ( .x(n368), .a(tc_a[18]) );
    inv_1 U59 ( .x(n244), .a(tc_wd_43) );
    inv_1 U60 ( .x(n251), .a(tc_wd[15]) );
    inv_1 U61 ( .x(n250), .a(tc_wd_44) );
    inv_1 U62 ( .x(n280), .a(tc_wd[29]) );
    inv_1 U63 ( .x(n267), .a(tc_wd_52) );
    inv_1 U64 ( .x(n274), .a(tc_wd[24]) );
    inv_1 U65 ( .x(n271), .a(tc_wd[25]) );
    inv_1 U66 ( .x(n212), .a(tc_wd[26]) );
    inv_1 U67 ( .x(n210), .a(tc_wd_54) );
    inv_1 U68 ( .x(n216), .a(tc_wd_62) );
    inv_1 U69 ( .x(n201), .a(tc_wd_38) );
    inv_1 U70 ( .x(n427), .a(n196) );
    inv_1 U71 ( .x(n207), .a(tc_wd_50) );
    inv_1 U72 ( .x(n424), .a(n202) );
    inv_1 U73 ( .x(n236), .a(tc_wd_39) );
    inv_1 U74 ( .x(n233), .a(tc_wd_36) );
    inv_1 U75 ( .x(n240), .a(tc_wd[8]) );
    inv_1 U76 ( .x(n237), .a(tc_wd[9]) );
    inv_1 U77 ( .x(n224), .a(tc_wd_32) );
    inv_1 U78 ( .x(n413), .a(n219) );
    nand2_1 U79 ( .x(n421), .a(n418), .b(n416) );
    nand2_1 U80 ( .x(n428), .a(n425), .b(n422) );
    nand2_1 U81 ( .x(n414), .a(n411), .b(n408) );
    inv_1 U82 ( .x(n238), .a(tc_wd[41]) );
    inv_1 U83 ( .x(n272), .a(tc_wd[57]) );
    inv_1 U84 ( .x(n350), .a(tc_a[44]) );
    inv_1 U85 ( .x(n351), .a(tc_a[43]) );
    inv_1 U86 ( .x(n366), .a(tc_a[41]) );
    inv_1 U87 ( .x(n335), .a(tc_a[39]) );
    inv_1 U88 ( .x(n310), .a(tc_a[38]) );
    inv_1 U89 ( .x(n355), .a(tc_a[52]) );
    and3_1 U90 ( .x(tc_ok), .a(n531), .b(n532), .c(respond) );
    and2_1 U91 ( .x(tc_slow), .a(respond), .b(acc_o) );
    inv_1 U94 ( .x(n313), .a(tc_itag[5]) );
    and2_1 U95 ( .x(n121), .a(n334), .b(n335) );
    and2_1 U96 ( .x(n122), .a(n359), .b(n360) );
    and2_1 U97 ( .x(n123), .a(n336), .b(n337) );
    and2_1 U98 ( .x(n124), .a(n237), .b(n238) );
    and2_1 U99 ( .x(n125), .a(n251), .b(n252) );
    and2_1 U100 ( .x(n126), .a(n271), .b(n272) );
    and2_1 U101 ( .x(n127), .a(n217), .b(n218) );
    and2_1 U102 ( .x(n128), .a(n311), .b(n312) );
    nor2_1 U103 ( .x(n130), .a(tc_size[3]), .b(tc_size[2]) );
    nand2i_1 U105 ( .x(n284), .a(tc_wd[31]), .b(n285) );
    oa22_1 U106 ( .x(n449), .a(tc_a[27]), .b(tc_a[59]), .c(tc_a[54]), .d(tc_a
        [22]) );
    inv_1 U107 ( .x(n359), .a(tc_a[27]) );
    inv_1 U108 ( .x(n360), .a(tc_a[59]) );
    nand2i_1 U109 ( .x(n282), .a(tc_wd[28]), .b(n283) );
    nor2_1 U110 ( .x(n479), .a(tc_itag[0]), .b(tc_itag[5]) );
    nand4_1 U112 ( .x(n380), .a(n279), .b(n276), .c(n284), .d(n282) );
    aoi21_1 U113 ( .x(n425), .a(n200), .b(n201), .c(n427) );
    oa22_1 U114 ( .x(n397), .a(tc_wd[13]), .b(tc_wd_45), .c(tc_wd[11]), .d(
        tc_wd_43) );
    nor2_1 U115 ( .x(n454), .a(tc_a[20]), .b(tc_a[52]) );
    aoi21_1 U116 ( .x(n422), .a(n206), .b(n207), .c(n424) );
    oa22_1 U117 ( .x(n418), .a(tc_wd[26]), .b(tc_wd_58), .c(tc_wd[22]), .d(
        tc_wd_54) );
    oa22_1 U118 ( .x(n416), .a(tc_wd[14]), .b(tc_wd_46), .c(tc_wd[30]), .d(
        tc_wd_62) );
    inv_1 U119 ( .x(n217), .a(tc_wd[14]) );
    aoi22_1 U120 ( .x(n463), .a(n336), .b(n337), .c(n334), .d(n335) );
    nor2_1 U121 ( .x(n453), .a(tc_a[11]), .b(tc_a[43]) );
    oa22_1 U122 ( .x(n395), .a(tc_wd[15]), .b(tc_wd_47), .c(tc_wd[12]), .d(
        tc_wd_44) );
    oa22_1 U123 ( .x(n404), .a(tc_wd[7]), .b(tc_wd_39), .c(tc_wd[4]), .d(
        tc_wd_36) );
    oa22_1 U124 ( .x(n383), .a(tc_wd[23]), .b(tc_wd_55), .c(tc_wd[20]), .d(
        tc_wd_52) );
    aoi21_1 U125 ( .x(n411), .a(n223), .b(n224), .c(n413) );
    nor2_1 U126 ( .x(n443), .a(tc_a[49]), .b(tc_a[17]) );
    aoi22_1 U127 ( .x(n477), .a(n311), .b(n312), .c(n309), .d(n310) );
    oa21_1 U128 ( .x(n455), .a(tc_a[12]), .b(tc_a[44]), .c(n345) );
    inv_1 U129 ( .x(dat_i[5]), .a(n230) );
    inv_1 U130 ( .x(dat_i[9]), .a(n238) );
    inv_1 U131 ( .x(dat_i[25]), .a(n272) );
    buf_1 U132 ( .x(sel_i_3), .a(tc_size[3]) );
    buf_1 U133 ( .x(adr_i[16]), .a(tc_a[48]) );
    nor2_1 U134 ( .x(n135), .a(tc_a[14]), .b(tc_a[46]) );
    inv_1 U135 ( .x(n305), .a(tc_a[46]) );
    inv_1 U136 ( .x(n487), .a(n302) );
    nand2i_1 U137 ( .x(n445), .a(n446), .b(n442) );
    nor2_1 U138 ( .x(n136), .a(tc_a[29]), .b(tc_a[61]) );
    inv_1 U139 ( .x(n320), .a(tc_a[61]) );
    nand2_1 U140 ( .x(n400), .a(n397), .b(n395) );
    inv_1 U141 ( .x(n137), .a(n340) );
    inv_1 U142 ( .x(dat_i[2]), .a(n198) );
    nand2_1 U143 ( .x(n386), .a(n383), .b(n381) );
    nand3i_1 U144 ( .x(n478), .a(n479), .b(n477), .c(n475) );
    nand2_1 U145 ( .x(n407), .a(n404), .b(n402) );
    inv_1 U146 ( .x(dat_i[10]), .a(n204) );
    inv_1 U147 ( .x(dat_i[1]), .a(n221) );
    nor2_1 U148 ( .x(n141), .a(tc_a[3]), .b(tc_a[35]) );
    inv_1 U149 ( .x(n321), .a(tc_a[35]) );
    nor2_1 U151 ( .x(n483), .a(n484), .b(n485) );
    nor2_1 U152 ( .x(n480), .a(n474), .b(n478) );
    inv_1 U153 ( .x(dat_i[3]), .a(n227) );
    nor2_1 U154 ( .x(n188), .a(n517), .b(n525) );
    nand2_1 U155 ( .x(n180), .a(n401), .b(n387) );
    nor2_1 U156 ( .x(n401), .a(n394), .b(n400) );
    nor2_1 U157 ( .x(n387), .a(n380), .b(n386) );
    nor2_1 U158 ( .x(n481), .a(n482), .b(n135) );
    nor2_1 U159 ( .x(n491), .a(n195), .b(n492) );
    nor2_1 U160 ( .x(n195), .a(tc_size[1]), .b(tc_size[3]) );
    inv_1 U161 ( .x(adr_i[18]), .a(n369) );
    nand2_1 U162 ( .x(n181), .a(n429), .b(n415) );
    nor2_1 U163 ( .x(n429), .a(n421), .b(n428) );
    nor2_1 U164 ( .x(n415), .a(n407), .b(n414) );
    inv_1 U165 ( .x(adr_i[0]), .a(n324) );
    inv_1 U166 ( .x(n324), .a(tc_a[32]) );
    inv_1 U167 ( .x(sel_i[1]), .a(n130) );
    inv_1 U168 ( .x(st_i[2]), .a(n343) );
    inv_1 U169 ( .x(adr_i[9]), .a(n366) );
    inv_1 U170 ( .x(adr_i[24]), .a(n363) );
    inv_1 U171 ( .x(adr_i[19]), .a(n319) );
    inv_1 U172 ( .x(n319), .a(tc_a[51]) );
    inv_1 U173 ( .x(n369), .a(tc_a[50]) );
    inv_1 U174 ( .x(st_i[3]), .a(n344) );
    inv_1 U175 ( .x(adr_i[13]), .a(n354) );
    inv_1 U176 ( .x(adr_i[12]), .a(n350) );
    inv_1 U177 ( .x(adr_i[8]), .a(n304) );
    inv_1 U178 ( .x(n304), .a(tc_a[40]) );
    inv_1 U179 ( .x(adr_i[2]), .a(n330) );
    buf_1 U180 ( .x(adr_i[17]), .a(tc_a[49]) );
    nand2_1 U181 ( .x(n497), .a(n496), .b(n130) );
    inv_1 U182 ( .x(adr_i[10]), .a(n291) );
    and2_1 U183 ( .x(n438), .a(n373), .b(n367) );
    inv_1 U184 ( .x(n439), .a(n373) );
    inv_1 U185 ( .x(n440), .a(n367) );
    inv_1 U186 ( .x(adr_i[20]), .a(n355) );
    inv_1 U187 ( .x(adr_i[27]), .a(n360) );
    inv_1 U188 ( .x(adr_i[4]), .a(n333) );
    inv_1 U189 ( .x(adr_i[25]), .a(n308) );
    inv_1 U190 ( .x(adr_i[30]), .a(n337) );
    inv_1 U191 ( .x(adr_i[31]), .a(n297) );
    inv_1 U192 ( .x(n297), .a(tc_a[63]) );
    inv_1 U193 ( .x(adr_i[15]), .a(n347) );
    inv_1 U194 ( .x(adr_i[11]), .a(n351) );
    inv_1 U195 ( .x(adr_i[1]), .a(n301) );
    inv_1 U196 ( .x(n301), .a(tc_a[33]) );
    nand2_1 U197 ( .x(n503), .a(n499), .b(n502) );
    nor2_1 U198 ( .x(n499), .a(n497), .b(n498) );
    inv_1 U199 ( .x(adr_i[21]), .a(n312) );
    inv_1 U200 ( .x(n312), .a(tc_a[53]) );
    inv_1 U201 ( .x(seq_i), .a(n288) );
    inv_1 U202 ( .x(adr_i[5]), .a(n327) );
    inv_1 U203 ( .x(st_i[4]), .a(n316) );
    inv_1 U204 ( .x(n316), .a(tc_itag[9]) );
    inv_1 U205 ( .x(st_i[1]), .a(n298) );
    inv_1 U206 ( .x(adr_i[23]), .a(n294) );
    inv_1 U207 ( .x(adr_i[22]), .a(n358) );
    nand2_1 U208 ( .x(complb0), .a(n188), .b(n189) );
    nor2_1 U209 ( .x(n189), .a(n503), .b(n510) );
    inv_1 U210 ( .x(adr_i[29]), .a(n320) );
    inv_1 U211 ( .x(adr_i[7]), .a(n335) );
    inv_1 U212 ( .x(adr_i[14]), .a(n305) );
    inv_1 U213 ( .x(adr_i[6]), .a(n310) );
    inv_1 U214 ( .x(st_i[0]), .a(n313) );
    inv_1 U215 ( .x(adr_i[3]), .a(n321) );
    nand3_1 U218 ( .x(n507), .a(n192), .b(n136), .c(n473) );
    nand2_1 U219 ( .x(n508), .a(n471), .b(n141) );
    nor2_1 U220 ( .x(n488), .a(n489), .b(n490) );
    nand4_1 U222 ( .x(complw0), .a(n182), .b(n183), .c(n184), .d(n185) );
    nor2_1 U223 ( .x(n192), .a(tc_a_58), .b(tc_a[26]) );
    nor2_1 U224 ( .x(n193), .a(tc_a[48]), .b(tc_a[16]) );
    nand2_1 U225 ( .x(n364), .a(n365), .b(n366) );
    nand2_1 U226 ( .x(n394), .a(n391), .b(n388) );
    nand4_1 U227 ( .x(n430), .a(n423), .b(n424), .c(n426), .d(n427) );
    nand4_1 U228 ( .x(n431), .a(n127), .b(n417), .c(n419), .d(n420) );
    nor2_1 U229 ( .x(n185), .a(n430), .b(n431) );
    nand4_1 U230 ( .x(n432), .a(n409), .b(n410), .c(n412), .d(n413) );
    nand4_1 U231 ( .x(n433), .a(n403), .b(n124), .c(n405), .d(n406) );
    nor2_1 U232 ( .x(n184), .a(n432), .b(n433) );
    nand4_1 U233 ( .x(n434), .a(n125), .b(n396), .c(n398), .d(n399) );
    nand4_1 U234 ( .x(n435), .a(n389), .b(n390), .c(n392), .d(n393) );
    nor2_1 U235 ( .x(n183), .a(n434), .b(n435) );
    nand4_1 U236 ( .x(n436), .a(n382), .b(n126), .c(n384), .d(n385) );
    nand4_1 U237 ( .x(n437), .a(n376), .b(n377), .c(n378), .d(n379) );
    nor2_1 U238 ( .x(n182), .a(n436), .b(n437) );
    nand2_1 U239 ( .x(n441), .a(n438), .b(n370) );
    nor2_1 U240 ( .x(n442), .a(n443), .b(n444) );
    nor3_1 U241 ( .x(n470), .a(n471), .b(n136), .c(n141) );
    nor3_1 U242 ( .x(n472), .a(n473), .b(n192), .c(n193) );
    nand2_1 U243 ( .x(n474), .a(n472), .b(n470) );
    nor2_1 U244 ( .x(n475), .a(n476), .b(n194) );
    nand3i_1 U245 ( .x(n486), .a(n487), .b(n481), .c(n483) );
    nand3i_1 U246 ( .x(n493), .a(n494), .b(n488), .c(n491) );
    nor2_1 U247 ( .x(n495), .a(n493), .b(n486) );
    nand2_1 U248 ( .x(n191), .a(n495), .b(n480) );
    nand3_1 U249 ( .x(n498), .a(n489), .b(n492), .c(n490) );
    nand3_1 U250 ( .x(n500), .a(n485), .b(n494), .c(n484) );
    nand2_1 U251 ( .x(n501), .a(n135), .b(n487) );
    nor2_1 U252 ( .x(n502), .a(n500), .b(n501) );
    nand3_1 U253 ( .x(n504), .a(n128), .b(n482), .c(n129) );
    nor2_1 U254 ( .x(n506), .a(n504), .b(n505) );
    nor2_1 U255 ( .x(n509), .a(n507), .b(n508) );
    nand2_1 U256 ( .x(n510), .a(n509), .b(n506) );
    nand3_1 U257 ( .x(n511), .a(n465), .b(n466), .c(n468) );
    nand3_1 U258 ( .x(n512), .a(n123), .b(n121), .c(n460) );
    nor2_1 U259 ( .x(n513), .a(n511), .b(n512) );
    nand3_1 U260 ( .x(n514), .a(n462), .b(n459), .c(n457) );
    nand2_1 U261 ( .x(n515), .a(n453), .b(n456) );
    nor2_1 U262 ( .x(n516), .a(n514), .b(n515) );
    nand2_1 U263 ( .x(n517), .a(n516), .b(n513) );
    nand2_1 U264 ( .x(n518), .a(n454), .b(n452) );
    nor2i_1 U265 ( .x(n519), .a(n450), .b(n518) );
    nand2_1 U266 ( .x(n520), .a(n444), .b(n122) );
    nor2i_1 U267 ( .x(n522), .a(n446), .b(n521) );
    nand2_1 U268 ( .x(n523), .a(n439), .b(n524) );
    inv_1 U270 ( .x(n365), .a(tc_a[9]) );
    inv_1 U271 ( .x(n371), .a(tc_a_60) );
    inv_1 U272 ( .x(n446), .a(n364) );
    nor2_1 U273 ( .x(complb1), .a(n190), .b(n191) );
    nor2_1 U274 ( .x(complw1), .a(n180), .b(n181) );
    nand3i_1 U276 ( .x(n190), .a(n441), .b(n447), .c(n469) );
    and4_1 U277 ( .x(n5), .a(n3), .b(n4), .c(n519), .d(n522) );
    inv_1 U216 ( .x(n3), .a(n520) );
    inv_1 U217 ( .x(n4), .a(n523) );
    inv_1 U428 ( .x(n525), .a(n5) );
    nor2_1 U278 ( .x(n447), .a(n448), .b(n445) );
    nor2_1 U279 ( .x(n469), .a(n467), .b(n461) );
    nand2_1 U280 ( .x(n370), .a(n371), .b(n372) );
    nand3i_1 U281 ( .x(n448), .a(n454), .b(n449), .c(n451) );
    nand3i_1 U282 ( .x(n461), .a(n462), .b(n455), .c(n458) );
    nand3i_1 U283 ( .x(n467), .a(n468), .b(n463), .c(n464) );
    inv_1 U284 ( .x(n382), .a(n273) );
    inv_1 U285 ( .x(n384), .a(n268) );
    inv_1 U286 ( .x(n385), .a(n265) );
    inv_1 U287 ( .x(n376), .a(n284) );
    inv_1 U288 ( .x(n377), .a(n282) );
    inv_1 U289 ( .x(n378), .a(n279) );
    inv_1 U290 ( .x(n379), .a(n276) );
    inv_1 U291 ( .x(n396), .a(n248) );
    inv_1 U292 ( .x(n398), .a(n245) );
    inv_1 U293 ( .x(n399), .a(n242) );
    inv_1 U294 ( .x(n389), .a(n262) );
    inv_1 U295 ( .x(n390), .a(n259) );
    inv_1 U296 ( .x(n392), .a(n256) );
    inv_1 U297 ( .x(n393), .a(n253) );
    inv_1 U298 ( .x(n409), .a(n228) );
    inv_1 U299 ( .x(n410), .a(n225) );
    inv_1 U300 ( .x(n412), .a(n222) );
    inv_1 U301 ( .x(n403), .a(n239) );
    inv_1 U302 ( .x(n405), .a(n234) );
    inv_1 U303 ( .x(n406), .a(n231) );
    inv_1 U304 ( .x(n423), .a(n205) );
    inv_1 U305 ( .x(n426), .a(n199) );
    inv_1 U306 ( .x(n417), .a(n214) );
    inv_1 U307 ( .x(n419), .a(n211) );
    inv_1 U308 ( .x(n420), .a(n208) );
    inv_1 U309 ( .x(n444), .a(n361) );
    inv_1 U310 ( .x(n524), .a(n370) );
    inv_1 U311 ( .x(n450), .a(n356) );
    nand2_1 U312 ( .x(n521), .a(n443), .b(n440) );
    inv_1 U313 ( .x(n372), .a(tc_a[28]) );
    nor2_1 U314 ( .x(n451), .a(n452), .b(n453) );
    nor2_1 U315 ( .x(n458), .a(n459), .b(n460) );
    inv_1 U316 ( .x(n468), .a(n331) );
    nor2_1 U317 ( .x(n464), .a(n465), .b(n466) );
    inv_1 U318 ( .x(n494), .a(n295) );
    nand2_1 U319 ( .x(n273), .a(n274), .b(n275) );
    nand2_1 U320 ( .x(n279), .a(n280), .b(n281) );
    nand2_1 U321 ( .x(n276), .a(n277), .b(n278) );
    nand2_1 U322 ( .x(n262), .a(n263), .b(n264) );
    nand2_1 U323 ( .x(n259), .a(n260), .b(n261) );
    nand2_1 U324 ( .x(n256), .a(n257), .b(n258) );
    nand2_1 U325 ( .x(n253), .a(n254), .b(n255) );
    nand2_1 U326 ( .x(n228), .a(n229), .b(n230) );
    nand2_1 U327 ( .x(n225), .a(n226), .b(n227) );
    nand2_1 U328 ( .x(n219), .a(n220), .b(n221) );
    nand2_1 U329 ( .x(n239), .a(n240), .b(n241) );
    nand2_1 U330 ( .x(n202), .a(n203), .b(n204) );
    nand2_1 U331 ( .x(n196), .a(n197), .b(n198) );
    nor2_1 U332 ( .x(n391), .a(n392), .b(n393) );
    nor2_1 U333 ( .x(n388), .a(n389), .b(n390) );
    nor2_1 U334 ( .x(n381), .a(n382), .b(n126) );
    nor2_1 U335 ( .x(n402), .a(n403), .b(n124) );
    nor2_1 U336 ( .x(n408), .a(n409), .b(n410) );
    inv_1 U337 ( .x(n459), .a(n341) );
    inv_1 U338 ( .x(n465), .a(n328) );
    inv_1 U339 ( .x(n466), .a(n325) );
    inv_1 U340 ( .x(n460), .a(n338) );
    nand2_1 U341 ( .x(n361), .a(n362), .b(n363) );
    nand2_1 U342 ( .x(n373), .a(n374), .b(n375) );
    nand2_1 U343 ( .x(n356), .a(n358), .b(n357) );
    inv_1 U344 ( .x(n452), .a(n352) );
    inv_1 U345 ( .x(n484), .a(n299) );
    inv_1 U346 ( .x(n489), .a(n289) );
    inv_1 U347 ( .x(n492), .a(n286) );
    inv_1 U348 ( .x(n490), .a(n292) );
    inv_1 U349 ( .x(n473), .a(n317) );
    inv_1 U350 ( .x(n471), .a(n322) );
    inv_1 U351 ( .x(n482), .a(n306) );
    inv_1 U352 ( .x(n476), .a(n314) );
    nand2_1 U353 ( .x(n367), .a(n368), .b(n369) );
    nand2_1 U354 ( .x(n331), .a(n332), .b(n333) );
    nand2_1 U355 ( .x(n302), .a(n303), .b(n304) );
    nand2_1 U356 ( .x(n295), .a(n296), .b(n297) );
    inv_1 U357 ( .x(n275), .a(tc_wd_56) );
    inv_1 U358 ( .x(n285), .a(tc_wd_63) );
    inv_1 U359 ( .x(n283), .a(tc_wd_60) );
    inv_1 U360 ( .x(n281), .a(tc_wd_61) );
    inv_1 U361 ( .x(n278), .a(tc_wd_59) );
    inv_1 U362 ( .x(n264), .a(tc_wd_53) );
    inv_1 U363 ( .x(n261), .a(tc_wd_51) );
    inv_1 U364 ( .x(n258), .a(tc_wd_48) );
    inv_1 U365 ( .x(n254), .a(tc_wd[17]) );
    inv_1 U366 ( .x(n255), .a(tc_wd_49) );
    inv_1 U367 ( .x(n230), .a(tc_wd[37]) );
    inv_1 U368 ( .x(n227), .a(tc_wd[35]) );
    inv_1 U369 ( .x(n221), .a(tc_wd[33]) );
    inv_1 U370 ( .x(n241), .a(tc_wd_40) );
    inv_1 U371 ( .x(n204), .a(tc_wd[42]) );
    inv_1 U372 ( .x(n198), .a(tc_wd[34]) );
    nand2_1 U373 ( .x(n341), .a(n342), .b(n343) );
    nand2_1 U374 ( .x(n345), .a(n347), .b(n346) );
    nand2_1 U375 ( .x(n328), .a(n329), .b(n330) );
    nand2_1 U376 ( .x(n325), .a(n326), .b(n327) );
    nand2_1 U377 ( .x(n338), .a(n340), .b(n339) );
    inv_1 U378 ( .x(n362), .a(tc_a[24]) );
    inv_1 U379 ( .x(n363), .a(tc_a[56]) );
    inv_1 U380 ( .x(n357), .a(tc_a[22]) );
    inv_1 U381 ( .x(n358), .a(tc_a[54]) );
    nand2_1 U382 ( .x(n352), .a(n353), .b(n354) );
    nand2_1 U383 ( .x(n299), .a(n300), .b(n301) );
    nand2_1 U384 ( .x(n289), .a(n290), .b(n291) );
    nand2_1 U385 ( .x(n286), .a(n287), .b(n288) );
    nand2_1 U386 ( .x(n292), .a(n293), .b(n294) );
    nand2_1 U387 ( .x(n317), .a(n318), .b(n319) );
    nand2_1 U388 ( .x(n322), .a(n323), .b(n324) );
    nand2_1 U389 ( .x(n306), .a(n307), .b(n308) );
    nand2_1 U390 ( .x(n314), .a(n315), .b(n316) );
    inv_1 U391 ( .x(n332), .a(tc_a[4]) );
    inv_1 U392 ( .x(n333), .a(tc_a[36]) );
    inv_1 U393 ( .x(n296), .a(tc_a[31]) );
    inv_1 U394 ( .x(n342), .a(tc_itag[2]) );
    inv_1 U395 ( .x(n343), .a(tc_itag[7]) );
    inv_1 U396 ( .x(n346), .a(tc_a[15]) );
    inv_1 U397 ( .x(n347), .a(tc_a[47]) );
    inv_1 U398 ( .x(n329), .a(tc_a[2]) );
    inv_1 U399 ( .x(n330), .a(tc_a[34]) );
    inv_1 U400 ( .x(n326), .a(tc_a[5]) );
    inv_1 U401 ( .x(n327), .a(tc_a[37]) );
    inv_1 U402 ( .x(n337), .a(tc_a[62]) );
    inv_1 U403 ( .x(n339), .a(tc_lock[0]) );
    inv_1 U404 ( .x(n340), .a(tc_lock[1]) );
    inv_1 U405 ( .x(n353), .a(tc_a[13]) );
    inv_1 U406 ( .x(n354), .a(tc_a[45]) );
    inv_1 U407 ( .x(n300), .a(tc_a[1]) );
    inv_1 U408 ( .x(n290), .a(tc_a[10]) );
    inv_1 U409 ( .x(n291), .a(tc_a[42]) );
    inv_1 U410 ( .x(n287), .a(tc_seq[0]) );
    inv_1 U411 ( .x(n288), .a(tc_seq[1]) );
    inv_1 U412 ( .x(n293), .a(tc_a[23]) );
    inv_1 U413 ( .x(n294), .a(tc_a[55]) );
    inv_1 U414 ( .x(n318), .a(tc_a[19]) );
    inv_1 U415 ( .x(n323), .a(tc_a[0]) );
    inv_1 U416 ( .x(n307), .a(tc_a[25]) );
    inv_1 U417 ( .x(n308), .a(tc_a[57]) );
    buf_1 U418 ( .x(we_i), .a(tc_rnw[0]) );
    matched_delay_cp2slave_resp_dmem U419 ( .x(req_out_delayed), .a(req_out)
         );
    and4_1 U420 ( .x(_25_net_), .a(sel_o[0]), .b(sel_o[1]), .c(n529), .d(n530)
         );
    inv_1 U421 ( .x(_24_net_), .a(we_i) );
    and2_1 U422 ( .x(tc_defer), .a(rty_o), .b(respond) );
    and4_1 U423 ( .x(_26_net_), .a(sel_o[0]), .b(sel_o[1]), .c(sel_o[3]), .d(
        sel_o[2]) );
    inv_1 U424 ( .x(n532), .a(acc_o) );
    inv_1 U425 ( .x(n531), .a(rty_o) );
    inv_1 U426 ( .x(n529), .a(sel_o[2]) );
    inv_1 U427 ( .x(n530), .a(sel_o[3]) );
    buf_1 U150 ( .x(n142), .a(req_in_i) );
    matched_delay_cp2slave_comdmem matchDelCom ( .x(req_in), .a(req_in_i) );
    nand2_1 U275 ( .x(req_in_i), .a(n186), .b(n187) );
    inv_1 U221 ( .x(n186), .a(all_w) );
    inv_1 U269 ( .x(n187), .a(all_r) );
    dffp_1 mult_i_reg ( .q(mult_i), .d(n137), .ck(n142) );
    ao222_1 \cg_respond/__tmp99/U1  ( .x(respond), .a(req_out), .b(tc_ack), 
        .c(req_out), .d(respond), .e(tc_ack), .f(respond) );
    oa21_1 \cg_all_r/__tmp99/U1  ( .x(all_r), .a(tc_rnw[1]), .b(all_r), .c(
        comp_basic) );
    ao31_1 \cg_all_w/__tmp99/aoi  ( .x(\cg_all_w/__tmp99/loop ), .a(comp_basic
        ), .b(comp_wd), .c(we_i), .d(all_w) );
    oa21_1 \cg_all_w/__tmp99/outGate  ( .x(all_w), .a(comp_basic), .b(comp_wd), 
        .c(\cg_all_w/__tmp99/loop ) );
    ao222_1 \cg_wd/__tmp99/U1  ( .x(comp_wd), .a(complw0), .b(complw1), .c(
        complw0), .d(comp_wd), .e(complw1), .f(comp_wd) );
    ao222_1 \cg_basic/__tmp99/U1  ( .x(comp_basic), .a(complb0), .b(complb1), 
        .c(complb0), .d(comp_basic), .e(complb1), .f(comp_basic) );
    inv_1 \Usze1/Uii  ( .x(\Usze1/ni ), .a(_26_net_) );
    inv_1 \Usze1/Uih  ( .x(\Usze1/nh ), .a(tr_size[3]) );
    inv_1 \Usze1/Uil  ( .x(\Usze1/nl ), .a(tr_size[1]) );
    ao23_1 \Usze1/Ucl/U1/U1  ( .x(tr_size[1]), .a(n2), .b(tr_size[1]), .c(n1), 
        .d(\Usze1/ni ), .e(\Usze1/nh ) );
    ao23_1 \Usze1/Uch/U1/U1  ( .x(tr_size[3]), .a(n1), .b(tr_size[3]), .c(n1), 
        .d(_26_net_), .e(\Usze1/nl ) );
    inv_1 \Usze0/Uii  ( .x(\Usze0/ni ), .a(_25_net_) );
    inv_1 \Usze0/Uih  ( .x(\Usze0/nh ), .a(tr_size[2]) );
    inv_1 \Usze0/Uil  ( .x(\Usze0/nl ), .a(tr_size[0]) );
    ao23_1 \Usze0/Ucl/U1/U1  ( .x(tr_size[0]), .a(n2), .b(tr_size[0]), .c(n1), 
        .d(\Usze0/ni ), .e(\Usze0/nh ) );
    ao23_1 \Usze0/Uch/U1/U1  ( .x(tr_size[2]), .a(n2), .b(tr_size[2]), .c(n1), 
        .d(_25_net_), .e(\Usze0/nl ) );
    inv_1 \Urnw/Uii  ( .x(\Urnw/ni ), .a(_24_net_) );
    inv_1 \Urnw/Uih  ( .x(\Urnw/nh ), .a(tr_rnw[1]) );
    inv_1 \Urnw/Uil  ( .x(\Urnw/nl ), .a(tr_rnw[0]) );
    ao23_1 \Urnw/Ucl/U1/U1  ( .x(tr_rnw[0]), .a(n1), .b(tr_rnw[0]), .c(n1), 
        .d(\Urnw/ni ), .e(\Urnw/nh ) );
    ao23_1 \Urnw/Uch/U1/U1  ( .x(tr_rnw[1]), .a(n1), .b(tr_rnw[1]), .c(n1), 
        .d(_24_net_), .e(\Urnw/nl ) );
    inv_1 \Uerr/Uii  ( .x(\Uerr/ni ), .a(err_o) );
    inv_1 \Uerr/Uih  ( .x(\Uerr/nh ), .a(tr_err[1]) );
    inv_1 \Uerr/Uil  ( .x(\Uerr/nl ), .a(tr_err[0]) );
    ao23_1 \Uerr/Ucl/U1/U1  ( .x(tr_err[0]), .a(n1), .b(tr_err[0]), .c(n1), 
        .d(\Uerr/ni ), .e(\Uerr/nh ) );
    ao23_1 \Uerr/Uch/U1/U1  ( .x(tr_err[1]), .a(n1), .b(tr_err[1]), .c(n1), 
        .d(err_o), .e(\Uerr/nl ) );
    inv_0 U1 ( .x(n298), .a(tc_itag[6]) );
    nor2_0 U2 ( .x(n485), .a(tc_itag[1]), .b(tc_itag[6]) );
    inv_0 U4 ( .x(n344), .a(tc_itag[8]) );
    nor2_0 U8 ( .x(n462), .a(tc_itag[3]), .b(tc_itag[8]) );
    nor2_0 U92 ( .x(n496), .a(tc_size[0]), .b(tc_size[1]) );
    nor2_0 U93 ( .x(n194), .a(tc_size[0]), .b(tc_size[2]) );
    buf_16 U104 ( .x(n1), .a(req_out_delayed) );
    buf_16 U111 ( .x(n2), .a(req_out_delayed) );
endmodule


module slave_if_dmem ( nReset, sc_req, sc_we, sc_mult, sc_seq, sc_prd, sc_ts, 
    sc_st, sc_sel, sc_adr, sc_dat, sc_ack, sr_req, sr_err, sr_rty, sr_acc, 
    sr_mult, sr_ts, sr_rt, sr_sel, sr_dat, sr_ack, chaincommand, 
    nchaincommandack, chainresponse, nchainresponseack, e_dp, e_ip, e_tic, 
    r_dp, r_ip, r_tic );
output [2:0] sc_ts;
output [4:0] sc_st;
output [3:0] sc_sel;
output [31:0] sc_adr;
output [31:0] sc_dat;
input  [2:0] sr_ts;
input  [4:0] sr_rt;
input  [3:0] sr_sel;
input  [31:0] sr_dat;
input  [4:0] chaincommand;
output [4:0] chainresponse;
input  [2:0] e_dp;
input  [2:0] e_ip;
input  [2:0] e_tic;
input  [2:0] r_dp;
input  [2:0] r_ip;
input  [2:0] r_tic;
input  nReset, sc_ack, sr_req, sr_err, sr_rty, sr_acc, sr_mult, 
    nchainresponseack;
output sc_req, sc_we, sc_mult, sc_seq, sc_prd, sr_ack, nchaincommandack;
    wire nroute_ack, rt_ack, routetx_req, ct_ack, ct_defer, ct_slow, ct_ok, 
        routetx_ack, \route[4] , \route[1] , \route[0] , \rt_rd[63] , 
        \rt_rd[62] , \rt_rd[61] , \rt_rd[60] , \rt_rd[59] , \rt_rd[58] , 
        \rt_rd[57] , \rt_rd[56] , \rt_rd[55] , \rt_rd[54] , \rt_rd[53] , 
        \rt_rd[52] , \rt_rd[51] , \rt_rd[50] , \rt_rd[49] , \rt_rd[48] , 
        \rt_rd[47] , \rt_rd[46] , \rt_rd[45] , \rt_rd[44] , \rt_rd[43] , 
        \rt_rd[42] , \rt_rd[41] , \rt_rd[40] , \rt_rd[39] , \rt_rd[38] , 
        \rt_rd[37] , \rt_rd[36] , \rt_rd[35] , \rt_rd[34] , \rt_rd[33] , 
        \rt_rd[32] , \rt_rd[31] , \rt_rd[30] , \rt_rd[29] , \rt_rd[28] , 
        \rt_rd[27] , \rt_rd[26] , \rt_rd[25] , \rt_rd[24] , \rt_rd[23] , 
        \rt_rd[22] , \rt_rd[21] , \rt_rd[20] , \rt_rd[19] , \rt_rd[18] , 
        \rt_rd[17] , \rt_rd[16] , \rt_rd[15] , \rt_rd[14] , \rt_rd[13] , 
        \rt_rd[12] , \rt_rd[11] , \rt_rd[10] , \rt_rd[9] , \rt_rd[8] , 
        \rt_rd[7] , \rt_rd[6] , \rt_rd[5] , \rt_rd[4] , \rt_rd[3] , \rt_rd[2] , 
        \rt_rd[1] , \rt_rd[0] , \rt_err[1] , \rt_err[0] , \ct_wd[63] , 
        \ct_wd[62] , \ct_wd[61] , \ct_wd[60] , \ct_wd[59] , \ct_wd[58] , 
        \ct_wd[57] , \ct_wd[56] , \ct_wd[55] , \ct_wd[54] , \ct_wd[53] , 
        \ct_wd[52] , \ct_wd[51] , \ct_wd[50] , \ct_wd[49] , \ct_wd[48] , 
        \ct_wd[47] , \ct_wd[46] , \ct_wd[45] , \ct_wd[44] , \ct_wd[43] , 
        \ct_wd[42] , \ct_wd[41] , \ct_wd[40] , \ct_wd[39] , \ct_wd[38] , 
        \ct_wd[37] , \ct_wd[36] , \ct_wd[35] , \ct_wd[34] , \ct_wd[33] , 
        \ct_wd[32] , \ct_wd[31] , \ct_wd[30] , \ct_wd[29] , \ct_wd[28] , 
        \ct_wd[27] , \ct_wd[26] , \ct_wd[25] , \ct_wd[24] , \ct_wd[23] , 
        \ct_wd[22] , \ct_wd[21] , \ct_wd[20] , \ct_wd[19] , \ct_wd[18] , 
        \ct_wd[17] , \ct_wd[16] , \ct_wd[15] , \ct_wd[14] , \ct_wd[13] , 
        \ct_wd[12] , \ct_wd[11] , \ct_wd[10] , \ct_wd[9] , \ct_wd[8] , 
        \ct_wd[7] , \ct_wd[6] , \ct_wd[5] , \ct_wd[4] , \ct_wd[3] , \ct_wd[2] , 
        \ct_wd[1] , \ct_wd[0] , \tag_l[4] , \tag_l[3] , \tag_l[2] , \tag_l[1] , 
        \tag_l[0] , \tag_h[4] , \tag_h[3] , \tag_h[2] , \tag_h[1] , \tag_h[0] , 
        \ct_seq[1] , \ct_seq[0] , \ct_lock[1] , \ct_lock[0] , \ct_itag[9] , 
        \ct_itag[8] , \ct_itag[7] , \ct_itag[6] , \ct_itag[5] , \ct_itag[4] , 
        \ct_itag[3] , \ct_itag[2] , \ct_itag[1] , \ct_itag[0] , \ct_size[3] , 
        \ct_size[2] , \ct_size[1] , \ct_size[0] , \ct_rnw[1] , \ct_rnw[0] , 
        \ct_a[63] , \ct_a[62] , \ct_a[61] , \ct_a[60] , \ct_a[59] , \ct_a[58] , 
        \ct_a[57] , \ct_a[56] , \ct_a[55] , \ct_a[54] , \ct_a[53] , \ct_a[52] , 
        \ct_a[51] , \ct_a[50] , \ct_a[49] , \ct_a[48] , \ct_a[47] , \ct_a[46] , 
        \ct_a[45] , \ct_a[44] , \ct_a[43] , \ct_a[42] , \ct_a[41] , \ct_a[40] , 
        \ct_a[39] , \ct_a[38] , \ct_a[37] , \ct_a[36] , \ct_a[35] , \ct_a[34] , 
        \ct_a[33] , \ct_a[32] , \ct_a[31] , \ct_a[30] , \ct_a[29] , \ct_a[28] , 
        \ct_a[27] , \ct_a[26] , \ct_a[25] , \ct_a[24] , \ct_a[23] , \ct_a[22] , 
        \ct_a[21] , \ct_a[20] , \ct_a[19] , \ct_a[18] , \ct_a[17] , \ct_a[16] , 
        \ct_a[15] , \ct_a[14] , \ct_a[13] , \ct_a[12] , \ct_a[11] , \ct_a[10] , 
        \ct_a[9] , \ct_a[8] , \ct_a[7] , \ct_a[6] , \ct_a[5] , \ct_a[4] , 
        \ct_a[3] , \ct_a[2] , \ct_a[1] , \ct_a[0] , \rl[2] , \rl[1] , \rl[0] , 
        \rh[2] , \rh[1] , SYNOPSYS_UNCONNECTED_2, \el[2] , \el[1] , \el[0] , 
        SYNOPSYS_UNCONNECTED_1, \eh[1] , \eh[0] , SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4, reset, SYNOPSYS_UNCONNECTED_5;
    assign sc_prd = 1'b0;
    assign sc_ts[2] = 1'b0;
    assign sc_ts[1] = 1'b0;
    assign sc_ts[0] = 1'b0;
    assign sc_sel[0] = 1'b1;
    target_dmem tg ( .addr({\ct_a[63] , \ct_a[62] , \ct_a[61] , \ct_a[60] , 
        \ct_a[59] , \ct_a[58] , \ct_a[57] , \ct_a[56] , \ct_a[55] , \ct_a[54] , 
        \ct_a[53] , \ct_a[52] , \ct_a[51] , \ct_a[50] , \ct_a[49] , \ct_a[48] , 
        \ct_a[47] , \ct_a[46] , \ct_a[45] , \ct_a[44] , \ct_a[43] , \ct_a[42] , 
        \ct_a[41] , \ct_a[40] , \ct_a[39] , \ct_a[38] , \ct_a[37] , \ct_a[36] , 
        \ct_a[35] , \ct_a[34] , \ct_a[33] , \ct_a[32] , \ct_a[31] , \ct_a[30] , 
        \ct_a[29] , \ct_a[28] , \ct_a[27] , \ct_a[26] , \ct_a[25] , \ct_a[24] , 
        \ct_a[23] , \ct_a[22] , \ct_a[21] , \ct_a[20] , \ct_a[19] , \ct_a[18] , 
        \ct_a[17] , \ct_a[16] , \ct_a[15] , \ct_a[14] , \ct_a[13] , \ct_a[12] , 
        \ct_a[11] , \ct_a[10] , \ct_a[9] , \ct_a[8] , \ct_a[7] , \ct_a[6] , 
        \ct_a[5] , \ct_a[4] , \ct_a[3] , \ct_a[2] , \ct_a[1] , \ct_a[0] }), 
        .chainresponse(chainresponse), .crnw({\ct_rnw[1] , \ct_rnw[0] }), 
        .csize({\ct_size[3] , \ct_size[2] , \ct_size[1] , \ct_size[0] }), 
        .ctag({\ct_itag[9] , \ct_itag[8] , \ct_itag[7] , \ct_itag[6] , 
        \ct_itag[5] , \ct_itag[4] , \ct_itag[3] , \ct_itag[2] , \ct_itag[1] , 
        \ct_itag[0] }), .lock({\ct_lock[1] , \ct_lock[0] }), 
        .nchaincommandack(nchaincommandack), .nrouteack(nroute_ack), .rack(
        rt_ack), .routetxreq(routetx_req), .seq({\ct_seq[1] , \ct_seq[0] }), 
        .tag_h({\tag_h[4] , \tag_h[3] , \tag_h[2] , \tag_h[1] , \tag_h[0] }), 
        .tag_l({\tag_l[4] , \tag_l[3] , \tag_l[2] , \tag_l[1] , \tag_l[0] }), 
        .wd({\ct_wd[63] , \ct_wd[62] , \ct_wd[61] , \ct_wd[60] , \ct_wd[59] , 
        \ct_wd[58] , \ct_wd[57] , \ct_wd[56] , \ct_wd[55] , \ct_wd[54] , 
        \ct_wd[53] , \ct_wd[52] , \ct_wd[51] , \ct_wd[50] , \ct_wd[49] , 
        \ct_wd[48] , \ct_wd[47] , \ct_wd[46] , \ct_wd[45] , \ct_wd[44] , 
        \ct_wd[43] , \ct_wd[42] , \ct_wd[41] , \ct_wd[40] , \ct_wd[39] , 
        \ct_wd[38] , \ct_wd[37] , \ct_wd[36] , \ct_wd[35] , \ct_wd[34] , 
        \ct_wd[33] , \ct_wd[32] , \ct_wd[31] , \ct_wd[30] , \ct_wd[29] , 
        \ct_wd[28] , \ct_wd[27] , \ct_wd[26] , \ct_wd[25] , \ct_wd[24] , 
        \ct_wd[23] , \ct_wd[22] , \ct_wd[21] , \ct_wd[20] , \ct_wd[19] , 
        \ct_wd[18] , \ct_wd[17] , \ct_wd[16] , \ct_wd[15] , \ct_wd[14] , 
        \ct_wd[13] , \ct_wd[12] , \ct_wd[11] , \ct_wd[10] , \ct_wd[9] , 
        \ct_wd[8] , \ct_wd[7] , \ct_wd[6] , \ct_wd[5] , \ct_wd[4] , \ct_wd[3] , 
        \ct_wd[2] , \ct_wd[1] , \ct_wd[0] }), .cack(ct_ack), .cdefer(ct_defer), 
        .chaincommand(chaincommand), .cndefer(ct_slow), .cok(ct_ok), .err({
        \rt_err[1] , \rt_err[0] }), .nReset(nReset), .nchainresponseack(
        nchainresponseack), .rd({\rt_rd[63] , \rt_rd[62] , \rt_rd[61] , 
        \rt_rd[60] , \rt_rd[59] , \rt_rd[58] , \rt_rd[57] , \rt_rd[56] , 
        \rt_rd[55] , \rt_rd[54] , \rt_rd[53] , \rt_rd[52] , \rt_rd[51] , 
        \rt_rd[50] , \rt_rd[49] , \rt_rd[48] , \rt_rd[47] , \rt_rd[46] , 
        \rt_rd[45] , \rt_rd[44] , \rt_rd[43] , \rt_rd[42] , \rt_rd[41] , 
        \rt_rd[40] , \rt_rd[39] , \rt_rd[38] , \rt_rd[37] , \rt_rd[36] , 
        \rt_rd[35] , \rt_rd[34] , \rt_rd[33] , \rt_rd[32] , \rt_rd[31] , 
        \rt_rd[30] , \rt_rd[29] , \rt_rd[28] , \rt_rd[27] , \rt_rd[26] , 
        \rt_rd[25] , \rt_rd[24] , \rt_rd[23] , \rt_rd[22] , \rt_rd[21] , 
        \rt_rd[20] , \rt_rd[19] , \rt_rd[18] , \rt_rd[17] , \rt_rd[16] , 
        \rt_rd[15] , \rt_rd[14] , \rt_rd[13] , \rt_rd[12] , \rt_rd[11] , 
        \rt_rd[10] , \rt_rd[9] , \rt_rd[8] , \rt_rd[7] , \rt_rd[6] , 
        \rt_rd[5] , \rt_rd[4] , \rt_rd[3] , \rt_rd[2] , \rt_rd[1] , \rt_rd[0] 
        }), .route({\route[4] , 1'b0, 1'b0, \route[1] , \route[0] }), 
        .routetxack(routetx_ack) );
    t_adec_dmem dec ( .e_h({SYNOPSYS_UNCONNECTED_1, \eh[1] , \eh[0] }), .e_l({
        \el[2] , \el[1] , \el[0] }), .r_h({\rh[2] , \rh[1] , 
        SYNOPSYS_UNCONNECTED_2}), .r_l({\rl[2] , \rl[1] , \rl[0] }), .e_dp(
        e_dp), .e_ip(e_ip), .e_tic(e_tic), .r_dp(r_dp), .r_ip(r_ip), .r_tic(
        r_tic), .tag_h({\tag_h[4] , \tag_h[3] , \tag_h[2] , \tag_h[1] , 
        \tag_h[0] }), .tag_l({\tag_l[4] , \tag_l[3] , \tag_l[2] , \tag_l[1] , 
        \tag_l[0] }) );
    resp_route_tx_dmem rt ( .o({\route[4] , SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4, \route[1] , \route[0] }), .rtxack(routetx_ack), 
        .e_h({1'b0, \eh[1] , \eh[0] }), .e_l({\el[2] , \el[1] , \el[0] }), 
        .noa(nroute_ack), .r_h({\rh[2] , \rh[1] , 1'b0}), .r_l({\rl[2] , 
        \rl[1] , \rl[0] }), .rtxreq(routetx_req) );
    inv_2 U1 ( .x(reset), .a(nReset) );
    cp2slave_dmem chainif2slave ( .tc_seq({\ct_seq[1] , \ct_seq[0] }), 
        .tc_size({\ct_size[3] , \ct_size[2] , \ct_size[1] , \ct_size[0] }), 
        .tc_itag({\ct_itag[9] , \ct_itag[8] , \ct_itag[7] , \ct_itag[6] , 
        \ct_itag[5] , \ct_itag[4] , \ct_itag[3] , \ct_itag[2] , \ct_itag[1] , 
        \ct_itag[0] }), .tc_wd({\ct_wd[63] , \ct_wd[62] , \ct_wd[61] , 
        \ct_wd[60] , \ct_wd[59] , \ct_wd[58] , \ct_wd[57] , \ct_wd[56] , 
        \ct_wd[55] , \ct_wd[54] , \ct_wd[53] , \ct_wd[52] , \ct_wd[51] , 
        \ct_wd[50] , \ct_wd[49] , \ct_wd[48] , \ct_wd[47] , \ct_wd[46] , 
        \ct_wd[45] , \ct_wd[44] , \ct_wd[43] , \ct_wd[42] , \ct_wd[41] , 
        \ct_wd[40] , \ct_wd[39] , \ct_wd[38] , \ct_wd[37] , \ct_wd[36] , 
        \ct_wd[35] , \ct_wd[34] , \ct_wd[33] , \ct_wd[32] , \ct_wd[31] , 
        \ct_wd[30] , \ct_wd[29] , \ct_wd[28] , \ct_wd[27] , \ct_wd[26] , 
        \ct_wd[25] , \ct_wd[24] , \ct_wd[23] , \ct_wd[22] , \ct_wd[21] , 
        \ct_wd[20] , \ct_wd[19] , \ct_wd[18] , \ct_wd[17] , \ct_wd[16] , 
        \ct_wd[15] , \ct_wd[14] , \ct_wd[13] , \ct_wd[12] , \ct_wd[11] , 
        \ct_wd[10] , \ct_wd[9] , \ct_wd[8] , \ct_wd[7] , \ct_wd[6] , 
        \ct_wd[5] , \ct_wd[4] , \ct_wd[3] , \ct_wd[2] , \ct_wd[1] , \ct_wd[0] 
        }), .tc_lock({\ct_lock[1] , \ct_lock[0] }), .tc_a({\ct_a[63] , 
        \ct_a[62] , \ct_a[61] , \ct_a[60] , \ct_a[59] , \ct_a[58] , \ct_a[57] , 
        \ct_a[56] , \ct_a[55] , \ct_a[54] , \ct_a[53] , \ct_a[52] , \ct_a[51] , 
        \ct_a[50] , \ct_a[49] , \ct_a[48] , \ct_a[47] , \ct_a[46] , \ct_a[45] , 
        \ct_a[44] , \ct_a[43] , \ct_a[42] , \ct_a[41] , \ct_a[40] , \ct_a[39] , 
        \ct_a[38] , \ct_a[37] , \ct_a[36] , \ct_a[35] , \ct_a[34] , \ct_a[33] , 
        \ct_a[32] , \ct_a[31] , \ct_a[30] , \ct_a[29] , \ct_a[28] , \ct_a[27] , 
        \ct_a[26] , \ct_a[25] , \ct_a[24] , \ct_a[23] , \ct_a[22] , \ct_a[21] , 
        \ct_a[20] , \ct_a[19] , \ct_a[18] , \ct_a[17] , \ct_a[16] , \ct_a[15] , 
        \ct_a[14] , \ct_a[13] , \ct_a[12] , \ct_a[11] , \ct_a[10] , \ct_a[9] , 
        \ct_a[8] , \ct_a[7] , \ct_a[6] , \ct_a[5] , \ct_a[4] , \ct_a[3] , 
        \ct_a[2] , \ct_a[1] , \ct_a[0] }), .tc_rnw({\ct_rnw[1] , \ct_rnw[0] }), 
        .tc_ok(ct_ok), .tc_defer(ct_defer), .tc_slow(ct_slow), .tc_ack(ct_ack), 
        .req_in(sc_req), .st_i(sc_st), .we_i(sc_we), .mult_i(sc_mult), .adr_i(
        sc_adr), .dat_i(sc_dat), .seq_i(sc_seq), .sel_i({sc_sel[3], sc_sel[2], 
        sc_sel[1], SYNOPSYS_UNCONNECTED_5}), .ack_in(sc_ack), .tr_rd({
        \rt_rd[63] , \rt_rd[62] , \rt_rd[61] , \rt_rd[60] , \rt_rd[59] , 
        \rt_rd[58] , \rt_rd[57] , \rt_rd[56] , \rt_rd[55] , \rt_rd[54] , 
        \rt_rd[53] , \rt_rd[52] , \rt_rd[51] , \rt_rd[50] , \rt_rd[49] , 
        \rt_rd[48] , \rt_rd[47] , \rt_rd[46] , \rt_rd[45] , \rt_rd[44] , 
        \rt_rd[43] , \rt_rd[42] , \rt_rd[41] , \rt_rd[40] , \rt_rd[39] , 
        \rt_rd[38] , \rt_rd[37] , \rt_rd[36] , \rt_rd[35] , \rt_rd[34] , 
        \rt_rd[33] , \rt_rd[32] , \rt_rd[31] , \rt_rd[30] , \rt_rd[29] , 
        \rt_rd[28] , \rt_rd[27] , \rt_rd[26] , \rt_rd[25] , \rt_rd[24] , 
        \rt_rd[23] , \rt_rd[22] , \rt_rd[21] , \rt_rd[20] , \rt_rd[19] , 
        \rt_rd[18] , \rt_rd[17] , \rt_rd[16] , \rt_rd[15] , \rt_rd[14] , 
        \rt_rd[13] , \rt_rd[12] , \rt_rd[11] , \rt_rd[10] , \rt_rd[9] , 
        \rt_rd[8] , \rt_rd[7] , \rt_rd[6] , \rt_rd[5] , \rt_rd[4] , \rt_rd[3] , 
        \rt_rd[2] , \rt_rd[1] , \rt_rd[0] }), .tr_err({\rt_err[1] , 
        \rt_err[0] }), .tr_ack(rt_ack), .req_out(sr_req), .dat_o(sr_dat), 
        .err_o(sr_err), .rty_o(sr_rty), .acc_o(sr_acc), .sel_o(sr_sel), 
        .mult_o(sr_mult), .rt_o(sr_rt), .ack_out(sr_ack), .reset(reset) );
endmodule


module chain_sendmux8_10 ( ctrlack, oh, ol, i_h, i_l, ctrlreq, oa );
output [7:0] oh;
output [7:0] ol;
input  [7:0] i_h;
input  [7:0] i_l;
input  ctrlreq, oa;
output ctrlack;
    wire \drive[1] , \drive[0] , \U1693/drivemonitor , \U1693/naa , 
        \U1693/net2 , \U1693/net3 , \U1693/bdone , \U1693/U1702/Z ;
    and2_1 \U33_0_/U8  ( .x(oh[0]), .a(i_h[0]), .b(\drive[1] ) );
    and2_1 \U33_1_/U8  ( .x(oh[1]), .a(i_h[1]), .b(\drive[1] ) );
    and2_1 \U33_2_/U8  ( .x(oh[2]), .a(i_h[2]), .b(\drive[1] ) );
    and2_1 \U33_3_/U8  ( .x(oh[3]), .a(i_h[3]), .b(\drive[1] ) );
    and2_1 \U33_4_/U8  ( .x(oh[4]), .a(i_h[4]), .b(\drive[1] ) );
    and2_1 \U33_5_/U8  ( .x(oh[5]), .a(i_h[5]), .b(\drive[1] ) );
    and2_1 \U33_6_/U8  ( .x(oh[6]), .a(i_h[6]), .b(\drive[1] ) );
    and2_1 \U33_7_/U8  ( .x(oh[7]), .a(i_h[7]), .b(\drive[1] ) );
    and2_1 \U1670_0_/U8  ( .x(ol[0]), .a(\drive[0] ), .b(i_l[0]) );
    and2_1 \U1670_1_/U8  ( .x(ol[1]), .a(\drive[0] ), .b(i_l[1]) );
    and2_1 \U1670_2_/U8  ( .x(ol[2]), .a(\drive[0] ), .b(i_l[2]) );
    and2_1 \U1670_3_/U8  ( .x(ol[3]), .a(\drive[0] ), .b(i_l[3]) );
    and2_1 \U1670_4_/U8  ( .x(ol[4]), .a(\drive[0] ), .b(i_l[4]) );
    and2_1 \U1670_5_/U8  ( .x(ol[5]), .a(\drive[0] ), .b(i_l[5]) );
    and2_1 \U1670_6_/U8  ( .x(ol[6]), .a(\drive[0] ), .b(i_l[6]) );
    and2_1 \U1670_7_/U8  ( .x(ol[7]), .a(\drive[0] ), .b(i_l[7]) );
    nor2_2 \U1693/U1703/U6  ( .x(ctrlack), .a(\U1693/drivemonitor ), .b(
        \U1693/naa ) );
    inv_2 \U1693/U1699/U3  ( .x(\U1693/net2 ), .a(\U1693/net3 ) );
    and2_4 \U1693/U2_0_/U8  ( .x(\drive[0] ), .a(ctrlreq), .b(\U1693/net2 ) );
    and2_4 \U1693/U2_1_/U8  ( .x(\drive[1] ), .a(ctrlreq), .b(\U1693/net2 ) );
    inv_1 \U1693/U1701/U3  ( .x(\U1693/naa ), .a(\U1693/bdone ) );
    ao222_1 \U1693/U13/U18/U1/U1  ( .x(\U1693/drivemonitor ), .a(\drive[1] ), 
        .b(\drive[0] ), .c(\drive[1] ), .d(\U1693/drivemonitor ), .e(
        \drive[0] ), .f(\U1693/drivemonitor ) );
    aoi21_1 \U1693/U1702/U30/U1/U1  ( .x(\U1693/bdone ), .a(\U1693/U1702/Z ), 
        .b(oa), .c(\U1693/net2 ) );
    inv_1 \U1693/U1702/U30/U1/U2  ( .x(\U1693/U1702/Z ), .a(\U1693/bdone ) );
    ao23_1 \U1693/U1693/U21/U1/U1  ( .x(\U1693/net3 ), .a(ctrlreq), .b(
        \U1693/net3 ), .c(ctrlreq), .d(\U1693/drivemonitor ), .e(oa) );
endmodule


module chain_sendmux8_9 ( ctrlack, oh, ol, i_h, i_l, ctrlreq, oa );
output [7:0] oh;
output [7:0] ol;
input  [7:0] i_h;
input  [7:0] i_l;
input  ctrlreq, oa;
output ctrlack;
    wire \drive[1] , \drive[0] , \U1693/drivemonitor , \U1693/naa , 
        \U1693/net2 , \U1693/net3 , \U1693/bdone , \U1693/U1702/Z ;
    and2_1 \U33_0_/U8  ( .x(oh[0]), .a(i_h[0]), .b(\drive[1] ) );
    and2_1 \U33_1_/U8  ( .x(oh[1]), .a(i_h[1]), .b(\drive[1] ) );
    and2_1 \U33_2_/U8  ( .x(oh[2]), .a(i_h[2]), .b(\drive[1] ) );
    and2_1 \U33_3_/U8  ( .x(oh[3]), .a(i_h[3]), .b(\drive[1] ) );
    and2_1 \U33_4_/U8  ( .x(oh[4]), .a(i_h[4]), .b(\drive[1] ) );
    and2_1 \U33_5_/U8  ( .x(oh[5]), .a(i_h[5]), .b(\drive[1] ) );
    and2_1 \U33_6_/U8  ( .x(oh[6]), .a(i_h[6]), .b(\drive[1] ) );
    and2_1 \U33_7_/U8  ( .x(oh[7]), .a(i_h[7]), .b(\drive[1] ) );
    and2_1 \U1670_0_/U8  ( .x(ol[0]), .a(\drive[0] ), .b(i_l[0]) );
    and2_1 \U1670_1_/U8  ( .x(ol[1]), .a(\drive[0] ), .b(i_l[1]) );
    and2_1 \U1670_2_/U8  ( .x(ol[2]), .a(\drive[0] ), .b(i_l[2]) );
    and2_1 \U1670_3_/U8  ( .x(ol[3]), .a(\drive[0] ), .b(i_l[3]) );
    and2_1 \U1670_4_/U8  ( .x(ol[4]), .a(\drive[0] ), .b(i_l[4]) );
    and2_1 \U1670_5_/U8  ( .x(ol[5]), .a(\drive[0] ), .b(i_l[5]) );
    and2_1 \U1670_6_/U8  ( .x(ol[6]), .a(\drive[0] ), .b(i_l[6]) );
    and2_1 \U1670_7_/U8  ( .x(ol[7]), .a(\drive[0] ), .b(i_l[7]) );
    nor2_2 \U1693/U1703/U6  ( .x(ctrlack), .a(\U1693/drivemonitor ), .b(
        \U1693/naa ) );
    inv_2 \U1693/U1699/U3  ( .x(\U1693/net2 ), .a(\U1693/net3 ) );
    and2_4 \U1693/U2_0_/U8  ( .x(\drive[0] ), .a(ctrlreq), .b(\U1693/net2 ) );
    and2_4 \U1693/U2_1_/U8  ( .x(\drive[1] ), .a(ctrlreq), .b(\U1693/net2 ) );
    inv_1 \U1693/U1701/U3  ( .x(\U1693/naa ), .a(\U1693/bdone ) );
    ao222_1 \U1693/U13/U18/U1/U1  ( .x(\U1693/drivemonitor ), .a(\drive[1] ), 
        .b(\drive[0] ), .c(\drive[1] ), .d(\U1693/drivemonitor ), .e(
        \drive[0] ), .f(\U1693/drivemonitor ) );
    aoi21_1 \U1693/U1702/U30/U1/U1  ( .x(\U1693/bdone ), .a(\U1693/U1702/Z ), 
        .b(oa), .c(\U1693/net2 ) );
    inv_1 \U1693/U1702/U30/U1/U2  ( .x(\U1693/U1702/Z ), .a(\U1693/bdone ) );
    ao23_1 \U1693/U1693/U21/U1/U1  ( .x(\U1693/net3 ), .a(ctrlreq), .b(
        \U1693/net3 ), .c(ctrlreq), .d(\U1693/drivemonitor ), .e(oa) );
endmodule


module chain_sendmux8_8 ( ctrlack, oh, ol, i_h, i_l, ctrlreq, oa );
output [7:0] oh;
output [7:0] ol;
input  [7:0] i_h;
input  [7:0] i_l;
input  ctrlreq, oa;
output ctrlack;
    wire \drive[1] , \drive[0] , \U1693/drivemonitor , \U1693/naa , 
        \U1693/net2 , \U1693/net3 , \U1693/bdone , \U1693/U1702/Z ;
    and2_1 \U33_0_/U8  ( .x(oh[0]), .a(i_h[0]), .b(\drive[1] ) );
    and2_1 \U33_1_/U8  ( .x(oh[1]), .a(i_h[1]), .b(\drive[1] ) );
    and2_1 \U33_2_/U8  ( .x(oh[2]), .a(i_h[2]), .b(\drive[1] ) );
    and2_1 \U33_3_/U8  ( .x(oh[3]), .a(i_h[3]), .b(\drive[1] ) );
    and2_1 \U33_4_/U8  ( .x(oh[4]), .a(i_h[4]), .b(\drive[1] ) );
    and2_1 \U33_5_/U8  ( .x(oh[5]), .a(i_h[5]), .b(\drive[1] ) );
    and2_1 \U33_6_/U8  ( .x(oh[6]), .a(i_h[6]), .b(\drive[1] ) );
    and2_1 \U33_7_/U8  ( .x(oh[7]), .a(i_h[7]), .b(\drive[1] ) );
    and2_1 \U1670_0_/U8  ( .x(ol[0]), .a(\drive[0] ), .b(i_l[0]) );
    and2_1 \U1670_1_/U8  ( .x(ol[1]), .a(\drive[0] ), .b(i_l[1]) );
    and2_1 \U1670_2_/U8  ( .x(ol[2]), .a(\drive[0] ), .b(i_l[2]) );
    and2_1 \U1670_3_/U8  ( .x(ol[3]), .a(\drive[0] ), .b(i_l[3]) );
    and2_1 \U1670_4_/U8  ( .x(ol[4]), .a(\drive[0] ), .b(i_l[4]) );
    and2_1 \U1670_5_/U8  ( .x(ol[5]), .a(\drive[0] ), .b(i_l[5]) );
    and2_1 \U1670_6_/U8  ( .x(ol[6]), .a(\drive[0] ), .b(i_l[6]) );
    and2_1 \U1670_7_/U8  ( .x(ol[7]), .a(\drive[0] ), .b(i_l[7]) );
    nor2_2 \U1693/U1703/U6  ( .x(ctrlack), .a(\U1693/drivemonitor ), .b(
        \U1693/naa ) );
    inv_2 \U1693/U1699/U3  ( .x(\U1693/net2 ), .a(\U1693/net3 ) );
    and2_4 \U1693/U2_0_/U8  ( .x(\drive[0] ), .a(ctrlreq), .b(\U1693/net2 ) );
    and2_4 \U1693/U2_1_/U8  ( .x(\drive[1] ), .a(ctrlreq), .b(\U1693/net2 ) );
    inv_1 \U1693/U1701/U3  ( .x(\U1693/naa ), .a(\U1693/bdone ) );
    ao222_1 \U1693/U13/U18/U1/U1  ( .x(\U1693/drivemonitor ), .a(\drive[1] ), 
        .b(\drive[0] ), .c(\drive[1] ), .d(\U1693/drivemonitor ), .e(
        \drive[0] ), .f(\U1693/drivemonitor ) );
    aoi21_1 \U1693/U1702/U30/U1/U1  ( .x(\U1693/bdone ), .a(\U1693/U1702/Z ), 
        .b(oa), .c(\U1693/net2 ) );
    inv_1 \U1693/U1702/U30/U1/U2  ( .x(\U1693/U1702/Z ), .a(\U1693/bdone ) );
    ao23_1 \U1693/U1693/U21/U1/U1  ( .x(\U1693/net3 ), .a(ctrlreq), .b(
        \U1693/net3 ), .c(ctrlreq), .d(\U1693/drivemonitor ), .e(oa) );
endmodule


module chain_sendmux8_11 ( ctrlack, oh, ol, i_h, i_l, ctrlreq, oa );
output [7:0] oh;
output [7:0] ol;
input  [7:0] i_h;
input  [7:0] i_l;
input  ctrlreq, oa;
output ctrlack;
    wire \drive[1] , \drive[0] , \U1693/drivemonitor , \U1693/naa , 
        \U1693/net2 , \U1693/net3 , \U1693/bdone , \U1693/U1702/Z ;
    and2_1 \U33_0_/U8  ( .x(oh[0]), .a(i_h[0]), .b(\drive[1] ) );
    and2_1 \U33_1_/U8  ( .x(oh[1]), .a(i_h[1]), .b(\drive[1] ) );
    and2_1 \U33_2_/U8  ( .x(oh[2]), .a(i_h[2]), .b(\drive[1] ) );
    and2_1 \U33_3_/U8  ( .x(oh[3]), .a(i_h[3]), .b(\drive[1] ) );
    and2_1 \U33_4_/U8  ( .x(oh[4]), .a(i_h[4]), .b(\drive[1] ) );
    and2_1 \U33_5_/U8  ( .x(oh[5]), .a(i_h[5]), .b(\drive[1] ) );
    and2_1 \U33_6_/U8  ( .x(oh[6]), .a(i_h[6]), .b(\drive[1] ) );
    and2_1 \U33_7_/U8  ( .x(oh[7]), .a(i_h[7]), .b(\drive[1] ) );
    and2_1 \U1670_0_/U8  ( .x(ol[0]), .a(\drive[0] ), .b(i_l[0]) );
    and2_1 \U1670_1_/U8  ( .x(ol[1]), .a(\drive[0] ), .b(i_l[1]) );
    and2_1 \U1670_2_/U8  ( .x(ol[2]), .a(\drive[0] ), .b(i_l[2]) );
    and2_1 \U1670_3_/U8  ( .x(ol[3]), .a(\drive[0] ), .b(i_l[3]) );
    and2_1 \U1670_4_/U8  ( .x(ol[4]), .a(\drive[0] ), .b(i_l[4]) );
    and2_1 \U1670_5_/U8  ( .x(ol[5]), .a(\drive[0] ), .b(i_l[5]) );
    and2_1 \U1670_6_/U8  ( .x(ol[6]), .a(\drive[0] ), .b(i_l[6]) );
    and2_1 \U1670_7_/U8  ( .x(ol[7]), .a(\drive[0] ), .b(i_l[7]) );
    nor2_2 \U1693/U1703/U6  ( .x(ctrlack), .a(\U1693/drivemonitor ), .b(
        \U1693/naa ) );
    inv_2 \U1693/U1699/U3  ( .x(\U1693/net2 ), .a(\U1693/net3 ) );
    and2_4 \U1693/U2_0_/U8  ( .x(\drive[0] ), .a(ctrlreq), .b(\U1693/net2 ) );
    and2_4 \U1693/U2_1_/U8  ( .x(\drive[1] ), .a(ctrlreq), .b(\U1693/net2 ) );
    inv_1 \U1693/U1701/U3  ( .x(\U1693/naa ), .a(\U1693/bdone ) );
    ao222_1 \U1693/U13/U18/U1/U1  ( .x(\U1693/drivemonitor ), .a(\drive[1] ), 
        .b(\drive[0] ), .c(\drive[1] ), .d(\U1693/drivemonitor ), .e(
        \drive[0] ), .f(\U1693/drivemonitor ) );
    aoi21_1 \U1693/U1702/U30/U1/U1  ( .x(\U1693/bdone ), .a(\U1693/U1702/Z ), 
        .b(oa), .c(\U1693/net2 ) );
    inv_1 \U1693/U1702/U30/U1/U2  ( .x(\U1693/U1702/Z ), .a(\U1693/bdone ) );
    ao23_1 \U1693/U1693/U21/U1/U1  ( .x(\U1693/net3 ), .a(ctrlreq), .b(
        \U1693/net3 ), .c(ctrlreq), .d(\U1693/drivemonitor ), .e(oa) );
endmodule


module chain_sendword_1 ( ctrlack, oh, ol, chainackff, ctrlreq, ih, il );
output [7:0] oh;
output [7:0] ol;
input  [31:0] ih;
input  [31:0] il;
input  chainackff, ctrlreq;
output ctrlack;
    wire net44, \fourth_ol[7] , \fourth_ol[6] , \fourth_ol[5] , \fourth_ol[4] , 
        \fourth_ol[3] , \fourth_ol[2] , \fourth_ol[1] , \fourth_ol[0] , 
        \fourth_oh[7] , \fourth_oh[6] , \fourth_oh[5] , \fourth_oh[4] , 
        \fourth_oh[3] , \fourth_oh[2] , \fourth_oh[1] , \fourth_oh[0] , net51, 
        \third_ol[7] , \third_ol[6] , \third_ol[5] , \third_ol[4] , 
        \third_ol[3] , \third_ol[2] , \third_ol[1] , \third_ol[0] , 
        \third_oh[7] , \third_oh[6] , \third_oh[5] , \third_oh[4] , 
        \third_oh[3] , \third_oh[2] , \third_oh[1] , \third_oh[0] , net58, 
        \second_ol[7] , \second_ol[6] , \second_ol[5] , \second_ol[4] , 
        \second_ol[3] , \second_ol[2] , \second_ol[1] , \second_ol[0] , 
        \second_oh[7] , \second_oh[6] , \second_oh[5] , \second_oh[4] , 
        \second_oh[3] , \second_oh[2] , \second_oh[1] , \second_oh[0] , 
        bctrlreq, \first_ol[7] , \first_ol[6] , \first_ol[5] , \first_ol[4] , 
        \first_ol[3] , \first_ol[2] , \first_ol[1] , \first_ol[0] , 
        \first_oh[7] , \first_oh[6] , \first_oh[5] , \first_oh[4] , 
        \first_oh[3] , \first_oh[2] , \first_oh[1] , \first_oh[0] , 
        \U309_0_/n5 , \U309_0_/n1 , \U309_0_/n2 , \U309_0_/n3 , \U309_0_/n4 , 
        \U309_1_/n5 , \U309_1_/n1 , \U309_1_/n2 , \U309_1_/n3 , \U309_1_/n4 , 
        \U309_2_/n5 , \U309_2_/n1 , \U309_2_/n2 , \U309_2_/n3 , \U309_2_/n4 , 
        \U309_3_/n5 , \U309_3_/n1 , \U309_3_/n2 , \U309_3_/n3 , \U309_3_/n4 , 
        \U309_4_/n5 , \U309_4_/n1 , \U309_4_/n2 , \U309_4_/n3 , \U309_4_/n4 , 
        \U309_5_/n5 , \U309_5_/n1 , \U309_5_/n2 , \U309_5_/n3 , \U309_5_/n4 , 
        \U309_6_/n5 , \U309_6_/n1 , \U309_6_/n2 , \U309_6_/n3 , \U309_6_/n4 , 
        \U309_7_/n5 , \U309_7_/n1 , \U309_7_/n2 , \U309_7_/n3 , \U309_7_/n4 , 
        \U310_0_/n5 , \U310_0_/n1 , \U310_0_/n2 , \U310_0_/n3 , \U310_0_/n4 , 
        \U310_1_/n5 , \U310_1_/n1 , \U310_1_/n2 , \U310_1_/n3 , \U310_1_/n4 , 
        \U310_2_/n5 , \U310_2_/n1 , \U310_2_/n2 , \U310_2_/n3 , \U310_2_/n4 , 
        \U310_3_/n5 , \U310_3_/n1 , \U310_3_/n2 , \U310_3_/n3 , \U310_3_/n4 , 
        \U310_4_/n5 , \U310_4_/n1 , \U310_4_/n2 , \U310_4_/n3 , \U310_4_/n4 , 
        \U310_5_/n5 , \U310_5_/n1 , \U310_5_/n2 , \U310_5_/n3 , \U310_5_/n4 , 
        \U310_6_/n5 , \U310_6_/n1 , \U310_6_/n2 , \U310_6_/n3 , \U310_6_/n4 , 
        \U310_7_/n5 , \U310_7_/n1 , \U310_7_/n2 , \U310_7_/n3 , \U310_7_/n4 ;
    chain_sendmux8_10 I4 ( .ctrlack(ctrlack), .oh({\fourth_oh[7] , 
        \fourth_oh[6] , \fourth_oh[5] , \fourth_oh[4] , \fourth_oh[3] , 
        \fourth_oh[2] , \fourth_oh[1] , \fourth_oh[0] }), .ol({\fourth_ol[7] , 
        \fourth_ol[6] , \fourth_ol[5] , \fourth_ol[4] , \fourth_ol[3] , 
        \fourth_ol[2] , \fourth_ol[1] , \fourth_ol[0] }), .i_h(ih[7:0]), .i_l(
        il[7:0]), .ctrlreq(net44), .oa(chainackff) );
    chain_sendmux8_9 I3 ( .ctrlack(net44), .oh({\third_oh[7] , \third_oh[6] , 
        \third_oh[5] , \third_oh[4] , \third_oh[3] , \third_oh[2] , 
        \third_oh[1] , \third_oh[0] }), .ol({\third_ol[7] , \third_ol[6] , 
        \third_ol[5] , \third_ol[4] , \third_ol[3] , \third_ol[2] , 
        \third_ol[1] , \third_ol[0] }), .i_h(ih[15:8]), .i_l(il[15:8]), 
        .ctrlreq(net51), .oa(chainackff) );
    chain_sendmux8_8 I2 ( .ctrlack(net51), .oh({\second_oh[7] , \second_oh[6] , 
        \second_oh[5] , \second_oh[4] , \second_oh[3] , \second_oh[2] , 
        \second_oh[1] , \second_oh[0] }), .ol({\second_ol[7] , \second_ol[6] , 
        \second_ol[5] , \second_ol[4] , \second_ol[3] , \second_ol[2] , 
        \second_ol[1] , \second_ol[0] }), .i_h(ih[23:16]), .i_l(il[23:16]), 
        .ctrlreq(net58), .oa(chainackff) );
    chain_sendmux8_11 U320 ( .ctrlack(net58), .oh({\first_oh[7] , 
        \first_oh[6] , \first_oh[5] , \first_oh[4] , \first_oh[3] , 
        \first_oh[2] , \first_oh[1] , \first_oh[0] }), .ol({\first_ol[7] , 
        \first_ol[6] , \first_ol[5] , \first_ol[4] , \first_ol[3] , 
        \first_ol[2] , \first_ol[1] , \first_ol[0] }), .i_h(ih[31:24]), .i_l(
        il[31:24]), .ctrlreq(bctrlreq), .oa(chainackff) );
    buf_2 \U328/U7  ( .x(bctrlreq), .a(ctrlreq) );
    and4_2 \U309_0_/U24  ( .x(\U309_0_/n5 ), .a(\U309_0_/n1 ), .b(\U309_0_/n2 
        ), .c(\U309_0_/n3 ), .d(\U309_0_/n4 ) );
    inv_1 \U309_0_/U1  ( .x(\U309_0_/n1 ), .a(\fourth_oh[0] ) );
    inv_1 \U309_0_/U2  ( .x(\U309_0_/n2 ), .a(\third_oh[0] ) );
    inv_1 \U309_0_/U3  ( .x(\U309_0_/n3 ), .a(\second_oh[0] ) );
    inv_1 \U309_0_/U4  ( .x(\U309_0_/n4 ), .a(\first_oh[0] ) );
    inv_4 \U309_0_/U5  ( .x(oh[0]), .a(\U309_0_/n5 ) );
    and4_2 \U309_1_/U24  ( .x(\U309_1_/n5 ), .a(\U309_1_/n1 ), .b(\U309_1_/n2 
        ), .c(\U309_1_/n3 ), .d(\U309_1_/n4 ) );
    inv_1 \U309_1_/U1  ( .x(\U309_1_/n1 ), .a(\fourth_oh[1] ) );
    inv_1 \U309_1_/U2  ( .x(\U309_1_/n2 ), .a(\third_oh[1] ) );
    inv_1 \U309_1_/U3  ( .x(\U309_1_/n3 ), .a(\second_oh[1] ) );
    inv_1 \U309_1_/U4  ( .x(\U309_1_/n4 ), .a(\first_oh[1] ) );
    inv_4 \U309_1_/U5  ( .x(oh[1]), .a(\U309_1_/n5 ) );
    and4_2 \U309_2_/U24  ( .x(\U309_2_/n5 ), .a(\U309_2_/n1 ), .b(\U309_2_/n2 
        ), .c(\U309_2_/n3 ), .d(\U309_2_/n4 ) );
    inv_1 \U309_2_/U1  ( .x(\U309_2_/n1 ), .a(\fourth_oh[2] ) );
    inv_1 \U309_2_/U2  ( .x(\U309_2_/n2 ), .a(\third_oh[2] ) );
    inv_1 \U309_2_/U3  ( .x(\U309_2_/n3 ), .a(\second_oh[2] ) );
    inv_1 \U309_2_/U4  ( .x(\U309_2_/n4 ), .a(\first_oh[2] ) );
    inv_4 \U309_2_/U5  ( .x(oh[2]), .a(\U309_2_/n5 ) );
    and4_2 \U309_3_/U24  ( .x(\U309_3_/n5 ), .a(\U309_3_/n1 ), .b(\U309_3_/n2 
        ), .c(\U309_3_/n3 ), .d(\U309_3_/n4 ) );
    inv_1 \U309_3_/U1  ( .x(\U309_3_/n1 ), .a(\fourth_oh[3] ) );
    inv_1 \U309_3_/U2  ( .x(\U309_3_/n2 ), .a(\third_oh[3] ) );
    inv_1 \U309_3_/U3  ( .x(\U309_3_/n3 ), .a(\second_oh[3] ) );
    inv_1 \U309_3_/U4  ( .x(\U309_3_/n4 ), .a(\first_oh[3] ) );
    inv_4 \U309_3_/U5  ( .x(oh[3]), .a(\U309_3_/n5 ) );
    and4_2 \U309_4_/U24  ( .x(\U309_4_/n5 ), .a(\U309_4_/n1 ), .b(\U309_4_/n2 
        ), .c(\U309_4_/n3 ), .d(\U309_4_/n4 ) );
    inv_1 \U309_4_/U1  ( .x(\U309_4_/n1 ), .a(\fourth_oh[4] ) );
    inv_1 \U309_4_/U2  ( .x(\U309_4_/n2 ), .a(\third_oh[4] ) );
    inv_1 \U309_4_/U3  ( .x(\U309_4_/n3 ), .a(\second_oh[4] ) );
    inv_1 \U309_4_/U4  ( .x(\U309_4_/n4 ), .a(\first_oh[4] ) );
    inv_4 \U309_4_/U5  ( .x(oh[4]), .a(\U309_4_/n5 ) );
    and4_2 \U309_5_/U24  ( .x(\U309_5_/n5 ), .a(\U309_5_/n1 ), .b(\U309_5_/n2 
        ), .c(\U309_5_/n3 ), .d(\U309_5_/n4 ) );
    inv_1 \U309_5_/U1  ( .x(\U309_5_/n1 ), .a(\fourth_oh[5] ) );
    inv_1 \U309_5_/U2  ( .x(\U309_5_/n2 ), .a(\third_oh[5] ) );
    inv_1 \U309_5_/U3  ( .x(\U309_5_/n3 ), .a(\second_oh[5] ) );
    inv_1 \U309_5_/U4  ( .x(\U309_5_/n4 ), .a(\first_oh[5] ) );
    inv_4 \U309_5_/U5  ( .x(oh[5]), .a(\U309_5_/n5 ) );
    and4_2 \U309_6_/U24  ( .x(\U309_6_/n5 ), .a(\U309_6_/n1 ), .b(\U309_6_/n2 
        ), .c(\U309_6_/n3 ), .d(\U309_6_/n4 ) );
    inv_1 \U309_6_/U1  ( .x(\U309_6_/n1 ), .a(\fourth_oh[6] ) );
    inv_1 \U309_6_/U2  ( .x(\U309_6_/n2 ), .a(\third_oh[6] ) );
    inv_1 \U309_6_/U3  ( .x(\U309_6_/n3 ), .a(\second_oh[6] ) );
    inv_1 \U309_6_/U4  ( .x(\U309_6_/n4 ), .a(\first_oh[6] ) );
    inv_4 \U309_6_/U5  ( .x(oh[6]), .a(\U309_6_/n5 ) );
    and4_2 \U309_7_/U24  ( .x(\U309_7_/n5 ), .a(\U309_7_/n1 ), .b(\U309_7_/n2 
        ), .c(\U309_7_/n3 ), .d(\U309_7_/n4 ) );
    inv_1 \U309_7_/U1  ( .x(\U309_7_/n1 ), .a(\fourth_oh[7] ) );
    inv_1 \U309_7_/U2  ( .x(\U309_7_/n2 ), .a(\third_oh[7] ) );
    inv_1 \U309_7_/U3  ( .x(\U309_7_/n3 ), .a(\second_oh[7] ) );
    inv_1 \U309_7_/U4  ( .x(\U309_7_/n4 ), .a(\first_oh[7] ) );
    inv_4 \U309_7_/U5  ( .x(oh[7]), .a(\U309_7_/n5 ) );
    and4_2 \U310_0_/U24  ( .x(\U310_0_/n5 ), .a(\U310_0_/n1 ), .b(\U310_0_/n2 
        ), .c(\U310_0_/n3 ), .d(\U310_0_/n4 ) );
    inv_1 \U310_0_/U1  ( .x(\U310_0_/n1 ), .a(\fourth_ol[0] ) );
    inv_1 \U310_0_/U2  ( .x(\U310_0_/n2 ), .a(\third_ol[0] ) );
    inv_1 \U310_0_/U3  ( .x(\U310_0_/n3 ), .a(\second_ol[0] ) );
    inv_1 \U310_0_/U4  ( .x(\U310_0_/n4 ), .a(\first_ol[0] ) );
    inv_4 \U310_0_/U5  ( .x(ol[0]), .a(\U310_0_/n5 ) );
    and4_2 \U310_1_/U24  ( .x(\U310_1_/n5 ), .a(\U310_1_/n1 ), .b(\U310_1_/n2 
        ), .c(\U310_1_/n3 ), .d(\U310_1_/n4 ) );
    inv_1 \U310_1_/U1  ( .x(\U310_1_/n1 ), .a(\fourth_ol[1] ) );
    inv_1 \U310_1_/U2  ( .x(\U310_1_/n2 ), .a(\third_ol[1] ) );
    inv_1 \U310_1_/U3  ( .x(\U310_1_/n3 ), .a(\second_ol[1] ) );
    inv_1 \U310_1_/U4  ( .x(\U310_1_/n4 ), .a(\first_ol[1] ) );
    inv_4 \U310_1_/U5  ( .x(ol[1]), .a(\U310_1_/n5 ) );
    and4_2 \U310_2_/U24  ( .x(\U310_2_/n5 ), .a(\U310_2_/n1 ), .b(\U310_2_/n2 
        ), .c(\U310_2_/n3 ), .d(\U310_2_/n4 ) );
    inv_1 \U310_2_/U1  ( .x(\U310_2_/n1 ), .a(\fourth_ol[2] ) );
    inv_1 \U310_2_/U2  ( .x(\U310_2_/n2 ), .a(\third_ol[2] ) );
    inv_1 \U310_2_/U3  ( .x(\U310_2_/n3 ), .a(\second_ol[2] ) );
    inv_1 \U310_2_/U4  ( .x(\U310_2_/n4 ), .a(\first_ol[2] ) );
    inv_4 \U310_2_/U5  ( .x(ol[2]), .a(\U310_2_/n5 ) );
    and4_2 \U310_3_/U24  ( .x(\U310_3_/n5 ), .a(\U310_3_/n1 ), .b(\U310_3_/n2 
        ), .c(\U310_3_/n3 ), .d(\U310_3_/n4 ) );
    inv_1 \U310_3_/U1  ( .x(\U310_3_/n1 ), .a(\fourth_ol[3] ) );
    inv_1 \U310_3_/U2  ( .x(\U310_3_/n2 ), .a(\third_ol[3] ) );
    inv_1 \U310_3_/U3  ( .x(\U310_3_/n3 ), .a(\second_ol[3] ) );
    inv_1 \U310_3_/U4  ( .x(\U310_3_/n4 ), .a(\first_ol[3] ) );
    inv_4 \U310_3_/U5  ( .x(ol[3]), .a(\U310_3_/n5 ) );
    and4_2 \U310_4_/U24  ( .x(\U310_4_/n5 ), .a(\U310_4_/n1 ), .b(\U310_4_/n2 
        ), .c(\U310_4_/n3 ), .d(\U310_4_/n4 ) );
    inv_1 \U310_4_/U1  ( .x(\U310_4_/n1 ), .a(\fourth_ol[4] ) );
    inv_1 \U310_4_/U2  ( .x(\U310_4_/n2 ), .a(\third_ol[4] ) );
    inv_1 \U310_4_/U3  ( .x(\U310_4_/n3 ), .a(\second_ol[4] ) );
    inv_1 \U310_4_/U4  ( .x(\U310_4_/n4 ), .a(\first_ol[4] ) );
    inv_4 \U310_4_/U5  ( .x(ol[4]), .a(\U310_4_/n5 ) );
    and4_2 \U310_5_/U24  ( .x(\U310_5_/n5 ), .a(\U310_5_/n1 ), .b(\U310_5_/n2 
        ), .c(\U310_5_/n3 ), .d(\U310_5_/n4 ) );
    inv_1 \U310_5_/U1  ( .x(\U310_5_/n1 ), .a(\fourth_ol[5] ) );
    inv_1 \U310_5_/U2  ( .x(\U310_5_/n2 ), .a(\third_ol[5] ) );
    inv_1 \U310_5_/U3  ( .x(\U310_5_/n3 ), .a(\second_ol[5] ) );
    inv_1 \U310_5_/U4  ( .x(\U310_5_/n4 ), .a(\first_ol[5] ) );
    inv_4 \U310_5_/U5  ( .x(ol[5]), .a(\U310_5_/n5 ) );
    and4_2 \U310_6_/U24  ( .x(\U310_6_/n5 ), .a(\U310_6_/n1 ), .b(\U310_6_/n2 
        ), .c(\U310_6_/n3 ), .d(\U310_6_/n4 ) );
    inv_1 \U310_6_/U1  ( .x(\U310_6_/n1 ), .a(\fourth_ol[6] ) );
    inv_1 \U310_6_/U2  ( .x(\U310_6_/n2 ), .a(\third_ol[6] ) );
    inv_1 \U310_6_/U3  ( .x(\U310_6_/n3 ), .a(\second_ol[6] ) );
    inv_1 \U310_6_/U4  ( .x(\U310_6_/n4 ), .a(\first_ol[6] ) );
    inv_4 \U310_6_/U5  ( .x(ol[6]), .a(\U310_6_/n5 ) );
    and4_2 \U310_7_/U24  ( .x(\U310_7_/n5 ), .a(\U310_7_/n1 ), .b(\U310_7_/n2 
        ), .c(\U310_7_/n3 ), .d(\U310_7_/n4 ) );
    inv_1 \U310_7_/U1  ( .x(\U310_7_/n1 ), .a(\fourth_ol[7] ) );
    inv_1 \U310_7_/U2  ( .x(\U310_7_/n2 ), .a(\third_ol[7] ) );
    inv_1 \U310_7_/U3  ( .x(\U310_7_/n3 ), .a(\second_ol[7] ) );
    inv_1 \U310_7_/U4  ( .x(\U310_7_/n4 ), .a(\first_ol[7] ) );
    inv_4 \U310_7_/U5  ( .x(ol[7]), .a(\U310_7_/n5 ) );
endmodule


module chain_dr8bit_completion_40 ( o, i );
input  [15:0] i;
output o;
    wire \nx[0] , \nx[1] , \nx[2] , \nx[3] , \ny[0] , \ny[1] , \ny[2] , 
        \ny[3] , y, x, \U6/Z , \U3/net3 , \U3/U20/Z , \U3/net2 , \U3/U21/Z , 
        \U3/U19/Z , \U5/net3 , \U5/U20/Z , \U5/net2 , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_43 ( o, i );
input  [15:0] i;
output o;
    wire \nx[0] , \nx[1] , \nx[2] , \nx[3] , \ny[0] , \ny[1] , \ny[2] , 
        \ny[3] , y, x, \U6/Z , \U3/net3 , \U3/U20/Z , \U3/net2 , \U3/U21/Z , 
        \U3/U19/Z , \U5/net3 , \U5/U20/Z , \U5/net2 , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_42 ( o, i );
input  [15:0] i;
output o;
    wire \nx[0] , \nx[1] , \nx[2] , \nx[3] , \ny[0] , \ny[1] , \ny[2] , 
        \ny[3] , y, x, \U6/Z , \U3/net3 , \U3/U20/Z , \U3/net2 , \U3/U21/Z , 
        \U3/U19/Z , \U5/net3 , \U5/U20/Z , \U5/net2 , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr8bit_completion_41 ( o, i );
input  [15:0] i;
output o;
    wire \nx[0] , \nx[1] , \nx[2] , \nx[3] , \ny[0] , \ny[1] , \ny[2] , 
        \ny[3] , y, x, \U6/Z , \U3/net3 , \U3/U20/Z , \U3/net2 , \U3/U21/Z , 
        \U3/U19/Z , \U5/net3 , \U5/U20/Z , \U5/net2 , \U5/U21/Z , \U5/U19/Z ;
    nor2_1 \U2_0_/U5  ( .x(\nx[0] ), .a(i[4]), .b(i[12]) );
    nor2_1 \U2_1_/U5  ( .x(\nx[1] ), .a(i[5]), .b(i[13]) );
    nor2_1 \U2_2_/U5  ( .x(\nx[2] ), .a(i[6]), .b(i[14]) );
    nor2_1 \U2_3_/U5  ( .x(\nx[3] ), .a(i[7]), .b(i[15]) );
    nor2_1 \U4_0_/U5  ( .x(\ny[0] ), .a(i[0]), .b(i[8]) );
    nor2_1 \U4_1_/U5  ( .x(\ny[1] ), .a(i[1]), .b(i[9]) );
    nor2_1 \U4_2_/U5  ( .x(\ny[2] ), .a(i[2]), .b(i[10]) );
    nor2_1 \U4_3_/U5  ( .x(\ny[3] ), .a(i[3]), .b(i[11]) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(y), .b(x), .c(y), .d(\U6/Z ), .e(x), .f(
        \U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U3/U20/U30/U1  ( .x(\U3/net3 ), .a(\nx[3] ), .b(\nx[2] ), .c(
        \nx[3] ), .d(\U3/U20/Z ), .e(\nx[2] ), .f(\U3/U20/Z ) );
    inv_1 \U3/U20/U30/Uinv  ( .x(\U3/U20/Z ), .a(\U3/net3 ) );
    aoi222_1 \U3/U21/U30/U1  ( .x(x), .a(\U3/net3 ), .b(\U3/net2 ), .c(
        \U3/net3 ), .d(\U3/U21/Z ), .e(\U3/net2 ), .f(\U3/U21/Z ) );
    inv_1 \U3/U21/U30/Uinv  ( .x(\U3/U21/Z ), .a(x) );
    aoi222_1 \U3/U19/U30/U1  ( .x(\U3/net2 ), .a(\nx[1] ), .b(\nx[0] ), .c(
        \nx[1] ), .d(\U3/U19/Z ), .e(\nx[0] ), .f(\U3/U19/Z ) );
    inv_1 \U3/U19/U30/Uinv  ( .x(\U3/U19/Z ), .a(\U3/net2 ) );
    aoi222_1 \U5/U20/U30/U1  ( .x(\U5/net3 ), .a(\ny[3] ), .b(\ny[2] ), .c(
        \ny[3] ), .d(\U5/U20/Z ), .e(\ny[2] ), .f(\U5/U20/Z ) );
    inv_1 \U5/U20/U30/Uinv  ( .x(\U5/U20/Z ), .a(\U5/net3 ) );
    aoi222_1 \U5/U21/U30/U1  ( .x(y), .a(\U5/net3 ), .b(\U5/net2 ), .c(
        \U5/net3 ), .d(\U5/U21/Z ), .e(\U5/net2 ), .f(\U5/U21/Z ) );
    inv_1 \U5/U21/U30/Uinv  ( .x(\U5/U21/Z ), .a(y) );
    aoi222_1 \U5/U19/U30/U1  ( .x(\U5/net2 ), .a(\ny[1] ), .b(\ny[0] ), .c(
        \ny[1] ), .d(\U5/U19/Z ), .e(\ny[0] ), .f(\U5/U19/Z ) );
    inv_1 \U5/U19/U30/Uinv  ( .x(\U5/U19/Z ), .a(\U5/net2 ) );
endmodule


module chain_dr32bit_completion_9 ( o, i );
input  [63:0] i;
output o;
    wire \cd[3] , \cd[2] , \cd[1] , \cd[0] , ny, \U16/Z , nx, \U6/Z , \U15/Z ;
    chain_dr8bit_completion_40 U11 ( .o(\cd[3] ), .i({i[63], i[62], i[61], 
        i[60], i[59], i[58], i[57], i[56], i[31], i[30], i[29], i[28], i[27], 
        i[26], i[25], i[24]}) );
    chain_dr8bit_completion_43 U14 ( .o(\cd[2] ), .i({i[55], i[54], i[53], 
        i[52], i[51], i[50], i[49], i[48], i[23], i[22], i[21], i[20], i[19], 
        i[18], i[17], i[16]}) );
    chain_dr8bit_completion_42 U13 ( .o(\cd[1] ), .i({i[47], i[46], i[45], 
        i[44], i[43], i[42], i[41], i[40], i[15], i[14], i[13], i[12], i[11], 
        i[10], i[9], i[8]}) );
    chain_dr8bit_completion_41 U12 ( .o(\cd[0] ), .i({i[39], i[38], i[37], 
        i[36], i[35], i[34], i[33], i[32], i[7], i[6], i[5], i[4], i[3], i[2], 
        i[1], i[0]}) );
    aoi222_1 \U16/U30/U1  ( .x(ny), .a(\cd[0] ), .b(\cd[1] ), .c(\cd[0] ), .d(
        \U16/Z ), .e(\cd[1] ), .f(\U16/Z ) );
    inv_1 \U16/U30/Uinv  ( .x(\U16/Z ), .a(ny) );
    aoi222_1 \U6/U30/U1  ( .x(o), .a(ny), .b(nx), .c(ny), .d(\U6/Z ), .e(nx), 
        .f(\U6/Z ) );
    inv_1 \U6/U30/Uinv  ( .x(\U6/Z ), .a(o) );
    aoi222_1 \U15/U30/U1  ( .x(nx), .a(\cd[3] ), .b(\cd[2] ), .c(\cd[3] ), .d(
        \U15/Z ), .e(\cd[2] ), .f(\U15/Z ) );
    inv_1 \U15/U30/Uinv  ( .x(\U15/Z ), .a(nx) );
endmodule


module chain_selement_ga_64 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_trhdr_1 ( chainff_ack, chainh, chainl, eop, hdrack, normal_ack, 
    notify_ack, read_req, routereq, chain_ff_h, chainack, chainff_l, eopack, 
    err, nReset, normal_response, notify_accept, notify_defer, rcol_h, rcol_l, 
    read_ack, rnw_h, rnw_l, routeack, rsize_h, rsize_l, rtag_h, rtag_l );
output [7:0] chainh;
output [7:0] chainl;
input  [7:0] chain_ff_h;
input  [7:0] chainff_l;
input  [1:0] err;
input  [2:0] rcol_h;
input  [2:0] rcol_l;
input  [1:0] rsize_h;
input  [1:0] rsize_l;
input  [4:0] rtag_h;
input  [4:0] rtag_l;
input  chainack, eopack, nReset, normal_response, notify_accept, notify_defer, 
    read_ack, rnw_h, rnw_l, routeack;
output chainff_ack, eop, hdrack, normal_ack, notify_ack, read_req, routereq;
    wire done_eop, done_pl, \net413[15] , \hdr[16] , \hdr[0] , \net413[14] , 
        \hdr[17] , \hdr[1] , \net413[13] , \net413[12] , \net413[11] , 
        \net413[10] , \net413[9] , \net413[8] , \net413[7] , \net413[6] , 
        \net413[5] , \net413[4] , \net413[3] , \net413[2] , \net413[1] , 
        \net413[0] , net364, donotify, dowrite, net383, done_defer, done_write, 
        done_read, \net343[7] , \drive_l[0] , \net343[6] , \net343[5] , 
        \net343[3] , \net343[2] , \net343[1] , \net343[0] , net340, net337, 
        \net334[7] , \drive_l[1] , \net334[6] , \net334[4] , \net334[2] , 
        \net334[1] , \net334[0] , \net284[7] , \drive_h[1] , \net284[6] , 
        \net284[5] , \net284[4] , \net284[3] , \net284[2] , \net284[1] , 
        \net284[0] , \net288[7] , \drive_h[0] , \net288[6] , \net288[5] , 
        \net288[4] , \net288[3] , \net288[2] , \net288[1] , \net288[0] , 
        net332, done_accept, net321, net359, net362, ctrl_cd, \U311/nz[0] , 
        \U311/nz[1] , \U311/x[3] , \U311/U28/Z , \U311/x[0] , \U311/U32/Z , 
        \U311/x[5] , \U311/U20/Z , \U311/x[2] , \U311/U29/Z , \U311/x[7] , 
        \U311/U25/Z , \U311/y[0] , \U311/x[1] , \U311/U33/Z , \U311/y[2] , 
        \U311/x[4] , \U311/U21/Z , \U311/x[6] , \U311/U26/Z , \U311/y[1] , 
        \U311/U34/Z , \U311/U30/Z , \U311/U19/Z , \U311/y[3] , \U311/U27/Z , 
        \U311/U35/Z , \U311/U31/Z , net407, \U151/Z , done_hdr, 
        \U319/U21/U1/loop , \U323/U21/U1/loop , \U320/U21/U1/loop , 
        \U321/U21/U1/loop , \U322/U21/U1/loop , \U210/drivemonitor , 
        \U210/naa , \U210/net2 , \U210/net3 , net0230, \U210/bdone , 
        \U210/U1702/Z , \I0/drivemonitor , \I0/naa , \I0/net2 , \I0/net3 , 
        \I0/bdone , \I0/U1702/Z ;
    chain_selement_ga_64 U215 ( .Aa(done_eop), .Br(eop), .Ar(done_pl), .Ba(
        eopack) );
    nor2_1 \U308_0_/U5  ( .x(\net413[15] ), .a(\hdr[16] ), .b(\hdr[0] ) );
    nor2_1 \U308_1_/U5  ( .x(\net413[14] ), .a(\hdr[17] ), .b(\hdr[1] ) );
    nor2_1 \U308_2_/U5  ( .x(\net413[13] ), .a(1'b0), .b(routereq) );
    nor2_1 \U308_3_/U5  ( .x(\net413[12] ), .a(routereq), .b(1'b0) );
    nor2_1 \U308_4_/U5  ( .x(\net413[11] ), .a(1'b0), .b(routereq) );
    nor2_1 \U308_5_/U5  ( .x(\net413[10] ), .a(rnw_h), .b(rnw_l) );
    nor2_1 \U308_6_/U5  ( .x(\net413[9] ), .a(rsize_h[0]), .b(rsize_l[0]) );
    nor2_1 \U308_7_/U5  ( .x(\net413[8] ), .a(rsize_h[1]), .b(rsize_l[1]) );
    nor2_1 \U308_8_/U5  ( .x(\net413[7] ), .a(rtag_h[0]), .b(rtag_l[0]) );
    nor2_1 \U308_9_/U5  ( .x(\net413[6] ), .a(rtag_h[1]), .b(rtag_l[1]) );
    nor2_1 \U308_10_/U5  ( .x(\net413[5] ), .a(rtag_h[2]), .b(rtag_l[2]) );
    nor2_1 \U308_11_/U5  ( .x(\net413[4] ), .a(rtag_h[3]), .b(rtag_l[3]) );
    nor2_1 \U308_12_/U5  ( .x(\net413[3] ), .a(rtag_h[4]), .b(rtag_l[4]) );
    nor2_1 \U308_13_/U5  ( .x(\net413[2] ), .a(rcol_h[0]), .b(rcol_l[0]) );
    nor2_1 \U308_14_/U5  ( .x(\net413[1] ), .a(rcol_h[1]), .b(rcol_l[1]) );
    nor2_1 \U308_15_/U5  ( .x(\net413[0] ), .a(rcol_h[2]), .b(rcol_l[2]) );
    or3_1 \U257/U12  ( .x(net364), .a(donotify), .b(dowrite), .c(read_ack) );
    or3_1 \U297/U12  ( .x(net383), .a(done_defer), .b(done_write), .c(
        done_read) );
    and2_2 \U237/U8  ( .x(\hdr[1] ), .a(nReset), .b(normal_response) );
    and2_1 \U307_0_/U8  ( .x(\net343[7] ), .a(\drive_l[0] ), .b(\hdr[0] ) );
    and2_1 \U307_1_/U8  ( .x(\net343[6] ), .a(\drive_l[0] ), .b(\hdr[1] ) );
    and2_1 \U307_2_/U8  ( .x(\net343[5] ), .a(\drive_l[0] ), .b(routereq) );
    and2_1 \U307_4_/U8  ( .x(\net343[3] ), .a(\drive_l[0] ), .b(routereq) );
    and2_1 \U307_5_/U8  ( .x(\net343[2] ), .a(\drive_l[0] ), .b(rnw_l) );
    and2_1 \U307_6_/U8  ( .x(\net343[1] ), .a(\drive_l[0] ), .b(rsize_l[0]) );
    and2_1 \U307_7_/U8  ( .x(\net343[0] ), .a(\drive_l[0] ), .b(rsize_l[1]) );
    and2_1 \U235/U8  ( .x(net340), .a(err[1]), .b(nReset) );
    and2_1 \U236/U8  ( .x(net337), .a(nReset), .b(err[0]) );
    and2_1 \U306_0_/U8  ( .x(\net334[7] ), .a(\hdr[16] ), .b(\drive_l[1] ) );
    and2_1 \U306_1_/U8  ( .x(\net334[6] ), .a(\hdr[17] ), .b(\drive_l[1] ) );
    and2_1 \U306_3_/U8  ( .x(\net334[4] ), .a(routereq), .b(\drive_l[1] ) );
    and2_1 \U306_5_/U8  ( .x(\net334[2] ), .a(rnw_h), .b(\drive_l[1] ) );
    and2_1 \U306_6_/U8  ( .x(\net334[1] ), .a(rsize_h[0]), .b(\drive_l[1] ) );
    and2_1 \U306_7_/U8  ( .x(\net334[0] ), .a(rsize_h[1]), .b(\drive_l[1] ) );
    and2_1 \I1_0_/U8  ( .x(\net284[7] ), .a(rtag_h[0]), .b(\drive_h[1] ) );
    and2_1 \I1_1_/U8  ( .x(\net284[6] ), .a(rtag_h[1]), .b(\drive_h[1] ) );
    and2_1 \I1_2_/U8  ( .x(\net284[5] ), .a(rtag_h[2]), .b(\drive_h[1] ) );
    and2_1 \I1_3_/U8  ( .x(\net284[4] ), .a(rtag_h[3]), .b(\drive_h[1] ) );
    and2_1 \I1_4_/U8  ( .x(\net284[3] ), .a(rtag_h[4]), .b(\drive_h[1] ) );
    and2_1 \I1_5_/U8  ( .x(\net284[2] ), .a(rcol_h[0]), .b(\drive_h[1] ) );
    and2_1 \I1_6_/U8  ( .x(\net284[1] ), .a(rcol_h[1]), .b(\drive_h[1] ) );
    and2_1 \I1_7_/U8  ( .x(\net284[0] ), .a(rcol_h[2]), .b(\drive_h[1] ) );
    and2_1 \I2_0_/U8  ( .x(\net288[7] ), .a(\drive_h[0] ), .b(rtag_l[0]) );
    and2_1 \I2_1_/U8  ( .x(\net288[6] ), .a(\drive_h[0] ), .b(rtag_l[1]) );
    and2_1 \I2_2_/U8  ( .x(\net288[5] ), .a(\drive_h[0] ), .b(rtag_l[2]) );
    and2_1 \I2_3_/U8  ( .x(\net288[4] ), .a(\drive_h[0] ), .b(rtag_l[3]) );
    and2_1 \I2_4_/U8  ( .x(\net288[3] ), .a(\drive_h[0] ), .b(rtag_l[4]) );
    and2_1 \I2_5_/U8  ( .x(\net288[2] ), .a(\drive_h[0] ), .b(rcol_l[0]) );
    and2_1 \I2_6_/U8  ( .x(\net288[1] ), .a(\drive_h[0] ), .b(rcol_l[1]) );
    and2_1 \I2_7_/U8  ( .x(\net288[0] ), .a(\drive_h[0] ), .b(rcol_l[2]) );
    inv_1 \U318/U3  ( .x(net332), .a(routereq) );
    or2_4 \U255/U12  ( .x(notify_ack), .a(done_accept), .b(done_defer) );
    or2_4 \U228/U12  ( .x(\hdr[17] ), .a(notify_defer), .b(notify_accept) );
    or2_4 \U204/U12  ( .x(net321), .a(net359), .b(net362) );
    or2_4 \U221/U12  ( .x(\hdr[16] ), .a(net359), .b(notify_defer) );
    or2_4 \U252/U12  ( .x(normal_ack), .a(done_write), .b(done_read) );
    or2_4 \U280/U12  ( .x(\hdr[0] ), .a(net362), .b(notify_accept) );
    or2_4 \U317/U12  ( .x(routereq), .a(\hdr[17] ), .b(net321) );
    or3_4 \U309_0_/U12  ( .x(chainh[0]), .a(\net334[7] ), .b(\net284[7] ), .c(
        chain_ff_h[0]) );
    or3_4 \U309_1_/U12  ( .x(chainh[1]), .a(\net334[6] ), .b(\net284[6] ), .c(
        chain_ff_h[1]) );
    or3_4 \U309_3_/U12  ( .x(chainh[3]), .a(\net334[4] ), .b(\net284[4] ), .c(
        chain_ff_h[3]) );
    or3_4 \U309_5_/U12  ( .x(chainh[5]), .a(\net334[2] ), .b(\net284[2] ), .c(
        chain_ff_h[5]) );
    or3_4 \U309_6_/U12  ( .x(chainh[6]), .a(\net334[1] ), .b(\net284[1] ), .c(
        chain_ff_h[6]) );
    or3_4 \U309_7_/U12  ( .x(chainh[7]), .a(\net334[0] ), .b(\net284[0] ), .c(
        chain_ff_h[7]) );
    or3_4 \U310_0_/U12  ( .x(chainl[0]), .a(\net343[7] ), .b(\net288[7] ), .c(
        chainff_l[0]) );
    or3_4 \U310_1_/U12  ( .x(chainl[1]), .a(\net343[6] ), .b(\net288[6] ), .c(
        chainff_l[1]) );
    or3_4 \U310_2_/U12  ( .x(chainl[2]), .a(\net343[5] ), .b(\net288[5] ), .c(
        chainff_l[2]) );
    or3_4 \U310_4_/U12  ( .x(chainl[4]), .a(\net343[3] ), .b(\net288[3] ), .c(
        chainff_l[4]) );
    or3_4 \U310_5_/U12  ( .x(chainl[5]), .a(\net343[2] ), .b(\net288[2] ), .c(
        chainff_l[5]) );
    or3_4 \U310_6_/U12  ( .x(chainl[6]), .a(\net343[1] ), .b(\net288[1] ), .c(
        chainff_l[6]) );
    or3_4 \U310_7_/U12  ( .x(chainl[7]), .a(\net343[0] ), .b(\net288[0] ), .c(
        chainff_l[7]) );
    ao222_1 \U311/U37/U18/U1/U1  ( .x(ctrl_cd), .a(\U311/nz[0] ), .b(
        \U311/nz[1] ), .c(\U311/nz[0] ), .d(ctrl_cd), .e(\U311/nz[1] ), .f(
        ctrl_cd) );
    aoi222_1 \U311/U28/U30/U1  ( .x(\U311/x[3] ), .a(\net413[8] ), .b(
        \net413[9] ), .c(\net413[8] ), .d(\U311/U28/Z ), .e(\net413[9] ), .f(
        \U311/U28/Z ) );
    inv_1 \U311/U28/U30/Uinv  ( .x(\U311/U28/Z ), .a(\U311/x[3] ) );
    aoi222_1 \U311/U32/U30/U1  ( .x(\U311/x[0] ), .a(\net413[14] ), .b(
        \net413[15] ), .c(\net413[14] ), .d(\U311/U32/Z ), .e(\net413[15] ), 
        .f(\U311/U32/Z ) );
    inv_1 \U311/U32/U30/Uinv  ( .x(\U311/U32/Z ), .a(\U311/x[0] ) );
    aoi222_1 \U311/U20/U30/U1  ( .x(\U311/x[5] ), .a(\net413[4] ), .b(
        \net413[5] ), .c(\net413[4] ), .d(\U311/U20/Z ), .e(\net413[5] ), .f(
        \U311/U20/Z ) );
    inv_1 \U311/U20/U30/Uinv  ( .x(\U311/U20/Z ), .a(\U311/x[5] ) );
    aoi222_1 \U311/U29/U30/U1  ( .x(\U311/x[2] ), .a(\net413[10] ), .b(
        \net413[11] ), .c(\net413[10] ), .d(\U311/U29/Z ), .e(\net413[11] ), 
        .f(\U311/U29/Z ) );
    inv_1 \U311/U29/U30/Uinv  ( .x(\U311/U29/Z ), .a(\U311/x[2] ) );
    aoi222_1 \U311/U25/U30/U1  ( .x(\U311/x[7] ), .a(\net413[0] ), .b(
        \net413[1] ), .c(\net413[0] ), .d(\U311/U25/Z ), .e(\net413[1] ), .f(
        \U311/U25/Z ) );
    inv_1 \U311/U25/U30/Uinv  ( .x(\U311/U25/Z ), .a(\U311/x[7] ) );
    aoi222_1 \U311/U33/U30/U1  ( .x(\U311/y[0] ), .a(\U311/x[1] ), .b(
        \U311/x[0] ), .c(\U311/x[1] ), .d(\U311/U33/Z ), .e(\U311/x[0] ), .f(
        \U311/U33/Z ) );
    inv_1 \U311/U33/U30/Uinv  ( .x(\U311/U33/Z ), .a(\U311/y[0] ) );
    aoi222_1 \U311/U21/U30/U1  ( .x(\U311/y[2] ), .a(\U311/x[5] ), .b(
        \U311/x[4] ), .c(\U311/x[5] ), .d(\U311/U21/Z ), .e(\U311/x[4] ), .f(
        \U311/U21/Z ) );
    inv_1 \U311/U21/U30/Uinv  ( .x(\U311/U21/Z ), .a(\U311/y[2] ) );
    aoi222_1 \U311/U26/U30/U1  ( .x(\U311/x[6] ), .a(\net413[2] ), .b(
        \net413[3] ), .c(\net413[2] ), .d(\U311/U26/Z ), .e(\net413[3] ), .f(
        \U311/U26/Z ) );
    inv_1 \U311/U26/U30/Uinv  ( .x(\U311/U26/Z ), .a(\U311/x[6] ) );
    aoi222_1 \U311/U34/U30/U1  ( .x(\U311/nz[0] ), .a(\U311/y[1] ), .b(
        \U311/y[0] ), .c(\U311/y[1] ), .d(\U311/U34/Z ), .e(\U311/y[0] ), .f(
        \U311/U34/Z ) );
    inv_1 \U311/U34/U30/Uinv  ( .x(\U311/U34/Z ), .a(\U311/nz[0] ) );
    aoi222_1 \U311/U30/U30/U1  ( .x(\U311/y[1] ), .a(\U311/x[3] ), .b(
        \U311/x[2] ), .c(\U311/x[3] ), .d(\U311/U30/Z ), .e(\U311/x[2] ), .f(
        \U311/U30/Z ) );
    inv_1 \U311/U30/U30/Uinv  ( .x(\U311/U30/Z ), .a(\U311/y[1] ) );
    aoi222_1 \U311/U19/U30/U1  ( .x(\U311/x[4] ), .a(\net413[6] ), .b(
        \net413[7] ), .c(\net413[6] ), .d(\U311/U19/Z ), .e(\net413[7] ), .f(
        \U311/U19/Z ) );
    inv_1 \U311/U19/U30/Uinv  ( .x(\U311/U19/Z ), .a(\U311/x[4] ) );
    aoi222_1 \U311/U27/U30/U1  ( .x(\U311/y[3] ), .a(\U311/x[7] ), .b(
        \U311/x[6] ), .c(\U311/x[7] ), .d(\U311/U27/Z ), .e(\U311/x[6] ), .f(
        \U311/U27/Z ) );
    inv_1 \U311/U27/U30/Uinv  ( .x(\U311/U27/Z ), .a(\U311/y[3] ) );
    aoi222_1 \U311/U35/U30/U1  ( .x(\U311/nz[1] ), .a(\U311/y[3] ), .b(
        \U311/y[2] ), .c(\U311/y[3] ), .d(\U311/U35/Z ), .e(\U311/y[2] ), .f(
        \U311/U35/Z ) );
    inv_1 \U311/U35/U30/Uinv  ( .x(\U311/U35/Z ), .a(\U311/nz[1] ) );
    aoi222_1 \U311/U31/U30/U1  ( .x(\U311/x[1] ), .a(\net413[12] ), .b(
        \net413[13] ), .c(\net413[12] ), .d(\U311/U31/Z ), .e(\net413[13] ), 
        .f(\U311/U31/Z ) );
    inv_1 \U311/U31/U30/Uinv  ( .x(\U311/U31/Z ), .a(\U311/x[1] ) );
    aoi21_1 \U151/U30/U1/U1  ( .x(net407), .a(\U151/Z ), .b(chainff_ack), .c(
        net332) );
    inv_1 \U151/U30/U1/U2  ( .x(\U151/Z ), .a(net407) );
    ao222_1 \U324/U18/U1/U1  ( .x(hdrack), .a(ctrl_cd), .b(net383), .c(ctrl_cd
        ), .d(hdrack), .e(net383), .f(hdrack) );
    ao222_1 \U244/U18/U1/U1  ( .x(donotify), .a(done_hdr), .b(\hdr[17] ), .c(
        done_hdr), .d(donotify), .e(\hdr[17] ), .f(donotify) );
    ao222_1 \U260/U18/U1/U1  ( .x(net362), .a(net337), .b(\hdr[1] ), .c(net337
        ), .d(net362), .e(\hdr[1] ), .f(net362) );
    ao222_1 \U296/U18/U1/U1  ( .x(done_accept), .a(done_eop), .b(notify_accept
        ), .c(done_eop), .d(done_accept), .e(notify_accept), .f(done_accept)
         );
    ao222_1 \U261/U18/U1/U1  ( .x(net359), .a(net340), .b(\hdr[1] ), .c(net340
        ), .d(net359), .e(\hdr[1] ), .f(net359) );
    ao222_1 \U316/U18/U1/U1  ( .x(done_pl), .a(net364), .b(routeack), .c(
        net364), .d(done_pl), .e(routeack), .f(done_pl) );
    ao31_1 \U319/U21/U1/aoi  ( .x(\U319/U21/U1/loop ), .a(\hdr[1] ), .b(
        done_hdr), .c(rnw_h), .d(read_req) );
    oa21_1 \U319/U21/U1/outGate  ( .x(read_req), .a(\hdr[1] ), .b(done_hdr), 
        .c(\U319/U21/U1/loop ) );
    ao31_1 \U323/U21/U1/aoi  ( .x(\U323/U21/U1/loop ), .a(done_eop), .b(
        notify_defer), .c(ctrl_cd), .d(done_defer) );
    oa21_1 \U323/U21/U1/outGate  ( .x(done_defer), .a(done_eop), .b(
        notify_defer), .c(\U323/U21/U1/loop ) );
    ao31_1 \U320/U21/U1/aoi  ( .x(\U320/U21/U1/loop ), .a(\hdr[1] ), .b(
        done_hdr), .c(rnw_l), .d(dowrite) );
    oa21_1 \U320/U21/U1/outGate  ( .x(dowrite), .a(\hdr[1] ), .b(done_hdr), 
        .c(\U320/U21/U1/loop ) );
    ao31_1 \U321/U21/U1/aoi  ( .x(\U321/U21/U1/loop ), .a(read_req), .b(
        done_eop), .c(ctrl_cd), .d(done_read) );
    oa21_1 \U321/U21/U1/outGate  ( .x(done_read), .a(read_req), .b(done_eop), 
        .c(\U321/U21/U1/loop ) );
    ao31_1 \U322/U21/U1/aoi  ( .x(\U322/U21/U1/loop ), .a(dowrite), .b(
        done_eop), .c(ctrl_cd), .d(done_write) );
    oa21_1 \U322/U21/U1/outGate  ( .x(done_write), .a(dowrite), .b(done_eop), 
        .c(\U322/U21/U1/loop ) );
    nor2_2 \U210/U1703/U6  ( .x(done_hdr), .a(\U210/drivemonitor ), .b(
        \U210/naa ) );
    inv_2 \U210/U1699/U3  ( .x(\U210/net2 ), .a(\U210/net3 ) );
    and2_4 \U210/U2_0_/U8  ( .x(\drive_l[0] ), .a(net0230), .b(\U210/net2 ) );
    and2_4 \U210/U2_1_/U8  ( .x(\drive_l[1] ), .a(net0230), .b(\U210/net2 ) );
    inv_1 \U210/U1701/U3  ( .x(\U210/naa ), .a(\U210/bdone ) );
    ao222_1 \U210/U13/U18/U1/U1  ( .x(\U210/drivemonitor ), .a(\drive_l[1] ), 
        .b(\drive_l[0] ), .c(\drive_l[1] ), .d(\U210/drivemonitor ), .e(
        \drive_l[0] ), .f(\U210/drivemonitor ) );
    aoi21_1 \U210/U1702/U30/U1/U1  ( .x(\U210/bdone ), .a(\U210/U1702/Z ), .b(
        chainff_ack), .c(\U210/net2 ) );
    inv_1 \U210/U1702/U30/U1/U2  ( .x(\U210/U1702/Z ), .a(\U210/bdone ) );
    ao23_1 \U210/U1693/U21/U1/U1  ( .x(\U210/net3 ), .a(net0230), .b(
        \U210/net3 ), .c(net0230), .d(\U210/drivemonitor ), .e(chainff_ack) );
    nor2_2 \I0/U1703/U6  ( .x(net0230), .a(\I0/drivemonitor ), .b(\I0/naa ) );
    inv_2 \I0/U1699/U3  ( .x(\I0/net2 ), .a(\I0/net3 ) );
    and2_4 \I0/U2_0_/U8  ( .x(\drive_h[0] ), .a(net407), .b(\I0/net2 ) );
    and2_4 \I0/U2_1_/U8  ( .x(\drive_h[1] ), .a(net407), .b(\I0/net2 ) );
    inv_1 \I0/U1701/U3  ( .x(\I0/naa ), .a(\I0/bdone ) );
    ao222_1 \I0/U13/U18/U1/U1  ( .x(\I0/drivemonitor ), .a(\drive_h[1] ), .b(
        \drive_h[0] ), .c(\drive_h[1] ), .d(\I0/drivemonitor ), .e(
        \drive_h[0] ), .f(\I0/drivemonitor ) );
    aoi21_1 \I0/U1702/U30/U1/U1  ( .x(\I0/bdone ), .a(\I0/U1702/Z ), .b(
        chainff_ack), .c(\I0/net2 ) );
    inv_1 \I0/U1702/U30/U1/U2  ( .x(\I0/U1702/Z ), .a(\I0/bdone ) );
    ao23_1 \I0/U1693/U21/U1/U1  ( .x(\I0/net3 ), .a(net407), .b(\I0/net3 ), 
        .c(net407), .d(\I0/drivemonitor ), .e(chainff_ack) );
    buf_3 U1 ( .x(chainff_ack), .a(chainack) );
    or2_1 U2 ( .x(chainh[4]), .a(chain_ff_h[4]), .b(\net284[3] ) );
    or2_1 U3 ( .x(chainh[2]), .a(chain_ff_h[2]), .b(\net284[5] ) );
    or2_1 U4 ( .x(chainl[3]), .a(chainff_l[3]), .b(\net288[4] ) );
endmodule


module chain_dr2fr_byte_4 ( eop_ack, ia, o, eop, ih, il, nReset, noa );
output [4:0] o;
input  [7:0] ih;
input  [7:0] il;
input  eop, nReset, noa;
output eop_ack, ia;
    wire eop_ack_wire, nbReset, eop_pass, nxa, naa, nlowack, \twobitack[0] , 
        \twobitack[1] , nhighack, \twobitack[2] , \twobitack[3] , \U1018/Z , 
        \U1270/net189 , \U1270/net192 , \U1270/net191 , net199, \U1270/net190 , 
        \U1270/U1141/Z , \U1268/net189 , \U1268/net192 , \U1268/net191 , 
        net194, \U1268/net190 , \U1268/U1141/Z , \U1224/nack[0] , \x[3] , 
        \x[2] , \U1224/nack[1] , \x[1] , \U1224/net4 , \x[0] , 
        \U1224/U1125/U28/U1/clr , asel, \U1224/U1125/U28/U1/set , 
        \U1224/U1122/U28/U1/clr , csel, nca, \U1224/U1122/U28/U1/set , 
        \U1224/U916_0_/U25/U1/clr , \a[0] , \c[0] , \U1224/U916_0_/U25/U1/ob , 
        \U1224/U916_1_/U25/U1/clr , \a[1] , \c[1] , \U1224/U916_1_/U25/U1/ob , 
        \U1224/U916_2_/U25/U1/clr , \a[2] , \c[2] , \U1224/U916_2_/U25/U1/ob , 
        \U1224/U916_3_/U25/U1/clr , \a[3] , \c[3] , \U1224/U916_3_/U25/U1/ob , 
        \U1209/nack[0] , \U1209/nack[1] , \U1209/net4 , 
        \U1209/U1125/U28/U1/clr , xsel, \U1209/U1125/U28/U1/set , 
        \U1209/U1122/U28/U1/clr , ysel, nyla, \U1209/U1122/U28/U1/set , 
        \U1209/U916_0_/U25/U1/clr , \yl[0] , \U1209/U916_0_/U25/U1/ob , 
        \U1209/U916_1_/U25/U1/clr , \yl[1] , \U1209/U916_1_/U25/U1/ob , 
        \U1209/U916_2_/U25/U1/clr , \yl[2] , \U1209/U916_2_/U25/U1/ob , 
        \U1209/U916_3_/U25/U1/clr , \yl[3] , \U1209/U916_3_/U25/U1/ob , 
        \U1213/nack[0] , \y[3] , \y[2] , \U1213/nack[1] , \y[1] , \U1213/net4 , 
        \y[0] , \U1213/U1125/U28/U1/clr , bsel, nba, \U1213/U1125/U28/U1/set , 
        \U1213/U1122/U28/U1/clr , dsel, nda, \U1213/U1122/U28/U1/set , 
        \U1213/U916_0_/U25/U1/clr , nya, \b[0] , \d[0] , 
        \U1213/U916_0_/U25/U1/ob , \U1213/U916_1_/U25/U1/clr , \b[1] , \d[1] , 
        \U1213/U916_1_/U25/U1/ob , \U1213/U916_2_/U25/U1/clr , \b[2] , \d[2] , 
        \U1213/U916_2_/U25/U1/ob , \U1213/U916_3_/U25/U1/clr , \b[3] , \d[3] , 
        \U1213/U916_3_/U25/U1/ob , \cdh[0] , \cdh[1] , \cdl[0] , \cdl[1] , 
        \cdh[2] , \cdh[3] , \cdl[2] , \cdl[3] , cg, \U1296/ng , net195, 
        \U1296/U1384/Z , \U1296/U1386/U25/U1/clr , \U1296/U1386/U25/U1/ob , dg, 
        \U1298/ng , net193, \U1298/U1384/Z , \U1298/U1386/U25/U1/clr , 
        \U1298/U1386/U25/U1/ob , bg, \U1306/ng , \U1306/U1384/Z , 
        \U1306/U1386/U25/U1/clr , \U1306/U1386/U25/U1/ob , ag, \U1295/ng , 
        \U1295/U1384/Z , \U1295/U1386/U25/U1/clr , \U1295/U1386/U25/U1/ob , 
        \U1297/s , \U1297/r , \U1297/nback , \U1297/naack , \U1297/reset , 
        \U1297/U1128/U28/U1/clr , \U1297/U1128/U28/U1/set , 
        \U1297/U1127/U28/U1/clr , \U1297/U1127/U28/U1/set , \U1300/s , 
        \U1300/r , \U1300/nback , \U1300/naack , \U1300/reset , 
        \U1300/U1128/U28/U1/clr , \U1300/U1128/U28/U1/set , 
        \U1300/U1127/U28/U1/clr , \U1300/U1127/U28/U1/set , 
        \U1289/U1150/U28/U1/clr , \U1289/bnreset , \U1289/U1150/U28/U1/set , 
        \U1289/U1152/U28/U1/clr , \U1289/U1152/U28/U1/set , 
        \U1289/U1149/U28/U1/clr , \U1289/U1149/U28/U1/set , 
        \U1289/U1151/U28/U1/clr , \U1289/U1151/U28/U1/set , 
        \U1289/U1148/net189 , \U1289/U1148/net192 , \U1289/U1148/net191 , 
        \U1289/U1148/net190 , \U1289/U1148/U1141/Z , \U1271/U1150/U28/U1/clr , 
        \U1271/bnreset , \U1271/U1150/U28/U1/set , \U1271/U1152/U28/U1/clr , 
        \U1271/U1152/U28/U1/set , \U1271/U1149/U28/U1/clr , 
        \U1271/U1149/U28/U1/set , \U1271/U1151/U28/U1/clr , 
        \U1271/U1151/U28/U1/set , \U1271/U1148/net189 , \U1271/U1148/net192 , 
        \U1271/U1148/net191 , \U1271/U1148/net190 , \U1271/U1148/U1141/Z , 
        \U1225/s , \U1225/r , \U1225/nback , \U1225/naack , \U1225/reset , 
        \U1308/nack[1] , \U1308/nack[0] ;
    assign eop_ack = eop_ack_wire;
    assign o[4] = eop_ack_wire;
    buf_2 U1231 ( .x(nbReset), .a(nReset) );
    and3_1 \U1194/U9  ( .x(eop_pass), .a(nxa), .b(naa), .c(eop) );
    ao222_1 \U1301/U18/U1/U1  ( .x(nlowack), .a(\twobitack[0] ), .b(
        \twobitack[1] ), .c(\twobitack[0] ), .d(nlowack), .e(\twobitack[1] ), 
        .f(nlowack) );
    ao222_1 \U1302/U18/U1/U1  ( .x(nhighack), .a(\twobitack[2] ), .b(
        \twobitack[3] ), .c(\twobitack[2] ), .d(nhighack), .e(\twobitack[3] ), 
        .f(nhighack) );
    aoi222_1 \U1018/U30/U1  ( .x(ia), .a(nhighack), .b(nlowack), .c(nhighack), 
        .d(\U1018/Z ), .e(nlowack), .f(\U1018/Z ) );
    inv_1 \U1018/U30/Uinv  ( .x(\U1018/Z ), .a(ia) );
    ao222_2 \U1038/U19/U1/U1  ( .x(eop_ack_wire), .a(eop_pass), .b(noa), .c(
        eop_pass), .d(eop_ack_wire), .e(noa), .f(eop_ack_wire) );
    inv_1 \U1270/U1147/U3  ( .x(\U1270/net189 ), .a(nbReset) );
    nor2_1 \U1270/U582/U5  ( .x(\U1270/net192 ), .a(il[4]), .b(ih[4]) );
    nor2_1 \U1270/U580/U5  ( .x(\U1270/net191 ), .a(il[5]), .b(ih[5]) );
    nor2_2 \U1270/U1146/U6  ( .x(net199), .a(\U1270/net190 ), .b(
        \U1270/net189 ) );
    aoi222_1 \U1270/U1141/U30/U1  ( .x(\U1270/net190 ), .a(\U1270/net191 ), 
        .b(\U1270/net192 ), .c(\U1270/net191 ), .d(\U1270/U1141/Z ), .e(
        \U1270/net192 ), .f(\U1270/U1141/Z ) );
    inv_1 \U1270/U1141/U30/Uinv  ( .x(\U1270/U1141/Z ), .a(\U1270/net190 ) );
    inv_1 \U1268/U1147/U3  ( .x(\U1268/net189 ), .a(nbReset) );
    nor2_1 \U1268/U582/U5  ( .x(\U1268/net192 ), .a(il[6]), .b(ih[6]) );
    nor2_1 \U1268/U580/U5  ( .x(\U1268/net191 ), .a(il[7]), .b(ih[7]) );
    nor2_2 \U1268/U1146/U6  ( .x(net194), .a(\U1268/net190 ), .b(
        \U1268/net189 ) );
    aoi222_1 \U1268/U1141/U30/U1  ( .x(\U1268/net190 ), .a(\U1268/net191 ), 
        .b(\U1268/net192 ), .c(\U1268/net191 ), .d(\U1268/U1141/Z ), .e(
        \U1268/net192 ), .f(\U1268/U1141/Z ) );
    inv_1 \U1268/U1141/U30/Uinv  ( .x(\U1268/U1141/Z ), .a(\U1268/net190 ) );
    nor2_1 \U1224/U1128/U5  ( .x(\U1224/nack[0] ), .a(\x[3] ), .b(\x[2] ) );
    nor3_1 \U1224/U1127/U7  ( .x(\U1224/nack[1] ), .a(\x[1] ), .b(\U1224/net4 
        ), .c(\x[0] ) );
    inv_1 \U1224/U907/U3  ( .x(\U1224/net4 ), .a(nbReset) );
    aoai211_1 \U1224/U1125/U28/U1/U1  ( .x(\U1224/U1125/U28/U1/clr ), .a(
        \U1224/nack[1] ), .b(\U1224/nack[0] ), .c(asel), .d(naa) );
    nand3_1 \U1224/U1125/U28/U1/U2  ( .x(\U1224/U1125/U28/U1/set ), .a(asel), 
        .b(\U1224/nack[1] ), .c(\U1224/nack[0] ) );
    nand2_2 \U1224/U1125/U28/U1/U3  ( .x(naa), .a(\U1224/U1125/U28/U1/clr ), 
        .b(\U1224/U1125/U28/U1/set ) );
    aoai211_1 \U1224/U1122/U28/U1/U1  ( .x(\U1224/U1122/U28/U1/clr ), .a(
        \U1224/nack[0] ), .b(\U1224/nack[1] ), .c(csel), .d(nca) );
    nand3_1 \U1224/U1122/U28/U1/U2  ( .x(\U1224/U1122/U28/U1/set ), .a(csel), 
        .b(\U1224/nack[0] ), .c(\U1224/nack[1] ) );
    nand2_2 \U1224/U1122/U28/U1/U3  ( .x(nca), .a(\U1224/U1122/U28/U1/clr ), 
        .b(\U1224/U1122/U28/U1/set ) );
    oa31_1 \U1224/U916_0_/U25/U1/Uclr  ( .x(\U1224/U916_0_/U25/U1/clr ), .a(
        nxa), .b(\a[0] ), .c(\c[0] ), .d(\x[0] ) );
    oaoi211_1 \U1224/U916_0_/U25/U1/Uaoi  ( .x(\U1224/U916_0_/U25/U1/ob ), .a(
        \a[0] ), .b(\c[0] ), .c(nxa), .d(\U1224/U916_0_/U25/U1/clr ) );
    inv_2 \U1224/U916_0_/U25/U1/Ui  ( .x(\x[0] ), .a(\U1224/U916_0_/U25/U1/ob 
        ) );
    oa31_1 \U1224/U916_1_/U25/U1/Uclr  ( .x(\U1224/U916_1_/U25/U1/clr ), .a(
        nxa), .b(\a[1] ), .c(\c[1] ), .d(\x[1] ) );
    oaoi211_1 \U1224/U916_1_/U25/U1/Uaoi  ( .x(\U1224/U916_1_/U25/U1/ob ), .a(
        \a[1] ), .b(\c[1] ), .c(nxa), .d(\U1224/U916_1_/U25/U1/clr ) );
    inv_2 \U1224/U916_1_/U25/U1/Ui  ( .x(\x[1] ), .a(\U1224/U916_1_/U25/U1/ob 
        ) );
    oa31_1 \U1224/U916_2_/U25/U1/Uclr  ( .x(\U1224/U916_2_/U25/U1/clr ), .a(
        nxa), .b(\a[2] ), .c(\c[2] ), .d(\x[2] ) );
    oaoi211_1 \U1224/U916_2_/U25/U1/Uaoi  ( .x(\U1224/U916_2_/U25/U1/ob ), .a(
        \a[2] ), .b(\c[2] ), .c(nxa), .d(\U1224/U916_2_/U25/U1/clr ) );
    inv_2 \U1224/U916_2_/U25/U1/Ui  ( .x(\x[2] ), .a(\U1224/U916_2_/U25/U1/ob 
        ) );
    oa31_1 \U1224/U916_3_/U25/U1/Uclr  ( .x(\U1224/U916_3_/U25/U1/clr ), .a(
        nxa), .b(\a[3] ), .c(\c[3] ), .d(\x[3] ) );
    oaoi211_1 \U1224/U916_3_/U25/U1/Uaoi  ( .x(\U1224/U916_3_/U25/U1/ob ), .a(
        \a[3] ), .b(\c[3] ), .c(nxa), .d(\U1224/U916_3_/U25/U1/clr ) );
    inv_2 \U1224/U916_3_/U25/U1/Ui  ( .x(\x[3] ), .a(\U1224/U916_3_/U25/U1/ob 
        ) );
    nor2_1 \U1209/U1128/U5  ( .x(\U1209/nack[0] ), .a(o[3]), .b(o[2]) );
    nor3_1 \U1209/U1127/U7  ( .x(\U1209/nack[1] ), .a(o[1]), .b(\U1209/net4 ), 
        .c(o[0]) );
    inv_1 \U1209/U907/U3  ( .x(\U1209/net4 ), .a(nbReset) );
    aoai211_1 \U1209/U1125/U28/U1/U1  ( .x(\U1209/U1125/U28/U1/clr ), .a(
        \U1209/nack[1] ), .b(\U1209/nack[0] ), .c(xsel), .d(nxa) );
    nand3_1 \U1209/U1125/U28/U1/U2  ( .x(\U1209/U1125/U28/U1/set ), .a(xsel), 
        .b(\U1209/nack[1] ), .c(\U1209/nack[0] ) );
    nand2_2 \U1209/U1125/U28/U1/U3  ( .x(nxa), .a(\U1209/U1125/U28/U1/clr ), 
        .b(\U1209/U1125/U28/U1/set ) );
    aoai211_1 \U1209/U1122/U28/U1/U1  ( .x(\U1209/U1122/U28/U1/clr ), .a(
        \U1209/nack[0] ), .b(\U1209/nack[1] ), .c(ysel), .d(nyla) );
    nand3_1 \U1209/U1122/U28/U1/U2  ( .x(\U1209/U1122/U28/U1/set ), .a(ysel), 
        .b(\U1209/nack[0] ), .c(\U1209/nack[1] ) );
    nand2_2 \U1209/U1122/U28/U1/U3  ( .x(nyla), .a(\U1209/U1122/U28/U1/clr ), 
        .b(\U1209/U1122/U28/U1/set ) );
    oa31_1 \U1209/U916_0_/U25/U1/Uclr  ( .x(\U1209/U916_0_/U25/U1/clr ), .a(
        noa), .b(\x[0] ), .c(\yl[0] ), .d(o[0]) );
    oaoi211_1 \U1209/U916_0_/U25/U1/Uaoi  ( .x(\U1209/U916_0_/U25/U1/ob ), .a(
        \x[0] ), .b(\yl[0] ), .c(noa), .d(\U1209/U916_0_/U25/U1/clr ) );
    inv_2 \U1209/U916_0_/U25/U1/Ui  ( .x(o[0]), .a(\U1209/U916_0_/U25/U1/ob )
         );
    oa31_1 \U1209/U916_1_/U25/U1/Uclr  ( .x(\U1209/U916_1_/U25/U1/clr ), .a(
        noa), .b(\x[1] ), .c(\yl[1] ), .d(o[1]) );
    oaoi211_1 \U1209/U916_1_/U25/U1/Uaoi  ( .x(\U1209/U916_1_/U25/U1/ob ), .a(
        \x[1] ), .b(\yl[1] ), .c(noa), .d(\U1209/U916_1_/U25/U1/clr ) );
    inv_2 \U1209/U916_1_/U25/U1/Ui  ( .x(o[1]), .a(\U1209/U916_1_/U25/U1/ob )
         );
    oa31_1 \U1209/U916_2_/U25/U1/Uclr  ( .x(\U1209/U916_2_/U25/U1/clr ), .a(
        noa), .b(\x[2] ), .c(\yl[2] ), .d(o[2]) );
    oaoi211_1 \U1209/U916_2_/U25/U1/Uaoi  ( .x(\U1209/U916_2_/U25/U1/ob ), .a(
        \x[2] ), .b(\yl[2] ), .c(noa), .d(\U1209/U916_2_/U25/U1/clr ) );
    inv_2 \U1209/U916_2_/U25/U1/Ui  ( .x(o[2]), .a(\U1209/U916_2_/U25/U1/ob )
         );
    oa31_1 \U1209/U916_3_/U25/U1/Uclr  ( .x(\U1209/U916_3_/U25/U1/clr ), .a(
        noa), .b(\x[3] ), .c(\yl[3] ), .d(o[3]) );
    oaoi211_1 \U1209/U916_3_/U25/U1/Uaoi  ( .x(\U1209/U916_3_/U25/U1/ob ), .a(
        \x[3] ), .b(\yl[3] ), .c(noa), .d(\U1209/U916_3_/U25/U1/clr ) );
    inv_2 \U1209/U916_3_/U25/U1/Ui  ( .x(o[3]), .a(\U1209/U916_3_/U25/U1/ob )
         );
    nor2_1 \U1213/U1128/U5  ( .x(\U1213/nack[0] ), .a(\y[3] ), .b(\y[2] ) );
    nor3_1 \U1213/U1127/U7  ( .x(\U1213/nack[1] ), .a(\y[1] ), .b(\U1213/net4 
        ), .c(\y[0] ) );
    inv_1 \U1213/U907/U3  ( .x(\U1213/net4 ), .a(nbReset) );
    aoai211_1 \U1213/U1125/U28/U1/U1  ( .x(\U1213/U1125/U28/U1/clr ), .a(
        \U1213/nack[1] ), .b(\U1213/nack[0] ), .c(bsel), .d(nba) );
    nand3_1 \U1213/U1125/U28/U1/U2  ( .x(\U1213/U1125/U28/U1/set ), .a(bsel), 
        .b(\U1213/nack[1] ), .c(\U1213/nack[0] ) );
    nand2_2 \U1213/U1125/U28/U1/U3  ( .x(nba), .a(\U1213/U1125/U28/U1/clr ), 
        .b(\U1213/U1125/U28/U1/set ) );
    aoai211_1 \U1213/U1122/U28/U1/U1  ( .x(\U1213/U1122/U28/U1/clr ), .a(
        \U1213/nack[0] ), .b(\U1213/nack[1] ), .c(dsel), .d(nda) );
    nand3_1 \U1213/U1122/U28/U1/U2  ( .x(\U1213/U1122/U28/U1/set ), .a(dsel), 
        .b(\U1213/nack[0] ), .c(\U1213/nack[1] ) );
    nand2_2 \U1213/U1122/U28/U1/U3  ( .x(nda), .a(\U1213/U1122/U28/U1/clr ), 
        .b(\U1213/U1122/U28/U1/set ) );
    oa31_1 \U1213/U916_0_/U25/U1/Uclr  ( .x(\U1213/U916_0_/U25/U1/clr ), .a(
        nya), .b(\b[0] ), .c(\d[0] ), .d(\y[0] ) );
    oaoi211_1 \U1213/U916_0_/U25/U1/Uaoi  ( .x(\U1213/U916_0_/U25/U1/ob ), .a(
        \b[0] ), .b(\d[0] ), .c(nya), .d(\U1213/U916_0_/U25/U1/clr ) );
    inv_2 \U1213/U916_0_/U25/U1/Ui  ( .x(\y[0] ), .a(\U1213/U916_0_/U25/U1/ob 
        ) );
    oa31_1 \U1213/U916_1_/U25/U1/Uclr  ( .x(\U1213/U916_1_/U25/U1/clr ), .a(
        nya), .b(\b[1] ), .c(\d[1] ), .d(\y[1] ) );
    oaoi211_1 \U1213/U916_1_/U25/U1/Uaoi  ( .x(\U1213/U916_1_/U25/U1/ob ), .a(
        \b[1] ), .b(\d[1] ), .c(nya), .d(\U1213/U916_1_/U25/U1/clr ) );
    inv_2 \U1213/U916_1_/U25/U1/Ui  ( .x(\y[1] ), .a(\U1213/U916_1_/U25/U1/ob 
        ) );
    oa31_1 \U1213/U916_2_/U25/U1/Uclr  ( .x(\U1213/U916_2_/U25/U1/clr ), .a(
        nya), .b(\b[2] ), .c(\d[2] ), .d(\y[2] ) );
    oaoi211_1 \U1213/U916_2_/U25/U1/Uaoi  ( .x(\U1213/U916_2_/U25/U1/ob ), .a(
        \b[2] ), .b(\d[2] ), .c(nya), .d(\U1213/U916_2_/U25/U1/clr ) );
    inv_2 \U1213/U916_2_/U25/U1/Ui  ( .x(\y[2] ), .a(\U1213/U916_2_/U25/U1/ob 
        ) );
    oa31_1 \U1213/U916_3_/U25/U1/Uclr  ( .x(\U1213/U916_3_/U25/U1/clr ), .a(
        nya), .b(\b[3] ), .c(\d[3] ), .d(\y[3] ) );
    oaoi211_1 \U1213/U916_3_/U25/U1/Uaoi  ( .x(\U1213/U916_3_/U25/U1/ob ), .a(
        \b[3] ), .b(\d[3] ), .c(nya), .d(\U1213/U916_3_/U25/U1/clr ) );
    inv_2 \U1213/U916_3_/U25/U1/Ui  ( .x(\y[3] ), .a(\U1213/U916_3_/U25/U1/ob 
        ) );
    and3_2 \U1210/U1138/U9  ( .x(\d[3] ), .a(\cdh[0] ), .b(nda), .c(\cdh[1] )
         );
    and3_2 \U1210/U1137/U9  ( .x(\d[2] ), .a(\cdl[0] ), .b(nda), .c(\cdh[1] )
         );
    and3_2 \U1210/U1139/U9  ( .x(\d[1] ), .a(\cdh[0] ), .b(nda), .c(\cdl[1] )
         );
    and3_2 \U1210/U1136/U9  ( .x(\d[0] ), .a(\cdl[0] ), .b(nda), .c(\cdl[1] )
         );
    and3_2 \U1162/U1138/U9  ( .x(\a[3] ), .a(ih[6]), .b(naa), .c(ih[7]) );
    and3_2 \U1162/U1137/U9  ( .x(\a[2] ), .a(il[6]), .b(naa), .c(ih[7]) );
    and3_2 \U1162/U1139/U9  ( .x(\a[1] ), .a(ih[6]), .b(naa), .c(il[7]) );
    and3_2 \U1162/U1136/U9  ( .x(\a[0] ), .a(il[6]), .b(naa), .c(il[7]) );
    and3_2 \U1211/U1138/U9  ( .x(\b[3] ), .a(ih[4]), .b(nba), .c(ih[5]) );
    and3_2 \U1211/U1137/U9  ( .x(\b[2] ), .a(il[4]), .b(nba), .c(ih[5]) );
    and3_2 \U1211/U1139/U9  ( .x(\b[1] ), .a(ih[4]), .b(nba), .c(il[5]) );
    and3_2 \U1211/U1136/U9  ( .x(\b[0] ), .a(il[4]), .b(nba), .c(il[5]) );
    and3_2 \U1163/U1138/U9  ( .x(\c[3] ), .a(\cdh[2] ), .b(nca), .c(\cdh[3] )
         );
    and3_2 \U1163/U1137/U9  ( .x(\c[2] ), .a(\cdl[2] ), .b(nca), .c(\cdh[3] )
         );
    and3_2 \U1163/U1139/U9  ( .x(\c[1] ), .a(\cdh[2] ), .b(nca), .c(\cdl[3] )
         );
    and3_2 \U1163/U1136/U9  ( .x(\c[0] ), .a(\cdl[2] ), .b(nca), .c(\cdl[3] )
         );
    and2_1 \U1296/U1385/U8  ( .x(cg), .a(nbReset), .b(\U1296/ng ) );
    aoi222_1 \U1296/U1384/U30/U1  ( .x(\U1296/ng ), .a(nca), .b(net195), .c(
        nca), .d(\U1296/U1384/Z ), .e(net195), .f(\U1296/U1384/Z ) );
    inv_1 \U1296/U1384/U30/Uinv  ( .x(\U1296/U1384/Z ), .a(\U1296/ng ) );
    oa31_1 \U1296/U1386/U25/U1/Uclr  ( .x(\U1296/U1386/U25/U1/clr ), .a(
        \twobitack[2] ), .b(cg), .c(nca), .d(net195) );
    oaoi211_1 \U1296/U1386/U25/U1/Uaoi  ( .x(\U1296/U1386/U25/U1/ob ), .a(cg), 
        .b(nca), .c(\twobitack[2] ), .d(\U1296/U1386/U25/U1/clr ) );
    inv_2 \U1296/U1386/U25/U1/Ui  ( .x(net195), .a(\U1296/U1386/U25/U1/ob ) );
    and2_1 \U1298/U1385/U8  ( .x(dg), .a(nbReset), .b(\U1298/ng ) );
    aoi222_1 \U1298/U1384/U30/U1  ( .x(\U1298/ng ), .a(nda), .b(net193), .c(
        nda), .d(\U1298/U1384/Z ), .e(net193), .f(\U1298/U1384/Z ) );
    inv_1 \U1298/U1384/U30/Uinv  ( .x(\U1298/U1384/Z ), .a(\U1298/ng ) );
    oa31_1 \U1298/U1386/U25/U1/Uclr  ( .x(\U1298/U1386/U25/U1/clr ), .a(
        \twobitack[0] ), .b(dg), .c(nda), .d(net193) );
    oaoi211_1 \U1298/U1386/U25/U1/Uaoi  ( .x(\U1298/U1386/U25/U1/ob ), .a(dg), 
        .b(nda), .c(\twobitack[0] ), .d(\U1298/U1386/U25/U1/clr ) );
    inv_2 \U1298/U1386/U25/U1/Ui  ( .x(net193), .a(\U1298/U1386/U25/U1/ob ) );
    and2_1 \U1306/U1385/U8  ( .x(bg), .a(nbReset), .b(\U1306/ng ) );
    aoi222_1 \U1306/U1384/U30/U1  ( .x(\U1306/ng ), .a(nba), .b(\twobitack[1] 
        ), .c(nba), .d(\U1306/U1384/Z ), .e(\twobitack[1] ), .f(
        \U1306/U1384/Z ) );
    inv_1 \U1306/U1384/U30/Uinv  ( .x(\U1306/U1384/Z ), .a(\U1306/ng ) );
    oa31_1 \U1306/U1386/U25/U1/Uclr  ( .x(\U1306/U1386/U25/U1/clr ), .a(net199
        ), .b(bg), .c(nba), .d(\twobitack[1] ) );
    oaoi211_1 \U1306/U1386/U25/U1/Uaoi  ( .x(\U1306/U1386/U25/U1/ob ), .a(bg), 
        .b(nba), .c(net199), .d(\U1306/U1386/U25/U1/clr ) );
    inv_2 \U1306/U1386/U25/U1/Ui  ( .x(\twobitack[1] ), .a(
        \U1306/U1386/U25/U1/ob ) );
    and2_1 \U1295/U1385/U8  ( .x(ag), .a(nbReset), .b(\U1295/ng ) );
    aoi222_1 \U1295/U1384/U30/U1  ( .x(\U1295/ng ), .a(naa), .b(\twobitack[3] 
        ), .c(naa), .d(\U1295/U1384/Z ), .e(\twobitack[3] ), .f(
        \U1295/U1384/Z ) );
    inv_1 \U1295/U1384/U30/Uinv  ( .x(\U1295/U1384/Z ), .a(\U1295/ng ) );
    oa31_1 \U1295/U1386/U25/U1/Uclr  ( .x(\U1295/U1386/U25/U1/clr ), .a(net194
        ), .b(ag), .c(naa), .d(\twobitack[3] ) );
    oaoi211_1 \U1295/U1386/U25/U1/Uaoi  ( .x(\U1295/U1386/U25/U1/ob ), .a(ag), 
        .b(naa), .c(net194), .d(\U1295/U1386/U25/U1/clr ) );
    inv_2 \U1295/U1386/U25/U1/Ui  ( .x(\twobitack[3] ), .a(
        \U1295/U1386/U25/U1/ob ) );
    nand2_1 \U1297/U1131/U5  ( .x(\U1297/s ), .a(\U1297/r ), .b(\U1297/nback )
         );
    nand2_1 \U1297/U1103/U5  ( .x(\U1297/r ), .a(\U1297/naack ), .b(\U1297/s )
         );
    inv_1 \U1297/U1111/U3  ( .x(\U1297/reset ), .a(nbReset) );
    inv_1 \U1297/U1112/U3  ( .x(\U1297/naack ), .a(naa) );
    nor2_1 \U1297/U1130/U5  ( .x(\U1297/nback ), .a(nca), .b(\U1297/reset ) );
    aoai211_1 \U1297/U1128/U28/U1/U1  ( .x(\U1297/U1128/U28/U1/clr ), .a(
        \U1297/r ), .b(\U1297/naack ), .c(cg), .d(csel) );
    nand3_1 \U1297/U1128/U28/U1/U2  ( .x(\U1297/U1128/U28/U1/set ), .a(cg), 
        .b(\U1297/r ), .c(\U1297/naack ) );
    nand2_2 \U1297/U1128/U28/U1/U3  ( .x(csel), .a(\U1297/U1128/U28/U1/clr ), 
        .b(\U1297/U1128/U28/U1/set ) );
    aoai211_1 \U1297/U1127/U28/U1/U1  ( .x(\U1297/U1127/U28/U1/clr ), .a(
        \U1297/s ), .b(\U1297/nback ), .c(ag), .d(asel) );
    nand3_1 \U1297/U1127/U28/U1/U2  ( .x(\U1297/U1127/U28/U1/set ), .a(ag), 
        .b(\U1297/s ), .c(\U1297/nback ) );
    nand2_2 \U1297/U1127/U28/U1/U3  ( .x(asel), .a(\U1297/U1127/U28/U1/clr ), 
        .b(\U1297/U1127/U28/U1/set ) );
    nand2_1 \U1300/U1131/U5  ( .x(\U1300/s ), .a(\U1300/r ), .b(\U1300/nback )
         );
    nand2_1 \U1300/U1103/U5  ( .x(\U1300/r ), .a(\U1300/naack ), .b(\U1300/s )
         );
    inv_1 \U1300/U1111/U3  ( .x(\U1300/reset ), .a(nbReset) );
    inv_1 \U1300/U1112/U3  ( .x(\U1300/naack ), .a(nba) );
    nor2_1 \U1300/U1130/U5  ( .x(\U1300/nback ), .a(nda), .b(\U1300/reset ) );
    aoai211_1 \U1300/U1128/U28/U1/U1  ( .x(\U1300/U1128/U28/U1/clr ), .a(
        \U1300/r ), .b(\U1300/naack ), .c(dg), .d(dsel) );
    nand3_1 \U1300/U1128/U28/U1/U2  ( .x(\U1300/U1128/U28/U1/set ), .a(dg), 
        .b(\U1300/r ), .c(\U1300/naack ) );
    nand2_2 \U1300/U1128/U28/U1/U3  ( .x(dsel), .a(\U1300/U1128/U28/U1/clr ), 
        .b(\U1300/U1128/U28/U1/set ) );
    aoai211_1 \U1300/U1127/U28/U1/U1  ( .x(\U1300/U1127/U28/U1/clr ), .a(
        \U1300/s ), .b(\U1300/nback ), .c(bg), .d(bsel) );
    nand3_1 \U1300/U1127/U28/U1/U2  ( .x(\U1300/U1127/U28/U1/set ), .a(bg), 
        .b(\U1300/s ), .c(\U1300/nback ) );
    nand2_2 \U1300/U1127/U28/U1/U3  ( .x(bsel), .a(\U1300/U1127/U28/U1/clr ), 
        .b(\U1300/U1127/U28/U1/set ) );
    aoai211_1 \U1289/U1150/U28/U1/U1  ( .x(\U1289/U1150/U28/U1/clr ), .a(il[2]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdl[2] ) );
    nand3_1 \U1289/U1150/U28/U1/U2  ( .x(\U1289/U1150/U28/U1/set ), .a(net195), 
        .b(il[2]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1150/U28/U1/U3  ( .x(\cdl[2] ), .a(
        \U1289/U1150/U28/U1/clr ), .b(\U1289/U1150/U28/U1/set ) );
    aoai211_1 \U1289/U1152/U28/U1/U1  ( .x(\U1289/U1152/U28/U1/clr ), .a(il[3]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdl[3] ) );
    nand3_1 \U1289/U1152/U28/U1/U2  ( .x(\U1289/U1152/U28/U1/set ), .a(net195), 
        .b(il[3]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1152/U28/U1/U3  ( .x(\cdl[3] ), .a(
        \U1289/U1152/U28/U1/clr ), .b(\U1289/U1152/U28/U1/set ) );
    aoai211_1 \U1289/U1149/U28/U1/U1  ( .x(\U1289/U1149/U28/U1/clr ), .a(ih[2]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdh[2] ) );
    nand3_1 \U1289/U1149/U28/U1/U2  ( .x(\U1289/U1149/U28/U1/set ), .a(net195), 
        .b(ih[2]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1149/U28/U1/U3  ( .x(\cdh[2] ), .a(
        \U1289/U1149/U28/U1/clr ), .b(\U1289/U1149/U28/U1/set ) );
    aoai211_1 \U1289/U1151/U28/U1/U1  ( .x(\U1289/U1151/U28/U1/clr ), .a(ih[3]
        ), .b(\U1289/bnreset ), .c(net195), .d(\cdh[3] ) );
    nand3_1 \U1289/U1151/U28/U1/U2  ( .x(\U1289/U1151/U28/U1/set ), .a(net195), 
        .b(ih[3]), .c(\U1289/bnreset ) );
    nand2_2 \U1289/U1151/U28/U1/U3  ( .x(\cdh[3] ), .a(
        \U1289/U1151/U28/U1/clr ), .b(\U1289/U1151/U28/U1/set ) );
    inv_1 \U1289/U1148/U1147/U3  ( .x(\U1289/U1148/net189 ), .a(
        \U1289/bnreset ) );
    nor2_1 \U1289/U1148/U582/U5  ( .x(\U1289/U1148/net192 ), .a(\cdl[3] ), .b(
        \cdh[3] ) );
    nor2_1 \U1289/U1148/U580/U5  ( .x(\U1289/U1148/net191 ), .a(\cdl[2] ), .b(
        \cdh[2] ) );
    nor2_2 \U1289/U1148/U1146/U6  ( .x(\twobitack[2] ), .a(
        \U1289/U1148/net190 ), .b(\U1289/U1148/net189 ) );
    aoi222_1 \U1289/U1148/U1141/U30/U1  ( .x(\U1289/U1148/net190 ), .a(
        \U1289/U1148/net191 ), .b(\U1289/U1148/net192 ), .c(
        \U1289/U1148/net191 ), .d(\U1289/U1148/U1141/Z ), .e(
        \U1289/U1148/net192 ), .f(\U1289/U1148/U1141/Z ) );
    inv_1 \U1289/U1148/U1141/U30/Uinv  ( .x(\U1289/U1148/U1141/Z ), .a(
        \U1289/U1148/net190 ) );
    aoai211_1 \U1271/U1150/U28/U1/U1  ( .x(\U1271/U1150/U28/U1/clr ), .a(il[0]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdl[0] ) );
    nand3_1 \U1271/U1150/U28/U1/U2  ( .x(\U1271/U1150/U28/U1/set ), .a(net193), 
        .b(il[0]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1150/U28/U1/U3  ( .x(\cdl[0] ), .a(
        \U1271/U1150/U28/U1/clr ), .b(\U1271/U1150/U28/U1/set ) );
    aoai211_1 \U1271/U1152/U28/U1/U1  ( .x(\U1271/U1152/U28/U1/clr ), .a(il[1]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdl[1] ) );
    nand3_1 \U1271/U1152/U28/U1/U2  ( .x(\U1271/U1152/U28/U1/set ), .a(net193), 
        .b(il[1]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1152/U28/U1/U3  ( .x(\cdl[1] ), .a(
        \U1271/U1152/U28/U1/clr ), .b(\U1271/U1152/U28/U1/set ) );
    aoai211_1 \U1271/U1149/U28/U1/U1  ( .x(\U1271/U1149/U28/U1/clr ), .a(ih[0]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdh[0] ) );
    nand3_1 \U1271/U1149/U28/U1/U2  ( .x(\U1271/U1149/U28/U1/set ), .a(net193), 
        .b(ih[0]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1149/U28/U1/U3  ( .x(\cdh[0] ), .a(
        \U1271/U1149/U28/U1/clr ), .b(\U1271/U1149/U28/U1/set ) );
    aoai211_1 \U1271/U1151/U28/U1/U1  ( .x(\U1271/U1151/U28/U1/clr ), .a(ih[1]
        ), .b(\U1271/bnreset ), .c(net193), .d(\cdh[1] ) );
    nand3_1 \U1271/U1151/U28/U1/U2  ( .x(\U1271/U1151/U28/U1/set ), .a(net193), 
        .b(ih[1]), .c(\U1271/bnreset ) );
    nand2_2 \U1271/U1151/U28/U1/U3  ( .x(\cdh[1] ), .a(
        \U1271/U1151/U28/U1/clr ), .b(\U1271/U1151/U28/U1/set ) );
    inv_1 \U1271/U1148/U1147/U3  ( .x(\U1271/U1148/net189 ), .a(
        \U1271/bnreset ) );
    nor2_1 \U1271/U1148/U582/U5  ( .x(\U1271/U1148/net192 ), .a(\cdl[1] ), .b(
        \cdh[1] ) );
    nor2_1 \U1271/U1148/U580/U5  ( .x(\U1271/U1148/net191 ), .a(\cdl[0] ), .b(
        \cdh[0] ) );
    nor2_2 \U1271/U1148/U1146/U6  ( .x(\twobitack[0] ), .a(
        \U1271/U1148/net190 ), .b(\U1271/U1148/net189 ) );
    aoi222_1 \U1271/U1148/U1141/U30/U1  ( .x(\U1271/U1148/net190 ), .a(
        \U1271/U1148/net191 ), .b(\U1271/U1148/net192 ), .c(
        \U1271/U1148/net191 ), .d(\U1271/U1148/U1141/Z ), .e(
        \U1271/U1148/net192 ), .f(\U1271/U1148/U1141/Z ) );
    inv_1 \U1271/U1148/U1141/U30/Uinv  ( .x(\U1271/U1148/U1141/Z ), .a(
        \U1271/U1148/net190 ) );
    nand2_1 \U1225/U1128/U5  ( .x(\U1225/s ), .a(\U1225/r ), .b(\U1225/nback )
         );
    nand2_1 \U1225/U1103/U5  ( .x(\U1225/r ), .a(\U1225/naack ), .b(\U1225/s )
         );
    inv_1 \U1225/U1111/U3  ( .x(\U1225/reset ), .a(nbReset) );
    inv_1 \U1225/U1112/U3  ( .x(\U1225/naack ), .a(nxa) );
    nor2_1 \U1225/U1127/U5  ( .x(\U1225/nback ), .a(nyla), .b(\U1225/reset )
         );
    and2_2 \U1225/U1129/U8  ( .x(xsel), .a(\U1225/nback ), .b(\U1225/s ) );
    and2_2 \U1225/U1124/U8  ( .x(ysel), .a(\U1225/r ), .b(\U1225/naack ) );
    and3_4 \U1308/U20/U9  ( .x(nya), .a(\U1308/nack[1] ), .b(\U1308/nack[0] ), 
        .c(nbReset) );
    nor2_1 \U1308/U18/U5  ( .x(\U1308/nack[0] ), .a(\yl[3] ), .b(\yl[0] ) );
    nor2_1 \U1308/U19/U5  ( .x(\U1308/nack[1] ), .a(\yl[1] ), .b(\yl[2] ) );
    ao222_2 \U1308/U15_0_/U19/U1/U1  ( .x(\yl[0] ), .a(\y[0] ), .b(nyla), .c(
        \y[0] ), .d(\yl[0] ), .e(nyla), .f(\yl[0] ) );
    ao222_2 \U1308/U15_1_/U19/U1/U1  ( .x(\yl[1] ), .a(\y[1] ), .b(nyla), .c(
        \y[1] ), .d(\yl[1] ), .e(nyla), .f(\yl[1] ) );
    ao222_2 \U1308/U15_2_/U19/U1/U1  ( .x(\yl[2] ), .a(\y[2] ), .b(nyla), .c(
        \y[2] ), .d(\yl[2] ), .e(nyla), .f(\yl[2] ) );
    ao222_2 \U1308/U15_3_/U19/U1/U1  ( .x(\yl[3] ), .a(\y[3] ), .b(nyla), .c(
        \y[3] ), .d(\yl[3] ), .e(nyla), .f(\yl[3] ) );
    buf_3 U1 ( .x(\U1271/bnreset ), .a(nbReset) );
    buf_3 U2 ( .x(\U1289/bnreset ), .a(nbReset) );
endmodule


module chain_mergepackets_4 ( naa, nba, o, a, b, nReset, noa );
output [4:0] o;
input  [4:0] a;
input  [4:0] b;
input  nReset, noa;
output naa, nba;
    wire as, seta, asel, bsel, setb, reset, \noack[1] , \noack[0] , 
        \U916_0_/U25/U1/clr , \U916_0_/U25/U1/ob , \U916_1_/U25/U1/clr , 
        \U916_1_/U25/U1/ob , \U916_2_/U25/U1/clr , \U916_2_/U25/U1/ob , 
        \U916_3_/U25/U1/clr , \U916_3_/U25/U1/ob ;
    and2_1 \U1155/U8  ( .x(as), .a(seta), .b(asel) );
    nand2_1 \U1145/U5  ( .x(asel), .a(bsel), .b(seta) );
    nand2_1 \U1103/U5  ( .x(bsel), .a(setb), .b(asel) );
    inv_1 \U1135/U3  ( .x(reset), .a(nReset) );
    inv_1 \U1134/U3  ( .x(setb), .a(a[4]) );
    and3_2 \U1154/U9  ( .x(naa), .a(\noack[1] ), .b(\noack[0] ), .c(as) );
    nor3_1 \U1127/U7  ( .x(\noack[0] ), .a(o[1]), .b(reset), .c(o[0]) );
    nor2_1 \U1132/U5  ( .x(\noack[1] ), .a(o[3]), .b(o[2]) );
    oa31_1 \U916_0_/U25/U1/Uclr  ( .x(\U916_0_/U25/U1/clr ), .a(noa), .b(a[0]), 
        .c(b[0]), .d(o[0]) );
    oaoi211_1 \U916_0_/U25/U1/Uaoi  ( .x(\U916_0_/U25/U1/ob ), .a(a[0]), .b(b
        [0]), .c(noa), .d(\U916_0_/U25/U1/clr ) );
    inv_2 \U916_0_/U25/U1/Ui  ( .x(o[0]), .a(\U916_0_/U25/U1/ob ) );
    oa31_1 \U916_1_/U25/U1/Uclr  ( .x(\U916_1_/U25/U1/clr ), .a(noa), .b(a[1]), 
        .c(b[1]), .d(o[1]) );
    oaoi211_1 \U916_1_/U25/U1/Uaoi  ( .x(\U916_1_/U25/U1/ob ), .a(a[1]), .b(b
        [1]), .c(noa), .d(\U916_1_/U25/U1/clr ) );
    inv_2 \U916_1_/U25/U1/Ui  ( .x(o[1]), .a(\U916_1_/U25/U1/ob ) );
    oa31_1 \U916_2_/U25/U1/Uclr  ( .x(\U916_2_/U25/U1/clr ), .a(noa), .b(a[2]), 
        .c(b[2]), .d(o[2]) );
    oaoi211_1 \U916_2_/U25/U1/Uaoi  ( .x(\U916_2_/U25/U1/ob ), .a(a[2]), .b(b
        [2]), .c(noa), .d(\U916_2_/U25/U1/clr ) );
    inv_2 \U916_2_/U25/U1/Ui  ( .x(o[2]), .a(\U916_2_/U25/U1/ob ) );
    oa31_1 \U916_3_/U25/U1/Uclr  ( .x(\U916_3_/U25/U1/clr ), .a(noa), .b(a[3]), 
        .c(b[3]), .d(o[3]) );
    oaoi211_1 \U916_3_/U25/U1/Uaoi  ( .x(\U916_3_/U25/U1/ob ), .a(a[3]), .b(b
        [3]), .c(noa), .d(\U916_3_/U25/U1/clr ) );
    inv_2 \U916_3_/U25/U1/Ui  ( .x(o[3]), .a(\U916_3_/U25/U1/ob ) );
    ao222_2 \U1148/U19/U1/U1  ( .x(o[4]), .a(noa), .b(b[4]), .c(noa), .d(o[4]), 
        .e(b[4]), .f(o[4]) );
    aoi21_1 \U1153/U11  ( .x(seta), .a(o[4]), .b(setb), .c(reset) );
    and3_3 U1 ( .x(nba), .a(bsel), .b(\noack[0] ), .c(\noack[1] ) );
endmodule


module chain_tchdr_1 ( addr_req, col_h, col_l, itag_h, itag_l, lock, ncback, 
    neop, pred, pullcd, reset, rnw_h, rnw_l, seq, size_h, size_l, write_req, 
    chwh, chwl, addr_ack, addr_pull, nReset, nack, write_ack, write_pull );
output [2:0] col_h;
output [2:0] col_l;
output [4:0] itag_h;
output [4:0] itag_l;
output [1:0] lock;
output [1:0] pred;
output [1:0] seq;
output [1:0] size_h;
output [1:0] size_l;
input  [7:0] chwh;
input  [7:0] chwl;
input  addr_ack, addr_pull, nReset, nack, write_ack, write_pull;
output addr_req, ncback, neop, pullcd, reset, rnw_h, rnw_l, write_req;
    wire n9, pullcdwk, net94, net88, \ncd[0] , \ncd[1] , \ncd[2] , \ncd[3] , 
        \ncd[4] , \ncd[5] , \ncd[6] , \ncd[7] , read, ack, net83, \U1664/x[3] , 
        \U1664/U28/Z , \U1664/x[0] , \U1664/U32/Z , \U1664/x[2] , 
        \U1664/U29/Z , \U1664/y[0] , \U1664/x[1] , \U1664/U33/Z , \U1664/y[1] , 
        \U1664/U30/Z , \U1664/U31/Z , \U1664/U37/Z , receive, \U473/Z , 
        \hdr_hld/net32 , \hdr_hld/net33 , \hdr_hld/low/latch , 
        \hdr_hld/low/nlocalcd , \hdr_hld/low/localcd , \hdr_hld/low/ncd[0] , 
        \hdr_hld/low/ncd[1] , \hdr_hld/low/ncd[2] , \hdr_hld/low/ncd[3] , 
        \hdr_hld/ol[3] , \hdr_hld/oh[3] , \hdr_hld/low/ncd[4] , 
        \hdr_hld/ol[4] , \hdr_hld/oh[4] , \hdr_hld/low/ncd[5] , 
        \hdr_hld/low/ncd[6] , \hdr_hld/low/ncd[7] , 
        \hdr_hld/low/ctrlack_internal , \hdr_hld/low/acb , \hdr_hld/low/ba , 
        \hdr_hld/low/driveh , \hdr_hld/net20 , \hdr_hld/low/drivel , n2, n3, 
        n1, \hdr_hld/low/U4/U28/U1/clr , \hdr_hld/low/U4/U28/U1/set , 
        \hdr_hld/low/U1/Z , \hdr_hld/low/U1664/x[3] , 
        \hdr_hld/low/U1664/U28/Z , \hdr_hld/low/U1664/x[0] , 
        \hdr_hld/low/U1664/U32/Z , \hdr_hld/low/U1664/x[2] , 
        \hdr_hld/low/U1664/U29/Z , \hdr_hld/low/U1664/y[0] , 
        \hdr_hld/low/U1664/x[1] , \hdr_hld/low/U1664/U33/Z , 
        \hdr_hld/low/U1664/y[1] , \hdr_hld/low/U1664/U30/Z , 
        \hdr_hld/low/U1664/U31/Z , \hdr_hld/low/U1664/U37/Z , 
        \hdr_hld/low/U1669/nr , \hdr_hld/low/U1669/nd , \hdr_hld/low/U1669/n2 , 
        \hdr_hld/high/latch , \hdr_hld/high/nlocalcd , \hdr_hld/high/localcd , 
        \hdr_hld/high/ncd[0] , \hdr_hld/high/ncd[1] , \hdr_hld/high/ncd[2] , 
        \hdr_hld/high/ncd[3] , \hdr_hld/high/ncd[4] , \hdr_hld/high/ncd[5] , 
        \hdr_hld/high/ncd[6] , \hdr_hld/high/ncd[7] , 
        \hdr_hld/high/ctrlack_internal , \hdr_hld/high/acb , \hdr_hld/high/ba , 
        \hdr_hld/high/driveh , \hdr_hld/high/drivel , n7, n4, n5, n6, 
        \hdr_hld/high/U4/U28/U1/clr , \hdr_hld/high/U4/U28/U1/set , 
        \hdr_hld/high/U1/Z , \hdr_hld/high/U1664/x[3] , 
        \hdr_hld/high/U1664/U28/Z , \hdr_hld/high/U1664/x[0] , 
        \hdr_hld/high/U1664/U32/Z , \hdr_hld/high/U1664/x[2] , 
        \hdr_hld/high/U1664/U29/Z , \hdr_hld/high/U1664/y[0] , 
        \hdr_hld/high/U1664/x[1] , \hdr_hld/high/U1664/U33/Z , 
        \hdr_hld/high/U1664/y[1] , \hdr_hld/high/U1664/U30/Z , 
        \hdr_hld/high/U1664/U31/Z , \hdr_hld/high/U1664/U37/Z , 
        \hdr_hld/high/U1669/nr , \hdr_hld/high/U1669/nd , 
        \hdr_hld/high/U1669/n2 ;
    buf_1 U262 ( .x(n9), .a(pullcdwk) );
    or3_2 \U1668/U12  ( .x(ncback), .a(net94), .b(addr_pull), .c(write_pull)
         );
    inv_1 \I0/U3  ( .x(net94), .a(net88) );
    nor2_1 \U514_0_/U5  ( .x(\ncd[0] ), .a(chwh[0]), .b(chwl[0]) );
    nor2_1 \U514_1_/U5  ( .x(\ncd[1] ), .a(chwh[1]), .b(chwl[1]) );
    nor2_1 \U514_2_/U5  ( .x(\ncd[2] ), .a(chwh[2]), .b(chwl[2]) );
    nor2_1 \U514_3_/U5  ( .x(\ncd[3] ), .a(chwh[3]), .b(chwl[3]) );
    nor2_1 \U514_4_/U5  ( .x(\ncd[4] ), .a(chwh[4]), .b(chwl[4]) );
    nor2_1 \U514_5_/U5  ( .x(\ncd[5] ), .a(chwh[5]), .b(chwl[5]) );
    nor2_1 \U514_6_/U5  ( .x(\ncd[6] ), .a(chwh[6]), .b(chwl[6]) );
    nor2_1 \U514_7_/U5  ( .x(\ncd[7] ), .a(chwh[7]), .b(chwl[7]) );
    nor2_1 \U1669/U5  ( .x(neop), .a(read), .b(write_ack) );
    nand2_1 \U303/U5  ( .x(ack), .a(nack), .b(nReset) );
    nand2_1 \U1670/U5  ( .x(net83), .a(neop), .b(nReset) );
    ao222_1 \U47/U18/U1/U1  ( .x(read), .a(addr_ack), .b(rnw_h), .c(addr_ack), 
        .d(read), .e(rnw_h), .f(read) );
    ao222_1 \U48/U18/U1/U1  ( .x(write_req), .a(rnw_l), .b(addr_ack), .c(rnw_l
        ), .d(write_req), .e(addr_ack), .f(write_req) );
    aoi222_1 \U1664/U28/U30/U1  ( .x(\U1664/x[3] ), .a(\ncd[7] ), .b(\ncd[6] ), 
        .c(\ncd[7] ), .d(\U1664/U28/Z ), .e(\ncd[6] ), .f(\U1664/U28/Z ) );
    inv_1 \U1664/U28/U30/Uinv  ( .x(\U1664/U28/Z ), .a(\U1664/x[3] ) );
    aoi222_1 \U1664/U32/U30/U1  ( .x(\U1664/x[0] ), .a(\ncd[1] ), .b(\ncd[0] ), 
        .c(\ncd[1] ), .d(\U1664/U32/Z ), .e(\ncd[0] ), .f(\U1664/U32/Z ) );
    inv_1 \U1664/U32/U30/Uinv  ( .x(\U1664/U32/Z ), .a(\U1664/x[0] ) );
    aoi222_1 \U1664/U29/U30/U1  ( .x(\U1664/x[2] ), .a(\ncd[5] ), .b(\ncd[4] ), 
        .c(\ncd[5] ), .d(\U1664/U29/Z ), .e(\ncd[4] ), .f(\U1664/U29/Z ) );
    inv_1 \U1664/U29/U30/Uinv  ( .x(\U1664/U29/Z ), .a(\U1664/x[2] ) );
    aoi222_1 \U1664/U33/U30/U1  ( .x(\U1664/y[0] ), .a(\U1664/x[1] ), .b(
        \U1664/x[0] ), .c(\U1664/x[1] ), .d(\U1664/U33/Z ), .e(\U1664/x[0] ), 
        .f(\U1664/U33/Z ) );
    inv_1 \U1664/U33/U30/Uinv  ( .x(\U1664/U33/Z ), .a(\U1664/y[0] ) );
    aoi222_1 \U1664/U30/U30/U1  ( .x(\U1664/y[1] ), .a(\U1664/x[3] ), .b(
        \U1664/x[2] ), .c(\U1664/x[3] ), .d(\U1664/U30/Z ), .e(\U1664/x[2] ), 
        .f(\U1664/U30/Z ) );
    inv_1 \U1664/U30/U30/Uinv  ( .x(\U1664/U30/Z ), .a(\U1664/y[1] ) );
    aoi222_1 \U1664/U31/U30/U1  ( .x(\U1664/x[1] ), .a(\ncd[3] ), .b(\ncd[2] ), 
        .c(\ncd[3] ), .d(\U1664/U31/Z ), .e(\ncd[2] ), .f(\U1664/U31/Z ) );
    inv_1 \U1664/U31/U30/Uinv  ( .x(\U1664/U31/Z ), .a(\U1664/x[1] ) );
    aoi222_1 \U1664/U37/U30/U1  ( .x(pullcdwk), .a(\U1664/y[0] ), .b(
        \U1664/y[1] ), .c(\U1664/y[0] ), .d(\U1664/U37/Z ), .e(\U1664/y[1] ), 
        .f(\U1664/U37/Z ) );
    inv_1 \U1664/U37/U30/Uinv  ( .x(\U1664/U37/Z ), .a(pullcdwk) );
    aoi222_1 \U473/U30/U1  ( .x(receive), .a(net83), .b(ack), .c(net83), .d(
        \U473/Z ), .e(ack), .f(\U473/Z ) );
    inv_1 \U473/U30/Uinv  ( .x(\U473/Z ), .a(receive) );
    nor2_1 \hdr_hld/U3/U5  ( .x(net88), .a(\hdr_hld/net32 ), .b(
        \hdr_hld/net33 ) );
    buf_2 \hdr_hld/low/U1653  ( .x(\hdr_hld/low/latch ), .a(\hdr_hld/net32 )
         );
    nor2_1 \hdr_hld/low/U264/U5  ( .x(\hdr_hld/low/nlocalcd ), .a(reset), .b(
        \hdr_hld/low/localcd ) );
    nor2_1 \hdr_hld/low/U1659_0_/U5  ( .x(\hdr_hld/low/ncd[0] ), .a(seq[0]), 
        .b(seq[1]) );
    nor2_1 \hdr_hld/low/U1659_1_/U5  ( .x(\hdr_hld/low/ncd[1] ), .a(pred[0]), 
        .b(pred[1]) );
    nor2_1 \hdr_hld/low/U1659_2_/U5  ( .x(\hdr_hld/low/ncd[2] ), .a(lock[0]), 
        .b(lock[1]) );
    nor2_1 \hdr_hld/low/U1659_3_/U5  ( .x(\hdr_hld/low/ncd[3] ), .a(
        \hdr_hld/ol[3] ), .b(\hdr_hld/oh[3] ) );
    nor2_1 \hdr_hld/low/U1659_4_/U5  ( .x(\hdr_hld/low/ncd[4] ), .a(
        \hdr_hld/ol[4] ), .b(\hdr_hld/oh[4] ) );
    nor2_1 \hdr_hld/low/U1659_5_/U5  ( .x(\hdr_hld/low/ncd[5] ), .a(rnw_l), 
        .b(rnw_h) );
    nor2_1 \hdr_hld/low/U1659_6_/U5  ( .x(\hdr_hld/low/ncd[6] ), .a(size_l[0]), 
        .b(size_h[0]) );
    nor2_1 \hdr_hld/low/U1659_7_/U5  ( .x(\hdr_hld/low/ncd[7] ), .a(size_l[1]), 
        .b(size_h[1]) );
    nor2_1 \hdr_hld/low/U3/U5  ( .x(\hdr_hld/low/ctrlack_internal ), .a(
        \hdr_hld/low/acb ), .b(\hdr_hld/low/ba ) );
    buf_2 \hdr_hld/low/U1665/U7  ( .x(\hdr_hld/low/driveh ), .a(
        \hdr_hld/net20 ) );
    buf_2 \hdr_hld/low/U1666/U7  ( .x(\hdr_hld/low/drivel ), .a(
        \hdr_hld/net20 ) );
    ao23_1 \hdr_hld/low/U1658_0_/U21/U1/U1  ( .x(seq[0]), .a(n2), .b(seq[0]), 
        .c(\hdr_hld/low/drivel ), .d(chwl[0]), .e(n3) );
    ao23_1 \hdr_hld/low/U1658_1_/U21/U1/U1  ( .x(pred[0]), .a(n1), .b(pred[0]), 
        .c(\hdr_hld/low/drivel ), .d(chwl[1]), .e(n3) );
    ao23_1 \hdr_hld/low/U1658_2_/U21/U1/U1  ( .x(lock[0]), .a(n1), .b(lock[0]), 
        .c(\hdr_hld/low/driveh ), .d(chwl[2]), .e(n3) );
    ao23_1 \hdr_hld/low/U1658_3_/U21/U1/U1  ( .x(\hdr_hld/ol[3] ), .a(n1), .b(
        \hdr_hld/ol[3] ), .c(\hdr_hld/low/driveh ), .d(chwl[3]), .e(
        \hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1658_4_/U21/U1/U1  ( .x(\hdr_hld/ol[4] ), .a(n2), .b(
        \hdr_hld/ol[4] ), .c(\hdr_hld/low/drivel ), .d(chwl[4]), .e(
        \hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1658_5_/U21/U1/U1  ( .x(rnw_l), .a(
        \hdr_hld/low/driveh ), .b(rnw_l), .c(\hdr_hld/low/driveh ), .d(chwl[5]
        ), .e(\hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1658_6_/U21/U1/U1  ( .x(size_l[0]), .a(
        \hdr_hld/low/drivel ), .b(size_l[0]), .c(n2), .d(chwl[6]), .e(
        \hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1658_7_/U21/U1/U1  ( .x(size_l[1]), .a(
        \hdr_hld/low/drivel ), .b(size_l[1]), .c(\hdr_hld/low/drivel ), .d(
        chwl[7]), .e(\hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1651_0_/U21/U1/U1  ( .x(seq[1]), .a(
        \hdr_hld/low/drivel ), .b(seq[1]), .c(\hdr_hld/low/driveh ), .d(chwh
        [0]), .e(\hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1651_1_/U21/U1/U1  ( .x(pred[1]), .a(
        \hdr_hld/low/driveh ), .b(pred[1]), .c(n1), .d(chwh[1]), .e(
        \hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1651_2_/U21/U1/U1  ( .x(lock[1]), .a(
        \hdr_hld/low/driveh ), .b(lock[1]), .c(n1), .d(chwh[2]), .e(
        \hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1651_3_/U21/U1/U1  ( .x(\hdr_hld/oh[3] ), .a(
        \hdr_hld/low/drivel ), .b(\hdr_hld/oh[3] ), .c(n2), .d(chwh[3]), .e(
        \hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1651_4_/U21/U1/U1  ( .x(\hdr_hld/oh[4] ), .a(n2), .b(
        \hdr_hld/oh[4] ), .c(n1), .d(chwh[4]), .e(\hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1651_5_/U21/U1/U1  ( .x(rnw_h), .a(n2), .b(rnw_h), 
        .c(n1), .d(chwh[5]), .e(\hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1651_6_/U21/U1/U1  ( .x(size_h[0]), .a(n1), .b(size_h
        [0]), .c(n2), .d(chwh[6]), .e(\hdr_hld/low/latch ) );
    ao23_1 \hdr_hld/low/U1651_7_/U21/U1/U1  ( .x(size_h[1]), .a(
        \hdr_hld/low/driveh ), .b(size_h[1]), .c(n2), .d(chwh[7]), .e(
        \hdr_hld/low/latch ) );
    aoai211_1 \hdr_hld/low/U4/U28/U1/U1  ( .x(\hdr_hld/low/U4/U28/U1/clr ), 
        .a(\hdr_hld/net20 ), .b(\hdr_hld/low/acb ), .c(\hdr_hld/low/nlocalcd ), 
        .d(\hdr_hld/net32 ) );
    nand3_1 \hdr_hld/low/U4/U28/U1/U2  ( .x(\hdr_hld/low/U4/U28/U1/set ), .a(
        \hdr_hld/low/nlocalcd ), .b(\hdr_hld/net20 ), .c(\hdr_hld/low/acb ) );
    nand2_2 \hdr_hld/low/U4/U28/U1/U3  ( .x(\hdr_hld/net32 ), .a(
        \hdr_hld/low/U4/U28/U1/clr ), .b(\hdr_hld/low/U4/U28/U1/set ) );
    oai21_1 \hdr_hld/low/U1/U30/U1/U1  ( .x(\hdr_hld/low/acb ), .a(
        \hdr_hld/low/U1/Z ), .b(\hdr_hld/low/ba ), .c(\hdr_hld/net20 ) );
    inv_1 \hdr_hld/low/U1/U30/U1/U2  ( .x(\hdr_hld/low/U1/Z ), .a(
        \hdr_hld/low/acb ) );
    ao222_1 \hdr_hld/low/U5/U18/U1/U1  ( .x(\hdr_hld/low/ba ), .a(
        \hdr_hld/low/latch ), .b(n9), .c(\hdr_hld/low/latch ), .d(
        \hdr_hld/low/ba ), .e(n9), .f(\hdr_hld/low/ba ) );
    aoi222_1 \hdr_hld/low/U1664/U28/U30/U1  ( .x(\hdr_hld/low/U1664/x[3] ), 
        .a(\hdr_hld/low/ncd[7] ), .b(\hdr_hld/low/ncd[6] ), .c(
        \hdr_hld/low/ncd[7] ), .d(\hdr_hld/low/U1664/U28/Z ), .e(
        \hdr_hld/low/ncd[6] ), .f(\hdr_hld/low/U1664/U28/Z ) );
    inv_1 \hdr_hld/low/U1664/U28/U30/Uinv  ( .x(\hdr_hld/low/U1664/U28/Z ), 
        .a(\hdr_hld/low/U1664/x[3] ) );
    aoi222_1 \hdr_hld/low/U1664/U32/U30/U1  ( .x(\hdr_hld/low/U1664/x[0] ), 
        .a(\hdr_hld/low/ncd[1] ), .b(\hdr_hld/low/ncd[0] ), .c(
        \hdr_hld/low/ncd[1] ), .d(\hdr_hld/low/U1664/U32/Z ), .e(
        \hdr_hld/low/ncd[0] ), .f(\hdr_hld/low/U1664/U32/Z ) );
    inv_1 \hdr_hld/low/U1664/U32/U30/Uinv  ( .x(\hdr_hld/low/U1664/U32/Z ), 
        .a(\hdr_hld/low/U1664/x[0] ) );
    aoi222_1 \hdr_hld/low/U1664/U29/U30/U1  ( .x(\hdr_hld/low/U1664/x[2] ), 
        .a(\hdr_hld/low/ncd[5] ), .b(\hdr_hld/low/ncd[4] ), .c(
        \hdr_hld/low/ncd[5] ), .d(\hdr_hld/low/U1664/U29/Z ), .e(
        \hdr_hld/low/ncd[4] ), .f(\hdr_hld/low/U1664/U29/Z ) );
    inv_1 \hdr_hld/low/U1664/U29/U30/Uinv  ( .x(\hdr_hld/low/U1664/U29/Z ), 
        .a(\hdr_hld/low/U1664/x[2] ) );
    aoi222_1 \hdr_hld/low/U1664/U33/U30/U1  ( .x(\hdr_hld/low/U1664/y[0] ), 
        .a(\hdr_hld/low/U1664/x[1] ), .b(\hdr_hld/low/U1664/x[0] ), .c(
        \hdr_hld/low/U1664/x[1] ), .d(\hdr_hld/low/U1664/U33/Z ), .e(
        \hdr_hld/low/U1664/x[0] ), .f(\hdr_hld/low/U1664/U33/Z ) );
    inv_1 \hdr_hld/low/U1664/U33/U30/Uinv  ( .x(\hdr_hld/low/U1664/U33/Z ), 
        .a(\hdr_hld/low/U1664/y[0] ) );
    aoi222_1 \hdr_hld/low/U1664/U30/U30/U1  ( .x(\hdr_hld/low/U1664/y[1] ), 
        .a(\hdr_hld/low/U1664/x[3] ), .b(\hdr_hld/low/U1664/x[2] ), .c(
        \hdr_hld/low/U1664/x[3] ), .d(\hdr_hld/low/U1664/U30/Z ), .e(
        \hdr_hld/low/U1664/x[2] ), .f(\hdr_hld/low/U1664/U30/Z ) );
    inv_1 \hdr_hld/low/U1664/U30/U30/Uinv  ( .x(\hdr_hld/low/U1664/U30/Z ), 
        .a(\hdr_hld/low/U1664/y[1] ) );
    aoi222_1 \hdr_hld/low/U1664/U31/U30/U1  ( .x(\hdr_hld/low/U1664/x[1] ), 
        .a(\hdr_hld/low/ncd[3] ), .b(\hdr_hld/low/ncd[2] ), .c(
        \hdr_hld/low/ncd[3] ), .d(\hdr_hld/low/U1664/U31/Z ), .e(
        \hdr_hld/low/ncd[2] ), .f(\hdr_hld/low/U1664/U31/Z ) );
    inv_1 \hdr_hld/low/U1664/U31/U30/Uinv  ( .x(\hdr_hld/low/U1664/U31/Z ), 
        .a(\hdr_hld/low/U1664/x[1] ) );
    aoi222_1 \hdr_hld/low/U1664/U37/U30/U1  ( .x(\hdr_hld/low/localcd ), .a(
        \hdr_hld/low/U1664/y[0] ), .b(\hdr_hld/low/U1664/y[1] ), .c(
        \hdr_hld/low/U1664/y[0] ), .d(\hdr_hld/low/U1664/U37/Z ), .e(
        \hdr_hld/low/U1664/y[1] ), .f(\hdr_hld/low/U1664/U37/Z ) );
    inv_1 \hdr_hld/low/U1664/U37/U30/Uinv  ( .x(\hdr_hld/low/U1664/U37/Z ), 
        .a(\hdr_hld/low/localcd ) );
    nor3_1 \hdr_hld/low/U1669/Unr  ( .x(\hdr_hld/low/U1669/nr ), .a(
        \hdr_hld/low/ctrlack_internal ), .b(\hdr_hld/low/driveh ), .c(n1) );
    nand3_1 \hdr_hld/low/U1669/Und  ( .x(\hdr_hld/low/U1669/nd ), .a(
        \hdr_hld/low/ctrlack_internal ), .b(n2), .c(\hdr_hld/low/drivel ) );
    oa21_1 \hdr_hld/low/U1669/U1  ( .x(\hdr_hld/low/U1669/n2 ), .a(
        \hdr_hld/low/U1669/n2 ), .b(\hdr_hld/low/U1669/nr ), .c(
        \hdr_hld/low/U1669/nd ) );
    inv_2 \hdr_hld/low/U1669/U3  ( .x(addr_req), .a(\hdr_hld/low/U1669/n2 ) );
    buf_2 \hdr_hld/high/U1653  ( .x(\hdr_hld/high/latch ), .a(\hdr_hld/net33 )
         );
    nor2_1 \hdr_hld/high/U264/U5  ( .x(\hdr_hld/high/nlocalcd ), .a(reset), 
        .b(\hdr_hld/high/localcd ) );
    nor2_1 \hdr_hld/high/U1659_0_/U5  ( .x(\hdr_hld/high/ncd[0] ), .a(itag_l
        [0]), .b(itag_h[0]) );
    nor2_1 \hdr_hld/high/U1659_1_/U5  ( .x(\hdr_hld/high/ncd[1] ), .a(itag_l
        [1]), .b(itag_h[1]) );
    nor2_1 \hdr_hld/high/U1659_2_/U5  ( .x(\hdr_hld/high/ncd[2] ), .a(itag_l
        [2]), .b(itag_h[2]) );
    nor2_1 \hdr_hld/high/U1659_3_/U5  ( .x(\hdr_hld/high/ncd[3] ), .a(itag_l
        [3]), .b(itag_h[3]) );
    nor2_1 \hdr_hld/high/U1659_4_/U5  ( .x(\hdr_hld/high/ncd[4] ), .a(itag_l
        [4]), .b(itag_h[4]) );
    nor2_1 \hdr_hld/high/U1659_5_/U5  ( .x(\hdr_hld/high/ncd[5] ), .a(col_l[0]
        ), .b(col_h[0]) );
    nor2_1 \hdr_hld/high/U1659_6_/U5  ( .x(\hdr_hld/high/ncd[6] ), .a(col_l[1]
        ), .b(col_h[1]) );
    nor2_1 \hdr_hld/high/U1659_7_/U5  ( .x(\hdr_hld/high/ncd[7] ), .a(col_l[2]
        ), .b(col_h[2]) );
    nor2_1 \hdr_hld/high/U3/U5  ( .x(\hdr_hld/high/ctrlack_internal ), .a(
        \hdr_hld/high/acb ), .b(\hdr_hld/high/ba ) );
    buf_2 \hdr_hld/high/U1665/U7  ( .x(\hdr_hld/high/driveh ), .a(receive) );
    buf_2 \hdr_hld/high/U1666/U7  ( .x(\hdr_hld/high/drivel ), .a(receive) );
    ao23_1 \hdr_hld/high/U1658_0_/U21/U1/U1  ( .x(itag_l[0]), .a(
        \hdr_hld/high/drivel ), .b(itag_l[0]), .c(\hdr_hld/high/drivel ), .d(
        chwl[0]), .e(n7) );
    ao23_1 \hdr_hld/high/U1658_1_/U21/U1/U1  ( .x(itag_l[1]), .a(
        \hdr_hld/high/drivel ), .b(itag_l[1]), .c(\hdr_hld/high/drivel ), .d(
        chwl[1]), .e(n7) );
    ao23_1 \hdr_hld/high/U1658_2_/U21/U1/U1  ( .x(itag_l[2]), .a(
        \hdr_hld/high/drivel ), .b(itag_l[2]), .c(\hdr_hld/high/drivel ), .d(
        chwl[2]), .e(n7) );
    ao23_1 \hdr_hld/high/U1658_3_/U21/U1/U1  ( .x(itag_l[3]), .a(
        \hdr_hld/high/drivel ), .b(itag_l[3]), .c(\hdr_hld/high/drivel ), .d(
        chwl[3]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1658_4_/U21/U1/U1  ( .x(itag_l[4]), .a(n4), .b(
        itag_l[4]), .c(\hdr_hld/high/drivel ), .d(chwl[4]), .e(
        \hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1658_5_/U21/U1/U1  ( .x(col_l[0]), .a(n4), .b(col_l
        [0]), .c(\hdr_hld/high/drivel ), .d(chwl[5]), .e(\hdr_hld/high/latch )
         );
    ao23_1 \hdr_hld/high/U1658_6_/U21/U1/U1  ( .x(col_l[1]), .a(
        \hdr_hld/high/drivel ), .b(col_l[1]), .c(\hdr_hld/high/drivel ), .d(
        chwl[6]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1658_7_/U21/U1/U1  ( .x(col_l[2]), .a(n4), .b(col_l
        [2]), .c(\hdr_hld/high/drivel ), .d(chwl[7]), .e(\hdr_hld/high/latch )
         );
    ao23_1 \hdr_hld/high/U1651_0_/U21/U1/U1  ( .x(itag_h[0]), .a(n5), .b(
        itag_h[0]), .c(n5), .d(chwh[0]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1651_1_/U21/U1/U1  ( .x(itag_h[1]), .a(n5), .b(
        itag_h[1]), .c(n6), .d(chwh[1]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1651_2_/U21/U1/U1  ( .x(itag_h[2]), .a(n5), .b(
        itag_h[2]), .c(n6), .d(chwh[2]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1651_3_/U21/U1/U1  ( .x(itag_h[3]), .a(n5), .b(
        itag_h[3]), .c(n6), .d(chwh[3]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1651_4_/U21/U1/U1  ( .x(itag_h[4]), .a(n5), .b(
        itag_h[4]), .c(n6), .d(chwh[4]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1651_5_/U21/U1/U1  ( .x(col_h[0]), .a(n5), .b(col_h
        [0]), .c(n6), .d(chwh[5]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1651_6_/U21/U1/U1  ( .x(col_h[1]), .a(n5), .b(col_h
        [1]), .c(n5), .d(chwh[6]), .e(\hdr_hld/high/latch ) );
    ao23_1 \hdr_hld/high/U1651_7_/U21/U1/U1  ( .x(col_h[2]), .a(n5), .b(col_h
        [2]), .c(n5), .d(chwh[7]), .e(\hdr_hld/high/latch ) );
    aoai211_1 \hdr_hld/high/U4/U28/U1/U1  ( .x(\hdr_hld/high/U4/U28/U1/clr ), 
        .a(receive), .b(\hdr_hld/high/acb ), .c(\hdr_hld/high/nlocalcd ), .d(
        \hdr_hld/net33 ) );
    nand3_1 \hdr_hld/high/U4/U28/U1/U2  ( .x(\hdr_hld/high/U4/U28/U1/set ), 
        .a(\hdr_hld/high/nlocalcd ), .b(receive), .c(\hdr_hld/high/acb ) );
    nand2_2 \hdr_hld/high/U4/U28/U1/U3  ( .x(\hdr_hld/net33 ), .a(
        \hdr_hld/high/U4/U28/U1/clr ), .b(\hdr_hld/high/U4/U28/U1/set ) );
    oai21_1 \hdr_hld/high/U1/U30/U1/U1  ( .x(\hdr_hld/high/acb ), .a(
        \hdr_hld/high/U1/Z ), .b(\hdr_hld/high/ba ), .c(receive) );
    inv_1 \hdr_hld/high/U1/U30/U1/U2  ( .x(\hdr_hld/high/U1/Z ), .a(
        \hdr_hld/high/acb ) );
    ao222_1 \hdr_hld/high/U5/U18/U1/U1  ( .x(\hdr_hld/high/ba ), .a(
        \hdr_hld/high/latch ), .b(n9), .c(\hdr_hld/high/latch ), .d(
        \hdr_hld/high/ba ), .e(n9), .f(\hdr_hld/high/ba ) );
    aoi222_1 \hdr_hld/high/U1664/U28/U30/U1  ( .x(\hdr_hld/high/U1664/x[3] ), 
        .a(\hdr_hld/high/ncd[7] ), .b(\hdr_hld/high/ncd[6] ), .c(
        \hdr_hld/high/ncd[7] ), .d(\hdr_hld/high/U1664/U28/Z ), .e(
        \hdr_hld/high/ncd[6] ), .f(\hdr_hld/high/U1664/U28/Z ) );
    inv_1 \hdr_hld/high/U1664/U28/U30/Uinv  ( .x(\hdr_hld/high/U1664/U28/Z ), 
        .a(\hdr_hld/high/U1664/x[3] ) );
    aoi222_1 \hdr_hld/high/U1664/U32/U30/U1  ( .x(\hdr_hld/high/U1664/x[0] ), 
        .a(\hdr_hld/high/ncd[1] ), .b(\hdr_hld/high/ncd[0] ), .c(
        \hdr_hld/high/ncd[1] ), .d(\hdr_hld/high/U1664/U32/Z ), .e(
        \hdr_hld/high/ncd[0] ), .f(\hdr_hld/high/U1664/U32/Z ) );
    inv_1 \hdr_hld/high/U1664/U32/U30/Uinv  ( .x(\hdr_hld/high/U1664/U32/Z ), 
        .a(\hdr_hld/high/U1664/x[0] ) );
    aoi222_1 \hdr_hld/high/U1664/U29/U30/U1  ( .x(\hdr_hld/high/U1664/x[2] ), 
        .a(\hdr_hld/high/ncd[5] ), .b(\hdr_hld/high/ncd[4] ), .c(
        \hdr_hld/high/ncd[5] ), .d(\hdr_hld/high/U1664/U29/Z ), .e(
        \hdr_hld/high/ncd[4] ), .f(\hdr_hld/high/U1664/U29/Z ) );
    inv_1 \hdr_hld/high/U1664/U29/U30/Uinv  ( .x(\hdr_hld/high/U1664/U29/Z ), 
        .a(\hdr_hld/high/U1664/x[2] ) );
    aoi222_1 \hdr_hld/high/U1664/U33/U30/U1  ( .x(\hdr_hld/high/U1664/y[0] ), 
        .a(\hdr_hld/high/U1664/x[1] ), .b(\hdr_hld/high/U1664/x[0] ), .c(
        \hdr_hld/high/U1664/x[1] ), .d(\hdr_hld/high/U1664/U33/Z ), .e(
        \hdr_hld/high/U1664/x[0] ), .f(\hdr_hld/high/U1664/U33/Z ) );
    inv_1 \hdr_hld/high/U1664/U33/U30/Uinv  ( .x(\hdr_hld/high/U1664/U33/Z ), 
        .a(\hdr_hld/high/U1664/y[0] ) );
    aoi222_1 \hdr_hld/high/U1664/U30/U30/U1  ( .x(\hdr_hld/high/U1664/y[1] ), 
        .a(\hdr_hld/high/U1664/x[3] ), .b(\hdr_hld/high/U1664/x[2] ), .c(
        \hdr_hld/high/U1664/x[3] ), .d(\hdr_hld/high/U1664/U30/Z ), .e(
        \hdr_hld/high/U1664/x[2] ), .f(\hdr_hld/high/U1664/U30/Z ) );
    inv_1 \hdr_hld/high/U1664/U30/U30/Uinv  ( .x(\hdr_hld/high/U1664/U30/Z ), 
        .a(\hdr_hld/high/U1664/y[1] ) );
    aoi222_1 \hdr_hld/high/U1664/U31/U30/U1  ( .x(\hdr_hld/high/U1664/x[1] ), 
        .a(\hdr_hld/high/ncd[3] ), .b(\hdr_hld/high/ncd[2] ), .c(
        \hdr_hld/high/ncd[3] ), .d(\hdr_hld/high/U1664/U31/Z ), .e(
        \hdr_hld/high/ncd[2] ), .f(\hdr_hld/high/U1664/U31/Z ) );
    inv_1 \hdr_hld/high/U1664/U31/U30/Uinv  ( .x(\hdr_hld/high/U1664/U31/Z ), 
        .a(\hdr_hld/high/U1664/x[1] ) );
    aoi222_1 \hdr_hld/high/U1664/U37/U30/U1  ( .x(\hdr_hld/high/localcd ), .a(
        \hdr_hld/high/U1664/y[0] ), .b(\hdr_hld/high/U1664/y[1] ), .c(
        \hdr_hld/high/U1664/y[0] ), .d(\hdr_hld/high/U1664/U37/Z ), .e(
        \hdr_hld/high/U1664/y[1] ), .f(\hdr_hld/high/U1664/U37/Z ) );
    inv_1 \hdr_hld/high/U1664/U37/U30/Uinv  ( .x(\hdr_hld/high/U1664/U37/Z ), 
        .a(\hdr_hld/high/localcd ) );
    nor3_1 \hdr_hld/high/U1669/Unr  ( .x(\hdr_hld/high/U1669/nr ), .a(
        \hdr_hld/high/ctrlack_internal ), .b(\hdr_hld/high/drivel ), .c(n6) );
    nand3_1 \hdr_hld/high/U1669/Und  ( .x(\hdr_hld/high/U1669/nd ), .a(
        \hdr_hld/high/ctrlack_internal ), .b(\hdr_hld/high/drivel ), .c(n6) );
    oa21_1 \hdr_hld/high/U1669/U1  ( .x(\hdr_hld/high/U1669/n2 ), .a(
        \hdr_hld/high/U1669/n2 ), .b(\hdr_hld/high/U1669/nr ), .c(
        \hdr_hld/high/U1669/nd ) );
    inv_2 \hdr_hld/high/U1669/U3  ( .x(\hdr_hld/net20 ), .a(
        \hdr_hld/high/U1669/n2 ) );
    buf_2 U1 ( .x(n2), .a(\hdr_hld/net20 ) );
    buf_2 U2 ( .x(n1), .a(\hdr_hld/net20 ) );
    buf_1 U3 ( .x(n3), .a(\hdr_hld/low/latch ) );
    buf_1 U4 ( .x(n4), .a(\hdr_hld/high/drivel ) );
    buf_3 U5 ( .x(n5), .a(\hdr_hld/high/driveh ) );
    buf_3 U6 ( .x(n6), .a(\hdr_hld/high/driveh ) );
    buf_1 U7 ( .x(n7), .a(\hdr_hld/high/latch ) );
    inv_2 U8 ( .x(reset), .a(nReset) );
    buf_3 U9 ( .x(pullcd), .a(n9) );
endmodule


module chain_irdemux_32new_3 ( ctrlack, oh, ol, pullreq, pull_h, pull_l, 
    pullcd, reset, ctrlreq );
output [31:0] oh;
output [31:0] ol;
input  [7:0] pull_h;
input  [7:0] pull_l;
input  pullcd, reset, ctrlreq;
output ctrlack, pullreq;
    wire net30, net31, \I0/net32 , \I0/net33 , \I0/low/latch , 
        \I0/low/nlocalcd , \I0/low/localcd , \I0/low/ncd[0] , \I0/low/ncd[1] , 
        \I0/low/ncd[2] , \I0/low/ncd[3] , \I0/low/ncd[4] , \I0/low/ncd[5] , 
        \I0/low/ncd[6] , \I0/low/ncd[7] , \I0/low/ctrlack_internal , 
        \I0/low/acb , \I0/low/ba , \I0/low/driveh , \I0/net20 , 
        \I0/low/drivel , n1, n2, \I0/low/U4/U28/U1/clr , 
        \I0/low/U4/U28/U1/set , \I0/low/U1/Z , \I0/low/U1664/x[3] , 
        \I0/low/U1664/U28/Z , \I0/low/U1664/x[0] , \I0/low/U1664/U32/Z , 
        \I0/low/U1664/x[2] , \I0/low/U1664/U29/Z , \I0/low/U1664/y[0] , 
        \I0/low/U1664/x[1] , \I0/low/U1664/U33/Z , \I0/low/U1664/y[1] , 
        \I0/low/U1664/U30/Z , \I0/low/U1664/U31/Z , \I0/low/U1664/U37/Z , 
        \I0/low/U1669/nr , \I0/low/U1669/nd , \I0/low/U1669/n2 , 
        \I0/high/latch , \I0/high/nlocalcd , \I0/high/localcd , 
        \I0/high/ncd[0] , \I0/high/ncd[1] , \I0/high/ncd[2] , \I0/high/ncd[3] , 
        \I0/high/ncd[4] , \I0/high/ncd[5] , \I0/high/ncd[6] , \I0/high/ncd[7] , 
        \I0/high/ctrlack_internal , \I0/high/acb , \I0/high/ba , 
        \I0/high/driveh , net17, \I0/high/drivel , n3, n4, 
        \I0/high/U4/U28/U1/clr , \I0/high/U4/U28/U1/set , \I0/high/U1/Z , 
        \I0/high/U1664/x[3] , \I0/high/U1664/U28/Z , \I0/high/U1664/x[0] , 
        \I0/high/U1664/U32/Z , \I0/high/U1664/x[2] , \I0/high/U1664/U29/Z , 
        \I0/high/U1664/y[0] , \I0/high/U1664/x[1] , \I0/high/U1664/U33/Z , 
        \I0/high/U1664/y[1] , \I0/high/U1664/U30/Z , \I0/high/U1664/U31/Z , 
        \I0/high/U1664/U37/Z , \I0/high/U1669/nr , \I0/high/U1669/nd , 
        \I0/high/U1669/n2 , \I1/net32 , \I1/net33 , \I1/low/latch , 
        \I1/low/nlocalcd , \I1/low/localcd , \I1/low/ncd[0] , \I1/low/ncd[1] , 
        \I1/low/ncd[2] , \I1/low/ncd[3] , \I1/low/ncd[4] , \I1/low/ncd[5] , 
        \I1/low/ncd[6] , \I1/low/ncd[7] , \I1/low/ctrlack_internal , 
        \I1/low/acb , \I1/low/ba , \I1/low/driveh , \I1/net20 , 
        \I1/low/drivel , n5, n6, \I1/low/U4/U28/U1/clr , 
        \I1/low/U4/U28/U1/set , \I1/low/U1/Z , \I1/low/U1664/x[3] , 
        \I1/low/U1664/U28/Z , \I1/low/U1664/x[0] , \I1/low/U1664/U32/Z , 
        \I1/low/U1664/x[2] , \I1/low/U1664/U29/Z , \I1/low/U1664/y[0] , 
        \I1/low/U1664/x[1] , \I1/low/U1664/U33/Z , \I1/low/U1664/y[1] , 
        \I1/low/U1664/U30/Z , \I1/low/U1664/U31/Z , \I1/low/U1664/U37/Z , 
        \I1/low/U1669/nr , \I1/low/U1669/nd , \I1/low/U1669/n2 , 
        \I1/high/latch , \I1/high/nlocalcd , \I1/high/localcd , 
        \I1/high/ncd[0] , \I1/high/ncd[1] , \I1/high/ncd[2] , \I1/high/ncd[3] , 
        \I1/high/ncd[4] , \I1/high/ncd[5] , \I1/high/ncd[6] , \I1/high/ncd[7] , 
        \I1/high/ctrlack_internal , \I1/high/acb , \I1/high/ba , n7, n8, n12, 
        n10, n11, \I1/high/U4/U28/U1/clr , \I1/high/U4/U28/U1/set , 
        \I1/high/U1/Z , \I1/high/U1664/x[3] , \I1/high/U1664/U28/Z , 
        \I1/high/U1664/x[0] , \I1/high/U1664/U32/Z , \I1/high/U1664/x[2] , 
        \I1/high/U1664/U29/Z , \I1/high/U1664/y[0] , \I1/high/U1664/x[1] , 
        \I1/high/U1664/U33/Z , \I1/high/U1664/y[1] , \I1/high/U1664/U30/Z , 
        \I1/high/U1664/U31/Z , \I1/high/U1664/U37/Z , \I1/high/U1669/nr , 
        \I1/high/U1669/nd , \I1/high/U1669/n2 , n9;
    nand2_1 \U3/U5  ( .x(pullreq), .a(net30), .b(net31) );
    nor2_1 \I0/U3/U5  ( .x(net30), .a(\I0/net32 ), .b(\I0/net33 ) );
    buf_2 \I0/low/U1653  ( .x(\I0/low/latch ), .a(\I0/net32 ) );
    nor2_1 \I0/low/U264/U5  ( .x(\I0/low/nlocalcd ), .a(reset), .b(
        \I0/low/localcd ) );
    nor2_1 \I0/low/U1659_0_/U5  ( .x(\I0/low/ncd[0] ), .a(ol[0]), .b(oh[0]) );
    nor2_1 \I0/low/U1659_1_/U5  ( .x(\I0/low/ncd[1] ), .a(ol[1]), .b(oh[1]) );
    nor2_1 \I0/low/U1659_2_/U5  ( .x(\I0/low/ncd[2] ), .a(ol[2]), .b(oh[2]) );
    nor2_1 \I0/low/U1659_3_/U5  ( .x(\I0/low/ncd[3] ), .a(ol[3]), .b(oh[3]) );
    nor2_1 \I0/low/U1659_4_/U5  ( .x(\I0/low/ncd[4] ), .a(ol[4]), .b(oh[4]) );
    nor2_1 \I0/low/U1659_5_/U5  ( .x(\I0/low/ncd[5] ), .a(ol[5]), .b(oh[5]) );
    nor2_1 \I0/low/U1659_6_/U5  ( .x(\I0/low/ncd[6] ), .a(ol[6]), .b(oh[6]) );
    nor2_1 \I0/low/U1659_7_/U5  ( .x(\I0/low/ncd[7] ), .a(ol[7]), .b(oh[7]) );
    nor2_1 \I0/low/U3/U5  ( .x(\I0/low/ctrlack_internal ), .a(\I0/low/acb ), 
        .b(\I0/low/ba ) );
    buf_2 \I0/low/U1665/U7  ( .x(\I0/low/driveh ), .a(\I0/net20 ) );
    buf_2 \I0/low/U1666/U7  ( .x(\I0/low/drivel ), .a(\I0/net20 ) );
    ao23_1 \I0/low/U1658_0_/U21/U1/U1  ( .x(ol[0]), .a(\I0/low/driveh ), .b(ol
        [0]), .c(n1), .d(pull_l[0]), .e(n2) );
    ao23_1 \I0/low/U1658_1_/U21/U1/U1  ( .x(ol[1]), .a(\I0/low/drivel ), .b(ol
        [1]), .c(\I0/low/driveh ), .d(pull_l[1]), .e(n2) );
    ao23_1 \I0/low/U1658_2_/U21/U1/U1  ( .x(ol[2]), .a(\I0/low/drivel ), .b(ol
        [2]), .c(\I0/low/driveh ), .d(pull_l[2]), .e(n2) );
    ao23_1 \I0/low/U1658_3_/U21/U1/U1  ( .x(ol[3]), .a(\I0/low/driveh ), .b(ol
        [3]), .c(\I0/low/drivel ), .d(pull_l[3]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_4_/U21/U1/U1  ( .x(ol[4]), .a(n1), .b(ol[4]), .c(
        \I0/low/drivel ), .d(pull_l[4]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_5_/U21/U1/U1  ( .x(ol[5]), .a(\I0/low/driveh ), .b(ol
        [5]), .c(n1), .d(pull_l[5]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_6_/U21/U1/U1  ( .x(ol[6]), .a(\I0/low/drivel ), .b(ol
        [6]), .c(\I0/low/driveh ), .d(pull_l[6]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_7_/U21/U1/U1  ( .x(ol[7]), .a(n1), .b(ol[7]), .c(n1), 
        .d(pull_l[7]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_0_/U21/U1/U1  ( .x(oh[0]), .a(\I0/low/driveh ), .b(oh
        [0]), .c(n1), .d(pull_h[0]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_1_/U21/U1/U1  ( .x(oh[1]), .a(n1), .b(oh[1]), .c(
        \I0/low/drivel ), .d(pull_h[1]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_2_/U21/U1/U1  ( .x(oh[2]), .a(\I0/low/drivel ), .b(oh
        [2]), .c(\I0/low/drivel ), .d(pull_h[2]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_3_/U21/U1/U1  ( .x(oh[3]), .a(n1), .b(oh[3]), .c(
        \I0/low/driveh ), .d(pull_h[3]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_4_/U21/U1/U1  ( .x(oh[4]), .a(n1), .b(oh[4]), .c(n1), 
        .d(pull_h[4]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_5_/U21/U1/U1  ( .x(oh[5]), .a(\I0/low/drivel ), .b(oh
        [5]), .c(n1), .d(pull_h[5]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_6_/U21/U1/U1  ( .x(oh[6]), .a(\I0/low/drivel ), .b(oh
        [6]), .c(\I0/low/driveh ), .d(pull_h[6]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_7_/U21/U1/U1  ( .x(oh[7]), .a(\I0/low/driveh ), .b(oh
        [7]), .c(\I0/low/drivel ), .d(pull_h[7]), .e(\I0/low/latch ) );
    aoai211_1 \I0/low/U4/U28/U1/U1  ( .x(\I0/low/U4/U28/U1/clr ), .a(
        \I0/net20 ), .b(\I0/low/acb ), .c(\I0/low/nlocalcd ), .d(\I0/net32 )
         );
    nand3_1 \I0/low/U4/U28/U1/U2  ( .x(\I0/low/U4/U28/U1/set ), .a(
        \I0/low/nlocalcd ), .b(\I0/net20 ), .c(\I0/low/acb ) );
    nand2_2 \I0/low/U4/U28/U1/U3  ( .x(\I0/net32 ), .a(\I0/low/U4/U28/U1/clr ), 
        .b(\I0/low/U4/U28/U1/set ) );
    oai21_1 \I0/low/U1/U30/U1/U1  ( .x(\I0/low/acb ), .a(\I0/low/U1/Z ), .b(
        \I0/low/ba ), .c(\I0/net20 ) );
    inv_1 \I0/low/U1/U30/U1/U2  ( .x(\I0/low/U1/Z ), .a(\I0/low/acb ) );
    ao222_1 \I0/low/U5/U18/U1/U1  ( .x(\I0/low/ba ), .a(\I0/low/latch ), .b(
        pullcd), .c(\I0/low/latch ), .d(\I0/low/ba ), .e(pullcd), .f(
        \I0/low/ba ) );
    aoi222_1 \I0/low/U1664/U28/U30/U1  ( .x(\I0/low/U1664/x[3] ), .a(
        \I0/low/ncd[7] ), .b(\I0/low/ncd[6] ), .c(\I0/low/ncd[7] ), .d(
        \I0/low/U1664/U28/Z ), .e(\I0/low/ncd[6] ), .f(\I0/low/U1664/U28/Z )
         );
    inv_1 \I0/low/U1664/U28/U30/Uinv  ( .x(\I0/low/U1664/U28/Z ), .a(
        \I0/low/U1664/x[3] ) );
    aoi222_1 \I0/low/U1664/U32/U30/U1  ( .x(\I0/low/U1664/x[0] ), .a(
        \I0/low/ncd[1] ), .b(\I0/low/ncd[0] ), .c(\I0/low/ncd[1] ), .d(
        \I0/low/U1664/U32/Z ), .e(\I0/low/ncd[0] ), .f(\I0/low/U1664/U32/Z )
         );
    inv_1 \I0/low/U1664/U32/U30/Uinv  ( .x(\I0/low/U1664/U32/Z ), .a(
        \I0/low/U1664/x[0] ) );
    aoi222_1 \I0/low/U1664/U29/U30/U1  ( .x(\I0/low/U1664/x[2] ), .a(
        \I0/low/ncd[5] ), .b(\I0/low/ncd[4] ), .c(\I0/low/ncd[5] ), .d(
        \I0/low/U1664/U29/Z ), .e(\I0/low/ncd[4] ), .f(\I0/low/U1664/U29/Z )
         );
    inv_1 \I0/low/U1664/U29/U30/Uinv  ( .x(\I0/low/U1664/U29/Z ), .a(
        \I0/low/U1664/x[2] ) );
    aoi222_1 \I0/low/U1664/U33/U30/U1  ( .x(\I0/low/U1664/y[0] ), .a(
        \I0/low/U1664/x[1] ), .b(\I0/low/U1664/x[0] ), .c(\I0/low/U1664/x[1] ), 
        .d(\I0/low/U1664/U33/Z ), .e(\I0/low/U1664/x[0] ), .f(
        \I0/low/U1664/U33/Z ) );
    inv_1 \I0/low/U1664/U33/U30/Uinv  ( .x(\I0/low/U1664/U33/Z ), .a(
        \I0/low/U1664/y[0] ) );
    aoi222_1 \I0/low/U1664/U30/U30/U1  ( .x(\I0/low/U1664/y[1] ), .a(
        \I0/low/U1664/x[3] ), .b(\I0/low/U1664/x[2] ), .c(\I0/low/U1664/x[3] ), 
        .d(\I0/low/U1664/U30/Z ), .e(\I0/low/U1664/x[2] ), .f(
        \I0/low/U1664/U30/Z ) );
    inv_1 \I0/low/U1664/U30/U30/Uinv  ( .x(\I0/low/U1664/U30/Z ), .a(
        \I0/low/U1664/y[1] ) );
    aoi222_1 \I0/low/U1664/U31/U30/U1  ( .x(\I0/low/U1664/x[1] ), .a(
        \I0/low/ncd[3] ), .b(\I0/low/ncd[2] ), .c(\I0/low/ncd[3] ), .d(
        \I0/low/U1664/U31/Z ), .e(\I0/low/ncd[2] ), .f(\I0/low/U1664/U31/Z )
         );
    inv_1 \I0/low/U1664/U31/U30/Uinv  ( .x(\I0/low/U1664/U31/Z ), .a(
        \I0/low/U1664/x[1] ) );
    aoi222_1 \I0/low/U1664/U37/U30/U1  ( .x(\I0/low/localcd ), .a(
        \I0/low/U1664/y[0] ), .b(\I0/low/U1664/y[1] ), .c(\I0/low/U1664/y[0] ), 
        .d(\I0/low/U1664/U37/Z ), .e(\I0/low/U1664/y[1] ), .f(
        \I0/low/U1664/U37/Z ) );
    inv_1 \I0/low/U1664/U37/U30/Uinv  ( .x(\I0/low/U1664/U37/Z ), .a(
        \I0/low/localcd ) );
    nor3_1 \I0/low/U1669/Unr  ( .x(\I0/low/U1669/nr ), .a(
        \I0/low/ctrlack_internal ), .b(n1), .c(\I0/low/driveh ) );
    nand3_1 \I0/low/U1669/Und  ( .x(\I0/low/U1669/nd ), .a(
        \I0/low/ctrlack_internal ), .b(\I0/low/drivel ), .c(\I0/low/driveh )
         );
    oa21_1 \I0/low/U1669/U1  ( .x(\I0/low/U1669/n2 ), .a(\I0/low/U1669/n2 ), 
        .b(\I0/low/U1669/nr ), .c(\I0/low/U1669/nd ) );
    inv_2 \I0/low/U1669/U3  ( .x(ctrlack), .a(\I0/low/U1669/n2 ) );
    buf_2 \I0/high/U1653  ( .x(\I0/high/latch ), .a(\I0/net33 ) );
    nor2_1 \I0/high/U264/U5  ( .x(\I0/high/nlocalcd ), .a(reset), .b(
        \I0/high/localcd ) );
    nor2_1 \I0/high/U1659_0_/U5  ( .x(\I0/high/ncd[0] ), .a(ol[8]), .b(oh[8])
         );
    nor2_1 \I0/high/U1659_1_/U5  ( .x(\I0/high/ncd[1] ), .a(ol[9]), .b(oh[9])
         );
    nor2_1 \I0/high/U1659_2_/U5  ( .x(\I0/high/ncd[2] ), .a(ol[10]), .b(oh[10]
        ) );
    nor2_1 \I0/high/U1659_3_/U5  ( .x(\I0/high/ncd[3] ), .a(ol[11]), .b(oh[11]
        ) );
    nor2_1 \I0/high/U1659_4_/U5  ( .x(\I0/high/ncd[4] ), .a(ol[12]), .b(oh[12]
        ) );
    nor2_1 \I0/high/U1659_5_/U5  ( .x(\I0/high/ncd[5] ), .a(ol[13]), .b(oh[13]
        ) );
    nor2_1 \I0/high/U1659_6_/U5  ( .x(\I0/high/ncd[6] ), .a(ol[14]), .b(oh[14]
        ) );
    nor2_1 \I0/high/U1659_7_/U5  ( .x(\I0/high/ncd[7] ), .a(ol[15]), .b(oh[15]
        ) );
    nor2_1 \I0/high/U3/U5  ( .x(\I0/high/ctrlack_internal ), .a(\I0/high/acb ), 
        .b(\I0/high/ba ) );
    buf_2 \I0/high/U1665/U7  ( .x(\I0/high/driveh ), .a(net17) );
    buf_2 \I0/high/U1666/U7  ( .x(\I0/high/drivel ), .a(net17) );
    ao23_1 \I0/high/U1658_0_/U21/U1/U1  ( .x(ol[8]), .a(\I0/high/driveh ), .b(
        ol[8]), .c(n3), .d(pull_l[0]), .e(n4) );
    ao23_1 \I0/high/U1658_1_/U21/U1/U1  ( .x(ol[9]), .a(\I0/high/drivel ), .b(
        ol[9]), .c(\I0/high/driveh ), .d(pull_l[1]), .e(n4) );
    ao23_1 \I0/high/U1658_2_/U21/U1/U1  ( .x(ol[10]), .a(\I0/high/drivel ), 
        .b(ol[10]), .c(\I0/high/driveh ), .d(pull_l[2]), .e(n4) );
    ao23_1 \I0/high/U1658_3_/U21/U1/U1  ( .x(ol[11]), .a(\I0/high/driveh ), 
        .b(ol[11]), .c(\I0/high/drivel ), .d(pull_l[3]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1658_4_/U21/U1/U1  ( .x(ol[12]), .a(n3), .b(ol[12]), .c(
        \I0/high/drivel ), .d(pull_l[4]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1658_5_/U21/U1/U1  ( .x(ol[13]), .a(\I0/high/driveh ), 
        .b(ol[13]), .c(n3), .d(pull_l[5]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1658_6_/U21/U1/U1  ( .x(ol[14]), .a(\I0/high/drivel ), 
        .b(ol[14]), .c(\I0/high/driveh ), .d(pull_l[6]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1658_7_/U21/U1/U1  ( .x(ol[15]), .a(n3), .b(ol[15]), .c(
        n3), .d(pull_l[7]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_0_/U21/U1/U1  ( .x(oh[8]), .a(\I0/high/driveh ), .b(
        oh[8]), .c(n3), .d(pull_h[0]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_1_/U21/U1/U1  ( .x(oh[9]), .a(n3), .b(oh[9]), .c(
        \I0/high/drivel ), .d(pull_h[1]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_2_/U21/U1/U1  ( .x(oh[10]), .a(\I0/high/drivel ), 
        .b(oh[10]), .c(\I0/high/drivel ), .d(pull_h[2]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1651_3_/U21/U1/U1  ( .x(oh[11]), .a(n3), .b(oh[11]), .c(
        \I0/high/driveh ), .d(pull_h[3]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_4_/U21/U1/U1  ( .x(oh[12]), .a(n3), .b(oh[12]), .c(
        n3), .d(pull_h[4]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_5_/U21/U1/U1  ( .x(oh[13]), .a(\I0/high/drivel ), 
        .b(oh[13]), .c(n3), .d(pull_h[5]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_6_/U21/U1/U1  ( .x(oh[14]), .a(\I0/high/drivel ), 
        .b(oh[14]), .c(\I0/high/driveh ), .d(pull_h[6]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1651_7_/U21/U1/U1  ( .x(oh[15]), .a(\I0/high/driveh ), 
        .b(oh[15]), .c(\I0/high/drivel ), .d(pull_h[7]), .e(\I0/high/latch )
         );
    aoai211_1 \I0/high/U4/U28/U1/U1  ( .x(\I0/high/U4/U28/U1/clr ), .a(net17), 
        .b(\I0/high/acb ), .c(\I0/high/nlocalcd ), .d(\I0/net33 ) );
    nand3_1 \I0/high/U4/U28/U1/U2  ( .x(\I0/high/U4/U28/U1/set ), .a(
        \I0/high/nlocalcd ), .b(net17), .c(\I0/high/acb ) );
    nand2_2 \I0/high/U4/U28/U1/U3  ( .x(\I0/net33 ), .a(
        \I0/high/U4/U28/U1/clr ), .b(\I0/high/U4/U28/U1/set ) );
    oai21_1 \I0/high/U1/U30/U1/U1  ( .x(\I0/high/acb ), .a(\I0/high/U1/Z ), 
        .b(\I0/high/ba ), .c(net17) );
    inv_1 \I0/high/U1/U30/U1/U2  ( .x(\I0/high/U1/Z ), .a(\I0/high/acb ) );
    ao222_1 \I0/high/U5/U18/U1/U1  ( .x(\I0/high/ba ), .a(\I0/high/latch ), 
        .b(pullcd), .c(\I0/high/latch ), .d(\I0/high/ba ), .e(pullcd), .f(
        \I0/high/ba ) );
    aoi222_1 \I0/high/U1664/U28/U30/U1  ( .x(\I0/high/U1664/x[3] ), .a(
        \I0/high/ncd[7] ), .b(\I0/high/ncd[6] ), .c(\I0/high/ncd[7] ), .d(
        \I0/high/U1664/U28/Z ), .e(\I0/high/ncd[6] ), .f(\I0/high/U1664/U28/Z 
        ) );
    inv_1 \I0/high/U1664/U28/U30/Uinv  ( .x(\I0/high/U1664/U28/Z ), .a(
        \I0/high/U1664/x[3] ) );
    aoi222_1 \I0/high/U1664/U32/U30/U1  ( .x(\I0/high/U1664/x[0] ), .a(
        \I0/high/ncd[1] ), .b(\I0/high/ncd[0] ), .c(\I0/high/ncd[1] ), .d(
        \I0/high/U1664/U32/Z ), .e(\I0/high/ncd[0] ), .f(\I0/high/U1664/U32/Z 
        ) );
    inv_1 \I0/high/U1664/U32/U30/Uinv  ( .x(\I0/high/U1664/U32/Z ), .a(
        \I0/high/U1664/x[0] ) );
    aoi222_1 \I0/high/U1664/U29/U30/U1  ( .x(\I0/high/U1664/x[2] ), .a(
        \I0/high/ncd[5] ), .b(\I0/high/ncd[4] ), .c(\I0/high/ncd[5] ), .d(
        \I0/high/U1664/U29/Z ), .e(\I0/high/ncd[4] ), .f(\I0/high/U1664/U29/Z 
        ) );
    inv_1 \I0/high/U1664/U29/U30/Uinv  ( .x(\I0/high/U1664/U29/Z ), .a(
        \I0/high/U1664/x[2] ) );
    aoi222_1 \I0/high/U1664/U33/U30/U1  ( .x(\I0/high/U1664/y[0] ), .a(
        \I0/high/U1664/x[1] ), .b(\I0/high/U1664/x[0] ), .c(
        \I0/high/U1664/x[1] ), .d(\I0/high/U1664/U33/Z ), .e(
        \I0/high/U1664/x[0] ), .f(\I0/high/U1664/U33/Z ) );
    inv_1 \I0/high/U1664/U33/U30/Uinv  ( .x(\I0/high/U1664/U33/Z ), .a(
        \I0/high/U1664/y[0] ) );
    aoi222_1 \I0/high/U1664/U30/U30/U1  ( .x(\I0/high/U1664/y[1] ), .a(
        \I0/high/U1664/x[3] ), .b(\I0/high/U1664/x[2] ), .c(
        \I0/high/U1664/x[3] ), .d(\I0/high/U1664/U30/Z ), .e(
        \I0/high/U1664/x[2] ), .f(\I0/high/U1664/U30/Z ) );
    inv_1 \I0/high/U1664/U30/U30/Uinv  ( .x(\I0/high/U1664/U30/Z ), .a(
        \I0/high/U1664/y[1] ) );
    aoi222_1 \I0/high/U1664/U31/U30/U1  ( .x(\I0/high/U1664/x[1] ), .a(
        \I0/high/ncd[3] ), .b(\I0/high/ncd[2] ), .c(\I0/high/ncd[3] ), .d(
        \I0/high/U1664/U31/Z ), .e(\I0/high/ncd[2] ), .f(\I0/high/U1664/U31/Z 
        ) );
    inv_1 \I0/high/U1664/U31/U30/Uinv  ( .x(\I0/high/U1664/U31/Z ), .a(
        \I0/high/U1664/x[1] ) );
    aoi222_1 \I0/high/U1664/U37/U30/U1  ( .x(\I0/high/localcd ), .a(
        \I0/high/U1664/y[0] ), .b(\I0/high/U1664/y[1] ), .c(
        \I0/high/U1664/y[0] ), .d(\I0/high/U1664/U37/Z ), .e(
        \I0/high/U1664/y[1] ), .f(\I0/high/U1664/U37/Z ) );
    inv_1 \I0/high/U1664/U37/U30/Uinv  ( .x(\I0/high/U1664/U37/Z ), .a(
        \I0/high/localcd ) );
    nor3_1 \I0/high/U1669/Unr  ( .x(\I0/high/U1669/nr ), .a(
        \I0/high/ctrlack_internal ), .b(n3), .c(\I0/high/driveh ) );
    nand3_1 \I0/high/U1669/Und  ( .x(\I0/high/U1669/nd ), .a(
        \I0/high/ctrlack_internal ), .b(\I0/high/drivel ), .c(\I0/high/driveh 
        ) );
    oa21_1 \I0/high/U1669/U1  ( .x(\I0/high/U1669/n2 ), .a(\I0/high/U1669/n2 ), 
        .b(\I0/high/U1669/nr ), .c(\I0/high/U1669/nd ) );
    inv_2 \I0/high/U1669/U3  ( .x(\I0/net20 ), .a(\I0/high/U1669/n2 ) );
    nor2_1 \I1/U3/U5  ( .x(net31), .a(\I1/net32 ), .b(\I1/net33 ) );
    buf_2 \I1/low/U1653  ( .x(\I1/low/latch ), .a(\I1/net32 ) );
    nor2_1 \I1/low/U264/U5  ( .x(\I1/low/nlocalcd ), .a(reset), .b(
        \I1/low/localcd ) );
    nor2_1 \I1/low/U1659_0_/U5  ( .x(\I1/low/ncd[0] ), .a(ol[16]), .b(oh[16])
         );
    nor2_1 \I1/low/U1659_1_/U5  ( .x(\I1/low/ncd[1] ), .a(ol[17]), .b(oh[17])
         );
    nor2_1 \I1/low/U1659_2_/U5  ( .x(\I1/low/ncd[2] ), .a(ol[18]), .b(oh[18])
         );
    nor2_1 \I1/low/U1659_3_/U5  ( .x(\I1/low/ncd[3] ), .a(ol[19]), .b(oh[19])
         );
    nor2_1 \I1/low/U1659_4_/U5  ( .x(\I1/low/ncd[4] ), .a(ol[20]), .b(oh[20])
         );
    nor2_1 \I1/low/U1659_5_/U5  ( .x(\I1/low/ncd[5] ), .a(ol[21]), .b(oh[21])
         );
    nor2_1 \I1/low/U1659_6_/U5  ( .x(\I1/low/ncd[6] ), .a(ol[22]), .b(oh[22])
         );
    nor2_1 \I1/low/U1659_7_/U5  ( .x(\I1/low/ncd[7] ), .a(ol[23]), .b(oh[23])
         );
    nor2_1 \I1/low/U3/U5  ( .x(\I1/low/ctrlack_internal ), .a(\I1/low/acb ), 
        .b(\I1/low/ba ) );
    buf_2 \I1/low/U1665/U7  ( .x(\I1/low/driveh ), .a(\I1/net20 ) );
    buf_2 \I1/low/U1666/U7  ( .x(\I1/low/drivel ), .a(\I1/net20 ) );
    ao23_1 \I1/low/U1658_0_/U21/U1/U1  ( .x(ol[16]), .a(\I1/low/drivel ), .b(
        ol[16]), .c(n5), .d(pull_l[0]), .e(n6) );
    ao23_1 \I1/low/U1658_1_/U21/U1/U1  ( .x(ol[17]), .a(\I1/low/driveh ), .b(
        ol[17]), .c(n5), .d(pull_l[1]), .e(n6) );
    ao23_1 \I1/low/U1658_2_/U21/U1/U1  ( .x(ol[18]), .a(\I1/low/drivel ), .b(
        ol[18]), .c(\I1/low/driveh ), .d(pull_l[2]), .e(n6) );
    ao23_1 \I1/low/U1658_3_/U21/U1/U1  ( .x(ol[19]), .a(n5), .b(ol[19]), .c(
        \I1/low/driveh ), .d(pull_l[3]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_4_/U21/U1/U1  ( .x(ol[20]), .a(\I1/low/driveh ), .b(
        ol[20]), .c(\I1/low/drivel ), .d(pull_l[4]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_5_/U21/U1/U1  ( .x(ol[21]), .a(n5), .b(ol[21]), .c(
        \I1/low/drivel ), .d(pull_l[5]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_6_/U21/U1/U1  ( .x(ol[22]), .a(\I1/low/driveh ), .b(
        ol[22]), .c(n5), .d(pull_l[6]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_7_/U21/U1/U1  ( .x(ol[23]), .a(\I1/low/drivel ), .b(
        ol[23]), .c(\I1/low/driveh ), .d(pull_l[7]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_0_/U21/U1/U1  ( .x(oh[16]), .a(\I1/low/driveh ), .b(
        oh[16]), .c(\I1/low/drivel ), .d(pull_h[0]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_1_/U21/U1/U1  ( .x(oh[17]), .a(\I1/low/drivel ), .b(
        oh[17]), .c(n5), .d(pull_h[1]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_2_/U21/U1/U1  ( .x(oh[18]), .a(\I1/low/drivel ), .b(
        oh[18]), .c(\I1/low/driveh ), .d(pull_h[2]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_3_/U21/U1/U1  ( .x(oh[19]), .a(n5), .b(oh[19]), .c(n5
        ), .d(pull_h[3]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_4_/U21/U1/U1  ( .x(oh[20]), .a(n5), .b(oh[20]), .c(n5
        ), .d(pull_h[4]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_5_/U21/U1/U1  ( .x(oh[21]), .a(\I1/low/drivel ), .b(
        oh[21]), .c(\I1/low/driveh ), .d(pull_h[5]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_6_/U21/U1/U1  ( .x(oh[22]), .a(n5), .b(oh[22]), .c(
        \I1/low/drivel ), .d(pull_h[6]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_7_/U21/U1/U1  ( .x(oh[23]), .a(\I1/low/driveh ), .b(
        oh[23]), .c(\I1/low/drivel ), .d(pull_h[7]), .e(\I1/low/latch ) );
    aoai211_1 \I1/low/U4/U28/U1/U1  ( .x(\I1/low/U4/U28/U1/clr ), .a(
        \I1/net20 ), .b(\I1/low/acb ), .c(\I1/low/nlocalcd ), .d(\I1/net32 )
         );
    nand3_1 \I1/low/U4/U28/U1/U2  ( .x(\I1/low/U4/U28/U1/set ), .a(
        \I1/low/nlocalcd ), .b(\I1/net20 ), .c(\I1/low/acb ) );
    nand2_2 \I1/low/U4/U28/U1/U3  ( .x(\I1/net32 ), .a(\I1/low/U4/U28/U1/clr ), 
        .b(\I1/low/U4/U28/U1/set ) );
    oai21_1 \I1/low/U1/U30/U1/U1  ( .x(\I1/low/acb ), .a(\I1/low/U1/Z ), .b(
        \I1/low/ba ), .c(\I1/net20 ) );
    inv_1 \I1/low/U1/U30/U1/U2  ( .x(\I1/low/U1/Z ), .a(\I1/low/acb ) );
    ao222_1 \I1/low/U5/U18/U1/U1  ( .x(\I1/low/ba ), .a(\I1/low/latch ), .b(
        pullcd), .c(\I1/low/latch ), .d(\I1/low/ba ), .e(pullcd), .f(
        \I1/low/ba ) );
    aoi222_1 \I1/low/U1664/U28/U30/U1  ( .x(\I1/low/U1664/x[3] ), .a(
        \I1/low/ncd[7] ), .b(\I1/low/ncd[6] ), .c(\I1/low/ncd[7] ), .d(
        \I1/low/U1664/U28/Z ), .e(\I1/low/ncd[6] ), .f(\I1/low/U1664/U28/Z )
         );
    inv_1 \I1/low/U1664/U28/U30/Uinv  ( .x(\I1/low/U1664/U28/Z ), .a(
        \I1/low/U1664/x[3] ) );
    aoi222_1 \I1/low/U1664/U32/U30/U1  ( .x(\I1/low/U1664/x[0] ), .a(
        \I1/low/ncd[1] ), .b(\I1/low/ncd[0] ), .c(\I1/low/ncd[1] ), .d(
        \I1/low/U1664/U32/Z ), .e(\I1/low/ncd[0] ), .f(\I1/low/U1664/U32/Z )
         );
    inv_1 \I1/low/U1664/U32/U30/Uinv  ( .x(\I1/low/U1664/U32/Z ), .a(
        \I1/low/U1664/x[0] ) );
    aoi222_1 \I1/low/U1664/U29/U30/U1  ( .x(\I1/low/U1664/x[2] ), .a(
        \I1/low/ncd[5] ), .b(\I1/low/ncd[4] ), .c(\I1/low/ncd[5] ), .d(
        \I1/low/U1664/U29/Z ), .e(\I1/low/ncd[4] ), .f(\I1/low/U1664/U29/Z )
         );
    inv_1 \I1/low/U1664/U29/U30/Uinv  ( .x(\I1/low/U1664/U29/Z ), .a(
        \I1/low/U1664/x[2] ) );
    aoi222_1 \I1/low/U1664/U33/U30/U1  ( .x(\I1/low/U1664/y[0] ), .a(
        \I1/low/U1664/x[1] ), .b(\I1/low/U1664/x[0] ), .c(\I1/low/U1664/x[1] ), 
        .d(\I1/low/U1664/U33/Z ), .e(\I1/low/U1664/x[0] ), .f(
        \I1/low/U1664/U33/Z ) );
    inv_1 \I1/low/U1664/U33/U30/Uinv  ( .x(\I1/low/U1664/U33/Z ), .a(
        \I1/low/U1664/y[0] ) );
    aoi222_1 \I1/low/U1664/U30/U30/U1  ( .x(\I1/low/U1664/y[1] ), .a(
        \I1/low/U1664/x[3] ), .b(\I1/low/U1664/x[2] ), .c(\I1/low/U1664/x[3] ), 
        .d(\I1/low/U1664/U30/Z ), .e(\I1/low/U1664/x[2] ), .f(
        \I1/low/U1664/U30/Z ) );
    inv_1 \I1/low/U1664/U30/U30/Uinv  ( .x(\I1/low/U1664/U30/Z ), .a(
        \I1/low/U1664/y[1] ) );
    aoi222_1 \I1/low/U1664/U31/U30/U1  ( .x(\I1/low/U1664/x[1] ), .a(
        \I1/low/ncd[3] ), .b(\I1/low/ncd[2] ), .c(\I1/low/ncd[3] ), .d(
        \I1/low/U1664/U31/Z ), .e(\I1/low/ncd[2] ), .f(\I1/low/U1664/U31/Z )
         );
    inv_1 \I1/low/U1664/U31/U30/Uinv  ( .x(\I1/low/U1664/U31/Z ), .a(
        \I1/low/U1664/x[1] ) );
    aoi222_1 \I1/low/U1664/U37/U30/U1  ( .x(\I1/low/localcd ), .a(
        \I1/low/U1664/y[0] ), .b(\I1/low/U1664/y[1] ), .c(\I1/low/U1664/y[0] ), 
        .d(\I1/low/U1664/U37/Z ), .e(\I1/low/U1664/y[1] ), .f(
        \I1/low/U1664/U37/Z ) );
    inv_1 \I1/low/U1664/U37/U30/Uinv  ( .x(\I1/low/U1664/U37/Z ), .a(
        \I1/low/localcd ) );
    nor3_1 \I1/low/U1669/Unr  ( .x(\I1/low/U1669/nr ), .a(
        \I1/low/ctrlack_internal ), .b(n5), .c(\I1/low/driveh ) );
    nand3_1 \I1/low/U1669/Und  ( .x(\I1/low/U1669/nd ), .a(
        \I1/low/ctrlack_internal ), .b(\I1/low/drivel ), .c(\I1/low/driveh )
         );
    oa21_1 \I1/low/U1669/U1  ( .x(\I1/low/U1669/n2 ), .a(\I1/low/U1669/n2 ), 
        .b(\I1/low/U1669/nr ), .c(\I1/low/U1669/nd ) );
    inv_2 \I1/low/U1669/U3  ( .x(net17), .a(\I1/low/U1669/n2 ) );
    buf_2 \I1/high/U1653  ( .x(\I1/high/latch ), .a(\I1/net33 ) );
    nor2_1 \I1/high/U264/U5  ( .x(\I1/high/nlocalcd ), .a(reset), .b(
        \I1/high/localcd ) );
    nor2_1 \I1/high/U1659_0_/U5  ( .x(\I1/high/ncd[0] ), .a(ol[24]), .b(oh[24]
        ) );
    nor2_1 \I1/high/U1659_1_/U5  ( .x(\I1/high/ncd[1] ), .a(ol[25]), .b(oh[25]
        ) );
    nor2_1 \I1/high/U1659_2_/U5  ( .x(\I1/high/ncd[2] ), .a(ol[26]), .b(oh[26]
        ) );
    nor2_1 \I1/high/U1659_3_/U5  ( .x(\I1/high/ncd[3] ), .a(ol[27]), .b(oh[27]
        ) );
    nor2_1 \I1/high/U1659_4_/U5  ( .x(\I1/high/ncd[4] ), .a(ol[28]), .b(oh[28]
        ) );
    nor2_1 \I1/high/U1659_5_/U5  ( .x(\I1/high/ncd[5] ), .a(ol[29]), .b(oh[29]
        ) );
    nor2_1 \I1/high/U1659_6_/U5  ( .x(\I1/high/ncd[6] ), .a(ol[30]), .b(oh[30]
        ) );
    nor2_1 \I1/high/U1659_7_/U5  ( .x(\I1/high/ncd[7] ), .a(ol[31]), .b(oh[31]
        ) );
    nor2_1 \I1/high/U3/U5  ( .x(\I1/high/ctrlack_internal ), .a(\I1/high/acb ), 
        .b(\I1/high/ba ) );
    ao23_1 \I1/high/U1658_0_/U21/U1/U1  ( .x(ol[24]), .a(n7), .b(ol[24]), .c(
        n8), .d(pull_l[0]), .e(n12) );
    ao23_1 \I1/high/U1658_1_/U21/U1/U1  ( .x(ol[25]), .a(n7), .b(ol[25]), .c(
        n8), .d(pull_l[1]), .e(n12) );
    ao23_1 \I1/high/U1658_2_/U21/U1/U1  ( .x(ol[26]), .a(n7), .b(ol[26]), .c(
        n7), .d(pull_l[2]), .e(n12) );
    ao23_1 \I1/high/U1658_3_/U21/U1/U1  ( .x(ol[27]), .a(n7), .b(ol[27]), .c(
        n7), .d(pull_l[3]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1658_4_/U21/U1/U1  ( .x(ol[28]), .a(n7), .b(ol[28]), .c(
        n7), .d(pull_l[4]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1658_5_/U21/U1/U1  ( .x(ol[29]), .a(n7), .b(ol[29]), .c(
        n8), .d(pull_l[5]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1658_6_/U21/U1/U1  ( .x(ol[30]), .a(n7), .b(ol[30]), .c(
        n8), .d(pull_l[6]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1658_7_/U21/U1/U1  ( .x(ol[31]), .a(n7), .b(ol[31]), .c(
        n8), .d(pull_l[7]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_0_/U21/U1/U1  ( .x(oh[24]), .a(n10), .b(oh[24]), .c(
        n10), .d(pull_h[0]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_1_/U21/U1/U1  ( .x(oh[25]), .a(n10), .b(oh[25]), .c(
        n11), .d(pull_h[1]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_2_/U21/U1/U1  ( .x(oh[26]), .a(n10), .b(oh[26]), .c(
        n11), .d(pull_h[2]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_3_/U21/U1/U1  ( .x(oh[27]), .a(n10), .b(oh[27]), .c(
        n10), .d(pull_h[3]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_4_/U21/U1/U1  ( .x(oh[28]), .a(n10), .b(oh[28]), .c(
        n11), .d(pull_h[4]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_5_/U21/U1/U1  ( .x(oh[29]), .a(n10), .b(oh[29]), .c(
        n11), .d(pull_h[5]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_6_/U21/U1/U1  ( .x(oh[30]), .a(n10), .b(oh[30]), .c(
        n11), .d(pull_h[6]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_7_/U21/U1/U1  ( .x(oh[31]), .a(n10), .b(oh[31]), .c(
        n10), .d(pull_h[7]), .e(\I1/high/latch ) );
    aoai211_1 \I1/high/U4/U28/U1/U1  ( .x(\I1/high/U4/U28/U1/clr ), .a(ctrlreq
        ), .b(\I1/high/acb ), .c(\I1/high/nlocalcd ), .d(\I1/net33 ) );
    nand3_1 \I1/high/U4/U28/U1/U2  ( .x(\I1/high/U4/U28/U1/set ), .a(
        \I1/high/nlocalcd ), .b(ctrlreq), .c(\I1/high/acb ) );
    nand2_2 \I1/high/U4/U28/U1/U3  ( .x(\I1/net33 ), .a(
        \I1/high/U4/U28/U1/clr ), .b(\I1/high/U4/U28/U1/set ) );
    oai21_1 \I1/high/U1/U30/U1/U1  ( .x(\I1/high/acb ), .a(\I1/high/U1/Z ), 
        .b(\I1/high/ba ), .c(ctrlreq) );
    inv_1 \I1/high/U1/U30/U1/U2  ( .x(\I1/high/U1/Z ), .a(\I1/high/acb ) );
    ao222_1 \I1/high/U5/U18/U1/U1  ( .x(\I1/high/ba ), .a(\I1/high/latch ), 
        .b(pullcd), .c(\I1/high/latch ), .d(\I1/high/ba ), .e(pullcd), .f(
        \I1/high/ba ) );
    aoi222_1 \I1/high/U1664/U28/U30/U1  ( .x(\I1/high/U1664/x[3] ), .a(
        \I1/high/ncd[7] ), .b(\I1/high/ncd[6] ), .c(\I1/high/ncd[7] ), .d(
        \I1/high/U1664/U28/Z ), .e(\I1/high/ncd[6] ), .f(\I1/high/U1664/U28/Z 
        ) );
    inv_1 \I1/high/U1664/U28/U30/Uinv  ( .x(\I1/high/U1664/U28/Z ), .a(
        \I1/high/U1664/x[3] ) );
    aoi222_1 \I1/high/U1664/U32/U30/U1  ( .x(\I1/high/U1664/x[0] ), .a(
        \I1/high/ncd[1] ), .b(\I1/high/ncd[0] ), .c(\I1/high/ncd[1] ), .d(
        \I1/high/U1664/U32/Z ), .e(\I1/high/ncd[0] ), .f(\I1/high/U1664/U32/Z 
        ) );
    inv_1 \I1/high/U1664/U32/U30/Uinv  ( .x(\I1/high/U1664/U32/Z ), .a(
        \I1/high/U1664/x[0] ) );
    aoi222_1 \I1/high/U1664/U29/U30/U1  ( .x(\I1/high/U1664/x[2] ), .a(
        \I1/high/ncd[5] ), .b(\I1/high/ncd[4] ), .c(\I1/high/ncd[5] ), .d(
        \I1/high/U1664/U29/Z ), .e(\I1/high/ncd[4] ), .f(\I1/high/U1664/U29/Z 
        ) );
    inv_1 \I1/high/U1664/U29/U30/Uinv  ( .x(\I1/high/U1664/U29/Z ), .a(
        \I1/high/U1664/x[2] ) );
    aoi222_1 \I1/high/U1664/U33/U30/U1  ( .x(\I1/high/U1664/y[0] ), .a(
        \I1/high/U1664/x[1] ), .b(\I1/high/U1664/x[0] ), .c(
        \I1/high/U1664/x[1] ), .d(\I1/high/U1664/U33/Z ), .e(
        \I1/high/U1664/x[0] ), .f(\I1/high/U1664/U33/Z ) );
    inv_1 \I1/high/U1664/U33/U30/Uinv  ( .x(\I1/high/U1664/U33/Z ), .a(
        \I1/high/U1664/y[0] ) );
    aoi222_1 \I1/high/U1664/U30/U30/U1  ( .x(\I1/high/U1664/y[1] ), .a(
        \I1/high/U1664/x[3] ), .b(\I1/high/U1664/x[2] ), .c(
        \I1/high/U1664/x[3] ), .d(\I1/high/U1664/U30/Z ), .e(
        \I1/high/U1664/x[2] ), .f(\I1/high/U1664/U30/Z ) );
    inv_1 \I1/high/U1664/U30/U30/Uinv  ( .x(\I1/high/U1664/U30/Z ), .a(
        \I1/high/U1664/y[1] ) );
    aoi222_1 \I1/high/U1664/U31/U30/U1  ( .x(\I1/high/U1664/x[1] ), .a(
        \I1/high/ncd[3] ), .b(\I1/high/ncd[2] ), .c(\I1/high/ncd[3] ), .d(
        \I1/high/U1664/U31/Z ), .e(\I1/high/ncd[2] ), .f(\I1/high/U1664/U31/Z 
        ) );
    inv_1 \I1/high/U1664/U31/U30/Uinv  ( .x(\I1/high/U1664/U31/Z ), .a(
        \I1/high/U1664/x[1] ) );
    aoi222_1 \I1/high/U1664/U37/U30/U1  ( .x(\I1/high/localcd ), .a(
        \I1/high/U1664/y[0] ), .b(\I1/high/U1664/y[1] ), .c(
        \I1/high/U1664/y[0] ), .d(\I1/high/U1664/U37/Z ), .e(
        \I1/high/U1664/y[1] ), .f(\I1/high/U1664/U37/Z ) );
    inv_1 \I1/high/U1664/U37/U30/Uinv  ( .x(\I1/high/U1664/U37/Z ), .a(
        \I1/high/localcd ) );
    nor3_1 \I1/high/U1669/Unr  ( .x(\I1/high/U1669/nr ), .a(
        \I1/high/ctrlack_internal ), .b(n8), .c(n11) );
    nand3_1 \I1/high/U1669/Und  ( .x(\I1/high/U1669/nd ), .a(
        \I1/high/ctrlack_internal ), .b(n8), .c(n11) );
    oa21_1 \I1/high/U1669/U1  ( .x(\I1/high/U1669/n2 ), .a(\I1/high/U1669/n2 ), 
        .b(\I1/high/U1669/nr ), .c(\I1/high/U1669/nd ) );
    inv_2 \I1/high/U1669/U3  ( .x(\I1/net20 ), .a(\I1/high/U1669/n2 ) );
    buf_2 U1 ( .x(n1), .a(\I0/net20 ) );
    buf_1 U2 ( .x(n2), .a(\I0/low/latch ) );
    buf_2 U3 ( .x(n3), .a(net17) );
    buf_1 U4 ( .x(n4), .a(\I0/high/latch ) );
    buf_2 U5 ( .x(n5), .a(\I1/net20 ) );
    buf_1 U6 ( .x(n6), .a(\I1/low/latch ) );
    inv_2 U7 ( .x(n7), .a(n9) );
    inv_1 U8 ( .x(n8), .a(n9) );
    inv_0 U9 ( .x(n9), .a(ctrlreq) );
    inv_2 U10 ( .x(n10), .a(n9) );
    inv_1 U11 ( .x(n11), .a(n9) );
    buf_1 U12 ( .x(n12), .a(\I1/high/latch ) );
endmodule


module chain_irdemux_32new_2 ( ctrlack, oh, ol, pullreq, pull_h, pull_l, 
    pullcd, reset, ctrlreq );
output [31:0] oh;
output [31:0] ol;
input  [7:0] pull_h;
input  [7:0] pull_l;
input  pullcd, reset, ctrlreq;
output ctrlack, pullreq;
    wire net30, net31, \I0/net32 , \I0/net33 , \I0/low/latch , 
        \I0/low/nlocalcd , \I0/low/localcd , \I0/low/ncd[0] , \I0/low/ncd[1] , 
        \I0/low/ncd[2] , \I0/low/ncd[3] , \I0/low/ncd[4] , \I0/low/ncd[5] , 
        \I0/low/ncd[6] , \I0/low/ncd[7] , \I0/low/ctrlack_internal , 
        \I0/low/acb , \I0/low/ba , \I0/low/driveh , \I0/net20 , 
        \I0/low/drivel , n1, n2, \I0/low/U4/U28/U1/clr , 
        \I0/low/U4/U28/U1/set , \I0/low/U1/Z , \I0/low/U1664/x[3] , 
        \I0/low/U1664/U28/Z , \I0/low/U1664/x[0] , \I0/low/U1664/U32/Z , 
        \I0/low/U1664/x[2] , \I0/low/U1664/U29/Z , \I0/low/U1664/y[0] , 
        \I0/low/U1664/x[1] , \I0/low/U1664/U33/Z , \I0/low/U1664/y[1] , 
        \I0/low/U1664/U30/Z , \I0/low/U1664/U31/Z , \I0/low/U1664/U37/Z , 
        \I0/low/U1669/nr , \I0/low/U1669/nd , \I0/low/U1669/n2 , 
        \I0/high/latch , \I0/high/nlocalcd , \I0/high/localcd , 
        \I0/high/ncd[0] , \I0/high/ncd[1] , \I0/high/ncd[2] , \I0/high/ncd[3] , 
        \I0/high/ncd[4] , \I0/high/ncd[5] , \I0/high/ncd[6] , \I0/high/ncd[7] , 
        \I0/high/ctrlack_internal , \I0/high/acb , \I0/high/ba , 
        \I0/high/driveh , net17, \I0/high/drivel , n3, n4, 
        \I0/high/U4/U28/U1/clr , \I0/high/U4/U28/U1/set , \I0/high/U1/Z , 
        \I0/high/U1664/x[3] , \I0/high/U1664/U28/Z , \I0/high/U1664/x[0] , 
        \I0/high/U1664/U32/Z , \I0/high/U1664/x[2] , \I0/high/U1664/U29/Z , 
        \I0/high/U1664/y[0] , \I0/high/U1664/x[1] , \I0/high/U1664/U33/Z , 
        \I0/high/U1664/y[1] , \I0/high/U1664/U30/Z , \I0/high/U1664/U31/Z , 
        \I0/high/U1664/U37/Z , \I0/high/U1669/nr , \I0/high/U1669/nd , 
        \I0/high/U1669/n2 , \I1/net32 , \I1/net33 , \I1/low/latch , 
        \I1/low/nlocalcd , \I1/low/localcd , \I1/low/ncd[0] , \I1/low/ncd[1] , 
        \I1/low/ncd[2] , \I1/low/ncd[3] , \I1/low/ncd[4] , \I1/low/ncd[5] , 
        \I1/low/ncd[6] , \I1/low/ncd[7] , \I1/low/ctrlack_internal , 
        \I1/low/acb , \I1/low/ba , \I1/low/driveh , \I1/net20 , 
        \I1/low/drivel , n5, n6, \I1/low/U4/U28/U1/clr , 
        \I1/low/U4/U28/U1/set , \I1/low/U1/Z , \I1/low/U1664/x[3] , 
        \I1/low/U1664/U28/Z , \I1/low/U1664/x[0] , \I1/low/U1664/U32/Z , 
        \I1/low/U1664/x[2] , \I1/low/U1664/U29/Z , \I1/low/U1664/y[0] , 
        \I1/low/U1664/x[1] , \I1/low/U1664/U33/Z , \I1/low/U1664/y[1] , 
        \I1/low/U1664/U30/Z , \I1/low/U1664/U31/Z , \I1/low/U1664/U37/Z , 
        \I1/low/U1669/nr , \I1/low/U1669/nd , \I1/low/U1669/n2 , 
        \I1/high/latch , \I1/high/nlocalcd , \I1/high/localcd , 
        \I1/high/ncd[0] , \I1/high/ncd[1] , \I1/high/ncd[2] , \I1/high/ncd[3] , 
        \I1/high/ncd[4] , \I1/high/ncd[5] , \I1/high/ncd[6] , \I1/high/ncd[7] , 
        \I1/high/ctrlack_internal , \I1/high/acb , \I1/high/ba , 
        \I1/high/driveh , \I1/high/drivel , n7, n8, \I1/high/U4/U28/U1/clr , 
        \I1/high/U4/U28/U1/set , \I1/high/U1/Z , \I1/high/U1664/x[3] , 
        \I1/high/U1664/U28/Z , \I1/high/U1664/x[0] , \I1/high/U1664/U32/Z , 
        \I1/high/U1664/x[2] , \I1/high/U1664/U29/Z , \I1/high/U1664/y[0] , 
        \I1/high/U1664/x[1] , \I1/high/U1664/U33/Z , \I1/high/U1664/y[1] , 
        \I1/high/U1664/U30/Z , \I1/high/U1664/U31/Z , \I1/high/U1664/U37/Z , 
        \I1/high/U1669/nr , \I1/high/U1669/nd , \I1/high/U1669/n2 ;
    nand2_1 \U3/U5  ( .x(pullreq), .a(net30), .b(net31) );
    nor2_1 \I0/U3/U5  ( .x(net30), .a(\I0/net32 ), .b(\I0/net33 ) );
    buf_2 \I0/low/U1653  ( .x(\I0/low/latch ), .a(\I0/net32 ) );
    nor2_1 \I0/low/U264/U5  ( .x(\I0/low/nlocalcd ), .a(reset), .b(
        \I0/low/localcd ) );
    nor2_1 \I0/low/U1659_0_/U5  ( .x(\I0/low/ncd[0] ), .a(ol[0]), .b(oh[0]) );
    nor2_1 \I0/low/U1659_1_/U5  ( .x(\I0/low/ncd[1] ), .a(ol[1]), .b(oh[1]) );
    nor2_1 \I0/low/U1659_2_/U5  ( .x(\I0/low/ncd[2] ), .a(ol[2]), .b(oh[2]) );
    nor2_1 \I0/low/U1659_3_/U5  ( .x(\I0/low/ncd[3] ), .a(ol[3]), .b(oh[3]) );
    nor2_1 \I0/low/U1659_4_/U5  ( .x(\I0/low/ncd[4] ), .a(ol[4]), .b(oh[4]) );
    nor2_1 \I0/low/U1659_5_/U5  ( .x(\I0/low/ncd[5] ), .a(ol[5]), .b(oh[5]) );
    nor2_1 \I0/low/U1659_6_/U5  ( .x(\I0/low/ncd[6] ), .a(ol[6]), .b(oh[6]) );
    nor2_1 \I0/low/U1659_7_/U5  ( .x(\I0/low/ncd[7] ), .a(ol[7]), .b(oh[7]) );
    nor2_1 \I0/low/U3/U5  ( .x(\I0/low/ctrlack_internal ), .a(\I0/low/acb ), 
        .b(\I0/low/ba ) );
    buf_2 \I0/low/U1665/U7  ( .x(\I0/low/driveh ), .a(\I0/net20 ) );
    buf_2 \I0/low/U1666/U7  ( .x(\I0/low/drivel ), .a(\I0/net20 ) );
    ao23_1 \I0/low/U1658_0_/U21/U1/U1  ( .x(ol[0]), .a(\I0/low/driveh ), .b(ol
        [0]), .c(n1), .d(pull_l[0]), .e(n2) );
    ao23_1 \I0/low/U1658_1_/U21/U1/U1  ( .x(ol[1]), .a(\I0/low/drivel ), .b(ol
        [1]), .c(\I0/low/driveh ), .d(pull_l[1]), .e(n2) );
    ao23_1 \I0/low/U1658_2_/U21/U1/U1  ( .x(ol[2]), .a(\I0/low/drivel ), .b(ol
        [2]), .c(\I0/low/driveh ), .d(pull_l[2]), .e(n2) );
    ao23_1 \I0/low/U1658_3_/U21/U1/U1  ( .x(ol[3]), .a(\I0/low/driveh ), .b(ol
        [3]), .c(\I0/low/drivel ), .d(pull_l[3]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_4_/U21/U1/U1  ( .x(ol[4]), .a(n1), .b(ol[4]), .c(
        \I0/low/drivel ), .d(pull_l[4]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_5_/U21/U1/U1  ( .x(ol[5]), .a(\I0/low/driveh ), .b(ol
        [5]), .c(n1), .d(pull_l[5]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_6_/U21/U1/U1  ( .x(ol[6]), .a(\I0/low/drivel ), .b(ol
        [6]), .c(\I0/low/driveh ), .d(pull_l[6]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1658_7_/U21/U1/U1  ( .x(ol[7]), .a(n1), .b(ol[7]), .c(n1), 
        .d(pull_l[7]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_0_/U21/U1/U1  ( .x(oh[0]), .a(\I0/low/driveh ), .b(oh
        [0]), .c(n1), .d(pull_h[0]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_1_/U21/U1/U1  ( .x(oh[1]), .a(n1), .b(oh[1]), .c(
        \I0/low/drivel ), .d(pull_h[1]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_2_/U21/U1/U1  ( .x(oh[2]), .a(\I0/low/drivel ), .b(oh
        [2]), .c(\I0/low/drivel ), .d(pull_h[2]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_3_/U21/U1/U1  ( .x(oh[3]), .a(n1), .b(oh[3]), .c(
        \I0/low/driveh ), .d(pull_h[3]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_4_/U21/U1/U1  ( .x(oh[4]), .a(n1), .b(oh[4]), .c(n1), 
        .d(pull_h[4]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_5_/U21/U1/U1  ( .x(oh[5]), .a(\I0/low/drivel ), .b(oh
        [5]), .c(n1), .d(pull_h[5]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_6_/U21/U1/U1  ( .x(oh[6]), .a(\I0/low/drivel ), .b(oh
        [6]), .c(\I0/low/driveh ), .d(pull_h[6]), .e(\I0/low/latch ) );
    ao23_1 \I0/low/U1651_7_/U21/U1/U1  ( .x(oh[7]), .a(\I0/low/driveh ), .b(oh
        [7]), .c(\I0/low/drivel ), .d(pull_h[7]), .e(\I0/low/latch ) );
    aoai211_1 \I0/low/U4/U28/U1/U1  ( .x(\I0/low/U4/U28/U1/clr ), .a(
        \I0/net20 ), .b(\I0/low/acb ), .c(\I0/low/nlocalcd ), .d(\I0/net32 )
         );
    nand3_1 \I0/low/U4/U28/U1/U2  ( .x(\I0/low/U4/U28/U1/set ), .a(
        \I0/low/nlocalcd ), .b(\I0/net20 ), .c(\I0/low/acb ) );
    nand2_2 \I0/low/U4/U28/U1/U3  ( .x(\I0/net32 ), .a(\I0/low/U4/U28/U1/clr ), 
        .b(\I0/low/U4/U28/U1/set ) );
    oai21_1 \I0/low/U1/U30/U1/U1  ( .x(\I0/low/acb ), .a(\I0/low/U1/Z ), .b(
        \I0/low/ba ), .c(\I0/net20 ) );
    inv_1 \I0/low/U1/U30/U1/U2  ( .x(\I0/low/U1/Z ), .a(\I0/low/acb ) );
    ao222_1 \I0/low/U5/U18/U1/U1  ( .x(\I0/low/ba ), .a(\I0/low/latch ), .b(
        pullcd), .c(\I0/low/latch ), .d(\I0/low/ba ), .e(pullcd), .f(
        \I0/low/ba ) );
    aoi222_1 \I0/low/U1664/U28/U30/U1  ( .x(\I0/low/U1664/x[3] ), .a(
        \I0/low/ncd[7] ), .b(\I0/low/ncd[6] ), .c(\I0/low/ncd[7] ), .d(
        \I0/low/U1664/U28/Z ), .e(\I0/low/ncd[6] ), .f(\I0/low/U1664/U28/Z )
         );
    inv_1 \I0/low/U1664/U28/U30/Uinv  ( .x(\I0/low/U1664/U28/Z ), .a(
        \I0/low/U1664/x[3] ) );
    aoi222_1 \I0/low/U1664/U32/U30/U1  ( .x(\I0/low/U1664/x[0] ), .a(
        \I0/low/ncd[1] ), .b(\I0/low/ncd[0] ), .c(\I0/low/ncd[1] ), .d(
        \I0/low/U1664/U32/Z ), .e(\I0/low/ncd[0] ), .f(\I0/low/U1664/U32/Z )
         );
    inv_1 \I0/low/U1664/U32/U30/Uinv  ( .x(\I0/low/U1664/U32/Z ), .a(
        \I0/low/U1664/x[0] ) );
    aoi222_1 \I0/low/U1664/U29/U30/U1  ( .x(\I0/low/U1664/x[2] ), .a(
        \I0/low/ncd[5] ), .b(\I0/low/ncd[4] ), .c(\I0/low/ncd[5] ), .d(
        \I0/low/U1664/U29/Z ), .e(\I0/low/ncd[4] ), .f(\I0/low/U1664/U29/Z )
         );
    inv_1 \I0/low/U1664/U29/U30/Uinv  ( .x(\I0/low/U1664/U29/Z ), .a(
        \I0/low/U1664/x[2] ) );
    aoi222_1 \I0/low/U1664/U33/U30/U1  ( .x(\I0/low/U1664/y[0] ), .a(
        \I0/low/U1664/x[1] ), .b(\I0/low/U1664/x[0] ), .c(\I0/low/U1664/x[1] ), 
        .d(\I0/low/U1664/U33/Z ), .e(\I0/low/U1664/x[0] ), .f(
        \I0/low/U1664/U33/Z ) );
    inv_1 \I0/low/U1664/U33/U30/Uinv  ( .x(\I0/low/U1664/U33/Z ), .a(
        \I0/low/U1664/y[0] ) );
    aoi222_1 \I0/low/U1664/U30/U30/U1  ( .x(\I0/low/U1664/y[1] ), .a(
        \I0/low/U1664/x[3] ), .b(\I0/low/U1664/x[2] ), .c(\I0/low/U1664/x[3] ), 
        .d(\I0/low/U1664/U30/Z ), .e(\I0/low/U1664/x[2] ), .f(
        \I0/low/U1664/U30/Z ) );
    inv_1 \I0/low/U1664/U30/U30/Uinv  ( .x(\I0/low/U1664/U30/Z ), .a(
        \I0/low/U1664/y[1] ) );
    aoi222_1 \I0/low/U1664/U31/U30/U1  ( .x(\I0/low/U1664/x[1] ), .a(
        \I0/low/ncd[3] ), .b(\I0/low/ncd[2] ), .c(\I0/low/ncd[3] ), .d(
        \I0/low/U1664/U31/Z ), .e(\I0/low/ncd[2] ), .f(\I0/low/U1664/U31/Z )
         );
    inv_1 \I0/low/U1664/U31/U30/Uinv  ( .x(\I0/low/U1664/U31/Z ), .a(
        \I0/low/U1664/x[1] ) );
    aoi222_1 \I0/low/U1664/U37/U30/U1  ( .x(\I0/low/localcd ), .a(
        \I0/low/U1664/y[0] ), .b(\I0/low/U1664/y[1] ), .c(\I0/low/U1664/y[0] ), 
        .d(\I0/low/U1664/U37/Z ), .e(\I0/low/U1664/y[1] ), .f(
        \I0/low/U1664/U37/Z ) );
    inv_1 \I0/low/U1664/U37/U30/Uinv  ( .x(\I0/low/U1664/U37/Z ), .a(
        \I0/low/localcd ) );
    nor3_1 \I0/low/U1669/Unr  ( .x(\I0/low/U1669/nr ), .a(
        \I0/low/ctrlack_internal ), .b(n1), .c(\I0/low/driveh ) );
    nand3_1 \I0/low/U1669/Und  ( .x(\I0/low/U1669/nd ), .a(
        \I0/low/ctrlack_internal ), .b(\I0/low/drivel ), .c(\I0/low/driveh )
         );
    oa21_1 \I0/low/U1669/U1  ( .x(\I0/low/U1669/n2 ), .a(\I0/low/U1669/n2 ), 
        .b(\I0/low/U1669/nr ), .c(\I0/low/U1669/nd ) );
    inv_2 \I0/low/U1669/U3  ( .x(ctrlack), .a(\I0/low/U1669/n2 ) );
    buf_2 \I0/high/U1653  ( .x(\I0/high/latch ), .a(\I0/net33 ) );
    nor2_1 \I0/high/U264/U5  ( .x(\I0/high/nlocalcd ), .a(reset), .b(
        \I0/high/localcd ) );
    nor2_1 \I0/high/U1659_0_/U5  ( .x(\I0/high/ncd[0] ), .a(ol[8]), .b(oh[8])
         );
    nor2_1 \I0/high/U1659_1_/U5  ( .x(\I0/high/ncd[1] ), .a(ol[9]), .b(oh[9])
         );
    nor2_1 \I0/high/U1659_2_/U5  ( .x(\I0/high/ncd[2] ), .a(ol[10]), .b(oh[10]
        ) );
    nor2_1 \I0/high/U1659_3_/U5  ( .x(\I0/high/ncd[3] ), .a(ol[11]), .b(oh[11]
        ) );
    nor2_1 \I0/high/U1659_4_/U5  ( .x(\I0/high/ncd[4] ), .a(ol[12]), .b(oh[12]
        ) );
    nor2_1 \I0/high/U1659_5_/U5  ( .x(\I0/high/ncd[5] ), .a(ol[13]), .b(oh[13]
        ) );
    nor2_1 \I0/high/U1659_6_/U5  ( .x(\I0/high/ncd[6] ), .a(ol[14]), .b(oh[14]
        ) );
    nor2_1 \I0/high/U1659_7_/U5  ( .x(\I0/high/ncd[7] ), .a(ol[15]), .b(oh[15]
        ) );
    nor2_1 \I0/high/U3/U5  ( .x(\I0/high/ctrlack_internal ), .a(\I0/high/acb ), 
        .b(\I0/high/ba ) );
    buf_2 \I0/high/U1665/U7  ( .x(\I0/high/driveh ), .a(net17) );
    buf_2 \I0/high/U1666/U7  ( .x(\I0/high/drivel ), .a(net17) );
    ao23_1 \I0/high/U1658_0_/U21/U1/U1  ( .x(ol[8]), .a(\I0/high/driveh ), .b(
        ol[8]), .c(n3), .d(pull_l[0]), .e(n4) );
    ao23_1 \I0/high/U1658_1_/U21/U1/U1  ( .x(ol[9]), .a(\I0/high/drivel ), .b(
        ol[9]), .c(\I0/high/driveh ), .d(pull_l[1]), .e(n4) );
    ao23_1 \I0/high/U1658_2_/U21/U1/U1  ( .x(ol[10]), .a(\I0/high/drivel ), 
        .b(ol[10]), .c(\I0/high/driveh ), .d(pull_l[2]), .e(n4) );
    ao23_1 \I0/high/U1658_3_/U21/U1/U1  ( .x(ol[11]), .a(\I0/high/driveh ), 
        .b(ol[11]), .c(\I0/high/drivel ), .d(pull_l[3]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1658_4_/U21/U1/U1  ( .x(ol[12]), .a(n3), .b(ol[12]), .c(
        \I0/high/drivel ), .d(pull_l[4]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1658_5_/U21/U1/U1  ( .x(ol[13]), .a(\I0/high/driveh ), 
        .b(ol[13]), .c(n3), .d(pull_l[5]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1658_6_/U21/U1/U1  ( .x(ol[14]), .a(\I0/high/drivel ), 
        .b(ol[14]), .c(\I0/high/driveh ), .d(pull_l[6]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1658_7_/U21/U1/U1  ( .x(ol[15]), .a(n3), .b(ol[15]), .c(
        n3), .d(pull_l[7]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_0_/U21/U1/U1  ( .x(oh[8]), .a(\I0/high/driveh ), .b(
        oh[8]), .c(n3), .d(pull_h[0]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_1_/U21/U1/U1  ( .x(oh[9]), .a(n3), .b(oh[9]), .c(
        \I0/high/drivel ), .d(pull_h[1]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_2_/U21/U1/U1  ( .x(oh[10]), .a(\I0/high/drivel ), 
        .b(oh[10]), .c(\I0/high/drivel ), .d(pull_h[2]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1651_3_/U21/U1/U1  ( .x(oh[11]), .a(n3), .b(oh[11]), .c(
        \I0/high/driveh ), .d(pull_h[3]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_4_/U21/U1/U1  ( .x(oh[12]), .a(n3), .b(oh[12]), .c(
        n3), .d(pull_h[4]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_5_/U21/U1/U1  ( .x(oh[13]), .a(\I0/high/drivel ), 
        .b(oh[13]), .c(n3), .d(pull_h[5]), .e(\I0/high/latch ) );
    ao23_1 \I0/high/U1651_6_/U21/U1/U1  ( .x(oh[14]), .a(\I0/high/drivel ), 
        .b(oh[14]), .c(\I0/high/driveh ), .d(pull_h[6]), .e(\I0/high/latch )
         );
    ao23_1 \I0/high/U1651_7_/U21/U1/U1  ( .x(oh[15]), .a(\I0/high/driveh ), 
        .b(oh[15]), .c(\I0/high/drivel ), .d(pull_h[7]), .e(\I0/high/latch )
         );
    aoai211_1 \I0/high/U4/U28/U1/U1  ( .x(\I0/high/U4/U28/U1/clr ), .a(net17), 
        .b(\I0/high/acb ), .c(\I0/high/nlocalcd ), .d(\I0/net33 ) );
    nand3_1 \I0/high/U4/U28/U1/U2  ( .x(\I0/high/U4/U28/U1/set ), .a(
        \I0/high/nlocalcd ), .b(net17), .c(\I0/high/acb ) );
    nand2_2 \I0/high/U4/U28/U1/U3  ( .x(\I0/net33 ), .a(
        \I0/high/U4/U28/U1/clr ), .b(\I0/high/U4/U28/U1/set ) );
    oai21_1 \I0/high/U1/U30/U1/U1  ( .x(\I0/high/acb ), .a(\I0/high/U1/Z ), 
        .b(\I0/high/ba ), .c(net17) );
    inv_1 \I0/high/U1/U30/U1/U2  ( .x(\I0/high/U1/Z ), .a(\I0/high/acb ) );
    ao222_1 \I0/high/U5/U18/U1/U1  ( .x(\I0/high/ba ), .a(\I0/high/latch ), 
        .b(pullcd), .c(\I0/high/latch ), .d(\I0/high/ba ), .e(pullcd), .f(
        \I0/high/ba ) );
    aoi222_1 \I0/high/U1664/U28/U30/U1  ( .x(\I0/high/U1664/x[3] ), .a(
        \I0/high/ncd[7] ), .b(\I0/high/ncd[6] ), .c(\I0/high/ncd[7] ), .d(
        \I0/high/U1664/U28/Z ), .e(\I0/high/ncd[6] ), .f(\I0/high/U1664/U28/Z 
        ) );
    inv_1 \I0/high/U1664/U28/U30/Uinv  ( .x(\I0/high/U1664/U28/Z ), .a(
        \I0/high/U1664/x[3] ) );
    aoi222_1 \I0/high/U1664/U32/U30/U1  ( .x(\I0/high/U1664/x[0] ), .a(
        \I0/high/ncd[1] ), .b(\I0/high/ncd[0] ), .c(\I0/high/ncd[1] ), .d(
        \I0/high/U1664/U32/Z ), .e(\I0/high/ncd[0] ), .f(\I0/high/U1664/U32/Z 
        ) );
    inv_1 \I0/high/U1664/U32/U30/Uinv  ( .x(\I0/high/U1664/U32/Z ), .a(
        \I0/high/U1664/x[0] ) );
    aoi222_1 \I0/high/U1664/U29/U30/U1  ( .x(\I0/high/U1664/x[2] ), .a(
        \I0/high/ncd[5] ), .b(\I0/high/ncd[4] ), .c(\I0/high/ncd[5] ), .d(
        \I0/high/U1664/U29/Z ), .e(\I0/high/ncd[4] ), .f(\I0/high/U1664/U29/Z 
        ) );
    inv_1 \I0/high/U1664/U29/U30/Uinv  ( .x(\I0/high/U1664/U29/Z ), .a(
        \I0/high/U1664/x[2] ) );
    aoi222_1 \I0/high/U1664/U33/U30/U1  ( .x(\I0/high/U1664/y[0] ), .a(
        \I0/high/U1664/x[1] ), .b(\I0/high/U1664/x[0] ), .c(
        \I0/high/U1664/x[1] ), .d(\I0/high/U1664/U33/Z ), .e(
        \I0/high/U1664/x[0] ), .f(\I0/high/U1664/U33/Z ) );
    inv_1 \I0/high/U1664/U33/U30/Uinv  ( .x(\I0/high/U1664/U33/Z ), .a(
        \I0/high/U1664/y[0] ) );
    aoi222_1 \I0/high/U1664/U30/U30/U1  ( .x(\I0/high/U1664/y[1] ), .a(
        \I0/high/U1664/x[3] ), .b(\I0/high/U1664/x[2] ), .c(
        \I0/high/U1664/x[3] ), .d(\I0/high/U1664/U30/Z ), .e(
        \I0/high/U1664/x[2] ), .f(\I0/high/U1664/U30/Z ) );
    inv_1 \I0/high/U1664/U30/U30/Uinv  ( .x(\I0/high/U1664/U30/Z ), .a(
        \I0/high/U1664/y[1] ) );
    aoi222_1 \I0/high/U1664/U31/U30/U1  ( .x(\I0/high/U1664/x[1] ), .a(
        \I0/high/ncd[3] ), .b(\I0/high/ncd[2] ), .c(\I0/high/ncd[3] ), .d(
        \I0/high/U1664/U31/Z ), .e(\I0/high/ncd[2] ), .f(\I0/high/U1664/U31/Z 
        ) );
    inv_1 \I0/high/U1664/U31/U30/Uinv  ( .x(\I0/high/U1664/U31/Z ), .a(
        \I0/high/U1664/x[1] ) );
    aoi222_1 \I0/high/U1664/U37/U30/U1  ( .x(\I0/high/localcd ), .a(
        \I0/high/U1664/y[0] ), .b(\I0/high/U1664/y[1] ), .c(
        \I0/high/U1664/y[0] ), .d(\I0/high/U1664/U37/Z ), .e(
        \I0/high/U1664/y[1] ), .f(\I0/high/U1664/U37/Z ) );
    inv_1 \I0/high/U1664/U37/U30/Uinv  ( .x(\I0/high/U1664/U37/Z ), .a(
        \I0/high/localcd ) );
    nor3_1 \I0/high/U1669/Unr  ( .x(\I0/high/U1669/nr ), .a(
        \I0/high/ctrlack_internal ), .b(n3), .c(\I0/high/driveh ) );
    nand3_1 \I0/high/U1669/Und  ( .x(\I0/high/U1669/nd ), .a(
        \I0/high/ctrlack_internal ), .b(\I0/high/drivel ), .c(\I0/high/driveh 
        ) );
    oa21_1 \I0/high/U1669/U1  ( .x(\I0/high/U1669/n2 ), .a(\I0/high/U1669/n2 ), 
        .b(\I0/high/U1669/nr ), .c(\I0/high/U1669/nd ) );
    inv_2 \I0/high/U1669/U3  ( .x(\I0/net20 ), .a(\I0/high/U1669/n2 ) );
    nor2_1 \I1/U3/U5  ( .x(net31), .a(\I1/net32 ), .b(\I1/net33 ) );
    buf_2 \I1/low/U1653  ( .x(\I1/low/latch ), .a(\I1/net32 ) );
    nor2_1 \I1/low/U264/U5  ( .x(\I1/low/nlocalcd ), .a(reset), .b(
        \I1/low/localcd ) );
    nor2_1 \I1/low/U1659_0_/U5  ( .x(\I1/low/ncd[0] ), .a(ol[16]), .b(oh[16])
         );
    nor2_1 \I1/low/U1659_1_/U5  ( .x(\I1/low/ncd[1] ), .a(ol[17]), .b(oh[17])
         );
    nor2_1 \I1/low/U1659_2_/U5  ( .x(\I1/low/ncd[2] ), .a(ol[18]), .b(oh[18])
         );
    nor2_1 \I1/low/U1659_3_/U5  ( .x(\I1/low/ncd[3] ), .a(ol[19]), .b(oh[19])
         );
    nor2_1 \I1/low/U1659_4_/U5  ( .x(\I1/low/ncd[4] ), .a(ol[20]), .b(oh[20])
         );
    nor2_1 \I1/low/U1659_5_/U5  ( .x(\I1/low/ncd[5] ), .a(ol[21]), .b(oh[21])
         );
    nor2_1 \I1/low/U1659_6_/U5  ( .x(\I1/low/ncd[6] ), .a(ol[22]), .b(oh[22])
         );
    nor2_1 \I1/low/U1659_7_/U5  ( .x(\I1/low/ncd[7] ), .a(ol[23]), .b(oh[23])
         );
    nor2_1 \I1/low/U3/U5  ( .x(\I1/low/ctrlack_internal ), .a(\I1/low/acb ), 
        .b(\I1/low/ba ) );
    buf_2 \I1/low/U1665/U7  ( .x(\I1/low/driveh ), .a(\I1/net20 ) );
    buf_2 \I1/low/U1666/U7  ( .x(\I1/low/drivel ), .a(\I1/net20 ) );
    ao23_1 \I1/low/U1658_0_/U21/U1/U1  ( .x(ol[16]), .a(\I1/low/driveh ), .b(
        ol[16]), .c(n5), .d(pull_l[0]), .e(n6) );
    ao23_1 \I1/low/U1658_1_/U21/U1/U1  ( .x(ol[17]), .a(\I1/low/drivel ), .b(
        ol[17]), .c(\I1/low/driveh ), .d(pull_l[1]), .e(n6) );
    ao23_1 \I1/low/U1658_2_/U21/U1/U1  ( .x(ol[18]), .a(\I1/low/drivel ), .b(
        ol[18]), .c(\I1/low/driveh ), .d(pull_l[2]), .e(n6) );
    ao23_1 \I1/low/U1658_3_/U21/U1/U1  ( .x(ol[19]), .a(\I1/low/driveh ), .b(
        ol[19]), .c(\I1/low/drivel ), .d(pull_l[3]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_4_/U21/U1/U1  ( .x(ol[20]), .a(n5), .b(ol[20]), .c(
        \I1/low/drivel ), .d(pull_l[4]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_5_/U21/U1/U1  ( .x(ol[21]), .a(\I1/low/driveh ), .b(
        ol[21]), .c(n5), .d(pull_l[5]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_6_/U21/U1/U1  ( .x(ol[22]), .a(\I1/low/drivel ), .b(
        ol[22]), .c(\I1/low/driveh ), .d(pull_l[6]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1658_7_/U21/U1/U1  ( .x(ol[23]), .a(n5), .b(ol[23]), .c(n5
        ), .d(pull_l[7]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_0_/U21/U1/U1  ( .x(oh[16]), .a(\I1/low/driveh ), .b(
        oh[16]), .c(n5), .d(pull_h[0]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_1_/U21/U1/U1  ( .x(oh[17]), .a(n5), .b(oh[17]), .c(
        \I1/low/drivel ), .d(pull_h[1]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_2_/U21/U1/U1  ( .x(oh[18]), .a(\I1/low/drivel ), .b(
        oh[18]), .c(\I1/low/drivel ), .d(pull_h[2]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_3_/U21/U1/U1  ( .x(oh[19]), .a(n5), .b(oh[19]), .c(
        \I1/low/driveh ), .d(pull_h[3]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_4_/U21/U1/U1  ( .x(oh[20]), .a(n5), .b(oh[20]), .c(n5
        ), .d(pull_h[4]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_5_/U21/U1/U1  ( .x(oh[21]), .a(\I1/low/drivel ), .b(
        oh[21]), .c(n5), .d(pull_h[5]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_6_/U21/U1/U1  ( .x(oh[22]), .a(\I1/low/drivel ), .b(
        oh[22]), .c(\I1/low/driveh ), .d(pull_h[6]), .e(\I1/low/latch ) );
    ao23_1 \I1/low/U1651_7_/U21/U1/U1  ( .x(oh[23]), .a(\I1/low/driveh ), .b(
        oh[23]), .c(\I1/low/drivel ), .d(pull_h[7]), .e(\I1/low/latch ) );
    aoai211_1 \I1/low/U4/U28/U1/U1  ( .x(\I1/low/U4/U28/U1/clr ), .a(
        \I1/net20 ), .b(\I1/low/acb ), .c(\I1/low/nlocalcd ), .d(\I1/net32 )
         );
    nand3_1 \I1/low/U4/U28/U1/U2  ( .x(\I1/low/U4/U28/U1/set ), .a(
        \I1/low/nlocalcd ), .b(\I1/net20 ), .c(\I1/low/acb ) );
    nand2_2 \I1/low/U4/U28/U1/U3  ( .x(\I1/net32 ), .a(\I1/low/U4/U28/U1/clr ), 
        .b(\I1/low/U4/U28/U1/set ) );
    oai21_1 \I1/low/U1/U30/U1/U1  ( .x(\I1/low/acb ), .a(\I1/low/U1/Z ), .b(
        \I1/low/ba ), .c(\I1/net20 ) );
    inv_1 \I1/low/U1/U30/U1/U2  ( .x(\I1/low/U1/Z ), .a(\I1/low/acb ) );
    ao222_1 \I1/low/U5/U18/U1/U1  ( .x(\I1/low/ba ), .a(\I1/low/latch ), .b(
        pullcd), .c(\I1/low/latch ), .d(\I1/low/ba ), .e(pullcd), .f(
        \I1/low/ba ) );
    aoi222_1 \I1/low/U1664/U28/U30/U1  ( .x(\I1/low/U1664/x[3] ), .a(
        \I1/low/ncd[7] ), .b(\I1/low/ncd[6] ), .c(\I1/low/ncd[7] ), .d(
        \I1/low/U1664/U28/Z ), .e(\I1/low/ncd[6] ), .f(\I1/low/U1664/U28/Z )
         );
    inv_1 \I1/low/U1664/U28/U30/Uinv  ( .x(\I1/low/U1664/U28/Z ), .a(
        \I1/low/U1664/x[3] ) );
    aoi222_1 \I1/low/U1664/U32/U30/U1  ( .x(\I1/low/U1664/x[0] ), .a(
        \I1/low/ncd[1] ), .b(\I1/low/ncd[0] ), .c(\I1/low/ncd[1] ), .d(
        \I1/low/U1664/U32/Z ), .e(\I1/low/ncd[0] ), .f(\I1/low/U1664/U32/Z )
         );
    inv_1 \I1/low/U1664/U32/U30/Uinv  ( .x(\I1/low/U1664/U32/Z ), .a(
        \I1/low/U1664/x[0] ) );
    aoi222_1 \I1/low/U1664/U29/U30/U1  ( .x(\I1/low/U1664/x[2] ), .a(
        \I1/low/ncd[5] ), .b(\I1/low/ncd[4] ), .c(\I1/low/ncd[5] ), .d(
        \I1/low/U1664/U29/Z ), .e(\I1/low/ncd[4] ), .f(\I1/low/U1664/U29/Z )
         );
    inv_1 \I1/low/U1664/U29/U30/Uinv  ( .x(\I1/low/U1664/U29/Z ), .a(
        \I1/low/U1664/x[2] ) );
    aoi222_1 \I1/low/U1664/U33/U30/U1  ( .x(\I1/low/U1664/y[0] ), .a(
        \I1/low/U1664/x[1] ), .b(\I1/low/U1664/x[0] ), .c(\I1/low/U1664/x[1] ), 
        .d(\I1/low/U1664/U33/Z ), .e(\I1/low/U1664/x[0] ), .f(
        \I1/low/U1664/U33/Z ) );
    inv_1 \I1/low/U1664/U33/U30/Uinv  ( .x(\I1/low/U1664/U33/Z ), .a(
        \I1/low/U1664/y[0] ) );
    aoi222_1 \I1/low/U1664/U30/U30/U1  ( .x(\I1/low/U1664/y[1] ), .a(
        \I1/low/U1664/x[3] ), .b(\I1/low/U1664/x[2] ), .c(\I1/low/U1664/x[3] ), 
        .d(\I1/low/U1664/U30/Z ), .e(\I1/low/U1664/x[2] ), .f(
        \I1/low/U1664/U30/Z ) );
    inv_1 \I1/low/U1664/U30/U30/Uinv  ( .x(\I1/low/U1664/U30/Z ), .a(
        \I1/low/U1664/y[1] ) );
    aoi222_1 \I1/low/U1664/U31/U30/U1  ( .x(\I1/low/U1664/x[1] ), .a(
        \I1/low/ncd[3] ), .b(\I1/low/ncd[2] ), .c(\I1/low/ncd[3] ), .d(
        \I1/low/U1664/U31/Z ), .e(\I1/low/ncd[2] ), .f(\I1/low/U1664/U31/Z )
         );
    inv_1 \I1/low/U1664/U31/U30/Uinv  ( .x(\I1/low/U1664/U31/Z ), .a(
        \I1/low/U1664/x[1] ) );
    aoi222_1 \I1/low/U1664/U37/U30/U1  ( .x(\I1/low/localcd ), .a(
        \I1/low/U1664/y[0] ), .b(\I1/low/U1664/y[1] ), .c(\I1/low/U1664/y[0] ), 
        .d(\I1/low/U1664/U37/Z ), .e(\I1/low/U1664/y[1] ), .f(
        \I1/low/U1664/U37/Z ) );
    inv_1 \I1/low/U1664/U37/U30/Uinv  ( .x(\I1/low/U1664/U37/Z ), .a(
        \I1/low/localcd ) );
    nor3_1 \I1/low/U1669/Unr  ( .x(\I1/low/U1669/nr ), .a(
        \I1/low/ctrlack_internal ), .b(n5), .c(\I1/low/driveh ) );
    nand3_1 \I1/low/U1669/Und  ( .x(\I1/low/U1669/nd ), .a(
        \I1/low/ctrlack_internal ), .b(\I1/low/drivel ), .c(\I1/low/driveh )
         );
    oa21_1 \I1/low/U1669/U1  ( .x(\I1/low/U1669/n2 ), .a(\I1/low/U1669/n2 ), 
        .b(\I1/low/U1669/nr ), .c(\I1/low/U1669/nd ) );
    inv_2 \I1/low/U1669/U3  ( .x(net17), .a(\I1/low/U1669/n2 ) );
    buf_2 \I1/high/U1653  ( .x(\I1/high/latch ), .a(\I1/net33 ) );
    nor2_1 \I1/high/U264/U5  ( .x(\I1/high/nlocalcd ), .a(reset), .b(
        \I1/high/localcd ) );
    nor2_1 \I1/high/U1659_0_/U5  ( .x(\I1/high/ncd[0] ), .a(ol[24]), .b(oh[24]
        ) );
    nor2_1 \I1/high/U1659_1_/U5  ( .x(\I1/high/ncd[1] ), .a(ol[25]), .b(oh[25]
        ) );
    nor2_1 \I1/high/U1659_2_/U5  ( .x(\I1/high/ncd[2] ), .a(ol[26]), .b(oh[26]
        ) );
    nor2_1 \I1/high/U1659_3_/U5  ( .x(\I1/high/ncd[3] ), .a(ol[27]), .b(oh[27]
        ) );
    nor2_1 \I1/high/U1659_4_/U5  ( .x(\I1/high/ncd[4] ), .a(ol[28]), .b(oh[28]
        ) );
    nor2_1 \I1/high/U1659_5_/U5  ( .x(\I1/high/ncd[5] ), .a(ol[29]), .b(oh[29]
        ) );
    nor2_1 \I1/high/U1659_6_/U5  ( .x(\I1/high/ncd[6] ), .a(ol[30]), .b(oh[30]
        ) );
    nor2_1 \I1/high/U1659_7_/U5  ( .x(\I1/high/ncd[7] ), .a(ol[31]), .b(oh[31]
        ) );
    nor2_1 \I1/high/U3/U5  ( .x(\I1/high/ctrlack_internal ), .a(\I1/high/acb ), 
        .b(\I1/high/ba ) );
    buf_2 \I1/high/U1665/U7  ( .x(\I1/high/driveh ), .a(ctrlreq) );
    buf_2 \I1/high/U1666/U7  ( .x(\I1/high/drivel ), .a(ctrlreq) );
    ao23_1 \I1/high/U1658_0_/U21/U1/U1  ( .x(ol[24]), .a(\I1/high/driveh ), 
        .b(ol[24]), .c(n7), .d(pull_l[0]), .e(n8) );
    ao23_1 \I1/high/U1658_1_/U21/U1/U1  ( .x(ol[25]), .a(\I1/high/drivel ), 
        .b(ol[25]), .c(\I1/high/driveh ), .d(pull_l[1]), .e(n8) );
    ao23_1 \I1/high/U1658_2_/U21/U1/U1  ( .x(ol[26]), .a(\I1/high/drivel ), 
        .b(ol[26]), .c(\I1/high/driveh ), .d(pull_l[2]), .e(n8) );
    ao23_1 \I1/high/U1658_3_/U21/U1/U1  ( .x(ol[27]), .a(\I1/high/driveh ), 
        .b(ol[27]), .c(\I1/high/drivel ), .d(pull_l[3]), .e(\I1/high/latch )
         );
    ao23_1 \I1/high/U1658_4_/U21/U1/U1  ( .x(ol[28]), .a(n7), .b(ol[28]), .c(
        \I1/high/drivel ), .d(pull_l[4]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1658_5_/U21/U1/U1  ( .x(ol[29]), .a(\I1/high/driveh ), 
        .b(ol[29]), .c(n7), .d(pull_l[5]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1658_6_/U21/U1/U1  ( .x(ol[30]), .a(\I1/high/drivel ), 
        .b(ol[30]), .c(\I1/high/driveh ), .d(pull_l[6]), .e(\I1/high/latch )
         );
    ao23_1 \I1/high/U1658_7_/U21/U1/U1  ( .x(ol[31]), .a(n7), .b(ol[31]), .c(
        n7), .d(pull_l[7]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_0_/U21/U1/U1  ( .x(oh[24]), .a(\I1/high/driveh ), 
        .b(oh[24]), .c(n7), .d(pull_h[0]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_1_/U21/U1/U1  ( .x(oh[25]), .a(n7), .b(oh[25]), .c(
        \I1/high/drivel ), .d(pull_h[1]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_2_/U21/U1/U1  ( .x(oh[26]), .a(\I1/high/drivel ), 
        .b(oh[26]), .c(\I1/high/drivel ), .d(pull_h[2]), .e(\I1/high/latch )
         );
    ao23_1 \I1/high/U1651_3_/U21/U1/U1  ( .x(oh[27]), .a(n7), .b(oh[27]), .c(
        \I1/high/driveh ), .d(pull_h[3]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_4_/U21/U1/U1  ( .x(oh[28]), .a(n7), .b(oh[28]), .c(
        n7), .d(pull_h[4]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_5_/U21/U1/U1  ( .x(oh[29]), .a(\I1/high/drivel ), 
        .b(oh[29]), .c(n7), .d(pull_h[5]), .e(\I1/high/latch ) );
    ao23_1 \I1/high/U1651_6_/U21/U1/U1  ( .x(oh[30]), .a(\I1/high/drivel ), 
        .b(oh[30]), .c(\I1/high/driveh ), .d(pull_h[6]), .e(\I1/high/latch )
         );
    ao23_1 \I1/high/U1651_7_/U21/U1/U1  ( .x(oh[31]), .a(\I1/high/driveh ), 
        .b(oh[31]), .c(\I1/high/drivel ), .d(pull_h[7]), .e(\I1/high/latch )
         );
    aoai211_1 \I1/high/U4/U28/U1/U1  ( .x(\I1/high/U4/U28/U1/clr ), .a(ctrlreq
        ), .b(\I1/high/acb ), .c(\I1/high/nlocalcd ), .d(\I1/net33 ) );
    nand3_1 \I1/high/U4/U28/U1/U2  ( .x(\I1/high/U4/U28/U1/set ), .a(
        \I1/high/nlocalcd ), .b(ctrlreq), .c(\I1/high/acb ) );
    nand2_2 \I1/high/U4/U28/U1/U3  ( .x(\I1/net33 ), .a(
        \I1/high/U4/U28/U1/clr ), .b(\I1/high/U4/U28/U1/set ) );
    oai21_1 \I1/high/U1/U30/U1/U1  ( .x(\I1/high/acb ), .a(\I1/high/U1/Z ), 
        .b(\I1/high/ba ), .c(ctrlreq) );
    inv_1 \I1/high/U1/U30/U1/U2  ( .x(\I1/high/U1/Z ), .a(\I1/high/acb ) );
    ao222_1 \I1/high/U5/U18/U1/U1  ( .x(\I1/high/ba ), .a(\I1/high/latch ), 
        .b(pullcd), .c(\I1/high/latch ), .d(\I1/high/ba ), .e(pullcd), .f(
        \I1/high/ba ) );
    aoi222_1 \I1/high/U1664/U28/U30/U1  ( .x(\I1/high/U1664/x[3] ), .a(
        \I1/high/ncd[7] ), .b(\I1/high/ncd[6] ), .c(\I1/high/ncd[7] ), .d(
        \I1/high/U1664/U28/Z ), .e(\I1/high/ncd[6] ), .f(\I1/high/U1664/U28/Z 
        ) );
    inv_1 \I1/high/U1664/U28/U30/Uinv  ( .x(\I1/high/U1664/U28/Z ), .a(
        \I1/high/U1664/x[3] ) );
    aoi222_1 \I1/high/U1664/U32/U30/U1  ( .x(\I1/high/U1664/x[0] ), .a(
        \I1/high/ncd[1] ), .b(\I1/high/ncd[0] ), .c(\I1/high/ncd[1] ), .d(
        \I1/high/U1664/U32/Z ), .e(\I1/high/ncd[0] ), .f(\I1/high/U1664/U32/Z 
        ) );
    inv_1 \I1/high/U1664/U32/U30/Uinv  ( .x(\I1/high/U1664/U32/Z ), .a(
        \I1/high/U1664/x[0] ) );
    aoi222_1 \I1/high/U1664/U29/U30/U1  ( .x(\I1/high/U1664/x[2] ), .a(
        \I1/high/ncd[5] ), .b(\I1/high/ncd[4] ), .c(\I1/high/ncd[5] ), .d(
        \I1/high/U1664/U29/Z ), .e(\I1/high/ncd[4] ), .f(\I1/high/U1664/U29/Z 
        ) );
    inv_1 \I1/high/U1664/U29/U30/Uinv  ( .x(\I1/high/U1664/U29/Z ), .a(
        \I1/high/U1664/x[2] ) );
    aoi222_1 \I1/high/U1664/U33/U30/U1  ( .x(\I1/high/U1664/y[0] ), .a(
        \I1/high/U1664/x[1] ), .b(\I1/high/U1664/x[0] ), .c(
        \I1/high/U1664/x[1] ), .d(\I1/high/U1664/U33/Z ), .e(
        \I1/high/U1664/x[0] ), .f(\I1/high/U1664/U33/Z ) );
    inv_1 \I1/high/U1664/U33/U30/Uinv  ( .x(\I1/high/U1664/U33/Z ), .a(
        \I1/high/U1664/y[0] ) );
    aoi222_1 \I1/high/U1664/U30/U30/U1  ( .x(\I1/high/U1664/y[1] ), .a(
        \I1/high/U1664/x[3] ), .b(\I1/high/U1664/x[2] ), .c(
        \I1/high/U1664/x[3] ), .d(\I1/high/U1664/U30/Z ), .e(
        \I1/high/U1664/x[2] ), .f(\I1/high/U1664/U30/Z ) );
    inv_1 \I1/high/U1664/U30/U30/Uinv  ( .x(\I1/high/U1664/U30/Z ), .a(
        \I1/high/U1664/y[1] ) );
    aoi222_1 \I1/high/U1664/U31/U30/U1  ( .x(\I1/high/U1664/x[1] ), .a(
        \I1/high/ncd[3] ), .b(\I1/high/ncd[2] ), .c(\I1/high/ncd[3] ), .d(
        \I1/high/U1664/U31/Z ), .e(\I1/high/ncd[2] ), .f(\I1/high/U1664/U31/Z 
        ) );
    inv_1 \I1/high/U1664/U31/U30/Uinv  ( .x(\I1/high/U1664/U31/Z ), .a(
        \I1/high/U1664/x[1] ) );
    aoi222_1 \I1/high/U1664/U37/U30/U1  ( .x(\I1/high/localcd ), .a(
        \I1/high/U1664/y[0] ), .b(\I1/high/U1664/y[1] ), .c(
        \I1/high/U1664/y[0] ), .d(\I1/high/U1664/U37/Z ), .e(
        \I1/high/U1664/y[1] ), .f(\I1/high/U1664/U37/Z ) );
    inv_1 \I1/high/U1664/U37/U30/Uinv  ( .x(\I1/high/U1664/U37/Z ), .a(
        \I1/high/localcd ) );
    nor3_1 \I1/high/U1669/Unr  ( .x(\I1/high/U1669/nr ), .a(
        \I1/high/ctrlack_internal ), .b(n7), .c(\I1/high/driveh ) );
    nand3_1 \I1/high/U1669/Und  ( .x(\I1/high/U1669/nd ), .a(
        \I1/high/ctrlack_internal ), .b(\I1/high/drivel ), .c(\I1/high/driveh 
        ) );
    oa21_1 \I1/high/U1669/U1  ( .x(\I1/high/U1669/n2 ), .a(\I1/high/U1669/n2 ), 
        .b(\I1/high/U1669/nr ), .c(\I1/high/U1669/nd ) );
    inv_2 \I1/high/U1669/U3  ( .x(\I1/net20 ), .a(\I1/high/U1669/n2 ) );
    buf_2 U1 ( .x(n1), .a(\I0/net20 ) );
    buf_1 U2 ( .x(n2), .a(\I0/low/latch ) );
    buf_2 U3 ( .x(n3), .a(net17) );
    buf_1 U4 ( .x(n4), .a(\I0/high/latch ) );
    buf_2 U5 ( .x(n5), .a(\I1/net20 ) );
    buf_1 U6 ( .x(n6), .a(\I1/low/latch ) );
    buf_2 U7 ( .x(n7), .a(ctrlreq) );
    buf_1 U8 ( .x(n8), .a(\I1/high/latch ) );
endmodule


module chain_fr2dr_byte_1 ( nia, oh, ol, i, nReset, noa );
output [7:0] oh;
output [7:0] ol;
input  [4:0] i;
input  nReset, noa;
output nia;
    wire nbReset, eop, ncla, csela, asela, \U891/reset , \U891/neopack , 
        \U891/iay , \U891/naack[0] , \U891/naack[1] , \U891/U1128/nb , \b[3] , 
        \b[2] , \U891/U1128/na , \b[1] , \b[0] , \U891/ackb , \a[3] , \a[2] , 
        \U891/nack , \U891/acka , \a[1] , \a[0] , bsela, bsel, asel, 
        \U891/U1118_0_/nr , naa, \U891/U1118_0_/nd , \U891/U1118_0_/n2 , 
        \U891/U1118_1_/nr , \U891/U1118_1_/nd , \U891/U1118_1_/n2 , 
        \U891/U1118_2_/nr , \U891/U1118_2_/nd , \U891/U1118_2_/n2 , 
        \U891/U1118_3_/nr , \U891/U1118_3_/nd , \U891/U1118_3_/n2 , 
        \U891/U1117_0_/nr , nba, \U891/U1117_0_/nd , \U891/U1117_0_/n2 , 
        \U891/U1117_1_/nr , \U891/U1117_1_/nd , \U891/U1117_1_/n2 , 
        \U891/U1117_2_/nr , \U891/U1117_2_/nd , \U891/U1117_2_/n2 , 
        \U891/U1117_3_/nr , \U891/U1117_3_/nd , \U891/U1117_3_/n2 , 
        \U886/reset , \U886/U1128/nb , \f[3] , \f[2] , \U886/U1128/na , \f[1] , 
        \f[0] , \U886/ackb , \U886/nack , \U886/acka , \U886/U1127/n5 , 
        \U886/U1127/n1 , \U886/U1127/n2 , \U886/U1127/n3 , \U886/U1127/n4 , 
        \e[3] , \e[2] , \e[1] , \e[0] , fsela, fsel, esela, esel, 
        \U886/U1118_0_/nr , nea, \U886/U1118_0_/nd , \U886/U1118_0_/n2 , 
        \U886/U1118_1_/nr , \U886/U1118_1_/nd , \U886/U1118_1_/n2 , 
        \U886/U1118_2_/nr , \U886/U1118_2_/nd , \U886/U1118_2_/n2 , 
        \U886/U1118_3_/nr , \U886/U1118_3_/nd , \U886/U1118_3_/n2 , 
        \U886/U1117_0_/nr , nfa, \U886/U1117_0_/nd , \U886/U1117_0_/n2 , 
        \U886/U1117_1_/nr , \U886/U1117_1_/nd , \U886/U1117_1_/n2 , 
        \U886/U1117_2_/nr , \U886/U1117_2_/nd , \U886/U1117_2_/n2 , 
        \U886/U1117_3_/nr , \U886/U1117_3_/nd , \U886/U1117_3_/n2 , 
        \U884/reset , \U884/U1128/nb , \d[3] , \d[2] , \U884/U1128/na , \d[1] , 
        \d[0] , \U884/ackb , \U884/nack , \U884/acka , \U884/U1127/n5 , 
        \U884/U1127/n1 , \U884/U1127/n2 , \U884/U1127/n3 , \U884/U1127/n4 , 
        \c[3] , \c[2] , \c[1] , \c[0] , dsela, dsel, csel, \U884/U1118_0_/nr , 
        nca, \U884/U1118_0_/nd , \U884/U1118_0_/n2 , \U884/U1118_1_/nr , 
        \U884/U1118_1_/nd , \U884/U1118_1_/n2 , \U884/U1118_2_/nr , 
        \U884/U1118_2_/nd , \U884/U1118_2_/n2 , \U884/U1118_3_/nr , 
        \U884/U1118_3_/nd , \U884/U1118_3_/n2 , \U884/U1117_0_/nr , nda, 
        \U884/U1117_0_/nd , \U884/U1117_0_/n2 , \U884/U1117_1_/nr , 
        \U884/U1117_1_/nd , \U884/U1117_1_/n2 , \U884/U1117_2_/nr , 
        \U884/U1117_2_/nd , \U884/U1117_2_/n2 , \U884/U1117_3_/nr , 
        \U884/U1117_3_/nd , \U884/U1117_3_/n2 , \U888/s , \U888/r , 
        \U888/nback , \U888/naack , \U888/reset , \U887/s , \U887/r , 
        \U887/nback , \U887/naack , \U887/reset , \U885/s , \U885/r , 
        \U885/nback , \U885/naack , \U885/reset , \U877/x , \U877/reset , 
        \U877/y , \U877/U590/U25/U1/clr , net135, \cl[3] , \cl[1] , 
        \U877/U590/U25/U1/ob , n1, \U877/U589/U25/U1/clr , \cl[0] , 
        \U877/U589/U25/U1/ob , \U877/U588/U25/U1/clr , \cl[2] , 
        \U877/U588/U25/U1/ob , \U877/U591/U25/U1/clr , \U877/U591/U25/U1/ob , 
        \U876/x , \U876/reset , \U876/y , \U876/U590/U25/U1/clr , 
        \U876/U590/U25/U1/ob , \U876/U589/U25/U1/clr , \U876/U589/U25/U1/ob , 
        \U876/U588/U25/U1/clr , \U876/U588/U25/U1/ob , \U876/U591/U25/U1/clr , 
        \U876/U591/U25/U1/ob , \U2/x , \U2/reset , \U2/y , 
        \U2/U590/U25/U1/clr , \U2/U590/U25/U1/ob , \U2/U589/U25/U1/clr , 
        \U2/U589/U25/U1/ob , \U2/U588/U25/U1/clr , \U2/U588/U25/U1/ob , 
        \U2/U591/U25/U1/clr , \U2/U591/U25/U1/ob , \U1/x , \U1/reset , \U1/y , 
        \U1/U590/U25/U1/clr , \U1/U590/U25/U1/ob , \U1/U589/U25/U1/clr , 
        \U1/U589/U25/U1/ob , \U1/U588/U25/U1/clr , \U1/U588/U25/U1/ob , 
        \U1/U591/U25/U1/clr , \U1/U591/U25/U1/ob , \U881/nack[1] , 
        \U881/nack[0] ;
    buf_2 U897 ( .x(nbReset), .a(nReset) );
    and4_1 \U894/U12  ( .x(eop), .a(ncla), .b(csela), .c(asela), .d(i[4]) );
    inv_1 \U891/U1126/U3  ( .x(\U891/reset ), .a(nbReset) );
    inv_1 \U891/U1139/U3  ( .x(\U891/neopack ), .a(eop) );
    nand3_1 \U891/U1131/U9  ( .x(\U891/iay ), .a(\U891/neopack ), .b(
        \U891/naack[0] ), .c(\U891/naack[1] ) );
    nor3_1 \U891/U1128/U27  ( .x(\U891/U1128/nb ), .a(\U891/reset ), .b(\b[3] 
        ), .c(\b[2] ) );
    nor2_1 \U891/U1128/U26  ( .x(\U891/U1128/na ), .a(\b[1] ), .b(\b[0] ) );
    nand2_2 \U891/U1128/U29  ( .x(\U891/ackb ), .a(\U891/U1128/nb ), .b(
        \U891/U1128/na ) );
    nor2_1 \U891/U1133/U5  ( .x(\U891/naack[0] ), .a(\a[3] ), .b(\a[2] ) );
    nor2_1 \U891/U1108/U5  ( .x(\U891/nack ), .a(\U891/acka ), .b(\U891/ackb )
         );
    nor2_1 \U891/U1134/U5  ( .x(\U891/naack[1] ), .a(\a[1] ), .b(\a[0] ) );
    nor2_2 \U891/U914/U6  ( .x(nia), .a(\U891/iay ), .b(\U891/ackb ) );
    nand2_1 \U891/U1130/U5  ( .x(\U891/acka ), .a(\U891/naack[0] ), .b(
        \U891/naack[1] ) );
    ao222_4 \U891/U1121/U1/U1  ( .x(bsela), .a(\U891/nack ), .b(bsel), .c(
        \U891/nack ), .d(bsela), .e(bsel), .f(bsela) );
    ao222_4 \U891/U1120/U1/U1  ( .x(asela), .a(asel), .b(\U891/nack ), .c(asel
        ), .d(asela), .e(\U891/nack ), .f(asela) );
    nor3_1 \U891/U1118_0_/Unr  ( .x(\U891/U1118_0_/nr ), .a(i[0]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_0_/Und  ( .x(\U891/U1118_0_/nd ), .a(i[0]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_0_/U1  ( .x(\U891/U1118_0_/n2 ), .a(\U891/U1118_0_/n2 ), 
        .b(\U891/U1118_0_/nr ), .c(\U891/U1118_0_/nd ) );
    inv_2 \U891/U1118_0_/U3  ( .x(\a[0] ), .a(\U891/U1118_0_/n2 ) );
    nor3_1 \U891/U1118_1_/Unr  ( .x(\U891/U1118_1_/nr ), .a(i[1]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_1_/Und  ( .x(\U891/U1118_1_/nd ), .a(i[1]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_1_/U1  ( .x(\U891/U1118_1_/n2 ), .a(\U891/U1118_1_/n2 ), 
        .b(\U891/U1118_1_/nr ), .c(\U891/U1118_1_/nd ) );
    inv_2 \U891/U1118_1_/U3  ( .x(\a[1] ), .a(\U891/U1118_1_/n2 ) );
    nor3_1 \U891/U1118_2_/Unr  ( .x(\U891/U1118_2_/nr ), .a(i[2]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_2_/Und  ( .x(\U891/U1118_2_/nd ), .a(i[2]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_2_/U1  ( .x(\U891/U1118_2_/n2 ), .a(\U891/U1118_2_/n2 ), 
        .b(\U891/U1118_2_/nr ), .c(\U891/U1118_2_/nd ) );
    inv_2 \U891/U1118_2_/U3  ( .x(\a[2] ), .a(\U891/U1118_2_/n2 ) );
    nor3_1 \U891/U1118_3_/Unr  ( .x(\U891/U1118_3_/nr ), .a(i[3]), .b(asela), 
        .c(naa) );
    nand3_1 \U891/U1118_3_/Und  ( .x(\U891/U1118_3_/nd ), .a(i[3]), .b(asela), 
        .c(naa) );
    oa21_1 \U891/U1118_3_/U1  ( .x(\U891/U1118_3_/n2 ), .a(\U891/U1118_3_/n2 ), 
        .b(\U891/U1118_3_/nr ), .c(\U891/U1118_3_/nd ) );
    inv_2 \U891/U1118_3_/U3  ( .x(\a[3] ), .a(\U891/U1118_3_/n2 ) );
    nor3_1 \U891/U1117_0_/Unr  ( .x(\U891/U1117_0_/nr ), .a(i[0]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_0_/Und  ( .x(\U891/U1117_0_/nd ), .a(i[0]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_0_/U1  ( .x(\U891/U1117_0_/n2 ), .a(\U891/U1117_0_/n2 ), 
        .b(\U891/U1117_0_/nr ), .c(\U891/U1117_0_/nd ) );
    inv_2 \U891/U1117_0_/U3  ( .x(\b[0] ), .a(\U891/U1117_0_/n2 ) );
    nor3_1 \U891/U1117_1_/Unr  ( .x(\U891/U1117_1_/nr ), .a(i[1]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_1_/Und  ( .x(\U891/U1117_1_/nd ), .a(i[1]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_1_/U1  ( .x(\U891/U1117_1_/n2 ), .a(\U891/U1117_1_/n2 ), 
        .b(\U891/U1117_1_/nr ), .c(\U891/U1117_1_/nd ) );
    inv_2 \U891/U1117_1_/U3  ( .x(\b[1] ), .a(\U891/U1117_1_/n2 ) );
    nor3_1 \U891/U1117_2_/Unr  ( .x(\U891/U1117_2_/nr ), .a(i[2]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_2_/Und  ( .x(\U891/U1117_2_/nd ), .a(i[2]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_2_/U1  ( .x(\U891/U1117_2_/n2 ), .a(\U891/U1117_2_/n2 ), 
        .b(\U891/U1117_2_/nr ), .c(\U891/U1117_2_/nd ) );
    inv_2 \U891/U1117_2_/U3  ( .x(\b[2] ), .a(\U891/U1117_2_/n2 ) );
    nor3_1 \U891/U1117_3_/Unr  ( .x(\U891/U1117_3_/nr ), .a(i[3]), .b(bsela), 
        .c(nba) );
    nand3_1 \U891/U1117_3_/Und  ( .x(\U891/U1117_3_/nd ), .a(i[3]), .b(bsela), 
        .c(nba) );
    oa21_1 \U891/U1117_3_/U1  ( .x(\U891/U1117_3_/n2 ), .a(\U891/U1117_3_/n2 ), 
        .b(\U891/U1117_3_/nr ), .c(\U891/U1117_3_/nd ) );
    inv_2 \U891/U1117_3_/U3  ( .x(\b[3] ), .a(\U891/U1117_3_/n2 ) );
    inv_1 \U886/U1126/U3  ( .x(\U886/reset ), .a(nbReset) );
    nor3_1 \U886/U1128/U27  ( .x(\U886/U1128/nb ), .a(\U886/reset ), .b(\f[3] 
        ), .c(\f[2] ) );
    nor2_1 \U886/U1128/U26  ( .x(\U886/U1128/na ), .a(\f[1] ), .b(\f[0] ) );
    nand2_2 \U886/U1128/U29  ( .x(\U886/ackb ), .a(\U886/U1128/nb ), .b(
        \U886/U1128/na ) );
    nor2_1 \U886/U1108/U5  ( .x(\U886/nack ), .a(\U886/acka ), .b(\U886/ackb )
         );
    nor2_2 \U886/U914/U6  ( .x(nba), .a(\U886/acka ), .b(\U886/ackb ) );
    and4_1 \U886/U1127/U25  ( .x(\U886/U1127/n5 ), .a(\U886/U1127/n1 ), .b(
        \U886/U1127/n2 ), .c(\U886/U1127/n3 ), .d(\U886/U1127/n4 ) );
    inv_1 \U886/U1127/U1  ( .x(\U886/U1127/n1 ), .a(\e[3] ) );
    inv_1 \U886/U1127/U2  ( .x(\U886/U1127/n2 ), .a(\e[2] ) );
    inv_1 \U886/U1127/U3  ( .x(\U886/U1127/n3 ), .a(\e[1] ) );
    inv_1 \U886/U1127/U4  ( .x(\U886/U1127/n4 ), .a(\e[0] ) );
    inv_2 \U886/U1127/U5  ( .x(\U886/acka ), .a(\U886/U1127/n5 ) );
    ao222_2 \U886/U1121/U19/U1/U1  ( .x(fsela), .a(\U886/nack ), .b(fsel), .c(
        \U886/nack ), .d(fsela), .e(fsel), .f(fsela) );
    ao222_2 \U886/U1120/U19/U1/U1  ( .x(esela), .a(esel), .b(\U886/nack ), .c(
        esel), .d(esela), .e(\U886/nack ), .f(esela) );
    nor3_1 \U886/U1118_0_/Unr  ( .x(\U886/U1118_0_/nr ), .a(\b[0] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_0_/Und  ( .x(\U886/U1118_0_/nd ), .a(\b[0] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_0_/U1  ( .x(\U886/U1118_0_/n2 ), .a(\U886/U1118_0_/n2 ), 
        .b(\U886/U1118_0_/nr ), .c(\U886/U1118_0_/nd ) );
    inv_2 \U886/U1118_0_/U3  ( .x(\e[0] ), .a(\U886/U1118_0_/n2 ) );
    nor3_1 \U886/U1118_1_/Unr  ( .x(\U886/U1118_1_/nr ), .a(\b[1] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_1_/Und  ( .x(\U886/U1118_1_/nd ), .a(\b[1] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_1_/U1  ( .x(\U886/U1118_1_/n2 ), .a(\U886/U1118_1_/n2 ), 
        .b(\U886/U1118_1_/nr ), .c(\U886/U1118_1_/nd ) );
    inv_2 \U886/U1118_1_/U3  ( .x(\e[1] ), .a(\U886/U1118_1_/n2 ) );
    nor3_1 \U886/U1118_2_/Unr  ( .x(\U886/U1118_2_/nr ), .a(\b[2] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_2_/Und  ( .x(\U886/U1118_2_/nd ), .a(\b[2] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_2_/U1  ( .x(\U886/U1118_2_/n2 ), .a(\U886/U1118_2_/n2 ), 
        .b(\U886/U1118_2_/nr ), .c(\U886/U1118_2_/nd ) );
    inv_2 \U886/U1118_2_/U3  ( .x(\e[2] ), .a(\U886/U1118_2_/n2 ) );
    nor3_1 \U886/U1118_3_/Unr  ( .x(\U886/U1118_3_/nr ), .a(\b[3] ), .b(esela), 
        .c(nea) );
    nand3_1 \U886/U1118_3_/Und  ( .x(\U886/U1118_3_/nd ), .a(\b[3] ), .b(esela
        ), .c(nea) );
    oa21_1 \U886/U1118_3_/U1  ( .x(\U886/U1118_3_/n2 ), .a(\U886/U1118_3_/n2 ), 
        .b(\U886/U1118_3_/nr ), .c(\U886/U1118_3_/nd ) );
    inv_2 \U886/U1118_3_/U3  ( .x(\e[3] ), .a(\U886/U1118_3_/n2 ) );
    nor3_1 \U886/U1117_0_/Unr  ( .x(\U886/U1117_0_/nr ), .a(\b[0] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_0_/Und  ( .x(\U886/U1117_0_/nd ), .a(\b[0] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_0_/U1  ( .x(\U886/U1117_0_/n2 ), .a(\U886/U1117_0_/n2 ), 
        .b(\U886/U1117_0_/nr ), .c(\U886/U1117_0_/nd ) );
    inv_2 \U886/U1117_0_/U3  ( .x(\f[0] ), .a(\U886/U1117_0_/n2 ) );
    nor3_1 \U886/U1117_1_/Unr  ( .x(\U886/U1117_1_/nr ), .a(\b[1] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_1_/Und  ( .x(\U886/U1117_1_/nd ), .a(\b[1] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_1_/U1  ( .x(\U886/U1117_1_/n2 ), .a(\U886/U1117_1_/n2 ), 
        .b(\U886/U1117_1_/nr ), .c(\U886/U1117_1_/nd ) );
    inv_2 \U886/U1117_1_/U3  ( .x(\f[1] ), .a(\U886/U1117_1_/n2 ) );
    nor3_1 \U886/U1117_2_/Unr  ( .x(\U886/U1117_2_/nr ), .a(\b[2] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_2_/Und  ( .x(\U886/U1117_2_/nd ), .a(\b[2] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_2_/U1  ( .x(\U886/U1117_2_/n2 ), .a(\U886/U1117_2_/n2 ), 
        .b(\U886/U1117_2_/nr ), .c(\U886/U1117_2_/nd ) );
    inv_2 \U886/U1117_2_/U3  ( .x(\f[2] ), .a(\U886/U1117_2_/n2 ) );
    nor3_1 \U886/U1117_3_/Unr  ( .x(\U886/U1117_3_/nr ), .a(\b[3] ), .b(fsela), 
        .c(nfa) );
    nand3_1 \U886/U1117_3_/Und  ( .x(\U886/U1117_3_/nd ), .a(\b[3] ), .b(fsela
        ), .c(nfa) );
    oa21_1 \U886/U1117_3_/U1  ( .x(\U886/U1117_3_/n2 ), .a(\U886/U1117_3_/n2 ), 
        .b(\U886/U1117_3_/nr ), .c(\U886/U1117_3_/nd ) );
    inv_2 \U886/U1117_3_/U3  ( .x(\f[3] ), .a(\U886/U1117_3_/n2 ) );
    inv_1 \U884/U1126/U3  ( .x(\U884/reset ), .a(nbReset) );
    nor3_1 \U884/U1128/U27  ( .x(\U884/U1128/nb ), .a(\U884/reset ), .b(\d[3] 
        ), .c(\d[2] ) );
    nor2_1 \U884/U1128/U26  ( .x(\U884/U1128/na ), .a(\d[1] ), .b(\d[0] ) );
    nand2_2 \U884/U1128/U29  ( .x(\U884/ackb ), .a(\U884/U1128/nb ), .b(
        \U884/U1128/na ) );
    nor2_1 \U884/U1108/U5  ( .x(\U884/nack ), .a(\U884/acka ), .b(\U884/ackb )
         );
    nor2_2 \U884/U914/U6  ( .x(naa), .a(\U884/acka ), .b(\U884/ackb ) );
    and4_1 \U884/U1127/U25  ( .x(\U884/U1127/n5 ), .a(\U884/U1127/n1 ), .b(
        \U884/U1127/n2 ), .c(\U884/U1127/n3 ), .d(\U884/U1127/n4 ) );
    inv_1 \U884/U1127/U1  ( .x(\U884/U1127/n1 ), .a(\c[3] ) );
    inv_1 \U884/U1127/U2  ( .x(\U884/U1127/n2 ), .a(\c[2] ) );
    inv_1 \U884/U1127/U3  ( .x(\U884/U1127/n3 ), .a(\c[1] ) );
    inv_1 \U884/U1127/U4  ( .x(\U884/U1127/n4 ), .a(\c[0] ) );
    inv_2 \U884/U1127/U5  ( .x(\U884/acka ), .a(\U884/U1127/n5 ) );
    ao222_2 \U884/U1121/U19/U1/U1  ( .x(dsela), .a(\U884/nack ), .b(dsel), .c(
        \U884/nack ), .d(dsela), .e(dsel), .f(dsela) );
    ao222_2 \U884/U1120/U19/U1/U1  ( .x(csela), .a(csel), .b(\U884/nack ), .c(
        csel), .d(csela), .e(\U884/nack ), .f(csela) );
    nor3_1 \U884/U1118_0_/Unr  ( .x(\U884/U1118_0_/nr ), .a(\a[0] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_0_/Und  ( .x(\U884/U1118_0_/nd ), .a(\a[0] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_0_/U1  ( .x(\U884/U1118_0_/n2 ), .a(\U884/U1118_0_/n2 ), 
        .b(\U884/U1118_0_/nr ), .c(\U884/U1118_0_/nd ) );
    inv_2 \U884/U1118_0_/U3  ( .x(\c[0] ), .a(\U884/U1118_0_/n2 ) );
    nor3_1 \U884/U1118_1_/Unr  ( .x(\U884/U1118_1_/nr ), .a(\a[1] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_1_/Und  ( .x(\U884/U1118_1_/nd ), .a(\a[1] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_1_/U1  ( .x(\U884/U1118_1_/n2 ), .a(\U884/U1118_1_/n2 ), 
        .b(\U884/U1118_1_/nr ), .c(\U884/U1118_1_/nd ) );
    inv_2 \U884/U1118_1_/U3  ( .x(\c[1] ), .a(\U884/U1118_1_/n2 ) );
    nor3_1 \U884/U1118_2_/Unr  ( .x(\U884/U1118_2_/nr ), .a(\a[2] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_2_/Und  ( .x(\U884/U1118_2_/nd ), .a(\a[2] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_2_/U1  ( .x(\U884/U1118_2_/n2 ), .a(\U884/U1118_2_/n2 ), 
        .b(\U884/U1118_2_/nr ), .c(\U884/U1118_2_/nd ) );
    inv_2 \U884/U1118_2_/U3  ( .x(\c[2] ), .a(\U884/U1118_2_/n2 ) );
    nor3_1 \U884/U1118_3_/Unr  ( .x(\U884/U1118_3_/nr ), .a(\a[3] ), .b(csela), 
        .c(nca) );
    nand3_1 \U884/U1118_3_/Und  ( .x(\U884/U1118_3_/nd ), .a(\a[3] ), .b(csela
        ), .c(nca) );
    oa21_1 \U884/U1118_3_/U1  ( .x(\U884/U1118_3_/n2 ), .a(\U884/U1118_3_/n2 ), 
        .b(\U884/U1118_3_/nr ), .c(\U884/U1118_3_/nd ) );
    inv_2 \U884/U1118_3_/U3  ( .x(\c[3] ), .a(\U884/U1118_3_/n2 ) );
    nor3_1 \U884/U1117_0_/Unr  ( .x(\U884/U1117_0_/nr ), .a(\a[0] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_0_/Und  ( .x(\U884/U1117_0_/nd ), .a(\a[0] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_0_/U1  ( .x(\U884/U1117_0_/n2 ), .a(\U884/U1117_0_/n2 ), 
        .b(\U884/U1117_0_/nr ), .c(\U884/U1117_0_/nd ) );
    inv_2 \U884/U1117_0_/U3  ( .x(\d[0] ), .a(\U884/U1117_0_/n2 ) );
    nor3_1 \U884/U1117_1_/Unr  ( .x(\U884/U1117_1_/nr ), .a(\a[1] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_1_/Und  ( .x(\U884/U1117_1_/nd ), .a(\a[1] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_1_/U1  ( .x(\U884/U1117_1_/n2 ), .a(\U884/U1117_1_/n2 ), 
        .b(\U884/U1117_1_/nr ), .c(\U884/U1117_1_/nd ) );
    inv_2 \U884/U1117_1_/U3  ( .x(\d[1] ), .a(\U884/U1117_1_/n2 ) );
    nor3_1 \U884/U1117_2_/Unr  ( .x(\U884/U1117_2_/nr ), .a(\a[2] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_2_/Und  ( .x(\U884/U1117_2_/nd ), .a(\a[2] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_2_/U1  ( .x(\U884/U1117_2_/n2 ), .a(\U884/U1117_2_/n2 ), 
        .b(\U884/U1117_2_/nr ), .c(\U884/U1117_2_/nd ) );
    inv_2 \U884/U1117_2_/U3  ( .x(\d[2] ), .a(\U884/U1117_2_/n2 ) );
    nor3_1 \U884/U1117_3_/Unr  ( .x(\U884/U1117_3_/nr ), .a(\a[3] ), .b(dsela), 
        .c(nda) );
    nand3_1 \U884/U1117_3_/Und  ( .x(\U884/U1117_3_/nd ), .a(\a[3] ), .b(dsela
        ), .c(nda) );
    oa21_1 \U884/U1117_3_/U1  ( .x(\U884/U1117_3_/n2 ), .a(\U884/U1117_3_/n2 ), 
        .b(\U884/U1117_3_/nr ), .c(\U884/U1117_3_/nd ) );
    inv_2 \U884/U1117_3_/U3  ( .x(\d[3] ), .a(\U884/U1117_3_/n2 ) );
    nand2_1 \U888/U1128/U5  ( .x(\U888/s ), .a(\U888/r ), .b(\U888/nback ) );
    nand2_1 \U888/U1103/U5  ( .x(\U888/r ), .a(\U888/naack ), .b(\U888/s ) );
    inv_1 \U888/U1111/U3  ( .x(\U888/reset ), .a(nbReset) );
    inv_1 \U888/U1112/U3  ( .x(\U888/naack ), .a(esela) );
    nor2_1 \U888/U1127/U5  ( .x(\U888/nback ), .a(fsela), .b(\U888/reset ) );
    and2_2 \U888/U1129/U8  ( .x(esel), .a(\U888/nback ), .b(\U888/s ) );
    and2_2 \U888/U1124/U8  ( .x(fsel), .a(\U888/r ), .b(\U888/naack ) );
    nand2_1 \U887/U1128/U5  ( .x(\U887/s ), .a(\U887/r ), .b(\U887/nback ) );
    nand2_1 \U887/U1103/U5  ( .x(\U887/r ), .a(\U887/naack ), .b(\U887/s ) );
    inv_1 \U887/U1111/U3  ( .x(\U887/reset ), .a(nbReset) );
    inv_1 \U887/U1112/U3  ( .x(\U887/naack ), .a(csela) );
    nor2_1 \U887/U1127/U5  ( .x(\U887/nback ), .a(dsela), .b(\U887/reset ) );
    and2_2 \U887/U1129/U8  ( .x(csel), .a(\U887/nback ), .b(\U887/s ) );
    and2_2 \U887/U1124/U8  ( .x(dsel), .a(\U887/r ), .b(\U887/naack ) );
    nand2_1 \U885/U1128/U5  ( .x(\U885/s ), .a(\U885/r ), .b(\U885/nback ) );
    nand2_1 \U885/U1103/U5  ( .x(\U885/r ), .a(\U885/naack ), .b(\U885/s ) );
    inv_1 \U885/U1111/U3  ( .x(\U885/reset ), .a(nbReset) );
    inv_1 \U885/U1112/U3  ( .x(\U885/naack ), .a(asela) );
    nor2_1 \U885/U1127/U5  ( .x(\U885/nback ), .a(bsela), .b(\U885/reset ) );
    and2_2 \U885/U1129/U8  ( .x(asel), .a(\U885/nback ), .b(\U885/s ) );
    and2_2 \U885/U1124/U8  ( .x(bsel), .a(\U885/r ), .b(\U885/naack ) );
    nor3_1 \U877/U594/U7  ( .x(\U877/x ), .a(ol[7]), .b(\U877/reset ), .c(oh
        [7]) );
    nor3_1 \U877/U593/U7  ( .x(\U877/y ), .a(ol[6]), .b(\U877/reset ), .c(oh
        [6]) );
    inv_1 \U877/U604/U3  ( .x(\U877/reset ), .a(nbReset) );
    oa31_1 \U877/U590/U25/U1/Uclr  ( .x(\U877/U590/U25/U1/clr ), .a(net135), 
        .b(\cl[3] ), .c(\cl[1] ), .d(oh[6]) );
    oaoi211_1 \U877/U590/U25/U1/Uaoi  ( .x(\U877/U590/U25/U1/ob ), .a(\cl[3] ), 
        .b(\cl[1] ), .c(n1), .d(\U877/U590/U25/U1/clr ) );
    inv_2 \U877/U590/U25/U1/Ui  ( .x(oh[6]), .a(\U877/U590/U25/U1/ob ) );
    oa31_1 \U877/U589/U25/U1/Uclr  ( .x(\U877/U589/U25/U1/clr ), .a(net135), 
        .b(\cl[1] ), .c(\cl[0] ), .d(ol[7]) );
    oaoi211_1 \U877/U589/U25/U1/Uaoi  ( .x(\U877/U589/U25/U1/ob ), .a(\cl[1] ), 
        .b(\cl[0] ), .c(n1), .d(\U877/U589/U25/U1/clr ) );
    inv_2 \U877/U589/U25/U1/Ui  ( .x(ol[7]), .a(\U877/U589/U25/U1/ob ) );
    oa31_1 \U877/U588/U25/U1/Uclr  ( .x(\U877/U588/U25/U1/clr ), .a(net135), 
        .b(\cl[3] ), .c(\cl[2] ), .d(oh[7]) );
    oaoi211_1 \U877/U588/U25/U1/Uaoi  ( .x(\U877/U588/U25/U1/ob ), .a(\cl[3] ), 
        .b(\cl[2] ), .c(n1), .d(\U877/U588/U25/U1/clr ) );
    inv_2 \U877/U588/U25/U1/Ui  ( .x(oh[7]), .a(\U877/U588/U25/U1/ob ) );
    oa31_1 \U877/U591/U25/U1/Uclr  ( .x(\U877/U591/U25/U1/clr ), .a(net135), 
        .b(\cl[2] ), .c(\cl[0] ), .d(ol[6]) );
    oaoi211_1 \U877/U591/U25/U1/Uaoi  ( .x(\U877/U591/U25/U1/ob ), .a(\cl[2] ), 
        .b(\cl[0] ), .c(n1), .d(\U877/U591/U25/U1/clr ) );
    inv_2 \U877/U591/U25/U1/Ui  ( .x(ol[6]), .a(\U877/U591/U25/U1/ob ) );
    ao222_2 \U877/U592/U19/U1/U1  ( .x(ncla), .a(\U877/x ), .b(\U877/y ), .c(
        \U877/x ), .d(ncla), .e(\U877/y ), .f(ncla) );
    nor3_1 \U876/U594/U7  ( .x(\U876/x ), .a(ol[3]), .b(\U876/reset ), .c(oh
        [3]) );
    nor3_1 \U876/U593/U7  ( .x(\U876/y ), .a(ol[2]), .b(\U876/reset ), .c(oh
        [2]) );
    inv_1 \U876/U604/U3  ( .x(\U876/reset ), .a(nbReset) );
    oa31_1 \U876/U590/U25/U1/Uclr  ( .x(\U876/U590/U25/U1/clr ), .a(net135), 
        .b(\d[3] ), .c(\d[1] ), .d(oh[2]) );
    oaoi211_1 \U876/U590/U25/U1/Uaoi  ( .x(\U876/U590/U25/U1/ob ), .a(\d[3] ), 
        .b(\d[1] ), .c(n1), .d(\U876/U590/U25/U1/clr ) );
    inv_2 \U876/U590/U25/U1/Ui  ( .x(oh[2]), .a(\U876/U590/U25/U1/ob ) );
    oa31_1 \U876/U589/U25/U1/Uclr  ( .x(\U876/U589/U25/U1/clr ), .a(net135), 
        .b(\d[1] ), .c(\d[0] ), .d(ol[3]) );
    oaoi211_1 \U876/U589/U25/U1/Uaoi  ( .x(\U876/U589/U25/U1/ob ), .a(\d[1] ), 
        .b(\d[0] ), .c(n1), .d(\U876/U589/U25/U1/clr ) );
    inv_2 \U876/U589/U25/U1/Ui  ( .x(ol[3]), .a(\U876/U589/U25/U1/ob ) );
    oa31_1 \U876/U588/U25/U1/Uclr  ( .x(\U876/U588/U25/U1/clr ), .a(net135), 
        .b(\d[3] ), .c(\d[2] ), .d(oh[3]) );
    oaoi211_1 \U876/U588/U25/U1/Uaoi  ( .x(\U876/U588/U25/U1/ob ), .a(\d[3] ), 
        .b(\d[2] ), .c(n1), .d(\U876/U588/U25/U1/clr ) );
    inv_2 \U876/U588/U25/U1/Ui  ( .x(oh[3]), .a(\U876/U588/U25/U1/ob ) );
    oa31_1 \U876/U591/U25/U1/Uclr  ( .x(\U876/U591/U25/U1/clr ), .a(net135), 
        .b(\d[2] ), .c(\d[0] ), .d(ol[2]) );
    oaoi211_1 \U876/U591/U25/U1/Uaoi  ( .x(\U876/U591/U25/U1/ob ), .a(\d[2] ), 
        .b(\d[0] ), .c(n1), .d(\U876/U591/U25/U1/clr ) );
    inv_2 \U876/U591/U25/U1/Ui  ( .x(ol[2]), .a(\U876/U591/U25/U1/ob ) );
    ao222_2 \U876/U592/U19/U1/U1  ( .x(nda), .a(\U876/x ), .b(\U876/y ), .c(
        \U876/x ), .d(nda), .e(\U876/y ), .f(nda) );
    nor3_1 \U2/U594/U7  ( .x(\U2/x ), .a(ol[1]), .b(\U2/reset ), .c(oh[1]) );
    nor3_1 \U2/U593/U7  ( .x(\U2/y ), .a(ol[0]), .b(\U2/reset ), .c(oh[0]) );
    inv_1 \U2/U604/U3  ( .x(\U2/reset ), .a(nbReset) );
    oa31_1 \U2/U590/U25/U1/Uclr  ( .x(\U2/U590/U25/U1/clr ), .a(net135), .b(
        \f[3] ), .c(\f[1] ), .d(oh[0]) );
    oaoi211_1 \U2/U590/U25/U1/Uaoi  ( .x(\U2/U590/U25/U1/ob ), .a(\f[3] ), .b(
        \f[1] ), .c(n1), .d(\U2/U590/U25/U1/clr ) );
    inv_2 \U2/U590/U25/U1/Ui  ( .x(oh[0]), .a(\U2/U590/U25/U1/ob ) );
    oa31_1 \U2/U589/U25/U1/Uclr  ( .x(\U2/U589/U25/U1/clr ), .a(net135), .b(
        \f[1] ), .c(\f[0] ), .d(ol[1]) );
    oaoi211_1 \U2/U589/U25/U1/Uaoi  ( .x(\U2/U589/U25/U1/ob ), .a(\f[1] ), .b(
        \f[0] ), .c(n1), .d(\U2/U589/U25/U1/clr ) );
    inv_2 \U2/U589/U25/U1/Ui  ( .x(ol[1]), .a(\U2/U589/U25/U1/ob ) );
    oa31_1 \U2/U588/U25/U1/Uclr  ( .x(\U2/U588/U25/U1/clr ), .a(net135), .b(
        \f[3] ), .c(\f[2] ), .d(oh[1]) );
    oaoi211_1 \U2/U588/U25/U1/Uaoi  ( .x(\U2/U588/U25/U1/ob ), .a(\f[3] ), .b(
        \f[2] ), .c(n1), .d(\U2/U588/U25/U1/clr ) );
    inv_2 \U2/U588/U25/U1/Ui  ( .x(oh[1]), .a(\U2/U588/U25/U1/ob ) );
    oa31_1 \U2/U591/U25/U1/Uclr  ( .x(\U2/U591/U25/U1/clr ), .a(net135), .b(
        \f[2] ), .c(\f[0] ), .d(ol[0]) );
    oaoi211_1 \U2/U591/U25/U1/Uaoi  ( .x(\U2/U591/U25/U1/ob ), .a(\f[2] ), .b(
        \f[0] ), .c(n1), .d(\U2/U591/U25/U1/clr ) );
    inv_2 \U2/U591/U25/U1/Ui  ( .x(ol[0]), .a(\U2/U591/U25/U1/ob ) );
    ao222_2 \U2/U592/U19/U1/U1  ( .x(nfa), .a(\U2/x ), .b(\U2/y ), .c(\U2/x ), 
        .d(nfa), .e(\U2/y ), .f(nfa) );
    nor3_1 \U1/U594/U7  ( .x(\U1/x ), .a(ol[5]), .b(\U1/reset ), .c(oh[5]) );
    nor3_1 \U1/U593/U7  ( .x(\U1/y ), .a(ol[4]), .b(\U1/reset ), .c(oh[4]) );
    inv_1 \U1/U604/U3  ( .x(\U1/reset ), .a(nbReset) );
    oa31_1 \U1/U590/U25/U1/Uclr  ( .x(\U1/U590/U25/U1/clr ), .a(net135), .b(
        \e[3] ), .c(\e[1] ), .d(oh[4]) );
    oaoi211_1 \U1/U590/U25/U1/Uaoi  ( .x(\U1/U590/U25/U1/ob ), .a(\e[3] ), .b(
        \e[1] ), .c(n1), .d(\U1/U590/U25/U1/clr ) );
    inv_2 \U1/U590/U25/U1/Ui  ( .x(oh[4]), .a(\U1/U590/U25/U1/ob ) );
    oa31_1 \U1/U589/U25/U1/Uclr  ( .x(\U1/U589/U25/U1/clr ), .a(net135), .b(
        \e[1] ), .c(\e[0] ), .d(ol[5]) );
    oaoi211_1 \U1/U589/U25/U1/Uaoi  ( .x(\U1/U589/U25/U1/ob ), .a(\e[1] ), .b(
        \e[0] ), .c(n1), .d(\U1/U589/U25/U1/clr ) );
    inv_2 \U1/U589/U25/U1/Ui  ( .x(ol[5]), .a(\U1/U589/U25/U1/ob ) );
    oa31_1 \U1/U588/U25/U1/Uclr  ( .x(\U1/U588/U25/U1/clr ), .a(net135), .b(
        \e[3] ), .c(\e[2] ), .d(oh[5]) );
    oaoi211_1 \U1/U588/U25/U1/Uaoi  ( .x(\U1/U588/U25/U1/ob ), .a(\e[3] ), .b(
        \e[2] ), .c(n1), .d(\U1/U588/U25/U1/clr ) );
    inv_2 \U1/U588/U25/U1/Ui  ( .x(oh[5]), .a(\U1/U588/U25/U1/ob ) );
    oa31_1 \U1/U591/U25/U1/Uclr  ( .x(\U1/U591/U25/U1/clr ), .a(net135), .b(
        \e[2] ), .c(\e[0] ), .d(ol[4]) );
    oaoi211_1 \U1/U591/U25/U1/Uaoi  ( .x(\U1/U591/U25/U1/ob ), .a(\e[2] ), .b(
        \e[0] ), .c(n1), .d(\U1/U591/U25/U1/clr ) );
    inv_2 \U1/U591/U25/U1/Ui  ( .x(ol[4]), .a(\U1/U591/U25/U1/ob ) );
    ao222_2 \U1/U592/U19/U1/U1  ( .x(nea), .a(\U1/x ), .b(\U1/y ), .c(\U1/x ), 
        .d(nea), .e(\U1/y ), .f(nea) );
    and3_4 \U881/U20/U9  ( .x(nca), .a(\U881/nack[1] ), .b(\U881/nack[0] ), 
        .c(nbReset) );
    nor2_1 \U881/U18/U5  ( .x(\U881/nack[0] ), .a(\cl[3] ), .b(\cl[0] ) );
    nor2_1 \U881/U19/U5  ( .x(\U881/nack[1] ), .a(\cl[1] ), .b(\cl[2] ) );
    ao222_2 \U881/U15_0_/U19/U1/U1  ( .x(\cl[0] ), .a(\c[0] ), .b(ncla), .c(
        \c[0] ), .d(\cl[0] ), .e(ncla), .f(\cl[0] ) );
    ao222_2 \U881/U15_1_/U19/U1/U1  ( .x(\cl[1] ), .a(\c[1] ), .b(ncla), .c(
        \c[1] ), .d(\cl[1] ), .e(ncla), .f(\cl[1] ) );
    ao222_2 \U881/U15_2_/U19/U1/U1  ( .x(\cl[2] ), .a(\c[2] ), .b(ncla), .c(
        \c[2] ), .d(\cl[2] ), .e(ncla), .f(\cl[2] ) );
    ao222_2 \U881/U15_3_/U19/U1/U1  ( .x(\cl[3] ), .a(\c[3] ), .b(ncla), .c(
        \c[3] ), .d(\cl[3] ), .e(ncla), .f(\cl[3] ) );
    and2_5 U1 ( .x(n1), .a(nbReset), .b(noa) );
    and2_3 U2 ( .x(net135), .a(nbReset), .b(noa) );
endmodule


module chain_selement_ga_71 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_70 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_t_ctrl_1 ( cack, fcdefer, fcslowack, screq, ack, defer, fcack, 
    nReset, scack, slowack );
input  ack, defer, fcack, nReset, scack, slowack;
output cack, fcdefer, fcslowack, screq;
    wire net269, net280, net275, net270, net268, net266, net274, net273, 
        net267, net264, net272, net271, net263, net277, net265, net278, net276, 
        net279, \U49/U28/U1/clr , \U49/U28/U1/set , \U50/U28/U1/clr , 
        \U50/U28/U1/set , \U51/U28/U1/clr , \U51/U28/U1/set , \U57/acb , 
        \U57/U1/Z ;
    chain_selement_ga_71 U55 ( .Aa(net269), .Br(fcdefer), .Ar(net280), .Ba(
        fcack) );
    chain_selement_ga_70 U54 ( .Aa(net275), .Br(fcslowack), .Ar(net270), .Ba(
        fcack) );
    or2_4 \U12/U12  ( .x(net268), .a(net266), .b(net270) );
    or2_4 \U56/U12  ( .x(net274), .a(net275), .b(net269) );
    or2_4 \U14/U12  ( .x(net273), .a(net274), .b(net266) );
    or3_1 \U36/U12  ( .x(cack), .a(net267), .b(net264), .c(net272) );
    nor3_1 \U21/U7  ( .x(net271), .a(net270), .b(net266), .c(net280) );
    and2_1 \U53/U8  ( .x(net263), .a(net271), .b(nReset) );
    and2_1 \U43/U8  ( .x(net277), .a(net265), .b(nReset) );
    nor2_1 \U22/U5  ( .x(net265), .a(net278), .b(net276) );
    ao222_2 \U44/U19/U1/U1  ( .x(net276), .a(net280), .b(net273), .c(net280), 
        .d(net276), .e(net273), .f(net276) );
    ao222_2 \U40/U19/U1/U1  ( .x(net280), .a(net272), .b(net277), .c(net272), 
        .d(net280), .e(net277), .f(net280) );
    ao222_2 \U45/U19/U1/U1  ( .x(net279), .a(net273), .b(net268), .c(net273), 
        .d(net279), .e(net268), .f(net279) );
    ao222_2 \U42/U19/U1/U1  ( .x(net266), .a(net277), .b(net267), .c(net277), 
        .d(net266), .e(net267), .f(net266) );
    ao222_2 \U39/U19/U1/U1  ( .x(net270), .a(net277), .b(net264), .c(net277), 
        .d(net270), .e(net264), .f(net270) );
    aoai211_1 \U49/U28/U1/U1  ( .x(\U49/U28/U1/clr ), .a(ack), .b(nReset), .c(
        net263), .d(net267) );
    nand3_1 \U49/U28/U1/U2  ( .x(\U49/U28/U1/set ), .a(net263), .b(ack), .c(
        nReset) );
    nand2_2 \U49/U28/U1/U3  ( .x(net267), .a(\U49/U28/U1/clr ), .b(
        \U49/U28/U1/set ) );
    aoai211_1 \U50/U28/U1/U1  ( .x(\U50/U28/U1/clr ), .a(slowack), .b(nReset), 
        .c(net263), .d(net264) );
    nand3_1 \U50/U28/U1/U2  ( .x(\U50/U28/U1/set ), .a(net263), .b(slowack), 
        .c(nReset) );
    nand2_2 \U50/U28/U1/U3  ( .x(net264), .a(\U50/U28/U1/clr ), .b(
        \U50/U28/U1/set ) );
    aoai211_1 \U51/U28/U1/U1  ( .x(\U51/U28/U1/clr ), .a(defer), .b(nReset), 
        .c(net263), .d(net272) );
    nand2_2 \U51/U28/U1/U3  ( .x(net272), .a(\U51/U28/U1/clr ), .b(
        \U51/U28/U1/set ) );
    and2_1 \U57/U2/U8  ( .x(screq), .a(net279), .b(\U57/acb ) );
    nor2_1 \U57/U3/U5  ( .x(net278), .a(\U57/acb ), .b(scack) );
    oai21_1 \U57/U1/U30/U1/U1  ( .x(\U57/acb ), .a(\U57/U1/Z ), .b(scack), .c(
        net279) );
    inv_1 \U57/U1/U30/U1/U2  ( .x(\U57/U1/Z ), .a(\U57/acb ) );
    nand3_0 U1 ( .x(\U51/U28/U1/set ), .a(net263), .b(defer), .c(nReset) );
endmodule


module target_imem ( addr, ccol, chainresponse, crnw, csize, ctag, lock, 
    nchaincommandack, nrouteack, pred, rack, routetxreq, seq, tag_h, tag_l, wd, 
    cack, cdefer, chaincommand, cndefer, cok, err, nReset, nchainresponseack, 
    rd, route, routetxack );
output [63:0] addr;
output [5:0] ccol;
output [4:0] chainresponse;
output [1:0] crnw;
output [3:0] csize;
output [9:0] ctag;
output [1:0] lock;
output [1:0] pred;
output [1:0] seq;
output [4:0] tag_h;
output [4:0] tag_l;
output [63:0] wd;
input  [4:0] chaincommand;
input  [1:0] err;
input  [63:0] rd;
input  [4:0] route;
input  cack, cdefer, cndefer, cok, nReset, nchainresponseack, routetxack;
output nchaincommandack, nrouteack, rack, routetxreq;
    wire read_ctrlack, chainff_ack, read_req, \chainff_l[7] , \chainff_l[6] , 
        \chainff_l[5] , \chainff_l[4] , \chainff_l[3] , \chainff_l[2] , 
        \chainff_l[1] , \chainff_l[0] , \chainff_h[7] , \chainff_h[6] , 
        \chainff_h[5] , \chainff_h[4] , \chainff_h[3] , \chainff_h[2] , 
        \chainff_h[1] , \chainff_h[0] , read_cd, teop, rhdrack, fcack, tcba, 
        net145, n5, screq, fcslowack, fcdefer, read_ack, \rhdr_h[7] , 
        \rhdr_l[7] , \rhdr_l[6] , \rhdr_l[5] , \rhdr_h[6] , \rhdr_h[5] , 
        \rhdr_l[15] , \rhdr_l[14] , \rhdr_l[13] , \rhdr_h[15] , \rhdr_h[14] , 
        \rhdr_h[13] , \tcbl[7] , \tcbl[6] , \tcbl[5] , \tcbl[4] , \tcbl[3] , 
        \tcbl[2] , \tcbl[1] , \tcbl[0] , \tcbh[7] , \tcbh[6] , \tcbh[5] , 
        \tcbh[4] , \tcbh[3] , \tcbh[2] , \tcbh[1] , \tcbh[0] , nbreset, 
        ntresponseack, \tresponse[4] , \tresponse[3] , \tresponse[2] , 
        \tresponse[1] , \tresponse[0] , net200, noba, pullcd, net168, n9, n10, 
        net188, net201, net194, net178, net189, net191, \obl[7] , \obl[6] , 
        \obl[5] , \obl[4] , \obl[3] , \obl[2] , \obl[1] , \obl[0] , \obh[7] , 
        \obh[6] , \obh[5] , \obh[4] , \obh[3] , \obh[2] , \obh[1] , \obh[0] , 
        n11, n12, net284, net265, \chdrack[0] , \U1761/y[0] , \U1761/y[1] , 
        chdrctrlack, hdrcd, \U1761/x[3] , \nchdr_ack[7] , \nchdr_ack[6] , 
        \U1761/U28/Z , \U1761/x[0] , \nchdr_ack[1] , \nchdr_ack[0] , 
        \U1761/U32/Z , \U1761/x[2] , \nchdr_ack[5] , \nchdr_ack[4] , 
        \U1761/U29/Z , \U1761/x[1] , \U1761/U33/Z , \U1761/U30/Z , 
        \nchdr_ack[3] , \nchdr_ack[2] , \U1761/U31/Z , \U1632/Z , \chdrack[1] , 
        \U1676/Z , \U1770/U21/nr , \nchdr_ack[10] , \nchdr_ack[9] , 
        \nchdr_ack[8] , \U1770/U21/nd , \U1770/U21/n2 , \net242[10] , 
        \net244[10] , \net243[10] , \net242[9] , \net244[9] , \net243[9] , 
        \net242[8] , \net244[8] , \net243[8] , \net242[7] , \net244[7] , 
        \net243[7] , \net242[6] , \net244[6] , \net243[6] , \net242[5] , 
        \net244[5] , \net243[5] , \net242[4] , \net244[4] , \net243[4] , 
        \net242[3] , \net244[3] , \net243[3] , \net242[2] , \net244[2] , 
        \net243[2] , \net242[1] , \net244[1] , \net243[1] , \net242[0] , 
        \net244[0] , \net243[0] , \U1574_0_/net231 , n8, n7, \U1574_1_/net231 , 
        n6, \U1574_2_/net231 , \U1574_3_/net231 , \U1574_4_/net231 , 
        \U1574_5_/net231 , \U1574_6_/net231 , \U1574_7_/net231 , 
        \U1574_8_/net231 , \U1574_9_/net231 , \U1574_10_/net231 , net248;
    chain_sendword_1 U1765 ( .ctrlack(read_ctrlack), .oh({\chainff_h[7] , 
        \chainff_h[6] , \chainff_h[5] , \chainff_h[4] , \chainff_h[3] , 
        \chainff_h[2] , \chainff_h[1] , \chainff_h[0] }), .ol({\chainff_l[7] , 
        \chainff_l[6] , \chainff_l[5] , \chainff_l[4] , \chainff_l[3] , 
        \chainff_l[2] , \chainff_l[1] , \chainff_l[0] }), .chainackff(
        chainff_ack), .ctrlreq(read_req), .ih(rd[63:32]), .il(rd[31:0]) );
    chain_dr32bit_completion_9 rd_cd ( .o(read_cd), .i(rd) );
    chain_trhdr_1 xmitHdr ( .chainff_ack(chainff_ack), .chainh({\tcbh[7] , 
        \tcbh[6] , \tcbh[5] , \tcbh[4] , \tcbh[3] , \tcbh[2] , \tcbh[1] , 
        \tcbh[0] }), .chainl({\tcbl[7] , \tcbl[6] , \tcbl[5] , \tcbl[4] , 
        \tcbl[3] , \tcbl[2] , \tcbl[1] , \tcbl[0] }), .eop(teop), .hdrack(
        rhdrack), .normal_ack(rack), .notify_ack(fcack), .read_req(read_req), 
        .routereq(routetxreq), .chain_ff_h({\chainff_h[7] , \chainff_h[6] , 
        \chainff_h[5] , \chainff_h[4] , \chainff_h[3] , \chainff_h[2] , 
        \chainff_h[1] , \chainff_h[0] }), .chainack(tcba), .chainff_l({
        \chainff_l[7] , \chainff_l[6] , \chainff_l[5] , \chainff_l[4] , 
        \chainff_l[3] , \chainff_l[2] , \chainff_l[1] , \chainff_l[0] }), 
        .eopack(net145), .err(err), .nReset(n5), .normal_response(screq), 
        .notify_accept(fcslowack), .notify_defer(fcdefer), .rcol_h({
        \rhdr_h[15] , \rhdr_h[14] , \rhdr_h[13] }), .rcol_l({\rhdr_l[15] , 
        \rhdr_l[14] , \rhdr_l[13] }), .read_ack(read_ack), .rnw_h(\rhdr_h[7] ), 
        .rnw_l(\rhdr_l[7] ), .routeack(routetxack), .rsize_h({\rhdr_h[6] , 
        \rhdr_h[5] }), .rsize_l({\rhdr_l[6] , \rhdr_l[5] }), .rtag_h(tag_h), 
        .rtag_l(tag_l) );
    chain_dr2fr_byte_4 dr2fr ( .eop_ack(net145), .ia(tcba), .o({\tresponse[4] , 
        \tresponse[3] , \tresponse[2] , \tresponse[1] , \tresponse[0] }), 
        .eop(teop), .ih({\tcbh[7] , \tcbh[6] , \tcbh[5] , \tcbh[4] , \tcbh[3] , 
        \tcbh[2] , \tcbh[1] , \tcbh[0] }), .il({\tcbl[7] , \tcbl[6] , 
        \tcbl[5] , \tcbl[4] , \tcbl[3] , \tcbl[2] , \tcbl[1] , \tcbl[0] }), 
        .nReset(nbreset), .noa(ntresponseack) );
    chain_mergepackets_4 merger ( .naa(nrouteack), .nba(ntresponseack), .o(
        chainresponse), .a(route), .b({\tresponse[4] , \tresponse[3] , 
        \tresponse[2] , \tresponse[1] , \tresponse[0] }), .nReset(nbreset), 
        .noa(nchainresponseack) );
    chain_tchdr_1 header ( .addr_req(net200), .col_h(ccol[5:3]), .col_l(ccol
        [2:0]), .itag_h(ctag[9:5]), .itag_l(ctag[4:0]), .lock(lock), .ncback(
        noba), .pred(pred), .pullcd(pullcd), .reset(net168), .rnw_h(n9), 
        .rnw_l(n10), .seq(seq), .size_h(csize[3:2]), .size_l({n11, n12}), 
        .write_req(net188), .chwh({\obh[7] , \obh[6] , \obh[5] , \obh[4] , 
        \obh[3] , \obh[2] , \obh[1] , \obh[0] }), .chwl({\obl[7] , \obl[6] , 
        \obl[5] , \obl[4] , \obl[3] , \obl[2] , \obl[1] , \obl[0] }), 
        .addr_ack(net201), .addr_pull(net194), .nReset(n5), .nack(net178), 
        .write_ack(net189), .write_pull(net191) );
    chain_irdemux_32new_3 wd_hld ( .ctrlack(net189), .oh(wd[63:32]), .ol(wd
        [31:0]), .pullreq(net191), .pull_h({\obh[7] , \obh[6] , \obh[5] , 
        \obh[4] , \obh[3] , \obh[2] , \obh[1] , \obh[0] }), .pull_l({\obl[7] , 
        \obl[6] , \obl[5] , \obl[4] , \obl[3] , \obl[2] , \obl[1] , \obl[0] }), 
        .pullcd(pullcd), .reset(net168), .ctrlreq(net188) );
    chain_irdemux_32new_2 adr_hld ( .ctrlack(net201), .oh(addr[63:32]), .ol(
        addr[31:0]), .pullreq(net194), .pull_h({\obh[7] , \obh[6] , \obh[5] , 
        \obh[4] , \obh[3] , \obh[2] , \obh[1] , \obh[0] }), .pull_l({\obl[7] , 
        \obl[6] , \obl[5] , \obl[4] , \obl[3] , \obl[2] , \obl[1] , \obl[0] }), 
        .pullcd(pullcd), .reset(net168), .ctrlreq(net200) );
    chain_fr2dr_byte_1 chain_decoder ( .nia(nchaincommandack), .oh({\obh[7] , 
        \obh[6] , \obh[5] , \obh[4] , \obh[3] , \obh[2] , \obh[1] , \obh[0] }), 
        .ol({\obl[7] , \obl[6] , \obl[5] , \obl[4] , \obl[3] , \obl[2] , 
        \obl[1] , \obl[0] }), .i(chaincommand), .nReset(nbreset), .noa(noba)
         );
    chain_t_ctrl_1 cmd_ctrl ( .cack(net284), .fcdefer(fcdefer), .fcslowack(
        fcslowack), .screq(screq), .ack(cok), .defer(cdefer), .fcack(fcack), 
        .nReset(n5), .scack(rack), .slowack(cndefer) );
    inv_1 \I4/U3  ( .x(net265), .a(nbreset) );
    ao222_1 \U1761/U37/U18/U1/U1  ( .x(\chdrack[0] ), .a(\U1761/y[0] ), .b(
        \U1761/y[1] ), .c(\U1761/y[0] ), .d(\chdrack[0] ), .e(\U1761/y[1] ), 
        .f(\chdrack[0] ) );
    ao222_1 \U1762/U18/U1/U1  ( .x(chdrctrlack), .a(hdrcd), .b(net284), .c(
        hdrcd), .d(chdrctrlack), .e(net284), .f(chdrctrlack) );
    ao222_1 \U1769/U18/U1/U1  ( .x(read_ack), .a(read_ctrlack), .b(read_cd), 
        .c(read_ctrlack), .d(read_ack), .e(read_cd), .f(read_ack) );
    aoi222_1 \U1761/U28/U30/U1  ( .x(\U1761/x[3] ), .a(\nchdr_ack[7] ), .b(
        \nchdr_ack[6] ), .c(\nchdr_ack[7] ), .d(\U1761/U28/Z ), .e(
        \nchdr_ack[6] ), .f(\U1761/U28/Z ) );
    inv_1 \U1761/U28/U30/Uinv  ( .x(\U1761/U28/Z ), .a(\U1761/x[3] ) );
    aoi222_1 \U1761/U32/U30/U1  ( .x(\U1761/x[0] ), .a(\nchdr_ack[1] ), .b(
        \nchdr_ack[0] ), .c(\nchdr_ack[1] ), .d(\U1761/U32/Z ), .e(
        \nchdr_ack[0] ), .f(\U1761/U32/Z ) );
    inv_1 \U1761/U32/U30/Uinv  ( .x(\U1761/U32/Z ), .a(\U1761/x[0] ) );
    aoi222_1 \U1761/U29/U30/U1  ( .x(\U1761/x[2] ), .a(\nchdr_ack[5] ), .b(
        \nchdr_ack[4] ), .c(\nchdr_ack[5] ), .d(\U1761/U29/Z ), .e(
        \nchdr_ack[4] ), .f(\U1761/U29/Z ) );
    inv_1 \U1761/U29/U30/Uinv  ( .x(\U1761/U29/Z ), .a(\U1761/x[2] ) );
    aoi222_1 \U1761/U33/U30/U1  ( .x(\U1761/y[0] ), .a(\U1761/x[1] ), .b(
        \U1761/x[0] ), .c(\U1761/x[1] ), .d(\U1761/U33/Z ), .e(\U1761/x[0] ), 
        .f(\U1761/U33/Z ) );
    inv_1 \U1761/U33/U30/Uinv  ( .x(\U1761/U33/Z ), .a(\U1761/y[0] ) );
    aoi222_1 \U1761/U30/U30/U1  ( .x(\U1761/y[1] ), .a(\U1761/x[3] ), .b(
        \U1761/x[2] ), .c(\U1761/x[3] ), .d(\U1761/U30/Z ), .e(\U1761/x[2] ), 
        .f(\U1761/U30/Z ) );
    inv_1 \U1761/U30/U30/Uinv  ( .x(\U1761/U30/Z ), .a(\U1761/y[1] ) );
    aoi222_1 \U1761/U31/U30/U1  ( .x(\U1761/x[1] ), .a(\nchdr_ack[3] ), .b(
        \nchdr_ack[2] ), .c(\nchdr_ack[3] ), .d(\U1761/U31/Z ), .e(
        \nchdr_ack[2] ), .f(\U1761/U31/Z ) );
    inv_1 \U1761/U31/U30/Uinv  ( .x(\U1761/U31/Z ), .a(\U1761/x[1] ) );
    aoi222_1 \U1632/U30/U1  ( .x(net178), .a(cack), .b(chdrctrlack), .c(cack), 
        .d(\U1632/Z ), .e(chdrctrlack), .f(\U1632/Z ) );
    inv_1 \U1632/U30/Uinv  ( .x(\U1632/Z ), .a(net178) );
    aoi222_1 \U1676/U30/U1  ( .x(hdrcd), .a(\chdrack[0] ), .b(\chdrack[1] ), 
        .c(\chdrack[0] ), .d(\U1676/Z ), .e(\chdrack[1] ), .f(\U1676/Z ) );
    inv_1 \U1676/U30/Uinv  ( .x(\U1676/Z ), .a(hdrcd) );
    nor3_1 \U1770/U21/Unr  ( .x(\U1770/U21/nr ), .a(\nchdr_ack[10] ), .b(
        \nchdr_ack[9] ), .c(\nchdr_ack[8] ) );
    nand3_1 \U1770/U21/Und  ( .x(\U1770/U21/nd ), .a(\nchdr_ack[10] ), .b(
        \nchdr_ack[9] ), .c(\nchdr_ack[8] ) );
    oa21_1 \U1770/U21/U1  ( .x(\U1770/U21/n2 ), .a(\U1770/U21/n2 ), .b(
        \U1770/U21/nr ), .c(\U1770/U21/nd ) );
    inv_1 \U1770/U21/U3  ( .x(\chdrack[1] ), .a(\U1770/U21/n2 ) );
    nor2_1 \U1652_0_/U2/U5  ( .x(\nchdr_ack[0] ), .a(\net242[10] ), .b(
        \net244[10] ) );
    ao222_2 \U1652_0_/U12/U19/U1/U1  ( .x(\net244[10] ), .a(\net243[10] ), .b(
        csize[0]), .c(\net243[10] ), .d(\net244[10] ), .e(csize[0]), .f(
        \net244[10] ) );
    ao222_2 \U1652_0_/U11/U19/U1/U1  ( .x(\net242[10] ), .a(csize[2]), .b(
        \net243[10] ), .c(csize[2]), .d(\net242[10] ), .e(\net243[10] ), .f(
        \net242[10] ) );
    nor2_1 \U1652_1_/U2/U5  ( .x(\nchdr_ack[1] ), .a(\net242[9] ), .b(
        \net244[9] ) );
    ao222_2 \U1652_1_/U12/U19/U1/U1  ( .x(\net244[9] ), .a(\net243[9] ), .b(
        csize[1]), .c(\net243[9] ), .d(\net244[9] ), .e(csize[1]), .f(
        \net244[9] ) );
    ao222_2 \U1652_1_/U11/U19/U1/U1  ( .x(\net242[9] ), .a(csize[3]), .b(
        \net243[9] ), .c(csize[3]), .d(\net242[9] ), .e(\net243[9] ), .f(
        \net242[9] ) );
    nor2_1 \U1652_2_/U2/U5  ( .x(\nchdr_ack[2] ), .a(\net242[8] ), .b(
        \net244[8] ) );
    ao222_2 \U1652_2_/U12/U19/U1/U1  ( .x(\net244[8] ), .a(\net243[8] ), .b(
        crnw[0]), .c(\net243[8] ), .d(\net244[8] ), .e(crnw[0]), .f(
        \net244[8] ) );
    ao222_2 \U1652_2_/U11/U19/U1/U1  ( .x(\net242[8] ), .a(crnw[1]), .b(
        \net243[8] ), .c(crnw[1]), .d(\net242[8] ), .e(\net243[8] ), .f(
        \net242[8] ) );
    nor2_1 \U1652_3_/U2/U5  ( .x(\nchdr_ack[3] ), .a(\net242[7] ), .b(
        \net244[7] ) );
    ao222_2 \U1652_3_/U12/U19/U1/U1  ( .x(\net244[7] ), .a(\net243[7] ), .b(
        ctag[0]), .c(\net243[7] ), .d(\net244[7] ), .e(ctag[0]), .f(
        \net244[7] ) );
    ao222_2 \U1652_3_/U11/U19/U1/U1  ( .x(\net242[7] ), .a(ctag[5]), .b(
        \net243[7] ), .c(ctag[5]), .d(\net242[7] ), .e(\net243[7] ), .f(
        \net242[7] ) );
    nor2_1 \U1652_4_/U2/U5  ( .x(\nchdr_ack[4] ), .a(\net242[6] ), .b(
        \net244[6] ) );
    ao222_2 \U1652_4_/U12/U19/U1/U1  ( .x(\net244[6] ), .a(\net243[6] ), .b(
        ctag[1]), .c(\net243[6] ), .d(\net244[6] ), .e(ctag[1]), .f(
        \net244[6] ) );
    ao222_2 \U1652_4_/U11/U19/U1/U1  ( .x(\net242[6] ), .a(ctag[6]), .b(
        \net243[6] ), .c(ctag[6]), .d(\net242[6] ), .e(\net243[6] ), .f(
        \net242[6] ) );
    nor2_1 \U1652_5_/U2/U5  ( .x(\nchdr_ack[5] ), .a(\net242[5] ), .b(
        \net244[5] ) );
    ao222_2 \U1652_5_/U12/U19/U1/U1  ( .x(\net244[5] ), .a(\net243[5] ), .b(
        ctag[2]), .c(\net243[5] ), .d(\net244[5] ), .e(ctag[2]), .f(
        \net244[5] ) );
    ao222_2 \U1652_5_/U11/U19/U1/U1  ( .x(\net242[5] ), .a(ctag[7]), .b(
        \net243[5] ), .c(ctag[7]), .d(\net242[5] ), .e(\net243[5] ), .f(
        \net242[5] ) );
    nor2_1 \U1652_6_/U2/U5  ( .x(\nchdr_ack[6] ), .a(\net242[4] ), .b(
        \net244[4] ) );
    ao222_2 \U1652_6_/U12/U19/U1/U1  ( .x(\net244[4] ), .a(\net243[4] ), .b(
        ctag[3]), .c(\net243[4] ), .d(\net244[4] ), .e(ctag[3]), .f(
        \net244[4] ) );
    ao222_2 \U1652_6_/U11/U19/U1/U1  ( .x(\net242[4] ), .a(ctag[8]), .b(
        \net243[4] ), .c(ctag[8]), .d(\net242[4] ), .e(\net243[4] ), .f(
        \net242[4] ) );
    nor2_1 \U1652_7_/U2/U5  ( .x(\nchdr_ack[7] ), .a(\net242[3] ), .b(
        \net244[3] ) );
    ao222_2 \U1652_7_/U12/U19/U1/U1  ( .x(\net244[3] ), .a(\net243[3] ), .b(
        ctag[4]), .c(\net243[3] ), .d(\net244[3] ), .e(ctag[4]), .f(
        \net244[3] ) );
    ao222_2 \U1652_7_/U11/U19/U1/U1  ( .x(\net242[3] ), .a(ctag[9]), .b(
        \net243[3] ), .c(ctag[9]), .d(\net242[3] ), .e(\net243[3] ), .f(
        \net242[3] ) );
    nor2_1 \U1652_8_/U2/U5  ( .x(\nchdr_ack[8] ), .a(\net242[2] ), .b(
        \net244[2] ) );
    ao222_2 \U1652_8_/U12/U19/U1/U1  ( .x(\net244[2] ), .a(\net243[2] ), .b(
        ccol[0]), .c(\net243[2] ), .d(\net244[2] ), .e(ccol[0]), .f(
        \net244[2] ) );
    ao222_2 \U1652_8_/U11/U19/U1/U1  ( .x(\net242[2] ), .a(ccol[3]), .b(
        \net243[2] ), .c(ccol[3]), .d(\net242[2] ), .e(\net243[2] ), .f(
        \net242[2] ) );
    nor2_1 \U1652_9_/U2/U5  ( .x(\nchdr_ack[9] ), .a(\net242[1] ), .b(
        \net244[1] ) );
    ao222_2 \U1652_9_/U12/U19/U1/U1  ( .x(\net244[1] ), .a(\net243[1] ), .b(
        ccol[1]), .c(\net243[1] ), .d(\net244[1] ), .e(ccol[1]), .f(
        \net244[1] ) );
    ao222_2 \U1652_9_/U11/U19/U1/U1  ( .x(\net242[1] ), .a(ccol[4]), .b(
        \net243[1] ), .c(ccol[4]), .d(\net242[1] ), .e(\net243[1] ), .f(
        \net242[1] ) );
    nor2_1 \U1652_10_/U2/U5  ( .x(\nchdr_ack[10] ), .a(\net242[0] ), .b(
        \net244[0] ) );
    ao222_2 \U1652_10_/U12/U19/U1/U1  ( .x(\net244[0] ), .a(\net243[0] ), .b(
        ccol[2]), .c(\net243[0] ), .d(\net244[0] ), .e(ccol[2]), .f(
        \net244[0] ) );
    ao222_2 \U1652_10_/U11/U19/U1/U1  ( .x(\net242[0] ), .a(ccol[5]), .b(
        \net243[0] ), .c(ccol[5]), .d(\net242[0] ), .e(\net243[0] ), .f(
        \net242[0] ) );
    nor2_1 \U1574_0_/U2/U5  ( .x(\U1574_0_/net231 ), .a(\rhdr_l[5] ), .b(
        \rhdr_h[5] ) );
    and2_1 \U1574_0_/U13/U8  ( .x(\net243[10] ), .a(\U1574_0_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_0_/U12/U19/U1/U1  ( .x(\rhdr_h[5] ), .a(n8), .b(
        \net242[10] ), .c(n8), .d(\rhdr_h[5] ), .e(\net242[10] ), .f(
        \rhdr_h[5] ) );
    ao222_2 \U1574_0_/U11/U19/U1/U1  ( .x(\rhdr_l[5] ), .a(\net244[10] ), .b(
        n7), .c(\net244[10] ), .d(\rhdr_l[5] ), .e(n8), .f(\rhdr_l[5] ) );
    nor2_1 \U1574_1_/U2/U5  ( .x(\U1574_1_/net231 ), .a(\rhdr_l[6] ), .b(
        \rhdr_h[6] ) );
    and2_1 \U1574_1_/U13/U8  ( .x(\net243[9] ), .a(\U1574_1_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_1_/U12/U19/U1/U1  ( .x(\rhdr_h[6] ), .a(n7), .b(\net242[9] 
        ), .c(n6), .d(\rhdr_h[6] ), .e(\net242[9] ), .f(\rhdr_h[6] ) );
    ao222_2 \U1574_1_/U11/U19/U1/U1  ( .x(\rhdr_l[6] ), .a(\net244[9] ), .b(n7
        ), .c(\net244[9] ), .d(\rhdr_l[6] ), .e(n8), .f(\rhdr_l[6] ) );
    nor2_1 \U1574_2_/U2/U5  ( .x(\U1574_2_/net231 ), .a(\rhdr_l[7] ), .b(
        \rhdr_h[7] ) );
    and2_1 \U1574_2_/U13/U8  ( .x(\net243[8] ), .a(\U1574_2_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_2_/U12/U19/U1/U1  ( .x(\rhdr_h[7] ), .a(n6), .b(\net242[8] 
        ), .c(n6), .d(\rhdr_h[7] ), .e(\net242[8] ), .f(\rhdr_h[7] ) );
    ao222_2 \U1574_2_/U11/U19/U1/U1  ( .x(\rhdr_l[7] ), .a(\net244[8] ), .b(n7
        ), .c(\net244[8] ), .d(\rhdr_l[7] ), .e(n8), .f(\rhdr_l[7] ) );
    nor2_1 \U1574_3_/U2/U5  ( .x(\U1574_3_/net231 ), .a(tag_l[0]), .b(tag_h[0]
        ) );
    and2_1 \U1574_3_/U13/U8  ( .x(\net243[7] ), .a(\U1574_3_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_3_/U12/U19/U1/U1  ( .x(tag_h[0]), .a(n8), .b(\net242[7] ), 
        .c(n6), .d(tag_h[0]), .e(\net242[7] ), .f(tag_h[0]) );
    ao222_2 \U1574_3_/U11/U19/U1/U1  ( .x(tag_l[0]), .a(\net244[7] ), .b(n7), 
        .c(\net244[7] ), .d(tag_l[0]), .e(n6), .f(tag_l[0]) );
    nor2_1 \U1574_4_/U2/U5  ( .x(\U1574_4_/net231 ), .a(tag_l[1]), .b(tag_h[1]
        ) );
    and2_1 \U1574_4_/U13/U8  ( .x(\net243[6] ), .a(\U1574_4_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_4_/U12/U19/U1/U1  ( .x(tag_h[1]), .a(n6), .b(\net242[6] ), 
        .c(n6), .d(tag_h[1]), .e(\net242[6] ), .f(tag_h[1]) );
    ao222_2 \U1574_4_/U11/U19/U1/U1  ( .x(tag_l[1]), .a(\net244[6] ), .b(n7), 
        .c(\net244[6] ), .d(tag_l[1]), .e(n6), .f(tag_l[1]) );
    nor2_1 \U1574_5_/U2/U5  ( .x(\U1574_5_/net231 ), .a(tag_l[2]), .b(tag_h[2]
        ) );
    and2_1 \U1574_5_/U13/U8  ( .x(\net243[5] ), .a(\U1574_5_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_5_/U12/U19/U1/U1  ( .x(tag_h[2]), .a(n7), .b(\net242[5] ), 
        .c(n6), .d(tag_h[2]), .e(\net242[5] ), .f(tag_h[2]) );
    ao222_2 \U1574_5_/U11/U19/U1/U1  ( .x(tag_l[2]), .a(\net244[5] ), .b(n7), 
        .c(\net244[5] ), .d(tag_l[2]), .e(n8), .f(tag_l[2]) );
    nor2_1 \U1574_6_/U2/U5  ( .x(\U1574_6_/net231 ), .a(tag_l[3]), .b(tag_h[3]
        ) );
    and2_1 \U1574_6_/U13/U8  ( .x(\net243[4] ), .a(\U1574_6_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_6_/U12/U19/U1/U1  ( .x(tag_h[3]), .a(n6), .b(\net242[4] ), 
        .c(n8), .d(tag_h[3]), .e(\net242[4] ), .f(tag_h[3]) );
    ao222_2 \U1574_6_/U11/U19/U1/U1  ( .x(tag_l[3]), .a(\net244[4] ), .b(n7), 
        .c(\net244[4] ), .d(tag_l[3]), .e(n6), .f(tag_l[3]) );
    nor2_1 \U1574_7_/U2/U5  ( .x(\U1574_7_/net231 ), .a(tag_l[4]), .b(tag_h[4]
        ) );
    and2_1 \U1574_7_/U13/U8  ( .x(\net243[3] ), .a(\U1574_7_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_7_/U12/U19/U1/U1  ( .x(tag_h[4]), .a(n6), .b(\net242[3] ), 
        .c(n8), .d(tag_h[4]), .e(\net242[3] ), .f(tag_h[4]) );
    ao222_2 \U1574_7_/U11/U19/U1/U1  ( .x(tag_l[4]), .a(\net244[3] ), .b(n7), 
        .c(\net244[3] ), .d(tag_l[4]), .e(n6), .f(tag_l[4]) );
    nor2_1 \U1574_8_/U2/U5  ( .x(\U1574_8_/net231 ), .a(\rhdr_l[13] ), .b(
        \rhdr_h[13] ) );
    and2_1 \U1574_8_/U13/U8  ( .x(\net243[2] ), .a(\U1574_8_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_8_/U12/U19/U1/U1  ( .x(\rhdr_h[13] ), .a(n7), .b(
        \net242[2] ), .c(n8), .d(\rhdr_h[13] ), .e(\net242[2] ), .f(
        \rhdr_h[13] ) );
    ao222_2 \U1574_8_/U11/U19/U1/U1  ( .x(\rhdr_l[13] ), .a(\net244[2] ), .b(
        n7), .c(\net244[2] ), .d(\rhdr_l[13] ), .e(n6), .f(\rhdr_l[13] ) );
    nor2_1 \U1574_9_/U2/U5  ( .x(\U1574_9_/net231 ), .a(\rhdr_l[14] ), .b(
        \rhdr_h[14] ) );
    and2_1 \U1574_9_/U13/U8  ( .x(\net243[1] ), .a(\U1574_9_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_9_/U12/U19/U1/U1  ( .x(\rhdr_h[14] ), .a(n8), .b(
        \net242[1] ), .c(n6), .d(\rhdr_h[14] ), .e(\net242[1] ), .f(
        \rhdr_h[14] ) );
    ao222_2 \U1574_9_/U11/U19/U1/U1  ( .x(\rhdr_l[14] ), .a(\net244[1] ), .b(
        n7), .c(\net244[1] ), .d(\rhdr_l[14] ), .e(n8), .f(\rhdr_l[14] ) );
    nor2_1 \U1574_10_/U2/U5  ( .x(\U1574_10_/net231 ), .a(\rhdr_l[15] ), .b(
        \rhdr_h[15] ) );
    and2_1 \U1574_10_/U13/U8  ( .x(\net243[0] ), .a(\U1574_10_/net231 ), .b(
        nbreset) );
    ao222_2 \U1574_10_/U12/U19/U1/U1  ( .x(\rhdr_h[15] ), .a(n8), .b(
        \net242[0] ), .c(n8), .d(\rhdr_h[15] ), .e(\net242[0] ), .f(
        \rhdr_h[15] ) );
    ao222_2 \U1574_10_/U11/U19/U1/U1  ( .x(\rhdr_l[15] ), .a(\net244[0] ), .b(
        n7), .c(\net244[0] ), .d(\rhdr_l[15] ), .e(n8), .f(\rhdr_l[15] ) );
    buf_1 U1 ( .x(csize[0]), .a(n12) );
    buf_1 U2 ( .x(csize[1]), .a(n11) );
    buf_1 U3 ( .x(crnw[0]), .a(n10) );
    buf_1 U4 ( .x(crnw[1]), .a(n9) );
    inv_5 U5 ( .x(n5), .a(net265) );
    buf_3 U6 ( .x(nbreset), .a(nReset) );
    buf_3 U7 ( .x(n6), .a(net248) );
    buf_3 U8 ( .x(n8), .a(net248) );
    buf_3 U9 ( .x(n7), .a(net248) );
    nor2_1 U10 ( .x(net248), .a(net265), .b(rhdrack) );
endmodule


module t_adec_imem ( e_h, e_l, r_h, r_l, e_dp, e_ip, e_tic, r_dp, r_ip, r_tic, 
    tag_h, tag_l );
output [2:0] e_h;
output [2:0] e_l;
output [2:0] r_h;
output [2:0] r_l;
input  [2:0] e_dp;
input  [2:0] e_ip;
input  [2:0] e_tic;
input  [2:0] r_dp;
input  [2:0] r_ip;
input  [2:0] r_tic;
input  [4:0] tag_h;
input  [4:0] tag_l;
    wire e_h_1, e_h_0, e_l_2, r_h_1;
    assign e_h[2] = 1'b0;
    assign e_h[1] = e_h_1;
    assign e_h[0] = e_h_0;
    assign e_l[2] = e_l_2;
    assign e_l[1] = e_h_0;
    assign e_l[0] = e_h_1;
    assign r_h[2] = e_h_0;
    assign r_h[1] = r_h_1;
    assign r_h[0] = 1'b0;
    assign r_l[2] = e_h_1;
    assign r_l[0] = e_l_2;
    assign r_h_1 = tag_h[4];
    or2_1 U3 ( .x(r_l[1]), .a(e_h_1), .b(tag_h[3]) );
    buf_3 U6 ( .x(e_h_1), .a(tag_h[2]) );
    or2_2 U7 ( .x(e_l_2), .a(r_h_1), .b(r_l[1]) );
    or2_2 U8 ( .x(e_h_0), .a(tag_h[3]), .b(r_h_1) );
endmodule


module chain_selement_ga_75 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module chain_selement_ga_17 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_symbol_16 ( o, txack, txack_last, e, oa, r, txreq );
output [2:0] o;
input  [1:0] e;
input  [1:0] r;
input  oa, txreq;
output txack, txack_last;
    wire ack, net10, \c[0] , \c[1] ;
    chain_selement_ga_17 U1239 ( .Aa(ack), .Br(net10), .Ar(txreq), .Ba(oa) );
    and2_1 \U1229_0_/U8  ( .x(o[0]), .a(\c[0] ), .b(net10) );
    and2_1 \U1229_1_/U8  ( .x(o[1]), .a(\c[1] ), .b(net10) );
    and2_1 \U1229_2_/U8  ( .x(o[2]), .a(e[1]), .b(net10) );
    ao23_1 \U1251/U19/U21/U1/U1  ( .x(txack_last), .a(ack), .b(txack_last), 
        .c(ack), .d(e[1]), .e(e[1]) );
    ao23_1 \U1250/U19/U21/U1/U1  ( .x(txack), .a(ack), .b(txack), .c(ack), .d(
        e[0]), .e(e[0]) );
    ao222_1 \U1210/U18/U1/U1  ( .x(\c[0] ), .a(e[0]), .b(r[0]), .c(e[0]), .d(
        \c[0] ), .e(r[0]), .f(\c[0] ) );
    ao222_1 \U1209/U18/U1/U1  ( .x(\c[1] ), .a(e[0]), .b(r[1]), .c(e[0]), .d(
        \c[1] ), .e(r[1]), .f(\c[1] ) );
endmodule


module chain_selement_ga_18 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_symbol_17 ( o, txack, txack_last, e, oa, r, txreq );
output [2:0] o;
input  [1:0] e;
input  [1:0] r;
input  oa, txreq;
output txack, txack_last;
    wire ack, net10, \c[0] , \c[1] , n2, n1;
    chain_selement_ga_18 U1239 ( .Aa(ack), .Br(net10), .Ar(txreq), .Ba(oa) );
    and2_1 \U1229_0_/U8  ( .x(o[0]), .a(\c[0] ), .b(net10) );
    and2_1 \U1229_1_/U8  ( .x(o[1]), .a(\c[1] ), .b(net10) );
    and2_1 \U1229_2_/U8  ( .x(o[2]), .a(e[1]), .b(net10) );
    ao23_1 \U1251/U19/U21/U1/U1  ( .x(txack_last), .a(ack), .b(txack_last), 
        .c(ack), .d(e[1]), .e(e[1]) );
    ao23_1 \U1250/U19/U21/U1/U1  ( .x(txack), .a(ack), .b(txack), .c(ack), .d(
        n2), .e(n2) );
    ao222_1 \U1210/U18/U1/U1  ( .x(\c[0] ), .a(n2), .b(r[0]), .c(n2), .d(
        \c[0] ), .e(r[0]), .f(\c[0] ) );
    ao222_1 \U1209/U18/U1/U1  ( .x(\c[1] ), .a(n2), .b(r[1]), .c(n2), .d(
        \c[1] ), .e(r[1]), .f(\c[1] ) );
    inv_0 U1 ( .x(n1), .a(e[0]) );
    inv_2 U2 ( .x(n2), .a(n1) );
endmodule


module chain_selement_ga_16 ( Aa, Br, Ar, Ba );
input  Ar, Ba;
output Aa, Br;
    wire net2, \U12/Z , \U11/Z ;
    and2_2 \U2/U8  ( .x(Br), .a(Ar), .b(net2) );
    oai21_1 \U12/U30/U1/U1  ( .x(net2), .a(\U12/Z ), .b(Ba), .c(Ar) );
    inv_1 \U12/U30/U1/U2  ( .x(\U12/Z ), .a(net2) );
    aoi21_1 \U11/U30/U1/U1  ( .x(Aa), .a(\U11/Z ), .b(Ba), .c(net2) );
    inv_1 \U11/U30/U1/U2  ( .x(\U11/Z ), .a(Aa) );
endmodule


module route_symbol_15 ( o, txack, txack_last, e, oa, r, txreq );
output [2:0] o;
input  [1:0] e;
input  [1:0] r;
input  oa, txreq;
output txack, txack_last;
    wire ack, net10, \c[0] , \c[1] ;
    chain_selement_ga_16 U1239 ( .Aa(ack), .Br(net10), .Ar(txreq), .Ba(oa) );
    and2_1 \U1229_0_/U8  ( .x(o[0]), .a(\c[0] ), .b(net10) );
    and2_1 \U1229_1_/U8  ( .x(o[1]), .a(\c[1] ), .b(net10) );
    and2_1 \U1229_2_/U8  ( .x(o[2]), .a(e[1]), .b(net10) );
    ao23_1 \U1251/U19/U21/U1/U1  ( .x(txack_last), .a(ack), .b(txack_last), 
        .c(ack), .d(e[1]), .e(e[1]) );
    ao23_1 \U1250/U19/U21/U1/U1  ( .x(txack), .a(ack), .b(txack), .c(ack), .d(
        e[0]), .e(e[0]) );
    ao222_1 \U1210/U18/U1/U1  ( .x(\c[0] ), .a(e[0]), .b(r[0]), .c(e[0]), .d(
        \c[0] ), .e(r[0]), .f(\c[0] ) );
    ao222_1 \U1209/U18/U1/U1  ( .x(\c[1] ), .a(e[0]), .b(r[1]), .c(e[0]), .d(
        \c[1] ), .e(r[1]), .f(\c[1] ) );
endmodule


module resp_route_tx_imem ( o, rtxack, e_h, e_l, noa, r_h, r_l, rtxreq );
output [4:0] o;
input  [2:0] e_h;
input  [2:0] e_l;
input  [2:0] r_h;
input  [2:0] r_l;
input  noa, rtxreq;
output rtxack;
    wire \last[0] , eopsym, net87, net66, net84, \last[2] , net77, \r1[2] , 
        \r1[1] , \r1[0] , \last[1] , \r0[2] , \r0[1] , \r0[0] , \last[3] , 
        \r2[2] , \r2[1] , \r2[0] , net106, net103, \net72[1] , \net72[0] , 
        \I8/nb , \I8/na , \I11/n5 , \I11/n1 , \I11/n2 , \I11/n3 , \I11/n4 , 
        net56, \I7_0_/U25/U1/clr , \I7_0_/U25/U1/ob , \I7_1_/U25/U1/clr , 
        \I7_1_/U25/U1/ob ;
    assign o[3] = 1'b0;
    assign o[2] = 1'b0;
    chain_selement_ga_75 I9 ( .Aa(\last[0] ), .Br(eopsym), .Ar(net87), .Ba(
        net66) );
    route_symbol_16 I2 ( .o({\r1[2] , \r1[1] , \r1[0] }), .txack(net84), 
        .txack_last(\last[2] ), .e({e_h[1], e_l[1]}), .oa(net66), .r({r_h[1], 
        r_l[1]}), .txreq(net77) );
    route_symbol_17 I3 ( .o({\r0[2] , \r0[1] , \r0[0] }), .txack(net87), 
        .txack_last(\last[1] ), .e({e_h[0], e_l[0]}), .oa(net66), .r({r_h[0], 
        r_l[0]}), .txreq(net84) );
    route_symbol_15 I1 ( .o({\r2[2] , \r2[1] , \r2[0] }), .txack(net77), 
        .txack_last(\last[3] ), .e({e_h[2], e_l[2]}), .oa(net66), .r({r_h[2], 
        r_l[2]}), .txreq(rtxreq) );
    nor2_1 \I5/U5  ( .x(net106), .a(eopsym), .b(\r2[2] ) );
    nor2_1 \I16/U5  ( .x(net103), .a(\r1[2] ), .b(\r0[2] ) );
    or2_1 \I14_0_/U12  ( .x(\net72[1] ), .a(\r2[0] ), .b(\r1[0] ) );
    or2_1 \I14_1_/U12  ( .x(\net72[0] ), .a(\r2[1] ), .b(\r1[1] ) );
    nor3_1 \I8/U27  ( .x(\I8/nb ), .a(o[4]), .b(1'b0), .c(1'b0) );
    nor2_1 \I8/U26  ( .x(\I8/na ), .a(o[1]), .b(o[0]) );
    nand2_2 \I8/U29  ( .x(net66), .a(\I8/nb ), .b(\I8/na ) );
    and4_1 \I11/U16  ( .x(\I11/n5 ), .a(\I11/n1 ), .b(\I11/n2 ), .c(\I11/n3 ), 
        .d(\I11/n4 ) );
    inv_1 \I11/U1  ( .x(\I11/n1 ), .a(\last[3] ) );
    inv_1 \I11/U2  ( .x(\I11/n2 ), .a(\last[2] ) );
    inv_1 \I11/U3  ( .x(\I11/n3 ), .a(\last[1] ) );
    inv_1 \I11/U4  ( .x(\I11/n4 ), .a(\last[0] ) );
    inv_1 \I11/U5  ( .x(rtxack), .a(\I11/n5 ) );
    nand2_1 \I17/U5  ( .x(net56), .a(net106), .b(net103) );
    ao222_1 \I15/U18/U1/U1  ( .x(o[4]), .a(noa), .b(net56), .c(noa), .d(o[4]), 
        .e(net56), .f(o[4]) );
    oa31_1 \I7_0_/U25/U1/Uclr  ( .x(\I7_0_/U25/U1/clr ), .a(noa), .b(\r0[0] ), 
        .c(\net72[1] ), .d(o[0]) );
    oaoi211_1 \I7_0_/U25/U1/Uaoi  ( .x(\I7_0_/U25/U1/ob ), .a(\r0[0] ), .b(
        \net72[1] ), .c(noa), .d(\I7_0_/U25/U1/clr ) );
    inv_2 \I7_0_/U25/U1/Ui  ( .x(o[0]), .a(\I7_0_/U25/U1/ob ) );
    oa31_1 \I7_1_/U25/U1/Uclr  ( .x(\I7_1_/U25/U1/clr ), .a(noa), .b(\r0[1] ), 
        .c(\net72[0] ), .d(o[1]) );
    oaoi211_1 \I7_1_/U25/U1/Uaoi  ( .x(\I7_1_/U25/U1/ob ), .a(\r0[1] ), .b(
        \net72[0] ), .c(noa), .d(\I7_1_/U25/U1/clr ) );
    inv_2 \I7_1_/U25/U1/Ui  ( .x(o[1]), .a(\I7_1_/U25/U1/ob ) );
endmodule


module sr2dr_word_7 ( i, req, h, l );
input  [31:0] i;
output [31:0] h;
output [31:0] l;
input  req;
    wire \U31/ni , \U31/nh , \U31/nl , n9, n1, n2, \U30/ni , \U30/nh , 
        \U30/nl , n8, \U29/ni , \U29/nh , \U29/nl , \U28/ni , \U28/nh , 
        \U28/nl , \U27/ni , \U27/nh , \U27/nl , \U26/ni , \U26/nh , \U26/nl , 
        n7, n4, \U25/ni , \U25/nh , \U25/nl , \U24/ni , \U24/nh , \U24/nl , 
        \U23/ni , \U23/nh , \U23/nl , n3, \U22/ni , \U22/nh , \U22/nl , n6, 
        \U21/ni , \U21/nh , \U21/nl , \U20/ni , \U20/nh , \U20/nl , n5, 
        \U19/ni , \U19/nh , \U19/nl , \U18/ni , \U18/nh , \U18/nl , \U17/ni , 
        \U17/nh , \U17/nl , \U16/ni , \U16/nh , \U16/nl , \U15/ni , \U15/nh , 
        \U15/nl , \U14/ni , \U14/nh , \U14/nl , \U13/ni , \U13/nh , \U13/nl , 
        \U12/ni , \U12/nh , \U12/nl , \U11/ni , \U11/nh , \U11/nl , \U10/ni , 
        \U10/nh , \U10/nl , \U9/ni , \U9/nh , \U9/nl , \U8/ni , \U8/nh , 
        \U8/nl , \U7/ni , \U7/nh , \U7/nl , \U6/ni , \U6/nh , \U6/nl , \U5/ni , 
        \U5/nh , \U5/nl , \U4/ni , \U4/nh , \U4/nl , \U3/ni , \U3/nh , \U3/nl , 
        \U2/ni , \U2/nh , \U2/nl , \U1/ni , \U1/nh , \U1/nl , \U0/ni , \U0/nh , 
        \U0/nl , n12, n11, n10;
    inv_1 \U31/Uii  ( .x(\U31/ni ), .a(i[31]) );
    inv_1 \U31/Uih  ( .x(\U31/nh ), .a(h[31]) );
    inv_1 \U31/Uil  ( .x(\U31/nl ), .a(l[31]) );
    ao23_1 \U31/Ucl/U1/U1  ( .x(l[31]), .a(n9), .b(l[31]), .c(n1), .d(\U31/ni 
        ), .e(\U31/nh ) );
    ao23_1 \U31/Uch/U1/U1  ( .x(h[31]), .a(n9), .b(h[31]), .c(n2), .d(i[31]), 
        .e(\U31/nl ) );
    inv_1 \U30/Uii  ( .x(\U30/ni ), .a(i[30]) );
    inv_1 \U30/Uih  ( .x(\U30/nh ), .a(h[30]) );
    inv_1 \U30/Uil  ( .x(\U30/nl ), .a(l[30]) );
    ao23_1 \U30/Ucl/U1/U1  ( .x(l[30]), .a(n8), .b(l[30]), .c(n1), .d(\U30/ni 
        ), .e(\U30/nh ) );
    ao23_1 \U30/Uch/U1/U1  ( .x(h[30]), .a(n8), .b(h[30]), .c(n1), .d(i[30]), 
        .e(\U30/nl ) );
    inv_1 \U29/Uii  ( .x(\U29/ni ), .a(i[29]) );
    inv_1 \U29/Uih  ( .x(\U29/nh ), .a(h[29]) );
    inv_1 \U29/Uil  ( .x(\U29/nl ), .a(l[29]) );
    ao23_1 \U29/Ucl/U1/U1  ( .x(l[29]), .a(n8), .b(l[29]), .c(n1), .d(\U29/ni 
        ), .e(\U29/nh ) );
    ao23_1 \U29/Uch/U1/U1  ( .x(h[29]), .a(n8), .b(h[29]), .c(n2), .d(i[29]), 
        .e(\U29/nl ) );
    inv_1 \U28/Uii  ( .x(\U28/ni ), .a(i[28]) );
    inv_1 \U28/Uih  ( .x(\U28/nh ), .a(h[28]) );
    inv_1 \U28/Uil  ( .x(\U28/nl ), .a(l[28]) );
    ao23_1 \U28/Ucl/U1/U1  ( .x(l[28]), .a(n8), .b(l[28]), .c(n2), .d(\U28/ni 
        ), .e(\U28/nh ) );
    ao23_1 \U28/Uch/U1/U1  ( .x(h[28]), .a(n8), .b(h[28]), .c(n2), .d(i[28]), 
        .e(\U28/nl ) );
    inv_1 \U27/Uii  ( .x(\U27/ni ), .a(i[27]) );
    inv_1 \U27/Uih  ( .x(\U27/nh ), .a(h[27]) );
    inv_1 \U27/Uil  ( .x(\U27/nl ), .a(l[27]) );
    ao23_1 \U27/Ucl/U1/U1  ( .x(l[27]), .a(n8), .b(l[27]), .c(n2), .d(\U27/ni 
        ), .e(\U27/nh ) );
    ao23_1 \U27/Uch/U1/U1  ( .x(h[27]), .a(n8), .b(h[27]), .c(n2), .d(i[27]), 
        .e(\U27/nl ) );
    inv_1 \U26/Uii  ( .x(\U26/ni ), .a(i[26]) );
    inv_1 \U26/Uih  ( .x(\U26/nh ), .a(h[26]) );
    inv_1 \U26/Uil  ( .x(\U26/nl ), .a(l[26]) );
    ao23_1 \U26/Ucl/U1/U1  ( .x(l[26]), .a(n7), .b(l[26]), .c(n2), .d(\U26/ni 
        ), .e(\U26/nh ) );
    ao23_1 \U26/Uch/U1/U1  ( .x(h[26]), .a(n7), .b(h[26]), .c(n4), .d(i[26]), 
        .e(\U26/nl ) );
    inv_1 \U25/Uii  ( .x(\U25/ni ), .a(i[25]) );
    inv_1 \U25/Uih  ( .x(\U25/nh ), .a(h[25]) );
    inv_1 \U25/Uil  ( .x(\U25/nl ), .a(l[25]) );
    ao23_1 \U25/Ucl/U1/U1  ( .x(l[25]), .a(n7), .b(l[25]), .c(n4), .d(\U25/ni 
        ), .e(\U25/nh ) );
    ao23_1 \U25/Uch/U1/U1  ( .x(h[25]), .a(n7), .b(h[25]), .c(n4), .d(i[25]), 
        .e(\U25/nl ) );
    inv_1 \U24/Uii  ( .x(\U24/ni ), .a(i[24]) );
    inv_1 \U24/Uih  ( .x(\U24/nh ), .a(h[24]) );
    inv_1 \U24/Uil  ( .x(\U24/nl ), .a(l[24]) );
    ao23_1 \U24/Ucl/U1/U1  ( .x(l[24]), .a(n7), .b(l[24]), .c(n4), .d(\U24/ni 
        ), .e(\U24/nh ) );
    ao23_1 \U24/Uch/U1/U1  ( .x(h[24]), .a(n7), .b(h[24]), .c(n4), .d(i[24]), 
        .e(\U24/nl ) );
    inv_1 \U23/Uii  ( .x(\U23/ni ), .a(i[23]) );
    inv_1 \U23/Uih  ( .x(\U23/nh ), .a(h[23]) );
    inv_1 \U23/Uil  ( .x(\U23/nl ), .a(l[23]) );
    ao23_1 \U23/Ucl/U1/U1  ( .x(l[23]), .a(n7), .b(l[23]), .c(n3), .d(\U23/ni 
        ), .e(\U23/nh ) );
    ao23_1 \U23/Uch/U1/U1  ( .x(h[23]), .a(n7), .b(h[23]), .c(n3), .d(i[23]), 
        .e(\U23/nl ) );
    inv_1 \U22/Uii  ( .x(\U22/ni ), .a(i[22]) );
    inv_1 \U22/Uih  ( .x(\U22/nh ), .a(h[22]) );
    inv_1 \U22/Uil  ( .x(\U22/nl ), .a(l[22]) );
    ao23_1 \U22/Ucl/U1/U1  ( .x(l[22]), .a(n6), .b(l[22]), .c(n3), .d(\U22/ni 
        ), .e(\U22/nh ) );
    ao23_1 \U22/Uch/U1/U1  ( .x(h[22]), .a(n6), .b(h[22]), .c(n3), .d(i[22]), 
        .e(\U22/nl ) );
    inv_1 \U21/Uii  ( .x(\U21/ni ), .a(i[21]) );
    inv_1 \U21/Uih  ( .x(\U21/nh ), .a(h[21]) );
    inv_1 \U21/Uil  ( .x(\U21/nl ), .a(l[21]) );
    ao23_1 \U21/Ucl/U1/U1  ( .x(l[21]), .a(n6), .b(l[21]), .c(n3), .d(\U21/ni 
        ), .e(\U21/nh ) );
    ao23_1 \U21/Uch/U1/U1  ( .x(h[21]), .a(n6), .b(h[21]), .c(n3), .d(i[21]), 
        .e(\U21/nl ) );
    inv_1 \U20/Uii  ( .x(\U20/ni ), .a(i[20]) );
    inv_1 \U20/Uih  ( .x(\U20/nh ), .a(h[20]) );
    inv_1 \U20/Uil  ( .x(\U20/nl ), .a(l[20]) );
    ao23_1 \U20/Ucl/U1/U1  ( .x(l[20]), .a(n6), .b(l[20]), .c(n5), .d(\U20/ni 
        ), .e(\U20/nh ) );
    ao23_1 \U20/Uch/U1/U1  ( .x(h[20]), .a(n6), .b(h[20]), .c(n4), .d(i[20]), 
        .e(\U20/nl ) );
    inv_1 \U19/Uii  ( .x(\U19/ni ), .a(i[19]) );
    inv_1 \U19/Uih  ( .x(\U19/nh ), .a(h[19]) );
    inv_1 \U19/Uil  ( .x(\U19/nl ), .a(l[19]) );
    ao23_1 \U19/Ucl/U1/U1  ( .x(l[19]), .a(n6), .b(l[19]), .c(n4), .d(\U19/ni 
        ), .e(\U19/nh ) );
    ao23_1 \U19/Uch/U1/U1  ( .x(h[19]), .a(n6), .b(h[19]), .c(n4), .d(i[19]), 
        .e(\U19/nl ) );
    inv_1 \U18/Uii  ( .x(\U18/ni ), .a(i[18]) );
    inv_1 \U18/Uih  ( .x(\U18/nh ), .a(h[18]) );
    inv_1 \U18/Uil  ( .x(\U18/nl ), .a(l[18]) );
    ao23_1 \U18/Ucl/U1/U1  ( .x(l[18]), .a(n5), .b(l[18]), .c(n5), .d(\U18/ni 
        ), .e(\U18/nh ) );
    ao23_1 \U18/Uch/U1/U1  ( .x(h[18]), .a(n5), .b(h[18]), .c(n5), .d(i[18]), 
        .e(\U18/nl ) );
    inv_1 \U17/Uii  ( .x(\U17/ni ), .a(i[17]) );
    inv_1 \U17/Uih  ( .x(\U17/nh ), .a(h[17]) );
    inv_1 \U17/Uil  ( .x(\U17/nl ), .a(l[17]) );
    ao23_1 \U17/Ucl/U1/U1  ( .x(l[17]), .a(n6), .b(l[17]), .c(n5), .d(\U17/ni 
        ), .e(\U17/nh ) );
    ao23_1 \U17/Uch/U1/U1  ( .x(h[17]), .a(n7), .b(h[17]), .c(n4), .d(i[17]), 
        .e(\U17/nl ) );
    inv_1 \U16/Uii  ( .x(\U16/ni ), .a(i[16]) );
    inv_1 \U16/Uih  ( .x(\U16/nh ), .a(h[16]) );
    inv_1 \U16/Uil  ( .x(\U16/nl ), .a(l[16]) );
    ao23_1 \U16/Ucl/U1/U1  ( .x(l[16]), .a(n9), .b(l[16]), .c(n3), .d(\U16/ni 
        ), .e(\U16/nh ) );
    ao23_1 \U16/Uch/U1/U1  ( .x(h[16]), .a(n9), .b(h[16]), .c(n1), .d(i[16]), 
        .e(\U16/nl ) );
    inv_1 \U15/Uii  ( .x(\U15/ni ), .a(i[15]) );
    inv_1 \U15/Uih  ( .x(\U15/nh ), .a(h[15]) );
    inv_1 \U15/Uil  ( .x(\U15/nl ), .a(l[15]) );
    ao23_1 \U15/Ucl/U1/U1  ( .x(l[15]), .a(n8), .b(l[15]), .c(n1), .d(\U15/ni 
        ), .e(\U15/nh ) );
    ao23_1 \U15/Uch/U1/U1  ( .x(h[15]), .a(n7), .b(h[15]), .c(n1), .d(i[15]), 
        .e(\U15/nl ) );
    inv_1 \U14/Uii  ( .x(\U14/ni ), .a(i[14]) );
    inv_1 \U14/Uih  ( .x(\U14/nh ), .a(h[14]) );
    inv_1 \U14/Uil  ( .x(\U14/nl ), .a(l[14]) );
    ao23_1 \U14/Ucl/U1/U1  ( .x(l[14]), .a(n6), .b(l[14]), .c(n1), .d(\U14/ni 
        ), .e(\U14/nh ) );
    ao23_1 \U14/Uch/U1/U1  ( .x(h[14]), .a(n6), .b(h[14]), .c(n3), .d(i[14]), 
        .e(\U14/nl ) );
    inv_1 \U13/Uii  ( .x(\U13/ni ), .a(i[13]) );
    inv_1 \U13/Uih  ( .x(\U13/nh ), .a(h[13]) );
    inv_1 \U13/Uil  ( .x(\U13/nl ), .a(l[13]) );
    ao23_1 \U13/Ucl/U1/U1  ( .x(l[13]), .a(n6), .b(l[13]), .c(n4), .d(\U13/ni 
        ), .e(\U13/nh ) );
    ao23_1 \U13/Uch/U1/U1  ( .x(h[13]), .a(n6), .b(h[13]), .c(n4), .d(i[13]), 
        .e(\U13/nl ) );
    inv_1 \U12/Uii  ( .x(\U12/ni ), .a(i[12]) );
    inv_1 \U12/Uih  ( .x(\U12/nh ), .a(h[12]) );
    inv_1 \U12/Uil  ( .x(\U12/nl ), .a(l[12]) );
    ao23_1 \U12/Ucl/U1/U1  ( .x(l[12]), .a(n5), .b(l[12]), .c(n4), .d(\U12/ni 
        ), .e(\U12/nh ) );
    ao23_1 \U12/Uch/U1/U1  ( .x(h[12]), .a(n5), .b(h[12]), .c(n4), .d(i[12]), 
        .e(\U12/nl ) );
    inv_1 \U11/Uii  ( .x(\U11/ni ), .a(i[11]) );
    inv_1 \U11/Uih  ( .x(\U11/nh ), .a(h[11]) );
    inv_1 \U11/Uil  ( .x(\U11/nl ), .a(l[11]) );
    ao23_1 \U11/Ucl/U1/U1  ( .x(l[11]), .a(n5), .b(l[11]), .c(n4), .d(\U11/ni 
        ), .e(\U11/nh ) );
    ao23_1 \U11/Uch/U1/U1  ( .x(h[11]), .a(n5), .b(h[11]), .c(n4), .d(i[11]), 
        .e(\U11/nl ) );
    inv_1 \U10/Uii  ( .x(\U10/ni ), .a(i[10]) );
    inv_1 \U10/Uih  ( .x(\U10/nh ), .a(h[10]) );
    inv_1 \U10/Uil  ( .x(\U10/nl ), .a(l[10]) );
    ao23_1 \U10/Ucl/U1/U1  ( .x(l[10]), .a(n5), .b(l[10]), .c(n3), .d(\U10/ni 
        ), .e(\U10/nh ) );
    ao23_1 \U10/Uch/U1/U1  ( .x(h[10]), .a(n5), .b(h[10]), .c(n3), .d(i[10]), 
        .e(\U10/nl ) );
    inv_1 \U9/Uii  ( .x(\U9/ni ), .a(i[9]) );
    inv_1 \U9/Uih  ( .x(\U9/nh ), .a(h[9]) );
    inv_1 \U9/Uil  ( .x(\U9/nl ), .a(l[9]) );
    ao23_1 \U9/Ucl/U1/U1  ( .x(l[9]), .a(n5), .b(l[9]), .c(n3), .d(\U9/ni ), 
        .e(\U9/nh ) );
    ao23_1 \U9/Uch/U1/U1  ( .x(h[9]), .a(n5), .b(h[9]), .c(n3), .d(i[9]), .e(
        \U9/nl ) );
    inv_1 \U8/Uii  ( .x(\U8/ni ), .a(i[8]) );
    inv_1 \U8/Uih  ( .x(\U8/nh ), .a(h[8]) );
    inv_1 \U8/Uil  ( .x(\U8/nl ), .a(l[8]) );
    ao23_1 \U8/Ucl/U1/U1  ( .x(l[8]), .a(n5), .b(l[8]), .c(n3), .d(\U8/ni ), 
        .e(\U8/nh ) );
    ao23_1 \U8/Uch/U1/U1  ( .x(h[8]), .a(n5), .b(h[8]), .c(n3), .d(i[8]), .e(
        \U8/nl ) );
    inv_1 \U7/Uii  ( .x(\U7/ni ), .a(i[7]) );
    inv_1 \U7/Uih  ( .x(\U7/nh ), .a(h[7]) );
    inv_1 \U7/Uil  ( .x(\U7/nl ), .a(l[7]) );
    ao23_1 \U7/Ucl/U1/U1  ( .x(l[7]), .a(n7), .b(l[7]), .c(n3), .d(\U7/ni ), 
        .e(\U7/nh ) );
    ao23_1 \U7/Uch/U1/U1  ( .x(h[7]), .a(n7), .b(h[7]), .c(n2), .d(i[7]), .e(
        \U7/nl ) );
    inv_1 \U6/Uii  ( .x(\U6/ni ), .a(i[6]) );
    inv_1 \U6/Uih  ( .x(\U6/nh ), .a(h[6]) );
    inv_1 \U6/Uil  ( .x(\U6/nl ), .a(l[6]) );
    ao23_1 \U6/Ucl/U1/U1  ( .x(l[6]), .a(n7), .b(l[6]), .c(n2), .d(\U6/ni ), 
        .e(\U6/nh ) );
    ao23_1 \U6/Uch/U1/U1  ( .x(h[6]), .a(n7), .b(h[6]), .c(n2), .d(i[6]), .e(
        \U6/nl ) );
    inv_1 \U5/Uii  ( .x(\U5/ni ), .a(i[5]) );
    inv_1 \U5/Uih  ( .x(\U5/nh ), .a(h[5]) );
    inv_1 \U5/Uil  ( .x(\U5/nl ), .a(l[5]) );
    ao23_1 \U5/Ucl/U1/U1  ( .x(l[5]), .a(n7), .b(l[5]), .c(n2), .d(\U5/ni ), 
        .e(\U5/nh ) );
    ao23_1 \U5/Uch/U1/U1  ( .x(h[5]), .a(n7), .b(h[5]), .c(n2), .d(i[5]), .e(
        \U5/nl ) );
    inv_1 \U4/Uii  ( .x(\U4/ni ), .a(i[4]) );
    inv_1 \U4/Uih  ( .x(\U4/nh ), .a(h[4]) );
    inv_1 \U4/Uil  ( .x(\U4/nl ), .a(l[4]) );
    ao23_1 \U4/Ucl/U1/U1  ( .x(l[4]), .a(n6), .b(l[4]), .c(n2), .d(\U4/ni ), 
        .e(\U4/nh ) );
    ao23_1 \U4/Uch/U1/U1  ( .x(h[4]), .a(n6), .b(h[4]), .c(n2), .d(i[4]), .e(
        \U4/nl ) );
    inv_1 \U3/Uii  ( .x(\U3/ni ), .a(i[3]) );
    inv_1 \U3/Uih  ( .x(\U3/nh ), .a(h[3]) );
    inv_1 \U3/Uil  ( .x(\U3/nl ), .a(l[3]) );
    ao23_1 \U3/Ucl/U1/U1  ( .x(l[3]), .a(n6), .b(l[3]), .c(n2), .d(\U3/ni ), 
        .e(\U3/nh ) );
    ao23_1 \U3/Uch/U1/U1  ( .x(h[3]), .a(n8), .b(h[3]), .c(n1), .d(i[3]), .e(
        \U3/nl ) );
    inv_1 \U2/Uii  ( .x(\U2/ni ), .a(i[2]) );
    inv_1 \U2/Uih  ( .x(\U2/nh ), .a(h[2]) );
    inv_1 \U2/Uil  ( .x(\U2/nl ), .a(l[2]) );
    ao23_1 \U2/Ucl/U1/U1  ( .x(l[2]), .a(n8), .b(l[2]), .c(n1), .d(\U2/ni ), 
        .e(\U2/nh ) );
    ao23_1 \U2/Uch/U1/U1  ( .x(h[2]), .a(n8), .b(h[2]), .c(n1), .d(i[2]), .e(
        \U2/nl ) );
    inv_1 \U1/Uii  ( .x(\U1/ni ), .a(i[1]) );
    inv_1 \U1/Uih  ( .x(\U1/nh ), .a(h[1]) );
    inv_1 \U1/Uil  ( .x(\U1/nl ), .a(l[1]) );
    ao23_1 \U1/Ucl/U1/U1  ( .x(l[1]), .a(n8), .b(l[1]), .c(n1), .d(\U1/ni ), 
        .e(\U1/nh ) );
    ao23_1 \U1/Uch/U1/U1  ( .x(h[1]), .a(n8), .b(h[1]), .c(n1), .d(i[1]), .e(
        \U1/nl ) );
    inv_1 \U0/Uii  ( .x(\U0/ni ), .a(i[0]) );
    inv_1 \U0/Uih  ( .x(\U0/nh ), .a(h[0]) );
    inv_1 \U0/Uil  ( .x(\U0/nl ), .a(l[0]) );
    ao23_1 \U0/Ucl/U1/U1  ( .x(l[0]), .a(n8), .b(l[0]), .c(n1), .d(\U0/ni ), 
        .e(\U0/nh ) );
    ao23_1 \U0/Uch/U1/U1  ( .x(h[0]), .a(n8), .b(h[0]), .c(n1), .d(i[0]), .e(
        \U0/nl ) );
    buf_16 U1 ( .x(n1), .a(n12) );
    buf_16 U2 ( .x(n2), .a(n12) );
    buf_16 U3 ( .x(n3), .a(n12) );
    buf_16 U4 ( .x(n4), .a(n11) );
    buf_16 U5 ( .x(n5), .a(n11) );
    buf_16 U6 ( .x(n6), .a(n11) );
    buf_16 U7 ( .x(n7), .a(n10) );
    buf_16 U8 ( .x(n8), .a(n10) );
    buf_16 U9 ( .x(n9), .a(n10) );
    buf_16 U10 ( .x(n10), .a(req) );
    buf_16 U11 ( .x(n11), .a(req) );
    buf_16 U12 ( .x(n12), .a(req) );
endmodule


module matched_delay_cp2slave_resp_imem ( x, a );
input  a;
output x;
    buf_1 I1 ( .x(x), .a(a) );
endmodule


module matched_delay_cp2slave_comimem ( x, a );
input  a;
output x;
    buf_1 I1 ( .x(x), .a(a) );
endmodule


module cp2slave_imem ( tc_seq, tc_size, tc_itag, tc_wd, tc_lock, tc_a, tc_rnw, 
    tc_ok, tc_defer, tc_slow, tc_ack, req_in, ts_i, st_i, we_i, mult_i, adr_i, 
    dat_i, seq_i, prd_i, sel_i, ack_in, tr_rd, tr_err, tr_size, tr_ack, tr_rnw, 
    req_out, dat_o, err_o, rty_o, acc_o, sel_o, mult_o, rt_o, ack_out, reset
     );
input  [1:0] tc_seq;
input  [3:0] tc_size;
input  [9:0] tc_itag;
input  [63:0] tc_wd;
input  [1:0] tc_lock;
input  [63:0] tc_a;
input  [1:0] tc_rnw;
output [2:0] ts_i;
output [4:0] st_i;
output [31:0] adr_i;
output [31:0] dat_i;
output [3:0] sel_i;
output [63:0] tr_rd;
output [1:0] tr_err;
output [3:0] tr_size;
output [1:0] tr_rnw;
input  [31:0] dat_o;
input  [3:0] sel_o;
input  [4:0] rt_o;
input  ack_in, tr_ack, req_out, err_o, rty_o, acc_o, mult_o, reset;
output tc_ok, tc_defer, tc_slow, tc_ack, req_in, we_i, mult_i, seq_i, prd_i, 
    ack_out;
    wire tc_wd_63, tc_wd_62, tc_wd_61, tc_wd_60, tc_wd_59, tc_wd_58, tc_wd_56, 
        tc_wd_55, tc_wd_54, tc_wd_53, tc_wd_52, tc_wd_51, tc_wd_50, tc_wd_49, 
        tc_wd_48, tc_wd_47, tc_wd_46, tc_wd_45, tc_wd_44, tc_wd_43, tc_wd_40, 
        tc_wd_39, tc_wd_38, tc_wd_36, tc_wd_32, tc_a_60, tc_a_58, sel_i_3, n2, 
        n334, n311, n129, n309, n310, n315, n348, n349, n350, n456, n336, n457, 
        n345, n303, n505, n193, n476, n479, n229, n226, n257, n263, n260, n268, 
        n269, n270, n265, n266, n267, n277, n252, n248, n249, n250, n245, n246, 
        n247, n242, n243, n244, n222, n223, n224, n220, n234, n235, n236, n231, 
        n232, n233, n205, n206, n207, n203, n199, n200, n201, n197, n218, n214, 
        n215, n216, n211, n212, n213, n208, n209, n210, n374, n375, n368, n251, 
        n280, n274, n271, n427, n196, n424, n202, n240, n237, n413, n219, n421, 
        n418, n416, n428, n425, n422, n414, n411, n408, n238, n272, n351, n366, 
        n335, n355, n531, n532, respond, n313, n121, n122, n359, n360, n123, 
        n337, n124, n125, n126, n127, n217, n128, n312, n130, n1, n284, n285, 
        n449, n282, n283, n380, n279, n276, n397, n454, n463, n453, n395, n404, 
        n383, n443, n477, n455, n230, n135, n305, n487, n302, n445, n446, n442, 
        n136, n320, n400, n137, n340, n198, n386, n381, n478, n475, n407, n402, 
        n204, n221, n141, n321, n483, n484, n485, n480, n474, n227, n188, n517, 
        n525, n180, n401, n387, n394, n481, n482, n491, n195, n492, n369, n181, 
        n429, n415, n324, n343, n363, n319, n344, n354, n304, n330, n497, n496, 
        n291, n438, n373, n367, n439, n440, n333, n308, n297, n347, n301, n503, 
        n499, n502, n498, n288, n327, n316, n298, n294, n358, complb0, n189, 
        n510, n507, n192, n473, n508, n471, n488, n489, n490, complw0, n182, 
        n183, n184, n185, n364, n365, n391, n388, n430, n423, n426, n431, n417, 
        n419, n420, n432, n409, n410, n412, n433, n403, n405, n406, n434, n396, 
        n398, n399, n435, n389, n390, n392, n393, n436, n382, n384, n385, n437, 
        n376, n377, n378, n379, n441, n370, n444, n470, n472, n194, n486, n493, 
        n494, n495, n191, n500, n501, n504, n506, n509, n511, n465, n466, n468, 
        n512, n460, n513, n514, n462, n459, n515, n516, n518, n452, n519, n450, 
        n520, n522, n521, n523, n524, n371, complb1, n190, complw1, n447, n469, 
        n5, n3, n4, n448, n467, n461, n372, n451, n458, n464, n273, n262, n259, 
        n256, n253, n228, n225, n239, n361, n356, n331, n295, n275, n281, n278, 
        n264, n261, n258, n254, n255, n241, n341, n328, n325, n338, n362, n357, 
        n352, n299, n289, n286, n292, n317, n322, n306, n314, n332, n296, n342, 
        n346, n329, n326, n339, n353, n300, n290, n287, n293, n318, n323, n307, 
        req_out_delayed, _25_net_, n529, n530, _24_net_, _26_net_, n142, 
        req_in_i, n186, n187, all_w, all_r, comp_basic, 
        \cg_all_w/__tmp99/loop , comp_wd, \Usze1/ni , \Usze1/nh , \Usze1/nl , 
        n6, \Usze0/ni , \Usze0/nh , \Usze0/nl , \Urnw/ni , \Urnw/nh , 
        \Urnw/nl , \Uerr/ni , \Uerr/nh , \Uerr/nl ;
    assign tc_wd_63 = tc_wd[63];
    assign tc_wd_62 = tc_wd[62];
    assign tc_wd_61 = tc_wd[61];
    assign tc_wd_60 = tc_wd[60];
    assign tc_wd_59 = tc_wd[59];
    assign tc_wd_58 = tc_wd[58];
    assign tc_wd_56 = tc_wd[56];
    assign tc_wd_55 = tc_wd[55];
    assign tc_wd_54 = tc_wd[54];
    assign tc_wd_53 = tc_wd[53];
    assign tc_wd_52 = tc_wd[52];
    assign tc_wd_51 = tc_wd[51];
    assign tc_wd_50 = tc_wd[50];
    assign tc_wd_49 = tc_wd[49];
    assign tc_wd_48 = tc_wd[48];
    assign tc_wd_47 = tc_wd[47];
    assign tc_wd_46 = tc_wd[46];
    assign tc_wd_45 = tc_wd[45];
    assign tc_wd_44 = tc_wd[44];
    assign tc_wd_43 = tc_wd[43];
    assign tc_wd_40 = tc_wd[40];
    assign tc_wd_39 = tc_wd[39];
    assign tc_wd_38 = tc_wd[38];
    assign tc_wd_36 = tc_wd[36];
    assign tc_wd_32 = tc_wd[32];
    assign tc_a_60 = tc_a[60];
    assign tc_a_58 = tc_a[58];
    assign ts_i[2] = 1'b0;
    assign ts_i[1] = 1'b0;
    assign ts_i[0] = 1'b0;
    assign adr_i[28] = tc_a_60;
    assign adr_i[26] = tc_a_58;
    assign dat_i[31] = tc_wd_63;
    assign dat_i[30] = tc_wd_62;
    assign dat_i[29] = tc_wd_61;
    assign dat_i[28] = tc_wd_60;
    assign dat_i[27] = tc_wd_59;
    assign dat_i[26] = tc_wd_58;
    assign dat_i[24] = tc_wd_56;
    assign dat_i[23] = tc_wd_55;
    assign dat_i[22] = tc_wd_54;
    assign dat_i[21] = tc_wd_53;
    assign dat_i[20] = tc_wd_52;
    assign dat_i[19] = tc_wd_51;
    assign dat_i[18] = tc_wd_50;
    assign dat_i[17] = tc_wd_49;
    assign dat_i[16] = tc_wd_48;
    assign dat_i[15] = tc_wd_47;
    assign dat_i[14] = tc_wd_46;
    assign dat_i[13] = tc_wd_45;
    assign dat_i[12] = tc_wd_44;
    assign dat_i[11] = tc_wd_43;
    assign dat_i[8] = tc_wd_40;
    assign dat_i[7] = tc_wd_39;
    assign dat_i[6] = tc_wd_38;
    assign dat_i[4] = tc_wd_36;
    assign dat_i[0] = tc_wd_32;
    assign prd_i = 1'b0;
    assign sel_i[3] = sel_i_3;
    assign sel_i[2] = sel_i_3;
    assign sel_i[0] = 1'b1;
    assign tc_ack = ack_in;
    assign ack_out = tr_ack;
    sr2dr_word_7 Urd ( .i(dat_o), .req(n2), .h(tr_rd[63:32]), .l(tr_rd[31:0])
         );
    inv_1 U3 ( .x(n334), .a(tc_a[7]) );
    inv_1 U5 ( .x(n311), .a(tc_a[21]) );
    and2_1 U6 ( .x(n129), .a(n309), .b(n310) );
    inv_1 U7 ( .x(n309), .a(tc_a[6]) );
    inv_1 U9 ( .x(n315), .a(tc_itag[4]) );
    nand2_1 U10 ( .x(n348), .a(n349), .b(n350) );
    inv_1 U11 ( .x(n349), .a(tc_a[12]) );
    inv_1 U12 ( .x(n456), .a(n348) );
    inv_1 U13 ( .x(n336), .a(tc_a[30]) );
    inv_1 U14 ( .x(n457), .a(n345) );
    inv_1 U15 ( .x(n303), .a(tc_a[8]) );
    nand3_1 U16 ( .x(n505), .a(n193), .b(n476), .c(n479) );
    inv_1 U17 ( .x(n229), .a(tc_wd[5]) );
    inv_1 U18 ( .x(n226), .a(tc_wd[3]) );
    inv_1 U19 ( .x(n257), .a(tc_wd[16]) );
    inv_1 U20 ( .x(n263), .a(tc_wd[21]) );
    inv_1 U21 ( .x(n260), .a(tc_wd[19]) );
    nand2_1 U22 ( .x(n268), .a(n269), .b(n270) );
    inv_1 U23 ( .x(n269), .a(tc_wd[23]) );
    inv_1 U24 ( .x(n270), .a(tc_wd_55) );
    nand2_1 U25 ( .x(n265), .a(n266), .b(n267) );
    inv_1 U26 ( .x(n266), .a(tc_wd[20]) );
    inv_1 U27 ( .x(n277), .a(tc_wd[27]) );
    inv_1 U28 ( .x(n252), .a(tc_wd_47) );
    nand2_1 U29 ( .x(n248), .a(n249), .b(n250) );
    inv_1 U30 ( .x(n249), .a(tc_wd[12]) );
    nand2_1 U31 ( .x(n245), .a(n246), .b(n247) );
    inv_1 U32 ( .x(n246), .a(tc_wd[13]) );
    inv_1 U33 ( .x(n247), .a(tc_wd_45) );
    nand2_1 U34 ( .x(n242), .a(n243), .b(n244) );
    inv_1 U35 ( .x(n243), .a(tc_wd[11]) );
    nand2_1 U36 ( .x(n222), .a(n223), .b(n224) );
    inv_1 U37 ( .x(n223), .a(tc_wd[0]) );
    inv_1 U38 ( .x(n220), .a(tc_wd[1]) );
    nand2_1 U39 ( .x(n234), .a(n235), .b(n236) );
    inv_1 U40 ( .x(n235), .a(tc_wd[7]) );
    nand2_1 U41 ( .x(n231), .a(n232), .b(n233) );
    inv_1 U42 ( .x(n232), .a(tc_wd[4]) );
    nand2_1 U43 ( .x(n205), .a(n206), .b(n207) );
    inv_1 U44 ( .x(n206), .a(tc_wd[18]) );
    inv_1 U45 ( .x(n203), .a(tc_wd[10]) );
    nand2_1 U46 ( .x(n199), .a(n200), .b(n201) );
    inv_1 U47 ( .x(n200), .a(tc_wd[6]) );
    inv_1 U48 ( .x(n197), .a(tc_wd[2]) );
    inv_1 U49 ( .x(n218), .a(tc_wd_46) );
    nand2_1 U50 ( .x(n214), .a(n215), .b(n216) );
    inv_1 U51 ( .x(n215), .a(tc_wd[30]) );
    nand2_1 U52 ( .x(n211), .a(n212), .b(n213) );
    inv_1 U53 ( .x(n213), .a(tc_wd_58) );
    nand2_1 U54 ( .x(n208), .a(n209), .b(n210) );
    inv_1 U55 ( .x(n209), .a(tc_wd[22]) );
    inv_1 U56 ( .x(n374), .a(tc_rnw[0]) );
    inv_1 U57 ( .x(n375), .a(tc_rnw[1]) );
    inv_1 U58 ( .x(n368), .a(tc_a[18]) );
    inv_1 U59 ( .x(n244), .a(tc_wd_43) );
    inv_1 U60 ( .x(n251), .a(tc_wd[15]) );
    inv_1 U61 ( .x(n250), .a(tc_wd_44) );
    inv_1 U62 ( .x(n280), .a(tc_wd[29]) );
    inv_1 U63 ( .x(n267), .a(tc_wd_52) );
    inv_1 U64 ( .x(n274), .a(tc_wd[24]) );
    inv_1 U65 ( .x(n271), .a(tc_wd[25]) );
    inv_1 U66 ( .x(n212), .a(tc_wd[26]) );
    inv_1 U67 ( .x(n210), .a(tc_wd_54) );
    inv_1 U68 ( .x(n216), .a(tc_wd_62) );
    inv_1 U69 ( .x(n201), .a(tc_wd_38) );
    inv_1 U70 ( .x(n427), .a(n196) );
    inv_1 U71 ( .x(n207), .a(tc_wd_50) );
    inv_1 U72 ( .x(n424), .a(n202) );
    inv_1 U73 ( .x(n236), .a(tc_wd_39) );
    inv_1 U74 ( .x(n233), .a(tc_wd_36) );
    inv_1 U75 ( .x(n240), .a(tc_wd[8]) );
    inv_1 U76 ( .x(n237), .a(tc_wd[9]) );
    inv_1 U77 ( .x(n224), .a(tc_wd_32) );
    inv_1 U78 ( .x(n413), .a(n219) );
    nand2_1 U79 ( .x(n421), .a(n418), .b(n416) );
    nand2_1 U80 ( .x(n428), .a(n425), .b(n422) );
    nand2_1 U81 ( .x(n414), .a(n411), .b(n408) );
    inv_1 U82 ( .x(n238), .a(tc_wd[41]) );
    inv_1 U83 ( .x(n272), .a(tc_wd[57]) );
    inv_1 U84 ( .x(n350), .a(tc_a[44]) );
    inv_1 U85 ( .x(n351), .a(tc_a[43]) );
    inv_1 U86 ( .x(n366), .a(tc_a[41]) );
    inv_1 U87 ( .x(n335), .a(tc_a[39]) );
    inv_1 U88 ( .x(n310), .a(tc_a[38]) );
    inv_1 U89 ( .x(n355), .a(tc_a[52]) );
    and3_1 U90 ( .x(tc_ok), .a(n531), .b(n532), .c(respond) );
    and2_1 U91 ( .x(tc_slow), .a(respond), .b(acc_o) );
    inv_1 U94 ( .x(n313), .a(tc_itag[5]) );
    and2_1 U95 ( .x(n121), .a(n334), .b(n335) );
    and2_1 U96 ( .x(n122), .a(n359), .b(n360) );
    and2_1 U97 ( .x(n123), .a(n336), .b(n337) );
    and2_1 U98 ( .x(n124), .a(n237), .b(n238) );
    and2_1 U99 ( .x(n125), .a(n251), .b(n252) );
    and2_1 U100 ( .x(n126), .a(n271), .b(n272) );
    and2_1 U101 ( .x(n127), .a(n217), .b(n218) );
    and2_1 U102 ( .x(n128), .a(n311), .b(n312) );
    nor2_1 U103 ( .x(n130), .a(n1), .b(tc_size[2]) );
    nand2i_1 U105 ( .x(n284), .a(tc_wd[31]), .b(n285) );
    oa22_1 U106 ( .x(n449), .a(tc_a[27]), .b(tc_a[59]), .c(tc_a[54]), .d(tc_a
        [22]) );
    inv_1 U107 ( .x(n359), .a(tc_a[27]) );
    inv_1 U108 ( .x(n360), .a(tc_a[59]) );
    nand2i_1 U109 ( .x(n282), .a(tc_wd[28]), .b(n283) );
    nor2_1 U110 ( .x(n479), .a(tc_itag[0]), .b(tc_itag[5]) );
    nand4_1 U112 ( .x(n380), .a(n279), .b(n276), .c(n284), .d(n282) );
    aoi21_1 U113 ( .x(n425), .a(n200), .b(n201), .c(n427) );
    oa22_1 U114 ( .x(n397), .a(tc_wd[13]), .b(tc_wd_45), .c(tc_wd[11]), .d(
        tc_wd_43) );
    nor2_1 U115 ( .x(n454), .a(tc_a[20]), .b(tc_a[52]) );
    aoi21_1 U116 ( .x(n422), .a(n206), .b(n207), .c(n424) );
    oa22_1 U117 ( .x(n418), .a(tc_wd[26]), .b(tc_wd_58), .c(tc_wd[22]), .d(
        tc_wd_54) );
    oa22_1 U118 ( .x(n416), .a(tc_wd[14]), .b(tc_wd_46), .c(tc_wd[30]), .d(
        tc_wd_62) );
    inv_1 U119 ( .x(n217), .a(tc_wd[14]) );
    aoi22_1 U120 ( .x(n463), .a(n336), .b(n337), .c(n334), .d(n335) );
    nor2_1 U121 ( .x(n453), .a(tc_a[11]), .b(tc_a[43]) );
    oa22_1 U122 ( .x(n395), .a(tc_wd[15]), .b(tc_wd_47), .c(tc_wd[12]), .d(
        tc_wd_44) );
    oa22_1 U123 ( .x(n404), .a(tc_wd[7]), .b(tc_wd_39), .c(tc_wd[4]), .d(
        tc_wd_36) );
    oa22_1 U124 ( .x(n383), .a(tc_wd[23]), .b(tc_wd_55), .c(tc_wd[20]), .d(
        tc_wd_52) );
    aoi21_1 U125 ( .x(n411), .a(n223), .b(n224), .c(n413) );
    nor2_1 U126 ( .x(n443), .a(tc_a[49]), .b(tc_a[17]) );
    aoi22_1 U127 ( .x(n477), .a(n311), .b(n312), .c(n309), .d(n310) );
    oa21_1 U128 ( .x(n455), .a(tc_a[12]), .b(tc_a[44]), .c(n345) );
    inv_1 U129 ( .x(dat_i[5]), .a(n230) );
    inv_1 U130 ( .x(dat_i[9]), .a(n238) );
    inv_1 U131 ( .x(dat_i[25]), .a(n272) );
    buf_1 U132 ( .x(sel_i_3), .a(n1) );
    buf_1 U133 ( .x(adr_i[16]), .a(tc_a[48]) );
    nor2_1 U134 ( .x(n135), .a(tc_a[14]), .b(tc_a[46]) );
    inv_1 U135 ( .x(n305), .a(tc_a[46]) );
    inv_1 U136 ( .x(n487), .a(n302) );
    nand2i_1 U137 ( .x(n445), .a(n446), .b(n442) );
    nor2_1 U138 ( .x(n136), .a(tc_a[29]), .b(tc_a[61]) );
    inv_1 U139 ( .x(n320), .a(tc_a[61]) );
    nand2_1 U140 ( .x(n400), .a(n397), .b(n395) );
    inv_1 U141 ( .x(n137), .a(n340) );
    inv_1 U142 ( .x(dat_i[2]), .a(n198) );
    nand2_1 U143 ( .x(n386), .a(n383), .b(n381) );
    nand3i_1 U144 ( .x(n478), .a(n479), .b(n477), .c(n475) );
    nand2_1 U145 ( .x(n407), .a(n404), .b(n402) );
    inv_1 U146 ( .x(dat_i[10]), .a(n204) );
    inv_1 U147 ( .x(dat_i[1]), .a(n221) );
    nor2_1 U148 ( .x(n141), .a(tc_a[3]), .b(tc_a[35]) );
    inv_1 U149 ( .x(n321), .a(tc_a[35]) );
    nor2_1 U151 ( .x(n483), .a(n484), .b(n485) );
    nor2_1 U152 ( .x(n480), .a(n474), .b(n478) );
    inv_1 U153 ( .x(dat_i[3]), .a(n227) );
    nor2_1 U154 ( .x(n188), .a(n517), .b(n525) );
    nand2_1 U155 ( .x(n180), .a(n401), .b(n387) );
    nor2_1 U156 ( .x(n401), .a(n394), .b(n400) );
    nor2_1 U157 ( .x(n387), .a(n380), .b(n386) );
    nor2_1 U158 ( .x(n481), .a(n482), .b(n135) );
    nor2_1 U159 ( .x(n491), .a(n195), .b(n492) );
    nor2_1 U160 ( .x(n195), .a(tc_size[1]), .b(n1) );
    inv_1 U161 ( .x(adr_i[18]), .a(n369) );
    nand2_1 U162 ( .x(n181), .a(n429), .b(n415) );
    nor2_1 U163 ( .x(n429), .a(n421), .b(n428) );
    nor2_1 U164 ( .x(n415), .a(n407), .b(n414) );
    inv_1 U165 ( .x(adr_i[0]), .a(n324) );
    inv_1 U166 ( .x(n324), .a(tc_a[32]) );
    inv_1 U167 ( .x(sel_i[1]), .a(n130) );
    inv_1 U168 ( .x(st_i[2]), .a(n343) );
    inv_1 U169 ( .x(adr_i[9]), .a(n366) );
    inv_1 U170 ( .x(adr_i[24]), .a(n363) );
    inv_1 U171 ( .x(adr_i[19]), .a(n319) );
    inv_1 U172 ( .x(n319), .a(tc_a[51]) );
    inv_1 U173 ( .x(n369), .a(tc_a[50]) );
    inv_1 U174 ( .x(st_i[3]), .a(n344) );
    inv_1 U175 ( .x(adr_i[13]), .a(n354) );
    inv_1 U176 ( .x(adr_i[12]), .a(n350) );
    inv_1 U177 ( .x(adr_i[8]), .a(n304) );
    inv_1 U178 ( .x(n304), .a(tc_a[40]) );
    inv_1 U179 ( .x(adr_i[2]), .a(n330) );
    buf_1 U180 ( .x(adr_i[17]), .a(tc_a[49]) );
    nand2_1 U181 ( .x(n497), .a(n496), .b(n130) );
    inv_1 U182 ( .x(adr_i[10]), .a(n291) );
    and2_1 U183 ( .x(n438), .a(n373), .b(n367) );
    inv_1 U184 ( .x(n439), .a(n373) );
    inv_1 U185 ( .x(n440), .a(n367) );
    inv_1 U186 ( .x(adr_i[20]), .a(n355) );
    inv_1 U187 ( .x(adr_i[27]), .a(n360) );
    inv_1 U188 ( .x(adr_i[4]), .a(n333) );
    inv_1 U189 ( .x(adr_i[25]), .a(n308) );
    inv_1 U190 ( .x(adr_i[30]), .a(n337) );
    inv_1 U191 ( .x(adr_i[31]), .a(n297) );
    inv_1 U192 ( .x(n297), .a(tc_a[63]) );
    inv_1 U193 ( .x(adr_i[15]), .a(n347) );
    inv_1 U194 ( .x(adr_i[11]), .a(n351) );
    inv_1 U195 ( .x(adr_i[1]), .a(n301) );
    inv_1 U196 ( .x(n301), .a(tc_a[33]) );
    nand2_1 U197 ( .x(n503), .a(n499), .b(n502) );
    nor2_1 U198 ( .x(n499), .a(n497), .b(n498) );
    inv_1 U199 ( .x(adr_i[21]), .a(n312) );
    inv_1 U200 ( .x(n312), .a(tc_a[53]) );
    inv_1 U201 ( .x(seq_i), .a(n288) );
    inv_1 U202 ( .x(adr_i[5]), .a(n327) );
    inv_1 U203 ( .x(st_i[4]), .a(n316) );
    inv_1 U204 ( .x(n316), .a(tc_itag[9]) );
    inv_1 U205 ( .x(st_i[1]), .a(n298) );
    inv_1 U206 ( .x(adr_i[23]), .a(n294) );
    inv_1 U207 ( .x(adr_i[22]), .a(n358) );
    nand2_1 U208 ( .x(complb0), .a(n188), .b(n189) );
    nor2_1 U209 ( .x(n189), .a(n503), .b(n510) );
    inv_1 U210 ( .x(adr_i[29]), .a(n320) );
    inv_1 U211 ( .x(adr_i[7]), .a(n335) );
    inv_1 U212 ( .x(adr_i[14]), .a(n305) );
    inv_1 U213 ( .x(adr_i[6]), .a(n310) );
    inv_1 U214 ( .x(st_i[0]), .a(n313) );
    inv_1 U215 ( .x(adr_i[3]), .a(n321) );
    nand3_1 U218 ( .x(n507), .a(n192), .b(n136), .c(n473) );
    nand2_1 U219 ( .x(n508), .a(n471), .b(n141) );
    nor2_1 U220 ( .x(n488), .a(n489), .b(n490) );
    nand4_1 U222 ( .x(complw0), .a(n182), .b(n183), .c(n184), .d(n185) );
    nor2_1 U223 ( .x(n192), .a(tc_a_58), .b(tc_a[26]) );
    nor2_1 U224 ( .x(n193), .a(tc_a[48]), .b(tc_a[16]) );
    nand2_1 U225 ( .x(n364), .a(n365), .b(n366) );
    nand2_1 U226 ( .x(n394), .a(n391), .b(n388) );
    nand4_1 U227 ( .x(n430), .a(n423), .b(n424), .c(n426), .d(n427) );
    nand4_1 U228 ( .x(n431), .a(n127), .b(n417), .c(n419), .d(n420) );
    nor2_1 U229 ( .x(n185), .a(n430), .b(n431) );
    nand4_1 U230 ( .x(n432), .a(n409), .b(n410), .c(n412), .d(n413) );
    nand4_1 U231 ( .x(n433), .a(n403), .b(n124), .c(n405), .d(n406) );
    nor2_1 U232 ( .x(n184), .a(n432), .b(n433) );
    nand4_1 U233 ( .x(n434), .a(n125), .b(n396), .c(n398), .d(n399) );
    nand4_1 U234 ( .x(n435), .a(n389), .b(n390), .c(n392), .d(n393) );
    nor2_1 U235 ( .x(n183), .a(n434), .b(n435) );
    nand4_1 U236 ( .x(n436), .a(n382), .b(n126), .c(n384), .d(n385) );
    nand4_1 U237 ( .x(n437), .a(n376), .b(n377), .c(n378), .d(n379) );
    nor2_1 U238 ( .x(n182), .a(n436), .b(n437) );
    nand2_1 U239 ( .x(n441), .a(n438), .b(n370) );
    nor2_1 U240 ( .x(n442), .a(n443), .b(n444) );
    nor3_1 U241 ( .x(n470), .a(n471), .b(n136), .c(n141) );
    nor3_1 U242 ( .x(n472), .a(n473), .b(n192), .c(n193) );
    nand2_1 U243 ( .x(n474), .a(n472), .b(n470) );
    nor2_1 U244 ( .x(n475), .a(n476), .b(n194) );
    nand3i_1 U245 ( .x(n486), .a(n487), .b(n481), .c(n483) );
    nand3i_1 U246 ( .x(n493), .a(n494), .b(n488), .c(n491) );
    nor2_1 U247 ( .x(n495), .a(n493), .b(n486) );
    nand2_1 U248 ( .x(n191), .a(n495), .b(n480) );
    nand3_1 U249 ( .x(n498), .a(n489), .b(n492), .c(n490) );
    nand3_1 U250 ( .x(n500), .a(n485), .b(n494), .c(n484) );
    nand2_1 U251 ( .x(n501), .a(n135), .b(n487) );
    nor2_1 U252 ( .x(n502), .a(n500), .b(n501) );
    nand3_1 U253 ( .x(n504), .a(n128), .b(n482), .c(n129) );
    nor2_1 U254 ( .x(n506), .a(n504), .b(n505) );
    nor2_1 U255 ( .x(n509), .a(n507), .b(n508) );
    nand2_1 U256 ( .x(n510), .a(n509), .b(n506) );
    nand3_1 U257 ( .x(n511), .a(n465), .b(n466), .c(n468) );
    nand3_1 U258 ( .x(n512), .a(n123), .b(n121), .c(n460) );
    nor2_1 U259 ( .x(n513), .a(n511), .b(n512) );
    nand3_1 U260 ( .x(n514), .a(n462), .b(n459), .c(n457) );
    nand2_1 U261 ( .x(n515), .a(n453), .b(n456) );
    nor2_1 U262 ( .x(n516), .a(n514), .b(n515) );
    nand2_1 U263 ( .x(n517), .a(n516), .b(n513) );
    nand2_1 U264 ( .x(n518), .a(n454), .b(n452) );
    nor2i_1 U265 ( .x(n519), .a(n450), .b(n518) );
    nand2_1 U266 ( .x(n520), .a(n444), .b(n122) );
    nor2i_1 U267 ( .x(n522), .a(n446), .b(n521) );
    nand2_1 U268 ( .x(n523), .a(n439), .b(n524) );
    inv_1 U270 ( .x(n365), .a(tc_a[9]) );
    inv_1 U271 ( .x(n371), .a(tc_a_60) );
    inv_1 U272 ( .x(n446), .a(n364) );
    nor2_1 U273 ( .x(complb1), .a(n190), .b(n191) );
    nor2_1 U274 ( .x(complw1), .a(n180), .b(n181) );
    nand3i_1 U276 ( .x(n190), .a(n441), .b(n447), .c(n469) );
    and4_1 U277 ( .x(n5), .a(n3), .b(n4), .c(n519), .d(n522) );
    inv_1 U216 ( .x(n3), .a(n520) );
    inv_1 U217 ( .x(n4), .a(n523) );
    inv_1 U428 ( .x(n525), .a(n5) );
    nor2_1 U278 ( .x(n447), .a(n448), .b(n445) );
    nor2_1 U279 ( .x(n469), .a(n467), .b(n461) );
    nand2_1 U280 ( .x(n370), .a(n371), .b(n372) );
    nand3i_1 U281 ( .x(n448), .a(n454), .b(n449), .c(n451) );
    nand3i_1 U282 ( .x(n461), .a(n462), .b(n455), .c(n458) );
    nand3i_1 U283 ( .x(n467), .a(n468), .b(n463), .c(n464) );
    inv_1 U284 ( .x(n382), .a(n273) );
    inv_1 U285 ( .x(n384), .a(n268) );
    inv_1 U286 ( .x(n385), .a(n265) );
    inv_1 U287 ( .x(n376), .a(n284) );
    inv_1 U288 ( .x(n377), .a(n282) );
    inv_1 U289 ( .x(n378), .a(n279) );
    inv_1 U290 ( .x(n379), .a(n276) );
    inv_1 U291 ( .x(n396), .a(n248) );
    inv_1 U292 ( .x(n398), .a(n245) );
    inv_1 U293 ( .x(n399), .a(n242) );
    inv_1 U294 ( .x(n389), .a(n262) );
    inv_1 U295 ( .x(n390), .a(n259) );
    inv_1 U296 ( .x(n392), .a(n256) );
    inv_1 U297 ( .x(n393), .a(n253) );
    inv_1 U298 ( .x(n409), .a(n228) );
    inv_1 U299 ( .x(n410), .a(n225) );
    inv_1 U300 ( .x(n412), .a(n222) );
    inv_1 U301 ( .x(n403), .a(n239) );
    inv_1 U302 ( .x(n405), .a(n234) );
    inv_1 U303 ( .x(n406), .a(n231) );
    inv_1 U304 ( .x(n423), .a(n205) );
    inv_1 U305 ( .x(n426), .a(n199) );
    inv_1 U306 ( .x(n417), .a(n214) );
    inv_1 U307 ( .x(n419), .a(n211) );
    inv_1 U308 ( .x(n420), .a(n208) );
    inv_1 U309 ( .x(n444), .a(n361) );
    inv_1 U310 ( .x(n524), .a(n370) );
    inv_1 U311 ( .x(n450), .a(n356) );
    nand2_1 U312 ( .x(n521), .a(n443), .b(n440) );
    inv_1 U313 ( .x(n372), .a(tc_a[28]) );
    nor2_1 U314 ( .x(n451), .a(n452), .b(n453) );
    nor2_1 U315 ( .x(n458), .a(n459), .b(n460) );
    inv_1 U316 ( .x(n468), .a(n331) );
    nor2_1 U317 ( .x(n464), .a(n465), .b(n466) );
    inv_1 U318 ( .x(n494), .a(n295) );
    nand2_1 U319 ( .x(n273), .a(n274), .b(n275) );
    nand2_1 U320 ( .x(n279), .a(n280), .b(n281) );
    nand2_1 U321 ( .x(n276), .a(n277), .b(n278) );
    nand2_1 U322 ( .x(n262), .a(n263), .b(n264) );
    nand2_1 U323 ( .x(n259), .a(n260), .b(n261) );
    nand2_1 U324 ( .x(n256), .a(n257), .b(n258) );
    nand2_1 U325 ( .x(n253), .a(n254), .b(n255) );
    nand2_1 U326 ( .x(n228), .a(n229), .b(n230) );
    nand2_1 U327 ( .x(n225), .a(n226), .b(n227) );
    nand2_1 U328 ( .x(n219), .a(n220), .b(n221) );
    nand2_1 U329 ( .x(n239), .a(n240), .b(n241) );
    nand2_1 U330 ( .x(n202), .a(n203), .b(n204) );
    nand2_1 U331 ( .x(n196), .a(n197), .b(n198) );
    nor2_1 U332 ( .x(n391), .a(n392), .b(n393) );
    nor2_1 U333 ( .x(n388), .a(n389), .b(n390) );
    nor2_1 U334 ( .x(n381), .a(n382), .b(n126) );
    nor2_1 U335 ( .x(n402), .a(n403), .b(n124) );
    nor2_1 U336 ( .x(n408), .a(n409), .b(n410) );
    inv_1 U337 ( .x(n459), .a(n341) );
    inv_1 U338 ( .x(n465), .a(n328) );
    inv_1 U339 ( .x(n466), .a(n325) );
    inv_1 U340 ( .x(n460), .a(n338) );
    nand2_1 U341 ( .x(n361), .a(n362), .b(n363) );
    nand2_1 U342 ( .x(n373), .a(n374), .b(n375) );
    nand2_1 U343 ( .x(n356), .a(n358), .b(n357) );
    inv_1 U344 ( .x(n452), .a(n352) );
    inv_1 U345 ( .x(n484), .a(n299) );
    inv_1 U346 ( .x(n489), .a(n289) );
    inv_1 U347 ( .x(n492), .a(n286) );
    inv_1 U348 ( .x(n490), .a(n292) );
    inv_1 U349 ( .x(n473), .a(n317) );
    inv_1 U350 ( .x(n471), .a(n322) );
    inv_1 U351 ( .x(n482), .a(n306) );
    inv_1 U352 ( .x(n476), .a(n314) );
    nand2_1 U353 ( .x(n367), .a(n368), .b(n369) );
    nand2_1 U354 ( .x(n331), .a(n332), .b(n333) );
    nand2_1 U355 ( .x(n302), .a(n303), .b(n304) );
    nand2_1 U356 ( .x(n295), .a(n296), .b(n297) );
    inv_1 U357 ( .x(n275), .a(tc_wd_56) );
    inv_1 U358 ( .x(n285), .a(tc_wd_63) );
    inv_1 U359 ( .x(n283), .a(tc_wd_60) );
    inv_1 U360 ( .x(n281), .a(tc_wd_61) );
    inv_1 U361 ( .x(n278), .a(tc_wd_59) );
    inv_1 U362 ( .x(n264), .a(tc_wd_53) );
    inv_1 U363 ( .x(n261), .a(tc_wd_51) );
    inv_1 U364 ( .x(n258), .a(tc_wd_48) );
    inv_1 U365 ( .x(n254), .a(tc_wd[17]) );
    inv_1 U366 ( .x(n255), .a(tc_wd_49) );
    inv_1 U367 ( .x(n230), .a(tc_wd[37]) );
    inv_1 U368 ( .x(n227), .a(tc_wd[35]) );
    inv_1 U369 ( .x(n221), .a(tc_wd[33]) );
    inv_1 U370 ( .x(n241), .a(tc_wd_40) );
    inv_1 U371 ( .x(n204), .a(tc_wd[42]) );
    inv_1 U372 ( .x(n198), .a(tc_wd[34]) );
    nand2_1 U373 ( .x(n341), .a(n342), .b(n343) );
    nand2_1 U374 ( .x(n345), .a(n347), .b(n346) );
    nand2_1 U375 ( .x(n328), .a(n329), .b(n330) );
    nand2_1 U376 ( .x(n325), .a(n326), .b(n327) );
    nand2_1 U377 ( .x(n338), .a(n340), .b(n339) );
    inv_1 U378 ( .x(n362), .a(tc_a[24]) );
    inv_1 U379 ( .x(n363), .a(tc_a[56]) );
    inv_1 U380 ( .x(n357), .a(tc_a[22]) );
    inv_1 U381 ( .x(n358), .a(tc_a[54]) );
    nand2_1 U382 ( .x(n352), .a(n353), .b(n354) );
    nand2_1 U383 ( .x(n299), .a(n300), .b(n301) );
    nand2_1 U384 ( .x(n289), .a(n290), .b(n291) );
    nand2_1 U385 ( .x(n286), .a(n287), .b(n288) );
    nand2_1 U386 ( .x(n292), .a(n293), .b(n294) );
    nand2_1 U387 ( .x(n317), .a(n318), .b(n319) );
    nand2_1 U388 ( .x(n322), .a(n323), .b(n324) );
    nand2_1 U389 ( .x(n306), .a(n307), .b(n308) );
    nand2_1 U390 ( .x(n314), .a(n315), .b(n316) );
    inv_1 U391 ( .x(n332), .a(tc_a[4]) );
    inv_1 U392 ( .x(n333), .a(tc_a[36]) );
    inv_1 U393 ( .x(n296), .a(tc_a[31]) );
    inv_1 U394 ( .x(n342), .a(tc_itag[2]) );
    inv_1 U395 ( .x(n343), .a(tc_itag[7]) );
    inv_1 U396 ( .x(n346), .a(tc_a[15]) );
    inv_1 U397 ( .x(n347), .a(tc_a[47]) );
    inv_1 U398 ( .x(n329), .a(tc_a[2]) );
    inv_1 U399 ( .x(n330), .a(tc_a[34]) );
    inv_1 U400 ( .x(n326), .a(tc_a[5]) );
    inv_1 U401 ( .x(n327), .a(tc_a[37]) );
    inv_1 U402 ( .x(n337), .a(tc_a[62]) );
    inv_1 U403 ( .x(n339), .a(tc_lock[0]) );
    inv_1 U404 ( .x(n340), .a(tc_lock[1]) );
    inv_1 U405 ( .x(n353), .a(tc_a[13]) );
    inv_1 U406 ( .x(n354), .a(tc_a[45]) );
    inv_1 U407 ( .x(n300), .a(tc_a[1]) );
    inv_1 U408 ( .x(n290), .a(tc_a[10]) );
    inv_1 U409 ( .x(n291), .a(tc_a[42]) );
    inv_1 U410 ( .x(n287), .a(tc_seq[0]) );
    inv_1 U411 ( .x(n288), .a(tc_seq[1]) );
    inv_1 U412 ( .x(n293), .a(tc_a[23]) );
    inv_1 U413 ( .x(n294), .a(tc_a[55]) );
    inv_1 U414 ( .x(n318), .a(tc_a[19]) );
    inv_1 U415 ( .x(n323), .a(tc_a[0]) );
    inv_1 U416 ( .x(n307), .a(tc_a[25]) );
    inv_1 U417 ( .x(n308), .a(tc_a[57]) );
    buf_1 U418 ( .x(we_i), .a(tc_rnw[0]) );
    matched_delay_cp2slave_resp_imem U419 ( .x(req_out_delayed), .a(req_out)
         );
    and4_1 U420 ( .x(_25_net_), .a(sel_o[0]), .b(sel_o[1]), .c(n529), .d(n530)
         );
    inv_1 U421 ( .x(_24_net_), .a(we_i) );
    and2_1 U422 ( .x(tc_defer), .a(rty_o), .b(respond) );
    and4_1 U423 ( .x(_26_net_), .a(sel_o[0]), .b(sel_o[1]), .c(sel_o[3]), .d(
        sel_o[2]) );
    inv_1 U424 ( .x(n532), .a(acc_o) );
    inv_1 U425 ( .x(n531), .a(rty_o) );
    inv_1 U426 ( .x(n529), .a(sel_o[2]) );
    inv_1 U427 ( .x(n530), .a(sel_o[3]) );
    buf_1 U150 ( .x(n142), .a(req_in_i) );
    matched_delay_cp2slave_comimem matchDelCom ( .x(req_in), .a(req_in_i) );
    nand2_1 U275 ( .x(req_in_i), .a(n186), .b(n187) );
    inv_1 U221 ( .x(n186), .a(all_w) );
    inv_1 U269 ( .x(n187), .a(all_r) );
    dffp_1 mult_i_reg ( .q(mult_i), .d(n137), .ck(n142) );
    ao222_1 \cg_respond/__tmp99/U1  ( .x(respond), .a(req_out), .b(tc_ack), 
        .c(req_out), .d(respond), .e(tc_ack), .f(respond) );
    oa21_1 \cg_all_r/__tmp99/U1  ( .x(all_r), .a(tc_rnw[1]), .b(all_r), .c(
        comp_basic) );
    ao31_1 \cg_all_w/__tmp99/aoi  ( .x(\cg_all_w/__tmp99/loop ), .a(comp_basic
        ), .b(comp_wd), .c(we_i), .d(all_w) );
    oa21_1 \cg_all_w/__tmp99/outGate  ( .x(all_w), .a(comp_basic), .b(comp_wd), 
        .c(\cg_all_w/__tmp99/loop ) );
    ao222_1 \cg_wd/__tmp99/U1  ( .x(comp_wd), .a(complw0), .b(complw1), .c(
        complw0), .d(comp_wd), .e(complw1), .f(comp_wd) );
    ao222_1 \cg_basic/__tmp99/U1  ( .x(comp_basic), .a(complb0), .b(complb1), 
        .c(complb0), .d(comp_basic), .e(complb1), .f(comp_basic) );
    inv_1 \Usze1/Uii  ( .x(\Usze1/ni ), .a(_26_net_) );
    inv_1 \Usze1/Uih  ( .x(\Usze1/nh ), .a(tr_size[3]) );
    inv_1 \Usze1/Uil  ( .x(\Usze1/nl ), .a(tr_size[1]) );
    ao23_1 \Usze1/Ucl/U1/U1  ( .x(tr_size[1]), .a(n6), .b(tr_size[1]), .c(n2), 
        .d(\Usze1/ni ), .e(\Usze1/nh ) );
    ao23_1 \Usze1/Uch/U1/U1  ( .x(tr_size[3]), .a(n2), .b(tr_size[3]), .c(n2), 
        .d(_26_net_), .e(\Usze1/nl ) );
    inv_1 \Usze0/Uii  ( .x(\Usze0/ni ), .a(_25_net_) );
    inv_1 \Usze0/Uih  ( .x(\Usze0/nh ), .a(tr_size[2]) );
    inv_1 \Usze0/Uil  ( .x(\Usze0/nl ), .a(tr_size[0]) );
    ao23_1 \Usze0/Ucl/U1/U1  ( .x(tr_size[0]), .a(n6), .b(tr_size[0]), .c(n2), 
        .d(\Usze0/ni ), .e(\Usze0/nh ) );
    ao23_1 \Usze0/Uch/U1/U1  ( .x(tr_size[2]), .a(n6), .b(tr_size[2]), .c(n2), 
        .d(_25_net_), .e(\Usze0/nl ) );
    inv_1 \Urnw/Uii  ( .x(\Urnw/ni ), .a(_24_net_) );
    inv_1 \Urnw/Uih  ( .x(\Urnw/nh ), .a(tr_rnw[1]) );
    inv_1 \Urnw/Uil  ( .x(\Urnw/nl ), .a(tr_rnw[0]) );
    ao23_1 \Urnw/Ucl/U1/U1  ( .x(tr_rnw[0]), .a(n2), .b(tr_rnw[0]), .c(n2), 
        .d(\Urnw/ni ), .e(\Urnw/nh ) );
    ao23_1 \Urnw/Uch/U1/U1  ( .x(tr_rnw[1]), .a(n2), .b(tr_rnw[1]), .c(n2), 
        .d(_24_net_), .e(\Urnw/nl ) );
    inv_1 \Uerr/Uii  ( .x(\Uerr/ni ), .a(err_o) );
    inv_1 \Uerr/Uih  ( .x(\Uerr/nh ), .a(tr_err[1]) );
    inv_1 \Uerr/Uil  ( .x(\Uerr/nl ), .a(tr_err[0]) );
    ao23_1 \Uerr/Ucl/U1/U1  ( .x(tr_err[0]), .a(n2), .b(tr_err[0]), .c(n2), 
        .d(\Uerr/ni ), .e(\Uerr/nh ) );
    ao23_1 \Uerr/Uch/U1/U1  ( .x(tr_err[1]), .a(n2), .b(tr_err[1]), .c(n2), 
        .d(err_o), .e(\Uerr/nl ) );
    inv_0 U1 ( .x(n344), .a(tc_itag[8]) );
    nor2_0 U2 ( .x(n462), .a(tc_itag[3]), .b(tc_itag[8]) );
    inv_0 U4 ( .x(n298), .a(tc_itag[6]) );
    nor2_0 U8 ( .x(n485), .a(tc_itag[1]), .b(tc_itag[6]) );
    nor2_0 U92 ( .x(n496), .a(tc_size[0]), .b(tc_size[1]) );
    nor2_0 U93 ( .x(n194), .a(tc_size[0]), .b(tc_size[2]) );
    buf_1 U104 ( .x(n1), .a(tc_size[3]) );
    buf_16 U111 ( .x(n2), .a(req_out_delayed) );
    buf_16 U429 ( .x(n6), .a(req_out_delayed) );
endmodule


module slave_if_imem ( nReset, sc_req, sc_we, sc_mult, sc_seq, sc_prd, sc_ts, 
    sc_st, sc_sel, sc_adr, sc_dat, sc_ack, sr_req, sr_err, sr_rty, sr_acc, 
    sr_mult, sr_ts, sr_rt, sr_sel, sr_dat, sr_ack, chaincommand, 
    nchaincommandack, chainresponse, nchainresponseack, e_dp, e_ip, e_tic, 
    r_dp, r_ip, r_tic );
output [2:0] sc_ts;
output [4:0] sc_st;
output [3:0] sc_sel;
output [31:0] sc_adr;
output [31:0] sc_dat;
input  [2:0] sr_ts;
input  [4:0] sr_rt;
input  [3:0] sr_sel;
input  [31:0] sr_dat;
input  [4:0] chaincommand;
output [4:0] chainresponse;
input  [2:0] e_dp;
input  [2:0] e_ip;
input  [2:0] e_tic;
input  [2:0] r_dp;
input  [2:0] r_ip;
input  [2:0] r_tic;
input  nReset, sc_ack, sr_req, sr_err, sr_rty, sr_acc, sr_mult, 
    nchainresponseack;
output sc_req, sc_we, sc_mult, sc_seq, sc_prd, sr_ack, nchaincommandack;
    wire nroute_ack, rt_ack, routetx_req, ct_ack, ct_defer, ct_slow, ct_ok, 
        routetx_ack, \route[4] , \route[1] , \route[0] , \rt_rd[63] , 
        \rt_rd[62] , \rt_rd[61] , \rt_rd[60] , \rt_rd[59] , \rt_rd[58] , 
        \rt_rd[57] , \rt_rd[56] , \rt_rd[55] , \rt_rd[54] , \rt_rd[53] , 
        \rt_rd[52] , \rt_rd[51] , \rt_rd[50] , \rt_rd[49] , \rt_rd[48] , 
        \rt_rd[47] , \rt_rd[46] , \rt_rd[45] , \rt_rd[44] , \rt_rd[43] , 
        \rt_rd[42] , \rt_rd[41] , \rt_rd[40] , \rt_rd[39] , \rt_rd[38] , 
        \rt_rd[37] , \rt_rd[36] , \rt_rd[35] , \rt_rd[34] , \rt_rd[33] , 
        \rt_rd[32] , \rt_rd[31] , \rt_rd[30] , \rt_rd[29] , \rt_rd[28] , 
        \rt_rd[27] , \rt_rd[26] , \rt_rd[25] , \rt_rd[24] , \rt_rd[23] , 
        \rt_rd[22] , \rt_rd[21] , \rt_rd[20] , \rt_rd[19] , \rt_rd[18] , 
        \rt_rd[17] , \rt_rd[16] , \rt_rd[15] , \rt_rd[14] , \rt_rd[13] , 
        \rt_rd[12] , \rt_rd[11] , \rt_rd[10] , \rt_rd[9] , \rt_rd[8] , 
        \rt_rd[7] , \rt_rd[6] , \rt_rd[5] , \rt_rd[4] , \rt_rd[3] , \rt_rd[2] , 
        \rt_rd[1] , \rt_rd[0] , \rt_err[1] , \rt_err[0] , \ct_wd[63] , 
        \ct_wd[62] , \ct_wd[61] , \ct_wd[60] , \ct_wd[59] , \ct_wd[58] , 
        \ct_wd[57] , \ct_wd[56] , \ct_wd[55] , \ct_wd[54] , \ct_wd[53] , 
        \ct_wd[52] , \ct_wd[51] , \ct_wd[50] , \ct_wd[49] , \ct_wd[48] , 
        \ct_wd[47] , \ct_wd[46] , \ct_wd[45] , \ct_wd[44] , \ct_wd[43] , 
        \ct_wd[42] , \ct_wd[41] , \ct_wd[40] , \ct_wd[39] , \ct_wd[38] , 
        \ct_wd[37] , \ct_wd[36] , \ct_wd[35] , \ct_wd[34] , \ct_wd[33] , 
        \ct_wd[32] , \ct_wd[31] , \ct_wd[30] , \ct_wd[29] , \ct_wd[28] , 
        \ct_wd[27] , \ct_wd[26] , \ct_wd[25] , \ct_wd[24] , \ct_wd[23] , 
        \ct_wd[22] , \ct_wd[21] , \ct_wd[20] , \ct_wd[19] , \ct_wd[18] , 
        \ct_wd[17] , \ct_wd[16] , \ct_wd[15] , \ct_wd[14] , \ct_wd[13] , 
        \ct_wd[12] , \ct_wd[11] , \ct_wd[10] , \ct_wd[9] , \ct_wd[8] , 
        \ct_wd[7] , \ct_wd[6] , \ct_wd[5] , \ct_wd[4] , \ct_wd[3] , \ct_wd[2] , 
        \ct_wd[1] , \ct_wd[0] , \tag_l[4] , \tag_l[3] , \tag_l[2] , \tag_l[1] , 
        \tag_l[0] , \tag_h[4] , \tag_h[3] , \tag_h[2] , \tag_h[1] , \tag_h[0] , 
        \ct_seq[1] , \ct_seq[0] , \ct_lock[1] , \ct_lock[0] , \ct_itag[9] , 
        \ct_itag[8] , \ct_itag[7] , \ct_itag[6] , \ct_itag[5] , \ct_itag[4] , 
        \ct_itag[3] , \ct_itag[2] , \ct_itag[1] , \ct_itag[0] , \ct_size[3] , 
        \ct_size[2] , \ct_size[1] , \ct_size[0] , \ct_rnw[1] , \ct_rnw[0] , 
        \ct_a[63] , \ct_a[62] , \ct_a[61] , \ct_a[60] , \ct_a[59] , \ct_a[58] , 
        \ct_a[57] , \ct_a[56] , \ct_a[55] , \ct_a[54] , \ct_a[53] , \ct_a[52] , 
        \ct_a[51] , \ct_a[50] , \ct_a[49] , \ct_a[48] , \ct_a[47] , \ct_a[46] , 
        \ct_a[45] , \ct_a[44] , \ct_a[43] , \ct_a[42] , \ct_a[41] , \ct_a[40] , 
        \ct_a[39] , \ct_a[38] , \ct_a[37] , \ct_a[36] , \ct_a[35] , \ct_a[34] , 
        \ct_a[33] , \ct_a[32] , \ct_a[31] , \ct_a[30] , \ct_a[29] , \ct_a[28] , 
        \ct_a[27] , \ct_a[26] , \ct_a[25] , \ct_a[24] , \ct_a[23] , \ct_a[22] , 
        \ct_a[21] , \ct_a[20] , \ct_a[19] , \ct_a[18] , \ct_a[17] , \ct_a[16] , 
        \ct_a[15] , \ct_a[14] , \ct_a[13] , \ct_a[12] , \ct_a[11] , \ct_a[10] , 
        \ct_a[9] , \ct_a[8] , \ct_a[7] , \ct_a[6] , \ct_a[5] , \ct_a[4] , 
        \ct_a[3] , \ct_a[2] , \ct_a[1] , \ct_a[0] , \rl[2] , \rl[1] , \rl[0] , 
        \rh[2] , \rh[1] , SYNOPSYS_UNCONNECTED_2, \el[2] , \el[1] , \el[0] , 
        SYNOPSYS_UNCONNECTED_1, \eh[1] , \eh[0] , SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4, reset, SYNOPSYS_UNCONNECTED_5;
    assign sc_prd = 1'b0;
    assign sc_ts[2] = 1'b0;
    assign sc_ts[1] = 1'b0;
    assign sc_ts[0] = 1'b0;
    assign sc_sel[0] = 1'b1;
    target_imem tg ( .addr({\ct_a[63] , \ct_a[62] , \ct_a[61] , \ct_a[60] , 
        \ct_a[59] , \ct_a[58] , \ct_a[57] , \ct_a[56] , \ct_a[55] , \ct_a[54] , 
        \ct_a[53] , \ct_a[52] , \ct_a[51] , \ct_a[50] , \ct_a[49] , \ct_a[48] , 
        \ct_a[47] , \ct_a[46] , \ct_a[45] , \ct_a[44] , \ct_a[43] , \ct_a[42] , 
        \ct_a[41] , \ct_a[40] , \ct_a[39] , \ct_a[38] , \ct_a[37] , \ct_a[36] , 
        \ct_a[35] , \ct_a[34] , \ct_a[33] , \ct_a[32] , \ct_a[31] , \ct_a[30] , 
        \ct_a[29] , \ct_a[28] , \ct_a[27] , \ct_a[26] , \ct_a[25] , \ct_a[24] , 
        \ct_a[23] , \ct_a[22] , \ct_a[21] , \ct_a[20] , \ct_a[19] , \ct_a[18] , 
        \ct_a[17] , \ct_a[16] , \ct_a[15] , \ct_a[14] , \ct_a[13] , \ct_a[12] , 
        \ct_a[11] , \ct_a[10] , \ct_a[9] , \ct_a[8] , \ct_a[7] , \ct_a[6] , 
        \ct_a[5] , \ct_a[4] , \ct_a[3] , \ct_a[2] , \ct_a[1] , \ct_a[0] }), 
        .chainresponse(chainresponse), .crnw({\ct_rnw[1] , \ct_rnw[0] }), 
        .csize({\ct_size[3] , \ct_size[2] , \ct_size[1] , \ct_size[0] }), 
        .ctag({\ct_itag[9] , \ct_itag[8] , \ct_itag[7] , \ct_itag[6] , 
        \ct_itag[5] , \ct_itag[4] , \ct_itag[3] , \ct_itag[2] , \ct_itag[1] , 
        \ct_itag[0] }), .lock({\ct_lock[1] , \ct_lock[0] }), 
        .nchaincommandack(nchaincommandack), .nrouteack(nroute_ack), .rack(
        rt_ack), .routetxreq(routetx_req), .seq({\ct_seq[1] , \ct_seq[0] }), 
        .tag_h({\tag_h[4] , \tag_h[3] , \tag_h[2] , \tag_h[1] , \tag_h[0] }), 
        .tag_l({\tag_l[4] , \tag_l[3] , \tag_l[2] , \tag_l[1] , \tag_l[0] }), 
        .wd({\ct_wd[63] , \ct_wd[62] , \ct_wd[61] , \ct_wd[60] , \ct_wd[59] , 
        \ct_wd[58] , \ct_wd[57] , \ct_wd[56] , \ct_wd[55] , \ct_wd[54] , 
        \ct_wd[53] , \ct_wd[52] , \ct_wd[51] , \ct_wd[50] , \ct_wd[49] , 
        \ct_wd[48] , \ct_wd[47] , \ct_wd[46] , \ct_wd[45] , \ct_wd[44] , 
        \ct_wd[43] , \ct_wd[42] , \ct_wd[41] , \ct_wd[40] , \ct_wd[39] , 
        \ct_wd[38] , \ct_wd[37] , \ct_wd[36] , \ct_wd[35] , \ct_wd[34] , 
        \ct_wd[33] , \ct_wd[32] , \ct_wd[31] , \ct_wd[30] , \ct_wd[29] , 
        \ct_wd[28] , \ct_wd[27] , \ct_wd[26] , \ct_wd[25] , \ct_wd[24] , 
        \ct_wd[23] , \ct_wd[22] , \ct_wd[21] , \ct_wd[20] , \ct_wd[19] , 
        \ct_wd[18] , \ct_wd[17] , \ct_wd[16] , \ct_wd[15] , \ct_wd[14] , 
        \ct_wd[13] , \ct_wd[12] , \ct_wd[11] , \ct_wd[10] , \ct_wd[9] , 
        \ct_wd[8] , \ct_wd[7] , \ct_wd[6] , \ct_wd[5] , \ct_wd[4] , \ct_wd[3] , 
        \ct_wd[2] , \ct_wd[1] , \ct_wd[0] }), .cack(ct_ack), .cdefer(ct_defer), 
        .chaincommand(chaincommand), .cndefer(ct_slow), .cok(ct_ok), .err({
        \rt_err[1] , \rt_err[0] }), .nReset(nReset), .nchainresponseack(
        nchainresponseack), .rd({\rt_rd[63] , \rt_rd[62] , \rt_rd[61] , 
        \rt_rd[60] , \rt_rd[59] , \rt_rd[58] , \rt_rd[57] , \rt_rd[56] , 
        \rt_rd[55] , \rt_rd[54] , \rt_rd[53] , \rt_rd[52] , \rt_rd[51] , 
        \rt_rd[50] , \rt_rd[49] , \rt_rd[48] , \rt_rd[47] , \rt_rd[46] , 
        \rt_rd[45] , \rt_rd[44] , \rt_rd[43] , \rt_rd[42] , \rt_rd[41] , 
        \rt_rd[40] , \rt_rd[39] , \rt_rd[38] , \rt_rd[37] , \rt_rd[36] , 
        \rt_rd[35] , \rt_rd[34] , \rt_rd[33] , \rt_rd[32] , \rt_rd[31] , 
        \rt_rd[30] , \rt_rd[29] , \rt_rd[28] , \rt_rd[27] , \rt_rd[26] , 
        \rt_rd[25] , \rt_rd[24] , \rt_rd[23] , \rt_rd[22] , \rt_rd[21] , 
        \rt_rd[20] , \rt_rd[19] , \rt_rd[18] , \rt_rd[17] , \rt_rd[16] , 
        \rt_rd[15] , \rt_rd[14] , \rt_rd[13] , \rt_rd[12] , \rt_rd[11] , 
        \rt_rd[10] , \rt_rd[9] , \rt_rd[8] , \rt_rd[7] , \rt_rd[6] , 
        \rt_rd[5] , \rt_rd[4] , \rt_rd[3] , \rt_rd[2] , \rt_rd[1] , \rt_rd[0] 
        }), .route({\route[4] , 1'b0, 1'b0, \route[1] , \route[0] }), 
        .routetxack(routetx_ack) );
    t_adec_imem dec ( .e_h({SYNOPSYS_UNCONNECTED_1, \eh[1] , \eh[0] }), .e_l({
        \el[2] , \el[1] , \el[0] }), .r_h({\rh[2] , \rh[1] , 
        SYNOPSYS_UNCONNECTED_2}), .r_l({\rl[2] , \rl[1] , \rl[0] }), .e_dp(
        e_dp), .e_ip(e_ip), .e_tic(e_tic), .r_dp(r_dp), .r_ip(r_ip), .r_tic(
        r_tic), .tag_h({\tag_h[4] , \tag_h[3] , \tag_h[2] , \tag_h[1] , 
        \tag_h[0] }), .tag_l({\tag_l[4] , \tag_l[3] , \tag_l[2] , \tag_l[1] , 
        \tag_l[0] }) );
    resp_route_tx_imem rt ( .o({\route[4] , SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4, \route[1] , \route[0] }), .rtxack(routetx_ack), 
        .e_h({1'b0, \eh[1] , \eh[0] }), .e_l({\el[2] , \el[1] , \el[0] }), 
        .noa(nroute_ack), .r_h({\rh[2] , \rh[1] , 1'b0}), .r_l({\rl[2] , 
        \rl[1] , \rl[0] }), .rtxreq(routetx_req) );
    inv_2 U1 ( .x(reset), .a(nReset) );
    cp2slave_imem chainif2slave ( .tc_seq({\ct_seq[1] , \ct_seq[0] }), 
        .tc_size({\ct_size[3] , \ct_size[2] , \ct_size[1] , \ct_size[0] }), 
        .tc_itag({\ct_itag[9] , \ct_itag[8] , \ct_itag[7] , \ct_itag[6] , 
        \ct_itag[5] , \ct_itag[4] , \ct_itag[3] , \ct_itag[2] , \ct_itag[1] , 
        \ct_itag[0] }), .tc_wd({\ct_wd[63] , \ct_wd[62] , \ct_wd[61] , 
        \ct_wd[60] , \ct_wd[59] , \ct_wd[58] , \ct_wd[57] , \ct_wd[56] , 
        \ct_wd[55] , \ct_wd[54] , \ct_wd[53] , \ct_wd[52] , \ct_wd[51] , 
        \ct_wd[50] , \ct_wd[49] , \ct_wd[48] , \ct_wd[47] , \ct_wd[46] , 
        \ct_wd[45] , \ct_wd[44] , \ct_wd[43] , \ct_wd[42] , \ct_wd[41] , 
        \ct_wd[40] , \ct_wd[39] , \ct_wd[38] , \ct_wd[37] , \ct_wd[36] , 
        \ct_wd[35] , \ct_wd[34] , \ct_wd[33] , \ct_wd[32] , \ct_wd[31] , 
        \ct_wd[30] , \ct_wd[29] , \ct_wd[28] , \ct_wd[27] , \ct_wd[26] , 
        \ct_wd[25] , \ct_wd[24] , \ct_wd[23] , \ct_wd[22] , \ct_wd[21] , 
        \ct_wd[20] , \ct_wd[19] , \ct_wd[18] , \ct_wd[17] , \ct_wd[16] , 
        \ct_wd[15] , \ct_wd[14] , \ct_wd[13] , \ct_wd[12] , \ct_wd[11] , 
        \ct_wd[10] , \ct_wd[9] , \ct_wd[8] , \ct_wd[7] , \ct_wd[6] , 
        \ct_wd[5] , \ct_wd[4] , \ct_wd[3] , \ct_wd[2] , \ct_wd[1] , \ct_wd[0] 
        }), .tc_lock({\ct_lock[1] , \ct_lock[0] }), .tc_a({\ct_a[63] , 
        \ct_a[62] , \ct_a[61] , \ct_a[60] , \ct_a[59] , \ct_a[58] , \ct_a[57] , 
        \ct_a[56] , \ct_a[55] , \ct_a[54] , \ct_a[53] , \ct_a[52] , \ct_a[51] , 
        \ct_a[50] , \ct_a[49] , \ct_a[48] , \ct_a[47] , \ct_a[46] , \ct_a[45] , 
        \ct_a[44] , \ct_a[43] , \ct_a[42] , \ct_a[41] , \ct_a[40] , \ct_a[39] , 
        \ct_a[38] , \ct_a[37] , \ct_a[36] , \ct_a[35] , \ct_a[34] , \ct_a[33] , 
        \ct_a[32] , \ct_a[31] , \ct_a[30] , \ct_a[29] , \ct_a[28] , \ct_a[27] , 
        \ct_a[26] , \ct_a[25] , \ct_a[24] , \ct_a[23] , \ct_a[22] , \ct_a[21] , 
        \ct_a[20] , \ct_a[19] , \ct_a[18] , \ct_a[17] , \ct_a[16] , \ct_a[15] , 
        \ct_a[14] , \ct_a[13] , \ct_a[12] , \ct_a[11] , \ct_a[10] , \ct_a[9] , 
        \ct_a[8] , \ct_a[7] , \ct_a[6] , \ct_a[5] , \ct_a[4] , \ct_a[3] , 
        \ct_a[2] , \ct_a[1] , \ct_a[0] }), .tc_rnw({\ct_rnw[1] , \ct_rnw[0] }), 
        .tc_ok(ct_ok), .tc_defer(ct_defer), .tc_slow(ct_slow), .tc_ack(ct_ack), 
        .req_in(sc_req), .st_i(sc_st), .we_i(sc_we), .mult_i(sc_mult), .adr_i(
        sc_adr), .dat_i(sc_dat), .seq_i(sc_seq), .sel_i({sc_sel[3], sc_sel[2], 
        sc_sel[1], SYNOPSYS_UNCONNECTED_5}), .ack_in(sc_ack), .tr_rd({
        \rt_rd[63] , \rt_rd[62] , \rt_rd[61] , \rt_rd[60] , \rt_rd[59] , 
        \rt_rd[58] , \rt_rd[57] , \rt_rd[56] , \rt_rd[55] , \rt_rd[54] , 
        \rt_rd[53] , \rt_rd[52] , \rt_rd[51] , \rt_rd[50] , \rt_rd[49] , 
        \rt_rd[48] , \rt_rd[47] , \rt_rd[46] , \rt_rd[45] , \rt_rd[44] , 
        \rt_rd[43] , \rt_rd[42] , \rt_rd[41] , \rt_rd[40] , \rt_rd[39] , 
        \rt_rd[38] , \rt_rd[37] , \rt_rd[36] , \rt_rd[35] , \rt_rd[34] , 
        \rt_rd[33] , \rt_rd[32] , \rt_rd[31] , \rt_rd[30] , \rt_rd[29] , 
        \rt_rd[28] , \rt_rd[27] , \rt_rd[26] , \rt_rd[25] , \rt_rd[24] , 
        \rt_rd[23] , \rt_rd[22] , \rt_rd[21] , \rt_rd[20] , \rt_rd[19] , 
        \rt_rd[18] , \rt_rd[17] , \rt_rd[16] , \rt_rd[15] , \rt_rd[14] , 
        \rt_rd[13] , \rt_rd[12] , \rt_rd[11] , \rt_rd[10] , \rt_rd[9] , 
        \rt_rd[8] , \rt_rd[7] , \rt_rd[6] , \rt_rd[5] , \rt_rd[4] , \rt_rd[3] , 
        \rt_rd[2] , \rt_rd[1] , \rt_rd[0] }), .tr_err({\rt_err[1] , 
        \rt_err[0] }), .tr_ack(rt_ack), .req_out(sr_req), .dat_o(sr_dat), 
        .err_o(sr_err), .rty_o(sr_rty), .acc_o(sr_acc), .sel_o(sr_sel), 
        .mult_o(sr_mult), .rt_o(sr_rt), .ack_out(sr_ack), .reset(reset) );
endmodule


module aspida_net_core ( nrst, clk, ip_c_req, ip_c_we, ip_c_mult, ip_c_prd, 
    ip_c_seq, ip_c_ts, ip_c_sel, ip_c_adr, ip_c_dat, ip_c_ack, ip_r_req, 
    ip_r_we, ip_r_err, ip_r_rty, ip_r_acc, ip_r_ts, ip_r_sel, ip_r_dat, 
    ip_r_ack, dp_c_req, dp_c_we, dp_c_mult, dp_c_prd, dp_c_seq, dp_c_ts, 
    dp_c_sel, dp_c_adr, dp_c_dat, dp_c_ack, dp_r_req, dp_r_we, dp_r_err, 
    dp_r_rty, dp_r_acc, dp_r_ts, dp_r_sel, dp_r_dat, dp_r_ack, ei_c_req, 
    ei_c_ack, ei_c_we, ei_c_addr, ei_r_req, ei_r_ack, ei_data_in, ei_data_out, 
    c_BC, c_BC_ack, r_BC, r_BC_ack, wish_we_o, wish_stb_cyc_o, wish_ack_i, 
    wish_adr_o, wish_dat_i, wish_dat_o, dm_c_req, dm_c_we, dm_c_mult, dm_c_seq, 
    dm_c_prd, dm_c_ts, dm_c_st, dm_c_sel, dm_c_adr, dm_c_dat, dm_c_ack, 
    dm_r_req, dm_r_err, dm_r_rty, dm_r_acc, dm_r_mult, dm_r_ts, dm_r_rt, 
    dm_r_sel, dm_r_dat, dm_r_ack, im_c_req, im_c_we, im_c_mult, im_c_seq, 
    im_c_prd, im_c_ts, im_c_st, im_c_sel, im_c_adr, im_c_dat, im_c_ack, 
    im_r_req, im_r_err, im_r_rty, im_r_acc, im_r_mult, im_r_ts, im_r_rt, 
    im_r_sel, im_r_dat, im_r_ack, test_si, test_so, test_se, phi1, phi2, phi3, 
    force_bare );
input  [2:0] ip_c_ts;
input  [3:0] ip_c_sel;
input  [31:0] ip_c_adr;
input  [31:0] ip_c_dat;
output [2:0] ip_r_ts;
output [3:0] ip_r_sel;
output [31:0] ip_r_dat;
input  [2:0] dp_c_ts;
input  [3:0] dp_c_sel;
input  [31:0] dp_c_adr;
input  [31:0] dp_c_dat;
output [2:0] dp_r_ts;
output [3:0] dp_r_sel;
output [31:0] dp_r_dat;
input  [10:0] ei_c_addr;
input  [7:0] ei_data_in;
output [7:0] ei_data_out;
output [4:0] c_BC;
input  [4:0] r_BC;
output [11:0] wish_adr_o;
input  [31:0] wish_dat_i;
output [31:0] wish_dat_o;
output [2:0] dm_c_ts;
output [4:0] dm_c_st;
output [3:0] dm_c_sel;
output [31:0] dm_c_adr;
output [31:0] dm_c_dat;
input  [2:0] dm_r_ts;
input  [4:0] dm_r_rt;
input  [3:0] dm_r_sel;
input  [31:0] dm_r_dat;
output [2:0] im_c_ts;
output [4:0] im_c_st;
output [3:0] im_c_sel;
output [31:0] im_c_adr;
output [31:0] im_c_dat;
input  [2:0] im_r_ts;
input  [4:0] im_r_rt;
input  [3:0] im_r_sel;
input  [31:0] im_r_dat;
input  nrst, clk, ip_c_req, ip_c_we, ip_c_mult, ip_c_prd, ip_c_seq, ip_r_ack, 
    dp_c_req, dp_c_we, dp_c_mult, dp_c_prd, dp_c_seq, dp_r_ack, ei_c_req, 
    ei_c_we, ei_r_ack, c_BC_ack, wish_ack_i, dm_c_ack, dm_r_req, dm_r_err, 
    dm_r_rty, dm_r_acc, dm_r_mult, im_c_ack, im_r_req, im_r_err, im_r_rty, 
    im_r_acc, im_r_mult, test_si, test_se, phi1, phi2, phi3, force_bare;
output ip_c_ack, ip_r_req, ip_r_we, ip_r_err, ip_r_rty, ip_r_acc, dp_c_ack, 
    dp_r_req, dp_r_we, dp_r_err, dp_r_rty, dp_r_acc, ei_c_ack, ei_r_req, 
    r_BC_ack, wish_we_o, wish_stb_cyc_o, dm_c_req, dm_c_we, dm_c_mult, 
    dm_c_seq, dm_c_prd, dm_r_ack, im_c_req, im_c_we, im_c_mult, im_c_seq, 
    im_c_prd, im_r_ack, test_so;
    wire n1, real_c_Iport_ack, r_Iport_ack, \r_Iport[4] , \r_Iport[3] , 
        \r_Iport[2] , \r_Iport[1] , \r_Iport[0] , \c_Iport[4] , \c_Iport[3] , 
        \c_Iport[2] , \c_Iport[1] , \c_Iport[0] , n3, real_c_Dport_ack, 
        r_Dport_ack, \r_Dport[4] , \r_Dport[3] , \r_Dport[2] , \r_Dport[1] , 
        \r_Dport[0] , \c_Dport[4] , \c_Dport[3] , \c_Dport[2] , \c_Dport[1] , 
        \c_Dport[0] , tic_c_req, tic_c_we, tic_c_ack, tic_r_req, tic_r_ack, 
        real_c_TIC_ack, r_TIC_ack, \r_TIC[4] , \r_TIC[3] , \r_TIC[2] , 
        \r_TIC[1] , \r_TIC[0] , \c_TIC[4] , \c_TIC[3] , \c_TIC[2] , \c_TIC[1] , 
        \c_TIC[0] , \tic_r_dat[31] , \tic_r_dat[30] , \tic_r_dat[29] , 
        \tic_r_dat[28] , \tic_r_dat[27] , \tic_r_dat[26] , \tic_r_dat[25] , 
        \tic_r_dat[24] , \tic_r_dat[23] , \tic_r_dat[22] , \tic_r_dat[21] , 
        \tic_r_dat[20] , \tic_r_dat[19] , \tic_r_dat[18] , \tic_r_dat[17] , 
        \tic_r_dat[16] , \tic_r_dat[15] , \tic_r_dat[14] , \tic_r_dat[13] , 
        \tic_r_dat[12] , \tic_r_dat[11] , \tic_r_dat[10] , \tic_r_dat[9] , 
        \tic_r_dat[8] , \tic_r_dat[7] , \tic_r_dat[6] , \tic_r_dat[5] , 
        \tic_r_dat[4] , \tic_r_dat[3] , \tic_r_dat[2] , \tic_r_dat[1] , 
        \tic_r_dat[0] , \tic_c_dat[31] , \tic_c_dat[30] , \tic_c_dat[29] , 
        \tic_c_dat[28] , \tic_c_dat[27] , \tic_c_dat[26] , \tic_c_dat[25] , 
        \tic_c_dat[24] , \tic_c_dat[23] , \tic_c_dat[22] , \tic_c_dat[21] , 
        \tic_c_dat[20] , \tic_c_dat[19] , \tic_c_dat[18] , \tic_c_dat[17] , 
        \tic_c_dat[16] , \tic_c_dat[15] , \tic_c_dat[14] , \tic_c_dat[13] , 
        \tic_c_dat[12] , \tic_c_dat[11] , \tic_c_dat[10] , \tic_c_dat[9] , 
        \tic_c_dat[8] , \tic_c_dat[7] , \tic_c_dat[6] , \tic_c_dat[5] , 
        \tic_c_dat[4] , \tic_c_dat[3] , \tic_c_dat[2] , \tic_c_dat[1] , 
        \tic_c_dat[0] , \tic_c_adr[31] , \tic_c_adr[30] , \tic_c_adr[11] , 
        \tic_c_adr[10] , \tic_c_adr[9] , \tic_c_adr[8] , \tic_c_adr[7] , 
        \tic_c_adr[6] , \tic_c_adr[5] , \tic_c_adr[4] , \tic_c_adr[3] , 
        \tic_c_adr[2] , n4, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, 
        SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, 
        SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, 
        SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10, 
        SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12, 
        SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14, 
        SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16, 
        SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18, 
        SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20, c_BC_ack_n, 
        c_WB_ack_n, c_WB_ack, c_IMEM_ack_n, c_IMEM_ack, c_DMEM_ack_n, 
        c_DMEM_ack, n2, c_Iport_ack, c_TIC_ack, c_Dport_ack, \c_WB[4] , 
        \c_WB[0] , \c_WB[1] , \c_WB[2] , \c_WB[3] , \c_IMEM[4] , \c_IMEM[0] , 
        \c_IMEM[1] , \c_IMEM[2] , \c_IMEM[3] , \c_DMEM[4] , \c_DMEM[0] , 
        \c_DMEM[1] , \c_DMEM[2] , \c_DMEM[3] , scan_o_cmd, n12, n9, n15, n6, 
        r_Iport_ack_n, r_TIC_ack_n, r_Dport_ack_n, \r_IMEM[4] , \r_IMEM[0] , 
        \r_IMEM[1] , \r_IMEM[2] , \r_IMEM[3] , r_IMEM_ack, \r_DMEM[4] , 
        \r_DMEM[0] , \r_DMEM[1] , \r_DMEM[2] , \r_DMEM[3] , r_DMEM_ack, 
        \r_WB[4] , \r_WB[0] , \r_WB[1] , \r_WB[2] , \r_WB[3] , r_WB_ack, n13, 
        n10, n16, n7, real_r_WB_ack, real_r_DMEM_ack, real_r_IMEM_ack, n5, n14, 
        n11, n8, rst;
    assign ip_r_sel[3] = 1'b0;
    assign ip_r_sel[2] = 1'b0;
    assign ip_r_sel[1] = 1'b0;
    assign ip_r_sel[0] = 1'b0;
    assign dp_r_sel[3] = 1'b0;
    assign dp_r_sel[2] = 1'b0;
    assign dp_r_sel[1] = 1'b0;
    assign dp_r_sel[0] = 1'b0;
    master_if_iport iport ( .nReset(n1), .mc_req(ip_c_req), .mc_we(ip_c_we), 
        .mc_mult(ip_c_mult), .mc_prd(ip_c_prd), .mc_seq(ip_c_seq), .mc_ts(
        ip_c_ts), .mc_sel(ip_c_sel), .mc_adr(ip_c_adr), .mc_dat(ip_c_dat), 
        .mc_ack(ip_c_ack), .mr_req(ip_r_req), .mr_we(ip_r_we), .mr_err(
        ip_r_err), .mr_rty(ip_r_rty), .mr_acc(ip_r_acc), .mr_ts(ip_r_ts), 
        .mr_dat(ip_r_dat), .mr_ack(ip_r_ack), .chaincommand({\c_Iport[4] , 
        \c_Iport[3] , \c_Iport[2] , \c_Iport[1] , \c_Iport[0] }), 
        .nchaincommandack(real_c_Iport_ack), .chainresponse({\r_Iport[4] , 
        \r_Iport[3] , \r_Iport[2] , \r_Iport[1] , \r_Iport[0] }), 
        .nchainresponseack(r_Iport_ack), .e_bare({1'b0, 1'b0, 1'b1, 1'b0}), 
        .e_dm({1'b0, 1'b0, 1'b0, 1'b1}), .e_im({1'b0, 1'b0, 1'b0, 1'b1}), 
        .e_wish({1'b0, 1'b1, 1'b0, 1'b0}), .r_bare({1'b1, 1'b0, 1'b0, 1'b0}), 
        .r_dm({1'b1, 1'b1, 1'b1, 1'b0}), .r_im({1'b1, 1'b1, 1'b0, 1'b0}), 
        .r_wish({1'b0, 1'b0, 1'b0, 1'b0}), .tag_id({1'b1, 1'b0, 1'b0, 1'b0, 
        1'b0}), .force_bare(force_bare) );
    master_if_dport dport ( .nReset(n3), .mc_req(dp_c_req), .mc_we(dp_c_we), 
        .mc_mult(dp_c_mult), .mc_prd(dp_c_prd), .mc_seq(dp_c_seq), .mc_ts(
        dp_c_ts), .mc_sel(dp_c_sel), .mc_adr(dp_c_adr), .mc_dat(dp_c_dat), 
        .mc_ack(dp_c_ack), .mr_req(dp_r_req), .mr_we(dp_r_we), .mr_err(
        dp_r_err), .mr_rty(dp_r_rty), .mr_acc(dp_r_acc), .mr_ts(dp_r_ts), 
        .mr_dat(dp_r_dat), .mr_ack(dp_r_ack), .chaincommand({\c_Dport[4] , 
        \c_Dport[3] , \c_Dport[2] , \c_Dport[1] , \c_Dport[0] }), 
        .nchaincommandack(real_c_Dport_ack), .chainresponse({\r_Dport[4] , 
        \r_Dport[3] , \r_Dport[2] , \r_Dport[1] , \r_Dport[0] }), 
        .nchainresponseack(r_Dport_ack), .e_bare({1'b0, 1'b0, 1'b1, 1'b0}), 
        .e_dm({1'b0, 1'b0, 1'b0, 1'b1}), .e_im({1'b0, 1'b0, 1'b0, 1'b1}), 
        .e_wish({1'b0, 1'b1, 1'b0, 1'b0}), .r_bare({1'b1, 1'b0, 1'b0, 1'b0}), 
        .r_dm({1'b1, 1'b1, 1'b1, 1'b0}), .r_im({1'b1, 1'b1, 1'b0, 1'b0}), 
        .r_wish({1'b0, 1'b0, 1'b0, 1'b0}), .tag_id({1'b0, 1'b1, 1'b0, 1'b0, 
        1'b0}), .force_bare(force_bare) );
    master_if_tic tic ( .nReset(n3), .mc_req(tic_c_req), .mc_we(tic_c_we), 
        .mc_mult(1'b0), .mc_prd(1'b0), .mc_seq(1'b0), .mc_ts({1'b0, 1'b0, 1'b0
        }), .mc_sel({1'b1, 1'b1, 1'b1, 1'b1}), .mc_adr({\tic_c_adr[31] , 
        \tic_c_adr[30] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \tic_c_adr[11] , 
        \tic_c_adr[10] , \tic_c_adr[9] , \tic_c_adr[8] , \tic_c_adr[7] , 
        \tic_c_adr[6] , \tic_c_adr[5] , \tic_c_adr[4] , \tic_c_adr[3] , 
        \tic_c_adr[2] , 1'b0, 1'b0}), .mc_dat({\tic_c_dat[31] , 
        \tic_c_dat[30] , \tic_c_dat[29] , \tic_c_dat[28] , \tic_c_dat[27] , 
        \tic_c_dat[26] , \tic_c_dat[25] , \tic_c_dat[24] , \tic_c_dat[23] , 
        \tic_c_dat[22] , \tic_c_dat[21] , \tic_c_dat[20] , \tic_c_dat[19] , 
        \tic_c_dat[18] , \tic_c_dat[17] , \tic_c_dat[16] , \tic_c_dat[15] , 
        \tic_c_dat[14] , \tic_c_dat[13] , \tic_c_dat[12] , \tic_c_dat[11] , 
        \tic_c_dat[10] , \tic_c_dat[9] , \tic_c_dat[8] , \tic_c_dat[7] , 
        \tic_c_dat[6] , \tic_c_dat[5] , \tic_c_dat[4] , \tic_c_dat[3] , 
        \tic_c_dat[2] , \tic_c_dat[1] , \tic_c_dat[0] }), .mc_ack(tic_c_ack), 
        .mr_req(tic_r_req), .mr_dat({\tic_r_dat[31] , \tic_r_dat[30] , 
        \tic_r_dat[29] , \tic_r_dat[28] , \tic_r_dat[27] , \tic_r_dat[26] , 
        \tic_r_dat[25] , \tic_r_dat[24] , \tic_r_dat[23] , \tic_r_dat[22] , 
        \tic_r_dat[21] , \tic_r_dat[20] , \tic_r_dat[19] , \tic_r_dat[18] , 
        \tic_r_dat[17] , \tic_r_dat[16] , \tic_r_dat[15] , \tic_r_dat[14] , 
        \tic_r_dat[13] , \tic_r_dat[12] , \tic_r_dat[11] , \tic_r_dat[10] , 
        \tic_r_dat[9] , \tic_r_dat[8] , \tic_r_dat[7] , \tic_r_dat[6] , 
        \tic_r_dat[5] , \tic_r_dat[4] , \tic_r_dat[3] , \tic_r_dat[2] , 
        \tic_r_dat[1] , \tic_r_dat[0] }), .mr_ack(tic_r_ack), .chaincommand({
        \c_TIC[4] , \c_TIC[3] , \c_TIC[2] , \c_TIC[1] , \c_TIC[0] }), 
        .nchaincommandack(real_c_TIC_ack), .chainresponse({\r_TIC[4] , 
        \r_TIC[3] , \r_TIC[2] , \r_TIC[1] , \r_TIC[0] }), .nchainresponseack(
        r_TIC_ack), .e_bare({1'b0, 1'b0, 1'b1, 1'b0}), .e_dm({1'b0, 1'b0, 1'b0, 
        1'b1}), .e_im({1'b0, 1'b0, 1'b0, 1'b1}), .e_wish({1'b0, 1'b1, 1'b0, 
        1'b0}), .r_bare({1'b1, 1'b0, 1'b0, 1'b0}), .r_dm({1'b1, 1'b1, 1'b1, 
        1'b0}), .r_im({1'b1, 1'b1, 1'b0, 1'b0}), .r_wish({1'b0, 1'b0, 1'b0, 
        1'b0}), .tag_id({1'b0, 1'b0, 1'b1, 1'b0, 1'b0}), .force_bare(
        force_bare) );
    tic ticBlock ( .c_req(ei_c_req), .c_ack(ei_c_ack), .c_we(ei_c_we), 
        .c_addr(ei_c_addr), .r_req(ei_r_req), .r_ack(ei_r_ack), .data_in(
        ei_data_in), .data_out(ei_data_out), .reset_b(n4), .mc_req(tic_c_req), 
        .mc_we(tic_c_we), .mc_adr({\tic_c_adr[31] , \tic_c_adr[30] , 
        SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, 
        SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, \tic_c_adr[11] , \tic_c_adr[10] , 
        \tic_c_adr[9] , \tic_c_adr[8] , \tic_c_adr[7] , \tic_c_adr[6] , 
        \tic_c_adr[5] , \tic_c_adr[4] , \tic_c_adr[3] , \tic_c_adr[2] , 
        SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20}), .mc_dat({
        \tic_c_dat[31] , \tic_c_dat[30] , \tic_c_dat[29] , \tic_c_dat[28] , 
        \tic_c_dat[27] , \tic_c_dat[26] , \tic_c_dat[25] , \tic_c_dat[24] , 
        \tic_c_dat[23] , \tic_c_dat[22] , \tic_c_dat[21] , \tic_c_dat[20] , 
        \tic_c_dat[19] , \tic_c_dat[18] , \tic_c_dat[17] , \tic_c_dat[16] , 
        \tic_c_dat[15] , \tic_c_dat[14] , \tic_c_dat[13] , \tic_c_dat[12] , 
        \tic_c_dat[11] , \tic_c_dat[10] , \tic_c_dat[9] , \tic_c_dat[8] , 
        \tic_c_dat[7] , \tic_c_dat[6] , \tic_c_dat[5] , \tic_c_dat[4] , 
        \tic_c_dat[3] , \tic_c_dat[2] , \tic_c_dat[1] , \tic_c_dat[0] }), 
        .mc_ack(tic_c_ack), .mr_req(tic_r_req), .mr_dat({\tic_r_dat[31] , 
        \tic_r_dat[30] , \tic_r_dat[29] , \tic_r_dat[28] , \tic_r_dat[27] , 
        \tic_r_dat[26] , \tic_r_dat[25] , \tic_r_dat[24] , \tic_r_dat[23] , 
        \tic_r_dat[22] , \tic_r_dat[21] , \tic_r_dat[20] , \tic_r_dat[19] , 
        \tic_r_dat[18] , \tic_r_dat[17] , \tic_r_dat[16] , \tic_r_dat[15] , 
        \tic_r_dat[14] , \tic_r_dat[13] , \tic_r_dat[12] , \tic_r_dat[11] , 
        \tic_r_dat[10] , \tic_r_dat[9] , \tic_r_dat[8] , \tic_r_dat[7] , 
        \tic_r_dat[6] , \tic_r_dat[5] , \tic_r_dat[4] , \tic_r_dat[3] , 
        \tic_r_dat[2] , \tic_r_dat[1] , \tic_r_dat[0] }), .mr_ack(tic_r_ack)
         );
    inv_2 U10 ( .x(c_BC_ack_n), .a(c_BC_ack) );
    inv_2 U12 ( .x(c_WB_ack_n), .a(c_WB_ack) );
    inv_2 U13 ( .x(c_IMEM_ack_n), .a(c_IMEM_ack) );
    inv_2 U14 ( .x(c_DMEM_ack_n), .a(c_DMEM_ack) );
    comm_fab_scan cmd_fab ( .nrst(n2), .I_port_eop_i(\c_Iport[4] ), 
        .I_port_d0_i(\c_Iport[0] ), .I_port_d1_i(\c_Iport[1] ), .I_port_d2_i(
        \c_Iport[2] ), .I_port_d3_i(\c_Iport[3] ), .I_port_ack(c_Iport_ack), 
        .TIC_eop_i(\c_TIC[4] ), .TIC_d0_i(\c_TIC[0] ), .TIC_d1_i(\c_TIC[1] ), 
        .TIC_d2_i(\c_TIC[2] ), .TIC_d3_i(\c_TIC[3] ), .TIC_ack(c_TIC_ack), 
        .D_port_eop_i(\c_Dport[4] ), .D_port_d0_i(\c_Dport[0] ), .D_port_d1_i(
        \c_Dport[1] ), .D_port_d2_i(\c_Dport[2] ), .D_port_d3_i(\c_Dport[3] ), 
        .D_port_ack(c_Dport_ack), .BC_eop_i(c_BC[4]), .BC_d0_i(c_BC[0]), 
        .BC_d1_i(c_BC[1]), .BC_d2_i(c_BC[2]), .BC_d3_i(c_BC[3]), .BC_ack(
        c_BC_ack_n), .WB_eop_i(\c_WB[4] ), .WB_d0_i(\c_WB[0] ), .WB_d1_i(
        \c_WB[1] ), .WB_d2_i(\c_WB[2] ), .WB_d3_i(\c_WB[3] ), .WB_ack(
        c_WB_ack_n), .IMEM_eop_i(\c_IMEM[4] ), .IMEM_d0_i(\c_IMEM[0] ), 
        .IMEM_d1_i(\c_IMEM[1] ), .IMEM_d2_i(\c_IMEM[2] ), .IMEM_d3_i(
        \c_IMEM[3] ), .IMEM_ack(c_IMEM_ack_n), .DMEM_eop_i(\c_DMEM[4] ), 
        .DMEM_d0_i(\c_DMEM[0] ), .DMEM_d1_i(\c_DMEM[1] ), .DMEM_d2_i(
        \c_DMEM[2] ), .DMEM_d3_i(\c_DMEM[3] ), .DMEM_ack(c_DMEM_ack_n), 
        .test_si(test_si), .test_so(scan_o_cmd), .test_se(n12), .phi1(n9), 
        .phi2(n15), .phi3(n6) );
    inv_2 U20 ( .x(r_Iport_ack_n), .a(r_Iport_ack) );
    inv_2 U21 ( .x(r_TIC_ack_n), .a(r_TIC_ack) );
    inv_2 U22 ( .x(r_Dport_ack_n), .a(r_Dport_ack) );
    resp_fab_scan rsp_fab ( .nrst(n3), .IMEM_eop_i(\r_IMEM[4] ), .IMEM_d0_i(
        \r_IMEM[0] ), .IMEM_d1_i(\r_IMEM[1] ), .IMEM_d2_i(\r_IMEM[2] ), 
        .IMEM_d3_i(\r_IMEM[3] ), .IMEM_ack(r_IMEM_ack), .DMEM_eop_i(
        \r_DMEM[4] ), .DMEM_d0_i(\r_DMEM[0] ), .DMEM_d1_i(\r_DMEM[1] ), 
        .DMEM_d2_i(\r_DMEM[2] ), .DMEM_d3_i(\r_DMEM[3] ), .DMEM_ack(r_DMEM_ack
        ), .WB_eop_i(\r_WB[4] ), .WB_d0_i(\r_WB[0] ), .WB_d1_i(\r_WB[1] ), 
        .WB_d2_i(\r_WB[2] ), .WB_d3_i(\r_WB[3] ), .WB_ack(r_WB_ack), 
        .BC_eop_i(r_BC[4]), .BC_d0_i(r_BC[0]), .BC_d1_i(r_BC[1]), .BC_d2_i(
        r_BC[2]), .BC_d3_i(r_BC[3]), .BC_ack(r_BC_ack), .I_port_eop_i(
        \r_Iport[4] ), .I_port_d0_i(\r_Iport[0] ), .I_port_d1_i(\r_Iport[1] ), 
        .I_port_d2_i(\r_Iport[2] ), .I_port_d3_i(\r_Iport[3] ), .I_port_ack(
        r_Iport_ack_n), .TIC_eop_i(\r_TIC[4] ), .TIC_d0_i(\r_TIC[0] ), 
        .TIC_d1_i(\r_TIC[1] ), .TIC_d2_i(\r_TIC[2] ), .TIC_d3_i(\r_TIC[3] ), 
        .TIC_ack(r_TIC_ack_n), .D_port_eop_i(\r_Dport[4] ), .D_port_d0_i(
        \r_Dport[0] ), .D_port_d1_i(\r_Dport[1] ), .D_port_d2_i(\r_Dport[2] ), 
        .D_port_d3_i(\r_Dport[3] ), .D_port_ack(r_Dport_ack_n), .test_si(
        scan_o_cmd), .test_so(test_so), .test_se(n13), .phi1(n10), .phi2(n16), 
        .phi3(n7) );
    wb_block wb ( .nReset(n1), .clk(clk), .chaincommand({\c_WB[4] , \c_WB[3] , 
        \c_WB[2] , \c_WB[1] , \c_WB[0] }), .nchaincommandack(c_WB_ack), 
        .chainresponse({\r_WB[4] , \r_WB[3] , \r_WB[2] , \r_WB[1] , \r_WB[0] }
        ), .nchainresponseack(real_r_WB_ack), .e_dp({1'b0, 1'b0, 1'b1}), 
        .e_ip({1'b0, 1'b0, 1'b1}), .e_tic({1'b0, 1'b1, 1'b0}), .r_dp({1'b1, 
        1'b0, 1'b0}), .r_ip({1'b1, 1'b1, 1'b0}), .r_tic({1'b0, 1'b0, 1'b0}), 
        .wb_we_o(wish_we_o), .wb_stb_cyc_o(wish_stb_cyc_o), .wb_ack_i(
        wish_ack_i), .wb_adr_o(wish_adr_o), .wb_dat_i(wish_dat_i), .wb_dat_o(
        wish_dat_o) );
    slave_if_dmem dmem ( .nReset(n1), .sc_req(dm_c_req), .sc_we(dm_c_we), 
        .sc_mult(dm_c_mult), .sc_seq(dm_c_seq), .sc_prd(dm_c_prd), .sc_ts(
        dm_c_ts), .sc_st(dm_c_st), .sc_sel(dm_c_sel), .sc_adr(dm_c_adr), 
        .sc_dat(dm_c_dat), .sc_ack(dm_c_ack), .sr_req(dm_r_req), .sr_err(
        dm_r_err), .sr_rty(dm_r_rty), .sr_acc(dm_r_acc), .sr_mult(dm_r_mult), 
        .sr_ts(dm_r_ts), .sr_rt(dm_r_rt), .sr_sel(dm_r_sel), .sr_dat(dm_r_dat), 
        .sr_ack(dm_r_ack), .chaincommand({\c_DMEM[4] , \c_DMEM[3] , 
        \c_DMEM[2] , \c_DMEM[1] , \c_DMEM[0] }), .nchaincommandack(c_DMEM_ack), 
        .chainresponse({\r_DMEM[4] , \r_DMEM[3] , \r_DMEM[2] , \r_DMEM[1] , 
        \r_DMEM[0] }), .nchainresponseack(real_r_DMEM_ack), .e_dp({1'b0, 1'b0, 
        1'b1}), .e_ip({1'b0, 1'b0, 1'b1}), .e_tic({1'b0, 1'b1, 1'b0}), .r_dp({
        1'b1, 1'b0, 1'b0}), .r_ip({1'b1, 1'b1, 1'b0}), .r_tic({1'b0, 1'b0, 
        1'b0}) );
    slave_if_imem imem ( .nReset(n4), .sc_req(im_c_req), .sc_we(im_c_we), 
        .sc_mult(im_c_mult), .sc_seq(im_c_seq), .sc_prd(im_c_prd), .sc_ts(
        im_c_ts), .sc_st(im_c_st), .sc_sel(im_c_sel), .sc_adr(im_c_adr), 
        .sc_dat(im_c_dat), .sc_ack(im_c_ack), .sr_req(im_r_req), .sr_err(
        im_r_err), .sr_rty(im_r_rty), .sr_acc(im_r_acc), .sr_mult(im_r_mult), 
        .sr_ts(im_r_ts), .sr_rt(im_r_rt), .sr_sel(im_r_sel), .sr_dat(im_r_dat), 
        .sr_ack(im_r_ack), .chaincommand({\c_IMEM[4] , \c_IMEM[3] , 
        \c_IMEM[2] , \c_IMEM[1] , \c_IMEM[0] }), .nchaincommandack(c_IMEM_ack), 
        .chainresponse({\r_IMEM[4] , \r_IMEM[3] , \r_IMEM[2] , \r_IMEM[1] , 
        \r_IMEM[0] }), .nchainresponseack(real_r_IMEM_ack), .e_dp({1'b0, 1'b0, 
        1'b1}), .e_ip({1'b0, 1'b0, 1'b1}), .e_tic({1'b0, 1'b1, 1'b0}), .r_dp({
        1'b1, 1'b0, 1'b0}), .r_ip({1'b1, 1'b1, 1'b0}), .r_tic({1'b0, 1'b0, 
        1'b0}) );
    inv_2 U8 ( .x(n6), .a(n5) );
    inv_2 U9 ( .x(n7), .a(n5) );
    inv_2 U11 ( .x(n15), .a(n14) );
    inv_2 U15 ( .x(n13), .a(n11) );
    inv_2 U16 ( .x(n9), .a(n8) );
    inv_2 U17 ( .x(n10), .a(n8) );
    inv_2 U18 ( .x(n12), .a(n11) );
    inv_2 U19 ( .x(n16), .a(n14) );
    buf_3 U23 ( .x(n1), .a(nrst) );
    buf_3 U24 ( .x(n4), .a(nrst) );
    buf_4 U25 ( .x(n2), .a(nrst) );
    buf_4 U26 ( .x(n3), .a(nrst) );
    inv_2 U27 ( .x(n5), .a(phi3) );
    inv_2 U28 ( .x(n8), .a(phi1) );
    inv_5 U29 ( .x(n11), .a(test_se) );
    inv_2 U30 ( .x(n14), .a(phi2) );
    inv_5 U31 ( .x(rst), .a(n4) );
    nor2_4 U32 ( .x(real_c_Dport_ack), .a(rst), .b(c_Dport_ack) );
    nor2_4 U33 ( .x(real_r_IMEM_ack), .a(rst), .b(r_IMEM_ack) );
    nor2_4 U34 ( .x(real_r_DMEM_ack), .a(rst), .b(r_DMEM_ack) );
    nor2_4 U35 ( .x(real_r_WB_ack), .a(rst), .b(r_WB_ack) );
    nor2_4 U36 ( .x(real_c_TIC_ack), .a(rst), .b(c_TIC_ack) );
    nor2_4 U37 ( .x(real_c_Iport_ack), .a(rst), .b(c_Iport_ack) );
endmodule


module ASPIDA_top ( reset_DLX_d_PAD, reset_DLX_c_PAD, sync_async_PAD, INT_PAD, 
    CLI_PAD, FREEZE_PAD, STOP_FETCH_PAD, reset_ctrl_PAD, test_si_DLX_PAD, 
    test_so_DLX_PAD, test_se_PAD, global_g1_PAD, global_g2_PAD, 
    memory_load_enable_PAD, scan_in_PAD, scan_out_PAD, shift_clk_PAD, read_PAD, 
    inst_ram_load_PAD, del_scan_en_PAD, del_scan_in_PAD, ei_c_req_PAD, 
    ei_c_ack_PAD, ei_c_we_PAD, ei_c_addr_PAD, ei_r_req_PAD, ei_r_ack_PAD, 
    ei_data_inout_PAD, r_BC_PAD, r_BC_ack_PAD, c_BC_PAD, c_BC_ack_PAD, 
    wish_clk_PAD, wish_ack_i_PAD, wish_we_o_PAD, wish_stb_cyc_o_PAD, 
    wish_adr_o_PAD, wish_dat_io_PAD, stuckAtVdd_PAD );
input  [10:0] ei_c_addr_PAD;
inout  [7:0] ei_data_inout_PAD;
input  [4:0] r_BC_PAD;
output [4:0] c_BC_PAD;
output [11:0] wish_adr_o_PAD;
inout  [31:0] wish_dat_io_PAD;
input  reset_DLX_d_PAD, reset_DLX_c_PAD, sync_async_PAD, INT_PAD, FREEZE_PAD, 
    STOP_FETCH_PAD, reset_ctrl_PAD, test_si_DLX_PAD, test_se_PAD, 
    global_g1_PAD, global_g2_PAD, memory_load_enable_PAD, scan_in_PAD, 
    shift_clk_PAD, read_PAD, inst_ram_load_PAD, del_scan_en_PAD, 
    del_scan_in_PAD, ei_c_req_PAD, ei_c_we_PAD, ei_r_ack_PAD, c_BC_ack_PAD, 
    wish_clk_PAD, wish_ack_i_PAD;
output CLI_PAD, test_so_DLX_PAD, scan_out_PAD, ei_c_ack_PAD, ei_r_req_PAD, 
    r_BC_ack_PAD, wish_we_o_PAD, wish_stb_cyc_o_PAD, stuckAtVdd_PAD;
    wire STOP_fetch, reset_ctrl, FREEZE, memory_load_enable, scan_in, scan_out, 
        shift_clk, read, inst_ram_load, del_scan_en, del_scan_in, reset_DLX_d, 
        reset_DLX_c, INT, test_si_DLX, test_se, global_g1, global_g2, r_BC_4, 
        r_BC_3, r_BC_2, r_BC_1, r_BC_0, r_BC_ack, c_BC_ack, c_BC_4, c_BC_3, 
        c_BC_2, c_BC_1, c_BC_0, ei_c_req, ei_c_we, ei_c_addr_10, ei_c_addr_9, 
        ei_c_addr_8, ei_c_addr_7, ei_c_addr_6, ei_c_addr_5, ei_c_addr_4, 
        ei_c_addr_3, ei_c_addr_2, ei_c_addr_1, ei_c_addr_0, ei_c_ack, ei_r_req, 
        ei_data_in_7, ei_data_in_6, ei_data_in_5, ei_data_in_4, ei_data_in_3, 
        ei_data_in_2, ei_data_in_1, ei_data_in_0, ei_data_out_7, ei_data_out_6, 
        ei_data_out_5, ei_data_out_4, ei_data_out_3, ei_data_out_2, 
        ei_data_out_1, ei_data_out_0, _17_net_, ei_r_ack, wish_ack_i, wish_clk, 
        wish_stb_cyc_o, wish_we_o, wish_adr_o_11, wish_adr_o_10, wish_adr_o_9, 
        wish_adr_o_8, wish_adr_o_7, wish_adr_o_6, wish_adr_o_5, wish_adr_o_4, 
        wish_adr_o_3, wish_adr_o_2, wish_adr_o_1, wish_adr_o_0, wish_dat_i_31, 
        wish_dat_i_30, wish_dat_i_29, wish_dat_i_28, wish_dat_i_27, 
        wish_dat_i_26, wish_dat_i_25, wish_dat_i_24, wish_dat_i_23, 
        wish_dat_i_22, wish_dat_i_21, wish_dat_i_20, wish_dat_i_19, 
        wish_dat_i_18, wish_dat_i_17, wish_dat_i_16, wish_dat_i_15, 
        wish_dat_i_14, wish_dat_i_13, wish_dat_i_12, wish_dat_i_11, 
        wish_dat_i_10, wish_dat_i_9, wish_dat_i_8, wish_dat_i_7, wish_dat_i_6, 
        wish_dat_i_5, wish_dat_i_4, wish_dat_i_3, wish_dat_i_2, wish_dat_i_1, 
        wish_dat_i_0, wish_dat_o_31, wish_dat_o_30, wish_dat_o_29, 
        wish_dat_o_28, wish_dat_o_27, wish_dat_o_26, wish_dat_o_25, 
        wish_dat_o_24, wish_dat_o_23, wish_dat_o_22, wish_dat_o_21, 
        wish_dat_o_20, wish_dat_o_19, wish_dat_o_18, wish_dat_o_17, 
        wish_dat_o_16, wish_dat_o_15, wish_dat_o_14, wish_dat_o_13, 
        wish_dat_o_12, wish_dat_o_11, wish_dat_o_10, wish_dat_o_9, 
        wish_dat_o_8, wish_dat_o_7, wish_dat_o_6, wish_dat_o_5, wish_dat_o_4, 
        wish_dat_o_3, wish_dat_o_2, wish_dat_o_1, wish_dat_o_0, CLI, 
        reset_DLX_d_ff2, reset_DLX_ctrl, reset_DLX_d_ff1, 
        reset_DLX_d_ff1_shift, IM_addr_31, IM_addr_30, IM_addr_29, IM_addr_28, 
        IM_addr_27, IM_addr_26, IM_addr_25, IM_addr_24, IM_addr_23, IM_addr_22, 
        IM_addr_21, IM_addr_20, IM_addr_19, IM_addr_18, IM_addr_17, IM_addr_16, 
        IM_addr_15, IM_addr_14, IM_addr_13, IM_addr_12, IM_addr_11, IM_addr_10, 
        IM_addr_9, IM_addr_8, IM_addr_7, IM_addr_6, IM_addr_5, IM_addr_4, 
        IM_addr_3, IM_addr_2, IM_addr_1, IM_addr_0, nrst, ip_r_req, ip_c_ack, 
        ip_complete, Ctrl__IFinst___Regs_1__ro, ip_local, ip_not_local, 
        IM_complete_latched, IM_read_data_mem_31, IM_read_data_mem_30, 
        IM_read_data_mem_29, IM_read_data_mem_28, IM_read_data_mem_27, 
        IM_read_data_mem_26, IM_read_data_mem_25, IM_read_data_mem_24, 
        IM_read_data_mem_23, IM_read_data_mem_22, IM_read_data_mem_21, 
        IM_read_data_mem_20, IM_read_data_mem_19, IM_read_data_mem_18, 
        IM_read_data_mem_17, IM_read_data_mem_16, IM_read_data_mem_15, 
        IM_read_data_mem_14, IM_read_data_mem_13, IM_read_data_mem_12, 
        IM_read_data_mem_11, IM_read_data_mem_10, IM_read_data_mem_9, 
        IM_read_data_mem_8, IM_read_data_mem_7, IM_read_data_mem_6, 
        IM_read_data_mem_5, IM_read_data_mem_4, IM_read_data_mem_3, 
        IM_read_data_mem_2, IM_read_data_mem_1, IM_read_data_mem_0, 
        IM_read_data_mem_latched_31, IM_read_data_mem_latched_30, 
        IM_read_data_mem_latched_29, IM_read_data_mem_latched_28, 
        IM_read_data_mem_latched_27, IM_read_data_mem_latched_26, 
        IM_read_data_mem_latched_25, IM_read_data_mem_latched_24, 
        IM_read_data_mem_latched_23, IM_read_data_mem_latched_22, 
        IM_read_data_mem_latched_21, IM_read_data_mem_latched_20, 
        IM_read_data_mem_latched_19, IM_read_data_mem_latched_18, 
        IM_read_data_mem_latched_17, IM_read_data_mem_latched_16, 
        IM_read_data_mem_latched_15, IM_read_data_mem_latched_14, 
        IM_read_data_mem_latched_13, IM_read_data_mem_latched_12, 
        IM_read_data_mem_latched_11, IM_read_data_mem_latched_10, 
        IM_read_data_mem_latched_9, IM_read_data_mem_latched_8, 
        IM_read_data_mem_latched_7, IM_read_data_mem_latched_6, 
        IM_read_data_mem_latched_5, IM_read_data_mem_latched_4, 
        IM_read_data_mem_latched_3, IM_read_data_mem_latched_2, 
        IM_read_data_mem_latched_1, IM_read_data_mem_latched_0, ip_r_dat_31, 
        ip_r_dat_30, ip_r_dat_29, ip_r_dat_28, ip_r_dat_27, ip_r_dat_26, 
        ip_r_dat_25, ip_r_dat_24, ip_r_dat_23, ip_r_dat_22, ip_r_dat_21, 
        ip_r_dat_20, ip_r_dat_19, ip_r_dat_18, ip_r_dat_17, ip_r_dat_16, 
        ip_r_dat_15, ip_r_dat_14, ip_r_dat_13, ip_r_dat_12, ip_r_dat_11, 
        ip_r_dat_10, ip_r_dat_9, ip_r_dat_8, ip_r_dat_7, ip_r_dat_6, 
        ip_r_dat_5, ip_r_dat_4, ip_r_dat_3, ip_r_dat_2, ip_r_dat_1, ip_r_dat_0, 
        IM_read_data_31, IM_read_data_30, IM_read_data_29, IM_read_data_28, 
        IM_read_data_27, IM_read_data_26, IM_read_data_25, IM_read_data_24, 
        IM_read_data_23, IM_read_data_22, IM_read_data_21, IM_read_data_20, 
        IM_read_data_19, IM_read_data_18, IM_read_data_17, IM_read_data_16, 
        IM_read_data_15, IM_read_data_14, IM_read_data_13, IM_read_data_12, 
        IM_read_data_11, IM_read_data_10, IM_read_data_9, IM_read_data_8, 
        IM_read_data_7, IM_read_data_6, IM_read_data_5, IM_read_data_4, 
        IM_read_data_3, IM_read_data_2, IM_read_data_1, IM_read_data_0, 
        Ctrl__IFinst___Regs_1__ai, ip_r_ack, _36_net_, IM_complete, 
        im_grant_local_d, Ctrl__IFinst___Regs_1__ri, dp_r_req, dp_c_ack, 
        dp_complete, DM_addr_CPU_31, DM_addr_CPU_30, DM_addr_CPU_29, 
        DM_addr_CPU_28, DM_addr_CPU_27, DM_addr_CPU_26, DM_addr_CPU_25, 
        DM_addr_CPU_24, DM_addr_CPU_23, DM_addr_CPU_22, DM_addr_CPU_21, 
        DM_addr_CPU_20, DM_addr_CPU_19, DM_addr_CPU_18, DM_addr_CPU_17, 
        DM_addr_CPU_16, DM_addr_CPU_15, DM_addr_CPU_14, DM_addr_CPU_13, 
        DM_addr_CPU_12, DM_addr_CPU_11, DM_addr_CPU_10, DM_addr_CPU_9, 
        DM_addr_CPU_8, DM_addr_CPU_7, DM_addr_CPU_6, DM_addr_CPU_5, 
        DM_addr_CPU_4, DM_addr_CPU_3, DM_addr_CPU_2, DM_addr_CPU_1, 
        DM_addr_CPU_0, Ctrl__EXinst___Regs_1__ro, DM_read, DM_write, dp_local, 
        dp_not_local, mask_to_mem_3, mask_to_mem_2, mask_to_mem_1, 
        mask_to_mem_0, DM_write_data_MIF_31, DM_write_data_MIF_30, 
        DM_write_data_MIF_29, DM_write_data_MIF_28, DM_write_data_MIF_27, 
        DM_write_data_MIF_26, DM_write_data_MIF_25, DM_write_data_MIF_24, 
        DM_write_data_MIF_23, DM_write_data_MIF_22, DM_write_data_MIF_21, 
        DM_write_data_MIF_20, DM_write_data_MIF_19, DM_write_data_MIF_18, 
        DM_write_data_MIF_17, DM_write_data_MIF_16, DM_write_data_MIF_15, 
        DM_write_data_MIF_14, DM_write_data_MIF_13, DM_write_data_MIF_12, 
        DM_write_data_MIF_11, DM_write_data_MIF_10, DM_write_data_MIF_9, 
        DM_write_data_MIF_8, DM_write_data_MIF_7, DM_write_data_MIF_6, 
        DM_write_data_MIF_5, DM_write_data_MIF_4, DM_write_data_MIF_3, 
        DM_write_data_MIF_2, DM_write_data_MIF_1, DM_write_data_MIF_0, 
        DM_complete_latched, DM_read_data_mem_31, DM_read_data_mem_30, 
        DM_read_data_mem_29, DM_read_data_mem_28, DM_read_data_mem_27, 
        DM_read_data_mem_26, DM_read_data_mem_25, DM_read_data_mem_24, 
        DM_read_data_mem_23, DM_read_data_mem_22, DM_read_data_mem_21, 
        DM_read_data_mem_20, DM_read_data_mem_19, DM_read_data_mem_18, 
        DM_read_data_mem_17, DM_read_data_mem_16, DM_read_data_mem_15, 
        DM_read_data_mem_14, DM_read_data_mem_13, DM_read_data_mem_12, 
        DM_read_data_mem_11, DM_read_data_mem_10, DM_read_data_mem_9, 
        DM_read_data_mem_8, DM_read_data_mem_7, DM_read_data_mem_6, 
        DM_read_data_mem_5, DM_read_data_mem_4, DM_read_data_mem_3, 
        DM_read_data_mem_2, DM_read_data_mem_1, DM_read_data_mem_0, 
        DM_read_data_mem_latched_31, DM_read_data_mem_latched_30, 
        DM_read_data_mem_latched_29, DM_read_data_mem_latched_28, 
        DM_read_data_mem_latched_27, DM_read_data_mem_latched_26, 
        DM_read_data_mem_latched_25, DM_read_data_mem_latched_24, 
        DM_read_data_mem_latched_23, DM_read_data_mem_latched_22, 
        DM_read_data_mem_latched_21, DM_read_data_mem_latched_20, 
        DM_read_data_mem_latched_19, DM_read_data_mem_latched_18, 
        DM_read_data_mem_latched_17, DM_read_data_mem_latched_16, 
        DM_read_data_mem_latched_15, DM_read_data_mem_latched_14, 
        DM_read_data_mem_latched_13, DM_read_data_mem_latched_12, 
        DM_read_data_mem_latched_11, DM_read_data_mem_latched_10, 
        DM_read_data_mem_latched_9, DM_read_data_mem_latched_8, 
        DM_read_data_mem_latched_7, DM_read_data_mem_latched_6, 
        DM_read_data_mem_latched_5, DM_read_data_mem_latched_4, 
        DM_read_data_mem_latched_3, DM_read_data_mem_latched_2, 
        DM_read_data_mem_latched_1, DM_read_data_mem_latched_0, dp_r_dat_31, 
        dp_r_dat_30, dp_r_dat_29, dp_r_dat_28, dp_r_dat_27, dp_r_dat_26, 
        dp_r_dat_25, dp_r_dat_24, dp_r_dat_23, dp_r_dat_22, dp_r_dat_21, 
        dp_r_dat_20, dp_r_dat_19, dp_r_dat_18, dp_r_dat_17, dp_r_dat_16, 
        dp_r_dat_15, dp_r_dat_14, dp_r_dat_13, dp_r_dat_12, dp_r_dat_11, 
        dp_r_dat_10, dp_r_dat_9, dp_r_dat_8, dp_r_dat_7, dp_r_dat_6, 
        dp_r_dat_5, dp_r_dat_4, dp_r_dat_3, dp_r_dat_2, dp_r_dat_1, dp_r_dat_0, 
        Ctrl__MEMinst___Regs_1__ai, dp_r_ack, _37_net_, DM_complete, 
        dm_grant_local_d, Ctrl__MEMinst___Regs_1__ri, im_c_req, _38_net_, 
        im_decup, im_r_ack, im_grant_local, _39_net_, im_grant_chain, _40_net_, 
        im_grant_chain_d, _41_net_, N315, im_c_we, im_c_sel_latched_3, 
        im_c_sel_latched_2, im_c_sel_latched_1, im_c_sel_latched_0, 
        IM_mask_oe_3, IM_mask_oe_2, IM_mask_oe_1, IM_mask_oe_0, im_c_sel_3, 
        im_c_sel_2, im_c_sel_1, im_c_sel_0, IM_mask_we_3, IM_mask_we_2, 
        IM_mask_we_1, IM_mask_we_0, im_c_adr_10, im_c_adr_9, im_c_adr_8, 
        im_c_adr_7, im_c_adr_6, im_c_adr_5, im_c_adr_4, im_c_adr_3, im_c_adr_2, 
        im_c_dat_31, im_c_dat_30, im_c_dat_29, im_c_dat_28, im_c_dat_27, 
        im_c_dat_26, im_c_dat_25, im_c_dat_24, im_c_dat_23, im_c_dat_22, 
        im_c_dat_21, im_c_dat_20, im_c_dat_19, im_c_dat_18, im_c_dat_17, 
        im_c_dat_16, im_c_dat_15, im_c_dat_14, im_c_dat_13, im_c_dat_12, 
        im_c_dat_11, im_c_dat_10, im_c_dat_9, im_c_dat_8, im_c_dat_7, 
        im_c_dat_6, im_c_dat_5, im_c_dat_4, im_c_dat_3, im_c_dat_2, im_c_dat_1, 
        im_c_dat_0, im_c_mult_latched, im_c_ts_latched_2, im_c_ts_latched_1, 
        im_c_ts_latched_0, im_c_mult, im_c_ts_2, im_c_ts_1, im_c_ts_0, 
        IM_start, sram_lat_select_1, sram_lat_select_0, im_r_req, dm_c_req, 
        _42_net_, dm_decup, dm_r_ack, _43_net_, dm_grant_local, dm_grant_chain, 
        N597, _44_net_, _45_net_, dm_grant_chain_d, dm_c_we, 
        dm_c_sel_latched_3, dm_c_sel_latched_2, dm_c_sel_latched_1, 
        dm_c_sel_latched_0, DM_mask_oe_3, DM_mask_oe_2, DM_mask_oe_1, 
        DM_mask_oe_0, dm_c_sel_3, dm_c_sel_2, dm_c_sel_1, dm_c_sel_0, 
        DM_mask_we_3, DM_mask_we_2, DM_mask_we_1, DM_mask_we_0, dm_c_adr_10, 
        dm_c_adr_9, dm_c_adr_8, dm_c_adr_7, dm_c_adr_6, dm_c_adr_5, dm_c_adr_4, 
        dm_c_adr_3, dm_c_adr_2, DM_addr_MEM_10, DM_addr_MEM_9, DM_addr_MEM_8, 
        DM_addr_MEM_7, DM_addr_MEM_6, DM_addr_MEM_5, DM_addr_MEM_4, 
        DM_addr_MEM_3, DM_addr_MEM_2, dm_c_dat_31, dm_c_dat_30, dm_c_dat_29, 
        dm_c_dat_28, dm_c_dat_27, dm_c_dat_26, dm_c_dat_25, dm_c_dat_24, 
        dm_c_dat_23, dm_c_dat_22, dm_c_dat_21, dm_c_dat_20, dm_c_dat_19, 
        dm_c_dat_18, dm_c_dat_17, dm_c_dat_16, dm_c_dat_15, dm_c_dat_14, 
        dm_c_dat_13, dm_c_dat_12, dm_c_dat_11, dm_c_dat_10, dm_c_dat_9, 
        dm_c_dat_8, dm_c_dat_7, dm_c_dat_6, dm_c_dat_5, dm_c_dat_4, dm_c_dat_3, 
        dm_c_dat_2, dm_c_dat_1, dm_c_dat_0, dm_c_mult_latched, 
        dm_c_ts_latched_2, dm_c_ts_latched_1, dm_c_ts_latched_0, dm_c_mult, 
        dm_c_ts_2, dm_c_ts_1, dm_c_ts_0, DM_start, dm_r_req, data_out_load_31, 
        data_out_load_30, data_out_load_29, data_out_load_28, data_out_load_27, 
        data_out_load_26, data_out_load_25, data_out_load_24, data_out_load_23, 
        data_out_load_22, data_out_load_21, data_out_load_20, data_out_load_19, 
        data_out_load_18, data_out_load_17, data_out_load_16, data_out_load_15, 
        data_out_load_14, data_out_load_13, data_out_load_12, data_out_load_11, 
        data_out_load_10, data_out_load_9, data_out_load_8, data_out_load_7, 
        data_out_load_6, data_out_load_5, data_out_load_4, data_out_load_3, 
        data_out_load_2, data_out_load_1, data_out_load_0, 
        IM_write_data_mem_31, IM_write_data_mem_30, IM_write_data_mem_29, 
        IM_write_data_mem_28, IM_write_data_mem_27, IM_write_data_mem_26, 
        IM_write_data_mem_25, IM_write_data_mem_24, IM_write_data_mem_23, 
        IM_write_data_mem_22, IM_write_data_mem_21, IM_write_data_mem_20, 
        IM_write_data_mem_19, IM_write_data_mem_18, IM_write_data_mem_17, 
        IM_write_data_mem_16, IM_write_data_mem_15, IM_write_data_mem_14, 
        IM_write_data_mem_13, IM_write_data_mem_12, IM_write_data_mem_11, 
        IM_write_data_mem_10, IM_write_data_mem_9, IM_write_data_mem_8, 
        IM_write_data_mem_7, IM_write_data_mem_6, IM_write_data_mem_5, 
        IM_write_data_mem_4, IM_write_data_mem_3, IM_write_data_mem_2, 
        IM_write_data_mem_1, IM_write_data_mem_0, DM_write_data_mem_31, 
        DM_write_data_mem_30, DM_write_data_mem_29, DM_write_data_mem_28, 
        DM_write_data_mem_27, DM_write_data_mem_26, DM_write_data_mem_25, 
        DM_write_data_mem_24, DM_write_data_mem_23, DM_write_data_mem_22, 
        DM_write_data_mem_21, DM_write_data_mem_20, DM_write_data_mem_19, 
        DM_write_data_mem_18, DM_write_data_mem_17, DM_write_data_mem_16, 
        DM_write_data_mem_15, DM_write_data_mem_14, DM_write_data_mem_13, 
        DM_write_data_mem_12, DM_write_data_mem_11, DM_write_data_mem_10, 
        DM_write_data_mem_9, DM_write_data_mem_8, DM_write_data_mem_7, 
        DM_write_data_mem_6, DM_write_data_mem_5, DM_write_data_mem_4, 
        DM_write_data_mem_3, DM_write_data_mem_2, DM_write_data_mem_1, 
        DM_write_data_mem_0, addr_out_load_10, addr_out_load_9, 
        addr_out_load_8, addr_out_load_7, addr_out_load_6, addr_out_load_5, 
        addr_out_load_4, addr_out_load_3, addr_out_load_2, IM_addr_MEM_mem_10, 
        IM_addr_MEM_mem_9, IM_addr_MEM_mem_8, IM_addr_MEM_mem_7, 
        IM_addr_MEM_mem_6, IM_addr_MEM_mem_5, IM_addr_MEM_mem_4, 
        IM_addr_MEM_mem_3, IM_addr_MEM_mem_2, DM_addr_MEM_mem_10, 
        DM_addr_MEM_mem_9, DM_addr_MEM_mem_8, DM_addr_MEM_mem_7, 
        DM_addr_MEM_mem_6, DM_addr_MEM_mem_5, DM_addr_MEM_mem_4, 
        DM_addr_MEM_mem_3, DM_addr_MEM_mem_2, 
        Ctrl__MEMinst___Regs_1__delay_mux_sel_1, 
        Ctrl__MEMinst___Regs_1__delay_mux_sel_0, 
        Ctrl__EXinst___Regs_1__delay_mux_sel_1, 
        Ctrl__EXinst___Regs_1__delay_mux_sel_0, 
        Ctrl__IDinst___Regs_1__delay_mux_sel_1, 
        Ctrl__IDinst___Regs_1__delay_mux_sel_0, 
        Ctrl__IFinst___Regs_1__delay_mux_sel_1, 
        Ctrl__IFinst___Regs_1__delay_mux_sel_0, force_bare, 
        DM_read_data_CPU_31, DM_read_data_CPU_30, DM_read_data_CPU_29, 
        DM_read_data_CPU_28, DM_read_data_CPU_27, DM_read_data_CPU_26, 
        DM_read_data_CPU_25, DM_read_data_CPU_24, DM_read_data_CPU_23, 
        DM_read_data_CPU_22, DM_read_data_CPU_21, DM_read_data_CPU_20, 
        DM_read_data_CPU_19, DM_read_data_CPU_18, DM_read_data_CPU_17, 
        DM_read_data_CPU_16, DM_read_data_CPU_15, DM_read_data_CPU_14, 
        DM_read_data_CPU_13, DM_read_data_CPU_12, DM_read_data_CPU_11, 
        DM_read_data_CPU_10, DM_read_data_CPU_9, DM_read_data_CPU_8, 
        DM_read_data_CPU_7, DM_read_data_CPU_6, DM_read_data_CPU_5, 
        DM_read_data_CPU_4, DM_read_data_CPU_3, DM_read_data_CPU_2, 
        DM_read_data_CPU_1, DM_read_data_CPU_0, DM_write_data_CPU_31, 
        DM_write_data_CPU_30, DM_write_data_CPU_29, DM_write_data_CPU_28, 
        DM_write_data_CPU_27, DM_write_data_CPU_26, DM_write_data_CPU_25, 
        DM_write_data_CPU_24, DM_write_data_CPU_23, DM_write_data_CPU_22, 
        DM_write_data_CPU_21, DM_write_data_CPU_20, DM_write_data_CPU_19, 
        DM_write_data_CPU_18, DM_write_data_CPU_17, DM_write_data_CPU_16, 
        DM_write_data_CPU_15, DM_write_data_CPU_14, DM_write_data_CPU_13, 
        DM_write_data_CPU_12, DM_write_data_CPU_11, DM_write_data_CPU_10, 
        DM_write_data_CPU_9, DM_write_data_CPU_8, DM_write_data_CPU_7, 
        DM_write_data_CPU_6, DM_write_data_CPU_5, DM_write_data_CPU_4, 
        DM_write_data_CPU_3, DM_write_data_CPU_2, DM_write_data_CPU_1, 
        DM_write_data_CPU_0, byte0, word, data_in_to_sh_reg_31, 
        data_in_to_sh_reg_30, data_in_to_sh_reg_29, data_in_to_sh_reg_28, 
        data_in_to_sh_reg_27, data_in_to_sh_reg_26, data_in_to_sh_reg_25, 
        data_in_to_sh_reg_24, data_in_to_sh_reg_23, data_in_to_sh_reg_22, 
        data_in_to_sh_reg_21, data_in_to_sh_reg_20, data_in_to_sh_reg_19, 
        data_in_to_sh_reg_18, data_in_to_sh_reg_17, data_in_to_sh_reg_16, 
        data_in_to_sh_reg_15, data_in_to_sh_reg_14, data_in_to_sh_reg_13, 
        data_in_to_sh_reg_12, data_in_to_sh_reg_11, data_in_to_sh_reg_10, 
        data_in_to_sh_reg_9, data_in_to_sh_reg_8, data_in_to_sh_reg_7, 
        data_in_to_sh_reg_6, data_in_to_sh_reg_5, data_in_to_sh_reg_4, 
        data_in_to_sh_reg_3, data_in_to_sh_reg_2, data_in_to_sh_reg_1, 
        data_in_to_sh_reg_0, data_write_load, data_write_load_im, 
        data_write_load_dm, N1107, IMem_clk, DMem_clk, N1429, N1431, n37, n40, 
        n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, 
        n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, 
        n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, 
        n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, 
        n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, 
        n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, 
        n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, 
        n155, n156, n157, n158, n159, n160, n39, n38;
    wire SYNOPSYS_UNCONNECTED_1 , SYNOPSYS_UNCONNECTED_2 , 
	SYNOPSYS_UNCONNECTED_3 , SYNOPSYS_UNCONNECTED_4 , SYNOPSYS_UNCONNECTED_5 , 
	SYNOPSYS_UNCONNECTED_6 , SYNOPSYS_UNCONNECTED_7 , SYNOPSYS_UNCONNECTED_8 , 
	SYNOPSYS_UNCONNECTED_9 , SYNOPSYS_UNCONNECTED_10 , SYNOPSYS_UNCONNECTED_11 , 
	SYNOPSYS_UNCONNECTED_12 , SYNOPSYS_UNCONNECTED_13 , SYNOPSYS_UNCONNECTED_14 , 
	SYNOPSYS_UNCONNECTED_15 , SYNOPSYS_UNCONNECTED_16 , SYNOPSYS_UNCONNECTED_17 , 
	SYNOPSYS_UNCONNECTED_18 , SYNOPSYS_UNCONNECTED_19 , SYNOPSYS_UNCONNECTED_20 , 
	SYNOPSYS_UNCONNECTED_21 , SYNOPSYS_UNCONNECTED_22 , SYNOPSYS_UNCONNECTED_23 , 
	SYNOPSYS_UNCONNECTED_24 , SYNOPSYS_UNCONNECTED_25 , SYNOPSYS_UNCONNECTED_26 , 
	SYNOPSYS_UNCONNECTED_27 , SYNOPSYS_UNCONNECTED_28 , SYNOPSYS_UNCONNECTED_29 , 
	SYNOPSYS_UNCONNECTED_30 , SYNOPSYS_UNCONNECTED_31 , SYNOPSYS_UNCONNECTED_32 , 
	SYNOPSYS_UNCONNECTED_33 , SYNOPSYS_UNCONNECTED_34 , SYNOPSYS_UNCONNECTED_35 , 
	SYNOPSYS_UNCONNECTED_36 , SYNOPSYS_UNCONNECTED_37 , SYNOPSYS_UNCONNECTED_38 , 
	SYNOPSYS_UNCONNECTED_39 , SYNOPSYS_UNCONNECTED_40 , SYNOPSYS_UNCONNECTED_41 , 
	SYNOPSYS_UNCONNECTED_42 , SYNOPSYS_UNCONNECTED_43 , SYNOPSYS_UNCONNECTED_44 , 
	SYNOPSYS_UNCONNECTED_45 , SYNOPSYS_UNCONNECTED_46 , SYNOPSYS_UNCONNECTED_47 , 
	SYNOPSYS_UNCONNECTED_48 ;
    inbuf3_16 stop_fetch_pad_ ( .di(STOP_fetch), .pad(STOP_FETCH_PAD) );
    inbuf3_16 reset_ctrl_pad_ ( .di(reset_ctrl), .pad(reset_ctrl_PAD) );
    inbuf3_16 freeze_pad_ ( .di(FREEZE), .pad(FREEZE_PAD) );
    inbuf3_16 memory_load_enable_pad_ ( .di(memory_load_enable), .pad(
        memory_load_enable_PAD) );
    inbuf3_16 scan_in_pad_ ( .di(scan_in), .pad(scan_in_PAD) );
    iobuf3_16_12 scan_out_pad_ ( .pad(scan_out_PAD), .\do (scan_out), .en(1'b1
        ) );
    inbuf3_16 shift_clk_pad_ ( .di(shift_clk), .pad(shift_clk_PAD) );
    inbuf3_16 read_pad_ ( .di(read), .pad(read_PAD) );
    inbuf3_16 inst_ram_load_pad_ ( .di(inst_ram_load), .pad(inst_ram_load_PAD)
         );
    inbuf3_16 del_scan_en_pad_ ( .di(del_scan_en), .pad(del_scan_en_PAD) );
    inbuf3_16 del_scan_in_pad_ ( .di(del_scan_in), .pad(del_scan_in_PAD) );
    inbuf3_16 reset_DLX_d_pad_ ( .di(reset_DLX_d), .pad(reset_DLX_d_PAD) );
    inbuf3_16 reset_DLX_c_pad_ ( .di(reset_DLX_c), .pad(reset_DLX_c_PAD) );
    inbuf3_16 sync_async_pad_ ( .di(N1107), .pad(sync_async_PAD) );
    inbuf3_16 int_pad_ ( .di(INT), .pad(INT_PAD) );
    inbuf3_16 test_si_DLX_pad_ ( .di(test_si_DLX), .pad(test_si_DLX_PAD) );
    inbuf3_16 test_se_pad_ ( .di(test_se), .pad(test_se_PAD) );
    inbuf3_16 global_g1_pad_ ( .di(global_g1), .pad(global_g1_PAD) );
    inbuf3_16 global_g2_pad_ ( .di(global_g2), .pad(global_g2_PAD) );
    inbuf3_16 r_BC_pad_0 ( .di(r_BC_0), .pad(r_BC_PAD[0]) );
    inbuf3_16 r_BC_pad_1 ( .di(r_BC_1), .pad(r_BC_PAD[1]) );
    inbuf3_16 r_BC_pad_2 ( .di(r_BC_2), .pad(r_BC_PAD[2]) );
    inbuf3_16 r_BC_pad_3 ( .di(r_BC_3), .pad(r_BC_PAD[3]) );
    inbuf3_16 r_BC_pad_4 ( .di(r_BC_4), .pad(r_BC_PAD[4]) );
    iobuf3_16_12 r_BC_ack_pad_ ( .pad(r_BC_ack_PAD), .\do (r_BC_ack), .en(1'b1
        ) );
    inbuf3_16 c_BC_ack_pad_ ( .di(c_BC_ack), .pad(c_BC_ack_PAD) );
    iobuf3_16_12 c_BC_pad_0 ( .pad(c_BC_PAD[0]), .\do (c_BC_0), .en(1'b1) );
    iobuf3_16_12 c_BC_pad_1 ( .pad(c_BC_PAD[1]), .\do (c_BC_1), .en(1'b1) );
    iobuf3_16_12 c_BC_pad_2 ( .pad(c_BC_PAD[2]), .\do (c_BC_2), .en(1'b1) );
    iobuf3_16_12 c_BC_pad_3 ( .pad(c_BC_PAD[3]), .\do (c_BC_3), .en(1'b1) );
    iobuf3_16_12 c_BC_pad_4 ( .pad(c_BC_PAD[4]), .\do (c_BC_4), .en(1'b1) );
    inbuf3_16 ei_c_req_pad_ ( .di(ei_c_req), .pad(ei_c_req_PAD) );
    inbuf3_16 ei_c_we_pad_ ( .di(ei_c_we), .pad(ei_c_we_PAD) );
    inbuf3_16 ei_c_addr_pad_0 ( .di(ei_c_addr_0), .pad(ei_c_addr_PAD[0]) );
    inbuf3_16 ei_c_addr_pad_1 ( .di(ei_c_addr_1), .pad(ei_c_addr_PAD[1]) );
    inbuf3_16 ei_c_addr_pad_2 ( .di(ei_c_addr_2), .pad(ei_c_addr_PAD[2]) );
    inbuf3_16 ei_c_addr_pad_3 ( .di(ei_c_addr_3), .pad(ei_c_addr_PAD[3]) );
    inbuf3_16 ei_c_addr_pad_4 ( .di(ei_c_addr_4), .pad(ei_c_addr_PAD[4]) );
    inbuf3_16 ei_c_addr_pad_5 ( .di(ei_c_addr_5), .pad(ei_c_addr_PAD[5]) );
    inbuf3_16 ei_c_addr_pad_6 ( .di(ei_c_addr_6), .pad(ei_c_addr_PAD[6]) );
    inbuf3_16 ei_c_addr_pad_7 ( .di(ei_c_addr_7), .pad(ei_c_addr_PAD[7]) );
    inbuf3_16 ei_c_addr_pad_8 ( .di(ei_c_addr_8), .pad(ei_c_addr_PAD[8]) );
    inbuf3_16 ei_c_addr_pad_9 ( .di(ei_c_addr_9), .pad(ei_c_addr_PAD[9]) );
    inbuf3_16 ei_c_addr_pad_10 ( .di(ei_c_addr_10), .pad(ei_c_addr_PAD[10]) );
    iobuf3_16_12 ei_c_ack_pad_ ( .pad(ei_c_ack_PAD), .\do (ei_c_ack), .en(1'b1
        ) );
    iobuf3_16_12 ei_r_req_pad_ ( .pad(ei_r_req_PAD), .\do (ei_r_req), .en(1'b1
        ) );
    iobuf3_16_12 ei_data_inout_pad_0 ( .di(ei_data_in_0), .pad(
        ei_data_inout_PAD[0]), .\do (ei_data_out_0), .en(_17_net_) );
    iobuf3_16_12 ei_data_inout_pad_1 ( .di(ei_data_in_1), .pad(
        ei_data_inout_PAD[1]), .\do (ei_data_out_1), .en(_17_net_) );
    iobuf3_16_12 ei_data_inout_pad_2 ( .di(ei_data_in_2), .pad(
        ei_data_inout_PAD[2]), .\do (ei_data_out_2), .en(_17_net_) );
    iobuf3_16_12 ei_data_inout_pad_3 ( .di(ei_data_in_3), .pad(
        ei_data_inout_PAD[3]), .\do (ei_data_out_3), .en(_17_net_) );
    iobuf3_16_12 ei_data_inout_pad_4 ( .di(ei_data_in_4), .pad(
        ei_data_inout_PAD[4]), .\do (ei_data_out_4), .en(_17_net_) );
    iobuf3_16_12 ei_data_inout_pad_5 ( .di(ei_data_in_5), .pad(
        ei_data_inout_PAD[5]), .\do (ei_data_out_5), .en(_17_net_) );
    iobuf3_16_12 ei_data_inout_pad_6 ( .di(ei_data_in_6), .pad(
        ei_data_inout_PAD[6]), .\do (ei_data_out_6), .en(_17_net_) );
    iobuf3_16_12 ei_data_inout_pad_7 ( .di(ei_data_in_7), .pad(
        ei_data_inout_PAD[7]), .\do (ei_data_out_7), .en(_17_net_) );
    inbuf3_16 ei_r_ack_pad_ ( .di(ei_r_ack), .pad(ei_r_ack_PAD) );
    inbuf3_16 wish_ack_i_pad ( .di(wish_ack_i), .pad(wish_ack_i_PAD) );
    inbuf3_16 wish_clk_pad ( .di(wish_clk), .pad(wish_clk_PAD) );
    iobuf3_16_12 wish_stb_cyc_o_pad ( .pad(wish_stb_cyc_o_PAD), .\do (
        wish_stb_cyc_o), .en(1'b1) );
    iobuf3_16_12 wish_we_o_pad ( .pad(wish_we_o_PAD), .\do (n107), .en(1'b1)
         );
    iobuf3_16_12 wish_adr_o_pad_0 ( .pad(wish_adr_o_PAD[0]), .\do (
        wish_adr_o_0), .en(1'b1) );
    iobuf3_16_12 wish_adr_o_pad_1 ( .pad(wish_adr_o_PAD[1]), .\do (
        wish_adr_o_1), .en(1'b1) );
    iobuf3_16_12 wish_adr_o_pad_2 ( .pad(wish_adr_o_PAD[2]), .\do (
        wish_adr_o_2), .en(1'b1) );
    iobuf3_16_12 wish_adr_o_pad_3 ( .pad(wish_adr_o_PAD[3]), .\do (
        wish_adr_o_3), .en(1'b1) );
    iobuf3_16_12 wish_adr_o_pad_4 ( .pad(wish_adr_o_PAD[4]), .\do (
        wish_adr_o_4), .en(1'b1) );
    iobuf3_16_12 wish_adr_o_pad_5 ( .pad(wish_adr_o_PAD[5]), .\do (
        wish_adr_o_5), .en(1'b1) );
    iobuf3_16_12 wish_adr_o_pad_6 ( .pad(wish_adr_o_PAD[6]), .\do (
        wish_adr_o_6), .en(1'b1) );
    iobuf3_16_12 wish_adr_o_pad_7 ( .pad(wish_adr_o_PAD[7]), .\do (
        wish_adr_o_7), .en(1'b1) );
    iobuf3_16_12 wish_adr_o_pad_8 ( .pad(wish_adr_o_PAD[8]), .\do (
        wish_adr_o_8), .en(1'b1) );
    iobuf3_16_12 wish_adr_o_pad_9 ( .pad(wish_adr_o_PAD[9]), .\do (
        wish_adr_o_9), .en(1'b1) );
    iobuf3_16_12 wish_adr_o_pad_10 ( .pad(wish_adr_o_PAD[10]), .\do (
        wish_adr_o_10), .en(1'b1) );
    iobuf3_16_12 wish_adr_o_pad_11 ( .pad(wish_adr_o_PAD[11]), .\do (
        wish_adr_o_11), .en(1'b1) );
    iobuf3_16_12 wish_dat_io_pad_0 ( .di(wish_dat_i_0), .pad(wish_dat_io_PAD
        [0]), .\do (wish_dat_o_0), .en(wish_we_o) );
    iobuf3_16_12 wish_dat_io_pad_1 ( .di(wish_dat_i_1), .pad(wish_dat_io_PAD
        [1]), .\do (wish_dat_o_1), .en(n107) );
    iobuf3_16_12 wish_dat_io_pad_2 ( .di(wish_dat_i_2), .pad(wish_dat_io_PAD
        [2]), .\do (wish_dat_o_2), .en(n107) );
    iobuf3_16_12 wish_dat_io_pad_3 ( .di(wish_dat_i_3), .pad(wish_dat_io_PAD
        [3]), .\do (wish_dat_o_3), .en(n107) );
    iobuf3_16_12 wish_dat_io_pad_4 ( .di(wish_dat_i_4), .pad(wish_dat_io_PAD
        [4]), .\do (wish_dat_o_4), .en(n107) );
    iobuf3_16_12 wish_dat_io_pad_5 ( .di(wish_dat_i_5), .pad(wish_dat_io_PAD
        [5]), .\do (wish_dat_o_5), .en(n107) );
    iobuf3_16_12 wish_dat_io_pad_6 ( .di(wish_dat_i_6), .pad(wish_dat_io_PAD
        [6]), .\do (wish_dat_o_6), .en(n107) );
    iobuf3_16_12 wish_dat_io_pad_7 ( .di(wish_dat_i_7), .pad(wish_dat_io_PAD
        [7]), .\do (wish_dat_o_7), .en(n107) );
    iobuf3_16_12 wish_dat_io_pad_8 ( .di(wish_dat_i_8), .pad(wish_dat_io_PAD
        [8]), .\do (wish_dat_o_8), .en(n107) );
    iobuf3_16_12 wish_dat_io_pad_9 ( .di(wish_dat_i_9), .pad(wish_dat_io_PAD
        [9]), .\do (wish_dat_o_9), .en(n107) );
    iobuf3_16_12 wish_dat_io_pad_10 ( .di(wish_dat_i_10), .pad(wish_dat_io_PAD
        [10]), .\do (wish_dat_o_10), .en(n107) );
    iobuf3_16_12 wish_dat_io_pad_11 ( .di(wish_dat_i_11), .pad(wish_dat_io_PAD
        [11]), .\do (wish_dat_o_11), .en(n107) );
    iobuf3_16_12 wish_dat_io_pad_12 ( .di(wish_dat_i_12), .pad(wish_dat_io_PAD
        [12]), .\do (wish_dat_o_12), .en(n107) );
    iobuf3_16_12 wish_dat_io_pad_13 ( .di(wish_dat_i_13), .pad(wish_dat_io_PAD
        [13]), .\do (wish_dat_o_13), .en(n107) );
    iobuf3_16_12 wish_dat_io_pad_14 ( .di(wish_dat_i_14), .pad(wish_dat_io_PAD
        [14]), .\do (wish_dat_o_14), .en(n107) );
    iobuf3_16_12 wish_dat_io_pad_15 ( .di(wish_dat_i_15), .pad(wish_dat_io_PAD
        [15]), .\do (wish_dat_o_15), .en(wish_we_o) );
    iobuf3_16_12 wish_dat_io_pad_16 ( .di(wish_dat_i_16), .pad(wish_dat_io_PAD
        [16]), .\do (wish_dat_o_16), .en(wish_we_o) );
    iobuf3_16_12 wish_dat_io_pad_17 ( .di(wish_dat_i_17), .pad(wish_dat_io_PAD
        [17]), .\do (wish_dat_o_17), .en(n107) );
    iobuf3_16_12 wish_dat_io_pad_18 ( .di(wish_dat_i_18), .pad(wish_dat_io_PAD
        [18]), .\do (wish_dat_o_18), .en(n107) );
    iobuf3_16_12 wish_dat_io_pad_19 ( .di(wish_dat_i_19), .pad(wish_dat_io_PAD
        [19]), .\do (wish_dat_o_19), .en(n107) );
    iobuf3_16_12 wish_dat_io_pad_20 ( .di(wish_dat_i_20), .pad(wish_dat_io_PAD
        [20]), .\do (wish_dat_o_20), .en(n107) );
    iobuf3_16_12 wish_dat_io_pad_21 ( .di(wish_dat_i_21), .pad(wish_dat_io_PAD
        [21]), .\do (wish_dat_o_21), .en(n107) );
    iobuf3_16_12 wish_dat_io_pad_22 ( .di(wish_dat_i_22), .pad(wish_dat_io_PAD
        [22]), .\do (wish_dat_o_22), .en(n107) );
    iobuf3_16_12 wish_dat_io_pad_23 ( .di(wish_dat_i_23), .pad(wish_dat_io_PAD
        [23]), .\do (wish_dat_o_23), .en(n107) );
    iobuf3_16_12 wish_dat_io_pad_24 ( .di(wish_dat_i_24), .pad(wish_dat_io_PAD
        [24]), .\do (wish_dat_o_24), .en(n107) );
    iobuf3_16_12 wish_dat_io_pad_25 ( .di(wish_dat_i_25), .pad(wish_dat_io_PAD
        [25]), .\do (wish_dat_o_25), .en(n107) );
    iobuf3_16_12 wish_dat_io_pad_26 ( .di(wish_dat_i_26), .pad(wish_dat_io_PAD
        [26]), .\do (wish_dat_o_26), .en(n107) );
    iobuf3_16_12 wish_dat_io_pad_27 ( .di(wish_dat_i_27), .pad(wish_dat_io_PAD
        [27]), .\do (wish_dat_o_27), .en(n107) );
    iobuf3_16_12 wish_dat_io_pad_28 ( .di(wish_dat_i_28), .pad(wish_dat_io_PAD
        [28]), .\do (wish_dat_o_28), .en(n107) );
    iobuf3_16_12 wish_dat_io_pad_29 ( .di(wish_dat_i_29), .pad(wish_dat_io_PAD
        [29]), .\do (wish_dat_o_29), .en(n107) );
    iobuf3_16_12 wish_dat_io_pad_30 ( .di(wish_dat_i_30), .pad(wish_dat_io_PAD
        [30]), .\do (wish_dat_o_30), .en(n107) );
    iobuf3_16_12 wish_dat_io_pad_31 ( .di(wish_dat_i_31), .pad(wish_dat_io_PAD
        [31]), .\do (wish_dat_o_31), .en(wish_we_o) );
    iobuf3_16_12 cli_pad_ ( .pad(CLI_PAD), .\do (CLI), .en(1'b1) );
    iobuf3_16_12 test_so_DLX_pad_ ( .pad(test_so_DLX_PAD), .\do (IM_addr_31), 
        .en(1'b1) );
    iobuf3_16_12 stuckAtVdd_pad_ ( .pad(stuckAtVdd_PAD), .\do (1'b1), .en(1'b1
        ) );
    dffn_1 sync1g2 ( .q(reset_DLX_d_ff1), .d(reset_DLX_d), .ckb(global_g2) );
    dffn_1 sync2g2 ( .q(reset_DLX_d_ff2), .d(reset_DLX_d_ff1), .ckb(global_g2)
         );
    dffp_1 sync1shift ( .q(reset_DLX_d_ff1_shift), .d(reset_DLX_d), .ck(
        shift_clk) );
    dffp_1 sync2shift ( .d(reset_DLX_d_ff1_shift), .ck(shift_clk) );
    C_gate2 sync_ip_complete ( .in1(ip_r_req), .in2(ip_c_ack), .out(
        ip_complete) );
    C_gate2 sync_im_complete ( .in1(ip_local), .in2(_36_net_), .out(
        IM_complete_latched) );
    C_gate2 sync_dp_complete ( .in1(dp_r_req), .in2(dp_c_ack), .out(
        dp_complete) );
    C_gate2 sync_dm_complete ( .in1(dp_local), .in2(_37_net_), .out(
        DM_complete_latched) );
    C_gate2 sync_im_decup ( .in1(im_c_req), .in2(_38_net_), .out(im_decup) );
    C_gate2 sync_dm_decup0 ( .in1(im_grant_local), .in2(_39_net_), .out(
        im_grant_local_d) );
    C_gate2 sync_dm_decup1 ( .in1(im_grant_chain), .in2(_40_net_), .out(
        im_grant_chain_d) );
    mutex arb_im0 ( .r1(_41_net_), .r2(im_decup), .g1(im_grant_local), .g2(
        im_grant_chain) );
    sram_latency sramlat_imem ( .in(IM_start), .out(IM_complete), .mux_sel({
        sram_lat_select_1, sram_lat_select_0}) );
    C_gate2 sync_dm_decup2 ( .in1(dm_c_req), .in2(_42_net_), .out(dm_decup) );
    mutex arb_im1 ( .r1(_43_net_), .r2(dm_decup), .g1(dm_grant_local), .g2(
        dm_grant_chain) );
    C_gate2 sync_dm_decup3 ( .in1(dm_grant_local), .in2(_44_net_), .out(
        dm_grant_local_d) );
    C_gate2 sync_dm_decup4 ( .in1(dm_grant_chain), .in2(_45_net_), .out(
        dm_grant_chain_d) );
    sram_latency sramlat_dmem ( .in(DM_start), .out(DM_complete), .mux_sel({
        sram_lat_select_1, sram_lat_select_0}) );
    delay_shifter delem_shift_reg ( .reset(reset_DLX_d), .enable(del_scan_en), 
        .shift_clk(shift_clk), .scan_in(del_scan_in), .par_out({
        Ctrl__MEMinst___Regs_1__delay_mux_sel_1, 
        Ctrl__MEMinst___Regs_1__delay_mux_sel_0, 
        Ctrl__EXinst___Regs_1__delay_mux_sel_1, 
        Ctrl__EXinst___Regs_1__delay_mux_sel_0, 
        Ctrl__IDinst___Regs_1__delay_mux_sel_1, 
        Ctrl__IDinst___Regs_1__delay_mux_sel_0, 
        Ctrl__IFinst___Regs_1__delay_mux_sel_1, 
        Ctrl__IFinst___Regs_1__delay_mux_sel_0, sram_lat_select_1, 
        sram_lat_select_0, force_bare}) );
    DLX_sync_desync_with_ctrls processor ( .DM_read_data({DM_read_data_CPU_31, 
        DM_read_data_CPU_30, DM_read_data_CPU_29, DM_read_data_CPU_28, 
        DM_read_data_CPU_27, DM_read_data_CPU_26, DM_read_data_CPU_25, 
        DM_read_data_CPU_24, DM_read_data_CPU_23, DM_read_data_CPU_22, 
        DM_read_data_CPU_21, DM_read_data_CPU_20, DM_read_data_CPU_19, 
        DM_read_data_CPU_18, DM_read_data_CPU_17, DM_read_data_CPU_16, 
        DM_read_data_CPU_15, DM_read_data_CPU_14, DM_read_data_CPU_13, 
        DM_read_data_CPU_12, DM_read_data_CPU_11, DM_read_data_CPU_10, 
        DM_read_data_CPU_9, DM_read_data_CPU_8, DM_read_data_CPU_7, 
        DM_read_data_CPU_6, DM_read_data_CPU_5, DM_read_data_CPU_4, 
        DM_read_data_CPU_3, DM_read_data_CPU_2, DM_read_data_CPU_1, 
        DM_read_data_CPU_0}), .DM_write_data({DM_write_data_CPU_31, 
        DM_write_data_CPU_30, DM_write_data_CPU_29, DM_write_data_CPU_28, 
        DM_write_data_CPU_27, DM_write_data_CPU_26, DM_write_data_CPU_25, 
        DM_write_data_CPU_24, DM_write_data_CPU_23, DM_write_data_CPU_22, 
        DM_write_data_CPU_21, DM_write_data_CPU_20, DM_write_data_CPU_19, 
        DM_write_data_CPU_18, DM_write_data_CPU_17, DM_write_data_CPU_16, 
        DM_write_data_CPU_15, DM_write_data_CPU_14, DM_write_data_CPU_13, 
        DM_write_data_CPU_12, DM_write_data_CPU_11, DM_write_data_CPU_10, 
        DM_write_data_CPU_9, DM_write_data_CPU_8, DM_write_data_CPU_7, 
        DM_write_data_CPU_6, DM_write_data_CPU_5, DM_write_data_CPU_4, 
        DM_write_data_CPU_3, DM_write_data_CPU_2, DM_write_data_CPU_1, 
        DM_write_data_CPU_0}), .DM_addr({DM_addr_CPU_31, DM_addr_CPU_30, 
        DM_addr_CPU_29, DM_addr_CPU_28, DM_addr_CPU_27, DM_addr_CPU_26, 
        DM_addr_CPU_25, DM_addr_CPU_24, DM_addr_CPU_23, DM_addr_CPU_22, 
        DM_addr_CPU_21, DM_addr_CPU_20, DM_addr_CPU_19, DM_addr_CPU_18, 
        DM_addr_CPU_17, DM_addr_CPU_16, DM_addr_CPU_15, DM_addr_CPU_14, 
        DM_addr_CPU_13, DM_addr_CPU_12, DM_addr_CPU_11, DM_addr_CPU_10, 
        DM_addr_CPU_9, DM_addr_CPU_8, DM_addr_CPU_7, DM_addr_CPU_6, 
        DM_addr_CPU_5, DM_addr_CPU_4, DM_addr_CPU_3, DM_addr_CPU_2, 
        DM_addr_CPU_1, DM_addr_CPU_0}), .DM_write(DM_write), .DM_read(DM_read), 
        .NPC({IM_addr_31, IM_addr_30, IM_addr_29, IM_addr_28, IM_addr_27, 
        IM_addr_26, IM_addr_25, IM_addr_24, IM_addr_23, IM_addr_22, IM_addr_21, 
        IM_addr_20, IM_addr_19, IM_addr_18, IM_addr_17, IM_addr_16, IM_addr_15, 
        IM_addr_14, IM_addr_13, IM_addr_12, IM_addr_11, IM_addr_10, IM_addr_9, 
        IM_addr_8, IM_addr_7, IM_addr_6, IM_addr_5, IM_addr_4, IM_addr_3, 
        IM_addr_2, IM_addr_1, IM_addr_0}), .reset(n103), .IR({IM_read_data_31, 
        IM_read_data_30, IM_read_data_29, IM_read_data_28, IM_read_data_27, 
        IM_read_data_26, IM_read_data_25, IM_read_data_24, IM_read_data_23, 
        IM_read_data_22, IM_read_data_21, IM_read_data_20, IM_read_data_19, 
        IM_read_data_18, IM_read_data_17, IM_read_data_16, IM_read_data_15, 
        IM_read_data_14, IM_read_data_13, IM_read_data_12, IM_read_data_11, 
        IM_read_data_10, IM_read_data_9, IM_read_data_8, IM_read_data_7, 
        IM_read_data_6, IM_read_data_5, IM_read_data_4, IM_read_data_3, 
        IM_read_data_2, IM_read_data_1, IM_read_data_0}), .byte0(byte0), 
        .word(word), .INT(INT), .CLI(CLI), .FREEZE(FREEZE), .test_si(
        test_si_DLX), .test_se(n120), .sync_sel(N1107), .global_g1(n106), 
        .global_g2(n116), .Ctrl__reset(reset_DLX_ctrl), 
        .Ctrl__IFinst___Regs_1__ri(Ctrl__IFinst___Regs_1__ri), 
        .Ctrl__IFinst___Regs_1__ai(Ctrl__IFinst___Regs_1__ai), 
        .Ctrl__MEMinst___Regs_1__ri(Ctrl__MEMinst___Regs_1__ri), 
        .Ctrl__MEMinst___Regs_1__ai(Ctrl__MEMinst___Regs_1__ai), 
        .Ctrl__EXinst___Regs_1__ro(Ctrl__EXinst___Regs_1__ro), 
        .Ctrl__EXinst___Regs_1__ao(Ctrl__MEMinst___Regs_1__ai), 
        .Ctrl__IFinst___Regs_1__ro(Ctrl__IFinst___Regs_1__ro), 
        .Ctrl__IFinst___Regs_1__ao(Ctrl__IFinst___Regs_1__ai), 
        .Ctrl__EXinst___Regs_1__delay_mux_sel({
        Ctrl__EXinst___Regs_1__delay_mux_sel_1, 
        Ctrl__EXinst___Regs_1__delay_mux_sel_0}), 
        .Ctrl__IDinst___Regs_1__delay_mux_sel({
        Ctrl__IDinst___Regs_1__delay_mux_sel_1, 
        Ctrl__IDinst___Regs_1__delay_mux_sel_0}), 
        .Ctrl__IFinst___Regs_1__delay_mux_sel({
        Ctrl__IFinst___Regs_1__delay_mux_sel_1, 
        Ctrl__IFinst___Regs_1__delay_mux_sel_0}), 
        .Ctrl__MEMinst___Regs_1__delay_mux_sel({
        Ctrl__MEMinst___Regs_1__delay_mux_sel_1, 
        Ctrl__MEMinst___Regs_1__delay_mux_sel_0}) );
    mem_if mem_iface ( .DM_addr_CPU({DM_addr_CPU_31, DM_addr_CPU_30, 
        DM_addr_CPU_29, DM_addr_CPU_28, DM_addr_CPU_27, DM_addr_CPU_26, 
        DM_addr_CPU_25, DM_addr_CPU_24, DM_addr_CPU_23, DM_addr_CPU_22, 
        DM_addr_CPU_21, DM_addr_CPU_20, DM_addr_CPU_19, DM_addr_CPU_18, 
        DM_addr_CPU_17, DM_addr_CPU_16, DM_addr_CPU_15, DM_addr_CPU_14, 
        DM_addr_CPU_13, DM_addr_CPU_12, DM_addr_CPU_11, DM_addr_CPU_10, 
        DM_addr_CPU_9, DM_addr_CPU_8, DM_addr_CPU_7, DM_addr_CPU_6, 
        DM_addr_CPU_5, DM_addr_CPU_4, DM_addr_CPU_3, DM_addr_CPU_2, 
        DM_addr_CPU_1, DM_addr_CPU_0}), .DM_read_data_CPU({DM_read_data_CPU_31, 
        DM_read_data_CPU_30, DM_read_data_CPU_29, DM_read_data_CPU_28, 
        DM_read_data_CPU_27, DM_read_data_CPU_26, DM_read_data_CPU_25, 
        DM_read_data_CPU_24, DM_read_data_CPU_23, DM_read_data_CPU_22, 
        DM_read_data_CPU_21, DM_read_data_CPU_20, DM_read_data_CPU_19, 
        DM_read_data_CPU_18, DM_read_data_CPU_17, DM_read_data_CPU_16, 
        DM_read_data_CPU_15, DM_read_data_CPU_14, DM_read_data_CPU_13, 
        DM_read_data_CPU_12, DM_read_data_CPU_11, DM_read_data_CPU_10, 
        DM_read_data_CPU_9, DM_read_data_CPU_8, DM_read_data_CPU_7, 
        DM_read_data_CPU_6, DM_read_data_CPU_5, DM_read_data_CPU_4, 
        DM_read_data_CPU_3, DM_read_data_CPU_2, DM_read_data_CPU_1, 
        DM_read_data_CPU_0}), .DM_write_data_CPU({DM_write_data_CPU_31, 
        DM_write_data_CPU_30, DM_write_data_CPU_29, DM_write_data_CPU_28, 
        DM_write_data_CPU_27, DM_write_data_CPU_26, DM_write_data_CPU_25, 
        DM_write_data_CPU_24, DM_write_data_CPU_23, DM_write_data_CPU_22, 
        DM_write_data_CPU_21, DM_write_data_CPU_20, DM_write_data_CPU_19, 
        DM_write_data_CPU_18, DM_write_data_CPU_17, DM_write_data_CPU_16, 
        DM_write_data_CPU_15, DM_write_data_CPU_14, DM_write_data_CPU_13, 
        DM_write_data_CPU_12, DM_write_data_CPU_11, DM_write_data_CPU_10, 
        DM_write_data_CPU_9, DM_write_data_CPU_8, DM_write_data_CPU_7, 
        DM_write_data_CPU_6, DM_write_data_CPU_5, DM_write_data_CPU_4, 
        DM_write_data_CPU_3, DM_write_data_CPU_2, DM_write_data_CPU_1, 
        DM_write_data_CPU_0}), .word(word), .\byte (byte0), .DM_addr_MEM({
        DM_addr_MEM_10, DM_addr_MEM_9, DM_addr_MEM_8, DM_addr_MEM_7, 
        DM_addr_MEM_6, DM_addr_MEM_5, DM_addr_MEM_4, DM_addr_MEM_3, 
        DM_addr_MEM_2}), .DM_read_data_MEM({n47, n48, n50, n51, n52, n53, n54, 
        n81, n82, n83, n84, n85, n87, n88, n89, n90, n91, n92, n93, n94, n95, 
        n96, n41, n42, n43, n44, n45, n46, n49, n86, n97, n98}), 
        .DM_write_data_MEM({DM_write_data_MIF_31, DM_write_data_MIF_30, 
        DM_write_data_MIF_29, DM_write_data_MIF_28, DM_write_data_MIF_27, 
        DM_write_data_MIF_26, DM_write_data_MIF_25, DM_write_data_MIF_24, 
        DM_write_data_MIF_23, DM_write_data_MIF_22, DM_write_data_MIF_21, 
        DM_write_data_MIF_20, DM_write_data_MIF_19, DM_write_data_MIF_18, 
        DM_write_data_MIF_17, DM_write_data_MIF_16, DM_write_data_MIF_15, 
        DM_write_data_MIF_14, DM_write_data_MIF_13, DM_write_data_MIF_12, 
        DM_write_data_MIF_11, DM_write_data_MIF_10, DM_write_data_MIF_9, 
        DM_write_data_MIF_8, DM_write_data_MIF_7, DM_write_data_MIF_6, 
        DM_write_data_MIF_5, DM_write_data_MIF_4, DM_write_data_MIF_3, 
        DM_write_data_MIF_2, DM_write_data_MIF_1, DM_write_data_MIF_0}), 
        .DM_write(DM_write), .mask({mask_to_mem_3, mask_to_mem_2, 
        mask_to_mem_1, mask_to_mem_0}) );
    mem_load mem_load_inst ( .start(memory_load_enable), .scan_in(scan_in), 
        .scan_out(scan_out), .scan_clk(shift_clk), .data_out({data_out_load_31, 
        data_out_load_30, data_out_load_29, data_out_load_28, data_out_load_27, 
        data_out_load_26, data_out_load_25, data_out_load_24, data_out_load_23, 
        data_out_load_22, data_out_load_21, data_out_load_20, data_out_load_19, 
        data_out_load_18, data_out_load_17, data_out_load_16, data_out_load_15, 
        data_out_load_14, data_out_load_13, data_out_load_12, data_out_load_11, 
        data_out_load_10, data_out_load_9, data_out_load_8, data_out_load_7, 
        data_out_load_6, data_out_load_5, data_out_load_4, data_out_load_3, 
        data_out_load_2, data_out_load_1, data_out_load_0}), .data_in({
        data_in_to_sh_reg_31, data_in_to_sh_reg_30, data_in_to_sh_reg_29, 
        data_in_to_sh_reg_28, data_in_to_sh_reg_27, data_in_to_sh_reg_26, 
        data_in_to_sh_reg_25, data_in_to_sh_reg_24, data_in_to_sh_reg_23, 
        data_in_to_sh_reg_22, data_in_to_sh_reg_21, data_in_to_sh_reg_20, 
        data_in_to_sh_reg_19, data_in_to_sh_reg_18, data_in_to_sh_reg_17, 
        data_in_to_sh_reg_16, data_in_to_sh_reg_15, data_in_to_sh_reg_14, 
        data_in_to_sh_reg_13, data_in_to_sh_reg_12, data_in_to_sh_reg_11, 
        data_in_to_sh_reg_10, data_in_to_sh_reg_9, data_in_to_sh_reg_8, 
        data_in_to_sh_reg_7, data_in_to_sh_reg_6, data_in_to_sh_reg_5, 
        data_in_to_sh_reg_4, data_in_to_sh_reg_3, data_in_to_sh_reg_2, 
        data_in_to_sh_reg_1, data_in_to_sh_reg_0}), .data_write(
        data_write_load), .read(read), .addr_out({addr_out_load_10, 
        addr_out_load_9, addr_out_load_8, addr_out_load_7, addr_out_load_6, 
        addr_out_load_5, addr_out_load_4, addr_out_load_3, addr_out_load_2, 
        SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2}) );
    aspida_net_core chain_inst ( .nrst(nrst), .clk(wish_clk), .ip_c_req(
        ip_not_local), .ip_c_we(1'b0), .ip_c_mult(1'b0), .ip_c_prd(1'b0), 
        .ip_c_seq(1'b0), .ip_c_ts({1'b0, 1'b0, 1'b0}), .ip_c_sel({1'b1, 1'b1, 
        1'b1, 1'b1}), .ip_c_adr({IM_addr_31, IM_addr_30, IM_addr_29, 
        IM_addr_28, IM_addr_27, IM_addr_26, IM_addr_25, IM_addr_24, IM_addr_23, 
        IM_addr_22, IM_addr_21, IM_addr_20, IM_addr_19, IM_addr_18, IM_addr_17, 
        IM_addr_16, IM_addr_15, IM_addr_14, IM_addr_13, IM_addr_12, IM_addr_11, 
        IM_addr_10, IM_addr_9, IM_addr_8, IM_addr_7, IM_addr_6, IM_addr_5, 
        IM_addr_4, IM_addr_3, IM_addr_2, IM_addr_1, IM_addr_0}), .ip_c_dat({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ip_c_ack(ip_c_ack), 
        .ip_r_req(ip_r_req), .ip_r_dat({ip_r_dat_31, ip_r_dat_30, ip_r_dat_29, 
        ip_r_dat_28, ip_r_dat_27, ip_r_dat_26, ip_r_dat_25, ip_r_dat_24, 
        ip_r_dat_23, ip_r_dat_22, ip_r_dat_21, ip_r_dat_20, ip_r_dat_19, 
        ip_r_dat_18, ip_r_dat_17, ip_r_dat_16, ip_r_dat_15, ip_r_dat_14, 
        ip_r_dat_13, ip_r_dat_12, ip_r_dat_11, ip_r_dat_10, ip_r_dat_9, 
        ip_r_dat_8, ip_r_dat_7, ip_r_dat_6, ip_r_dat_5, ip_r_dat_4, ip_r_dat_3, 
        ip_r_dat_2, ip_r_dat_1, ip_r_dat_0}), .ip_r_ack(ip_r_ack), .dp_c_req(
        dp_not_local), .dp_c_we(DM_write), .dp_c_mult(1'b0), .dp_c_prd(1'b0), 
        .dp_c_seq(1'b0), .dp_c_ts({1'b0, 1'b0, 1'b0}), .dp_c_sel({
        mask_to_mem_3, mask_to_mem_2, mask_to_mem_1, mask_to_mem_0}), 
        .dp_c_adr({DM_addr_CPU_31, DM_addr_CPU_30, DM_addr_CPU_29, 
        DM_addr_CPU_28, DM_addr_CPU_27, DM_addr_CPU_26, DM_addr_CPU_25, 
        DM_addr_CPU_24, DM_addr_CPU_23, DM_addr_CPU_22, DM_addr_CPU_21, 
        DM_addr_CPU_20, DM_addr_CPU_19, DM_addr_CPU_18, DM_addr_CPU_17, 
        DM_addr_CPU_16, DM_addr_CPU_15, DM_addr_CPU_14, DM_addr_CPU_13, 
        DM_addr_CPU_12, DM_addr_CPU_11, DM_addr_CPU_10, DM_addr_CPU_9, 
        DM_addr_CPU_8, DM_addr_CPU_7, DM_addr_CPU_6, DM_addr_CPU_5, 
        DM_addr_CPU_4, DM_addr_CPU_3, DM_addr_CPU_2, DM_addr_CPU_1, 
        DM_addr_CPU_0}), .dp_c_dat({DM_write_data_MIF_31, DM_write_data_MIF_30, 
        DM_write_data_MIF_29, DM_write_data_MIF_28, DM_write_data_MIF_27, 
        DM_write_data_MIF_26, DM_write_data_MIF_25, DM_write_data_MIF_24, 
        DM_write_data_MIF_23, DM_write_data_MIF_22, DM_write_data_MIF_21, 
        DM_write_data_MIF_20, DM_write_data_MIF_19, DM_write_data_MIF_18, 
        DM_write_data_MIF_17, DM_write_data_MIF_16, DM_write_data_MIF_15, 
        DM_write_data_MIF_14, DM_write_data_MIF_13, DM_write_data_MIF_12, 
        DM_write_data_MIF_11, DM_write_data_MIF_10, DM_write_data_MIF_9, 
        DM_write_data_MIF_8, DM_write_data_MIF_7, DM_write_data_MIF_6, 
        DM_write_data_MIF_5, DM_write_data_MIF_4, DM_write_data_MIF_3, 
        DM_write_data_MIF_2, DM_write_data_MIF_1, DM_write_data_MIF_0}), 
        .dp_c_ack(dp_c_ack), .dp_r_req(dp_r_req), .dp_r_dat({dp_r_dat_31, 
        dp_r_dat_30, dp_r_dat_29, dp_r_dat_28, dp_r_dat_27, dp_r_dat_26, 
        dp_r_dat_25, dp_r_dat_24, dp_r_dat_23, dp_r_dat_22, dp_r_dat_21, 
        dp_r_dat_20, dp_r_dat_19, dp_r_dat_18, dp_r_dat_17, dp_r_dat_16, 
        dp_r_dat_15, dp_r_dat_14, dp_r_dat_13, dp_r_dat_12, dp_r_dat_11, 
        dp_r_dat_10, dp_r_dat_9, dp_r_dat_8, dp_r_dat_7, dp_r_dat_6, 
        dp_r_dat_5, dp_r_dat_4, dp_r_dat_3, dp_r_dat_2, dp_r_dat_1, dp_r_dat_0
        }), .dp_r_ack(dp_r_ack), .ei_c_req(ei_c_req), .ei_c_ack(ei_c_ack), 
        .ei_c_we(ei_c_we), .ei_c_addr({ei_c_addr_10, ei_c_addr_9, ei_c_addr_8, 
        ei_c_addr_7, ei_c_addr_6, ei_c_addr_5, ei_c_addr_4, ei_c_addr_3, 
        ei_c_addr_2, ei_c_addr_1, ei_c_addr_0}), .ei_r_req(ei_r_req), 
        .ei_r_ack(ei_r_ack), .ei_data_in({ei_data_in_7, ei_data_in_6, 
        ei_data_in_5, ei_data_in_4, ei_data_in_3, ei_data_in_2, ei_data_in_1, 
        ei_data_in_0}), .ei_data_out({ei_data_out_7, ei_data_out_6, 
        ei_data_out_5, ei_data_out_4, ei_data_out_3, ei_data_out_2, 
        ei_data_out_1, ei_data_out_0}), .c_BC({c_BC_4, c_BC_3, c_BC_2, c_BC_1, 
        c_BC_0}), .c_BC_ack(c_BC_ack), .r_BC({r_BC_4, r_BC_3, r_BC_2, r_BC_1, 
        r_BC_0}), .r_BC_ack(r_BC_ack), .wish_we_o(wish_we_o), .wish_stb_cyc_o(
        wish_stb_cyc_o), .wish_ack_i(wish_ack_i), .wish_adr_o({wish_adr_o_11, 
        wish_adr_o_10, wish_adr_o_9, wish_adr_o_8, wish_adr_o_7, wish_adr_o_6, 
        wish_adr_o_5, wish_adr_o_4, wish_adr_o_3, wish_adr_o_2, wish_adr_o_1, 
        wish_adr_o_0}), .wish_dat_i({wish_dat_i_31, wish_dat_i_30, 
        wish_dat_i_29, wish_dat_i_28, wish_dat_i_27, wish_dat_i_26, 
        wish_dat_i_25, wish_dat_i_24, wish_dat_i_23, wish_dat_i_22, 
        wish_dat_i_21, wish_dat_i_20, wish_dat_i_19, wish_dat_i_18, 
        wish_dat_i_17, wish_dat_i_16, wish_dat_i_15, wish_dat_i_14, 
        wish_dat_i_13, wish_dat_i_12, wish_dat_i_11, wish_dat_i_10, 
        wish_dat_i_9, wish_dat_i_8, wish_dat_i_7, wish_dat_i_6, wish_dat_i_5, 
        wish_dat_i_4, wish_dat_i_3, wish_dat_i_2, wish_dat_i_1, wish_dat_i_0}), 
        .wish_dat_o({wish_dat_o_31, wish_dat_o_30, wish_dat_o_29, 
        wish_dat_o_28, wish_dat_o_27, wish_dat_o_26, wish_dat_o_25, 
        wish_dat_o_24, wish_dat_o_23, wish_dat_o_22, wish_dat_o_21, 
        wish_dat_o_20, wish_dat_o_19, wish_dat_o_18, wish_dat_o_17, 
        wish_dat_o_16, wish_dat_o_15, wish_dat_o_14, wish_dat_o_13, 
        wish_dat_o_12, wish_dat_o_11, wish_dat_o_10, wish_dat_o_9, 
        wish_dat_o_8, wish_dat_o_7, wish_dat_o_6, wish_dat_o_5, wish_dat_o_4, 
        wish_dat_o_3, wish_dat_o_2, wish_dat_o_1, wish_dat_o_0}), .dm_c_req(
        dm_c_req), .dm_c_we(dm_c_we), .dm_c_mult(dm_c_mult), .dm_c_ts({
        dm_c_ts_2, dm_c_ts_1, dm_c_ts_0}), .dm_c_sel({dm_c_sel_3, dm_c_sel_2, 
        dm_c_sel_1, dm_c_sel_0}), .dm_c_adr({SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, 
        SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, 
        SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21, 
        SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23, dm_c_adr_10, 
        dm_c_adr_9, dm_c_adr_8, dm_c_adr_7, dm_c_adr_6, dm_c_adr_5, dm_c_adr_4, 
        dm_c_adr_3, dm_c_adr_2, SYNOPSYS_UNCONNECTED_24, 
        SYNOPSYS_UNCONNECTED_25}), .dm_c_dat({dm_c_dat_31, dm_c_dat_30, 
        dm_c_dat_29, dm_c_dat_28, dm_c_dat_27, dm_c_dat_26, dm_c_dat_25, 
        dm_c_dat_24, dm_c_dat_23, dm_c_dat_22, dm_c_dat_21, dm_c_dat_20, 
        dm_c_dat_19, dm_c_dat_18, dm_c_dat_17, dm_c_dat_16, dm_c_dat_15, 
        dm_c_dat_14, dm_c_dat_13, dm_c_dat_12, dm_c_dat_11, dm_c_dat_10, 
        dm_c_dat_9, dm_c_dat_8, dm_c_dat_7, dm_c_dat_6, dm_c_dat_5, dm_c_dat_4, 
        dm_c_dat_3, dm_c_dat_2, dm_c_dat_1, dm_c_dat_0}), .dm_c_ack(
        dm_grant_chain_d), .dm_r_req(dm_r_req), .dm_r_err(1'b0), .dm_r_rty(
        1'b0), .dm_r_acc(1'b0), .dm_r_mult(dm_c_mult_latched), .dm_r_ts({
        dm_c_ts_latched_2, dm_c_ts_latched_1, dm_c_ts_latched_0}), .dm_r_rt({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .dm_r_sel({dm_c_sel_latched_3, 
        dm_c_sel_latched_2, dm_c_sel_latched_1, dm_c_sel_latched_0}), 
        .dm_r_dat({DM_read_data_mem_31, DM_read_data_mem_30, 
        DM_read_data_mem_29, DM_read_data_mem_28, DM_read_data_mem_27, 
        DM_read_data_mem_26, DM_read_data_mem_25, DM_read_data_mem_24, 
        DM_read_data_mem_23, DM_read_data_mem_22, DM_read_data_mem_21, 
        DM_read_data_mem_20, DM_read_data_mem_19, DM_read_data_mem_18, 
        DM_read_data_mem_17, DM_read_data_mem_16, DM_read_data_mem_15, 
        DM_read_data_mem_14, DM_read_data_mem_13, DM_read_data_mem_12, 
        DM_read_data_mem_11, DM_read_data_mem_10, DM_read_data_mem_9, 
        DM_read_data_mem_8, DM_read_data_mem_7, DM_read_data_mem_6, 
        DM_read_data_mem_5, DM_read_data_mem_4, DM_read_data_mem_3, 
        DM_read_data_mem_2, DM_read_data_mem_1, DM_read_data_mem_0}), 
        .dm_r_ack(dm_r_ack), .im_c_req(im_c_req), .im_c_we(im_c_we), 
        .im_c_mult(im_c_mult), .im_c_ts({im_c_ts_2, im_c_ts_1, im_c_ts_0}), 
        .im_c_sel({im_c_sel_3, im_c_sel_2, im_c_sel_1, im_c_sel_0}), 
        .im_c_adr({SYNOPSYS_UNCONNECTED_26, SYNOPSYS_UNCONNECTED_27, 
        SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29, 
        SYNOPSYS_UNCONNECTED_30, SYNOPSYS_UNCONNECTED_31, 
        SYNOPSYS_UNCONNECTED_32, SYNOPSYS_UNCONNECTED_33, 
        SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35, 
        SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37, 
        SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39, 
        SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_41, 
        SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_43, 
        SYNOPSYS_UNCONNECTED_44, SYNOPSYS_UNCONNECTED_45, 
        SYNOPSYS_UNCONNECTED_46, im_c_adr_10, im_c_adr_9, im_c_adr_8, 
        im_c_adr_7, im_c_adr_6, im_c_adr_5, im_c_adr_4, im_c_adr_3, im_c_adr_2, 
        SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48}), .im_c_dat({
        im_c_dat_31, im_c_dat_30, im_c_dat_29, im_c_dat_28, im_c_dat_27, 
        im_c_dat_26, im_c_dat_25, im_c_dat_24, im_c_dat_23, im_c_dat_22, 
        im_c_dat_21, im_c_dat_20, im_c_dat_19, im_c_dat_18, im_c_dat_17, 
        im_c_dat_16, im_c_dat_15, im_c_dat_14, im_c_dat_13, im_c_dat_12, 
        im_c_dat_11, im_c_dat_10, im_c_dat_9, im_c_dat_8, im_c_dat_7, 
        im_c_dat_6, im_c_dat_5, im_c_dat_4, im_c_dat_3, im_c_dat_2, im_c_dat_1, 
        im_c_dat_0}), .im_c_ack(im_grant_chain_d), .im_r_req(im_r_req), 
        .im_r_err(1'b0), .im_r_rty(1'b0), .im_r_acc(1'b0), .im_r_mult(
        im_c_mult_latched), .im_r_ts({im_c_ts_latched_2, im_c_ts_latched_1, 
        im_c_ts_latched_0}), .im_r_rt({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .im_r_sel({im_c_sel_latched_3, im_c_sel_latched_2, im_c_sel_latched_1, 
        im_c_sel_latched_0}), .im_r_dat({IM_read_data_mem_31, 
        IM_read_data_mem_30, IM_read_data_mem_29, IM_read_data_mem_28, 
        IM_read_data_mem_27, IM_read_data_mem_26, IM_read_data_mem_25, 
        IM_read_data_mem_24, IM_read_data_mem_23, IM_read_data_mem_22, 
        IM_read_data_mem_21, IM_read_data_mem_20, IM_read_data_mem_19, 
        IM_read_data_mem_18, IM_read_data_mem_17, IM_read_data_mem_16, 
        IM_read_data_mem_15, IM_read_data_mem_14, IM_read_data_mem_13, 
        IM_read_data_mem_12, IM_read_data_mem_11, IM_read_data_mem_10, 
        IM_read_data_mem_9, IM_read_data_mem_8, IM_read_data_mem_7, 
        IM_read_data_mem_6, IM_read_data_mem_5, IM_read_data_mem_4, 
        IM_read_data_mem_3, IM_read_data_mem_2, IM_read_data_mem_1, 
        IM_read_data_mem_0}), .im_r_ack(im_r_ack), .test_si(1'b0), .test_se(
        1'b0), .phi1(1'b1), .phi2(1'b0), .phi3(1'b1), .force_bare(force_bare)
         );
    sram2k_pin instr_ram ( .a0(IM_addr_MEM_mem_2), .a1(IM_addr_MEM_mem_3), 
        .a2(IM_addr_MEM_mem_4), .a3(IM_addr_MEM_mem_5), .a4(IM_addr_MEM_mem_6), 
        .a5(IM_addr_MEM_mem_7), .a6(IM_addr_MEM_mem_8), .a7(IM_addr_MEM_mem_9), 
        .a8(IM_addr_MEM_mem_10), .di0(IM_write_data_mem_0), .di1(
        IM_write_data_mem_1), .di2(IM_write_data_mem_2), .di3(
        IM_write_data_mem_3), .di4(IM_write_data_mem_4), .di5(
        IM_write_data_mem_5), .di6(IM_write_data_mem_6), .di7(
        IM_write_data_mem_7), .di8(IM_write_data_mem_8), .di9(
        IM_write_data_mem_9), .di10(IM_write_data_mem_10), .di11(
        IM_write_data_mem_11), .di12(IM_write_data_mem_12), .di13(
        IM_write_data_mem_13), .di14(IM_write_data_mem_14), .di15(
        IM_write_data_mem_15), .di16(IM_write_data_mem_16), .di17(
        IM_write_data_mem_17), .di18(IM_write_data_mem_18), .di19(
        IM_write_data_mem_19), .di20(IM_write_data_mem_20), .di21(
        IM_write_data_mem_21), .di22(IM_write_data_mem_22), .di23(
        IM_write_data_mem_23), .di24(IM_write_data_mem_24), .di25(
        IM_write_data_mem_25), .di26(IM_write_data_mem_26), .di27(
        IM_write_data_mem_27), .di28(IM_write_data_mem_28), .di29(
        IM_write_data_mem_29), .di30(IM_write_data_mem_30), .di31(
        IM_write_data_mem_31), .clk(IMem_clk), .wrb(data_write_load_im), .ceb(
        1'b0), .iwen3(IM_mask_we_3), .iwen2(IM_mask_we_2), .iwen1(IM_mask_we_1
        ), .iwen0(IM_mask_we_0), .oen3(IM_mask_oe_3), .oen2(IM_mask_oe_2), 
        .oen1(IM_mask_oe_1), .oen0(IM_mask_oe_0), .do0(IM_read_data_mem_0), 
        .do1(IM_read_data_mem_1), .do2(IM_read_data_mem_2), .do3(
        IM_read_data_mem_3), .do4(IM_read_data_mem_4), .do5(IM_read_data_mem_5
        ), .do6(IM_read_data_mem_6), .do7(IM_read_data_mem_7), .do8(
        IM_read_data_mem_8), .do9(IM_read_data_mem_9), .do10(
        IM_read_data_mem_10), .do11(IM_read_data_mem_11), .do12(
        IM_read_data_mem_12), .do13(IM_read_data_mem_13), .do14(
        IM_read_data_mem_14), .do15(IM_read_data_mem_15), .do16(
        IM_read_data_mem_16), .do17(IM_read_data_mem_17), .do18(
        IM_read_data_mem_18), .do19(IM_read_data_mem_19), .do20(
        IM_read_data_mem_20), .do21(IM_read_data_mem_21), .do22(
        IM_read_data_mem_22), .do23(IM_read_data_mem_23), .do24(
        IM_read_data_mem_24), .do25(IM_read_data_mem_25), .do26(
        IM_read_data_mem_26), .do27(IM_read_data_mem_27), .do28(
        IM_read_data_mem_28), .do29(IM_read_data_mem_29), .do30(
        IM_read_data_mem_30), .do31(IM_read_data_mem_31) );
    sram2k_pin data_ram ( .a0(DM_addr_MEM_mem_2), .a1(DM_addr_MEM_mem_3), .a2(
        DM_addr_MEM_mem_4), .a3(DM_addr_MEM_mem_5), .a4(DM_addr_MEM_mem_6), 
        .a5(DM_addr_MEM_mem_7), .a6(DM_addr_MEM_mem_8), .a7(DM_addr_MEM_mem_9), 
        .a8(DM_addr_MEM_mem_10), .di0(DM_write_data_mem_0), .di1(
        DM_write_data_mem_1), .di2(DM_write_data_mem_2), .di3(
        DM_write_data_mem_3), .di4(DM_write_data_mem_4), .di5(
        DM_write_data_mem_5), .di6(DM_write_data_mem_6), .di7(
        DM_write_data_mem_7), .di8(DM_write_data_mem_8), .di9(
        DM_write_data_mem_9), .di10(DM_write_data_mem_10), .di11(
        DM_write_data_mem_11), .di12(DM_write_data_mem_12), .di13(
        DM_write_data_mem_13), .di14(DM_write_data_mem_14), .di15(
        DM_write_data_mem_15), .di16(DM_write_data_mem_16), .di17(
        DM_write_data_mem_17), .di18(DM_write_data_mem_18), .di19(
        DM_write_data_mem_19), .di20(DM_write_data_mem_20), .di21(
        DM_write_data_mem_21), .di22(DM_write_data_mem_22), .di23(
        DM_write_data_mem_23), .di24(DM_write_data_mem_24), .di25(
        DM_write_data_mem_25), .di26(DM_write_data_mem_26), .di27(
        DM_write_data_mem_27), .di28(DM_write_data_mem_28), .di29(
        DM_write_data_mem_29), .di30(DM_write_data_mem_30), .di31(
        DM_write_data_mem_31), .clk(DMem_clk), .wrb(data_write_load_dm), .ceb(
        1'b0), .iwen3(DM_mask_we_3), .iwen2(DM_mask_we_2), .iwen1(DM_mask_we_1
        ), .iwen0(DM_mask_we_0), .oen3(DM_mask_oe_3), .oen2(DM_mask_oe_2), 
        .oen1(DM_mask_oe_1), .oen0(DM_mask_oe_0), .do0(DM_read_data_mem_0), 
        .do1(DM_read_data_mem_1), .do2(DM_read_data_mem_2), .do3(
        DM_read_data_mem_3), .do4(DM_read_data_mem_4), .do5(DM_read_data_mem_5
        ), .do6(DM_read_data_mem_6), .do7(DM_read_data_mem_7), .do8(
        DM_read_data_mem_8), .do9(DM_read_data_mem_9), .do10(
        DM_read_data_mem_10), .do11(DM_read_data_mem_11), .do12(
        DM_read_data_mem_12), .do13(DM_read_data_mem_13), .do14(
        DM_read_data_mem_14), .do15(DM_read_data_mem_15), .do16(
        DM_read_data_mem_16), .do17(DM_read_data_mem_17), .do18(
        DM_read_data_mem_18), .do19(DM_read_data_mem_19), .do20(
        DM_read_data_mem_20), .do21(DM_read_data_mem_21), .do22(
        DM_read_data_mem_22), .do23(DM_read_data_mem_23), .do24(
        DM_read_data_mem_24), .do25(DM_read_data_mem_25), .do26(
        DM_read_data_mem_26), .do27(DM_read_data_mem_27), .do28(
        DM_read_data_mem_28), .do29(DM_read_data_mem_29), .do30(
        DM_read_data_mem_30), .do31(DM_read_data_mem_31) );
    oai21_1 U3 ( .x(Ctrl__IFinst___Regs_1__ri), .a(STOP_fetch), .b(N315), .c(
        n127) );
    nand2i_2 U4 ( .x(Ctrl__MEMinst___Regs_1__ri), .a(dp_complete), .b(n124) );
    oa21_2 U5 ( .x(n124), .a(n138), .b(n125), .c(N597) );
    inv_2 U6 ( .x(n127), .a(ip_complete) );
    mux2_2 U7 ( .x(reset_DLX_ctrl), .d0(reset_DLX_c), .sl(reset_ctrl), .d1(
        n103) );
    inv_2 U8 ( .x(N597), .a(DM_complete_latched) );
    nor2i_1 U9 ( .x(_42_net_), .a(nrst), .b(dm_r_ack) );
    inv_2 U10 ( .x(N315), .a(IM_complete_latched) );
    nor2i_1 U11 ( .x(_38_net_), .a(nrst), .b(im_r_ack) );
    and2_1 U12 ( .x(_37_net_), .a(dm_grant_local_d), .b(DM_complete) );
    and3i_1 U13 ( .x(dp_local), .a(n126), .b(n125), .c(
        Ctrl__EXinst___Regs_1__ro) );
    nand2i_2 U14 ( .x(n125), .a(DM_read), .b(n145) );
    or3i_2 U15 ( .x(n126), .a(DM_addr_CPU_11), .b(DM_addr_CPU_31), .c(
        DM_addr_CPU_12) );
    inv_2 U16 ( .x(n138), .a(Ctrl__EXinst___Regs_1__ro) );
    and2_1 U17 ( .x(_36_net_), .a(im_grant_local_d), .b(IM_complete) );
    and2_1 U18 ( .x(ip_local), .a(n128), .b(Ctrl__IFinst___Regs_1__ro) );
    inv_2 U19 ( .x(n128), .a(n137) );
    or3_2 U20 ( .x(n137), .a(IM_addr_31), .b(IM_addr_11), .c(IM_addr_12) );
    mux2_2 U21 ( .x(IM_read_data_9), .d0(IM_read_data_mem_latched_9), .sl(
        ip_not_local), .d1(ip_r_dat_9) );
    mux2_2 U22 ( .x(IM_read_data_8), .d0(IM_read_data_mem_latched_8), .sl(
        ip_not_local), .d1(ip_r_dat_8) );
    mux2_2 U23 ( .x(IM_read_data_7), .d0(IM_read_data_mem_latched_7), .sl(
        ip_not_local), .d1(ip_r_dat_7) );
    mux2_2 U24 ( .x(IM_read_data_6), .d0(IM_read_data_mem_latched_6), .sl(
        ip_not_local), .d1(ip_r_dat_6) );
    mux2_2 U25 ( .x(IM_read_data_5), .d0(IM_read_data_mem_latched_5), .sl(
        ip_not_local), .d1(ip_r_dat_5) );
    mux2_2 U26 ( .x(IM_read_data_4), .d0(IM_read_data_mem_latched_4), .sl(
        ip_not_local), .d1(ip_r_dat_4) );
    mux2_2 U27 ( .x(IM_read_data_3), .d0(IM_read_data_mem_latched_3), .sl(
        ip_not_local), .d1(ip_r_dat_3) );
    mux2_2 U28 ( .x(IM_read_data_31), .d0(IM_read_data_mem_latched_31), .sl(
        ip_not_local), .d1(ip_r_dat_31) );
    mux2_2 U29 ( .x(IM_read_data_30), .d0(IM_read_data_mem_latched_30), .sl(
        ip_not_local), .d1(ip_r_dat_30) );
    mux2_2 U30 ( .x(IM_read_data_2), .d0(IM_read_data_mem_latched_2), .sl(
        ip_not_local), .d1(ip_r_dat_2) );
    mux2_2 U31 ( .x(IM_read_data_29), .d0(IM_read_data_mem_latched_29), .sl(
        ip_not_local), .d1(ip_r_dat_29) );
    mux2_2 U32 ( .x(IM_read_data_28), .d0(IM_read_data_mem_latched_28), .sl(
        ip_not_local), .d1(ip_r_dat_28) );
    mux2_2 U33 ( .x(IM_read_data_27), .d0(IM_read_data_mem_latched_27), .sl(
        ip_not_local), .d1(ip_r_dat_27) );
    mux2_2 U35 ( .x(IM_read_data_26), .d0(IM_read_data_mem_latched_26), .sl(
        ip_not_local), .d1(ip_r_dat_26) );
    mux2_2 U36 ( .x(IM_read_data_25), .d0(IM_read_data_mem_latched_25), .sl(
        ip_not_local), .d1(ip_r_dat_25) );
    mux2_2 U37 ( .x(IM_read_data_24), .d0(IM_read_data_mem_latched_24), .sl(
        n108), .d1(ip_r_dat_24) );
    mux2_2 U39 ( .x(IM_read_data_23), .d0(IM_read_data_mem_latched_23), .sl(
        ip_not_local), .d1(ip_r_dat_23) );
    mux2_2 U40 ( .x(IM_read_data_22), .d0(IM_read_data_mem_latched_22), .sl(
        ip_not_local), .d1(ip_r_dat_22) );
    mux2_2 U41 ( .x(IM_read_data_21), .d0(IM_read_data_mem_latched_21), .sl(
        ip_not_local), .d1(ip_r_dat_21) );
    mux2_2 U42 ( .x(IM_read_data_20), .d0(IM_read_data_mem_latched_20), .sl(
        ip_not_local), .d1(ip_r_dat_20) );
    mux2_2 U43 ( .x(IM_read_data_1), .d0(IM_read_data_mem_latched_1), .sl(
        ip_not_local), .d1(ip_r_dat_1) );
    mux2_2 U44 ( .x(IM_read_data_19), .d0(IM_read_data_mem_latched_19), .sl(
        ip_not_local), .d1(ip_r_dat_19) );
    mux2_2 U45 ( .x(IM_read_data_18), .d0(IM_read_data_mem_latched_18), .sl(
        ip_not_local), .d1(ip_r_dat_18) );
    mux2_2 U46 ( .x(IM_read_data_17), .d0(IM_read_data_mem_latched_17), .sl(
        ip_not_local), .d1(ip_r_dat_17) );
    mux2_2 U47 ( .x(IM_read_data_16), .d0(IM_read_data_mem_latched_16), .sl(
        ip_not_local), .d1(ip_r_dat_16) );
    mux2_2 U48 ( .x(IM_read_data_15), .d0(IM_read_data_mem_latched_15), .sl(
        ip_not_local), .d1(ip_r_dat_15) );
    mux2_2 U49 ( .x(IM_read_data_14), .d0(IM_read_data_mem_latched_14), .sl(
        ip_not_local), .d1(ip_r_dat_14) );
    mux2_2 U50 ( .x(IM_read_data_13), .d0(IM_read_data_mem_latched_13), .sl(
        ip_not_local), .d1(ip_r_dat_13) );
    mux2_2 U51 ( .x(IM_read_data_12), .d0(IM_read_data_mem_latched_12), .sl(
        ip_not_local), .d1(ip_r_dat_12) );
    mux2_2 U52 ( .x(IM_read_data_11), .d0(IM_read_data_mem_latched_11), .sl(
        ip_not_local), .d1(ip_r_dat_11) );
    mux2_2 U53 ( .x(IM_read_data_10), .d0(IM_read_data_mem_latched_10), .sl(
        ip_not_local), .d1(ip_r_dat_10) );
    mux2_2 U54 ( .x(IM_read_data_0), .d0(IM_read_data_mem_latched_0), .sl(
        ip_not_local), .d1(ip_r_dat_0) );
    and2_1 U55 ( .x(_44_net_), .a(nrst), .b(N1431) );
    inv_2 U56 ( .x(N1431), .a(DM_complete) );
    and2_1 U57 ( .x(_39_net_), .a(N1429), .b(nrst) );
    inv_2 U58 ( .x(N1429), .a(IM_complete) );
    nand2_2 U59 ( .x(n155), .a(data_write_load), .b(n140) );
    inv_2 U60 ( .x(n140), .a(n160) );
    nand2_2 U61 ( .x(n156), .a(DM_write), .b(n144) );
    mux2_2 U62 ( .x(n150), .d0(n154), .sl(dm_grant_chain), .d1(n153) );
    nand2_2 U63 ( .x(n154), .a(DM_write), .b(n160) );
    nand2_2 U64 ( .x(n153), .a(dm_c_we), .b(n160) );
    inv_2 U65 ( .x(n145), .a(DM_write) );
    inv_2 U66 ( .x(n38), .a(dm_grant_chain_d) );
    inv_2 U67 ( .x(n39), .a(im_grant_chain_d) );
    nor2i_1 U68 ( .x(n149), .a(n136), .b(global_g2) );
    inv_2 U69 ( .x(_17_net_), .a(ei_c_we) );
    mux2_2 U70 ( .x(data_in_to_sh_reg_0), .d0(n98), .sl(inst_ram_load), .d1(
        IM_read_data_mem_0) );
    mux2_2 U71 ( .x(data_in_to_sh_reg_1), .d0(n97), .sl(inst_ram_load), .d1(
        IM_read_data_mem_1) );
    mux2_2 U72 ( .x(data_in_to_sh_reg_2), .d0(n86), .sl(n160), .d1(
        IM_read_data_mem_2) );
    mux2_2 U73 ( .x(data_in_to_sh_reg_3), .d0(n49), .sl(n160), .d1(
        IM_read_data_mem_3) );
    mux2_2 U74 ( .x(data_in_to_sh_reg_4), .d0(n46), .sl(inst_ram_load), .d1(
        IM_read_data_mem_4) );
    mux2_2 U75 ( .x(data_in_to_sh_reg_5), .d0(n45), .sl(inst_ram_load), .d1(
        IM_read_data_mem_5) );
    mux2_2 U76 ( .x(data_in_to_sh_reg_6), .d0(n44), .sl(n160), .d1(
        IM_read_data_mem_6) );
    mux2_2 U77 ( .x(data_in_to_sh_reg_7), .d0(n43), .sl(inst_ram_load), .d1(
        IM_read_data_mem_7) );
    mux2_2 U78 ( .x(data_in_to_sh_reg_8), .d0(n42), .sl(inst_ram_load), .d1(
        IM_read_data_mem_8) );
    mux2_2 U79 ( .x(data_in_to_sh_reg_9), .d0(n41), .sl(inst_ram_load), .d1(
        IM_read_data_mem_9) );
    mux2_2 U80 ( .x(data_in_to_sh_reg_10), .d0(n96), .sl(inst_ram_load), .d1(
        IM_read_data_mem_10) );
    mux2_2 U81 ( .x(data_in_to_sh_reg_11), .d0(n95), .sl(n160), .d1(
        IM_read_data_mem_11) );
    mux2_2 U82 ( .x(data_in_to_sh_reg_12), .d0(n94), .sl(inst_ram_load), .d1(
        IM_read_data_mem_12) );
    mux2_2 U83 ( .x(data_in_to_sh_reg_13), .d0(n93), .sl(n160), .d1(
        IM_read_data_mem_13) );
    mux2_2 U84 ( .x(data_in_to_sh_reg_14), .d0(n92), .sl(inst_ram_load), .d1(
        IM_read_data_mem_14) );
    mux2_2 U85 ( .x(data_in_to_sh_reg_15), .d0(n91), .sl(n160), .d1(
        IM_read_data_mem_15) );
    mux2_2 U86 ( .x(data_in_to_sh_reg_16), .d0(n90), .sl(inst_ram_load), .d1(
        IM_read_data_mem_16) );
    mux2_2 U87 ( .x(data_in_to_sh_reg_17), .d0(n89), .sl(n160), .d1(
        IM_read_data_mem_17) );
    mux2_2 U88 ( .x(data_in_to_sh_reg_18), .d0(n88), .sl(n160), .d1(
        IM_read_data_mem_18) );
    mux2_2 U89 ( .x(data_in_to_sh_reg_19), .d0(n87), .sl(n160), .d1(
        IM_read_data_mem_19) );
    mux2_2 U90 ( .x(data_in_to_sh_reg_20), .d0(n85), .sl(n160), .d1(
        IM_read_data_mem_20) );
    mux2_2 U91 ( .x(data_in_to_sh_reg_21), .d0(n84), .sl(n160), .d1(
        IM_read_data_mem_21) );
    mux2_2 U92 ( .x(data_in_to_sh_reg_22), .d0(n83), .sl(n160), .d1(
        IM_read_data_mem_22) );
    mux2_2 U93 ( .x(data_in_to_sh_reg_23), .d0(n82), .sl(n160), .d1(
        IM_read_data_mem_23) );
    mux2_2 U94 ( .x(data_in_to_sh_reg_24), .d0(n81), .sl(inst_ram_load), .d1(
        IM_read_data_mem_24) );
    mux2_2 U95 ( .x(data_in_to_sh_reg_25), .d0(n54), .sl(n160), .d1(
        IM_read_data_mem_25) );
    mux2_2 U96 ( .x(data_in_to_sh_reg_26), .d0(n53), .sl(n160), .d1(
        IM_read_data_mem_26) );
    mux2_2 U97 ( .x(data_in_to_sh_reg_27), .d0(n52), .sl(n160), .d1(
        IM_read_data_mem_27) );
    mux2_2 U98 ( .x(data_in_to_sh_reg_28), .d0(n51), .sl(n160), .d1(
        IM_read_data_mem_28) );
    mux2_2 U99 ( .x(data_in_to_sh_reg_29), .d0(n50), .sl(n160), .d1(
        IM_read_data_mem_29) );
    mux2_2 U100 ( .x(data_in_to_sh_reg_30), .d0(n48), .sl(inst_ram_load), .d1(
        IM_read_data_mem_30) );
    mux2_2 U101 ( .x(data_in_to_sh_reg_31), .d0(n47), .sl(n160), .d1(
        IM_read_data_mem_31) );
    inv_2 U102 ( .x(nrst), .a(reset_DLX_c) );
    mux2_2 U103 ( .x(DM_mask_oe_0), .d0(mask_to_mem_0), .sl(dm_grant_chain), 
        .d1(dm_c_sel_latched_0) );
    mux2_2 U104 ( .x(DM_mask_oe_1), .d0(mask_to_mem_1), .sl(dm_grant_chain), 
        .d1(dm_c_sel_latched_1) );
    mux2_2 U105 ( .x(DM_mask_oe_2), .d0(mask_to_mem_2), .sl(dm_grant_chain), 
        .d1(dm_c_sel_latched_2) );
    mux2_2 U106 ( .x(DM_mask_oe_3), .d0(mask_to_mem_3), .sl(dm_grant_chain), 
        .d1(dm_c_sel_latched_3) );
    mux2_2 U107 ( .x(DM_mask_we_0), .d0(mask_to_mem_0), .sl(dm_grant_chain), 
        .d1(dm_c_sel_0) );
    mux2_2 U108 ( .x(DM_mask_we_1), .d0(mask_to_mem_1), .sl(dm_grant_chain), 
        .d1(dm_c_sel_1) );
    mux2_2 U109 ( .x(DM_mask_we_2), .d0(mask_to_mem_2), .sl(dm_grant_chain), 
        .d1(dm_c_sel_2) );
    mux2_2 U110 ( .x(DM_mask_we_3), .d0(mask_to_mem_3), .sl(dm_grant_chain), 
        .d1(dm_c_sel_3) );
    nand2_2 U111 ( .x(data_write_load_dm), .a(n131), .b(n132) );
    oa31_2 U112 ( .x(n131), .a(n111), .b(n143), .c(n144), .d(n150) );
    inv_2 U113 ( .x(n143), .a(dm_c_we) );
    mux2_2 U114 ( .x(n132), .d0(n156), .sl(n157), .d1(n155) );
    ao222_1 U115 ( .x(DM_write_data_mem_31), .a(data_out_load_31), .b(n158), 
        .c(DM_write_data_MIF_31), .d(n129), .e(dm_c_dat_31), .f(n130) );
    ao222_1 U116 ( .x(DM_write_data_mem_30), .a(data_out_load_30), .b(n158), 
        .c(DM_write_data_MIF_30), .d(n159), .e(dm_c_dat_30), .f(n130) );
    ao222_1 U117 ( .x(DM_write_data_mem_29), .a(data_out_load_29), .b(n158), 
        .c(DM_write_data_MIF_29), .d(n129), .e(dm_c_dat_29), .f(n130) );
    ao222_1 U118 ( .x(DM_write_data_mem_28), .a(data_out_load_28), .b(n157), 
        .c(DM_write_data_MIF_28), .d(n159), .e(dm_c_dat_28), .f(n130) );
    ao222_1 U119 ( .x(DM_write_data_mem_27), .a(data_out_load_27), .b(n157), 
        .c(DM_write_data_MIF_27), .d(n129), .e(dm_c_dat_27), .f(n130) );
    ao222_1 U120 ( .x(DM_write_data_mem_26), .a(data_out_load_26), .b(n158), 
        .c(DM_write_data_MIF_26), .d(n159), .e(dm_c_dat_26), .f(n130) );
    ao222_1 U121 ( .x(DM_write_data_mem_25), .a(data_out_load_25), .b(n111), 
        .c(DM_write_data_MIF_25), .d(n129), .e(dm_c_dat_25), .f(n130) );
    ao222_1 U122 ( .x(DM_write_data_mem_24), .a(data_out_load_24), .b(n158), 
        .c(DM_write_data_MIF_24), .d(n159), .e(dm_c_dat_24), .f(n110) );
    ao222_1 U123 ( .x(DM_write_data_mem_23), .a(data_out_load_23), .b(n157), 
        .c(DM_write_data_MIF_23), .d(n129), .e(dm_c_dat_23), .f(n130) );
    ao222_1 U124 ( .x(DM_write_data_mem_22), .a(data_out_load_22), .b(n111), 
        .c(DM_write_data_MIF_22), .d(n159), .e(dm_c_dat_22), .f(n130) );
    ao222_1 U125 ( .x(DM_write_data_mem_21), .a(data_out_load_21), .b(n158), 
        .c(DM_write_data_MIF_21), .d(n129), .e(dm_c_dat_21), .f(n130) );
    ao222_1 U126 ( .x(DM_write_data_mem_20), .a(data_out_load_20), .b(n157), 
        .c(DM_write_data_MIF_20), .d(n159), .e(dm_c_dat_20), .f(n110) );
    ao222_1 U127 ( .x(DM_write_data_mem_19), .a(data_out_load_19), .b(n111), 
        .c(DM_write_data_MIF_19), .d(n129), .e(dm_c_dat_19), .f(n130) );
    ao222_1 U128 ( .x(DM_write_data_mem_18), .a(data_out_load_18), .b(n158), 
        .c(DM_write_data_MIF_18), .d(n159), .e(dm_c_dat_18), .f(n130) );
    ao222_1 U129 ( .x(DM_write_data_mem_17), .a(data_out_load_17), .b(n157), 
        .c(DM_write_data_MIF_17), .d(n129), .e(dm_c_dat_17), .f(n130) );
    ao222_1 U130 ( .x(DM_write_data_mem_16), .a(data_out_load_16), .b(n158), 
        .c(DM_write_data_MIF_16), .d(n159), .e(dm_c_dat_16), .f(n110) );
    ao222_1 U131 ( .x(DM_write_data_mem_15), .a(data_out_load_15), .b(n157), 
        .c(DM_write_data_MIF_15), .d(n129), .e(dm_c_dat_15), .f(n130) );
    ao222_1 U132 ( .x(DM_write_data_mem_14), .a(data_out_load_14), .b(n157), 
        .c(DM_write_data_MIF_14), .d(n159), .e(dm_c_dat_14), .f(n130) );
    ao222_1 U133 ( .x(DM_write_data_mem_13), .a(data_out_load_13), .b(n157), 
        .c(DM_write_data_MIF_13), .d(n129), .e(dm_c_dat_13), .f(n130) );
    ao222_1 U134 ( .x(DM_write_data_mem_12), .a(data_out_load_12), .b(n111), 
        .c(DM_write_data_MIF_12), .d(n159), .e(dm_c_dat_12), .f(n110) );
    ao222_1 U135 ( .x(DM_write_data_mem_11), .a(data_out_load_11), .b(n111), 
        .c(DM_write_data_MIF_11), .d(n129), .e(dm_c_dat_11), .f(n130) );
    ao222_1 U136 ( .x(DM_write_data_mem_10), .a(data_out_load_10), .b(n111), 
        .c(DM_write_data_MIF_10), .d(n159), .e(dm_c_dat_10), .f(n130) );
    ao222_1 U137 ( .x(DM_write_data_mem_9), .a(data_out_load_9), .b(n111), .c(
        DM_write_data_MIF_9), .d(n129), .e(dm_c_dat_9), .f(n130) );
    ao222_1 U138 ( .x(DM_write_data_mem_8), .a(data_out_load_8), .b(n158), .c(
        DM_write_data_MIF_8), .d(n159), .e(dm_c_dat_8), .f(n130) );
    ao222_1 U139 ( .x(DM_write_data_mem_7), .a(data_out_load_7), .b(n158), .c(
        DM_write_data_MIF_7), .d(n129), .e(dm_c_dat_7), .f(n130) );
    ao222_1 U140 ( .x(DM_write_data_mem_6), .a(data_out_load_6), .b(n158), .c(
        DM_write_data_MIF_6), .d(n159), .e(dm_c_dat_6), .f(n130) );
    ao222_1 U141 ( .x(DM_write_data_mem_5), .a(data_out_load_5), .b(n111), .c(
        DM_write_data_MIF_5), .d(n129), .e(dm_c_dat_5), .f(n130) );
    ao222_1 U142 ( .x(DM_write_data_mem_4), .a(data_out_load_4), .b(n158), .c(
        DM_write_data_MIF_4), .d(n159), .e(dm_c_dat_4), .f(n130) );
    ao222_1 U143 ( .x(DM_write_data_mem_3), .a(data_out_load_3), .b(n157), .c(
        DM_write_data_MIF_3), .d(n129), .e(dm_c_dat_3), .f(n130) );
    ao222_1 U144 ( .x(DM_write_data_mem_2), .a(data_out_load_2), .b(n157), .c(
        DM_write_data_MIF_2), .d(n159), .e(dm_c_dat_2), .f(n130) );
    ao222_1 U145 ( .x(DM_write_data_mem_1), .a(data_out_load_1), .b(n111), .c(
        DM_write_data_MIF_1), .d(n129), .e(dm_c_dat_1), .f(n130) );
    ao222_1 U146 ( .x(DM_write_data_mem_0), .a(data_out_load_0), .b(n157), .c(
        DM_write_data_MIF_0), .d(n159), .e(dm_c_dat_0), .f(n130) );
    ao222_1 U147 ( .x(DM_addr_MEM_mem_10), .a(addr_out_load_10), .b(n111), .c(
        DM_addr_MEM_10), .d(n129), .e(dm_c_adr_10), .f(n130) );
    ao222_1 U148 ( .x(DM_addr_MEM_mem_9), .a(addr_out_load_9), .b(n111), .c(
        DM_addr_MEM_9), .d(n159), .e(dm_c_adr_9), .f(n130) );
    ao222_1 U149 ( .x(DM_addr_MEM_mem_8), .a(addr_out_load_8), .b(n158), .c(
        DM_addr_MEM_8), .d(n129), .e(dm_c_adr_8), .f(n130) );
    ao222_1 U150 ( .x(DM_addr_MEM_mem_7), .a(addr_out_load_7), .b(n157), .c(
        DM_addr_MEM_7), .d(n159), .e(dm_c_adr_7), .f(n130) );
    ao222_1 U151 ( .x(DM_addr_MEM_mem_6), .a(addr_out_load_6), .b(n157), .c(
        DM_addr_MEM_6), .d(n129), .e(dm_c_adr_6), .f(n110) );
    ao222_1 U152 ( .x(DM_addr_MEM_mem_5), .a(addr_out_load_5), .b(n158), .c(
        DM_addr_MEM_5), .d(n159), .e(dm_c_adr_5), .f(n110) );
    ao222_1 U153 ( .x(DM_addr_MEM_mem_4), .a(addr_out_load_4), .b(n158), .c(
        DM_addr_MEM_4), .d(n129), .e(dm_c_adr_4), .f(n110) );
    ao222_1 U154 ( .x(DM_addr_MEM_mem_3), .a(addr_out_load_3), .b(n111), .c(
        DM_addr_MEM_3), .d(n159), .e(dm_c_adr_3), .f(n110) );
    ao222_1 U155 ( .x(DM_addr_MEM_mem_2), .a(addr_out_load_2), .b(n111), .c(
        DM_addr_MEM_2), .d(n129), .e(dm_c_adr_2), .f(n110) );
    inv_2 U156 ( .x(n129), .a(n146) );
    nand2_2 U157 ( .x(n146), .a(n139), .b(n144) );
    inv_2 U158 ( .x(n144), .a(dm_grant_chain) );
    inv_2 U159 ( .x(n159), .a(n146) );
    nand2i_2 U160 ( .x(IM_mask_oe_0), .a(im_c_sel_latched_0), .b(
        im_grant_chain) );
    nand2i_2 U161 ( .x(IM_mask_oe_1), .a(im_c_sel_latched_1), .b(
        im_grant_chain) );
    nand2i_2 U162 ( .x(IM_mask_oe_2), .a(im_c_sel_latched_2), .b(
        im_grant_chain) );
    nand2i_2 U163 ( .x(IM_mask_oe_3), .a(im_c_sel_latched_3), .b(
        im_grant_chain) );
    nand2i_2 U164 ( .x(IM_mask_we_0), .a(im_c_sel_0), .b(im_grant_chain) );
    nand2i_2 U165 ( .x(IM_mask_we_1), .a(im_c_sel_1), .b(im_grant_chain) );
    nand2i_2 U166 ( .x(IM_mask_we_2), .a(im_c_sel_2), .b(im_grant_chain) );
    nand2i_2 U167 ( .x(IM_mask_we_3), .a(im_c_sel_3), .b(im_grant_chain) );
    mux2i_1 U168 ( .x(data_write_load_im), .d0(n148), .sl(n135), .d1(n141) );
    nand2_2 U169 ( .x(n148), .a(im_grant_chain), .b(im_c_we) );
    and2_1 U170 ( .x(n135), .a(n160), .b(n158) );
    mux2i_1 U171 ( .x(n133), .d0(n149), .sl(n111), .d1(shift_clk) );
    mux2_2 U172 ( .x(IM_write_data_mem_31), .d0(im_c_dat_31), .sl(n157), .d1(
        data_out_load_31) );
    mux2_2 U173 ( .x(IM_write_data_mem_30), .d0(im_c_dat_30), .sl(n111), .d1(
        data_out_load_30) );
    mux2_2 U174 ( .x(IM_write_data_mem_29), .d0(im_c_dat_29), .sl(n157), .d1(
        data_out_load_29) );
    mux2_2 U175 ( .x(IM_write_data_mem_28), .d0(im_c_dat_28), .sl(n158), .d1(
        data_out_load_28) );
    mux2_2 U176 ( .x(IM_write_data_mem_27), .d0(im_c_dat_27), .sl(n111), .d1(
        data_out_load_27) );
    mux2_2 U177 ( .x(IM_write_data_mem_26), .d0(im_c_dat_26), .sl(n111), .d1(
        data_out_load_26) );
    mux2_2 U178 ( .x(IM_write_data_mem_25), .d0(im_c_dat_25), .sl(n157), .d1(
        data_out_load_25) );
    mux2_2 U179 ( .x(IM_write_data_mem_24), .d0(im_c_dat_24), .sl(n111), .d1(
        data_out_load_24) );
    mux2_2 U180 ( .x(IM_write_data_mem_23), .d0(im_c_dat_23), .sl(n158), .d1(
        data_out_load_23) );
    mux2_2 U181 ( .x(IM_write_data_mem_22), .d0(im_c_dat_22), .sl(n157), .d1(
        data_out_load_22) );
    mux2_2 U182 ( .x(IM_write_data_mem_21), .d0(im_c_dat_21), .sl(n158), .d1(
        data_out_load_21) );
    mux2_2 U183 ( .x(IM_write_data_mem_20), .d0(im_c_dat_20), .sl(n111), .d1(
        data_out_load_20) );
    mux2_2 U184 ( .x(IM_write_data_mem_19), .d0(im_c_dat_19), .sl(n158), .d1(
        data_out_load_19) );
    mux2_2 U185 ( .x(IM_write_data_mem_18), .d0(im_c_dat_18), .sl(n157), .d1(
        data_out_load_18) );
    mux2_2 U186 ( .x(IM_write_data_mem_17), .d0(im_c_dat_17), .sl(n111), .d1(
        data_out_load_17) );
    mux2_2 U187 ( .x(IM_write_data_mem_16), .d0(im_c_dat_16), .sl(n157), .d1(
        data_out_load_16) );
    mux2_2 U188 ( .x(IM_write_data_mem_15), .d0(im_c_dat_15), .sl(n157), .d1(
        data_out_load_15) );
    mux2_2 U189 ( .x(IM_write_data_mem_14), .d0(im_c_dat_14), .sl(n111), .d1(
        data_out_load_14) );
    mux2_2 U190 ( .x(IM_write_data_mem_13), .d0(im_c_dat_13), .sl(n158), .d1(
        data_out_load_13) );
    mux2_2 U191 ( .x(IM_write_data_mem_12), .d0(im_c_dat_12), .sl(n157), .d1(
        data_out_load_12) );
    mux2_2 U192 ( .x(IM_write_data_mem_11), .d0(im_c_dat_11), .sl(n158), .d1(
        data_out_load_11) );
    mux2_2 U193 ( .x(IM_write_data_mem_10), .d0(im_c_dat_10), .sl(n158), .d1(
        data_out_load_10) );
    mux2_2 U194 ( .x(IM_write_data_mem_9), .d0(im_c_dat_9), .sl(n158), .d1(
        data_out_load_9) );
    mux2_2 U195 ( .x(IM_write_data_mem_8), .d0(im_c_dat_8), .sl(n111), .d1(
        data_out_load_8) );
    mux2_2 U196 ( .x(IM_write_data_mem_7), .d0(im_c_dat_7), .sl(n157), .d1(
        data_out_load_7) );
    mux2_2 U197 ( .x(IM_write_data_mem_6), .d0(im_c_dat_6), .sl(n157), .d1(
        data_out_load_6) );
    mux2_2 U198 ( .x(IM_write_data_mem_5), .d0(im_c_dat_5), .sl(n158), .d1(
        data_out_load_5) );
    mux2_2 U199 ( .x(IM_write_data_mem_4), .d0(im_c_dat_4), .sl(n111), .d1(
        data_out_load_4) );
    mux2_2 U200 ( .x(IM_write_data_mem_3), .d0(im_c_dat_3), .sl(n158), .d1(
        data_out_load_3) );
    mux2_2 U201 ( .x(IM_write_data_mem_2), .d0(im_c_dat_2), .sl(n111), .d1(
        data_out_load_2) );
    mux2_2 U202 ( .x(IM_write_data_mem_1), .d0(im_c_dat_1), .sl(n158), .d1(
        data_out_load_1) );
    mux2_2 U203 ( .x(IM_write_data_mem_0), .d0(im_c_dat_0), .sl(n157), .d1(
        data_out_load_0) );
    ao222_1 U204 ( .x(IM_addr_MEM_mem_10), .a(addr_out_load_10), .b(n157), .c(
        IM_addr_10), .d(n40), .e(im_c_adr_10), .f(n37) );
    ao222_1 U205 ( .x(IM_addr_MEM_mem_9), .a(addr_out_load_9), .b(n157), .c(
        IM_addr_9), .d(n40), .e(im_c_adr_9), .f(n37) );
    ao222_1 U206 ( .x(IM_addr_MEM_mem_8), .a(addr_out_load_8), .b(n111), .c(
        IM_addr_8), .d(n40), .e(im_c_adr_8), .f(n37) );
    ao222_1 U207 ( .x(IM_addr_MEM_mem_7), .a(addr_out_load_7), .b(n111), .c(
        IM_addr_7), .d(n40), .e(im_c_adr_7), .f(n37) );
    ao222_1 U208 ( .x(IM_addr_MEM_mem_6), .a(addr_out_load_6), .b(n158), .c(
        IM_addr_6), .d(n40), .e(im_c_adr_6), .f(n37) );
    ao222_1 U209 ( .x(IM_addr_MEM_mem_5), .a(addr_out_load_5), .b(n111), .c(
        IM_addr_5), .d(n40), .e(im_c_adr_5), .f(n37) );
    ao222_1 U210 ( .x(IM_addr_MEM_mem_4), .a(addr_out_load_4), .b(n157), .c(
        IM_addr_4), .d(n40), .e(im_c_adr_4), .f(n37) );
    ao222_1 U211 ( .x(IM_addr_MEM_mem_3), .a(addr_out_load_3), .b(n157), .c(
        IM_addr_3), .d(n40), .e(im_c_adr_3), .f(n37) );
    ao222_1 U212 ( .x(IM_addr_MEM_mem_2), .a(addr_out_load_2), .b(n111), .c(
        IM_addr_2), .d(n40), .e(im_c_adr_2), .f(n37) );
    inv_2 U213 ( .x(n142), .a(im_grant_chain) );
    inv_2 U214 ( .x(n141), .a(data_write_load) );
    dffpr_2 dm_c_sel_latched_reg_0 ( .q(dm_c_sel_latched_0), .rb(nrst), .d(
        dm_c_sel_0), .ck(dm_c_req) );
    dffpr_2 dm_c_sel_latched_reg_1 ( .q(dm_c_sel_latched_1), .rb(nrst), .d(
        dm_c_sel_1), .ck(dm_c_req) );
    dffpr_2 dm_c_sel_latched_reg_2 ( .q(dm_c_sel_latched_2), .rb(nrst), .d(
        dm_c_sel_2), .ck(dm_c_req) );
    dffpr_2 dm_c_sel_latched_reg_3 ( .q(dm_c_sel_latched_3), .rb(nrst), .d(
        dm_c_sel_3), .ck(dm_c_req) );
    dffpr_2 dm_c_ts_latched_reg_0 ( .q(dm_c_ts_latched_0), .rb(nrst), .d(
        dm_c_ts_0), .ck(dm_c_req) );
    dffpr_2 dm_c_ts_latched_reg_1 ( .q(dm_c_ts_latched_1), .rb(nrst), .d(
        dm_c_ts_1), .ck(dm_c_req) );
    dffpr_2 dm_c_ts_latched_reg_2 ( .q(dm_c_ts_latched_2), .rb(nrst), .d(
        dm_c_ts_2), .ck(dm_c_req) );
    dffpr_2 dm_c_mult_latched_reg ( .q(dm_c_mult_latched), .rb(nrst), .d(
        dm_c_mult), .ck(dm_c_req) );
    dffpr_2 im_c_sel_latched_reg_0 ( .q(im_c_sel_latched_0), .rb(nrst), .d(
        im_c_sel_0), .ck(im_c_req) );
    dffpr_2 im_c_sel_latched_reg_1 ( .q(im_c_sel_latched_1), .rb(nrst), .d(
        im_c_sel_1), .ck(im_c_req) );
    dffpr_2 im_c_sel_latched_reg_2 ( .q(im_c_sel_latched_2), .rb(nrst), .d(
        im_c_sel_2), .ck(im_c_req) );
    dffpr_2 im_c_sel_latched_reg_3 ( .q(im_c_sel_latched_3), .rb(nrst), .d(
        im_c_sel_3), .ck(im_c_req) );
    dffpr_2 im_c_ts_latched_reg_0 ( .q(im_c_ts_latched_0), .rb(nrst), .d(
        im_c_ts_0), .ck(im_c_req) );
    dffpr_2 im_c_ts_latched_reg_1 ( .q(im_c_ts_latched_1), .rb(nrst), .d(
        im_c_ts_1), .ck(im_c_req) );
    dffpr_2 im_c_ts_latched_reg_2 ( .q(im_c_ts_latched_2), .rb(nrst), .d(
        im_c_ts_2), .ck(im_c_req) );
    dffpr_2 im_c_mult_latched_reg ( .q(im_c_mult_latched), .rb(nrst), .d(
        im_c_mult), .ck(im_c_req) );
    latn_2 DM_read_data_mem_latched_reg_0 ( .q(DM_read_data_mem_latched_0), 
        .d(DM_read_data_mem_0), .g(n100) );
    latn_2 DM_read_data_mem_latched_reg_1 ( .q(DM_read_data_mem_latched_1), 
        .d(DM_read_data_mem_1), .g(n100) );
    latn_2 DM_read_data_mem_latched_reg_2 ( .q(DM_read_data_mem_latched_2), 
        .d(DM_read_data_mem_2), .g(n100) );
    latn_2 DM_read_data_mem_latched_reg_3 ( .q(DM_read_data_mem_latched_3), 
        .d(DM_read_data_mem_3), .g(n100) );
    latn_2 DM_read_data_mem_latched_reg_4 ( .q(DM_read_data_mem_latched_4), 
        .d(DM_read_data_mem_4), .g(n100) );
    latn_2 DM_read_data_mem_latched_reg_5 ( .q(DM_read_data_mem_latched_5), 
        .d(DM_read_data_mem_5), .g(n100) );
    latn_2 DM_read_data_mem_latched_reg_6 ( .q(DM_read_data_mem_latched_6), 
        .d(DM_read_data_mem_6), .g(n100) );
    latn_2 DM_read_data_mem_latched_reg_7 ( .q(DM_read_data_mem_latched_7), 
        .d(DM_read_data_mem_7), .g(n100) );
    latn_2 DM_read_data_mem_latched_reg_8 ( .q(DM_read_data_mem_latched_8), 
        .d(DM_read_data_mem_8), .g(n100) );
    latn_2 DM_read_data_mem_latched_reg_9 ( .q(DM_read_data_mem_latched_9), 
        .d(DM_read_data_mem_9), .g(n100) );
    latn_2 DM_read_data_mem_latched_reg_10 ( .q(DM_read_data_mem_latched_10), 
        .d(DM_read_data_mem_10), .g(n100) );
    latn_2 DM_read_data_mem_latched_reg_11 ( .q(DM_read_data_mem_latched_11), 
        .d(DM_read_data_mem_11), .g(n100) );
    latn_2 DM_read_data_mem_latched_reg_12 ( .q(DM_read_data_mem_latched_12), 
        .d(DM_read_data_mem_12), .g(n100) );
    latn_2 DM_read_data_mem_latched_reg_13 ( .q(DM_read_data_mem_latched_13), 
        .d(DM_read_data_mem_13), .g(n100) );
    latn_2 DM_read_data_mem_latched_reg_14 ( .q(DM_read_data_mem_latched_14), 
        .d(DM_read_data_mem_14), .g(n100) );
    latn_2 DM_read_data_mem_latched_reg_15 ( .q(DM_read_data_mem_latched_15), 
        .d(DM_read_data_mem_15), .g(n100) );
    latn_2 DM_read_data_mem_latched_reg_16 ( .q(DM_read_data_mem_latched_16), 
        .d(DM_read_data_mem_16), .g(n100) );
    latn_2 DM_read_data_mem_latched_reg_17 ( .q(DM_read_data_mem_latched_17), 
        .d(DM_read_data_mem_17), .g(n100) );
    latn_2 DM_read_data_mem_latched_reg_18 ( .q(DM_read_data_mem_latched_18), 
        .d(DM_read_data_mem_18), .g(n100) );
    latn_2 DM_read_data_mem_latched_reg_19 ( .q(DM_read_data_mem_latched_19), 
        .d(DM_read_data_mem_19), .g(n100) );
    latn_2 DM_read_data_mem_latched_reg_20 ( .q(DM_read_data_mem_latched_20), 
        .d(DM_read_data_mem_20), .g(n100) );
    latn_2 DM_read_data_mem_latched_reg_21 ( .q(DM_read_data_mem_latched_21), 
        .d(DM_read_data_mem_21), .g(n100) );
    latn_2 DM_read_data_mem_latched_reg_22 ( .q(DM_read_data_mem_latched_22), 
        .d(DM_read_data_mem_22), .g(n100) );
    latn_2 DM_read_data_mem_latched_reg_23 ( .q(DM_read_data_mem_latched_23), 
        .d(DM_read_data_mem_23), .g(n100) );
    latn_2 DM_read_data_mem_latched_reg_24 ( .q(DM_read_data_mem_latched_24), 
        .d(DM_read_data_mem_24), .g(n100) );
    latn_2 DM_read_data_mem_latched_reg_25 ( .q(DM_read_data_mem_latched_25), 
        .d(DM_read_data_mem_25), .g(n100) );
    latn_2 DM_read_data_mem_latched_reg_26 ( .q(DM_read_data_mem_latched_26), 
        .d(DM_read_data_mem_26), .g(n100) );
    latn_2 DM_read_data_mem_latched_reg_27 ( .q(DM_read_data_mem_latched_27), 
        .d(DM_read_data_mem_27), .g(n100) );
    latn_2 DM_read_data_mem_latched_reg_28 ( .q(DM_read_data_mem_latched_28), 
        .d(DM_read_data_mem_28), .g(n100) );
    latn_2 DM_read_data_mem_latched_reg_29 ( .q(DM_read_data_mem_latched_29), 
        .d(DM_read_data_mem_29), .g(n100) );
    latn_2 DM_read_data_mem_latched_reg_30 ( .q(DM_read_data_mem_latched_30), 
        .d(DM_read_data_mem_30), .g(n100) );
    latn_2 DM_read_data_mem_latched_reg_31 ( .q(DM_read_data_mem_latched_31), 
        .d(DM_read_data_mem_31), .g(n100) );
    latn_2 IM_read_data_mem_latched_reg_0 ( .q(IM_read_data_mem_latched_0), 
        .d(IM_read_data_mem_0), .g(n102) );
    latn_2 IM_read_data_mem_latched_reg_1 ( .q(IM_read_data_mem_latched_1), 
        .d(IM_read_data_mem_1), .g(n102) );
    latn_2 IM_read_data_mem_latched_reg_2 ( .q(IM_read_data_mem_latched_2), 
        .d(IM_read_data_mem_2), .g(n102) );
    latn_2 IM_read_data_mem_latched_reg_3 ( .q(IM_read_data_mem_latched_3), 
        .d(IM_read_data_mem_3), .g(n102) );
    latn_2 IM_read_data_mem_latched_reg_4 ( .q(IM_read_data_mem_latched_4), 
        .d(IM_read_data_mem_4), .g(n102) );
    latn_2 IM_read_data_mem_latched_reg_5 ( .q(IM_read_data_mem_latched_5), 
        .d(IM_read_data_mem_5), .g(n102) );
    latn_2 IM_read_data_mem_latched_reg_6 ( .q(IM_read_data_mem_latched_6), 
        .d(IM_read_data_mem_6), .g(n102) );
    latn_2 IM_read_data_mem_latched_reg_7 ( .q(IM_read_data_mem_latched_7), 
        .d(IM_read_data_mem_7), .g(n102) );
    latn_2 IM_read_data_mem_latched_reg_8 ( .q(IM_read_data_mem_latched_8), 
        .d(IM_read_data_mem_8), .g(n102) );
    latn_2 IM_read_data_mem_latched_reg_9 ( .q(IM_read_data_mem_latched_9), 
        .d(IM_read_data_mem_9), .g(n102) );
    latn_2 IM_read_data_mem_latched_reg_10 ( .q(IM_read_data_mem_latched_10), 
        .d(IM_read_data_mem_10), .g(n102) );
    latn_2 IM_read_data_mem_latched_reg_11 ( .q(IM_read_data_mem_latched_11), 
        .d(IM_read_data_mem_11), .g(n102) );
    latn_2 IM_read_data_mem_latched_reg_12 ( .q(IM_read_data_mem_latched_12), 
        .d(IM_read_data_mem_12), .g(n102) );
    latn_2 IM_read_data_mem_latched_reg_13 ( .q(IM_read_data_mem_latched_13), 
        .d(IM_read_data_mem_13), .g(n102) );
    latn_2 IM_read_data_mem_latched_reg_14 ( .q(IM_read_data_mem_latched_14), 
        .d(IM_read_data_mem_14), .g(n102) );
    latn_2 IM_read_data_mem_latched_reg_15 ( .q(IM_read_data_mem_latched_15), 
        .d(IM_read_data_mem_15), .g(n102) );
    latn_2 IM_read_data_mem_latched_reg_16 ( .q(IM_read_data_mem_latched_16), 
        .d(IM_read_data_mem_16), .g(n102) );
    latn_2 IM_read_data_mem_latched_reg_17 ( .q(IM_read_data_mem_latched_17), 
        .d(IM_read_data_mem_17), .g(n102) );
    latn_2 IM_read_data_mem_latched_reg_18 ( .q(IM_read_data_mem_latched_18), 
        .d(IM_read_data_mem_18), .g(n102) );
    latn_2 IM_read_data_mem_latched_reg_19 ( .q(IM_read_data_mem_latched_19), 
        .d(IM_read_data_mem_19), .g(n102) );
    latn_2 IM_read_data_mem_latched_reg_20 ( .q(IM_read_data_mem_latched_20), 
        .d(IM_read_data_mem_20), .g(n102) );
    latn_2 IM_read_data_mem_latched_reg_21 ( .q(IM_read_data_mem_latched_21), 
        .d(IM_read_data_mem_21), .g(n102) );
    latn_2 IM_read_data_mem_latched_reg_22 ( .q(IM_read_data_mem_latched_22), 
        .d(IM_read_data_mem_22), .g(n102) );
    latn_2 IM_read_data_mem_latched_reg_23 ( .q(IM_read_data_mem_latched_23), 
        .d(IM_read_data_mem_23), .g(n102) );
    latn_2 IM_read_data_mem_latched_reg_24 ( .q(IM_read_data_mem_latched_24), 
        .d(IM_read_data_mem_24), .g(n102) );
    latn_2 IM_read_data_mem_latched_reg_25 ( .q(IM_read_data_mem_latched_25), 
        .d(IM_read_data_mem_25), .g(n102) );
    latn_2 IM_read_data_mem_latched_reg_26 ( .q(IM_read_data_mem_latched_26), 
        .d(IM_read_data_mem_26), .g(n102) );
    latn_2 IM_read_data_mem_latched_reg_27 ( .q(IM_read_data_mem_latched_27), 
        .d(IM_read_data_mem_27), .g(n102) );
    latn_2 IM_read_data_mem_latched_reg_28 ( .q(IM_read_data_mem_latched_28), 
        .d(IM_read_data_mem_28), .g(n102) );
    latn_2 IM_read_data_mem_latched_reg_29 ( .q(IM_read_data_mem_latched_29), 
        .d(IM_read_data_mem_29), .g(n102) );
    latn_2 IM_read_data_mem_latched_reg_30 ( .q(IM_read_data_mem_latched_30), 
        .d(IM_read_data_mem_30), .g(n102) );
    latn_2 IM_read_data_mem_latched_reg_31 ( .q(IM_read_data_mem_latched_31), 
        .d(IM_read_data_mem_31), .g(n102) );
    and2_1 U215 ( .x(n37), .a(im_grant_chain), .b(n139) );
    and2_1 U216 ( .x(n40), .a(n139), .b(n142) );
    mux2_2 U217 ( .x(n41), .d0(DM_read_data_mem_latched_9), .sl(dp_not_local), 
        .d1(dp_r_dat_9) );
    mux2_2 U218 ( .x(n42), .d0(DM_read_data_mem_latched_8), .sl(dp_not_local), 
        .d1(dp_r_dat_8) );
    mux2_2 U219 ( .x(n43), .d0(DM_read_data_mem_latched_7), .sl(dp_not_local), 
        .d1(dp_r_dat_7) );
    mux2_2 U220 ( .x(n44), .d0(DM_read_data_mem_latched_6), .sl(dp_not_local), 
        .d1(dp_r_dat_6) );
    mux2_2 U221 ( .x(n45), .d0(DM_read_data_mem_latched_5), .sl(dp_not_local), 
        .d1(dp_r_dat_5) );
    mux2_2 U222 ( .x(n46), .d0(DM_read_data_mem_latched_4), .sl(dp_not_local), 
        .d1(dp_r_dat_4) );
    mux2_2 U223 ( .x(n47), .d0(DM_read_data_mem_latched_31), .sl(dp_not_local), 
        .d1(dp_r_dat_31) );
    mux2_2 U224 ( .x(n48), .d0(DM_read_data_mem_latched_30), .sl(dp_not_local), 
        .d1(dp_r_dat_30) );
    mux2_2 U225 ( .x(n49), .d0(DM_read_data_mem_latched_3), .sl(dp_not_local), 
        .d1(dp_r_dat_3) );
    mux2_2 U226 ( .x(n50), .d0(DM_read_data_mem_latched_29), .sl(dp_not_local), 
        .d1(dp_r_dat_29) );
    mux2_2 U227 ( .x(n51), .d0(DM_read_data_mem_latched_28), .sl(dp_not_local), 
        .d1(dp_r_dat_28) );
    mux2_2 U228 ( .x(n52), .d0(DM_read_data_mem_latched_27), .sl(dp_not_local), 
        .d1(dp_r_dat_27) );
    mux2_2 U229 ( .x(n53), .d0(DM_read_data_mem_latched_26), .sl(dp_not_local), 
        .d1(dp_r_dat_26) );
    mux2_2 U230 ( .x(n54), .d0(DM_read_data_mem_latched_25), .sl(dp_not_local), 
        .d1(dp_r_dat_25) );
    mux2_2 U231 ( .x(n81), .d0(DM_read_data_mem_latched_24), .sl(n109), .d1(
        dp_r_dat_24) );
    mux2_2 U232 ( .x(n82), .d0(DM_read_data_mem_latched_23), .sl(dp_not_local), 
        .d1(dp_r_dat_23) );
    mux2_2 U233 ( .x(n83), .d0(DM_read_data_mem_latched_22), .sl(dp_not_local), 
        .d1(dp_r_dat_22) );
    mux2_2 U234 ( .x(n84), .d0(DM_read_data_mem_latched_21), .sl(dp_not_local), 
        .d1(dp_r_dat_21) );
    mux2_2 U235 ( .x(n85), .d0(DM_read_data_mem_latched_20), .sl(dp_not_local), 
        .d1(dp_r_dat_20) );
    mux2_2 U236 ( .x(n86), .d0(DM_read_data_mem_latched_2), .sl(dp_not_local), 
        .d1(dp_r_dat_2) );
    mux2_2 U237 ( .x(n87), .d0(DM_read_data_mem_latched_19), .sl(dp_not_local), 
        .d1(dp_r_dat_19) );
    mux2_2 U238 ( .x(n88), .d0(DM_read_data_mem_latched_18), .sl(dp_not_local), 
        .d1(dp_r_dat_18) );
    mux2_2 U239 ( .x(n89), .d0(DM_read_data_mem_latched_17), .sl(dp_not_local), 
        .d1(dp_r_dat_17) );
    mux2_2 U240 ( .x(n90), .d0(DM_read_data_mem_latched_16), .sl(dp_not_local), 
        .d1(dp_r_dat_16) );
    mux2_2 U241 ( .x(n91), .d0(DM_read_data_mem_latched_15), .sl(dp_not_local), 
        .d1(dp_r_dat_15) );
    mux2_2 U242 ( .x(n92), .d0(DM_read_data_mem_latched_14), .sl(dp_not_local), 
        .d1(dp_r_dat_14) );
    mux2_2 U243 ( .x(n93), .d0(DM_read_data_mem_latched_13), .sl(dp_not_local), 
        .d1(dp_r_dat_13) );
    mux2_2 U244 ( .x(n94), .d0(DM_read_data_mem_latched_12), .sl(dp_not_local), 
        .d1(dp_r_dat_12) );
    mux2_2 U245 ( .x(n95), .d0(DM_read_data_mem_latched_11), .sl(dp_not_local), 
        .d1(dp_r_dat_11) );
    mux2_2 U246 ( .x(n96), .d0(DM_read_data_mem_latched_10), .sl(dp_not_local), 
        .d1(dp_r_dat_10) );
    mux2_2 U247 ( .x(n97), .d0(DM_read_data_mem_latched_1), .sl(dp_not_local), 
        .d1(dp_r_dat_1) );
    mux2_2 U248 ( .x(n98), .d0(DM_read_data_mem_latched_0), .sl(dp_not_local), 
        .d1(dp_r_dat_0) );
    buf_3 U249 ( .x(n160), .a(inst_ram_load) );
    inv_2 U250 ( .x(n102), .a(n101) );
    inv_2 U251 ( .x(n100), .a(n99) );
    and2_1 U252 ( .x(n99), .a(N1107), .b(DM_complete_latched) );
    and2_1 U253 ( .x(n101), .a(N1107), .b(IM_complete_latched) );
    mux2_1 U254 ( .x(n103), .d0(reset_DLX_d_ff2), .sl(N1107), .d1(reset_DLX_d)
         );
    and2_1 U255 ( .x(n104), .a(N1107), .b(n139) );
    inv_1 U256 ( .x(n105), .a(n118) );
    inv_16 U257 ( .x(n106), .a(n105) );
    inv_0 U258 ( .x(n118), .a(n117) );
    buf_7 U259 ( .x(n107), .a(wish_we_o) );
    inv_0 U260 ( .x(n108), .a(n151) );
    inv_2 U261 ( .x(ip_not_local), .a(n151) );
    nand2_2 U262 ( .x(n151), .a(Ctrl__IFinst___Regs_1__ro), .b(n137) );
    inv_0 U263 ( .x(n109), .a(n152) );
    inv_2 U264 ( .x(dp_not_local), .a(n152) );
    nand3_1 U265 ( .x(n152), .a(n125), .b(n126), .c(Ctrl__EXinst___Regs_1__ro)
         );
    inv_0 U266 ( .x(n110), .a(n147) );
    inv_2 U267 ( .x(n130), .a(n147) );
    nand2_2 U268 ( .x(n147), .a(dm_grant_chain), .b(n139) );
    buf_3 U269 ( .x(n111), .a(memory_load_enable) );
    buf_3 U270 ( .x(n157), .a(memory_load_enable) );
    buf_3 U271 ( .x(n158), .a(memory_load_enable) );
    inv_1 U272 ( .x(n123), .a(N1107) );
    and3_1 U273 ( .x(n112), .a(N1107), .b(n139), .c(DM_start) );
    inv_0 U274 ( .x(n113), .a(n112) );
    nand2_0 U275 ( .x(DMem_clk), .a(n133), .b(n113) );
    nand2_0 U276 ( .x(n134), .a(IM_start), .b(n104) );
    nand2_0 U277 ( .x(IMem_clk), .a(n133), .b(n134) );
    inv_2 U278 ( .x(n139), .a(n158) );
    inv_0 U279 ( .x(n114), .a(n123) );
    inv_1 U280 ( .x(n115), .a(global_g2) );
    inv_16 U281 ( .x(n116), .a(n115) );
    inv_1 U282 ( .x(n117), .a(global_g1) );
    inv_1 U283 ( .x(n119), .a(n122) );
    inv_16 U284 ( .x(n120), .a(n119) );
    inv_0 U285 ( .x(n122), .a(n121) );
    inv_1 U286 ( .x(n121), .a(test_se) );
    inv_0 U287 ( .x(n136), .a(n114) );
    nand2i_4 U38 ( .x(IM_start), .a(im_grant_local_d), .b(n39) );
    nand2i_4 U34 ( .x(DM_start), .a(dm_grant_local_d), .b(n38) );
    and2_8 C1247 ( .x(ip_r_ack), .a(Ctrl__IFinst___Regs_1__ai), .b(ip_complete
        ) );
    and2_8 C1271 ( .x(dp_r_ack), .a(Ctrl__MEMinst___Regs_1__ai), .b(
        dp_complete) );
    and2_8 C1278 ( .x(_40_net_), .a(N1429), .b(nrst) );
    and2_8 C1280 ( .x(_41_net_), .a(ip_local), .b(N315) );
    and2_8 C1286 ( .x(im_r_req), .a(IM_complete), .b(im_grant_chain_d) );
    and2_8 C1288 ( .x(_43_net_), .a(dp_local), .b(N597) );
    and2_8 C1291 ( .x(_45_net_), .a(N1431), .b(nrst) );
    and2_8 C1299 ( .x(dm_r_req), .a(DM_complete), .b(dm_grant_chain_d) );
endmodule

