// Xilinx Verilog netlist produced by netgen application (version G.29)
// Command      : -intstyle ise -s 7 -pcf DLX_top.pcf -ngm DLX_top.ngm -w -ofmt verilog -sim DLX_top.ncd DLX_top_timesim.v 
// Input file   : DLX_top.ncd
// Output file  : DLX_top_timesim.v
// Design name  : DLX_top
// # of Modules : 1
// Xilinx       : /usr/local/vlsi/Xilinx-ISE-6.2
// Device       : 2s200epq208-7 (PRODUCTION 1.17 2003-12-13)

// This verilog netlist is a simulation model and uses simulation 
// primitives which may not represent the true implementation of the 
// device, however the netlist is functionally correct and should not 
// be modified. This file cannot be synthesized and should only be used 
// with supported simulation tools.

`timescale 1 ns/1 ps

module DLX_top (
  stall, branch_sig, hsync, clk_IF_del, DM_write, DM_write_data_0, DM_read, clk_MEM, PIPEEMPTY, vsync, clk_IF, clk_ID, clk_EX, CLI, clk_DM, INT, 
STOP_fetch, clk_vga, FREEZE, reset, DM_addr_eff, mask, red, NPC_eff, IR_MSB, green, blue, delay_selectRF, delay_selectIF, delay_selectID, 
delay_selectEX, delay_selectDM, delay_selectMEM
);
  output stall;
  output branch_sig;
  output hsync;
  output clk_IF_del;
  output DM_write;
  output DM_write_data_0;
  output DM_read;
  output clk_MEM;
  output PIPEEMPTY;
  output vsync;
  output clk_IF;
  output clk_ID;
  output clk_EX;
  output CLI;
  output clk_DM;
  input INT;
  input STOP_fetch;
  input clk_vga;
  input FREEZE;
  input reset;
  output [14 : 0] DM_addr_eff;
  output [3 : 0] mask;
  output [1 : 0] red;
  output [15 : 0] NPC_eff;
  output [7 : 0] IR_MSB;
  output [2 : 0] green;
  output [2 : 0] blue;
  input [1 : 0] delay_selectRF;
  input [1 : 0] delay_selectIF;
  input [1 : 0] delay_selectID;
  input [1 : 0] delay_selectEX;
  input [1 : 0] delay_selectDM;
  input [1 : 0] delay_selectMEM;
  wire mask_1_OBUF;
  wire DLX_clk_EX;
  wire DLX_EXinst__n0012;
  wire reset_IBUF;
  wire mask_2_OBUF;
  wire PIPEEMPTY_OBUF;
  wire DLX_clk_IF_del;
  wire N116776;
  wire N113314;
  wire N112968;
  wire N115578;
  wire N115216;
  wire DLX_clk_ID;
  wire DLX_IDinst__n0422;
  wire N110516;
  wire reset_IBUF_5;
  wire clk_DM_OBUF;
  wire DLX_clk_IF;
  wire clkdiv_vga;
  wire vga_top_vga1__n0010;
  wire green_0_OBUF;
  wire green_1_OBUF;
  wire green_2_OBUF;
  wire red_0_OBUF;
  wire red_1_OBUF;
  wire reset_IBUF_2;
  wire DLX_IDinst__n0441;
  wire N110648;
  wire reset_IBUF_3;
  wire DLX_IDinst__n0421;
  wire DLX_IDinst__n0124;
  wire INT_IBUF;
  wire N125635;
  wire N124056;
  wire N123038;
  wire N120114;
  wire N113660;
  wire N116396;
  wire N115984;
  wire N112616;
  wire N111878;
  wire N117154;
  wire vga_top_vga1__n0011;
  wire FREEZE_IBUF;
  wire IR_MSB_0_OBUF;
  wire IR_MSB_1_OBUF;
  wire IR_MSB_2_OBUF;
  wire IR_MSB_3_OBUF;
  wire IR_MSB_4_OBUF;
  wire IR_MSB_5_OBUF;
  wire IR_MSB_6_OBUF;
  wire IR_MSB_7_OBUF;
  wire delay_selectDM_0_IBUF;
  wire delay_selectDM_1_IBUF;
  wire delay_selectID_0_IBUF;
  wire delay_selectID_1_IBUF;
  wire DLX_MEMlc_master_ctrlMEM_l;
  wire delay_selectIF_0_IBUF;
  wire delay_selectIF_1_IBUF;
  wire delay_selectMEM_0_IBUF;
  wire delay_selectMEM_1_IBUF;
  wire blue_0_OBUF;
  wire blue_1_OBUF;
  wire blue_2_OBUF;
  wire STOP_fetch_IBUF;
  wire delay_selectEX_0_IBUF;
  wire delay_selectEX_1_IBUF;
  wire mask_0_OBUF;
  wire delay_selectRF_0_IBUF;
  wire delay_selectRF_1_IBUF;
  wire DLX_EXinst__n0011;
  wire mask_3_OBUF;
  wire clkbuf;
  wire clk0;
  wire clkdivub;
  wire clk0buf;
  wire DLX_ackin_ID;
  wire DLX_ackin_EX;
  wire DLX_IDinst__n0000;
  wire DLX_IDinst__n0410;
  wire DLX_IDinst__n0002;
  wire DLX_MEMinst_reg_write_MEM;
  wire GLOBAL_LOGIC0;
  wire DLX_IDinst__n0003;
  wire DLX_IDinst__n0004;
  wire DLX_EXinst_mem_write_EX;
  wire reset_IBUF_1;
  wire vga_top_vga1_Madd_addressout_inst_lut2_331;
  wire DLX_IDinst_reg_out_B_3_1;
  wire N111221;
  wire CHOICE3139;
  wire CHOICE3145;
  wire CHOICE3152;
  wire N108593;
  wire DLX_IDinst_reg_out_B_2_1;
  wire CHOICE1306;
  wire CHOICE1312;
  wire DLX_EXinst_N66494;
  wire \DLX_EXinst_Mshift__n0026_Sh[21] ;
  wire \DLX_EXinst_Mshift__n0026_Sh[29] ;
  wire CHOICE3132;
  wire CHOICE3032;
  wire CHOICE3038;
  wire CHOICE3045;
  wire N107934;
  wire N126675;
  wire DLX_IDinst_N70909;
  wire DLX_IDinst__n0377;
  wire DLX_IDinst_N70985;
  wire CHOICE3311;
  wire DLX_EXinst_N66202;
  wire CHOICE1042;
  wire CHOICE1048;
  wire CHOICE5189;
  wire N97960;
  wire N126636;
  wire CHOICE1402;
  wire DLX_IFlc_md_wint30;
  wire DLX_IFlc_md_wint40;
  wire DLX_IFlc_md_wint26;
  wire DLX_IFlc_md_wint34;
  wire DLX_IFlc_md_outp2;
  wire DLX_IDlc_md_wint30;
  wire DLX_IDlc_md_wint40;
  wire DLX_IDlc_md_wint26;
  wire DLX_IDlc_md_wint34;
  wire DLX_IDlc_md_outp2;
  wire DLX_EXlc_md_wint30;
  wire DLX_EXlc_md_wint40;
  wire DLX_EXlc_md_wint26;
  wire DLX_EXlc_md_wint34;
  wire DLX_EXlc_md_outp2;
  wire DLX_EXinst_N62986;
  wire DLX_EXinst_N63489;
  wire DLX_EXinst_N65165;
  wire DLX_EXinst_N64474;
  wire CHOICE5509;
  wire DLX_MEMlc_md_wint10;
  wire DLX_MEMlc_md_wint20;
  wire DLX_MEMlc_md_wint8;
  wire DLX_MEMlc_md_wint14;
  wire DLX_MEMlc_md_outp2;
  wire N93279;
  wire DLX_EXinst_N62821;
  wire CHOICE5341;
  wire N97665;
  wire N126486;
  wire DLX_IDinst__n0135;
  wire N98613;
  wire DLX_IDinst_N70647;
  wire N98420;
  wire DLX_IDinst__n0136;
  wire DLX_IDinst__n0344;
  wire DLX_IDinst__n0347;
  wire DLX_IDinst__n0345;
  wire DLX_IDinst_N69963;
  wire DM_delay_inst_wint26;
  wire DM_delay_inst_wint40;
  wire DM_delay_inst_wint20;
  wire DM_delay_inst_wint34;
  wire clk_EX_del;
  wire DLX_IFinst__n0000;
  wire DLX_IDinst_branch_sig;
  wire DLX_IFinst_stalled;
  wire DLX_RF_delay_inst_wint20;
  wire DLX_RF_delay_inst_wint30;
  wire DLX_RF_delay_inst_wint14;
  wire DLX_RF_delay_inst_wint24;
  wire \DLX_EXinst_Mshift__n0025_Sh[8] ;
  wire CHOICE1084;
  wire CHOICE1078;
  wire \DLX_EXinst_Mshift__n0025_Sh[40] ;
  wire N94305;
  wire DLX_EXinst_N62851;
  wire \DLX_EXinst_Mshift__n0025_Sh[11] ;
  wire CHOICE1060;
  wire CHOICE1054;
  wire \DLX_EXinst_Mshift__n0025_Sh[43] ;
  wire N93331;
  wire DLX_EXinst_N62826;
  wire CHOICE5264;
  wire N98032;
  wire N126560;
  wire DLX_EXinst_N62631;
  wire DLX_EXinst_N64319;
  wire DLX_EXinst_N62727;
  wire N96153;
  wire CHOICE5866;
  wire CHOICE5871;
  wire \DLX_IDinst_Imm[5] ;
  wire N110065;
  wire DLX_EXinst_N63185;
  wire DLX_EXinst_N64565;
  wire DLX_EXinst_N62715;
  wire CHOICE5100;
  wire \DLX_EXinst_Mshift__n0027_Sh[4] ;
  wire \DLX_EXinst_Mshift__n0027_Sh[12] ;
  wire \DLX_EXinst_Mshift__n0027_Sh[8] ;
  wire N93179;
  wire CHOICE5125;
  wire DLX_EXinst__n0081;
  wire \DLX_EXinst_Mshift__n0027_Sh[9] ;
  wire \DLX_EXinst_Mshift__n0027_Sh[5] ;
  wire N93127;
  wire \DLX_EXinst_Mshift__n0027_Sh[13] ;
  wire CHOICE5598;
  wire CHOICE1270;
  wire CHOICE1276;
  wire \DLX_EXinst_Mshift__n0028_Sh[8] ;
  wire CHOICE5969;
  wire CHOICE5973;
  wire DLX_EXinst__n0030_1;
  wire CHOICE1771;
  wire CHOICE1919;
  wire CHOICE1926;
  wire CHOICE5696;
  wire CHOICE5706;
  wire CHOICE5709;
  wire \DLX_EXinst_Mshift__n0027_Sh[10] ;
  wire \DLX_EXinst_Mshift__n0027_Sh[6] ;
  wire N93229;
  wire \DLX_EXinst_Mshift__n0027_Sh[14] ;
  wire CHOICE5432;
  wire DLX_EXinst_N63036;
  wire DLX_EXinst_N64904;
  wire DLX_EXinst_N63329;
  wire DLX_EXinst_N64255;
  wire CHOICE5540;
  wire \DLX_EXinst_Mshift__n0027_Sh[11] ;
  wire \DLX_EXinst_Mshift__n0027_Sh[7] ;
  wire \DLX_EXinst_Mshift__n0027_Sh[19] ;
  wire \DLX_EXinst_Mshift__n0027_Sh[15] ;
  wire CHOICE4965;
  wire DLX_IDinst_IR_function_field_2_1;
  wire DLX_IDinst_IR_function_field_3_1;
  wire DLX_EXinst_N63129;
  wire DLX_EXinst_N66421;
  wire N125971;
  wire N101537;
  wire DLX_EXinst_N62740;
  wire \DLX_EXinst_Mshift__n0026_Sh[60] ;
  wire N95810;
  wire DLX_EXinst_N63157;
  wire DLX_EXinst_N66431;
  wire N126006;
  wire CHOICE2965;
  wire \DLX_EXinst_Mshift__n0024_Sh[61] ;
  wire DLX_EXinst_N62936;
  wire CHOICE3085;
  wire CHOICE3097;
  wire DLX_EXinst_N63374;
  wire CHOICE1184;
  wire DLX_EXinst_N62896;
  wire DLX_EXinst_N62876;
  wire N97089;
  wire DLX_EXinst_N63066;
  wire DLX_EXinst_N63780;
  wire DLX_EXinst_N63046;
  wire DLX_EXinst_N63419;
  wire N97449;
  wire DLX_EXinst_N63379;
  wire DLX_EXinst_N63274;
  wire CHOICE1825;
  wire DLX_EXinst_N62881;
  wire N100843;
  wire CHOICE1162;
  wire CHOICE1168;
  wire \DLX_EXinst_Mshift__n0026_Sh[11] ;
  wire CHOICE5073;
  wire CHOICE5077;
  wire DLX_EXinst_N63016;
  wire DLX_EXinst_N63279;
  wire DLX_EXinst_N62996;
  wire DLX_EXinst_N63504;
  wire N97305;
  wire Mmux__COND_2__net2;
  wire DLX_EXinst_N63429;
  wire DLX_EXinst_N63061;
  wire DLX_EXinst_N63409;
  wire DLX_EXinst_N63041;
  wire N97375;
  wire DLX_EXinst_N62891;
  wire DLX_EXinst_N62871;
  wire N97161;
  wire DLX_EXinst_N62796;
  wire DLX_EXinst_N63459;
  wire DLX_EXinst_N63309;
  wire CHOICE1838;
  wire N100919;
  wire DLX_EXinst_N64334;
  wire DLX_EXinst_N62971;
  wire N101009;
  wire \DLX_EXinst_Mshift__n0024_Sh[27] ;
  wire N101253;
  wire DLX_EXinst_N63499;
  wire DLX_EXinst_N63334;
  wire DLX_EXinst_N62921;
  wire N97521;
  wire CHOICE3196;
  wire CHOICE3198;
  wire \DLX_EXinst_Mshift__n0023_Sh[27] ;
  wire CHOICE2542;
  wire DLX_IDinst_IR_function_field_0_1;
  wire DLX_IDinst_IR_function_field_1_1;
  wire CHOICE1012;
  wire CHOICE1006;
  wire \DLX_EXinst_Mshift__n0027_Sh[40] ;
  wire \DLX_EXinst_Mshift__n0023_Sh[61] ;
  wire DLX_EXinst_N62966;
  wire CHOICE3112;
  wire CHOICE3124;
  wire \DLX_EXinst_Mshift__n0026_Sh[17] ;
  wire \DLX_EXinst_Mshift__n0023_Sh[9] ;
  wire \DLX_EXinst_Mshift__n0026_Sh[13] ;
  wire CHOICE4587;
  wire N94155;
  wire DLX_EXinst_N63479;
  wire \DLX_EXinst_Mshift__n0027_Sh[2] ;
  wire \DLX_EXinst_Mshift__n0027_Sh[42] ;
  wire DLX_EXinst_N62766;
  wire CHOICE1000;
  wire CHOICE994;
  wire \DLX_EXinst_Mshift__n0027_Sh[43] ;
  wire CHOICE2980;
  wire N126268;
  wire DLX_EXinst_N62721;
  wire DLX_EXinst_N65090;
  wire \DLX_EXinst_Mshift__n0026_Sh[24] ;
  wire DLX_EXinst_N64500;
  wire DLX_EXinst_N62709;
  wire N93799;
  wire \DLX_EXinst_Mshift__n0028_Sh[59] ;
  wire \DLX_EXinst_Mshift__n0026_Sh[18] ;
  wire \DLX_EXinst_Mshift__n0026_Sh[22] ;
  wire \DLX_EXinst_Mshift__n0026_Sh[10] ;
  wire \DLX_EXinst_Mshift__n0026_Sh[14] ;
  wire CHOICE4531;
  wire DLX_EXinst_N62916;
  wire N93695;
  wire DLX_EXinst__n0048;
  wire N126169;
  wire N126500;
  wire DLX_EXinst_N62911;
  wire N93747;
  wire CHOICE5291;
  wire N97017;
  wire CHOICE5297;
  wire DLX_EXinst_N62981;
  wire DLX_EXinst_N65135;
  wire N127444;
  wire N93383;
  wire DLX_EXinst_N62831;
  wire N126154;
  wire CHOICE5815;
  wire DLX_EXinst__n0079;
  wire CHOICE5839;
  wire DLX_EXinst__n0078;
  wire \DLX_IDinst_Imm[31] ;
  wire DLX_EXinst__n0080;
  wire CHOICE5842;
  wire DLX_EXinst_N64914;
  wire CHOICE5162;
  wire CHOICE5166;
  wire CHOICE5140;
  wire \DLX_EXinst_Mshift__n0025_Sh[9] ;
  wire \DLX_EXinst_Mshift__n0025_Sh[5] ;
  wire N93487;
  wire \DLX_EXinst_Mshift__n0025_Sh[13] ;
  wire CHOICE5637;
  wire \DLX_EXinst_Mshift__n0025_Sh[10] ;
  wire \DLX_EXinst_Mshift__n0025_Sh[6] ;
  wire N93537;
  wire \DLX_EXinst_Mshift__n0025_Sh[14] ;
  wire CHOICE5471;
  wire DLX_EXinst_N63920;
  wire CHOICE4990;
  wire CHOICE4994;
  wire DLX_EXinst_N62901;
  wire N93587;
  wire CHOICE5216;
  wire CHOICE5222;
  wire DLX_EXinst_N62906;
  wire N93641;
  wire CHOICE5368;
  wire CHOICE5374;
  wire DLX_EXinst_N63494;
  wire DLX_EXinst_N64909;
  wire N127440;
  wire CHOICE3007;
  wire N126272;
  wire vram_out_vga_eff;
  wire vga_top_vga1_Madd_addressout_inst_cy_466;
  wire vga_top_vga1_Madd_addressout_inst_cy_468;
  wire vga_top_vga1_Mmult__n0043_inst_lut2_317;
  wire vga_top_vga1_Madd_addressout_inst_cy_470;
  wire vga_top_vga1_Mmult__n0043_inst_lut2_318;
  wire vga_top_vga1_Mmult__n0043_inst_lut2_319;
  wire vga_top_vga1_Madd_addressout_inst_cy_472;
  wire vga_top_vga1_Mmult__n0043_inst_lut2_320;
  wire vga_top_vga1_Mmult__n0043_inst_lut2_321;
  wire vga_top_vga1_Mmult__n0043_inst_lut2_322;
  wire vga_top_vga1_Mmult__n0043_inst_lut2_323;
  wire DLX_EXinst_Mcompar__n0057_inst_cy_135;
  wire DLX_EXinst_Mcompar__n0057_inst_cy_137;
  wire DLX_EXinst_Mcompar__n0057_inst_cy_139;
  wire DLX_EXinst_Mcompar__n0057_inst_cy_141;
  wire DLX_EXinst_Mcompar__n0057_inst_cy_143;
  wire DLX_EXinst_Mcompar__n0057_inst_cy_145;
  wire DLX_EXinst_Mcompar__n0057_inst_cy_147;
  wire DLX_EXinst_Mcompar__n0057_inst_cy_149;
  wire DLX_EXinst_Mcompar__n0057_inst_cy_151;
  wire DLX_EXinst_Mcompar__n0057_inst_cy_153;
  wire DLX_EXinst_Mcompar__n0057_inst_cy_155;
  wire DLX_EXinst_Mcompar__n0057_inst_cy_157;
  wire DLX_EXinst_Mcompar__n0057_inst_cy_159;
  wire DLX_EXinst_Mcompar__n0057_inst_cy_161;
  wire DLX_EXinst_Mcompar__n0057_inst_cy_163;
  wire DLX_EXinst__n0047;
  wire DLX_EXinst__n0046;
  wire DLX_EXinst_Mcompar__n0057_inst_cy_164;
  wire CHOICE5306;
  wire DLX_IDinst_Mcompar__n0000_inst_cy_266;
  wire DLX_IDinst_Mcompar__n0073_inst_cy_263;
  wire DLX_IDinst_reg_dst;
  wire DLX_IDinst__n0073;
  wire DLX_IDinst_Mcompar__n0314_inst_cy_263;
  wire vga_top_vga1_Mmult__n0043_inst_cy_440;
  wire vga_top_vga1_Mmult__n0043_inst_cy_442;
  wire vga_top_vga1_Mmult__n0043_inst_cy_444;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_167;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_169;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_171;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_173;
  wire \DLX_IDinst_Imm[6] ;
  wire \DLX_IDinst_Imm[7] ;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_175;
  wire \DLX_IDinst_Imm[8] ;
  wire \DLX_IDinst_Imm[9] ;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_177;
  wire \DLX_IDinst_Imm[10] ;
  wire \DLX_IDinst_Imm[11] ;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_179;
  wire \DLX_IDinst_Imm[12] ;
  wire \DLX_IDinst_Imm[13] ;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_181;
  wire \DLX_IDinst_Imm[14] ;
  wire \DLX_IDinst_Imm[15] ;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_183;
  wire DLX_IDinst_Imm_31_1;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_185;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_187;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_189;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_191;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_193;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_195;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_196;
  wire N127408;
  wire DLX_EXinst_Mcompar__n0059_inst_cy_167;
  wire DLX_EXinst_Mcompar__n0059_inst_cy_169;
  wire DLX_EXinst_Mcompar__n0059_inst_cy_171;
  wire DLX_EXinst_Mcompar__n0059_inst_cy_173;
  wire DLX_EXinst_Mcompar__n0059_inst_cy_175;
  wire DLX_EXinst_Mcompar__n0059_inst_cy_177;
  wire DLX_EXinst_Mcompar__n0059_inst_cy_179;
  wire DLX_EXinst_Mcompar__n0059_inst_cy_181;
  wire DLX_EXinst_Mcompar__n0059_inst_cy_183;
  wire DLX_EXinst_Mcompar__n0059_inst_cy_185;
  wire DLX_EXinst_Mcompar__n0059_inst_cy_187;
  wire DLX_EXinst_Mcompar__n0059_inst_cy_189;
  wire DLX_EXinst_Mcompar__n0059_inst_cy_191;
  wire DLX_EXinst_Mcompar__n0059_inst_cy_193;
  wire DLX_EXinst_Mcompar__n0059_inst_cy_195;
  wire DLX_EXinst__n0045;
  wire DLX_EXinst_N64448;
  wire DLX_EXinst_Mcompar__n0059_inst_cy_196;
  wire CHOICE5313;
  wire DLX_IDinst_Mcompar__n0075_inst_cy_263;
  wire DLX_EXinst__n0149;
  wire DLX_IDinst__n0075;
  wire DLX_IDinst_Mcompar__n0315_inst_cy_263;
  wire DLX_IDinst_Madd__n0129_inst_cy_269;
  wire DLX_IDinst_Madd__n0129_inst_lut2_198;
  wire DLX_IDinst_Madd__n0129_inst_cy_271;
  wire DLX_IDinst_Madd__n0129_inst_cy_273;
  wire DLX_IDinst_Madd__n0129_inst_cy_275;
  wire DLX_IDinst_Madd__n0129_inst_cy_277;
  wire DLX_IDinst_Madd__n0129_inst_cy_279;
  wire DLX_IDinst_Madd__n0129_inst_cy_281;
  wire DLX_IDinst_Madd__n0129_inst_cy_283;
  wire DLX_IDinst_Madd__n0129_inst_cy_285;
  wire DLX_IDinst__n0456;
  wire DLX_IDinst_Madd__n0129_inst_cy_287;
  wire DLX_IDinst_Madd__n0129_inst_cy_289;
  wire DLX_IDinst_Madd__n0129_inst_cy_291;
  wire DLX_IDinst_Madd__n0129_inst_cy_293;
  wire DLX_IDinst_Madd__n0129_inst_cy_295;
  wire DLX_IDinst_Madd__n0129_inst_cy_297;
  wire DLX_IDinst_Mcompar__n0003_inst_cy_266;
  wire DLX_IDinst__n0364;
  wire DLX_IDinst_N70679;
  wire N90703;
  wire N108996;
  wire vga_top_vga1_vcounter_Madd__n0000_inst_cy_10;
  wire GLOBAL_LOGIC1;
  wire vga_top_vga1__n0007;
  wire vga_top_vga1_vcounter_Madd__n0000_inst_cy_12;
  wire vga_top_vga1_vcounter_Madd__n0000_inst_cy_14;
  wire vga_top_vga1_vcounter_Madd__n0000_inst_cy_16;
  wire vga_top_vga1_hcounter_Madd__n0000_inst_cy_20;
  wire vga_top_vga1__n0006;
  wire vga_top_vga1_hcounter_Madd__n0000_inst_cy_22;
  wire vga_top_vga1_hcounter_Madd__n0000_inst_cy_24;
  wire vga_top_vga1_hcounter_Madd__n0000_inst_cy_26;
  wire vga_top_vga1_hcounter_Madd__n0000_inst_cy_28;
  wire vga_top_vga1_hcounter_Madd__n0000_inst_cy_30;
  wire vga_top_vga1_hcounter_Madd__n0000_inst_cy_32;
  wire DLX_EXinst_Mcompar__n0085_inst_cy_103;
  wire DLX_EXinst_Mcompar__n0085_inst_cy_105;
  wire DLX_EXinst_Mcompar__n0085_inst_cy_107;
  wire DLX_EXinst_Mcompar__n0085_inst_cy_109;
  wire DLX_EXinst_Mcompar__n0085_inst_cy_111;
  wire DLX_EXinst_Mcompar__n0085_inst_cy_113;
  wire DLX_EXinst_Mcompar__n0085_inst_cy_115;
  wire DLX_EXinst__n0085;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_199;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_201;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_203;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_205;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_207;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_209;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_211;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_213;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_215;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_217;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_219;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_221;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_223;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_225;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_227;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_228;
  wire CHOICE1126;
  wire DLX_IDinst_Mcompar__n0077_inst_cy_263;
  wire DLX_IDinst__n0077;
  wire N108704;
  wire DLX_EXinst_Maddsub__n0016_inst_cy_71;
  wire DLX_EXinst_Maddsub__n0016_inst_cy_73;
  wire DLX_EXinst_Maddsub__n0016_inst_cy_75;
  wire DLX_EXinst_Maddsub__n0016_inst_cy_77;
  wire DLX_EXinst_Maddsub__n0016_inst_cy_79;
  wire DLX_EXinst_Maddsub__n0016_inst_cy_81;
  wire DLX_EXinst_Maddsub__n0016_inst_cy_83;
  wire DLX_EXinst_Maddsub__n0016_inst_cy_85;
  wire DLX_EXinst_Maddsub__n0016_inst_cy_87;
  wire DLX_EXinst_Maddsub__n0016_inst_cy_89;
  wire DLX_EXinst_Maddsub__n0016_inst_cy_91;
  wire DLX_EXinst_Maddsub__n0016_inst_cy_93;
  wire DLX_EXinst_Maddsub__n0016_inst_cy_95;
  wire DLX_EXinst_Maddsub__n0016_inst_cy_97;
  wire DLX_EXinst_Maddsub__n0016_inst_cy_99;
  wire DLX_IDinst_Mcompar__n0078_inst_cy_263;
  wire DLX_IDinst__n0078;
  wire DLX_EXinst_Mcompar__n0087_inst_cy_119;
  wire DLX_EXinst_Mcompar__n0087_inst_cy_121;
  wire DLX_EXinst_Mcompar__n0087_inst_cy_123;
  wire DLX_EXinst_Mcompar__n0087_inst_cy_125;
  wire DLX_EXinst_Mcompar__n0087_inst_cy_127;
  wire DLX_EXinst_Mcompar__n0087_inst_cy_129;
  wire DLX_EXinst_Mcompar__n0087_inst_cy_131;
  wire DLX_EXinst__n0087;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_231;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_233;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_235;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_237;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_239;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_241;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_243;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_245;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_247;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_249;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_251;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_253;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_255;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_257;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_259;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_260;
  wire CHOICE5769;
  wire vga_top_vga1_Mcompar__n0030_inst_cy_358;
  wire vga_top_vga1_Mcompar__n0030_inst_cy_360;
  wire vga_top_vga1_Mcompar__n0030_inst_cy_362;
  wire vga_top_vga1_Mcompar__n0030_inst_cy_364;
  wire vga_top_vga1_Mcompar__n0030_inst_cy_366;
  wire vga_top_vga1_Mcompar__n0030_inst_cy_368;
  wire vga_top_vga1_Mcompar__n0030_inst_cy_370;
  wire vga_top_vga1__n0030;
  wire DLX_IFinst_Madd__n0005_inst_cy_41;
  wire DLX_IFinst_Madd__n0005_inst_cy_43;
  wire DLX_IFinst_Madd__n0005_inst_cy_45;
  wire DLX_IFinst_Madd__n0005_inst_cy_47;
  wire DLX_IFinst_Madd__n0005_inst_cy_49;
  wire DLX_IFinst_Madd__n0005_inst_cy_51;
  wire DLX_IFinst_Madd__n0005_inst_cy_53;
  wire DLX_IFinst_Madd__n0005_inst_cy_55;
  wire DLX_IFinst_Madd__n0005_inst_cy_57;
  wire DLX_IFinst_Madd__n0005_inst_cy_59;
  wire DLX_IFinst_Madd__n0005_inst_cy_61;
  wire DLX_IFinst_Madd__n0005_inst_cy_63;
  wire DLX_IFinst_Madd__n0005_inst_cy_65;
  wire DLX_IFinst_Madd__n0005_inst_cy_67;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_135;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_137;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_139;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_141;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_143;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_145;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_147;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_149;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_151;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_153;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_155;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_157;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_159;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_161;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_163;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_164;
  wire CHOICE5806;
  wire vga_top_vga1_N73384;
  wire vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_1;
  wire vga_top_vga1__n0014;
  wire vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_3;
  wire vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_5;
  wire vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_7;
  wire vga_top_vga1_Mcompar__n0033_inst_cy_344;
  wire vga_top_vga1_Mcompar__n0033_inst_cy_346;
  wire vga_top_vga1_Mcompar__n0033_inst_cy_348;
  wire vga_top_vga1_Mcompar__n0033_inst_cy_350;
  wire vga_top_vga1_Mcompar__n0033_inst_cy_352;
  wire vga_top_vga1_Mcompar__n0033_inst_cy_354;
  wire vga_top_vga1__n0033;
  wire vga_top_vga1_Mcompar__n0034_inst_cy_332;
  wire vga_top_vga1_Mcompar__n0034_inst_cy_334;
  wire vga_top_vga1_Mcompar__n0034_inst_cy_336;
  wire vga_top_vga1_Mcompar__n0034_inst_cy_338;
  wire vga_top_vga1_Mcompar__n0034_inst_cy_340;
  wire vga_top_vga1__n0034;
  wire DLX_IDinst_Msub__n0128_inst_cy_300;
  wire DLX_IDinst_Msub__n0128_inst_cy_302;
  wire DLX_IDinst_Msub__n0128_inst_cy_304;
  wire DLX_IDinst_Msub__n0128_inst_cy_306;
  wire DLX_IDinst_Msub__n0128_inst_cy_308;
  wire DLX_IDinst_Msub__n0128_inst_cy_310;
  wire DLX_IDinst_Msub__n0128_inst_cy_312;
  wire DLX_IDinst_Msub__n0128_inst_cy_314;
  wire DLX_IDinst_Msub__n0128_inst_cy_316;
  wire DLX_IDinst_Msub__n0128_inst_cy_318;
  wire DLX_IDinst_Msub__n0128_inst_cy_320;
  wire DLX_IDinst_Msub__n0128_inst_cy_322;
  wire DLX_IDinst_Msub__n0128_inst_cy_324;
  wire DLX_IDinst_Msub__n0128_inst_cy_326;
  wire DLX_IDinst_Msub__n0128_inst_cy_328;
  wire DLX_EXinst_Mcompar__n0053_inst_cy_103;
  wire DLX_EXinst_Mcompar__n0053_inst_cy_105;
  wire DLX_EXinst_Mcompar__n0053_inst_cy_107;
  wire DLX_EXinst_Mcompar__n0053_inst_cy_109;
  wire DLX_EXinst_Mcompar__n0053_inst_cy_111;
  wire DLX_EXinst_Mcompar__n0053_inst_cy_113;
  wire DLX_EXinst_Mcompar__n0053_inst_cy_115;
  wire DLX_EXinst__n0053;
  wire DLX_EXinst_Mcompar__n0061_inst_cy_199;
  wire DLX_EXinst_Mcompar__n0061_inst_cy_201;
  wire DLX_EXinst_Mcompar__n0061_inst_cy_203;
  wire DLX_EXinst_Mcompar__n0061_inst_cy_205;
  wire DLX_EXinst_Mcompar__n0061_inst_cy_207;
  wire DLX_EXinst_Mcompar__n0061_inst_cy_209;
  wire DLX_EXinst_Mcompar__n0061_inst_cy_211;
  wire DLX_EXinst_Mcompar__n0061_inst_cy_213;
  wire DLX_EXinst_Mcompar__n0061_inst_cy_215;
  wire DLX_EXinst_Mcompar__n0061_inst_cy_217;
  wire DLX_EXinst_Mcompar__n0061_inst_cy_219;
  wire DLX_EXinst_Mcompar__n0061_inst_cy_221;
  wire DLX_EXinst_Mcompar__n0061_inst_cy_223;
  wire DLX_EXinst_Mcompar__n0061_inst_cy_225;
  wire DLX_EXinst_Mcompar__n0061_inst_cy_227;
  wire DLX_EXinst_N66271;
  wire DLX_EXinst_Mcompar__n0061_inst_cy_228;
  wire vga_top_vga1_Mcompar__n0029_inst_cy_374;
  wire vga_top_vga1_Mcompar__n0029_inst_cy_376;
  wire vga_top_vga1_Mcompar__n0029_inst_cy_378;
  wire vga_top_vga1__n0029;
  wire vga_top_vga1_Mcompar__n0037_inst_cy_475;
  wire vga_top_vga1_Mcompar__n0037_inst_cy_477;
  wire vga_top_vga1__n0037;
  wire DLX_EXinst_Mcompar__n0055_inst_cy_119;
  wire DLX_EXinst_Mcompar__n0055_inst_cy_121;
  wire DLX_EXinst_Mcompar__n0055_inst_cy_123;
  wire DLX_EXinst_Mcompar__n0055_inst_cy_125;
  wire DLX_EXinst_Mcompar__n0055_inst_cy_127;
  wire DLX_EXinst_Mcompar__n0055_inst_cy_129;
  wire DLX_EXinst_Mcompar__n0055_inst_cy_131;
  wire DLX_EXinst__n0055;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_231;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_233;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_235;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_237;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_239;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_241;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_243;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_245;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_247;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_249;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_251;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_253;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_255;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_257;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_259;
  wire \DLX_EXinst_Mshift__n0025_Sh[22] ;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_260;
  wire vga_top_vga1__n0013;
  wire vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_1;
  wire vga_top_vga1__n0012;
  wire vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_3;
  wire vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_5;
  wire vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_7;
  wire DLX_IDinst__n0420;
  wire DLX_IDinst_delay_slot;
  wire DLX_IDinst_slot_num_FFd3;
  wire DLX_IDinst_slot_num_FFd1;
  wire DLX_IDinst_slot_num_FFd2;
  wire N109741;
  wire DLX_IDinst_N70570;
  wire CHOICE2516;
  wire DLX_IDinst_Ker709161_1;
  wire DLX_IDinst__n03641_1;
  wire DLX_IDinst_N70918;
  wire reset_IBUF_4;
  wire DLX_IDinst_mem_to_reg;
  wire DLX_IDinst_mem_read;
  wire DLX_EXinst_mem_to_reg_EX;
  wire DLX_EXinst_mem_read_EX;
  wire vga_top_vga1__n0052;
  wire vga_top_vga1_clockcounter_FFd1;
  wire DLX_IDinst_N69711;
  wire CHOICE4311;
  wire CHOICE4343;
  wire DLX_EXinst_N63689;
  wire CHOICE3879;
  wire CHOICE3909;
  wire DLX_IDinst__n0315;
  wire CHOICE2398;
  wire DLX_IDinst_N70991;
  wire DLX_IDinst_N70006;
  wire DLX_IDinst__n0132;
  wire DLX_IDinst__n0338;
  wire DLX_IDinst__n0062;
  wire DLX_IDinst_N70658;
  wire DLX_IDinst__n0314;
  wire CHOICE2847;
  wire CHOICE1387;
  wire CHOICE1796;
  wire CHOICE1800;
  wire N100686;
  wire DLX_IDinst__n0440;
  wire DLX_IDinst_stall;
  wire N95693;
  wire DLX_IDinst_intr_slot;
  wire DLX_IFinst_IR_curr_N3638;
  wire DLX_IDinst_reg_write;
  wire DLX_IDinst_mem_write;
  wire DLX_EXinst_reg_write_EX;
  wire DLX_IDinst__n0085;
  wire DLX_EXinst_N66350;
  wire DLX_IDinst__n0105;
  wire DLX_IDinst__n0104;
  wire DLX_IDinst__n0103;
  wire DLX_IDinst__n0102;
  wire DLX_EXinst_N66078;
  wire CHOICE5522;
  wire CHOICE5567;
  wire N101921;
  wire N91278;
  wire DLX_EXinst_N66130;
  wire DLX_EXinst_word;
  wire DLX_EXinst_byte;
  wire DLX_IDinst__n0443;
  wire DLX_IDinst__n0331;
  wire DLX_IDinst__n0387;
  wire DLX_IDinst__n0071;
  wire DLX_IDinst__n0310;
  wire DLX_IFinst_PC_N3535;
  wire CHOICE3460;
  wire N102532;
  wire DLX_IDinst_N69568;
  wire DLX_IDinst__n0133;
  wire N90322;
  wire N100496;
  wire DLX_IDinst_N70673;
  wire DLX_IDinst_N70821;
  wire N100243;
  wire N127551;
  wire N110935;
  wire CHOICE3205;
  wire CHOICE3208;
  wire DLX_EXinst__n0049;
  wire CHOICE3210;
  wire N108909;
  wire N101161;
  wire CHOICE2458;
  wire DLX_IDinst_N69914;
  wire CHOICE2461;
  wire CHOICE2194;
  wire CHOICE2197;
  wire CHOICE2386;
  wire CHOICE2482;
  wire CHOICE2338;
  wire CHOICE2218;
  wire DLX_MEMlc_pd_wint1;
  wire DLX_MEMlc_md_wint1;
  wire DLX_MEMlc_ridp3;
  wire DLX_MEMlc_md_wint2;
  wire DLX_EXinst_N66535;
  wire CHOICE4276;
  wire \DLX_EXinst_Mshift__n0027_Sh[23] ;
  wire CHOICE5801;
  wire N127155;
  wire DLX_EXinst__n0077;
  wire N107780;
  wire N108266;
  wire N126593;
  wire N126451;
  wire CHOICE2485;
  wire DLX_EXinst_N63284;
  wire DLX_EXinst_N62946;
  wire \DLX_EXinst_Mshift__n0023_Sh[5] ;
  wire CHOICE4459;
  wire CHOICE2221;
  wire N127392;
  wire N127298;
  wire CHOICE2206;
  wire DLX_MEMlc_md_wint12;
  wire DLX_MEMlc_md_wint13;
  wire DLX_MEMlc_md_wint3;
  wire CHOICE2209;
  wire DLX_reqout_MEM;
  wire DLX_MEMlc_slave_ctrlMEM_l;
  wire DLX_MEMlc_master_ctrlMEM_nro;
  wire CHOICE39;
  wire CHOICE2422;
  wire CHOICE2230;
  wire DLX_MEMlc_md_wint11;
  wire DLX_MEMlc_md_wint4;
  wire DLX_EXinst_N66177;
  wire N108433;
  wire CHOICE5307;
  wire CHOICE5316;
  wire N95120;
  wire CHOICE5230;
  wire CHOICE5239;
  wire N126519;
  wire N126584;
  wire DLX_EXinst__n0030;
  wire CHOICE4944;
  wire CHOICE4973;
  wire CHOICE4941;
  wire N100490;
  wire CHOICE5011;
  wire N126461;
  wire DLX_reqout_ID;
  wire DLX_reqin_IF;
  wire CHOICE2233;
  wire CHOICE1090;
  wire CHOICE1096;
  wire N126297;
  wire N126393;
  wire DLX_IDinst_N70653;
  wire N90148;
  wire CHOICE2266;
  wire CHOICE2242;
  wire N127388;
  wire N127318;
  wire DLX_MEMlc_md_wint6;
  wire DLX_MEMlc_md_wint7;
  wire DLX_MEMlc_md_wint5;
  wire CHOICE2245;
  wire DLX_EXinst_N64062;
  wire CHOICE2997;
  wire N107613;
  wire CHOICE4087;
  wire CHOICE4088;
  wire CHOICE3493;
  wire CHOICE3494;
  wire CHOICE3499;
  wire CHOICE3500;
  wire N126293;
  wire DLX_EXinst_N62791;
  wire DLX_EXinst_N63454;
  wire DLX_reqout_EX;
  wire DLX_EXlc_slave_ctrlEX_l;
  wire CHOICE45;
  wire \DLX_EXinst_Mshift__n0025_Sh[15] ;
  wire \DLX_EXinst_Mshift__n0025_Sh[47] ;
  wire DLX_RF_delay_inst_wint9;
  wire DLX_RF_delay_inst_wint10;
  wire CHOICE3436;
  wire vga_top_vga1_N73394;
  wire vga_top_vga1_N73363;
  wire CHOICE3221;
  wire DLX_RF_delay_inst_wint11;
  wire N127098;
  wire DLX_RF_delay_inst_wint12;
  wire DLX_RF_delay_inst_wint19;
  wire DLX_RF_delay_inst_wint21;
  wire vga_top_vga1_N73379;
  wire vga_top_vga1_N73357;
  wire vga_top_vga1_N73389;
  wire DLX_RF_delay_inst_wint13;
  wire DM_delay_inst_wint1;
  wire vga_top_vga1_N73374;
  wire CHOICE3425;
  wire CHOICE3444;
  wire CHOICE3445;
  wire DLX_RF_delay_inst_wint15;
  wire DLX_RF_delay_inst_wint22;
  wire DLX_RF_delay_inst_wint29;
  wire DM_delay_inst_wint2;
  wire DLX_RF_delay_inst_wint23;
  wire DM_delay_inst_wint3;
  wire CHOICE3518;
  wire CHOICE3519;
  wire DLX_EXinst__n0114;
  wire N101725;
  wire CHOICE5746;
  wire CHOICE5850;
  wire DLX_RF_delay_inst_wint16;
  wire DLX_RF_delay_inst_wint25;
  wire DM_delay_inst_wint4;
  wire DLX_MEMlc_md_wint9;
  wire DLX_RF_delay_inst_wint17;
  wire DM_delay_inst_wint5;
  wire DLX_RF_delay_inst_wint18;
  wire DLX_RF_delay_inst_wint26;
  wire DM_delay_inst_wint6;
  wire DLX_IDinst_N70077;
  wire N126589;
  wire DLX_RF_delay_inst_wint27;
  wire DM_delay_inst_wint7;
  wire DLX_EXinst_N66525;
  wire \DLX_EXinst_Mshift__n0027_Sh[1] ;
  wire N109130;
  wire \DLX_EXinst_Mshift__n0028_Sh[49] ;
  wire DLX_EXinst_N66373;
  wire CHOICE5657;
  wire CHOICE5659;
  wire CHOICE2100;
  wire N95527;
  wire DLX_RF_delay_inst_wint28;
  wire DM_delay_inst_wint8;
  wire DLX_ackout_ID;
  wire DLX_IDlc_slave_ctrlID_l;
  wire DLX_IDlc_master_ctrlID_nro;
  wire CHOICE51;
  wire DM_delay_inst_wint9;
  wire DLX_EXinst_N66087;
  wire CHOICE5411;
  wire CHOICE5491;
  wire DLX_IDinst_N70610;
  wire DLX_IDinst__n0350;
  wire DLX_IDinst__n0348;
  wire N127139;
  wire CHOICE3523;
  wire DLX_IDinst_N70035;
  wire CHOICE3525;
  wire CHOICE3526;
  wire vga_top_vga1_N73399;
  wire CHOICE3224;
  wire \DLX_EXinst_Mshift__n0027_Sh[3] ;
  wire \DLX_EXinst_Mshift__n0028_Sh[51] ;
  wire CHOICE5020;
  wire CHOICE5022;
  wire N127378;
  wire N127370;
  wire DLX_IFlc_pd_wint1;
  wire DLX_IFlc_md_wint32;
  wire DLX_IFlc_md_wint9;
  wire DLX_IFlc_md_wint33;
  wire DLX_IFlc_md_wint10;
  wire DLX_IFlc_md_wint31;
  wire DLX_IFlc_md_wint11;
  wire CHOICE5169;
  wire DLX_EXinst__n0128;
  wire N126847;
  wire CHOICE5172;
  wire CHOICE3317;
  wire DLX_IFlc_md_wint28;
  wire DLX_IFlc_md_wint19;
  wire DLX_IFlc_md_wint29;
  wire DLX_IFlc_md_wint20;
  wire DLX_IFlc_md_wint27;
  wire DLX_IFlc_md_wint12;
  wire DLX_IDinst_N70924;
  wire N126580;
  wire CHOICE3470;
  wire N106726;
  wire N126776;
  wire CHOICE2849;
  wire \DLX_EXinst_Mshift__n0027_Sh[47] ;
  wire DLX_IDinst__n0250;
  wire CHOICE3480;
  wire DLX_EXinst_N63484;
  wire CHOICE3472;
  wire CHOICE3481;
  wire DLX_IFlc_md_wint24;
  wire DLX_IFlc_md_wint25;
  wire DLX_IFlc_md_wint21;
  wire DLX_IFlc_md_wint23;
  wire DLX_IFlc_md_wint13;
  wire CHOICE292;
  wire DLX_EXinst_N62806;
  wire DLX_EXinst_N63006;
  wire DLX_EXinst_N66226;
  wire CHOICE4396;
  wire DLX_IFlc_md_wint18;
  wire DLX_IFlc_md_wint22;
  wire DLX_IFlc_md_wint14;
  wire DLX_EXinst_N62811;
  wire DLX_EXinst_N66485;
  wire \DLX_EXinst_Mshift__n0028_Sh[22] ;
  wire \DLX_EXinst_Mshift__n0028_Sh[30] ;
  wire \DLX_EXinst_Mshift__n0024_Sh[26] ;
  wire DLX_EXinst_N63026;
  wire CHOICE3077;
  wire \DLX_EXinst_Mshift__n0028_Sh[52] ;
  wire CHOICE1324;
  wire DLX_EXinst_N63514;
  wire DLX_EXinst_N63011;
  wire N94007;
  wire CHOICE3246;
  wire CHOICE3249;
  wire N125959;
  wire DLX_MEMinst_noop;
  wire DLX_EXinst_noop;
  wire DLX_IFlc_md_wint17;
  wire DLX_IFlc_md_wint15;
  wire DLX_EXinst_N63790;
  wire N94205;
  wire \DLX_EXinst_Mshift__n0028_Sh[17] ;
  wire \DLX_EXinst_Mshift__n0024_Sh[25] ;
  wire DLX_EXinst_N64854;
  wire CHOICE3745;
  wire CHOICE3759;
  wire CHOICE3736;
  wire CHOICE3791;
  wire N126534;
  wire \DLX_EXinst_Mshift__n0028_Sh[19] ;
  wire DLX_EXinst_N64849;
  wire DLX_EXinst_N63414;
  wire DLX_IFlc_md_wint8;
  wire DLX_IFlc_md_wint16;
  wire DLX_IFlc_md_wint39;
  wire DLX_EXinst_N63424;
  wire DLX_EXinst_N63056;
  wire \DLX_EXinst_Mshift__n0025_Sh[7] ;
  wire \DLX_EXinst_Mshift__n0025_Sh[23] ;
  wire DLX_EXinst_N64104;
  wire DLX_EXinst_N63339;
  wire DLX_EXinst_N63304;
  wire CHOICE1030;
  wire \DLX_EXinst_Mshift__n0028_Sh[58] ;
  wire CHOICE3917;
  wire CHOICE4487;
  wire N127404;
  wire DLX_EXinst_N63051;
  wire DLX_EXinst_N62856;
  wire DLX_EXinst_N63404;
  wire N94057;
  wire N127322;
  wire N127374;
  wire DLX_IDinst__n0335;
  wire DLX_IDinst__n0442;
  wire N90101;
  wire N127126;
  wire N127189;
  wire N90255;
  wire DLX_IDinst_N70635;
  wire DLX_IDinst_N70885;
  wire N100191;
  wire DLX_IDinst_N70072;
  wire DM_delay_inst_wint10;
  wire DLX_IDinst__n0145;
  wire DLX_IDinst_N70716;
  wire DLX_IFlc_md_wint35;
  wire CHOICE3457;
  wire CHOICE2099;
  wire CHOICE3458;
  wire DM_delay_inst_wint11;
  wire N93955;
  wire \DLX_EXinst_Mshift__n0028_Sh[21] ;
  wire DLX_EXinst_N64560;
  wire DLX_EXinst_N64072;
  wire DM_delay_inst_wint12;
  wire DM_delay_inst_wint19;
  wire DM_delay_inst_wint21;
  wire DLX_EXlc_master_ctrlEX_nro;
  wire CHOICE3377;
  wire CHOICE3408;
  wire DLX_EXinst_N66507;
  wire N126811;
  wire \DLX_EXinst_Mshift__n0028_Sh[16] ;
  wire CHOICE1321;
  wire DLX_EXinst_N65105;
  wire DLX_EXinst_N63081;
  wire DLX_EXinst_N62951;
  wire CHOICE4164;
  wire DM_delay_inst_wint13;
  wire DLX_EXinst_N63434;
  wire DLX_EXinst_N64314;
  wire CHOICE4628;
  wire DM_delay_inst_wint14;
  wire DM_delay_inst_wint22;
  wire DM_delay_inst_wint29;
  wire DM_delay_inst_wint30;
  wire DLX_EXinst_N63712;
  wire CHOICE5244;
  wire CHOICE5247;
  wire CHOICE5204;
  wire N126576;
  wire CHOICE5333;
  wire CHOICE4098;
  wire DM_delay_inst_wint15;
  wire DM_delay_inst_wint23;
  wire DM_delay_inst_wint31;
  wire DLX_EXinst_N62976;
  wire DLX_EXinst_N62866;
  wire DLX_EXinst_N63364;
  wire \DLX_EXinst_Mshift__n0026_Sh[19] ;
  wire DLX_EXinst_N64324;
  wire CHOICE4842;
  wire N127396;
  wire DLX_EXinst_N63444;
  wire DLX_IFlc_master_ctrlIF_l;
  wire DLX_RF_delay_inst_wint3;
  wire DM_delay_inst_wint16;
  wire DM_delay_inst_wint24;
  wire DM_delay_inst_wint32;
  wire DM_delay_inst_wint39;
  wire DLX_EXinst_N62733;
  wire CHOICE2085;
  wire \DLX_EXinst_Mshift__n0028_Sh[29] ;
  wire DLX_EXinst_N63269;
  wire CHOICE1758;
  wire DLX_EXinst_N63001;
  wire DLX_EXinst_N63509;
  wire N126263;
  wire CHOICE5740;
  wire CHOICE4610;
  wire CHOICE4032;
  wire DM_delay_inst_wint17;
  wire DM_delay_inst_wint25;
  wire DM_delay_inst_wint33;
  wire N95569;
  wire \DLX_EXinst_Mshift__n0028_Sh[24] ;
  wire CHOICE1132;
  wire DLX_EXinst_N63294;
  wire CHOICE1356;
  wire CHOICE1138;
  wire CHOICE1144;
  wire DLX_EXinst_N64530;
  wire CHOICE4261;
  wire CHOICE1282;
  wire \DLX_EXinst_Mshift__n0025_Sh[21] ;
  wire DLX_EXinst_N64094;
  wire CHOICE4780;
  wire N127314;
  wire N127286;
  wire DM_delay_inst_wint18;
  wire DM_delay_inst_wint27;
  wire DM_delay_inst_wint35;
  wire DLX_EXinst_N64864;
  wire N126134;
  wire \DLX_EXinst_Mshift__n0023_Sh[8] ;
  wire CHOICE5864;
  wire DLX_IFlc_md_wint7;
  wire DLX_IFlc_ridp3;
  wire DLX_IFlc_md_wint1;
  wire DLX_EXinst_N64804;
  wire CHOICE4016;
  wire DLX_EXinst_N62861;
  wire DLX_EXinst_N63359;
  wire DLX_EXinst_N63474;
  wire DLX_EXinst_N63519;
  wire \DLX_EXinst_Mshift__n0026_Sh[16] ;
  wire CHOICE3889;
  wire DLX_EXinst_N62776;
  wire DLX_EXinst_N63439;
  wire N95202;
  wire N57312;
  wire DLX_IFlc_md_wint6;
  wire DLX_IFlc_md_wint36;
  wire DLX_EXinst_N66112;
  wire DLX_EXinst_N62886;
  wire DLX_EXinst_N63384;
  wire DLX_EXinst_N62801;
  wire DLX_EXinst_N63464;
  wire \DLX_EXinst_Mshift__n0027_Sh[21] ;
  wire DM_delay_inst_wint28;
  wire DM_delay_inst_wint36;
  wire vga_top_vga1_videoon;
  wire DLX_EXinst_N63369;
  wire DLX_EXinst_N66105;
  wire DLX_EXinst_N62786;
  wire DLX_EXinst_N63449;
  wire DLX_EXinst_N64545;
  wire DLX_EXinst_N64329;
  wire CHOICE4321;
  wire CHOICE5408;
  wire CHOICE4740;
  wire CHOICE4675;
  wire CHOICE5574;
  wire DM_delay_inst_wint37;
  wire \DLX_EXinst_Mshift__n0027_Sh[0] ;
  wire CHOICE5976;
  wire DM_delay_inst_wint38;
  wire DLX_IFlc_md_wint5;
  wire DLX_IFlc_md_wint2;
  wire \DLX_EXinst_Mshift__n0025_Sh[19] ;
  wire CHOICE3836;
  wire DLX_EXinst_N64099;
  wire CHOICE3818;
  wire CHOICE5663;
  wire DLX_IFlc_md_wint4;
  wire DLX_IFlc_md_wint37;
  wire CHOICE859;
  wire \DLX_EXinst_Mshift__n0028_Sh[50] ;
  wire CHOICE3692;
  wire CHOICE5493;
  wire CHOICE1018;
  wire CHOICE1024;
  wire CHOICE4432;
  wire CHOICE1294;
  wire DLX_EXinst_N63469;
  wire DLX_EXinst_N63389;
  wire CHOICE5256;
  wire \DLX_EXinst_Mshift__n0028_Sh[11] ;
  wire DLX_IFlc_md_wint38;
  wire DLX_IFlc_md_wint3;
  wire DLX_EXinst_N64587;
  wire CHOICE4438;
  wire CHOICE5497;
  wire N93905;
  wire \DLX_EXinst_Mshift__n0024_Sh[29] ;
  wire DLX_EXinst_N64550;
  wire \DLX_EXinst_Mshift__n0026_Sh[30] ;
  wire N94255;
  wire DLX_EXinst_N65160;
  wire \DLX_EXinst_Mshift__n0023_Sh[29] ;
  wire \DLX_EXinst_Mshift__n0028_Sh[9] ;
  wire N93435;
  wire DLX_EXinst__n0147;
  wire DLX_IDinst_Mmux__n0148__net123;
  wire DLX_EXinst_N63785;
  wire DLX_EXinst_N62771;
  wire DLX_EXinst_N62991;
  wire CHOICE4554;
  wire CHOICE5026;
  wire N97593;
  wire DLX_EXinst_N66152;
  wire CHOICE3978;
  wire CHOICE3980;
  wire vga_top_vga1_helpme;
  wire N100333;
  wire \DLX_EXinst_Mshift__n0027_Sh[20] ;
  wire CHOICE1364;
  wire DLX_EXinst_N65100;
  wire N101839;
  wire CHOICE4567;
  wire DLX_EXinst_N66060;
  wire DLX_EXinst_N63836;
  wire DLX_IDinst__n0147;
  wire \DLX_EXinst_Mshift__n0025_Sh[12] ;
  wire N127334;
  wire DLX_EXinst_N62781;
  wire \DLX_EXinst_Mshift__n0025_Sh[20] ;
  wire DLX_EXinst_N63925;
  wire N97233;
  wire CHOICE3869;
  wire \DLX_EXinst_Mshift__n0025_Sh[3] ;
  wire \DLX_EXinst_Mshift__n0028_Sh[10] ;
  wire \DLX_EXinst_Mshift__n0028_Sh[18] ;
  wire DLX_EXinst_N64067;
  wire DLX_EXinst_N64814;
  wire CHOICE5384;
  wire CHOICE5393;
  wire N126442;
  wire N127107;
  wire CHOICE1343;
  wire CHOICE5577;
  wire DLX_EXinst_N66096;
  wire CHOICE1359;
  wire DLX_EXinst_N64824;
  wire DLX_EXinst_N63915;
  wire CHOICE4504;
  wire CHOICE4422;
  wire \DLX_EXinst_Mshift__n0027_Sh[22] ;
  wire \DLX_EXinst_Mshift__n0025_Sh[0] ;
  wire CHOICE3990;
  wire CHOICE3992;
  wire CHOICE3994;
  wire N127306;
  wire CHOICE1066;
  wire CHOICE3666;
  wire CHOICE3673;
  wire CHOICE3642;
  wire CHOICE3651;
  wire CHOICE3658;
  wire CHOICE3674;
  wire N126289;
  wire DLX_EXinst_N66519;
  wire DLX_EXinst_N66072;
  wire N95300;
  wire \DLX_EXinst_Mshift__n0023_Sh[30] ;
  wire \DLX_EXinst_Mshift__n0023_Sh[26] ;
  wire N89980;
  wire DLX_EXinst_N66443;
  wire \DLX_EXinst_Mshift__n0025_Sh[4] ;
  wire N96585;
  wire CHOICE4429;
  wire CHOICE4439;
  wire CHOICE4175;
  wire CHOICE4189;
  wire CHOICE4223;
  wire N126415;
  wire CHOICE3620;
  wire CHOICE3627;
  wire CHOICE3635;
  wire DLX_IDinst_zflag;
  wire CHOICE3267;
  wire DLX_EXinst__n0082;
  wire DLX_EXinst_N63031;
  wire \DLX_EXinst_Mshift__n0024_Sh[127] ;
  wire CHOICE4806;
  wire DLX_EXinst_N66437;
  wire N126528;
  wire CHOICE3802;
  wire CHOICE4354;
  wire N90461;
  wire \DLX_EXinst_Mshift__n0025_Sh[1] ;
  wire CHOICE1072;
  wire N90557;
  wire \DLX_EXinst_Mshift__n0025_Sh[2] ;
  wire CHOICE5556;
  wire CHOICE5223;
  wire DLX_EXinst_N66383;
  wire DLX_EXinst__n0061;
  wire CHOICE5905;
  wire CHOICE3812;
  wire CHOICE4364;
  wire CHOICE4361;
  wire CHOICE4370;
  wire CHOICE4371;
  wire CHOICE4792;
  wire N126281;
  wire CHOICE4796;
  wire DLX_EXinst_N66392;
  wire CHOICE5377;
  wire CHOICE1300;
  wire CHOICE3610;
  wire CHOICE3534;
  wire CHOICE4492;
  wire \DLX_EXinst_Mshift__n0024_Sh[28] ;
  wire CHOICE2075;
  wire DLX_EXinst_N66475;
  wire N96513;
  wire CHOICE3809;
  wire CHOICE3819;
  wire CHOICE4599;
  wire CHOICE5229;
  wire N127302;
  wire CHOICE4119;
  wire CHOICE3684;
  wire N127412;
  wire CHOICE3540;
  wire CHOICE3556;
  wire N90344;
  wire DLX_IDinst_N70295;
  wire N127093;
  wire CHOICE3691;
  wire CHOICE3698;
  wire CHOICE3699;
  wire DLX_IDinst_N70786;
  wire CHOICE2558;
  wire CHOICE2679;
  wire CHOICE3603;
  wire CHOICE4560;
  wire CHOICE4566;
  wire CHOICE4569;
  wire CHOICE3876;
  wire CHOICE2523;
  wire CHOICE2525;
  wire CHOICE5107;
  wire CHOICE5128;
  wire CHOICE5129;
  wire CHOICE2635;
  wire CHOICE2690;
  wire CHOICE2877;
  wire CHOICE2778;
  wire N100440;
  wire DLX_IDinst_N70623;
  wire N126038;
  wire CHOICE283;
  wire CHOICE5181;
  wire CHOICE2712;
  wire CHOICE2800;
  wire CHOICE2756;
  wire CHOICE2701;
  wire N95654;
  wire N95611;
  wire CHOICE4954;
  wire CHOICE2811;
  wire CHOICE2822;
  wire CHOICE2657;
  wire CHOICE2789;
  wire CHOICE4507;
  wire CHOICE4549;
  wire CHOICE4508;
  wire CHOICE4570;
  wire CHOICE2569;
  wire CHOICE2723;
  wire CHOICE2562;
  wire N100609;
  wire CHOICE2563;
  wire CHOICE2591;
  wire CHOICE2833;
  wire CHOICE2888;
  wire CHOICE2734;
  wire CHOICE5606;
  wire CHOICE5648;
  wire N126601;
  wire CHOICE4741;
  wire CHOICE4766;
  wire CHOICE4798;
  wire N126276;
  wire CHOICE2580;
  wire CHOICE2745;
  wire CHOICE2899;
  wire CHOICE2855;
  wire CHOICE3412;
  wire CHOICE2584;
  wire CHOICE2585;
  wire CHOICE2602;
  wire CHOICE2767;
  wire vga_top_vga1_clockcounter_FFd2;
  wire CHOICE2613;
  wire CHOICE2866;
  wire N125999;
  wire CHOICE2573;
  wire CHOICE2574;
  wire CHOICE1410;
  wire CHOICE1411;
  wire N98127;
  wire N108101;
  wire N126597;
  wire N126524;
  wire CHOICE2881;
  wire CHOICE2595;
  wire DLX_IDinst_N70663;
  wire N98806;
  wire DLX_IDinst_CLI;
  wire DLX_IDinst_N70333;
  wire CHOICE2596;
  wire DLX_IDinst_N70328;
  wire N127435;
  wire CHOICE2606;
  wire CHOICE2607;
  wire DLX_IDinst__n0151;
  wire N100688;
  wire CHOICE2617;
  wire CHOICE2618;
  wire DLX_IDinst__n0070;
  wire CHOICE2639;
  wire CHOICE2640;
  wire CHOICE2627;
  wire N127423;
  wire DLX_IDinst__n0252;
  wire N127366;
  wire N127294;
  wire N127362;
  wire N127290;
  wire N90497;
  wire CHOICE1479;
  wire CHOICE1757;
  wire DLX_IDinst__n0144;
  wire N95818;
  wire CHOICE2650;
  wire CHOICE2646;
  wire CHOICE2651;
  wire CHOICE4498;
  wire CHOICE4505;
  wire CHOICE4248;
  wire CHOICE3922;
  wire CHOICE2661;
  wire CHOICE2662;
  wire CHOICE3928;
  wire CHOICE3934;
  wire CHOICE3935;
  wire CHOICE3937;
  wire \DLX_EXinst_Mshift__n0023_Sh[127] ;
  wire CHOICE4849;
  wire CHOICE5047;
  wire CHOICE4185;
  wire CHOICE3861;
  wire N90656;
  wire N126506;
  wire CHOICE2508;
  wire CHOICE2668;
  wire CHOICE1444;
  wire CHOICE4879;
  wire N102270;
  wire CHOICE2081;
  wire CHOICE4234;
  wire CHOICE3862;
  wire CHOICE4206;
  wire CHOICE4220;
  wire CHOICE4196;
  wire CHOICE4211;
  wire N126419;
  wire CHOICE4621;
  wire DLX_EXinst__n0063;
  wire CHOICE5899;
  wire CHOICE4018;
  wire CHOICE4000;
  wire CHOICE4004;
  wire CHOICE4021;
  wire N126239;
  wire CHOICE4023;
  wire CHOICE4878;
  wire N97892;
  wire CHOICE4611;
  wire CHOICE4882;
  wire N127354;
  wire N127400;
  wire CHOICE3870;
  wire CHOICE3877;
  wire CHOICE4676;
  wire CHOICE3938;
  wire N127358;
  wire N127326;
  wire CHOICE3755;
  wire CHOICE4293;
  wire CHOICE3297;
  wire N127182;
  wire CHOICE4242;
  wire CHOICE4302;
  wire N100282;
  wire \DLX_EXinst_Mshift__n0027_Sh[41] ;
  wire N102162;
  wire CHOICE4294;
  wire CHOICE4897;
  wire CHOICE4884;
  wire N127200;
  wire DLX_EXinst_N64304;
  wire CHOICE4173;
  wire DLX_EXinst_N64859;
  wire CHOICE4241;
  wire CHOICE4301;
  wire N127350;
  wire CHOICE5421;
  wire CHOICE4233;
  wire CHOICE4308;
  wire CHOICE4309;
  wire N127342;
  wire N127338;
  wire CHOICE4686;
  wire CHOICE4895;
  wire CHOICE4811;
  wire DLX_EXinst_N64309;
  wire CHOICE4107;
  wire CHOICE4109;
  wire CHOICE4249;
  wire CHOICE4251;
  wire CHOICE19;
  wire DLX_EXlc_md_wint32;
  wire DLX_EXlc_pd_wint5;
  wire DLX_EXlc_ridp3;
  wire DLX_EXlc_md_wint33;
  wire DLX_EXlc_md_wint1;
  wire CHOICE5753;
  wire CHOICE5754;
  wire CHOICE4817;
  wire CHOICE4823;
  wire CHOICE4828;
  wire CHOICE4830;
  wire CHOICE3353;
  wire N126482;
  wire CHOICE5617;
  wire CHOICE5891;
  wire CHOICE4041;
  wire CHOICE4043;
  wire N126054;
  wire CHOICE3274;
  wire CHOICE2548;
  wire CHOICE5764;
  wire DLX_EXinst_N64077;
  wire CHOICE3743;
  wire DLX_EXlc_md_wint2;
  wire CHOICE5875;
  wire CHOICE5877;
  wire CHOICE5276;
  wire CHOICE5278;
  wire CHOICE1991;
  wire N102453;
  wire CHOICE5915;
  wire CHOICE5917;
  wire N127252;
  wire CHOICE3068;
  wire CHOICE1861;
  wire N127346;
  wire CHOICE5046;
  wire N127330;
  wire CHOICE4751;
  wire CHOICE2060;
  wire CHOICE1951;
  wire CHOICE5587;
  wire CHOICE4053;
  wire DLX_MEMlc_md_wint19;
  wire CHOICE4980;
  wire CHOICE5883;
  wire DLX_EXinst_N62941;
  wire CHOICE1868;
  wire N101095;
  wire DLX_EXlc_md_wint31;
  wire DLX_EXlc_md_wint3;
  wire N127310;
  wire CHOICE5953;
  wire CHOICE5954;
  wire \DLX_EXinst_Mshift__n0024_Sh[30] ;
  wire CHOICE1904;
  wire CHOICE1911;
  wire CHOICE1957;
  wire CHOICE5684;
  wire CHOICE5704;
  wire CHOICE4123;
  wire \DLX_EXinst_Mshift__n0028_Sh[57] ;
  wire CHOICE4758;
  wire N126306;
  wire N126107;
  wire CHOICE5914;
  wire CHOICE5517;
  wire CHOICE5683;
  wire CHOICE1962;
  wire N101641;
  wire CHOICE2046;
  wire \DLX_EXinst_Mshift__n0023_Sh[25] ;
  wire DLX_EXlc_md_wint28;
  wire DLX_EXlc_md_wint29;
  wire DLX_EXlc_md_wint4;
  wire N94107;
  wire CHOICE1150;
  wire CHOICE1156;
  wire DLX_EXinst_N63299;
  wire N126571;
  wire CHOICE5686;
  wire CHOICE5688;
  wire N126092;
  wire CHOICE5928;
  wire CHOICE5934;
  wire CHOICE5943;
  wire CHOICE5944;
  wire CHOICE1985;
  wire \DLX_EXinst_Mshift__n0026_Sh[49] ;
  wire CHOICE5722;
  wire CHOICE5724;
  wire CHOICE5728;
  wire CHOICE5729;
  wire CHOICE1036;
  wire CHOICE4693;
  wire N126383;
  wire CHOICE4763;
  wire N126301;
  wire \DLX_EXinst_Mshift__n0026_Sh[50] ;
  wire N126370;
  wire CHOICE5716;
  wire CHOICE5730;
  wire N127163;
  wire N101338;
  wire CHOICE1972;
  wire CHOICE5714;
  wire CHOICE4520;
  wire DLX_EXlc_md_wint27;
  wire DLX_EXlc_md_wint5;
  wire CHOICE5518;
  wire N98808;
  wire CHOICE5983;
  wire N126252;
  wire CHOICE5991;
  wire CHOICE5921;
  wire CHOICE3058;
  wire CHOICE5982;
  wire CHOICE5733;
  wire CHOICE4453;
  wire CHOICE4698;
  wire N126375;
  wire N110183;
  wire N127223;
  wire CHOICE1379;
  wire N98218;
  wire CHOICE2069;
  wire CHOICE3060;
  wire DLX_EXlc_md_wint24;
  wire DLX_EXlc_md_wint25;
  wire DLX_EXlc_md_wint6;
  wire CHOICE5530;
  wire CHOICE5542;
  wire CHOICE5543;
  wire CHOICE4130;
  wire CHOICE5562;
  wire CHOICE4385;
  wire CHOICE5520;
  wire \DLX_EXinst_Mshift__n0024_Sh[80] ;
  wire CHOICE5988;
  wire CHOICE5558;
  wire CHOICE5563;
  wire CHOICE3069;
  wire N126469;
  wire DLX_EXlc_md_wint23;
  wire DLX_EXlc_md_wint7;
  wire \DLX_EXinst_Mshift__n0026_Sh[6] ;
  wire CHOICE4391;
  wire CHOICE5550;
  wire CHOICE4537;
  wire CHOICE5564;
  wire CHOICE5548;
  wire CHOICE5300;
  wire CHOICE1349;
  wire CHOICE1102;
  wire CHOICE1331;
  wire DLX_EXinst_N63071;
  wire DLX_EXlc_md_wint22;
  wire DLX_EXlc_md_wint8;
  wire CHOICE5201;
  wire CHOICE5203;
  wire CHOICE5049;
  wire CHOICE5051;
  wire CHOICE2971;
  wire CHOICE5080;
  wire CHOICE5085;
  wire CHOICE5058;
  wire CHOICE5062;
  wire CHOICE5086;
  wire CHOICE5088;
  wire CHOICE3283;
  wire CHOICE1337;
  wire N107444;
  wire N90062;
  wire CHOICE1174;
  wire DLX_EXlc_md_wint21;
  wire DLX_EXlc_md_wint9;
  wire CHOICE5353;
  wire CHOICE5355;
  wire CHOICE5089;
  wire CHOICE3214;
  wire CHOICE5056;
  wire CHOICE3275;
  wire N109350;
  wire \DLX_EXinst_Mshift__n0026_Sh[52] ;
  wire CHOICE4003;
  wire DLX_EXinst_N63021;
  wire CHOICE3104;
  wire CHOICE1180;
  wire N94921;
  wire CHOICE4464;
  wire CHOICE3844;
  wire CHOICE5613;
  wire CHOICE1288;
  wire N126424;
  wire CHOICE3564;
  wire CHOICE4025;
  wire CHOICE4017;
  wire CHOICE5236;
  wire CHOICE3572;
  wire CHOICE3415;
  wire CHOICE3416;
  wire CHOICE4064;
  wire CHOICE3579;
  wire CHOICE4446;
  wire CHOICE4448;
  wire CHOICE3547;
  wire CHOICE3588;
  wire CHOICE4465;
  wire CHOICE4475;
  wire N126556;
  wire CHOICE4440;
  wire CHOICE4479;
  wire CHOICE4481;
  wire CHOICE3551;
  wire CHOICE3595;
  wire CHOICE3024;
  wire DLX_IDinst_N69781;
  wire CHOICE4596;
  wire CHOICE4472;
  wire CHOICE1210;
  wire CHOICE1108;
  wire CHOICE2008;
  wire N94857;
  wire CHOICE4378;
  wire CHOICE4380;
  wire CHOICE4478;
  wire CHOICE4397;
  wire CHOICE1417;
  wire CHOICE1418;
  wire N126610;
  wire CHOICE1216;
  wire CHOICE4157;
  wire N126478;
  wire CHOICE4372;
  wire CHOICE4411;
  wire CHOICE4413;
  wire CHOICE4407;
  wire N126614;
  wire CHOICE5383;
  wire CHOICE4404;
  wire DLX_EXlc_md_wint20;
  wire DLX_EXlc_md_wint10;
  wire N101425;
  wire CHOICE4410;
  wire CHOICE3826;
  wire CHOICE3828;
  wire CHOICE3833;
  wire CHOICE3847;
  wire N126465;
  wire CHOICE3166;
  wire CHOICE3168;
  wire CHOICE2043;
  wire CHOICE2051;
  wire CHOICE5356;
  wire CHOICE1452;
  wire CHOICE1453;
  wire CHOICE12;
  wire DLX_EXlc_md_wint19;
  wire DLX_EXlc_md_wint11;
  wire N101919;
  wire CHOICE3700;
  wire CHOICE3539;
  wire N126546;
  wire N126354;
  wire N96945;
  wire CHOICE3957;
  wire CHOICE2077;
  wire CHOICE3850;
  wire CHOICE3851;
  wire DLX_EXlc_md_wint18;
  wire DLX_EXlc_md_wint12;
  wire N102358;
  wire CHOICE3706;
  wire CHOICE3708;
  wire CHOICE3820;
  wire CHOICE3853;
  wire CHOICE3399;
  wire CHOICE3554;
  wire N126510;
  wire DLX_EXlc_md_wint17;
  wire DLX_EXlc_md_wint13;
  wire CHOICE3717;
  wire CHOICE3726;
  wire CHOICE3728;
  wire CHOICE3729;
  wire CHOICE3713;
  wire CHOICE3722;
  wire DLX_EXlc_md_wint16;
  wire DLX_EXlc_md_wint14;
  wire CHOICE2672;
  wire CHOICE2673;
  wire CHOICE2064;
  wire CHOICE5279;
  wire CHOICE1977;
  wire CHOICE4862;
  wire CHOICE4863;
  wire CHOICE3731;
  wire CHOICE3725;
  wire CHOICE1976;
  wire CHOICE2815;
  wire CHOICE2683;
  wire CHOICE4576;
  wire CHOICE4578;
  wire DLX_IFlc_master_ctrlIF_nro;
  wire DLX_IFlc_slave_ctrlIF_l;
  wire DLX_reqout_IF;
  wire CHOICE25;
  wire CHOICE3491;
  wire CHOICE2684;
  wire DLX_EXlc_md_wint35;
  wire DLX_EXlc_md_wint36;
  wire DLX_EXlc_md_wint15;
  wire CHOICE5126;
  wire N127149;
  wire \DLX_EXinst_Mshift__n0025_Sh[41] ;
  wire CHOICE4588;
  wire N126457;
  wire CHOICE5440;
  wire CHOICE5482;
  wire N126358;
  wire CHOICE4701;
  wire CHOICE4733;
  wire N126349;
  wire CHOICE3295;
  wire DLX_RF_delay_inst_wint4;
  wire CHOICE2551;
  wire N105035;
  wire DLX_RF_delay_inst_wint5;
  wire CHOICE4602;
  wire CHOICE4603;
  wire CHOICE2694;
  wire CHOICE2695;
  wire DLX_EXlc_md_wint37;
  wire CHOICE2782;
  wire CHOICE2783;
  wire CHOICE4605;
  wire DLX_RF_delay_inst_wint6;
  wire DLX_RF_delay_inst_wint7;
  wire DLX_RF_delay_inst_wint8;
  wire CHOICE2804;
  wire CHOICE2805;
  wire CHOICE2705;
  wire CHOICE2706;
  wire DLX_IDlc_md_wint32;
  wire DLX_IDlc_pd_wint1;
  wire DLX_IDlc_md_wint33;
  wire DLX_IDlc_ridp3;
  wire CHOICE1436;
  wire N95411;
  wire DLX_IDinst__n0173;
  wire CHOICE2760;
  wire CHOICE2793;
  wire N127196;
  wire N126388;
  wire CHOICE2716;
  wire CHOICE2717;
  wire CHOICE2826;
  wire CHOICE2827;
  wire CHOICE2794;
  wire CHOICE2913;
  wire CHOICE2182;
  wire CHOICE2727;
  wire CHOICE3466;
  wire DLX_IFlc_ridp2;
  wire CHOICE2816;
  wire CHOICE2728;
  wire CHOICE2093;
  wire CHOICE3448;
  wire CHOICE2738;
  wire CHOICE2739;
  wire CHOICE2837;
  wire CHOICE2838;
  wire CHOICE1786;
  wire DLX_EXlc_pd_wint1;
  wire DLX_EXlc_pd_wint2;
  wire N127555;
  wire DLX_EXlc_pd_wint3;
  wire DLX_EXlc_pd_wint4;
  wire DLX_EXlc_md_wint39;
  wire CHOICE2749;
  wire CHOICE2750;
  wire CHOICE2859;
  wire CHOICE2860;
  wire N92607;
  wire CHOICE2870;
  wire CHOICE2871;
  wire CHOICE2771;
  wire CHOICE2772;
  wire CHOICE5;
  wire DLX_EXlc_md_wint38;
  wire N95259;
  wire DLX_EXinst_N63996;
  wire DLX_EXinst_N64181;
  wire CHOICE5401;
  wire CHOICE2882;
  wire CHOICE2761;
  wire CHOICE5390;
  wire CHOICE4633;
  wire N126428;
  wire CHOICE4636;
  wire CHOICE1790;
  wire CHOICE2892;
  wire CHOICE2893;
  wire DLX_EXinst_N63910;
  wire CHOICE4283;
  wire CHOICE5398;
  wire N126437;
  wire CHOICE2903;
  wire CHOICE2904;
  wire DLX_EXinst_N64919;
  wire CHOICE4140;
  wire CHOICE4154;
  wire CHOICE4145;
  wire N126490;
  wire N92503;
  wire DLX_IDlc_md_wint31;
  wire DLX_IDlc_md_wint9;
  wire DLX_IDlc_md_wint10;
  wire DLX_IDlc_md_wint28;
  wire DLX_IDlc_md_wint29;
  wire DLX_IDlc_md_wint11;
  wire CHOICE4217;
  wire N126257;
  wire N92087;
  wire N92555;
  wire DLX_IDlc_md_wint27;
  wire DLX_IDlc_md_wint19;
  wire DLX_IDlc_md_wint20;
  wire DLX_IDlc_md_wint24;
  wire DLX_IDlc_md_wint25;
  wire DLX_IDlc_md_wint12;
  wire N91463;
  wire DLX_IDlc_md_wint23;
  wire DLX_IDlc_md_wint21;
  wire DLX_IDlc_md_wint22;
  wire DLX_IDlc_md_wint13;
  wire N126048;
  wire DLX_IDlc_md_wint18;
  wire DLX_IDlc_md_wint17;
  wire DLX_IDlc_md_wint14;
  wire CHOICE32;
  wire CHOICE3328;
  wire CHOICE3329;
  wire N95327;
  wire DLX_IDlc_md_wint16;
  wire DLX_IDlc_md_wint15;
  wire N92451;
  wire N91983;
  wire CHOICE3343;
  wire DLX_IDlc_md_wint8;
  wire N93075;
  wire CHOICE4514;
  wire CHOICE4516;
  wire DLX_IDlc_md_wint35;
  wire CHOICE4538;
  wire CHOICE4540;
  wire CHOICE4541;
  wire \DLX_EXinst_Mshift__n0025_Sh[42] ;
  wire CHOICE4532;
  wire N126564;
  wire CHOICE4970;
  wire CHOICE4543;
  wire CHOICE3944;
  wire CHOICE3946;
  wire N91619;
  wire N92399;
  wire N92035;
  wire CHOICE3950;
  wire CHOICE3964;
  wire CHOICE3966;
  wire CHOICE3967;
  wire N126807;
  wire DLX_EXinst__n0093;
  wire CHOICE4643;
  wire DLX_IDlc_md_wint7;
  wire DLX_IDlc_md_wint36;
  wire CHOICE5451;
  wire CHOICE3958;
  wire CHOICE3969;
  wire N93023;
  wire CHOICE3963;
  wire DLX_IDlc_md_wint6;
  wire DLX_IDlc_md_wint37;
  wire CHOICE5321;
  wire CHOICE5324;
  wire N126514;
  wire CHOICE4934;
  wire CHOICE4935;
  wire CHOICE5447;
  wire CHOICE3884;
  wire CHOICE2521;
  wire CHOICE4926;
  wire CHOICE4928;
  wire CHOICE4930;
  wire CHOICE3906;
  wire CHOICE3908;
  wire CHOICE1120;
  wire CHOICE4925;
  wire DLX_IDlc_md_wint5;
  wire DLX_IDlc_md_wint38;
  wire CHOICE4909;
  wire CHOICE4057;
  wire CHOICE3895;
  wire CHOICE3897;
  wire CHOICE3905;
  wire CHOICE4256;
  wire CHOICE4904;
  wire \DLX_EXinst_Mshift__n0025_Sh[44] ;
  wire CHOICE3903;
  wire CHOICE4913;
  wire CHOICE4915;
  wire CHOICE4329;
  wire CHOICE4339;
  wire CHOICE4340;
  wire DLX_IDlc_md_wint4;
  wire DLX_IDlc_md_wint39;
  wire CHOICE4091;
  wire N126538;
  wire CHOICE4999;
  wire N92347;
  wire N91515;
  wire N91931;
  wire CHOICE4219;
  wire CHOICE4708;
  wire CHOICE4316;
  wire CHOICE4342;
  wire CHOICE4205;
  wire CHOICE4336;
  wire CHOICE4337;
  wire CHOICE4327;
  wire CHOICE4269;
  wire CHOICE4279;
  wire CHOICE4280;
  wire N92971;
  wire CHOICE4153;
  wire N126411;
  wire CHOICE4151;
  wire CHOICE2509;
  wire N127567;
  wire CHOICE4282;
  wire CHOICE4139;
  wire CHOICE4277;
  wire CHOICE4267;
  wire CHOICE4831;
  wire CHOICE5784;
  wire CHOICE5315;
  wire CHOICE4860;
  wire CHOICE5147;
  wire CHOICE5168;
  wire CHOICE4079;
  wire CHOICE4085;
  wire N91879;
  wire N92243;
  wire CHOICE5326;
  wire N127563;
  wire CHOICE3766;
  wire CHOICE4837;
  wire CHOICE4865;
  wire CHOICE4866;
  wire CHOICE4073;
  wire CHOICE4074;
  wire N126398;
  wire CHOICE5828;
  wire CHOICE5785;
  wire N126495;
  wire N92919;
  wire CHOICE4668;
  wire N126403;
  wire CHOICE4868;
  wire CHOICE5818;
  wire N126446;
  wire CHOICE5845;
  wire CHOICE5788;
  wire N126362;
  wire CHOICE3785;
  wire CHOICE3775;
  wire CHOICE3789;
  wire CHOICE5145;
  wire DLX_reqin_ID;
  wire CHOICE5824;
  wire CHOICE3427;
  wire N126344;
  wire CHOICE3773;
  wire N126631;
  wire CHOICE5603;
  wire N126627;
  wire N92295;
  wire N90373;
  wire CHOICE5642;
  wire N126606;
  wire N91827;
  wire CHOICE3783;
  wire CHOICE5173;
  wire CHOICE4790;
  wire CHOICE5625;
  wire CHOICE5627;
  wire N126029;
  wire CHOICE4773;
  wire CHOICE5646;
  wire N92815;
  wire CHOICE4782;
  wire CHOICE2937;
  wire CHOICE2941;
  wire N126407;
  wire CHOICE5437;
  wire CHOICE5476;
  wire N126366;
  wire CHOICE4725;
  wire CHOICE4727;
  wire CHOICE4717;
  wire CHOICE4731;
  wire DLX_MEMlc_md_wint15;
  wire CHOICE5459;
  wire CHOICE5461;
  wire CHOICE4715;
  wire CHOICE5480;
  wire N107291;
  wire N126542;
  wire DLX_EXinst__n0095;
  wire N91723;
  wire N126432;
  wire N92191;
  wire CHOICE4660;
  wire CHOICE4662;
  wire CHOICE4652;
  wire CHOICE4666;
  wire DLX_MEMlc_md_wint17;
  wire DLX_MEMlc_md_wint18;
  wire DLX_MEMlc_md_wint16;
  wire CHOICE4650;
  wire CHOICE5008;
  wire N92867;
  wire N127167;
  wire CHOICE2927;
  wire N126820;
  wire CHOICE5238;
  wire CHOICE5249;
  wire N126551;
  wire N92139;
  wire N91775;
  wire CHOICE1114;
  wire N92763;
  wire N94733;
  wire CHOICE5392;
  wire CHOICE5403;
  wire N126207;
  wire N126379;
  wire N91671;
  wire CHOICE1880;
  wire N92659;
  wire N94673;
  wire N126620;
  wire CHOICE2112;
  wire N126473;
  wire CHOICE3225;
  wire N91567;
  wire N90291;
  wire N92711;
  wire CHOICE2470;
  wire CHOICE2254;
  wire N95468;
  wire CHOICE1425;
  wire CHOICE1446;
  wire DLX_IDlc_md_wint3;
  wire DLX_IDlc_md_wint1;
  wire CHOICE2257;
  wire CHOICE2446;
  wire CHOICE2278;
  wire CHOICE2924;
  wire DLX_IDlc_md_wint2;
  wire CHOICE2281;
  wire CHOICE2326;
  wire CHOICE2374;
  wire N127257;
  wire CHOICE2269;
  wire CHOICE2377;
  wire CHOICE3406;
  wire CHOICE1424;
  wire CHOICE2494;
  wire CHOICE2290;
  wire N126205;
  wire CHOICE2401;
  wire CHOICE2293;
  wire CHOICE2170;
  wire CHOICE2302;
  wire N126816;
  wire CHOICE2389;
  wire CHOICE2305;
  wire CHOICE2497;
  wire CHOICE2158;
  wire CHOICE2410;
  wire CHOICE2122;
  wire CHOICE2314;
  wire CHOICE2362;
  wire CHOICE2146;
  wire CHOICE2413;
  wire CHOICE2125;
  wire CHOICE2317;
  wire CHOICE2149;
  wire CHOICE2350;
  wire CHOICE2434;
  wire CHOICE2134;
  wire CHOICE2437;
  wire CHOICE2341;
  wire CHOICE1459;
  wire CHOICE1460;
  wire CHOICE2137;
  wire CHOICE2329;
  wire CHOICE2425;
  wire CHOICE2161;
  wire CHOICE1471;
  wire CHOICE1481;
  wire CHOICE2449;
  wire CHOICE2353;
  wire CHOICE2185;
  wire CHOICE2473;
  wire CHOICE2365;
  wire CHOICE2173;
  wire N90186;
  wire GLOBAL_LOGIC1_0;
  wire GLOBAL_LOGIC1_1;
  wire GLOBAL_LOGIC1_2;
  wire GLOBAL_LOGIC1_3;
  wire GLOBAL_LOGIC0_0;
  wire GLOBAL_LOGIC0_1;
  wire GLOBAL_LOGIC0_2;
  wire GLOBAL_LOGIC0_3;
  wire GLOBAL_LOGIC0_4;
  wire GLOBAL_LOGIC0_5;
  wire GLOBAL_LOGIC0_6;
  wire GLOBAL_LOGIC0_7;
  wire GLOBAL_LOGIC0_8;
  wire GLOBAL_LOGIC0_9;
  wire GLOBAL_LOGIC0_10;
  wire GSR = glbl.GSR;
  wire GTS = glbl.GTS;
  wire \mask<1>/ENABLE ;
  wire \mask<1>/TORGTS ;
  wire \mask<1>/OUTMUX ;
  wire \DM_write/OFF/RST ;
  wire \DM_write/ENABLE ;
  wire \DM_write/TORGTS ;
  wire \DM_write/OUTMUX ;
  wire DLX_EXinst_mem_write_EX_1;
  wire \DM_write/OD ;
  wire \mask<2>/ENABLE ;
  wire \mask<2>/TORGTS ;
  wire \mask<2>/OUTMUX ;
  wire \PIPEEMPTY/ENABLE ;
  wire \PIPEEMPTY/TORGTS ;
  wire \PIPEEMPTY/OUTMUX ;
  wire \clk_IF_del/ENABLE ;
  wire \clk_IF_del/TORGTS ;
  wire \clk_IF_del/OUTMUX ;
  wire \DM_addr_eff<10>/OFF/RST ;
  wire \DM_addr_eff<10>/ENABLE ;
  wire \DM_addr_eff<10>/TORGTS ;
  wire \DM_addr_eff<10>/OUTMUX ;
  wire DLX_EXinst_ALU_result_10_1;
  wire \DM_addr_eff<10>/OD ;
  wire \DM_addr_eff<11>/OFF/RST ;
  wire \DM_addr_eff<11>/ENABLE ;
  wire \DM_addr_eff<11>/TORGTS ;
  wire \DM_addr_eff<11>/OUTMUX ;
  wire DLX_EXinst_ALU_result_11_1;
  wire \DM_addr_eff<11>/OD ;
  wire \DM_addr_eff<12>/OFF/RST ;
  wire \DM_addr_eff<12>/ENABLE ;
  wire \DM_addr_eff<12>/TORGTS ;
  wire \DM_addr_eff<12>/OUTMUX ;
  wire DLX_EXinst_ALU_result_12_1;
  wire \DM_addr_eff<12>/OD ;
  wire \DM_addr_eff<13>/ENABLE ;
  wire \DM_addr_eff<13>/TORGTS ;
  wire \DM_addr_eff<13>/OUTMUX ;
  wire DLX_EXinst_ALU_result_13_1;
  wire \DM_addr_eff<13>/OD ;
  wire \DM_addr_eff<14>/ENABLE ;
  wire \DM_addr_eff<14>/TORGTS ;
  wire \DM_addr_eff<14>/OUTMUX ;
  wire DLX_EXinst_ALU_result_14_1;
  wire \DM_addr_eff<14>/OD ;
  wire \branch_sig/ENABLE ;
  wire \branch_sig/TORGTS ;
  wire \branch_sig/OUTMUX ;
  wire DLX_IDinst_branch_sig_1;
  wire \branch_sig/OD ;
  wire \clk_DM/ENABLE ;
  wire \clk_DM/TORGTS ;
  wire \clk_DM/OUTMUX ;
  wire \clk_ID/ENABLE ;
  wire \clk_ID/TORGTS ;
  wire \clk_ID/OUTMUX ;
  wire \clk_IF/ENABLE ;
  wire \clk_IF/TORGTS ;
  wire \clk_IF/OUTMUX ;
  wire \clk_EX/ENABLE ;
  wire \clk_EX/TORGTS ;
  wire \clk_EX/OUTMUX ;
  wire \hsync/ENABLE ;
  wire \hsync/TORGTS ;
  wire \hsync/OUTMUX ;
  wire vga_top_vga1_hsyncout;
  wire \hsync/LOGIC_ZERO ;
  wire \green<0>/ENABLE ;
  wire \green<0>/TORGTS ;
  wire \green<0>/OUTMUX ;
  wire \green<1>/ENABLE ;
  wire \green<1>/TORGTS ;
  wire \green<1>/OUTMUX ;
  wire \green<2>/ENABLE ;
  wire \green<2>/TORGTS ;
  wire \green<2>/OUTMUX ;
  wire \reset/IBUF ;
  wire \red<0>/ENABLE ;
  wire \red<0>/TORGTS ;
  wire \red<0>/OUTMUX ;
  wire \red<1>/ENABLE ;
  wire \red<1>/TORGTS ;
  wire \red<1>/OUTMUX ;
  wire \NPC_eff<0>/ENABLE ;
  wire \NPC_eff<0>/TORGTS ;
  wire \NPC_eff<0>/OUTMUX ;
  wire DLX_IFinst_NPC_0_1;
  wire \NPC_eff<0>/OD ;
  wire \DM_addr_eff<13>/OFF/RST ;
  wire \NPC_eff<1>/ENABLE ;
  wire \NPC_eff<1>/TORGTS ;
  wire \NPC_eff<1>/OUTMUX ;
  wire DLX_IFinst_NPC_1_1;
  wire \NPC_eff<1>/OD ;
  wire \NPC_eff<2>/ENABLE ;
  wire \NPC_eff<2>/TORGTS ;
  wire \NPC_eff<2>/OUTMUX ;
  wire DLX_IFinst_NPC_2_1;
  wire \NPC_eff<2>/OD ;
  wire \NPC_eff<3>/ENABLE ;
  wire \NPC_eff<3>/TORGTS ;
  wire \NPC_eff<3>/OUTMUX ;
  wire DLX_IFinst_NPC_3_1;
  wire \NPC_eff<3>/OD ;
  wire \NPC_eff<4>/ENABLE ;
  wire \NPC_eff<4>/TORGTS ;
  wire \NPC_eff<4>/OUTMUX ;
  wire DLX_IFinst_NPC_4_1;
  wire \NPC_eff<4>/OD ;
  wire \NPC_eff<5>/ENABLE ;
  wire \NPC_eff<5>/TORGTS ;
  wire \NPC_eff<5>/OUTMUX ;
  wire DLX_IFinst_NPC_5_1;
  wire \NPC_eff<5>/OD ;
  wire \NPC_eff<6>/ENABLE ;
  wire \NPC_eff<6>/TORGTS ;
  wire \NPC_eff<6>/OUTMUX ;
  wire DLX_IFinst_NPC_6_1;
  wire \NPC_eff<6>/OD ;
  wire \NPC_eff<7>/ENABLE ;
  wire \NPC_eff<7>/TORGTS ;
  wire \NPC_eff<7>/OUTMUX ;
  wire DLX_IFinst_NPC_7_1;
  wire \NPC_eff<7>/OD ;
  wire \NPC_eff<8>/ENABLE ;
  wire \NPC_eff<8>/TORGTS ;
  wire \NPC_eff<8>/OUTMUX ;
  wire DLX_IFinst_NPC_8_1;
  wire \NPC_eff<8>/OD ;
  wire \NPC_eff<9>/ENABLE ;
  wire \NPC_eff<9>/TORGTS ;
  wire \NPC_eff<9>/OUTMUX ;
  wire DLX_IFinst_NPC_9_1;
  wire \NPC_eff<9>/OD ;
  wire \stall/ENABLE ;
  wire \stall/TORGTS ;
  wire \stall/OUTMUX ;
  wire DLX_IDinst_stall_1;
  wire \stall/OD ;
  wire \CLI/ENABLE ;
  wire \CLI/TORGTS ;
  wire \CLI/OUTMUX ;
  wire DLX_IDinst_CLI_1;
  wire \CLI/OD ;
  wire \INT/IBUF ;
  wire \DM_addr_eff<0>/ENABLE ;
  wire \DM_addr_eff<0>/TORGTS ;
  wire \DM_addr_eff<0>/OUTMUX ;
  wire DLX_EXinst_ALU_result_0_1;
  wire \DM_addr_eff<0>/OD ;
  wire \DM_addr_eff<1>/ENABLE ;
  wire \DM_addr_eff<1>/TORGTS ;
  wire \DM_addr_eff<1>/OUTMUX ;
  wire DLX_EXinst_ALU_result_1_1;
  wire \DM_addr_eff<1>/OD ;
  wire \DM_addr_eff<2>/ENABLE ;
  wire \DM_addr_eff<2>/TORGTS ;
  wire \DM_addr_eff<2>/OUTMUX ;
  wire DLX_EXinst_ALU_result_2_1;
  wire \DM_addr_eff<2>/OD ;
  wire \DM_addr_eff<3>/ENABLE ;
  wire \DM_addr_eff<3>/TORGTS ;
  wire \DM_addr_eff<3>/OUTMUX ;
  wire DLX_EXinst_ALU_result_3_1;
  wire \DM_addr_eff<3>/OD ;
  wire \DM_addr_eff<4>/ENABLE ;
  wire \DM_addr_eff<4>/TORGTS ;
  wire \DM_addr_eff<4>/OUTMUX ;
  wire DLX_EXinst_ALU_result_4_1;
  wire \DM_addr_eff<4>/OD ;
  wire \DM_addr_eff<14>/OFF/RST ;
  wire \DM_addr_eff<5>/ENABLE ;
  wire \DM_addr_eff<5>/TORGTS ;
  wire \DM_addr_eff<5>/OUTMUX ;
  wire DLX_EXinst_ALU_result_5_1;
  wire \DM_addr_eff<5>/OD ;
  wire \DM_addr_eff<6>/ENABLE ;
  wire \DM_addr_eff<6>/TORGTS ;
  wire \DM_addr_eff<6>/OUTMUX ;
  wire DLX_EXinst_ALU_result_6_1;
  wire \DM_addr_eff<6>/OD ;
  wire \DM_addr_eff<7>/ENABLE ;
  wire \DM_addr_eff<7>/TORGTS ;
  wire \DM_addr_eff<7>/OUTMUX ;
  wire DLX_EXinst_ALU_result_7_1;
  wire \DM_addr_eff<7>/OD ;
  wire \DM_addr_eff<8>/ENABLE ;
  wire \DM_addr_eff<8>/TORGTS ;
  wire \DM_addr_eff<8>/OUTMUX ;
  wire DLX_EXinst_ALU_result_8_1;
  wire \DM_addr_eff<8>/OD ;
  wire \DM_addr_eff<9>/ENABLE ;
  wire \DM_addr_eff<9>/TORGTS ;
  wire \DM_addr_eff<9>/OUTMUX ;
  wire DLX_EXinst_ALU_result_9_1;
  wire \DM_addr_eff<9>/OD ;
  wire \vsync/ENABLE ;
  wire \vsync/TORGTS ;
  wire \vsync/OUTMUX ;
  wire vga_top_vga1_vsyncout;
  wire \vsync/LOGIC_ZERO ;
  wire \FREEZE/IBUF ;
  wire \IR_MSB<0>/ENABLE ;
  wire \IR_MSB<0>/TORGTS ;
  wire \IR_MSB<0>/OUTMUX ;
  wire \IR_MSB<1>/ENABLE ;
  wire \IR_MSB<1>/TORGTS ;
  wire \IR_MSB<1>/OUTMUX ;
  wire \IR_MSB<2>/ENABLE ;
  wire \IR_MSB<2>/TORGTS ;
  wire \IR_MSB<2>/OUTMUX ;
  wire \IR_MSB<3>/ENABLE ;
  wire \IR_MSB<3>/TORGTS ;
  wire \IR_MSB<3>/OUTMUX ;
  wire \IR_MSB<4>/ENABLE ;
  wire \IR_MSB<4>/TORGTS ;
  wire \IR_MSB<4>/OUTMUX ;
  wire \IR_MSB<5>/ENABLE ;
  wire \IR_MSB<5>/TORGTS ;
  wire \IR_MSB<5>/OUTMUX ;
  wire \IR_MSB<6>/ENABLE ;
  wire \IR_MSB<6>/TORGTS ;
  wire \IR_MSB<6>/OUTMUX ;
  wire \IR_MSB<7>/ENABLE ;
  wire \IR_MSB<7>/TORGTS ;
  wire \IR_MSB<7>/OUTMUX ;
  wire \delay_selectDM<0>/IBUF ;
  wire \delay_selectDM<1>/IBUF ;
  wire \branch_sig/OFF/RST ;
  wire \delay_selectID<0>/IBUF ;
  wire \delay_selectID<1>/IBUF ;
  wire \clk_MEM/ENABLE ;
  wire \clk_MEM/TORGTS ;
  wire \clk_MEM/OUTMUX ;
  wire \clk_MEM/ODNOT ;
  wire \delay_selectIF<0>/IBUF ;
  wire \delay_selectIF<1>/IBUF ;
  wire \delay_selectMEM<0>/IBUF ;
  wire \delay_selectMEM<1>/IBUF ;
  wire \blue<0>/ENABLE ;
  wire \blue<0>/TORGTS ;
  wire \blue<0>/OUTMUX ;
  wire \blue<1>/ENABLE ;
  wire \blue<1>/TORGTS ;
  wire \blue<1>/OUTMUX ;
  wire \blue<2>/ENABLE ;
  wire \blue<2>/TORGTS ;
  wire \blue<2>/OUTMUX ;
  wire \STOP_fetch/IBUF ;
  wire \delay_selectEX<0>/IBUF ;
  wire \delay_selectEX<1>/IBUF ;
  wire \mask<0>/ENABLE ;
  wire \mask<0>/TORGTS ;
  wire \mask<0>/OUTMUX ;
  wire \delay_selectRF<0>/IBUF ;
  wire \delay_selectRF<1>/IBUF ;
  wire \DM_read/ENABLE ;
  wire \DM_read/TORGTS ;
  wire \DM_read/OUTMUX ;
  wire DLX_EXinst_mem_read_EX_1;
  wire \DM_read/OD ;
  wire \mask<3>/ENABLE ;
  wire \mask<3>/TORGTS ;
  wire \mask<3>/OUTMUX ;
  wire \NPC_eff<10>/ENABLE ;
  wire \NPC_eff<10>/TORGTS ;
  wire \NPC_eff<10>/OUTMUX ;
  wire DLX_IFinst_NPC_10_1;
  wire \NPC_eff<10>/OD ;
  wire \NPC_eff<11>/ENABLE ;
  wire \NPC_eff<11>/TORGTS ;
  wire \NPC_eff<11>/OUTMUX ;
  wire DLX_IFinst_NPC_11_1;
  wire \NPC_eff<11>/OD ;
  wire \NPC_eff<12>/ENABLE ;
  wire \NPC_eff<12>/TORGTS ;
  wire \NPC_eff<12>/OUTMUX ;
  wire DLX_IFinst_NPC_12_1;
  wire \NPC_eff<12>/OD ;
  wire \NPC_eff<13>/ENABLE ;
  wire \NPC_eff<13>/TORGTS ;
  wire \NPC_eff<13>/OUTMUX ;
  wire DLX_IFinst_NPC_13_1;
  wire \NPC_eff<13>/OD ;
  wire \NPC_eff<14>/ENABLE ;
  wire \NPC_eff<14>/TORGTS ;
  wire \NPC_eff<14>/OUTMUX ;
  wire DLX_IFinst_NPC_14_1;
  wire \NPC_eff<14>/OD ;
  wire \NPC_eff<15>/ENABLE ;
  wire \NPC_eff<15>/TORGTS ;
  wire \NPC_eff<15>/OUTMUX ;
  wire DLX_IFinst_NPC_15_1;
  wire \NPC_eff<15>/OD ;
  wire \DM_write_data<0>/ENABLE ;
  wire \DM_write_data<0>/TORGTS ;
  wire \DM_write_data<0>/OUTMUX ;
  wire DLX_EXinst_reg_out_B_EX_0_1;
  wire \DM_write_data<0>/OD ;
  wire \clkdivider/LOCKED ;
  wire \clkdivider/CLK2X180 ;
  wire \clkdivider/CLK2X ;
  wire \clkdivider/CLK270 ;
  wire \clkdivider/CLK180 ;
  wire \clkdivider/CLK90 ;
  wire \clkdivider/LOGIC_ZERO ;
  wire \DLX_IDinst_RF_block0s0/DOB15 ;
  wire \DLX_IDinst_RF_block0s0/DOB14 ;
  wire \DLX_IDinst_RF_block0s0/DOB13 ;
  wire \DLX_IDinst_RF_block0s0/DOB12 ;
  wire \DLX_IDinst_RF_block0s0/DOB11 ;
  wire \DLX_IDinst_RF_block0s0/DOB10 ;
  wire \DLX_IDinst_RF_block0s0/DOB9 ;
  wire \DLX_IDinst_RF_block0s0/DOB8 ;
  wire \DLX_IDinst_RF_block0s0/DOB7 ;
  wire \DLX_IDinst_RF_block0s0/DOB6 ;
  wire \DLX_IDinst_RF_block0s0/DOB5 ;
  wire \DLX_IDinst_RF_block0s0/DOB4 ;
  wire \DLX_IDinst_RF_block0s0/DOB3 ;
  wire \DLX_IDinst_RF_block0s0/DOB2 ;
  wire \DLX_IDinst_RF_block0s0/DOB1 ;
  wire \DLX_IDinst_RF_block0s0/DOB0 ;
  wire \DLX_IDinst_RF_block0s0/DIA15 ;
  wire \DLX_IDinst_RF_block0s0/DIA14 ;
  wire \DLX_IDinst_RF_block0s0/DIA13 ;
  wire \DLX_IDinst_RF_block0s0/DIA12 ;
  wire \DLX_IDinst_RF_block0s0/DIA11 ;
  wire \DLX_IDinst_RF_block0s0/DIA10 ;
  wire \DLX_IDinst_RF_block0s0/DIA9 ;
  wire \DLX_IDinst_RF_block0s0/DIA8 ;
  wire \DLX_IDinst_RF_block0s0/DIA7 ;
  wire \DLX_IDinst_RF_block0s0/DIA6 ;
  wire \DLX_IDinst_RF_block0s0/DIA5 ;
  wire \DLX_IDinst_RF_block0s0/DIA4 ;
  wire \DLX_IDinst_RF_block0s0/DIA3 ;
  wire \DLX_IDinst_RF_block0s0/DIA2 ;
  wire \DLX_IDinst_RF_block0s0/DIA1 ;
  wire \DLX_IDinst_RF_block0s0/DIA0 ;
  wire \DLX_IDinst_RF_block0s0/ADDRB3 ;
  wire \DLX_IDinst_RF_block0s0/ADDRB2 ;
  wire \DLX_IDinst_RF_block0s0/ADDRB1 ;
  wire \DLX_IDinst_RF_block0s0/ADDRB0 ;
  wire \DLX_IDinst_RF_block0s0/ADDRA3 ;
  wire \DLX_IDinst_RF_block0s0/ADDRA2 ;
  wire \DLX_IDinst_RF_block0s0/ADDRA1 ;
  wire \DLX_IDinst_RF_block0s0/ADDRA0 ;
  wire \DLX_IDinst_RF_block0s0/LOGIC_ZERO ;
  wire \DLX_IDinst_RF_block0s1/DOB15 ;
  wire \DLX_IDinst_RF_block0s1/DOB14 ;
  wire \DLX_IDinst_RF_block0s1/DOB13 ;
  wire \DLX_IDinst_RF_block0s1/DOB12 ;
  wire \DLX_IDinst_RF_block0s1/DOB11 ;
  wire \DLX_IDinst_RF_block0s1/DOB10 ;
  wire \DLX_IDinst_RF_block0s1/DOB9 ;
  wire \DLX_IDinst_RF_block0s1/DOB8 ;
  wire \DLX_IDinst_RF_block0s1/DOB7 ;
  wire \DLX_IDinst_RF_block0s1/DOB6 ;
  wire \DLX_IDinst_RF_block0s1/DOB5 ;
  wire \DLX_IDinst_RF_block0s1/DOB4 ;
  wire \DLX_IDinst_RF_block0s1/DOB3 ;
  wire \DLX_IDinst_RF_block0s1/DOB2 ;
  wire \DLX_IDinst_RF_block0s1/DOB1 ;
  wire \DLX_IDinst_RF_block0s1/DOB0 ;
  wire \DLX_IDinst_RF_block0s1/DIA15 ;
  wire \DLX_IDinst_RF_block0s1/DIA14 ;
  wire \DLX_IDinst_RF_block0s1/DIA13 ;
  wire \DLX_IDinst_RF_block0s1/DIA12 ;
  wire \DLX_IDinst_RF_block0s1/DIA11 ;
  wire \DLX_IDinst_RF_block0s1/DIA10 ;
  wire \DLX_IDinst_RF_block0s1/DIA9 ;
  wire \DLX_IDinst_RF_block0s1/DIA8 ;
  wire \DLX_IDinst_RF_block0s1/DIA7 ;
  wire \DLX_IDinst_RF_block0s1/DIA6 ;
  wire \DLX_IDinst_RF_block0s1/DIA5 ;
  wire \DLX_IDinst_RF_block0s1/DIA4 ;
  wire \DLX_IDinst_RF_block0s1/DIA3 ;
  wire \DLX_IDinst_RF_block0s1/DIA2 ;
  wire \DLX_IDinst_RF_block0s1/DIA1 ;
  wire \DLX_IDinst_RF_block0s1/DIA0 ;
  wire \DLX_IDinst_RF_block0s1/ADDRB3 ;
  wire \DLX_IDinst_RF_block0s1/ADDRB2 ;
  wire \DLX_IDinst_RF_block0s1/ADDRB1 ;
  wire \DLX_IDinst_RF_block0s1/ADDRB0 ;
  wire \DLX_IDinst_RF_block0s1/ADDRA3 ;
  wire \DLX_IDinst_RF_block0s1/ADDRA2 ;
  wire \DLX_IDinst_RF_block0s1/ADDRA1 ;
  wire \DLX_IDinst_RF_block0s1/ADDRA0 ;
  wire \DLX_IDinst_RF_block0s1/LOGIC_ZERO ;
  wire \DLX_IDinst_RF_block1s0/DOB15 ;
  wire \DLX_IDinst_RF_block1s0/DOB14 ;
  wire \DLX_IDinst_RF_block1s0/DOB13 ;
  wire \DLX_IDinst_RF_block1s0/DOB12 ;
  wire \DLX_IDinst_RF_block1s0/DOB11 ;
  wire \DLX_IDinst_RF_block1s0/DOB10 ;
  wire \DLX_IDinst_RF_block1s0/DOB9 ;
  wire \DLX_IDinst_RF_block1s0/DOB8 ;
  wire \DLX_IDinst_RF_block1s0/DOB7 ;
  wire \DLX_IDinst_RF_block1s0/DOB6 ;
  wire \DLX_IDinst_RF_block1s0/DOB5 ;
  wire \DLX_IDinst_RF_block1s0/DOB4 ;
  wire \DLX_IDinst_RF_block1s0/DOB3 ;
  wire \DLX_IDinst_RF_block1s0/DOB2 ;
  wire \DLX_IDinst_RF_block1s0/DOB1 ;
  wire \DLX_IDinst_RF_block1s0/DOB0 ;
  wire \DLX_IDinst_RF_block1s0/DIA15 ;
  wire \DLX_IDinst_RF_block1s0/DIA14 ;
  wire \DLX_IDinst_RF_block1s0/DIA13 ;
  wire \DLX_IDinst_RF_block1s0/DIA12 ;
  wire \DLX_IDinst_RF_block1s0/DIA11 ;
  wire \DLX_IDinst_RF_block1s0/DIA10 ;
  wire \DLX_IDinst_RF_block1s0/DIA9 ;
  wire \DLX_IDinst_RF_block1s0/DIA8 ;
  wire \DLX_IDinst_RF_block1s0/DIA7 ;
  wire \DLX_IDinst_RF_block1s0/DIA6 ;
  wire \DLX_IDinst_RF_block1s0/DIA5 ;
  wire \DLX_IDinst_RF_block1s0/DIA4 ;
  wire \DLX_IDinst_RF_block1s0/DIA3 ;
  wire \DLX_IDinst_RF_block1s0/DIA2 ;
  wire \DLX_IDinst_RF_block1s0/DIA1 ;
  wire \DLX_IDinst_RF_block1s0/DIA0 ;
  wire \DLX_IDinst_RF_block1s0/ADDRB3 ;
  wire \DLX_IDinst_RF_block1s0/ADDRB2 ;
  wire \DLX_IDinst_RF_block1s0/ADDRB1 ;
  wire \DLX_IDinst_RF_block1s0/ADDRB0 ;
  wire \DLX_IDinst_RF_block1s0/ADDRA3 ;
  wire \DLX_IDinst_RF_block1s0/ADDRA2 ;
  wire \DLX_IDinst_RF_block1s0/ADDRA1 ;
  wire \DLX_IDinst_RF_block1s0/ADDRA0 ;
  wire \DLX_IDinst_RF_block1s0/LOGIC_ZERO ;
  wire \DLX_IDinst_RF_block1s1/DOB15 ;
  wire \DLX_IDinst_RF_block1s1/DOB14 ;
  wire \DLX_IDinst_RF_block1s1/DOB13 ;
  wire \DLX_IDinst_RF_block1s1/DOB12 ;
  wire \DLX_IDinst_RF_block1s1/DOB11 ;
  wire \DLX_IDinst_RF_block1s1/DOB10 ;
  wire \DLX_IDinst_RF_block1s1/DOB9 ;
  wire \DLX_IDinst_RF_block1s1/DOB8 ;
  wire \DLX_IDinst_RF_block1s1/DOB7 ;
  wire \DLX_IDinst_RF_block1s1/DOB6 ;
  wire \DLX_IDinst_RF_block1s1/DOB5 ;
  wire \DLX_IDinst_RF_block1s1/DOB4 ;
  wire \DLX_IDinst_RF_block1s1/DOB3 ;
  wire \DLX_IDinst_RF_block1s1/DOB2 ;
  wire \DLX_IDinst_RF_block1s1/DOB1 ;
  wire \DLX_IDinst_RF_block1s1/DOB0 ;
  wire \DLX_IDinst_RF_block1s1/DIA15 ;
  wire \DLX_IDinst_RF_block1s1/DIA14 ;
  wire \DLX_IDinst_RF_block1s1/DIA13 ;
  wire \DLX_IDinst_RF_block1s1/DIA12 ;
  wire \DLX_IDinst_RF_block1s1/DIA11 ;
  wire \DLX_IDinst_RF_block1s1/DIA10 ;
  wire \DLX_IDinst_RF_block1s1/DIA9 ;
  wire \DLX_IDinst_RF_block1s1/DIA8 ;
  wire \DLX_IDinst_RF_block1s1/DIA7 ;
  wire \DLX_IDinst_RF_block1s1/DIA6 ;
  wire \DLX_IDinst_RF_block1s1/DIA5 ;
  wire \DLX_IDinst_RF_block1s1/DIA4 ;
  wire \DLX_IDinst_RF_block1s1/DIA3 ;
  wire \DLX_IDinst_RF_block1s1/DIA2 ;
  wire \DLX_IDinst_RF_block1s1/DIA1 ;
  wire \DLX_IDinst_RF_block1s1/DIA0 ;
  wire \DLX_IDinst_RF_block1s1/ADDRB3 ;
  wire \DLX_IDinst_RF_block1s1/ADDRB2 ;
  wire \DLX_IDinst_RF_block1s1/ADDRB1 ;
  wire \DLX_IDinst_RF_block1s1/ADDRB0 ;
  wire \DLX_IDinst_RF_block1s1/ADDRA3 ;
  wire \DLX_IDinst_RF_block1s1/ADDRA2 ;
  wire \DLX_IDinst_RF_block1s1/ADDRA1 ;
  wire \DLX_IDinst_RF_block1s1/ADDRA0 ;
  wire \DLX_IDinst_RF_block1s1/LOGIC_ZERO ;
  wire \block0/DOB15 ;
  wire \block0/DOB14 ;
  wire \block0/DOB13 ;
  wire \block0/DOB12 ;
  wire \block0/DOB11 ;
  wire \block0/DOB10 ;
  wire \block0/DOB9 ;
  wire \block0/DOB8 ;
  wire \block0/DOA15 ;
  wire \block0/DOA14 ;
  wire \block0/DOA13 ;
  wire \block0/DOA12 ;
  wire \block0/DOA11 ;
  wire \block0/DOA10 ;
  wire \block0/DOA9 ;
  wire \block0/DOA8 ;
  wire \block0/DIB15 ;
  wire \block0/DIB14 ;
  wire \block0/DIB13 ;
  wire \block0/DIB12 ;
  wire \block0/DIB11 ;
  wire \block0/DIB10 ;
  wire \block0/DIB9 ;
  wire \block0/DIB8 ;
  wire \block0/DIB7 ;
  wire \block0/DIB6 ;
  wire \block0/DIB5 ;
  wire \block0/DIB4 ;
  wire \block0/DIB3 ;
  wire \block0/DIB2 ;
  wire \block0/DIB1 ;
  wire \block0/DIB0 ;
  wire \block0/DIA15 ;
  wire \block0/DIA14 ;
  wire \block0/DIA13 ;
  wire \block0/DIA12 ;
  wire \block0/DIA11 ;
  wire \block0/DIA10 ;
  wire \block0/DIA9 ;
  wire \block0/DIA8 ;
  wire \block0/ADDRB2 ;
  wire \block0/ADDRB1 ;
  wire \block0/ADDRB0 ;
  wire \block0/ADDRA2 ;
  wire \block0/ADDRA1 ;
  wire \block0/ADDRA0 ;
  wire \block0/LOGIC_ZERO ;
  wire \block0/LOGIC_ONE ;
  wire \block1/DOB15 ;
  wire \block1/DOB14 ;
  wire \block1/DOB13 ;
  wire \block1/DOB12 ;
  wire \block1/DOB11 ;
  wire \block1/DOB10 ;
  wire \block1/DOB9 ;
  wire \block1/DOB8 ;
  wire \block1/DOA15 ;
  wire \block1/DOA14 ;
  wire \block1/DOA13 ;
  wire \block1/DOA12 ;
  wire \block1/DOA11 ;
  wire \block1/DOA10 ;
  wire \block1/DOA9 ;
  wire \block1/DOA8 ;
  wire \block1/DIB15 ;
  wire \block1/DIB14 ;
  wire \block1/DIB13 ;
  wire \block1/DIB12 ;
  wire \block1/DIB11 ;
  wire \block1/DIB10 ;
  wire \block1/DIB9 ;
  wire \block1/DIB8 ;
  wire \block1/DIB7 ;
  wire \block1/DIB6 ;
  wire \block1/DIB5 ;
  wire \block1/DIB4 ;
  wire \block1/DIB3 ;
  wire \block1/DIB2 ;
  wire \block1/DIB1 ;
  wire \block1/DIB0 ;
  wire \block1/DIA15 ;
  wire \block1/DIA14 ;
  wire \block1/DIA13 ;
  wire \block1/DIA12 ;
  wire \block1/DIA11 ;
  wire \block1/DIA10 ;
  wire \block1/DIA9 ;
  wire \block1/DIA8 ;
  wire \block1/ADDRB2 ;
  wire \block1/ADDRB1 ;
  wire \block1/ADDRB0 ;
  wire \block1/ADDRA2 ;
  wire \block1/ADDRA1 ;
  wire \block1/ADDRA0 ;
  wire \block1/LOGIC_ZERO ;
  wire \block1/LOGIC_ONE ;
  wire \block2/DOB15 ;
  wire \block2/DOB14 ;
  wire \block2/DOB13 ;
  wire \block2/DOB12 ;
  wire \block2/DOB11 ;
  wire \block2/DOB10 ;
  wire \block2/DOB9 ;
  wire \block2/DOB8 ;
  wire \block2/DOA15 ;
  wire \block2/DOA14 ;
  wire \block2/DOA13 ;
  wire \block2/DOA12 ;
  wire \block2/DOA11 ;
  wire \block2/DOA10 ;
  wire \block2/DOA9 ;
  wire \block2/DOA8 ;
  wire \block2/DIB15 ;
  wire \block2/DIB14 ;
  wire \block2/DIB13 ;
  wire \block2/DIB12 ;
  wire \block2/DIB11 ;
  wire \block2/DIB10 ;
  wire \block2/DIB9 ;
  wire \block2/DIB8 ;
  wire \block2/DIB7 ;
  wire \block2/DIB6 ;
  wire \block2/DIB5 ;
  wire \block2/DIB4 ;
  wire \block2/DIB3 ;
  wire \block2/DIB2 ;
  wire \block2/DIB1 ;
  wire \block2/DIB0 ;
  wire \block2/DIA15 ;
  wire \block2/DIA14 ;
  wire \block2/DIA13 ;
  wire \block2/DIA12 ;
  wire \block2/DIA11 ;
  wire \block2/DIA10 ;
  wire \block2/DIA9 ;
  wire \block2/DIA8 ;
  wire \block2/ADDRB2 ;
  wire \block2/ADDRB1 ;
  wire \block2/ADDRB0 ;
  wire \block2/ADDRA2 ;
  wire \block2/ADDRA1 ;
  wire \block2/ADDRA0 ;
  wire \block2/LOGIC_ZERO ;
  wire \block2/LOGIC_ONE ;
  wire \block3/DOB15 ;
  wire \block3/DOB14 ;
  wire \block3/DOB13 ;
  wire \block3/DOB12 ;
  wire \block3/DOB11 ;
  wire \block3/DOB10 ;
  wire \block3/DOB9 ;
  wire \block3/DOB8 ;
  wire \block3/DOA15 ;
  wire \block3/DOA14 ;
  wire \block3/DOA13 ;
  wire \block3/DOA12 ;
  wire \block3/DOA11 ;
  wire \block3/DOA10 ;
  wire \block3/DOA9 ;
  wire \block3/DOA8 ;
  wire \block3/DIB15 ;
  wire \block3/DIB14 ;
  wire \block3/DIB13 ;
  wire \block3/DIB12 ;
  wire \block3/DIB11 ;
  wire \block3/DIB10 ;
  wire \block3/DIB9 ;
  wire \block3/DIB8 ;
  wire \block3/DIB7 ;
  wire \block3/DIB6 ;
  wire \block3/DIB5 ;
  wire \block3/DIB4 ;
  wire \block3/DIB3 ;
  wire \block3/DIB2 ;
  wire \block3/DIB1 ;
  wire \block3/DIB0 ;
  wire \block3/DIA15 ;
  wire \block3/DIA14 ;
  wire \block3/DIA13 ;
  wire \block3/DIA12 ;
  wire \block3/DIA11 ;
  wire \block3/DIA10 ;
  wire \block3/DIA9 ;
  wire \block3/DIA8 ;
  wire \block3/ADDRB2 ;
  wire \block3/ADDRB1 ;
  wire \block3/ADDRB0 ;
  wire \block3/ADDRA2 ;
  wire \block3/ADDRA1 ;
  wire \block3/ADDRA0 ;
  wire \block3/LOGIC_ZERO ;
  wire \block3/LOGIC_ONE ;
  wire \vga0/DOB15 ;
  wire \vga0/DOB14 ;
  wire \vga0/DOB13 ;
  wire \vga0/DOB12 ;
  wire \vga0/DOB11 ;
  wire \vga0/DOB10 ;
  wire \vga0/DOB9 ;
  wire \vga0/DOB8 ;
  wire \vga0/DOB7 ;
  wire \vga0/DOB6 ;
  wire \vga0/DOB5 ;
  wire \vga0/DOB4 ;
  wire \vga0/DOB3 ;
  wire \vga0/DOB2 ;
  wire \vga0/DOB1 ;
  wire \vga0/DOA15 ;
  wire \vga0/DOA14 ;
  wire \vga0/DOA13 ;
  wire \vga0/DOA12 ;
  wire \vga0/DOA11 ;
  wire \vga0/DOA10 ;
  wire \vga0/DOA9 ;
  wire \vga0/DOA8 ;
  wire \vga0/DOA7 ;
  wire \vga0/DOA6 ;
  wire \vga0/DOA5 ;
  wire \vga0/DOA4 ;
  wire \vga0/DOA3 ;
  wire \vga0/DOA2 ;
  wire \vga0/DOA1 ;
  wire \vga0/DIB15 ;
  wire \vga0/DIB14 ;
  wire \vga0/DIB13 ;
  wire \vga0/DIB12 ;
  wire \vga0/DIB11 ;
  wire \vga0/DIB10 ;
  wire \vga0/DIB9 ;
  wire \vga0/DIB8 ;
  wire \vga0/DIB7 ;
  wire \vga0/DIB6 ;
  wire \vga0/DIB5 ;
  wire \vga0/DIB4 ;
  wire \vga0/DIB3 ;
  wire \vga0/DIB2 ;
  wire \vga0/DIB1 ;
  wire \vga0/DIB0 ;
  wire \vga0/DIA15 ;
  wire \vga0/DIA14 ;
  wire \vga0/DIA13 ;
  wire \vga0/DIA12 ;
  wire \vga0/DIA11 ;
  wire \vga0/DIA10 ;
  wire \vga0/DIA9 ;
  wire \vga0/DIA8 ;
  wire \vga0/DIA7 ;
  wire \vga0/DIA6 ;
  wire \vga0/DIA5 ;
  wire \vga0/DIA4 ;
  wire \vga0/DIA3 ;
  wire \vga0/DIA2 ;
  wire \vga0/DIA1 ;
  wire \vga0/LOGIC_ZERO ;
  wire \vga0/LOGIC_ONE ;
  wire \vga1/DOB15 ;
  wire \vga1/DOB14 ;
  wire \vga1/DOB13 ;
  wire \vga1/DOB12 ;
  wire \vga1/DOB11 ;
  wire \vga1/DOB10 ;
  wire \vga1/DOB9 ;
  wire \vga1/DOB8 ;
  wire \vga1/DOB7 ;
  wire \vga1/DOB6 ;
  wire \vga1/DOB5 ;
  wire \vga1/DOB4 ;
  wire \vga1/DOB3 ;
  wire \vga1/DOB2 ;
  wire \vga1/DOB1 ;
  wire \vga1/DOA15 ;
  wire \vga1/DOA14 ;
  wire \vga1/DOA13 ;
  wire \vga1/DOA12 ;
  wire \vga1/DOA11 ;
  wire \vga1/DOA10 ;
  wire \vga1/DOA9 ;
  wire \vga1/DOA8 ;
  wire \vga1/DOA7 ;
  wire \vga1/DOA6 ;
  wire \vga1/DOA5 ;
  wire \vga1/DOA4 ;
  wire \vga1/DOA3 ;
  wire \vga1/DOA2 ;
  wire \vga1/DOA1 ;
  wire \vga1/DIB15 ;
  wire \vga1/DIB14 ;
  wire \vga1/DIB13 ;
  wire \vga1/DIB12 ;
  wire \vga1/DIB11 ;
  wire \vga1/DIB10 ;
  wire \vga1/DIB9 ;
  wire \vga1/DIB8 ;
  wire \vga1/DIB7 ;
  wire \vga1/DIB6 ;
  wire \vga1/DIB5 ;
  wire \vga1/DIB4 ;
  wire \vga1/DIB3 ;
  wire \vga1/DIB2 ;
  wire \vga1/DIB1 ;
  wire \vga1/DIB0 ;
  wire \vga1/DIA15 ;
  wire \vga1/DIA14 ;
  wire \vga1/DIA13 ;
  wire \vga1/DIA12 ;
  wire \vga1/DIA11 ;
  wire \vga1/DIA10 ;
  wire \vga1/DIA9 ;
  wire \vga1/DIA8 ;
  wire \vga1/DIA7 ;
  wire \vga1/DIA6 ;
  wire \vga1/DIA5 ;
  wire \vga1/DIA4 ;
  wire \vga1/DIA3 ;
  wire \vga1/DIA2 ;
  wire \vga1/DIA1 ;
  wire \vga1/LOGIC_ZERO ;
  wire \vga1/LOGIC_ONE ;
  wire \vga2/DOB15 ;
  wire \vga2/DOB14 ;
  wire \vga2/DOB13 ;
  wire \vga2/DOB12 ;
  wire \vga2/DOB11 ;
  wire \vga2/DOB10 ;
  wire \vga2/DOB9 ;
  wire \vga2/DOB8 ;
  wire \vga2/DOB7 ;
  wire \vga2/DOB6 ;
  wire \vga2/DOB5 ;
  wire \vga2/DOB4 ;
  wire \vga2/DOB3 ;
  wire \vga2/DOB2 ;
  wire \vga2/DOB1 ;
  wire \vga2/DOA15 ;
  wire \vga2/DOA14 ;
  wire \vga2/DOA13 ;
  wire \vga2/DOA12 ;
  wire \vga2/DOA11 ;
  wire \vga2/DOA10 ;
  wire \vga2/DOA9 ;
  wire \vga2/DOA8 ;
  wire \vga2/DOA7 ;
  wire \vga2/DOA6 ;
  wire \vga2/DOA5 ;
  wire \vga2/DOA4 ;
  wire \vga2/DOA3 ;
  wire \vga2/DOA2 ;
  wire \vga2/DOA1 ;
  wire \vga2/DIB15 ;
  wire \vga2/DIB14 ;
  wire \vga2/DIB13 ;
  wire \vga2/DIB12 ;
  wire \vga2/DIB11 ;
  wire \vga2/DIB10 ;
  wire \vga2/DIB9 ;
  wire \vga2/DIB8 ;
  wire \vga2/DIB7 ;
  wire \vga2/DIB6 ;
  wire \vga2/DIB5 ;
  wire \vga2/DIB4 ;
  wire \vga2/DIB3 ;
  wire \vga2/DIB2 ;
  wire \vga2/DIB1 ;
  wire \vga2/DIB0 ;
  wire \vga2/DIA15 ;
  wire \vga2/DIA14 ;
  wire \vga2/DIA13 ;
  wire \vga2/DIA12 ;
  wire \vga2/DIA11 ;
  wire \vga2/DIA10 ;
  wire \vga2/DIA9 ;
  wire \vga2/DIA8 ;
  wire \vga2/DIA7 ;
  wire \vga2/DIA6 ;
  wire \vga2/DIA5 ;
  wire \vga2/DIA4 ;
  wire \vga2/DIA3 ;
  wire \vga2/DIA2 ;
  wire \vga2/DIA1 ;
  wire \vga2/LOGIC_ZERO ;
  wire \vga2/LOGIC_ONE ;
  wire \vga3/DOB15 ;
  wire \vga3/DOB14 ;
  wire \vga3/DOB13 ;
  wire \vga3/DOB12 ;
  wire \vga3/DOB11 ;
  wire \vga3/DOB10 ;
  wire \vga3/DOB9 ;
  wire \vga3/DOB8 ;
  wire \vga3/DOB7 ;
  wire \vga3/DOB6 ;
  wire \vga3/DOB5 ;
  wire \vga3/DOB4 ;
  wire \vga3/DOB3 ;
  wire \vga3/DOB2 ;
  wire \vga3/DOB1 ;
  wire \vga3/DOA15 ;
  wire \vga3/DOA14 ;
  wire \vga3/DOA13 ;
  wire \vga3/DOA12 ;
  wire \vga3/DOA11 ;
  wire \vga3/DOA10 ;
  wire \vga3/DOA9 ;
  wire \vga3/DOA8 ;
  wire \vga3/DOA7 ;
  wire \vga3/DOA6 ;
  wire \vga3/DOA5 ;
  wire \vga3/DOA4 ;
  wire \vga3/DOA3 ;
  wire \vga3/DOA2 ;
  wire \vga3/DOA1 ;
  wire \vga3/DIB15 ;
  wire \vga3/DIB14 ;
  wire \vga3/DIB13 ;
  wire \vga3/DIB12 ;
  wire \vga3/DIB11 ;
  wire \vga3/DIB10 ;
  wire \vga3/DIB9 ;
  wire \vga3/DIB8 ;
  wire \vga3/DIB7 ;
  wire \vga3/DIB6 ;
  wire \vga3/DIB5 ;
  wire \vga3/DIB4 ;
  wire \vga3/DIB3 ;
  wire \vga3/DIB2 ;
  wire \vga3/DIB1 ;
  wire \vga3/DIB0 ;
  wire \vga3/DIA15 ;
  wire \vga3/DIA14 ;
  wire \vga3/DIA13 ;
  wire \vga3/DIA12 ;
  wire \vga3/DIA11 ;
  wire \vga3/DIA10 ;
  wire \vga3/DIA9 ;
  wire \vga3/DIA8 ;
  wire \vga3/DIA7 ;
  wire \vga3/DIA6 ;
  wire \vga3/DIA5 ;
  wire \vga3/DIA4 ;
  wire \vga3/DIA3 ;
  wire \vga3/DIA2 ;
  wire \vga3/DIA1 ;
  wire \vga3/LOGIC_ZERO ;
  wire \vga3/LOGIC_ONE ;
  wire \vga4/DOB15 ;
  wire \vga4/DOB14 ;
  wire \vga4/DOB13 ;
  wire \vga4/DOB12 ;
  wire \vga4/DOB11 ;
  wire \vga4/DOB10 ;
  wire \vga4/DOB9 ;
  wire \vga4/DOB8 ;
  wire \vga4/DOB7 ;
  wire \vga4/DOB6 ;
  wire \vga4/DOB5 ;
  wire \vga4/DOB4 ;
  wire \vga4/DOB3 ;
  wire \vga4/DOB2 ;
  wire \vga4/DOB1 ;
  wire \vga4/DOA15 ;
  wire \vga4/DOA14 ;
  wire \vga4/DOA13 ;
  wire \vga4/DOA12 ;
  wire \vga4/DOA11 ;
  wire \vga4/DOA10 ;
  wire \vga4/DOA9 ;
  wire \vga4/DOA8 ;
  wire \vga4/DOA7 ;
  wire \vga4/DOA6 ;
  wire \vga4/DOA5 ;
  wire \vga4/DOA4 ;
  wire \vga4/DOA3 ;
  wire \vga4/DOA2 ;
  wire \vga4/DOA1 ;
  wire \vga4/DIB15 ;
  wire \vga4/DIB14 ;
  wire \vga4/DIB13 ;
  wire \vga4/DIB12 ;
  wire \vga4/DIB11 ;
  wire \vga4/DIB10 ;
  wire \vga4/DIB9 ;
  wire \vga4/DIB8 ;
  wire \vga4/DIB7 ;
  wire \vga4/DIB6 ;
  wire \vga4/DIB5 ;
  wire \vga4/DIB4 ;
  wire \vga4/DIB3 ;
  wire \vga4/DIB2 ;
  wire \vga4/DIB1 ;
  wire \vga4/DIB0 ;
  wire \vga4/DIA15 ;
  wire \vga4/DIA14 ;
  wire \vga4/DIA13 ;
  wire \vga4/DIA12 ;
  wire \vga4/DIA11 ;
  wire \vga4/DIA10 ;
  wire \vga4/DIA9 ;
  wire \vga4/DIA8 ;
  wire \vga4/DIA7 ;
  wire \vga4/DIA6 ;
  wire \vga4/DIA5 ;
  wire \vga4/DIA4 ;
  wire \vga4/DIA3 ;
  wire \vga4/DIA2 ;
  wire \vga4/DIA1 ;
  wire \vga4/LOGIC_ZERO ;
  wire \vga4/LOGIC_ONE ;
  wire N127641;
  wire N127639;
  wire \N108593/F5MUX ;
  wire N127701;
  wire N127699;
  wire \CHOICE3132/F5MUX ;
  wire N127686;
  wire N127684;
  wire \N107934/F5MUX ;
  wire N127926;
  wire N127924;
  wire \CHOICE3311/F5MUX ;
  wire N128066;
  wire N128064;
  wire \N126636/F5MUX ;
  wire N128096;
  wire N128094;
  wire \CHOICE1402/F5MUX ;
  wire N127946;
  wire N127944;
  wire \DLX_IFlc_md_outp2/F5MUX ;
  wire N127941;
  wire N127939;
  wire \DLX_IDlc_md_outp2/F5MUX ;
  wire N127936;
  wire N127934;
  wire \DLX_EXlc_md_outp2/F5MUX ;
  wire N127881;
  wire N127879;
  wire \CHOICE5509/F5MUX ;
  wire N127931;
  wire N127929;
  wire \DLX_MEMlc_md_outp2/F5MUX ;
  wire N127781;
  wire N127779;
  wire \N126486/F5MUX ;
  wire N127886;
  wire N127884;
  wire \DLX_IDinst_N69963/F5MUX ;
  wire N128001;
  wire N127999;
  wire \clk_EX_del/F5MUX ;
  wire N127696;
  wire N127694;
  wire N127786;
  wire N127784;
  wire N127906;
  wire N127904;
  wire N127676;
  wire N127674;
  wire N127996;
  wire N127994;
  wire \DLX_clk_IF_del/F5MUX ;
  wire N127756;
  wire N127754;
  wire N127666;
  wire N127664;
  wire N128101;
  wire N128099;
  wire N127841;
  wire N127839;
  wire N127706;
  wire N127704;
  wire N127861;
  wire N127859;
  wire N127851;
  wire N127849;
  wire N127751;
  wire N127749;
  wire N127921;
  wire N127919;
  wire \DLX_EXinst_Mshift__n0025_Sh<40>/F5MUX ;
  wire N128061;
  wire N128059;
  wire N127741;
  wire N127739;
  wire N127971;
  wire N127969;
  wire N127631;
  wire N127629;
  wire N127736;
  wire N127734;
  wire N127611;
  wire N127609;
  wire N127991;
  wire N127989;
  wire \DLX_EXinst_Mshift__n0025_Sh<43>/F5MUX ;
  wire N127811;
  wire N127809;
  wire N127651;
  wire N127649;
  wire N127916;
  wire N127914;
  wire N127836;
  wire N127834;
  wire N128086;
  wire N128084;
  wire \N126560/F5MUX ;
  wire N127791;
  wire N127789;
  wire \CHOICE5871/F5MUX ;
  wire N128046;
  wire N128044;
  wire \CHOICE5100/F5MUX ;
  wire N127721;
  wire N127719;
  wire \CHOICE5125/F5MUX ;
  wire N127866;
  wire N127864;
  wire \CHOICE5598/F5MUX ;
  wire N127896;
  wire N127894;
  wire \CHOICE5973/F5MUX ;
  wire N127656;
  wire N127654;
  wire \CHOICE1771/F5MUX ;
  wire N127766;
  wire N127764;
  wire \CHOICE5709/F5MUX ;
  wire N127826;
  wire N127824;
  wire \CHOICE5432/F5MUX ;
  wire N128011;
  wire N128009;
  wire \CHOICE5540/F5MUX ;
  wire N128071;
  wire N128069;
  wire \CHOICE4965/F5MUX ;
  wire N128021;
  wire N128019;
  wire \N101537/F5MUX ;
  wire N127726;
  wire N127724;
  wire \N95810/F5MUX ;
  wire N128036;
  wire N128034;
  wire \CHOICE2965/F5MUX ;
  wire N127621;
  wire N127619;
  wire \CHOICE3097/F5MUX ;
  wire N128056;
  wire N128054;
  wire \N97089/F5MUX ;
  wire N127801;
  wire N127799;
  wire \N97449/F5MUX ;
  wire N127616;
  wire N127614;
  wire \N100843/F5MUX ;
  wire N127856;
  wire N127854;
  wire \CHOICE5077/F5MUX ;
  wire N127761;
  wire N127759;
  wire \N97305/F5MUX ;
  wire Mmux__COND_2__net1;
  wire Mmux__COND_2__net0;
  wire \Mmux__COND_2__net2/F5MUX ;
  wire N128076;
  wire N128074;
  wire \N97375/F5MUX ;
  wire N127796;
  wire N127794;
  wire \N97161/F5MUX ;
  wire N127951;
  wire N127949;
  wire \N100919/F5MUX ;
  wire N128031;
  wire N128029;
  wire \N101009/F5MUX ;
  wire N127871;
  wire N127869;
  wire \N101253/F5MUX ;
  wire N127831;
  wire N127829;
  wire \N97521/F5MUX ;
  wire N127636;
  wire N127634;
  wire \CHOICE3198/F5MUX ;
  wire N127911;
  wire N127909;
  wire \CHOICE2542/F5MUX ;
  wire N127626;
  wire N127624;
  wire \DLX_EXinst_Mshift__n0027_Sh<40>/F5MUX ;
  wire N127891;
  wire N127889;
  wire \CHOICE3124/F5MUX ;
  wire N127691;
  wire N127689;
  wire \CHOICE4587/F5MUX ;
  wire N127596;
  wire N127594;
  wire \DLX_EXinst_Mshift__n0027_Sh<42>/F5MUX ;
  wire N127606;
  wire N127604;
  wire \DLX_EXinst_Mshift__n0027_Sh<43>/F5MUX ;
  wire N127806;
  wire N127804;
  wire \N126268/F5MUX ;
  wire N127816;
  wire N127814;
  wire \DLX_EXinst_N65090/F5MUX ;
  wire N127771;
  wire N127769;
  wire \DLX_EXinst_N64500/F5MUX ;
  wire N128081;
  wire N128079;
  wire N128006;
  wire N128004;
  wire N128041;
  wire N128039;
  wire N127981;
  wire N127979;
  wire N127961;
  wire N127959;
  wire N127986;
  wire N127984;
  wire N127876;
  wire N127874;
  wire N127966;
  wire N127964;
  wire N127746;
  wire N127744;
  wire N127776;
  wire N127774;
  wire N128091;
  wire N128089;
  wire \DLX_EXinst_Mshift__n0028_Sh<59>/F5MUX ;
  wire N127711;
  wire N127709;
  wire \CHOICE4531/F5MUX ;
  wire N127671;
  wire N127669;
  wire \N126500/F5MUX ;
  wire N127731;
  wire N127729;
  wire \CHOICE5297/F5MUX ;
  wire N127956;
  wire N127954;
  wire \N127444/F5MUX ;
  wire N127716;
  wire N127714;
  wire \CHOICE5815/F5MUX ;
  wire N127821;
  wire N127819;
  wire \CHOICE5842/F5MUX ;
  wire N128016;
  wire N128014;
  wire \CHOICE5166/F5MUX ;
  wire N127901;
  wire N127899;
  wire \CHOICE5140/F5MUX ;
  wire N128026;
  wire N128024;
  wire \CHOICE5637/F5MUX ;
  wire N127846;
  wire N127844;
  wire \CHOICE5471/F5MUX ;
  wire N127646;
  wire N127644;
  wire \CHOICE4994/F5MUX ;
  wire N127601;
  wire N127599;
  wire \CHOICE5222/F5MUX ;
  wire N127681;
  wire N127679;
  wire \CHOICE5374/F5MUX ;
  wire N127661;
  wire N127659;
  wire \N127440/F5MUX ;
  wire \NPC_eff<0>/OFF/RST ;
  wire N127976;
  wire N127974;
  wire \N126272/F5MUX ;
  wire \vram_out_vga_eff/LOGIC_ONE ;
  wire \vram_out_vga<4>_rt ;
  wire \vram_out_vga_eff/F6MUX ;
  wire \Mmux__COND_2_inst_mux_f6_0.F51 ;
  wire N128051;
  wire N128049;
  wire \DLX_EXinst_Mshift__n0023_Sh<27>/F5MUX ;
  wire \vga_top_vga1_Madd_addressout_inst_lut2_331/FROM ;
  wire \vga_top_vga1_Madd_addressout_inst_lut2_331/CYMUXG ;
  wire \vga_top_vga1_Madd_addressout_inst_lut2_331/XORG ;
  wire vga_top_vga1_Madd_addressout_inst_lut2_332;
  wire vga_top_vga1_Madd_addressout_inst_cy_465;
  wire \vga_top_vga1_Madd_addressout_inst_lut2_331/LOGIC_ZERO ;
  wire vga_top_vga1_Madd_addressout_inst_lut2_333;
  wire \vga_address<7>/XORF ;
  wire \vga_address<7>/CYMUXG ;
  wire \vga_address<7>/XORG ;
  wire vga_top_vga1_Madd_addressout_inst_lut2_334;
  wire vga_top_vga1_Madd_addressout_inst_cy_467;
  wire \vga_address<7>/CYINIT ;
  wire DLX_EXinst_Mcompar__n0061_inst_lut2_148;
  wire \DLX_EXinst_Mcompar__n0061_inst_cy_213/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0061_inst_lut2_149;
  wire DLX_EXinst_Mcompar__n0061_inst_cy_212;
  wire \DLX_EXinst_Mcompar__n0061_inst_cy_213/CYINIT ;
  wire DLX_EXinst_Mcompar__n0061_inst_lut2_150;
  wire \DLX_EXinst_Mcompar__n0061_inst_cy_215/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0061_inst_lut2_151;
  wire DLX_EXinst_Mcompar__n0061_inst_cy_214;
  wire \DLX_EXinst_Mcompar__n0061_inst_cy_215/CYINIT ;
  wire DLX_EXinst_Mcompar__n0061_inst_lut2_152;
  wire \DLX_EXinst_Mcompar__n0061_inst_cy_217/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0061_inst_lut2_153;
  wire DLX_EXinst_Mcompar__n0061_inst_cy_216;
  wire \DLX_EXinst_Mcompar__n0061_inst_cy_217/CYINIT ;
  wire DLX_EXinst_Mcompar__n0061_inst_lut2_154;
  wire \DLX_EXinst_Mcompar__n0061_inst_cy_219/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0061_inst_lut2_155;
  wire DLX_EXinst_Mcompar__n0061_inst_cy_218;
  wire \DLX_EXinst_Mcompar__n0061_inst_cy_219/CYINIT ;
  wire DLX_EXinst_Mcompar__n0061_inst_lut2_156;
  wire \DLX_EXinst_Mcompar__n0061_inst_cy_221/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0061_inst_lut2_157;
  wire DLX_EXinst_Mcompar__n0061_inst_cy_220;
  wire \DLX_EXinst_Mcompar__n0061_inst_cy_221/CYINIT ;
  wire DLX_EXinst_Mcompar__n0061_inst_lut2_158;
  wire \DLX_EXinst_Mcompar__n0061_inst_cy_223/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0061_inst_lut2_159;
  wire DLX_EXinst_Mcompar__n0061_inst_cy_222;
  wire \DLX_EXinst_Mcompar__n0061_inst_cy_223/CYINIT ;
  wire DLX_EXinst_Mcompar__n0061_inst_lut2_160;
  wire \DLX_EXinst_Mcompar__n0061_inst_cy_225/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0061_inst_lut2_161;
  wire DLX_EXinst_Mcompar__n0061_inst_cy_224;
  wire \DLX_EXinst_Mcompar__n0061_inst_cy_225/CYINIT ;
  wire DLX_EXinst_Mcompar__n0061_inst_lut2_162;
  wire \DLX_EXinst_Mcompar__n0061_inst_cy_227/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0061_inst_lut2_163;
  wire DLX_EXinst_Mcompar__n0061_inst_cy_226;
  wire \DLX_EXinst_Mcompar__n0061_inst_cy_227/CYINIT ;
  wire DLX_EXinst_Mcompar__n0061_inst_lut2_164;
  wire \DLX_EXinst_reg_out_B_EX<30>/CYMUXF ;
  wire \DLX_EXinst_reg_out_B_EX<30>/CYINIT ;
  wire vga_top_vga1_Mcompar__n0029_inst_lut1_22;
  wire \vga_top_vga1_Mcompar__n0029_inst_cy_374/CYMUXG ;
  wire vga_top_vga1_Mcompar__n0029_inst_lut1_23;
  wire vga_top_vga1_Mcompar__n0029_inst_cy_373;
  wire \vga_top_vga1_Mcompar__n0029_inst_cy_374/LOGIC_ZERO ;
  wire \vga_top_vga1_Mcompar__n0029_inst_cy_374/LOGIC_ONE ;
  wire \$SIG_13 ;
  wire \vga_top_vga1_Mcompar__n0029_inst_cy_376/CYMUXG ;
  wire \$SIG_14 ;
  wire vga_top_vga1_Mcompar__n0029_inst_cy_375;
  wire \vga_top_vga1_Mcompar__n0029_inst_cy_376/LOGIC_ONE ;
  wire \vga_top_vga1_Mcompar__n0029_inst_cy_376/CYINIT ;
  wire vga_top_vga1_Mcompar__n0029_inst_lut4_51;
  wire \vga_top_vga1_Mcompar__n0029_inst_cy_378/CYMUXG ;
  wire vga_top_vga1_Mcompar__n0029_inst_lut4_52;
  wire vga_top_vga1_Mcompar__n0029_inst_cy_377;
  wire \vga_top_vga1_Mcompar__n0029_inst_cy_378/LOGIC_ZERO ;
  wire \vga_top_vga1_Mcompar__n0029_inst_cy_378/CYINIT ;
  wire \DM_addr_eff<4>/OFF/RST ;
  wire vga_top_vga1_Mcompar__n0029_inst_lut4_53;
  wire \vga_top_vga1__n0029/CYMUXG ;
  wire vga_top_vga1_Mcompar__n0029_inst_lut2_275;
  wire vga_top_vga1_Mcompar__n0029_inst_cy_379;
  wire \vga_top_vga1__n0029/LOGIC_ZERO ;
  wire \vga_top_vga1__n0029/CYINIT ;
  wire vga_top_vga1_Mcompar__n0037_inst_lut2_341;
  wire \vga_top_vga1_Mcompar__n0037_inst_cy_475/CYMUXG ;
  wire vga_top_vga1_Mcompar__n0037_inst_lut2_342;
  wire vga_top_vga1_Mcompar__n0037_inst_cy_474;
  wire \vga_top_vga1_Mcompar__n0037_inst_cy_475/LOGIC_ZERO ;
  wire \vga_top_vga1_Mcompar__n0037_inst_cy_475/LOGIC_ONE ;
  wire vga_top_vga1_Mcompar__n0037_inst_lut4_86;
  wire \vga_top_vga1_Mcompar__n0037_inst_cy_477/CYMUXG ;
  wire vga_top_vga1_Mcompar__n0037_inst_lut4_87;
  wire vga_top_vga1_Mcompar__n0037_inst_cy_476;
  wire \vga_top_vga1_Mcompar__n0037_inst_cy_477/LOGIC_ONE ;
  wire \vga_top_vga1_Mcompar__n0037_inst_cy_477/CYINIT ;
  wire vga_top_vga1_Mcompar__n0037_inst_lut4_88;
  wire \vga_top_vga1__n0037/CYMUXG ;
  wire vga_top_vga1_Mcompar__n0037_inst_lut2_343;
  wire vga_top_vga1_Mcompar__n0037_inst_cy_478;
  wire \vga_top_vga1__n0037/LOGIC_ONE ;
  wire \vga_top_vga1__n0037/CYINIT ;
  wire DLX_EXinst_Mcompar__n0055_inst_lut4_16;
  wire \DLX_EXinst_Mcompar__n0055_inst_cy_119/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0055_inst_lut4_17;
  wire DLX_EXinst_Mcompar__n0055_inst_cy_118;
  wire \DLX_EXinst_Mcompar__n0055_inst_cy_119/LOGIC_ONE ;
  wire \DLX_EXinst_Mcompar__n0055_inst_cy_119/LOGIC_ZERO ;
  wire DLX_EXinst_Mcompar__n0055_inst_lut4_18;
  wire \DLX_EXinst_Mcompar__n0055_inst_cy_121/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0055_inst_lut4_19;
  wire DLX_EXinst_Mcompar__n0055_inst_cy_120;
  wire \DLX_EXinst_Mcompar__n0055_inst_cy_121/LOGIC_ONE ;
  wire \DLX_EXinst_Mcompar__n0055_inst_cy_121/CYINIT ;
  wire DLX_EXinst_Mcompar__n0055_inst_lut4_20;
  wire \DLX_EXinst_Mcompar__n0055_inst_cy_123/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0055_inst_lut4_21;
  wire DLX_EXinst_Mcompar__n0055_inst_cy_122;
  wire \DLX_EXinst_Mcompar__n0055_inst_cy_123/LOGIC_ONE ;
  wire \DLX_EXinst_Mcompar__n0055_inst_cy_123/CYINIT ;
  wire DLX_EXinst_Mcompar__n0055_inst_lut4_22;
  wire \DLX_EXinst_Mcompar__n0055_inst_cy_125/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0055_inst_lut4_23;
  wire DLX_EXinst_Mcompar__n0055_inst_cy_124;
  wire \DLX_EXinst_Mcompar__n0055_inst_cy_125/LOGIC_ONE ;
  wire \DLX_EXinst_Mcompar__n0055_inst_cy_125/CYINIT ;
  wire DLX_EXinst_Mcompar__n0055_inst_lut4_24;
  wire \DLX_EXinst_Mcompar__n0055_inst_cy_127/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0055_inst_lut4_25;
  wire DLX_EXinst_Mcompar__n0055_inst_cy_126;
  wire \DLX_EXinst_Mcompar__n0055_inst_cy_127/LOGIC_ONE ;
  wire \DLX_EXinst_Mcompar__n0055_inst_cy_127/CYINIT ;
  wire DLX_EXinst_Mcompar__n0055_inst_lut4_26;
  wire \DLX_EXinst_Mcompar__n0055_inst_cy_129/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0055_inst_lut4_27;
  wire DLX_EXinst_Mcompar__n0055_inst_cy_128;
  wire \DLX_EXinst_Mcompar__n0055_inst_cy_129/LOGIC_ONE ;
  wire \DLX_EXinst_Mcompar__n0055_inst_cy_129/CYINIT ;
  wire DLX_EXinst_Mcompar__n0055_inst_lut4_28;
  wire \DLX_EXinst_Mcompar__n0055_inst_cy_131/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0055_inst_lut4_29;
  wire DLX_EXinst_Mcompar__n0055_inst_cy_130;
  wire \DLX_EXinst_Mcompar__n0055_inst_cy_131/LOGIC_ONE ;
  wire \DLX_EXinst_Mcompar__n0055_inst_cy_131/CYINIT ;
  wire DLX_EXinst_Mcompar__n0055_inst_lut4_30;
  wire \DLX_EXinst__n0055/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0055_inst_lut4_31;
  wire DLX_EXinst_Mcompar__n0055_inst_cy_132;
  wire \DLX_EXinst__n0055/LOGIC_ONE ;
  wire \DLX_EXinst__n0055/CYINIT ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_166;
  wire \DLX_EXinst_Mcompar__n0063_inst_cy_231/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_167;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_230;
  wire \DLX_EXinst_Mcompar__n0063_inst_cy_231/LOGIC_ZERO ;
  wire \vga_address<9>/FROM ;
  wire \vga_address<9>/XORF ;
  wire \vga_address<9>/CYMUXG ;
  wire \vga_address<9>/LOGIC_ZERO ;
  wire \vga_address<9>/XORG ;
  wire \vga_address<9>/GROM ;
  wire vga_top_vga1_Madd_addressout_inst_cy_469;
  wire \vga_address<9>/CYINIT ;
  wire \vga_address<11>/FROM ;
  wire \vga_address<11>/XORF ;
  wire \vga_address<11>/CYMUXG ;
  wire \vga_address<11>/LOGIC_ZERO ;
  wire \vga_address<11>/XORG ;
  wire \vga_address<11>/GROM ;
  wire vga_top_vga1_Madd_addressout_inst_cy_471;
  wire \vga_address<11>/CYINIT ;
  wire \NPC_eff<1>/OFF/RST ;
  wire \vga_address<13>/LOGIC_ZERO ;
  wire \vga_address<13>/FROM ;
  wire \vga_address<13>/XORF ;
  wire \vga_address<13>/XORG ;
  wire vga_top_vga1_Mmult__n0043_inst_lut2_323_rt;
  wire vga_top_vga1_Madd_addressout_inst_cy_473;
  wire \vga_address<13>/CYINIT ;
  wire DLX_EXinst_Mcompar__n0057_inst_lut2_70;
  wire \DLX_EXinst_Mcompar__n0057_inst_cy_135/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0057_inst_lut2_71;
  wire DLX_EXinst_Mcompar__n0057_inst_cy_134;
  wire \DLX_EXinst_Mcompar__n0057_inst_cy_135/LOGIC_ZERO ;
  wire DLX_EXinst_Mcompar__n0057_inst_lut2_72;
  wire \DLX_EXinst_Mcompar__n0057_inst_cy_137/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0057_inst_lut2_73;
  wire DLX_EXinst_Mcompar__n0057_inst_cy_136;
  wire \DLX_EXinst_Mcompar__n0057_inst_cy_137/CYINIT ;
  wire DLX_EXinst_Mcompar__n0057_inst_lut2_74;
  wire \DLX_EXinst_Mcompar__n0057_inst_cy_139/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0057_inst_lut2_75;
  wire DLX_EXinst_Mcompar__n0057_inst_cy_138;
  wire \DLX_EXinst_Mcompar__n0057_inst_cy_139/CYINIT ;
  wire DLX_EXinst_Mcompar__n0057_inst_lut2_76;
  wire \DLX_EXinst_Mcompar__n0057_inst_cy_141/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0057_inst_lut2_77;
  wire DLX_EXinst_Mcompar__n0057_inst_cy_140;
  wire \DLX_EXinst_Mcompar__n0057_inst_cy_141/CYINIT ;
  wire DLX_EXinst_Mcompar__n0057_inst_lut2_78;
  wire \DLX_EXinst_Mcompar__n0057_inst_cy_143/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0057_inst_lut2_79;
  wire DLX_EXinst_Mcompar__n0057_inst_cy_142;
  wire \DLX_EXinst_Mcompar__n0057_inst_cy_143/CYINIT ;
  wire DLX_EXinst_Mcompar__n0057_inst_lut2_80;
  wire \DLX_EXinst_Mcompar__n0057_inst_cy_145/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0057_inst_lut2_81;
  wire DLX_EXinst_Mcompar__n0057_inst_cy_144;
  wire \DLX_EXinst_Mcompar__n0057_inst_cy_145/CYINIT ;
  wire DLX_EXinst_Mcompar__n0057_inst_lut2_82;
  wire \DLX_EXinst_Mcompar__n0057_inst_cy_147/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0057_inst_lut2_83;
  wire DLX_EXinst_Mcompar__n0057_inst_cy_146;
  wire \DLX_EXinst_Mcompar__n0057_inst_cy_147/CYINIT ;
  wire DLX_EXinst_Mcompar__n0057_inst_lut2_84;
  wire \DLX_EXinst_Mcompar__n0057_inst_cy_149/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0057_inst_lut2_85;
  wire DLX_EXinst_Mcompar__n0057_inst_cy_148;
  wire \DLX_EXinst_Mcompar__n0057_inst_cy_149/CYINIT ;
  wire DLX_EXinst_Mcompar__n0057_inst_lut2_86;
  wire \DLX_EXinst_Mcompar__n0057_inst_cy_151/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0057_inst_lut2_87;
  wire DLX_EXinst_Mcompar__n0057_inst_cy_150;
  wire \DLX_EXinst_Mcompar__n0057_inst_cy_151/CYINIT ;
  wire DLX_EXinst_Mcompar__n0057_inst_lut2_88;
  wire \DLX_EXinst_Mcompar__n0057_inst_cy_153/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0057_inst_lut2_89;
  wire DLX_EXinst_Mcompar__n0057_inst_cy_152;
  wire \DLX_EXinst_Mcompar__n0057_inst_cy_153/CYINIT ;
  wire DLX_EXinst_Mcompar__n0057_inst_lut2_90;
  wire \DLX_EXinst_Mcompar__n0057_inst_cy_155/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0057_inst_lut2_91;
  wire DLX_EXinst_Mcompar__n0057_inst_cy_154;
  wire \DLX_EXinst_Mcompar__n0057_inst_cy_155/CYINIT ;
  wire DLX_EXinst_Mcompar__n0057_inst_lut2_92;
  wire \DLX_EXinst_Mcompar__n0057_inst_cy_157/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0057_inst_lut2_93;
  wire DLX_EXinst_Mcompar__n0057_inst_cy_156;
  wire \DLX_EXinst_Mcompar__n0057_inst_cy_157/CYINIT ;
  wire DLX_EXinst_Mcompar__n0057_inst_lut2_94;
  wire \DLX_EXinst_Mcompar__n0057_inst_cy_159/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0057_inst_lut2_95;
  wire DLX_EXinst_Mcompar__n0057_inst_cy_158;
  wire \DLX_EXinst_Mcompar__n0057_inst_cy_159/CYINIT ;
  wire DLX_EXinst_Mcompar__n0057_inst_lut2_96;
  wire \DLX_EXinst_Mcompar__n0057_inst_cy_161/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0057_inst_lut2_97;
  wire DLX_EXinst_Mcompar__n0057_inst_cy_160;
  wire \DLX_EXinst_Mcompar__n0057_inst_cy_161/CYINIT ;
  wire DLX_EXinst_Mcompar__n0057_inst_lut2_98;
  wire \DLX_EXinst_Mcompar__n0057_inst_cy_163/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0057_inst_lut2_99;
  wire DLX_EXinst_Mcompar__n0057_inst_cy_162;
  wire \DLX_EXinst_Mcompar__n0057_inst_cy_163/CYINIT ;
  wire DLX_EXinst_Mcompar__n0057_inst_lut2_100;
  wire \CHOICE5306/CYMUXF ;
  wire \CHOICE5306/GROM ;
  wire \CHOICE5306/CYINIT ;
  wire \NPC_eff<2>/OFF/RST ;
  wire DLX_IDinst_Mcompar__n0000_inst_lut4_43;
  wire \DLX_IDinst_Mcompar__n0000_inst_cy_266/CYMUXG ;
  wire DLX_IDinst_Mcompar__n0000_inst_lut4_44;
  wire DLX_IDinst_Mcompar__n0000_inst_cy_265;
  wire \DLX_IDinst_Mcompar__n0000_inst_cy_266/LOGIC_ONE ;
  wire \DLX_IDinst_Mcompar__n0000_inst_cy_266/LOGIC_ZERO ;
  wire \DLX_IDinst__n0000/LOGIC_ONE ;
  wire DLX_IDinst_Mcompar__n0000_inst_lut4_45;
  wire \DLX_IDinst__n0000/CYMUXF ;
  wire \DLX_IDinst__n0000/CYINIT ;
  wire DLX_IDinst_Mcompar__n0073_inst_lut4_40;
  wire \DLX_IDinst_Mcompar__n0073_inst_cy_263/CYMUXG ;
  wire DLX_IDinst_Mcompar__n0073_inst_lut4_41;
  wire DLX_IDinst_Mcompar__n0073_inst_cy_262;
  wire \DLX_IDinst_Mcompar__n0073_inst_cy_263/LOGIC_ZERO ;
  wire \DLX_IDinst_Mcompar__n0073_inst_cy_263/LOGIC_ONE ;
  wire \DLX_reg_dst_of_MEM<4>/LOGIC_ZERO ;
  wire DLX_IDinst_Mcompar__n0073_inst_lut4_42;
  wire \DLX_reg_dst_of_MEM<4>/CYMUXF ;
  wire \DLX_reg_dst_of_MEM<4>/CYINIT ;
  wire DLX_IDinst_Mcompar__n0314_inst_lut4_40;
  wire \DLX_IDinst_Mcompar__n0314_inst_cy_263/CYMUXG ;
  wire DLX_IDinst_Mcompar__n0314_inst_lut4_41;
  wire DLX_IDinst_Mcompar__n0314_inst_cy_262;
  wire \DLX_IDinst_Mcompar__n0314_inst_cy_263/LOGIC_ZERO ;
  wire \DLX_IDinst_Mcompar__n0314_inst_cy_263/LOGIC_ONE ;
  wire vga_top_vga1_Mmult__n0043_inst_lut2_303;
  wire \vga_top_vga1_Mmult__n0043_inst_lut2_317/CYMUXG ;
  wire \vga_top_vga1_Mmult__n0043_inst_lut2_317/XORG ;
  wire vga_top_vga1_Mmult__n0043_inst_lut2_304;
  wire vga_top_vga1_Mmult__n0043_inst_cy_439;
  wire \vga_top_vga1_Mmult__n0043_inst_lut2_317/LOGIC_ZERO ;
  wire vga_top_vga1_Mmult__n0043_inst_lut2_305;
  wire \vga_top_vga1_Mmult__n0043_inst_lut2_318/XORF ;
  wire \vga_top_vga1_Mmult__n0043_inst_lut2_318/CYMUXG ;
  wire \vga_top_vga1_Mmult__n0043_inst_lut2_318/XORG ;
  wire vga_top_vga1_Mmult__n0043_inst_lut2_306;
  wire vga_top_vga1_Mmult__n0043_inst_cy_441;
  wire \vga_top_vga1_Mmult__n0043_inst_lut2_318/CYINIT ;
  wire vga_top_vga1_Mmult__n0043_inst_lut2_307;
  wire \vga_top_vga1_Mmult__n0043_inst_lut2_320/XORF ;
  wire \vga_top_vga1_Mmult__n0043_inst_lut2_320/CYMUXG ;
  wire \vga_top_vga1_Mmult__n0043_inst_lut2_320/XORG ;
  wire vga_top_vga1_Mmult__n0043_inst_lut2_308;
  wire vga_top_vga1_Mmult__n0043_inst_cy_443;
  wire \vga_top_vga1_Mmult__n0043_inst_lut2_320/CYINIT ;
  wire vga_top_vga1_Mmult__n0043_inst_lut2_309;
  wire \vga_top_vga1_Mmult__n0043_inst_lut2_322/XORF ;
  wire \vga_top_vga1_Mmult__n0043_inst_lut2_322/XORG ;
  wire \vga_top_vga1_gridvcounter<7>_rt ;
  wire vga_top_vga1_Mmult__n0043_inst_cy_445;
  wire \vga_top_vga1_Mmult__n0043_inst_lut2_322/CYINIT ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_102;
  wire \DLX_EXinst_Mcompar__n0091_inst_cy_167/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_103;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_166;
  wire \DLX_EXinst_Mcompar__n0091_inst_cy_167/LOGIC_ZERO ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_104;
  wire \DLX_EXinst_Mcompar__n0091_inst_cy_169/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_105;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_168;
  wire \DLX_EXinst_Mcompar__n0091_inst_cy_169/CYINIT ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_106;
  wire \DLX_EXinst_Mcompar__n0091_inst_cy_171/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_107;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_170;
  wire \DLX_EXinst_Mcompar__n0091_inst_cy_171/CYINIT ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_108;
  wire \DLX_EXinst_Mcompar__n0091_inst_cy_173/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_109;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_172;
  wire \DLX_EXinst_Mcompar__n0091_inst_cy_173/CYINIT ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_110;
  wire \DLX_EXinst_Mcompar__n0091_inst_cy_175/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_111;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_174;
  wire \DLX_EXinst_Mcompar__n0091_inst_cy_175/CYINIT ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_112;
  wire \DLX_EXinst_Mcompar__n0091_inst_cy_177/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_113;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_176;
  wire \DLX_EXinst_Mcompar__n0091_inst_cy_177/CYINIT ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_114;
  wire \DLX_EXinst_Mcompar__n0091_inst_cy_179/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_115;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_178;
  wire \DLX_EXinst_Mcompar__n0091_inst_cy_179/CYINIT ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_116;
  wire \DLX_EXinst_Mcompar__n0091_inst_cy_181/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_117;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_180;
  wire \DLX_EXinst_Mcompar__n0091_inst_cy_181/CYINIT ;
  wire \NPC_eff<3>/OFF/RST ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_118;
  wire \DLX_EXinst_Mcompar__n0091_inst_cy_183/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_119;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_182;
  wire \DLX_EXinst_Mcompar__n0091_inst_cy_183/CYINIT ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_120;
  wire \DLX_EXinst_Mcompar__n0091_inst_cy_185/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_121;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_184;
  wire \DLX_EXinst_Mcompar__n0091_inst_cy_185/CYINIT ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_122;
  wire \DLX_EXinst_Mcompar__n0091_inst_cy_187/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_123;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_186;
  wire \DLX_EXinst_Mcompar__n0091_inst_cy_187/CYINIT ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_124;
  wire \DLX_EXinst_Mcompar__n0091_inst_cy_189/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_125;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_188;
  wire \DLX_EXinst_Mcompar__n0091_inst_cy_189/CYINIT ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_126;
  wire \DLX_EXinst_Mcompar__n0091_inst_cy_191/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_127;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_190;
  wire \DLX_EXinst_Mcompar__n0091_inst_cy_191/CYINIT ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_128;
  wire \DLX_EXinst_Mcompar__n0091_inst_cy_193/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_129;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_192;
  wire \DLX_EXinst_Mcompar__n0091_inst_cy_193/CYINIT ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_130;
  wire \DLX_EXinst_Mcompar__n0091_inst_cy_195/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_131;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_194;
  wire \DLX_EXinst_Mcompar__n0091_inst_cy_195/CYINIT ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_132;
  wire \N127408/CYMUXF ;
  wire \N127408/GROM ;
  wire \N127408/CYINIT ;
  wire DLX_EXinst_Mcompar__n0059_inst_lut2_102;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_167/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0059_inst_lut2_103;
  wire DLX_EXinst_Mcompar__n0059_inst_cy_166;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_167/LOGIC_ZERO ;
  wire DLX_EXinst_Mcompar__n0059_inst_lut2_104;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_169/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0059_inst_lut2_105;
  wire DLX_EXinst_Mcompar__n0059_inst_cy_168;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_169/CYINIT ;
  wire DLX_EXinst_Mcompar__n0059_inst_lut2_106;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_171/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0059_inst_lut2_107;
  wire DLX_EXinst_Mcompar__n0059_inst_cy_170;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_171/CYINIT ;
  wire DLX_EXinst_Mcompar__n0059_inst_lut2_108;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_173/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0059_inst_lut2_109;
  wire DLX_EXinst_Mcompar__n0059_inst_cy_172;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_173/CYINIT ;
  wire DLX_EXinst_Mcompar__n0059_inst_lut2_110;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_175/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0059_inst_lut2_111;
  wire DLX_EXinst_Mcompar__n0059_inst_cy_174;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_175/CYINIT ;
  wire DLX_EXinst_Mcompar__n0059_inst_lut2_112;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_177/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0059_inst_lut2_113;
  wire DLX_EXinst_Mcompar__n0059_inst_cy_176;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_177/CYINIT ;
  wire DLX_EXinst_Mcompar__n0059_inst_lut2_114;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_179/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0059_inst_lut2_115;
  wire DLX_EXinst_Mcompar__n0059_inst_cy_178;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_179/CYINIT ;
  wire DLX_EXinst_Mcompar__n0059_inst_lut2_116;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_181/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0059_inst_lut2_117;
  wire DLX_EXinst_Mcompar__n0059_inst_cy_180;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_181/CYINIT ;
  wire DLX_EXinst_Mcompar__n0059_inst_lut2_118;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_183/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0059_inst_lut2_119;
  wire DLX_EXinst_Mcompar__n0059_inst_cy_182;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_183/CYINIT ;
  wire DLX_EXinst_Mcompar__n0059_inst_lut2_120;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_185/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0059_inst_lut2_121;
  wire DLX_EXinst_Mcompar__n0059_inst_cy_184;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_185/CYINIT ;
  wire DLX_EXinst_Mcompar__n0059_inst_lut2_122;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_187/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0059_inst_lut2_123;
  wire DLX_EXinst_Mcompar__n0059_inst_cy_186;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_187/CYINIT ;
  wire DLX_EXinst_Mcompar__n0059_inst_lut2_124;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_189/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0059_inst_lut2_125;
  wire DLX_EXinst_Mcompar__n0059_inst_cy_188;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_189/CYINIT ;
  wire DLX_EXinst_Mcompar__n0059_inst_lut2_126;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_191/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0059_inst_lut2_127;
  wire DLX_EXinst_Mcompar__n0059_inst_cy_190;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_191/CYINIT ;
  wire DLX_EXinst_Mcompar__n0059_inst_lut2_128;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_193/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0059_inst_lut2_129;
  wire DLX_EXinst_Mcompar__n0059_inst_cy_192;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_193/CYINIT ;
  wire \NPC_eff<4>/OFF/RST ;
  wire DLX_EXinst_Mcompar__n0059_inst_lut2_130;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_195/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0059_inst_lut2_131;
  wire DLX_EXinst_Mcompar__n0059_inst_cy_194;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_195/CYINIT ;
  wire DLX_EXinst_Mcompar__n0059_inst_lut2_132;
  wire \CHOICE5313/CYMUXF ;
  wire \CHOICE5313/GROM ;
  wire \CHOICE5313/CYINIT ;
  wire DLX_IDinst_Mcompar__n0075_inst_lut4_40;
  wire \DLX_IDinst_Mcompar__n0075_inst_cy_263/CYMUXG ;
  wire DLX_IDinst_Mcompar__n0075_inst_lut4_41;
  wire DLX_IDinst_Mcompar__n0075_inst_cy_262;
  wire \DLX_IDinst_Mcompar__n0075_inst_cy_263/LOGIC_ZERO ;
  wire \DLX_IDinst_Mcompar__n0075_inst_cy_263/LOGIC_ONE ;
  wire \DLX_EXinst_reg_dst_out<4>/LOGIC_ZERO ;
  wire DLX_IDinst_Mcompar__n0075_inst_lut4_42;
  wire \DLX_EXinst_reg_dst_out<4>/CYMUXF ;
  wire \DLX_EXinst_reg_dst_out<4>/CYINIT ;
  wire DLX_IDinst_Mcompar__n0315_inst_lut4_40;
  wire \DLX_IDinst_Mcompar__n0315_inst_cy_263/CYMUXG ;
  wire DLX_IDinst_Mcompar__n0315_inst_lut4_41;
  wire DLX_IDinst_Mcompar__n0315_inst_cy_262;
  wire \DLX_IDinst_Mcompar__n0315_inst_cy_263/LOGIC_ZERO ;
  wire \DLX_IDinst_Mcompar__n0315_inst_cy_263/LOGIC_ONE ;
  wire \DLX_IDinst_Madd__n0129_inst_lut2_198/FROM ;
  wire \DLX_IDinst_Madd__n0129_inst_lut2_198/CYMUXG ;
  wire \DLX_IDinst_Madd__n0129_inst_lut2_198/XORG ;
  wire DLX_IDinst_Madd__n0129_inst_lut2_199;
  wire DLX_IDinst_Madd__n0129_inst_cy_268;
  wire \DLX_IDinst_Madd__n0129_inst_lut2_198/LOGIC_ZERO ;
  wire DLX_IDinst_Madd__n0129_inst_lut2_200;
  wire \DLX_IDinst__n0129<2>/XORF ;
  wire \DLX_IDinst__n0129<2>/CYMUXG ;
  wire \DLX_IDinst__n0129<2>/XORG ;
  wire DLX_IDinst_Madd__n0129_inst_lut2_201;
  wire DLX_IDinst_Madd__n0129_inst_cy_270;
  wire \DLX_IDinst__n0129<2>/CYINIT ;
  wire DLX_IDinst_Madd__n0129_inst_lut2_202;
  wire \DLX_IDinst__n0129<4>/XORF ;
  wire \DLX_IDinst__n0129<4>/CYMUXG ;
  wire \DLX_IDinst__n0129<4>/XORG ;
  wire DLX_IDinst_Madd__n0129_inst_lut2_203;
  wire DLX_IDinst_Madd__n0129_inst_cy_272;
  wire \DLX_IDinst__n0129<4>/CYINIT ;
  wire DLX_IDinst_Madd__n0129_inst_lut2_204;
  wire \DLX_IDinst__n0129<6>/XORF ;
  wire \DLX_IDinst__n0129<6>/CYMUXG ;
  wire \DLX_IDinst__n0129<6>/XORG ;
  wire DLX_IDinst_Madd__n0129_inst_lut2_205;
  wire DLX_IDinst_Madd__n0129_inst_cy_274;
  wire \DLX_IDinst__n0129<6>/CYINIT ;
  wire DLX_IDinst_Madd__n0129_inst_lut2_206;
  wire \DLX_IDinst__n0129<8>/XORF ;
  wire \DLX_IDinst__n0129<8>/CYMUXG ;
  wire \DLX_IDinst__n0129<8>/XORG ;
  wire DLX_IDinst_Madd__n0129_inst_lut2_207;
  wire DLX_IDinst_Madd__n0129_inst_cy_276;
  wire \DLX_IDinst__n0129<8>/CYINIT ;
  wire DLX_IDinst_Madd__n0129_inst_lut2_208;
  wire \DLX_IDinst__n0129<10>/XORF ;
  wire \DLX_IDinst__n0129<10>/CYMUXG ;
  wire \DLX_IDinst__n0129<10>/XORG ;
  wire DLX_IDinst_Madd__n0129_inst_lut2_209;
  wire DLX_IDinst_Madd__n0129_inst_cy_278;
  wire \DLX_IDinst__n0129<10>/CYINIT ;
  wire DLX_IDinst_Madd__n0129_inst_lut2_210;
  wire \DLX_IDinst__n0129<12>/XORF ;
  wire \DLX_IDinst__n0129<12>/CYMUXG ;
  wire \DLX_IDinst__n0129<12>/XORG ;
  wire DLX_IDinst_Madd__n0129_inst_lut2_211;
  wire DLX_IDinst_Madd__n0129_inst_cy_280;
  wire \DLX_IDinst__n0129<12>/CYINIT ;
  wire \NPC_eff<5>/OFF/RST ;
  wire DLX_IDinst_Madd__n0129_inst_lut2_212;
  wire \DLX_IDinst__n0129<14>/XORF ;
  wire \DLX_IDinst__n0129<14>/CYMUXG ;
  wire \DLX_IDinst__n0129<14>/XORG ;
  wire DLX_IDinst_Madd__n0129_inst_lut2_213;
  wire DLX_IDinst_Madd__n0129_inst_cy_282;
  wire \DLX_IDinst__n0129<14>/CYINIT ;
  wire DLX_IDinst_Madd__n0129_inst_lut2_214;
  wire \DLX_IDinst__n0129<16>/XORF ;
  wire \DLX_IDinst__n0129<16>/CYMUXG ;
  wire \DLX_IDinst__n0129<16>/XORG ;
  wire DLX_IDinst_Madd__n0129_inst_lut2_215;
  wire DLX_IDinst_Madd__n0129_inst_cy_284;
  wire \DLX_IDinst__n0129<16>/CYINIT ;
  wire DLX_IDinst_Madd__n0129_inst_lut2_216;
  wire \DLX_IDinst__n0129<18>/XORF ;
  wire \DLX_IDinst__n0129<18>/CYMUXG ;
  wire \DLX_IDinst__n0129<18>/XORG ;
  wire DLX_IDinst_Madd__n0129_inst_lut2_217;
  wire DLX_IDinst_Madd__n0129_inst_cy_286;
  wire \DLX_IDinst__n0129<18>/CYINIT ;
  wire DLX_IDinst_Madd__n0129_inst_lut2_218;
  wire \DLX_IDinst__n0129<20>/XORF ;
  wire \DLX_IDinst__n0129<20>/CYMUXG ;
  wire \DLX_IDinst__n0129<20>/XORG ;
  wire DLX_IDinst_Madd__n0129_inst_lut2_219;
  wire DLX_IDinst_Madd__n0129_inst_cy_288;
  wire \DLX_IDinst__n0129<20>/CYINIT ;
  wire DLX_IDinst_Madd__n0129_inst_lut2_220;
  wire \DLX_IDinst__n0129<22>/XORF ;
  wire \DLX_IDinst__n0129<22>/CYMUXG ;
  wire \DLX_IDinst__n0129<22>/XORG ;
  wire DLX_IDinst_Madd__n0129_inst_lut2_221;
  wire DLX_IDinst_Madd__n0129_inst_cy_290;
  wire \DLX_IDinst__n0129<22>/CYINIT ;
  wire DLX_IDinst_Madd__n0129_inst_lut2_222;
  wire \DLX_IDinst__n0129<24>/XORF ;
  wire \DLX_IDinst__n0129<24>/CYMUXG ;
  wire \DLX_IDinst__n0129<24>/XORG ;
  wire DLX_IDinst_Madd__n0129_inst_lut2_223;
  wire DLX_IDinst_Madd__n0129_inst_cy_292;
  wire \DLX_IDinst__n0129<24>/CYINIT ;
  wire DLX_IDinst_Madd__n0129_inst_lut2_224;
  wire \DLX_IDinst__n0129<26>/XORF ;
  wire \DLX_IDinst__n0129<26>/CYMUXG ;
  wire \DLX_IDinst__n0129<26>/XORG ;
  wire DLX_IDinst_Madd__n0129_inst_lut2_225;
  wire DLX_IDinst_Madd__n0129_inst_cy_294;
  wire \DLX_IDinst__n0129<26>/CYINIT ;
  wire DLX_IDinst_Madd__n0129_inst_lut2_226;
  wire \DLX_IDinst__n0129<28>/XORF ;
  wire \DLX_IDinst__n0129<28>/CYMUXG ;
  wire \DLX_IDinst__n0129<28>/XORG ;
  wire DLX_IDinst_Madd__n0129_inst_lut2_227;
  wire DLX_IDinst_Madd__n0129_inst_cy_296;
  wire \DLX_IDinst__n0129<28>/CYINIT ;
  wire DLX_IDinst_Madd__n0129_inst_lut2_228;
  wire \DLX_IDinst__n0129<30>/XORF ;
  wire \DLX_IDinst__n0129<30>/XORG ;
  wire DLX_IDinst_Madd__n0129_inst_lut2_229;
  wire DLX_IDinst_Madd__n0129_inst_cy_298;
  wire \DLX_IDinst__n0129<30>/CYINIT ;
  wire DLX_IDinst_Mcompar__n0003_inst_lut4_43;
  wire \DLX_IDinst_Mcompar__n0003_inst_cy_266/CYMUXG ;
  wire DLX_IDinst_Mcompar__n0003_inst_lut4_44;
  wire DLX_IDinst_Mcompar__n0003_inst_cy_265;
  wire \DLX_IDinst_Mcompar__n0003_inst_cy_266/LOGIC_ONE ;
  wire \DLX_IDinst_Mcompar__n0003_inst_cy_266/LOGIC_ZERO ;
  wire \DLX_IDinst_rt_addr<4>/FFY/RST ;
  wire \DLX_IDinst_rt_addr<4>/LOGIC_ONE ;
  wire DLX_IDinst_Mcompar__n0003_inst_lut4_45;
  wire \DLX_IDinst_rt_addr<4>/CYMUXF ;
  wire \DLX_IDinst_rt_addr<4>/CYINIT ;
  wire vga_top_vga1_vcounter_Madd__n0000_inst_lut2_9;
  wire \vga_top_vga1_vcounter<0>/CYMUXG ;
  wire \vga_top_vga1_vcounter<0>/GROM ;
  wire vga_top_vga1_vcounter_Madd__n0000_inst_cy_9;
  wire \vga_top_vga1_vcounter<0>/LOGIC_ZERO ;
  wire \vga_top_vga1_vcounter<2>/FROM ;
  wire \vga_top_vga1_vcounter<2>/CYMUXG ;
  wire \vga_top_vga1_vcounter<2>/LOGIC_ZERO ;
  wire \vga_top_vga1_vcounter<2>/GROM ;
  wire vga_top_vga1_vcounter_Madd__n0000_inst_cy_11;
  wire \vga_top_vga1_vcounter<2>/CYINIT ;
  wire \vga_top_vga1_vcounter<4>/FROM ;
  wire \vga_top_vga1_vcounter<4>/CYMUXG ;
  wire \vga_top_vga1_vcounter<4>/LOGIC_ZERO ;
  wire \vga_top_vga1_vcounter<4>/GROM ;
  wire vga_top_vga1_vcounter_Madd__n0000_inst_cy_13;
  wire \vga_top_vga1_vcounter<4>/CYINIT ;
  wire \vga_top_vga1_vcounter<6>/FROM ;
  wire \vga_top_vga1_vcounter<6>/CYMUXG ;
  wire \vga_top_vga1_vcounter<6>/LOGIC_ZERO ;
  wire \vga_top_vga1_vcounter<6>/GROM ;
  wire vga_top_vga1_vcounter_Madd__n0000_inst_cy_15;
  wire \vga_top_vga1_vcounter<6>/CYINIT ;
  wire \vga_top_vga1_vcounter<8>/LOGIC_ZERO ;
  wire \vga_top_vga1_vcounter<8>/FROM ;
  wire \vga_top_vga1_vcounter<9>_rt ;
  wire vga_top_vga1_vcounter_Madd__n0000_inst_cy_17;
  wire \vga_top_vga1_vcounter<8>/CYINIT ;
  wire vga_top_vga1_hcounter_Madd__n0000_inst_lut2_19;
  wire \vga_top_vga1_hcounter<0>/CYMUXG ;
  wire \vga_top_vga1_hcounter<0>/GROM ;
  wire vga_top_vga1_hcounter_Madd__n0000_inst_cy_19;
  wire \vga_top_vga1_hcounter<0>/LOGIC_ZERO ;
  wire \vga_top_vga1_hcounter<2>/FROM ;
  wire \vga_top_vga1_hcounter<2>/CYMUXG ;
  wire \vga_top_vga1_hcounter<2>/LOGIC_ZERO ;
  wire \vga_top_vga1_hcounter<2>/GROM ;
  wire vga_top_vga1_hcounter_Madd__n0000_inst_cy_21;
  wire \vga_top_vga1_hcounter<2>/CYINIT ;
  wire \vga_top_vga1_hcounter<4>/FROM ;
  wire \vga_top_vga1_hcounter<4>/CYMUXG ;
  wire \vga_top_vga1_hcounter<4>/LOGIC_ZERO ;
  wire \vga_top_vga1_hcounter<4>/GROM ;
  wire vga_top_vga1_hcounter_Madd__n0000_inst_cy_23;
  wire \vga_top_vga1_hcounter<4>/CYINIT ;
  wire \vga_top_vga1_hcounter<6>/FROM ;
  wire \vga_top_vga1_hcounter<6>/CYMUXG ;
  wire \vga_top_vga1_hcounter<6>/LOGIC_ZERO ;
  wire \vga_top_vga1_hcounter<6>/GROM ;
  wire vga_top_vga1_hcounter_Madd__n0000_inst_cy_25;
  wire \vga_top_vga1_hcounter<6>/CYINIT ;
  wire \vga_top_vga1_hcounter<8>/FROM ;
  wire \vga_top_vga1_hcounter<8>/CYMUXG ;
  wire \vga_top_vga1_hcounter<8>/LOGIC_ZERO ;
  wire \vga_top_vga1_hcounter<8>/GROM ;
  wire vga_top_vga1_hcounter_Madd__n0000_inst_cy_27;
  wire \vga_top_vga1_hcounter<8>/CYINIT ;
  wire \vga_top_vga1_hcounter<10>/FROM ;
  wire \vga_top_vga1_hcounter<10>/CYMUXG ;
  wire \vga_top_vga1_hcounter<10>/LOGIC_ZERO ;
  wire \vga_top_vga1_hcounter<10>/GROM ;
  wire vga_top_vga1_hcounter_Madd__n0000_inst_cy_29;
  wire \vga_top_vga1_hcounter<10>/CYINIT ;
  wire \vga_top_vga1_hcounter<12>/FROM ;
  wire \vga_top_vga1_hcounter<12>/CYMUXG ;
  wire \vga_top_vga1_hcounter<12>/LOGIC_ZERO ;
  wire \vga_top_vga1_hcounter<12>/GROM ;
  wire vga_top_vga1_hcounter_Madd__n0000_inst_cy_31;
  wire \vga_top_vga1_hcounter<12>/CYINIT ;
  wire \vga_top_vga1_hcounter<14>/LOGIC_ZERO ;
  wire \vga_top_vga1_hcounter<14>/FROM ;
  wire \vga_top_vga1_hcounter<15>_rt ;
  wire vga_top_vga1_hcounter_Madd__n0000_inst_cy_33;
  wire \vga_top_vga1_hcounter<14>/CYINIT ;
  wire DLX_EXinst_Mcompar__n0085_inst_lut4_0;
  wire \DLX_EXinst_Mcompar__n0085_inst_cy_103/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0085_inst_lut4_1;
  wire DLX_EXinst_Mcompar__n0085_inst_cy_102;
  wire \DLX_EXinst_Mcompar__n0085_inst_cy_103/LOGIC_ZERO ;
  wire \DLX_EXinst_Mcompar__n0085_inst_cy_103/LOGIC_ONE ;
  wire DLX_EXinst_Mcompar__n0085_inst_lut4_2;
  wire \DLX_EXinst_Mcompar__n0085_inst_cy_105/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0085_inst_lut4_3;
  wire DLX_EXinst_Mcompar__n0085_inst_cy_104;
  wire \DLX_EXinst_Mcompar__n0085_inst_cy_105/LOGIC_ZERO ;
  wire \DLX_EXinst_Mcompar__n0085_inst_cy_105/CYINIT ;
  wire DLX_EXinst_Mcompar__n0085_inst_lut4_4;
  wire \DLX_EXinst_Mcompar__n0085_inst_cy_107/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0085_inst_lut4_5;
  wire DLX_EXinst_Mcompar__n0085_inst_cy_106;
  wire \DLX_EXinst_Mcompar__n0085_inst_cy_107/LOGIC_ZERO ;
  wire \DLX_EXinst_Mcompar__n0085_inst_cy_107/CYINIT ;
  wire \NPC_eff<6>/OFF/RST ;
  wire DLX_EXinst_Mcompar__n0085_inst_lut4_6;
  wire \DLX_EXinst_Mcompar__n0085_inst_cy_109/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0085_inst_lut4_7;
  wire DLX_EXinst_Mcompar__n0085_inst_cy_108;
  wire \DLX_EXinst_Mcompar__n0085_inst_cy_109/LOGIC_ZERO ;
  wire \DLX_EXinst_Mcompar__n0085_inst_cy_109/CYINIT ;
  wire DLX_EXinst_Mcompar__n0085_inst_lut4_8;
  wire \DLX_EXinst_Mcompar__n0085_inst_cy_111/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0085_inst_lut4_9;
  wire DLX_EXinst_Mcompar__n0085_inst_cy_110;
  wire \DLX_EXinst_Mcompar__n0085_inst_cy_111/LOGIC_ZERO ;
  wire \DLX_EXinst_Mcompar__n0085_inst_cy_111/CYINIT ;
  wire DLX_EXinst_Mcompar__n0085_inst_lut4_10;
  wire \DLX_EXinst_Mcompar__n0085_inst_cy_113/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0085_inst_lut4_11;
  wire DLX_EXinst_Mcompar__n0085_inst_cy_112;
  wire \DLX_EXinst_Mcompar__n0085_inst_cy_113/LOGIC_ZERO ;
  wire \DLX_EXinst_Mcompar__n0085_inst_cy_113/CYINIT ;
  wire DLX_EXinst_Mcompar__n0085_inst_lut4_12;
  wire \DLX_EXinst_Mcompar__n0085_inst_cy_115/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0085_inst_lut4_13;
  wire DLX_EXinst_Mcompar__n0085_inst_cy_114;
  wire \DLX_EXinst_Mcompar__n0085_inst_cy_115/LOGIC_ZERO ;
  wire \DLX_EXinst_Mcompar__n0085_inst_cy_115/CYINIT ;
  wire DLX_EXinst_Mcompar__n0085_inst_lut4_14;
  wire \DLX_EXinst__n0085/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0085_inst_lut4_15;
  wire DLX_EXinst_Mcompar__n0085_inst_cy_116;
  wire \DLX_EXinst__n0085/LOGIC_ZERO ;
  wire \DLX_EXinst__n0085/CYINIT ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_134;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_199/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_135;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_198;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_199/LOGIC_ZERO ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_136;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_201/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_137;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_200;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_201/CYINIT ;
  wire \NPC_eff<7>/OFF/RST ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_138;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_203/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_139;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_202;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_203/CYINIT ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_140;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_205/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_141;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_204;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_205/CYINIT ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_142;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_207/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_143;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_206;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_207/CYINIT ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_144;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_209/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_145;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_208;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_209/CYINIT ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_146;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_211/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_147;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_210;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_211/CYINIT ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_148;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_213/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_149;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_212;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_213/CYINIT ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_150;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_215/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_151;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_214;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_215/CYINIT ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_152;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_217/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_153;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_216;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_217/CYINIT ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_154;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_219/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_155;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_218;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_219/CYINIT ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_156;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_221/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_157;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_220;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_221/CYINIT ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_158;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_223/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_159;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_222;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_223/CYINIT ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_160;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_225/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_161;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_224;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_225/CYINIT ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_162;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_227/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_163;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_226;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_227/CYINIT ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_164;
  wire \CHOICE1126/CYMUXF ;
  wire \CHOICE1126/GROM ;
  wire \CHOICE1126/CYINIT ;
  wire DLX_IDinst_Mcompar__n0077_inst_lut4_40;
  wire \DLX_IDinst_Mcompar__n0077_inst_cy_263/CYMUXG ;
  wire DLX_IDinst_Mcompar__n0077_inst_lut4_41;
  wire DLX_IDinst_Mcompar__n0077_inst_cy_262;
  wire \DLX_IDinst_Mcompar__n0077_inst_cy_263/LOGIC_ZERO ;
  wire \DLX_IDinst_Mcompar__n0077_inst_cy_263/LOGIC_ONE ;
  wire \DLX_IDinst__n0077/LOGIC_ZERO ;
  wire DLX_IDinst_Mcompar__n0077_inst_lut4_42;
  wire \DLX_IDinst__n0077/CYMUXF ;
  wire \DLX_IDinst__n0077/CYINIT ;
  wire DLX_EXinst_Maddsub__n0016_inst_lut3_6;
  wire \DLX_EXinst__n0016<0>/XORF ;
  wire \DLX_EXinst__n0016<0>/CYMUXG ;
  wire \DLX_EXinst__n0016<0>/XORG ;
  wire DLX_EXinst_Maddsub__n0016_inst_lut3_7;
  wire DLX_EXinst_Maddsub__n0016_inst_cy_70;
  wire \DLX_EXinst__n0016<0>/CYINIT ;
  wire DLX_EXinst_Maddsub__n0016_inst_lut3_8;
  wire \DLX_EXinst__n0016<2>/XORF ;
  wire \DLX_EXinst__n0016<2>/CYMUXG ;
  wire \DLX_EXinst__n0016<2>/XORG ;
  wire DLX_EXinst_Maddsub__n0016_inst_lut3_9;
  wire DLX_EXinst_Maddsub__n0016_inst_cy_72;
  wire \DLX_EXinst__n0016<2>/CYINIT ;
  wire DLX_EXinst_Maddsub__n0016_inst_lut3_10;
  wire \DLX_EXinst__n0016<4>/XORF ;
  wire \DLX_EXinst__n0016<4>/CYMUXG ;
  wire \DLX_EXinst__n0016<4>/XORG ;
  wire DLX_EXinst_Maddsub__n0016_inst_lut3_11;
  wire DLX_EXinst_Maddsub__n0016_inst_cy_74;
  wire \DLX_EXinst__n0016<4>/CYINIT ;
  wire DLX_EXinst_Maddsub__n0016_inst_lut3_12;
  wire \DLX_EXinst__n0016<6>/XORF ;
  wire \DLX_EXinst__n0016<6>/CYMUXG ;
  wire \DLX_EXinst__n0016<6>/XORG ;
  wire DLX_EXinst_Maddsub__n0016_inst_lut3_13;
  wire DLX_EXinst_Maddsub__n0016_inst_cy_76;
  wire \DLX_EXinst__n0016<6>/CYINIT ;
  wire DLX_EXinst_Maddsub__n0016_inst_lut3_14;
  wire \DLX_EXinst__n0016<8>/XORF ;
  wire \DLX_EXinst__n0016<8>/CYMUXG ;
  wire \DLX_EXinst__n0016<8>/XORG ;
  wire DLX_EXinst_Maddsub__n0016_inst_lut3_15;
  wire DLX_EXinst_Maddsub__n0016_inst_cy_78;
  wire \DLX_EXinst__n0016<8>/CYINIT ;
  wire DLX_EXinst_Maddsub__n0016_inst_lut3_16;
  wire \DLX_EXinst__n0016<10>/XORF ;
  wire \DLX_EXinst__n0016<10>/CYMUXG ;
  wire \DLX_EXinst__n0016<10>/XORG ;
  wire DLX_EXinst_Maddsub__n0016_inst_lut3_17;
  wire DLX_EXinst_Maddsub__n0016_inst_cy_80;
  wire \DLX_EXinst__n0016<10>/CYINIT ;
  wire \NPC_eff<8>/OFF/RST ;
  wire DLX_EXinst_Maddsub__n0016_inst_lut3_18;
  wire \DLX_EXinst__n0016<12>/XORF ;
  wire \DLX_EXinst__n0016<12>/CYMUXG ;
  wire \DLX_EXinst__n0016<12>/XORG ;
  wire DLX_EXinst_Maddsub__n0016_inst_lut3_19;
  wire DLX_EXinst_Maddsub__n0016_inst_cy_82;
  wire \DLX_EXinst__n0016<12>/CYINIT ;
  wire DLX_EXinst_Maddsub__n0016_inst_lut3_20;
  wire \DLX_EXinst__n0016<14>/XORF ;
  wire \DLX_EXinst__n0016<14>/CYMUXG ;
  wire \DLX_EXinst__n0016<14>/XORG ;
  wire DLX_EXinst_Maddsub__n0016_inst_lut3_21;
  wire DLX_EXinst_Maddsub__n0016_inst_cy_84;
  wire \DLX_EXinst__n0016<14>/CYINIT ;
  wire DLX_EXinst_Maddsub__n0016_inst_lut3_22;
  wire \DLX_EXinst__n0016<16>/XORF ;
  wire \DLX_EXinst__n0016<16>/CYMUXG ;
  wire \DLX_EXinst__n0016<16>/XORG ;
  wire DLX_EXinst_Maddsub__n0016_inst_lut3_23;
  wire DLX_EXinst_Maddsub__n0016_inst_cy_86;
  wire \DLX_EXinst__n0016<16>/CYINIT ;
  wire DLX_EXinst_Maddsub__n0016_inst_lut3_24;
  wire \DLX_EXinst__n0016<18>/XORF ;
  wire \DLX_EXinst__n0016<18>/CYMUXG ;
  wire \DLX_EXinst__n0016<18>/XORG ;
  wire DLX_EXinst_Maddsub__n0016_inst_lut3_25;
  wire DLX_EXinst_Maddsub__n0016_inst_cy_88;
  wire \DLX_EXinst__n0016<18>/CYINIT ;
  wire DLX_EXinst_Maddsub__n0016_inst_lut3_26;
  wire \DLX_EXinst__n0016<20>/XORF ;
  wire \DLX_EXinst__n0016<20>/CYMUXG ;
  wire \DLX_EXinst__n0016<20>/XORG ;
  wire DLX_EXinst_Maddsub__n0016_inst_lut3_27;
  wire DLX_EXinst_Maddsub__n0016_inst_cy_90;
  wire \DLX_EXinst__n0016<20>/CYINIT ;
  wire DLX_EXinst_Maddsub__n0016_inst_lut3_28;
  wire \DLX_EXinst__n0016<22>/XORF ;
  wire \DLX_EXinst__n0016<22>/CYMUXG ;
  wire \DLX_EXinst__n0016<22>/XORG ;
  wire DLX_EXinst_Maddsub__n0016_inst_lut3_29;
  wire DLX_EXinst_Maddsub__n0016_inst_cy_92;
  wire \DLX_EXinst__n0016<22>/CYINIT ;
  wire DLX_EXinst_Maddsub__n0016_inst_lut3_30;
  wire \DLX_EXinst__n0016<24>/XORF ;
  wire \DLX_EXinst__n0016<24>/CYMUXG ;
  wire \DLX_EXinst__n0016<24>/XORG ;
  wire DLX_EXinst_Maddsub__n0016_inst_lut3_31;
  wire DLX_EXinst_Maddsub__n0016_inst_cy_94;
  wire \DLX_EXinst__n0016<24>/CYINIT ;
  wire DLX_EXinst_Maddsub__n0016_inst_lut3_32;
  wire \DLX_EXinst__n0016<26>/XORF ;
  wire \DLX_EXinst__n0016<26>/CYMUXG ;
  wire \DLX_EXinst__n0016<26>/XORG ;
  wire DLX_EXinst_Maddsub__n0016_inst_lut3_33;
  wire DLX_EXinst_Maddsub__n0016_inst_cy_96;
  wire \DLX_EXinst__n0016<26>/CYINIT ;
  wire DLX_EXinst_Maddsub__n0016_inst_lut3_34;
  wire \DLX_EXinst__n0016<28>/XORF ;
  wire \DLX_EXinst__n0016<28>/CYMUXG ;
  wire \DLX_EXinst__n0016<28>/XORG ;
  wire DLX_EXinst_Maddsub__n0016_inst_lut3_35;
  wire DLX_EXinst_Maddsub__n0016_inst_cy_98;
  wire \DLX_EXinst__n0016<28>/CYINIT ;
  wire DLX_EXinst_Maddsub__n0016_inst_lut3_36;
  wire \DLX_EXinst__n0016<30>/XORF ;
  wire \DLX_EXinst__n0016<30>/XORG ;
  wire DLX_EXinst_Maddsub__n0016_inst_lut3_37;
  wire DLX_EXinst_Maddsub__n0016_inst_cy_100;
  wire \DLX_EXinst__n0016<30>/CYINIT ;
  wire DLX_IDinst_Mcompar__n0078_inst_lut4_40;
  wire \DLX_IDinst_Mcompar__n0078_inst_cy_263/CYMUXG ;
  wire DLX_IDinst_Mcompar__n0078_inst_lut4_41;
  wire DLX_IDinst_Mcompar__n0078_inst_cy_262;
  wire \DLX_IDinst_Mcompar__n0078_inst_cy_263/LOGIC_ZERO ;
  wire \DLX_IDinst_Mcompar__n0078_inst_cy_263/LOGIC_ONE ;
  wire \DLX_IDinst__n0078/LOGIC_ZERO ;
  wire DLX_IDinst_Mcompar__n0078_inst_lut4_42;
  wire \DLX_IDinst__n0078/CYMUXF ;
  wire \DLX_IDinst__n0078/CYINIT ;
  wire \NPC_eff<9>/OFF/RST ;
  wire DLX_EXinst_Mcompar__n0087_inst_lut4_16;
  wire \DLX_EXinst_Mcompar__n0087_inst_cy_119/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0087_inst_lut4_17;
  wire DLX_EXinst_Mcompar__n0087_inst_cy_118;
  wire \DLX_EXinst_Mcompar__n0087_inst_cy_119/LOGIC_ONE ;
  wire \DLX_EXinst_Mcompar__n0087_inst_cy_119/LOGIC_ZERO ;
  wire DLX_EXinst_Mcompar__n0087_inst_lut4_18;
  wire \DLX_EXinst_Mcompar__n0087_inst_cy_121/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0087_inst_lut4_19;
  wire DLX_EXinst_Mcompar__n0087_inst_cy_120;
  wire \DLX_EXinst_Mcompar__n0087_inst_cy_121/LOGIC_ONE ;
  wire \DLX_EXinst_Mcompar__n0087_inst_cy_121/CYINIT ;
  wire DLX_EXinst_Mcompar__n0087_inst_lut4_20;
  wire \DLX_EXinst_Mcompar__n0087_inst_cy_123/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0087_inst_lut4_21;
  wire DLX_EXinst_Mcompar__n0087_inst_cy_122;
  wire \DLX_EXinst_Mcompar__n0087_inst_cy_123/LOGIC_ONE ;
  wire \DLX_EXinst_Mcompar__n0087_inst_cy_123/CYINIT ;
  wire DLX_EXinst_Mcompar__n0087_inst_lut4_22;
  wire \DLX_EXinst_Mcompar__n0087_inst_cy_125/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0087_inst_lut4_23;
  wire DLX_EXinst_Mcompar__n0087_inst_cy_124;
  wire \DLX_EXinst_Mcompar__n0087_inst_cy_125/LOGIC_ONE ;
  wire \DLX_EXinst_Mcompar__n0087_inst_cy_125/CYINIT ;
  wire DLX_EXinst_Mcompar__n0087_inst_lut4_24;
  wire \DLX_EXinst_Mcompar__n0087_inst_cy_127/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0087_inst_lut4_25;
  wire DLX_EXinst_Mcompar__n0087_inst_cy_126;
  wire \DLX_EXinst_Mcompar__n0087_inst_cy_127/LOGIC_ONE ;
  wire \DLX_EXinst_Mcompar__n0087_inst_cy_127/CYINIT ;
  wire DLX_EXinst_Mcompar__n0087_inst_lut4_26;
  wire \DLX_EXinst_Mcompar__n0087_inst_cy_129/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0087_inst_lut4_27;
  wire DLX_EXinst_Mcompar__n0087_inst_cy_128;
  wire \DLX_EXinst_Mcompar__n0087_inst_cy_129/LOGIC_ONE ;
  wire \DLX_EXinst_Mcompar__n0087_inst_cy_129/CYINIT ;
  wire DLX_EXinst_Mcompar__n0087_inst_lut4_28;
  wire \DLX_EXinst_Mcompar__n0087_inst_cy_131/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0087_inst_lut4_29;
  wire DLX_EXinst_Mcompar__n0087_inst_cy_130;
  wire \DLX_EXinst_Mcompar__n0087_inst_cy_131/LOGIC_ONE ;
  wire \DLX_EXinst_Mcompar__n0087_inst_cy_131/CYINIT ;
  wire DLX_EXinst_Mcompar__n0087_inst_lut4_30;
  wire \DLX_EXinst__n0087/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0087_inst_lut4_31;
  wire DLX_EXinst_Mcompar__n0087_inst_cy_132;
  wire \DLX_EXinst__n0087/LOGIC_ONE ;
  wire \DLX_EXinst__n0087/CYINIT ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_166;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_231/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_167;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_230;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_231/LOGIC_ZERO ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_168;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_233/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_169;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_232;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_233/CYINIT ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_170;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_235/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_171;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_234;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_235/CYINIT ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_172;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_237/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_173;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_236;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_237/CYINIT ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_174;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_239/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_175;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_238;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_239/CYINIT ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_176;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_241/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_177;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_240;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_241/CYINIT ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_178;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_243/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_179;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_242;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_243/CYINIT ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_180;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_245/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_181;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_244;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_245/CYINIT ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_182;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_247/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_183;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_246;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_247/CYINIT ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_184;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_249/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_185;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_248;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_249/CYINIT ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_186;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_251/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_187;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_250;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_251/CYINIT ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_188;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_253/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_189;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_252;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_253/CYINIT ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_190;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_255/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_191;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_254;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_255/CYINIT ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_192;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_257/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_193;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_256;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_257/CYINIT ;
  wire \stall/OFF/RST ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_194;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_259/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_195;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_258;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_259/CYINIT ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_196;
  wire \CHOICE5769/CYMUXF ;
  wire \CHOICE5769/GROM ;
  wire \CHOICE5769/CYINIT ;
  wire vga_top_vga1_Mcompar__n0030_inst_lut4_48;
  wire \vga_top_vga1_Mcompar__n0030_inst_cy_358/CYMUXG ;
  wire vga_top_vga1_Mcompar__n0030_inst_lut4_49;
  wire vga_top_vga1_Mcompar__n0030_inst_cy_357;
  wire \vga_top_vga1_Mcompar__n0030_inst_cy_358/LOGIC_ZERO ;
  wire \vga_top_vga1_Mcompar__n0030_inst_cy_358/LOGIC_ONE ;
  wire vga_top_vga1_Mcompar__n0030_inst_lut1_10;
  wire \vga_top_vga1_Mcompar__n0030_inst_cy_360/CYMUXG ;
  wire vga_top_vga1_Mcompar__n0030_inst_lut1_11;
  wire vga_top_vga1_Mcompar__n0030_inst_cy_359;
  wire \vga_top_vga1_Mcompar__n0030_inst_cy_360/LOGIC_ONE ;
  wire \vga_top_vga1_Mcompar__n0030_inst_cy_360/CYINIT ;
  wire \$SIG_0 ;
  wire \vga_top_vga1_Mcompar__n0030_inst_cy_362/CYMUXG ;
  wire \$SIG_1 ;
  wire vga_top_vga1_Mcompar__n0030_inst_cy_361;
  wire \vga_top_vga1_Mcompar__n0030_inst_cy_362/LOGIC_ZERO ;
  wire \vga_top_vga1_Mcompar__n0030_inst_cy_362/CYINIT ;
  wire vga_top_vga1_Mcompar__n0030_inst_lut1_14;
  wire \vga_top_vga1_Mcompar__n0030_inst_cy_364/CYMUXG ;
  wire vga_top_vga1_Mcompar__n0030_inst_lut1_15;
  wire vga_top_vga1_Mcompar__n0030_inst_cy_363;
  wire \vga_top_vga1_Mcompar__n0030_inst_cy_364/LOGIC_ONE ;
  wire \vga_top_vga1_Mcompar__n0030_inst_cy_364/CYINIT ;
  wire \$SIG_2 ;
  wire \vga_top_vga1_Mcompar__n0030_inst_cy_366/CYMUXG ;
  wire \$SIG_3 ;
  wire vga_top_vga1_Mcompar__n0030_inst_cy_365;
  wire \vga_top_vga1_Mcompar__n0030_inst_cy_366/LOGIC_ZERO ;
  wire \vga_top_vga1_Mcompar__n0030_inst_cy_366/CYINIT ;
  wire vga_top_vga1_Mcompar__n0030_inst_lut1_18;
  wire \vga_top_vga1_Mcompar__n0030_inst_cy_368/CYMUXG ;
  wire vga_top_vga1_Mcompar__n0030_inst_lut1_19;
  wire vga_top_vga1_Mcompar__n0030_inst_cy_367;
  wire \vga_top_vga1_Mcompar__n0030_inst_cy_368/LOGIC_ONE ;
  wire \vga_top_vga1_Mcompar__n0030_inst_cy_368/CYINIT ;
  wire \$SIG_4 ;
  wire \vga_top_vga1_Mcompar__n0030_inst_cy_370/CYMUXG ;
  wire \$SIG_5 ;
  wire vga_top_vga1_Mcompar__n0030_inst_cy_369;
  wire \vga_top_vga1_Mcompar__n0030_inst_cy_370/LOGIC_ZERO ;
  wire \vga_top_vga1_Mcompar__n0030_inst_cy_370/CYINIT ;
  wire vga_top_vga1_Mcompar__n0030_inst_lut4_50;
  wire \vga_top_vga1__n0030/CYMUXG ;
  wire vga_top_vga1_Mcompar__n0030_inst_lut2_274;
  wire vga_top_vga1_Mcompar__n0030_inst_cy_371;
  wire \vga_top_vga1__n0030/LOGIC_ONE ;
  wire \vga_top_vga1__n0030/CYINIT ;
  wire DLX_IFinst_Madd__n0005_inst_lut2_40;
  wire \DLX_IFinst__n0015<3>/CYMUXG ;
  wire \DLX_IFinst__n0015<3>/XORG ;
  wire \DLX_IFinst__n0015<3>/GROM ;
  wire DLX_IFinst_Madd__n0005_inst_cy_40;
  wire \DLX_IFinst__n0015<3>/LOGIC_ZERO ;
  wire \DLX_IFinst__n0015<4>/FROM ;
  wire \DLX_IFinst__n0015<4>/XORF ;
  wire \DLX_IFinst__n0015<4>/CYMUXG ;
  wire \DLX_IFinst__n0015<4>/LOGIC_ZERO ;
  wire \DLX_IFinst__n0015<4>/XORG ;
  wire \DLX_IFinst__n0015<4>/GROM ;
  wire DLX_IFinst_Madd__n0005_inst_cy_42;
  wire \DLX_IFinst__n0015<4>/CYINIT ;
  wire \DLX_IFinst__n0015<6>/FROM ;
  wire \DLX_IFinst__n0015<6>/XORF ;
  wire \DLX_IFinst__n0015<6>/CYMUXG ;
  wire \DLX_IFinst__n0015<6>/LOGIC_ZERO ;
  wire \DLX_IFinst__n0015<6>/XORG ;
  wire \DLX_IFinst__n0015<6>/GROM ;
  wire DLX_IFinst_Madd__n0005_inst_cy_44;
  wire \DLX_IFinst__n0015<6>/CYINIT ;
  wire \DLX_IFinst__n0015<8>/FROM ;
  wire \DLX_IFinst__n0015<8>/XORF ;
  wire \DLX_IFinst__n0015<8>/CYMUXG ;
  wire \DLX_IFinst__n0015<8>/LOGIC_ZERO ;
  wire \DLX_IFinst__n0015<8>/XORG ;
  wire \DLX_IFinst__n0015<8>/GROM ;
  wire DLX_IFinst_Madd__n0005_inst_cy_46;
  wire \DLX_IFinst__n0015<8>/CYINIT ;
  wire \DLX_IFinst__n0015<10>/FROM ;
  wire \DLX_IFinst__n0015<10>/XORF ;
  wire \DLX_IFinst__n0015<10>/CYMUXG ;
  wire \DLX_IFinst__n0015<10>/LOGIC_ZERO ;
  wire \DLX_IFinst__n0015<10>/XORG ;
  wire \DLX_IFinst__n0015<10>/GROM ;
  wire DLX_IFinst_Madd__n0005_inst_cy_48;
  wire \DLX_IFinst__n0015<10>/CYINIT ;
  wire \DLX_IFinst__n0015<12>/FROM ;
  wire \DLX_IFinst__n0015<12>/XORF ;
  wire \DLX_IFinst__n0015<12>/CYMUXG ;
  wire \DLX_IFinst__n0015<12>/LOGIC_ZERO ;
  wire \DLX_IFinst__n0015<12>/XORG ;
  wire \DLX_IFinst__n0015<12>/GROM ;
  wire DLX_IFinst_Madd__n0005_inst_cy_50;
  wire \DLX_IFinst__n0015<12>/CYINIT ;
  wire \DLX_IFinst__n0015<14>/FROM ;
  wire \DLX_IFinst__n0015<14>/XORF ;
  wire \DLX_IFinst__n0015<14>/CYMUXG ;
  wire \DLX_IFinst__n0015<14>/LOGIC_ZERO ;
  wire \DLX_IFinst__n0015<14>/XORG ;
  wire \DLX_IFinst__n0015<14>/GROM ;
  wire DLX_IFinst_Madd__n0005_inst_cy_52;
  wire \DLX_IFinst__n0015<14>/CYINIT ;
  wire \DLX_IFinst__n0015<16>/FROM ;
  wire \DLX_IFinst__n0015<16>/XORF ;
  wire \DLX_IFinst__n0015<16>/CYMUXG ;
  wire \DLX_IFinst__n0015<16>/LOGIC_ZERO ;
  wire \DLX_IFinst__n0015<16>/XORG ;
  wire \DLX_IFinst__n0015<16>/GROM ;
  wire DLX_IFinst_Madd__n0005_inst_cy_54;
  wire \DLX_IFinst__n0015<16>/CYINIT ;
  wire \CLI/OFF/RST ;
  wire \DLX_IFinst__n0015<18>/FROM ;
  wire \DLX_IFinst__n0015<18>/XORF ;
  wire \DLX_IFinst__n0015<18>/CYMUXG ;
  wire \DLX_IFinst__n0015<18>/LOGIC_ZERO ;
  wire \DLX_IFinst__n0015<18>/XORG ;
  wire \DLX_IFinst__n0015<18>/GROM ;
  wire DLX_IFinst_Madd__n0005_inst_cy_56;
  wire \DLX_IFinst__n0015<18>/CYINIT ;
  wire \DLX_IFinst__n0015<20>/FROM ;
  wire \DLX_IFinst__n0015<20>/XORF ;
  wire \DLX_IFinst__n0015<20>/CYMUXG ;
  wire \DLX_IFinst__n0015<20>/LOGIC_ZERO ;
  wire \DLX_IFinst__n0015<20>/XORG ;
  wire \DLX_IFinst__n0015<20>/GROM ;
  wire DLX_IFinst_Madd__n0005_inst_cy_58;
  wire \DLX_IFinst__n0015<20>/CYINIT ;
  wire \DLX_IFinst__n0015<22>/FROM ;
  wire \DLX_IFinst__n0015<22>/XORF ;
  wire \DLX_IFinst__n0015<22>/CYMUXG ;
  wire \DLX_IFinst__n0015<22>/LOGIC_ZERO ;
  wire \DLX_IFinst__n0015<22>/XORG ;
  wire \DLX_IFinst__n0015<22>/GROM ;
  wire DLX_IFinst_Madd__n0005_inst_cy_60;
  wire \DLX_IFinst__n0015<22>/CYINIT ;
  wire \DLX_IFinst__n0015<24>/FROM ;
  wire \DLX_IFinst__n0015<24>/XORF ;
  wire \DLX_IFinst__n0015<24>/CYMUXG ;
  wire \DLX_IFinst__n0015<24>/LOGIC_ZERO ;
  wire \DLX_IFinst__n0015<24>/XORG ;
  wire \DLX_IFinst__n0015<24>/GROM ;
  wire DLX_IFinst_Madd__n0005_inst_cy_62;
  wire \DLX_IFinst__n0015<24>/CYINIT ;
  wire \DLX_IFinst__n0015<26>/FROM ;
  wire \DLX_IFinst__n0015<26>/XORF ;
  wire \DLX_IFinst__n0015<26>/CYMUXG ;
  wire \DLX_IFinst__n0015<26>/LOGIC_ZERO ;
  wire \DLX_IFinst__n0015<26>/XORG ;
  wire \DLX_IFinst__n0015<26>/GROM ;
  wire DLX_IFinst_Madd__n0005_inst_cy_64;
  wire \DLX_IFinst__n0015<26>/CYINIT ;
  wire \DLX_IFinst__n0015<28>/FROM ;
  wire \DLX_IFinst__n0015<28>/XORF ;
  wire \DLX_IFinst__n0015<28>/CYMUXG ;
  wire \DLX_IFinst__n0015<28>/LOGIC_ZERO ;
  wire \DLX_IFinst__n0015<28>/XORG ;
  wire \DLX_IFinst__n0015<28>/GROM ;
  wire DLX_IFinst_Madd__n0005_inst_cy_66;
  wire \DLX_IFinst__n0015<28>/CYINIT ;
  wire \DLX_IFinst__n0015<30>/LOGIC_ZERO ;
  wire \DLX_IFinst__n0015<30>/FROM ;
  wire \DLX_IFinst__n0015<30>/XORF ;
  wire \DLX_IFinst__n0015<30>/XORG ;
  wire \DLX_IFinst_NPC<31>_rt ;
  wire DLX_IFinst_Madd__n0005_inst_cy_68;
  wire \DLX_IFinst__n0015<30>/CYINIT ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_70;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_135/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_71;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_134;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_135/LOGIC_ZERO ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_72;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_137/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_73;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_136;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_137/CYINIT ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_74;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_139/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_75;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_138;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_139/CYINIT ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_76;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_141/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_77;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_140;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_141/CYINIT ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_78;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_143/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_79;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_142;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_143/CYINIT ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_80;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_145/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_81;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_144;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_145/CYINIT ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_82;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_147/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_83;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_146;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_147/CYINIT ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_84;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_149/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_85;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_148;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_149/CYINIT ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_86;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_151/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_87;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_150;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_151/CYINIT ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_88;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_153/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_89;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_152;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_153/CYINIT ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_90;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_155/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_91;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_154;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_155/CYINIT ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_92;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_157/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_93;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_156;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_157/CYINIT ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_94;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_159/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_95;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_158;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_159/CYINIT ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_96;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_161/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_97;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_160;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_161/CYINIT ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_98;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_163/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_99;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_162;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_163/CYINIT ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_100;
  wire \CHOICE5806/CYMUXF ;
  wire \CHOICE5806/GROM ;
  wire \CHOICE5806/CYINIT ;
  wire vga_top_vga1_gridvcounter_Madd__n0000_inst_lut2_0;
  wire \vga_top_vga1_gridvcounter<0>/CYMUXG ;
  wire \vga_top_vga1_gridvcounter<0>/GROM ;
  wire vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_0;
  wire \vga_top_vga1_gridvcounter<0>/LOGIC_ZERO ;
  wire \vga_top_vga1_gridvcounter<2>/FROM ;
  wire \vga_top_vga1_gridvcounter<2>/CYMUXG ;
  wire \vga_top_vga1_gridvcounter<2>/LOGIC_ZERO ;
  wire \vga_top_vga1_gridvcounter<2>/GROM ;
  wire vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_2;
  wire \vga_top_vga1_gridvcounter<2>/CYINIT ;
  wire \vga_top_vga1_gridvcounter<4>/FROM ;
  wire \vga_top_vga1_gridvcounter<4>/CYMUXG ;
  wire \vga_top_vga1_gridvcounter<4>/LOGIC_ZERO ;
  wire \vga_top_vga1_gridvcounter<4>/GROM ;
  wire vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_4;
  wire \vga_top_vga1_gridvcounter<4>/CYINIT ;
  wire \DM_addr_eff<0>/OFF/RST ;
  wire \vga_top_vga1_gridvcounter<6>/FROM ;
  wire \vga_top_vga1_gridvcounter<6>/CYMUXG ;
  wire \vga_top_vga1_gridvcounter<6>/LOGIC_ZERO ;
  wire \vga_top_vga1_gridvcounter<6>/GROM ;
  wire vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_6;
  wire \vga_top_vga1_gridvcounter<6>/CYINIT ;
  wire \vga_top_vga1_gridvcounter<8>_rt ;
  wire \vga_top_vga1_gridvcounter<8>/CYINIT ;
  wire vga_top_vga1_Mcompar__n0033_inst_lut1_4;
  wire \vga_top_vga1_Mcompar__n0033_inst_cy_344/CYMUXG ;
  wire vga_top_vga1_Mcompar__n0033_inst_lut1_5;
  wire vga_top_vga1_Mcompar__n0033_inst_cy_343;
  wire \vga_top_vga1_Mcompar__n0033_inst_cy_344/LOGIC_ZERO ;
  wire \vga_top_vga1_Mcompar__n0033_inst_cy_344/LOGIC_ONE ;
  wire vga_top_vga1_Mcompar__n0033_inst_lut2_269;
  wire \vga_top_vga1_Mcompar__n0033_inst_cy_346/CYMUXG ;
  wire vga_top_vga1_Mcompar__n0033_inst_lut2_270;
  wire vga_top_vga1_Mcompar__n0033_inst_cy_345;
  wire \vga_top_vga1_Mcompar__n0033_inst_cy_346/LOGIC_ONE ;
  wire \vga_top_vga1_Mcompar__n0033_inst_cy_346/CYINIT ;
  wire vga_top_vga1_Mcompar__n0033_inst_lut3_110;
  wire \vga_top_vga1_Mcompar__n0033_inst_cy_348/CYMUXG ;
  wire vga_top_vga1_Mcompar__n0033_inst_lut3_111;
  wire vga_top_vga1_Mcompar__n0033_inst_cy_347;
  wire \vga_top_vga1_Mcompar__n0033_inst_cy_348/LOGIC_ZERO ;
  wire \vga_top_vga1_Mcompar__n0033_inst_cy_348/CYINIT ;
  wire vga_top_vga1_Mcompar__n0033_inst_lut2_271;
  wire \vga_top_vga1_Mcompar__n0033_inst_cy_350/CYMUXG ;
  wire vga_top_vga1_Mcompar__n0033_inst_lut2_272;
  wire vga_top_vga1_Mcompar__n0033_inst_cy_349;
  wire \vga_top_vga1_Mcompar__n0033_inst_cy_350/LOGIC_ONE ;
  wire \vga_top_vga1_Mcompar__n0033_inst_cy_350/CYINIT ;
  wire vga_top_vga1_Mcompar__n0033_inst_lut1_6;
  wire \vga_top_vga1_Mcompar__n0033_inst_cy_352/CYMUXG ;
  wire vga_top_vga1_Mcompar__n0033_inst_lut1_7;
  wire vga_top_vga1_Mcompar__n0033_inst_cy_351;
  wire \vga_top_vga1_Mcompar__n0033_inst_cy_352/LOGIC_ZERO ;
  wire \vga_top_vga1_Mcompar__n0033_inst_cy_352/CYINIT ;
  wire \$SIG_7 ;
  wire \vga_top_vga1_Mcompar__n0033_inst_cy_354/CYMUXG ;
  wire \$SIG_8 ;
  wire vga_top_vga1_Mcompar__n0033_inst_cy_353;
  wire \vga_top_vga1_Mcompar__n0033_inst_cy_354/LOGIC_ONE ;
  wire \vga_top_vga1_Mcompar__n0033_inst_cy_354/CYINIT ;
  wire vga_top_vga1_Mcompar__n0033_inst_lut4_47;
  wire \vga_top_vga1__n0033/CYMUXG ;
  wire vga_top_vga1_Mcompar__n0033_inst_lut2_273;
  wire vga_top_vga1_Mcompar__n0033_inst_cy_355;
  wire \vga_top_vga1__n0033/LOGIC_ZERO ;
  wire \vga_top_vga1__n0033/CYINIT ;
  wire \$SIG_9 ;
  wire \vga_top_vga1_Mcompar__n0034_inst_cy_332/CYMUXG ;
  wire \$SIG_10 ;
  wire vga_top_vga1_Mcompar__n0034_inst_cy_331;
  wire \vga_top_vga1_Mcompar__n0034_inst_cy_332/LOGIC_ZERO ;
  wire \vga_top_vga1_Mcompar__n0034_inst_cy_332/LOGIC_ONE ;
  wire \DM_addr_eff<1>/OFF/RST ;
  wire vga_top_vga1_Mcompar__n0034_inst_lut2_262;
  wire \vga_top_vga1_Mcompar__n0034_inst_cy_334/CYMUXG ;
  wire vga_top_vga1_Mcompar__n0034_inst_lut2_263;
  wire vga_top_vga1_Mcompar__n0034_inst_cy_333;
  wire \vga_top_vga1_Mcompar__n0034_inst_cy_334/LOGIC_ONE ;
  wire \vga_top_vga1_Mcompar__n0034_inst_cy_334/CYINIT ;
  wire \$SIG_11 ;
  wire \vga_top_vga1_Mcompar__n0034_inst_cy_336/CYMUXG ;
  wire \$SIG_12 ;
  wire vga_top_vga1_Mcompar__n0034_inst_cy_335;
  wire \vga_top_vga1_Mcompar__n0034_inst_cy_336/LOGIC_ZERO ;
  wire \vga_top_vga1_Mcompar__n0034_inst_cy_336/CYINIT ;
  wire vga_top_vga1_Mcompar__n0034_inst_lut2_264;
  wire \vga_top_vga1_Mcompar__n0034_inst_cy_338/CYMUXG ;
  wire vga_top_vga1_Mcompar__n0034_inst_lut2_265;
  wire vga_top_vga1_Mcompar__n0034_inst_cy_337;
  wire \vga_top_vga1_Mcompar__n0034_inst_cy_338/LOGIC_ONE ;
  wire \vga_top_vga1_Mcompar__n0034_inst_cy_338/CYINIT ;
  wire vga_top_vga1_Mcompar__n0034_inst_lut2_266;
  wire \vga_top_vga1_Mcompar__n0034_inst_cy_340/CYMUXG ;
  wire vga_top_vga1_Mcompar__n0034_inst_lut2_267;
  wire vga_top_vga1_Mcompar__n0034_inst_cy_339;
  wire \vga_top_vga1_Mcompar__n0034_inst_cy_340/LOGIC_ZERO ;
  wire \vga_top_vga1_Mcompar__n0034_inst_cy_340/CYINIT ;
  wire vga_top_vga1_Mcompar__n0034_inst_lut4_46;
  wire \vga_top_vga1__n0034/CYMUXG ;
  wire vga_top_vga1_Mcompar__n0034_inst_lut2_268;
  wire vga_top_vga1_Mcompar__n0034_inst_cy_341;
  wire \vga_top_vga1__n0034/LOGIC_ONE ;
  wire \vga_top_vga1__n0034/CYINIT ;
  wire DLX_IDinst_Msub__n0128_inst_lut2_230;
  wire \DLX_IDinst__n0128<0>/XORF ;
  wire \DLX_IDinst__n0128<0>/CYMUXG ;
  wire \DLX_IDinst__n0128<0>/XORG ;
  wire DLX_IDinst_Msub__n0128_inst_lut2_231;
  wire DLX_IDinst_Msub__n0128_inst_cy_299;
  wire \DLX_IDinst__n0128<0>/CYINIT ;
  wire \DLX_IDinst__n0128<0>/LOGIC_ONE ;
  wire \DLX_IDinst__n0128<2>/FROM ;
  wire \DLX_IDinst__n0128<2>/XORF ;
  wire \DLX_IDinst__n0128<2>/CYMUXG ;
  wire \DLX_IDinst__n0128<2>/XORG ;
  wire DLX_IDinst_Msub__n0128_inst_lut2_233;
  wire DLX_IDinst_Msub__n0128_inst_cy_301;
  wire \DLX_IDinst__n0128<2>/CYINIT ;
  wire DLX_IDinst_Msub__n0128_inst_lut2_234;
  wire \DLX_IDinst__n0128<4>/XORF ;
  wire \DLX_IDinst__n0128<4>/CYMUXG ;
  wire \DLX_IDinst__n0128<4>/XORG ;
  wire DLX_IDinst_Msub__n0128_inst_lut2_235;
  wire DLX_IDinst_Msub__n0128_inst_cy_303;
  wire \DLX_IDinst__n0128<4>/CYINIT ;
  wire DLX_IDinst_Msub__n0128_inst_lut2_236;
  wire \DLX_IDinst__n0128<6>/XORF ;
  wire \DLX_IDinst__n0128<6>/CYMUXG ;
  wire \DLX_IDinst__n0128<6>/XORG ;
  wire DLX_IDinst_Msub__n0128_inst_lut2_237;
  wire DLX_IDinst_Msub__n0128_inst_cy_305;
  wire \DLX_IDinst__n0128<6>/CYINIT ;
  wire DLX_IDinst_Msub__n0128_inst_lut2_238;
  wire \DLX_IDinst__n0128<8>/XORF ;
  wire \DLX_IDinst__n0128<8>/CYMUXG ;
  wire \DLX_IDinst__n0128<8>/XORG ;
  wire DLX_IDinst_Msub__n0128_inst_lut2_239;
  wire DLX_IDinst_Msub__n0128_inst_cy_307;
  wire \DLX_IDinst__n0128<8>/CYINIT ;
  wire DLX_IDinst_Msub__n0128_inst_lut2_240;
  wire \DLX_IDinst__n0128<10>/XORF ;
  wire \DLX_IDinst__n0128<10>/CYMUXG ;
  wire \DLX_IDinst__n0128<10>/XORG ;
  wire DLX_IDinst_Msub__n0128_inst_lut2_241;
  wire DLX_IDinst_Msub__n0128_inst_cy_309;
  wire \DLX_IDinst__n0128<10>/CYINIT ;
  wire DLX_IDinst_Msub__n0128_inst_lut2_242;
  wire \DLX_IDinst__n0128<12>/XORF ;
  wire \DLX_IDinst__n0128<12>/CYMUXG ;
  wire \DLX_IDinst__n0128<12>/XORG ;
  wire DLX_IDinst_Msub__n0128_inst_lut2_243;
  wire DLX_IDinst_Msub__n0128_inst_cy_311;
  wire \DLX_IDinst__n0128<12>/CYINIT ;
  wire DLX_IDinst_Msub__n0128_inst_lut2_244;
  wire \DLX_IDinst__n0128<14>/XORF ;
  wire \DLX_IDinst__n0128<14>/CYMUXG ;
  wire \DLX_IDinst__n0128<14>/XORG ;
  wire DLX_IDinst_Msub__n0128_inst_lut2_245;
  wire DLX_IDinst_Msub__n0128_inst_cy_313;
  wire \DLX_IDinst__n0128<14>/CYINIT ;
  wire DLX_IDinst_Msub__n0128_inst_lut2_246;
  wire \DLX_IDinst__n0128<16>/XORF ;
  wire \DLX_IDinst__n0128<16>/CYMUXG ;
  wire \DLX_IDinst__n0128<16>/XORG ;
  wire DLX_IDinst_Msub__n0128_inst_lut2_247;
  wire DLX_IDinst_Msub__n0128_inst_cy_315;
  wire \DLX_IDinst__n0128<16>/CYINIT ;
  wire \DM_addr_eff<2>/OFF/RST ;
  wire DLX_IDinst_Msub__n0128_inst_lut2_248;
  wire \DLX_IDinst__n0128<18>/XORF ;
  wire \DLX_IDinst__n0128<18>/CYMUXG ;
  wire \DLX_IDinst__n0128<18>/XORG ;
  wire DLX_IDinst_Msub__n0128_inst_lut2_249;
  wire DLX_IDinst_Msub__n0128_inst_cy_317;
  wire \DLX_IDinst__n0128<18>/CYINIT ;
  wire DLX_IDinst_Msub__n0128_inst_lut2_250;
  wire \DLX_IDinst__n0128<20>/XORF ;
  wire \DLX_IDinst__n0128<20>/CYMUXG ;
  wire \DLX_IDinst__n0128<20>/XORG ;
  wire DLX_IDinst_Msub__n0128_inst_lut2_251;
  wire DLX_IDinst_Msub__n0128_inst_cy_319;
  wire \DLX_IDinst__n0128<20>/CYINIT ;
  wire DLX_IDinst_Msub__n0128_inst_lut2_252;
  wire \DLX_IDinst__n0128<22>/XORF ;
  wire \DLX_IDinst__n0128<22>/CYMUXG ;
  wire \DLX_IDinst__n0128<22>/XORG ;
  wire DLX_IDinst_Msub__n0128_inst_lut2_253;
  wire DLX_IDinst_Msub__n0128_inst_cy_321;
  wire \DLX_IDinst__n0128<22>/CYINIT ;
  wire DLX_IDinst_Msub__n0128_inst_lut2_254;
  wire \DLX_IDinst__n0128<24>/XORF ;
  wire \DLX_IDinst__n0128<24>/CYMUXG ;
  wire \DLX_IDinst__n0128<24>/XORG ;
  wire DLX_IDinst_Msub__n0128_inst_lut2_255;
  wire DLX_IDinst_Msub__n0128_inst_cy_323;
  wire \DLX_IDinst__n0128<24>/CYINIT ;
  wire DLX_IDinst_Msub__n0128_inst_lut2_256;
  wire \DLX_IDinst__n0128<26>/XORF ;
  wire \DLX_IDinst__n0128<26>/CYMUXG ;
  wire \DLX_IDinst__n0128<26>/XORG ;
  wire DLX_IDinst_Msub__n0128_inst_lut2_257;
  wire DLX_IDinst_Msub__n0128_inst_cy_325;
  wire \DLX_IDinst__n0128<26>/CYINIT ;
  wire DLX_IDinst_Msub__n0128_inst_lut2_258;
  wire \DLX_IDinst__n0128<28>/XORF ;
  wire \DLX_IDinst__n0128<28>/CYMUXG ;
  wire \DLX_IDinst__n0128<28>/XORG ;
  wire DLX_IDinst_Msub__n0128_inst_lut2_259;
  wire DLX_IDinst_Msub__n0128_inst_cy_327;
  wire \DLX_IDinst__n0128<28>/CYINIT ;
  wire DLX_IDinst_Msub__n0128_inst_lut2_260;
  wire \DLX_IDinst__n0128<30>/XORF ;
  wire \DLX_IDinst__n0128<30>/XORG ;
  wire DLX_IDinst_Msub__n0128_inst_lut2_261;
  wire DLX_IDinst_Msub__n0128_inst_cy_329;
  wire \DLX_IDinst__n0128<30>/CYINIT ;
  wire DLX_EXinst_Mcompar__n0053_inst_lut4_0;
  wire \DLX_EXinst_Mcompar__n0053_inst_cy_103/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0053_inst_lut4_1;
  wire DLX_EXinst_Mcompar__n0053_inst_cy_102;
  wire \DLX_EXinst_Mcompar__n0053_inst_cy_103/LOGIC_ZERO ;
  wire \DLX_EXinst_Mcompar__n0053_inst_cy_103/LOGIC_ONE ;
  wire DLX_EXinst_Mcompar__n0053_inst_lut4_2;
  wire \DLX_EXinst_Mcompar__n0053_inst_cy_105/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0053_inst_lut4_3;
  wire DLX_EXinst_Mcompar__n0053_inst_cy_104;
  wire \DLX_EXinst_Mcompar__n0053_inst_cy_105/LOGIC_ZERO ;
  wire \DLX_EXinst_Mcompar__n0053_inst_cy_105/CYINIT ;
  wire DLX_EXinst_Mcompar__n0053_inst_lut4_4;
  wire \DLX_EXinst_Mcompar__n0053_inst_cy_107/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0053_inst_lut4_5;
  wire DLX_EXinst_Mcompar__n0053_inst_cy_106;
  wire \DLX_EXinst_Mcompar__n0053_inst_cy_107/LOGIC_ZERO ;
  wire \DLX_EXinst_Mcompar__n0053_inst_cy_107/CYINIT ;
  wire DLX_EXinst_Mcompar__n0053_inst_lut4_6;
  wire \DLX_EXinst_Mcompar__n0053_inst_cy_109/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0053_inst_lut4_7;
  wire DLX_EXinst_Mcompar__n0053_inst_cy_108;
  wire \DLX_EXinst_Mcompar__n0053_inst_cy_109/LOGIC_ZERO ;
  wire \DLX_EXinst_Mcompar__n0053_inst_cy_109/CYINIT ;
  wire DLX_EXinst_Mcompar__n0053_inst_lut4_8;
  wire \DLX_EXinst_Mcompar__n0053_inst_cy_111/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0053_inst_lut4_9;
  wire DLX_EXinst_Mcompar__n0053_inst_cy_110;
  wire \DLX_EXinst_Mcompar__n0053_inst_cy_111/LOGIC_ZERO ;
  wire \DLX_EXinst_Mcompar__n0053_inst_cy_111/CYINIT ;
  wire DLX_EXinst_Mcompar__n0053_inst_lut4_10;
  wire \DLX_EXinst_Mcompar__n0053_inst_cy_113/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0053_inst_lut4_11;
  wire DLX_EXinst_Mcompar__n0053_inst_cy_112;
  wire \DLX_EXinst_Mcompar__n0053_inst_cy_113/LOGIC_ZERO ;
  wire \DLX_EXinst_Mcompar__n0053_inst_cy_113/CYINIT ;
  wire DLX_EXinst_Mcompar__n0053_inst_lut4_12;
  wire \DLX_EXinst_Mcompar__n0053_inst_cy_115/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0053_inst_lut4_13;
  wire DLX_EXinst_Mcompar__n0053_inst_cy_114;
  wire \DLX_EXinst_Mcompar__n0053_inst_cy_115/LOGIC_ZERO ;
  wire \DLX_EXinst_Mcompar__n0053_inst_cy_115/CYINIT ;
  wire DLX_EXinst_Mcompar__n0053_inst_lut4_14;
  wire \DLX_EXinst__n0053/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0053_inst_lut4_15;
  wire DLX_EXinst_Mcompar__n0053_inst_cy_116;
  wire \DLX_EXinst__n0053/LOGIC_ZERO ;
  wire \DLX_EXinst__n0053/CYINIT ;
  wire DLX_EXinst_Mcompar__n0061_inst_lut2_134;
  wire \DLX_EXinst_Mcompar__n0061_inst_cy_199/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0061_inst_lut2_135;
  wire DLX_EXinst_Mcompar__n0061_inst_cy_198;
  wire \DLX_EXinst_Mcompar__n0061_inst_cy_199/LOGIC_ZERO ;
  wire DLX_EXinst_Mcompar__n0061_inst_lut2_136;
  wire \DLX_EXinst_Mcompar__n0061_inst_cy_201/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0061_inst_lut2_137;
  wire DLX_EXinst_Mcompar__n0061_inst_cy_200;
  wire \DLX_EXinst_Mcompar__n0061_inst_cy_201/CYINIT ;
  wire DLX_EXinst_Mcompar__n0061_inst_lut2_138;
  wire \DLX_EXinst_Mcompar__n0061_inst_cy_203/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0061_inst_lut2_139;
  wire DLX_EXinst_Mcompar__n0061_inst_cy_202;
  wire \DLX_EXinst_Mcompar__n0061_inst_cy_203/CYINIT ;
  wire DLX_EXinst_Mcompar__n0061_inst_lut2_140;
  wire \DLX_EXinst_Mcompar__n0061_inst_cy_205/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0061_inst_lut2_141;
  wire DLX_EXinst_Mcompar__n0061_inst_cy_204;
  wire \DLX_EXinst_Mcompar__n0061_inst_cy_205/CYINIT ;
  wire DLX_EXinst_Mcompar__n0061_inst_lut2_142;
  wire \DLX_EXinst_Mcompar__n0061_inst_cy_207/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0061_inst_lut2_143;
  wire DLX_EXinst_Mcompar__n0061_inst_cy_206;
  wire \DLX_EXinst_Mcompar__n0061_inst_cy_207/CYINIT ;
  wire \DM_addr_eff<3>/OFF/RST ;
  wire DLX_EXinst_Mcompar__n0061_inst_lut2_144;
  wire \DLX_EXinst_Mcompar__n0061_inst_cy_209/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0061_inst_lut2_145;
  wire DLX_EXinst_Mcompar__n0061_inst_cy_208;
  wire \DLX_EXinst_Mcompar__n0061_inst_cy_209/CYINIT ;
  wire DLX_EXinst_Mcompar__n0061_inst_lut2_146;
  wire \DLX_EXinst_Mcompar__n0061_inst_cy_211/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0061_inst_lut2_147;
  wire DLX_EXinst_Mcompar__n0061_inst_cy_210;
  wire \DLX_EXinst_Mcompar__n0061_inst_cy_211/CYINIT ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_168;
  wire \DLX_EXinst_Mcompar__n0063_inst_cy_233/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_169;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_232;
  wire \DLX_EXinst_Mcompar__n0063_inst_cy_233/CYINIT ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_170;
  wire \DLX_EXinst_Mcompar__n0063_inst_cy_235/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_171;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_234;
  wire \DLX_EXinst_Mcompar__n0063_inst_cy_235/CYINIT ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_172;
  wire \DLX_EXinst_Mcompar__n0063_inst_cy_237/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_173;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_236;
  wire \DLX_EXinst_Mcompar__n0063_inst_cy_237/CYINIT ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_174;
  wire \DLX_EXinst_Mcompar__n0063_inst_cy_239/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_175;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_238;
  wire \DLX_EXinst_Mcompar__n0063_inst_cy_239/CYINIT ;
  wire \DM_addr_eff<5>/OFF/RST ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_176;
  wire \DLX_EXinst_Mcompar__n0063_inst_cy_241/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_177;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_240;
  wire \DLX_EXinst_Mcompar__n0063_inst_cy_241/CYINIT ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_178;
  wire \DLX_EXinst_Mcompar__n0063_inst_cy_243/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_179;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_242;
  wire \DLX_EXinst_Mcompar__n0063_inst_cy_243/CYINIT ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_180;
  wire \DLX_EXinst_Mcompar__n0063_inst_cy_245/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_181;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_244;
  wire \DLX_EXinst_Mcompar__n0063_inst_cy_245/CYINIT ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_182;
  wire \DLX_EXinst_Mcompar__n0063_inst_cy_247/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_183;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_246;
  wire \DLX_EXinst_Mcompar__n0063_inst_cy_247/CYINIT ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_184;
  wire \DLX_EXinst_Mcompar__n0063_inst_cy_249/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_185;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_248;
  wire \DLX_EXinst_Mcompar__n0063_inst_cy_249/CYINIT ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_186;
  wire \DLX_EXinst_Mcompar__n0063_inst_cy_251/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_187;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_250;
  wire \DLX_EXinst_Mcompar__n0063_inst_cy_251/CYINIT ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_188;
  wire \DLX_EXinst_Mcompar__n0063_inst_cy_253/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_189;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_252;
  wire \DLX_EXinst_Mcompar__n0063_inst_cy_253/CYINIT ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_190;
  wire \DLX_EXinst_Mcompar__n0063_inst_cy_255/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_191;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_254;
  wire \DLX_EXinst_Mcompar__n0063_inst_cy_255/CYINIT ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_192;
  wire \DLX_EXinst_Mcompar__n0063_inst_cy_257/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_193;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_256;
  wire \DLX_EXinst_Mcompar__n0063_inst_cy_257/CYINIT ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_194;
  wire \DLX_EXinst_Mcompar__n0063_inst_cy_259/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_195;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_258;
  wire \DLX_EXinst_Mcompar__n0063_inst_cy_259/CYINIT ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_196;
  wire \CHOICE5291/CYMUXF ;
  wire \CHOICE5291/GROM ;
  wire \CHOICE5291/CYINIT ;
  wire vga_top_vga1_gridhcounter_Madd__n0000_inst_lut2_0;
  wire \vga_top_vga1_gridhcounter<0>/CYMUXG ;
  wire \vga_top_vga1_gridhcounter<0>/GROM ;
  wire vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_0;
  wire \vga_top_vga1_gridhcounter<0>/LOGIC_ZERO ;
  wire \vga_top_vga1_gridhcounter<2>/FROM ;
  wire \vga_top_vga1_gridhcounter<2>/CYMUXG ;
  wire \vga_top_vga1_gridhcounter<2>/LOGIC_ZERO ;
  wire \vga_top_vga1_gridhcounter<2>/GROM ;
  wire vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_2;
  wire \vga_top_vga1_gridhcounter<2>/CYINIT ;
  wire \vga_top_vga1_gridhcounter<4>/FROM ;
  wire \vga_top_vga1_gridhcounter<4>/CYMUXG ;
  wire \vga_top_vga1_gridhcounter<4>/LOGIC_ZERO ;
  wire \vga_top_vga1_gridhcounter<4>/GROM ;
  wire vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_4;
  wire \vga_top_vga1_gridhcounter<4>/CYINIT ;
  wire \vga_top_vga1_gridhcounter<6>/FROM ;
  wire \vga_top_vga1_gridhcounter<6>/CYMUXG ;
  wire \vga_top_vga1_gridhcounter<6>/LOGIC_ZERO ;
  wire \vga_top_vga1_gridhcounter<6>/GROM ;
  wire vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_6;
  wire \vga_top_vga1_gridhcounter<6>/CYINIT ;
  wire \vga_top_vga1_gridhcounter<8>_rt ;
  wire \vga_top_vga1_gridhcounter<8>/CYINIT ;
  wire \DLX_IDinst_current_IR<1>/FROM ;
  wire \DLX_IDinst_current_IR<1>/GROM ;
  wire \DLX_IDinst_current_IR<3>/FROM ;
  wire \DLX_IDinst_current_IR<3>/GROM ;
  wire \DLX_IDinst_current_IR<5>/FROM ;
  wire \DLX_IDinst_current_IR<5>/GROM ;
  wire \DLX_IDinst_current_IR<7>/FROM ;
  wire \DLX_IDinst_current_IR<7>/GROM ;
  wire \DM_addr_eff<6>/OFF/RST ;
  wire \DLX_IDinst_current_IR<9>/FROM ;
  wire \DLX_IDinst_current_IR<9>/GROM ;
  wire \DLX_IDinst_slot_num_FFd1/FROM ;
  wire \DLX_IDinst_slot_num_FFd1-In ;
  wire \DLX_EXinst_mem_to_reg_EX/FFY/RST ;
  wire DLX_EXinst__n0010;
  wire \DLX_EXinst_mem_to_reg_EX/GROM ;
  wire \vga_top_vga1_helpcounter<2>/FROM ;
  wire \DLX_IDinst_reg_out_B_2_1/GROM ;
  wire \DLX_IDinst_reg_out_B<3>/GROM ;
  wire \DLX_EXinst_ALU_result<13>/FROM ;
  wire \DLX_EXinst_ALU_result<13>/GROM ;
  wire \DLX_MEMinst_RF_data_in<11>/FFY/RST ;
  wire \DLX_MEMinst_RF_data_in<11>/CKMUXNOT ;
  wire \DLX_MEMinst_RF_data_in<21>/FFY/RST ;
  wire \DLX_MEMinst_RF_data_in<21>/CKMUXNOT ;
  wire \DM_addr_eff<7>/OFF/RST ;
  wire \DLX_MEMinst_RF_data_in<13>/FFY/RST ;
  wire \DLX_MEMinst_RF_data_in<13>/CKMUXNOT ;
  wire \DLX_MEMinst_RF_data_in<31>/FFY/RST ;
  wire \DLX_MEMinst_RF_data_in<31>/CKMUXNOT ;
  wire \DLX_MEMinst_RF_data_in<23>/FFY/RST ;
  wire \DLX_MEMinst_RF_data_in<23>/CKMUXNOT ;
  wire \DLX_MEMinst_RF_data_in<15>/FFY/RST ;
  wire \DLX_MEMinst_RF_data_in<15>/CKMUXNOT ;
  wire \DLX_MEMinst_RF_data_in<25>/FFY/RST ;
  wire \DLX_MEMinst_RF_data_in<25>/CKMUXNOT ;
  wire \DLX_MEMinst_RF_data_in<17>/FFY/RST ;
  wire \DLX_MEMinst_RF_data_in<17>/CKMUXNOT ;
  wire \DLX_MEMinst_RF_data_in<27>/FFY/RST ;
  wire \DLX_MEMinst_RF_data_in<27>/CKMUXNOT ;
  wire \DLX_MEMinst_RF_data_in<19>/FFY/RST ;
  wire \DLX_MEMinst_RF_data_in<19>/CKMUXNOT ;
  wire \DLX_MEMinst_RF_data_in<29>/FFY/RST ;
  wire \DLX_MEMinst_RF_data_in<29>/CKMUXNOT ;
  wire \DLX_IDinst_current_IR<11>/FFY/RST ;
  wire \DLX_IDinst_current_IR<11>/FROM ;
  wire \DLX_IDinst_current_IR<11>/GROM ;
  wire \DLX_IDinst_current_IR<20>/LOGIC_ZERO ;
  wire DLX_IDinst_Mcompar__n0315_inst_lut4_42;
  wire \DLX_IDinst_current_IR<20>/CYMUXF ;
  wire \DLX_IDinst_current_IR<20>/CYINIT ;
  wire \DLX_IDinst_current_IR<20>/GROM ;
  wire \DLX_IDinst_current_IR<13>/FROM ;
  wire \DLX_IDinst_current_IR<13>/GROM ;
  wire \DLX_IDinst_current_IR<21>/FROM ;
  wire \DLX_IDinst_current_IR<21>/GROM ;
  wire \DLX_IDinst_current_IR<15>/FROM ;
  wire \DLX_IDinst_current_IR<15>/GROM ;
  wire \DLX_IDinst_current_IR<23>/FROM ;
  wire \DLX_IDinst_current_IR<23>/GROM ;
  wire \DLX_IDinst_current_IR<30>/FROM ;
  wire \DLX_IDinst_current_IR<30>/GROM ;
  wire \DLX_IDinst_current_IR<31>/FROM ;
  wire \DLX_IDinst_current_IR<31>/GROM ;
  wire \DM_addr_eff<8>/OFF/RST ;
  wire \DLX_IDinst_current_IR<24>/FROM ;
  wire \DLX_IDinst_current_IR<24>/GROM ;
  wire \DLX_IDinst_current_IR<17>/FROM ;
  wire \DLX_IDinst_current_IR<17>/GROM ;
  wire \DLX_IDinst_current_IR<25>/LOGIC_ZERO ;
  wire DLX_IDinst_Mcompar__n0314_inst_lut4_42;
  wire \DLX_IDinst_current_IR<25>/CYMUXF ;
  wire \DLX_IDinst_current_IR<25>/CYINIT ;
  wire \DLX_IDinst_current_IR<25>/GROM ;
  wire \DLX_IDinst_current_IR<26>/FROM ;
  wire \DLX_IDinst_current_IR<26>/GROM ;
  wire \DLX_IDinst_current_IR<19>/FROM ;
  wire \DLX_IDinst_current_IR<19>/GROM ;
  wire \DLX_IDinst_current_IR<27>/FROM ;
  wire \DLX_IDinst_current_IR<27>/GROM ;
  wire \DLX_IDinst_current_IR<28>/FROM ;
  wire \DLX_IDinst_current_IR<28>/GROM ;
  wire \DLX_IDinst_current_IR<29>/FROM ;
  wire \DLX_IDinst_current_IR<29>/GROM ;
  wire \DLX_reg_dst_of_MEM<1>/FROM ;
  wire \DLX_reg_dst_of_MEM<1>/GROM ;
  wire \DLX_reg_dst_of_MEM<3>/FROM ;
  wire \DLX_reg_dst_of_MEM<3>/GROM ;
  wire \DLX_IDinst_counter<1>/FROM ;
  wire \DM_addr_eff<9>/OFF/RST ;
  wire DLX_EXinst__n0009;
  wire \DLX_EXinst_reg_write_EX/GROM ;
  wire \DLX_IDinst_IR_function_field<0>/GROM ;
  wire \DLX_EXinst_reg_out_B_EX<14>/FROM ;
  wire \DLX_IDinst_IR_function_field<1>/GROM ;
  wire \DLX_IDinst_IR_function_field<2>/GROM ;
  wire \DLX_IDinst_IR_function_field<3>/GROM ;
  wire \DLX_EXinst_ALU_result<2>/FROM ;
  wire \DLX_EXinst_ALU_result<2>/GROM ;
  wire DLX_IDinst__n0099;
  wire DLX_IDinst__n0097;
  wire DLX_IDinst__n0098;
  wire \DLX_RF_data_in<1>/CKMUXNOT ;
  wire DLX_IDinst__n0095;
  wire DLX_IDinst__n0096;
  wire \DLX_RF_data_in<3>/CKMUXNOT ;
  wire \DLX_RF_data_in<5>/CKMUXNOT ;
  wire \DLX_RF_data_in<7>/CKMUXNOT ;
  wire \DLX_MEMinst_RF_data_in<9>/CKMUXNOT ;
  wire \DLX_IDinst_IR_opcode_field<5>/FFY/RST ;
  wire DLX_EXinst__n0015;
  wire DLX_EXinst__n0014;
  wire \DLX_IDinst_intr_slot/FFY/RST ;
  wire \DLX_IDinst_intr_slot/FROM ;
  wire DLX_IDinst__n0126;
  wire \DLX_IFinst_stalled/FROM ;
  wire \DLX_IFinst_stalled/GROM ;
  wire \DLX_IFinst_stalled/CEMUXNOT ;
  wire \DLX_IDinst_rt_addr<1>/FROM ;
  wire \DLX_IDinst_mem_read/FROM ;
  wire DLX_IDinst__n0111;
  wire \DLX_IDinst_mem_write/FROM ;
  wire DLX_IDinst__n0112;
  wire \DLX_EXinst_reg_out_B_EX<1>/GROM ;
  wire \DLX_EXinst_reg_dst_out<3>/FFY/RST ;
  wire \DLX_IDinst_IR_function_field<5>/FFY/RST ;
  wire DLX_IDinst__n0101;
  wire \CHOICE3210/FROM ;
  wire \CHOICE3210/GROM ;
  wire \DLX_IDinst_reg_out_A<28>/FROM ;
  wire N104508;
  wire \DLX_IDinst_reg_out_A<5>/FROM ;
  wire N103012;
  wire \CHOICE2386/FROM ;
  wire \CHOICE2386/GROM ;
  wire \CHOICE2338/FROM ;
  wire \CHOICE2338/GROM ;
  wire \DLX_MEMlc_ridp3/FROM ;
  wire \DLX_MEMlc_ridp3/GROM ;
  wire \N93747/FROM ;
  wire \N93747/GROM ;
  wire \N127155/FROM ;
  wire \N127155/GROM ;
  wire \N126593/FROM ;
  wire \N126593/GROM ;
  wire \DLX_IDinst_reg_out_A<29>/FROM ;
  wire N104644;
  wire \DLX_EXinst_Mshift__n0023_Sh<5>/FROM ;
  wire \DLX_EXinst_Mshift__n0023_Sh<5>/GROM ;
  wire \DLX_IDinst_reg_out_A<6>/FFY/RST ;
  wire \DLX_IDinst_reg_out_A<6>/FROM ;
  wire N103148;
  wire \N127392/FROM ;
  wire \N127392/GROM ;
  wire \CHOICE2194/FROM ;
  wire \CHOICE2194/GROM ;
  wire \DLX_MEMlc_md_wint13/FROM ;
  wire \DLX_MEMlc_md_wint13/GROM ;
  wire \DLX_IDinst_reg_out_A<7>/FROM ;
  wire N103080;
  wire \CHOICE39/FROM ;
  wire \CHOICE39/GROM ;
  wire \CHOICE2422/FROM ;
  wire \CHOICE2422/GROM ;
  wire \DLX_MEMlc_md_wint12/FROM ;
  wire \DLX_MEMlc_md_wint12/GROM ;
  wire \DLX_EXinst_N66177/FROM ;
  wire \DLX_EXinst_N66177/GROM ;
  wire \N126519/FROM ;
  wire \N126519/GROM ;
  wire \DLX_EXinst_ALU_result<19>/FROM ;
  wire N119626;
  wire \DLX_reqin_IF/GROM ;
  wire \DLX_IDinst_reg_out_A<8>/FROM ;
  wire N103216;
  wire \N126297/FROM ;
  wire \N126297/GROM ;
  wire \DLX_IDinst_N70653/FROM ;
  wire \DLX_IDinst_N70653/GROM ;
  wire \CHOICE2266/FROM ;
  wire \CHOICE2266/GROM ;
  wire \N127388/FROM ;
  wire \N127388/GROM ;
  wire \DLX_MEMlc_md_wint7/FROM ;
  wire \DLX_MEMlc_md_wint7/GROM ;
  wire \DLX_IDinst_reg_out_A<9>/FROM ;
  wire N103284;
  wire \DLX_EXinst_N64062/FROM ;
  wire \DLX_EXinst_N64062/GROM ;
  wire \N107613/FROM ;
  wire \N107613/GROM ;
  wire \CHOICE3500/FROM ;
  wire \CHOICE3500/GROM ;
  wire \DLX_MEMlc_md_wint1/FROM ;
  wire \DLX_MEMlc_md_wint1/GROM ;
  wire \N93229/FROM ;
  wire \N93229/GROM ;
  wire \CHOICE45/FROM ;
  wire \CHOICE45/GROM ;
  wire \N93695/FROM ;
  wire \N93695/GROM ;
  wire \DLX_RF_delay_inst_wint10/GROM ;
  wire \CHOICE3436/FROM ;
  wire \CHOICE3436/GROM ;
  wire \vga_top_vga1_N73363/FROM ;
  wire \vga_top_vga1_N73363/GROM ;
  wire \DLX_RF_delay_inst_wint11/GROM ;
  wire \DLX_IDinst__n0421/FROM ;
  wire \DLX_IDinst__n0421/GROM ;
  wire \DLX_RF_delay_inst_wint12/GROM ;
  wire \DLX_RF_delay_inst_wint20/FROM ;
  wire \DLX_RF_delay_inst_wint20/GROM ;
  wire \vga_top_vga1_N73357/FROM ;
  wire \vga_top_vga1_N73357/GROM ;
  wire \DLX_RF_delay_inst_wint13/GROM ;
  wire \DM_delay_inst_wint1/GROM ;
  wire \vga_top_vga1_N73374/FROM ;
  wire \vga_top_vga1_N73374/GROM ;
  wire \CHOICE3444/FROM ;
  wire \CHOICE3444/GROM ;
  wire \DLX_RF_delay_inst_wint14/FROM ;
  wire \DLX_RF_delay_inst_wint14/GROM ;
  wire \DLX_RF_delay_inst_wint22/GROM ;
  wire \DLX_RF_delay_inst_wint30/GROM ;
  wire \DM_delay_inst_wint2/GROM ;
  wire \DLX_RF_delay_inst_wint23/GROM ;
  wire \DM_delay_inst_wint3/GROM ;
  wire \CHOICE3518/FROM ;
  wire \CHOICE3518/GROM ;
  wire \CHOICE3847/FROM ;
  wire \CHOICE3847/GROM ;
  wire \CHOICE3166/FROM ;
  wire \CHOICE3166/GROM ;
  wire \N102162/FROM ;
  wire \N102162/GROM ;
  wire \CHOICE1452/FROM ;
  wire \CHOICE1452/GROM ;
  wire \DLX_ackout_ID/FROM ;
  wire \DLX_ackout_ID/GROM ;
  wire \DLX_EXlc_md_wint20/FROM ;
  wire \DLX_EXlc_md_wint20/GROM ;
  wire \CHOICE5839/FROM ;
  wire \CHOICE5839/GROM ;
  wire \N98127/FROM ;
  wire \N98127/GROM ;
  wire \DLX_EXinst_Mshift__n0028_Sh<51>/FROM ;
  wire \DLX_EXinst_Mshift__n0028_Sh<51>/GROM ;
  wire \CHOICE3539/FROM ;
  wire \CHOICE3539/GROM ;
  wire \N126546/FROM ;
  wire \N126546/GROM ;
  wire \CHOICE3957/FROM ;
  wire \CHOICE3957/GROM ;
  wire \CHOICE2077/FROM ;
  wire \CHOICE2077/GROM ;
  wire \CHOICE3850/FROM ;
  wire \CHOICE3850/GROM ;
  wire \DLX_IDinst__n0445<47>/FROM ;
  wire \DLX_IDinst__n0445<47>/GROM ;
  wire \DLX_EXlc_md_wint19/FROM ;
  wire \DLX_EXlc_md_wint19/GROM ;
  wire \N102358/FROM ;
  wire \N102358/GROM ;
  wire \DLX_IDinst__n0445<40>/FROM ;
  wire \DLX_IDinst__n0445<40>/GROM ;
  wire \DLX_IDinst__n0445<41>/FROM ;
  wire \DLX_IDinst__n0445<41>/GROM ;
  wire \DLX_IDinst__n0002/FROM ;
  wire \DLX_IDinst__n0002/GROM ;
  wire \CHOICE3706/FROM ;
  wire \CHOICE3706/GROM ;
  wire \DLX_EXinst_ALU_result<7>/FROM ;
  wire \DLX_EXinst_ALU_result<7>/GROM ;
  wire \CHOICE3399/FROM ;
  wire \CHOICE3399/GROM ;
  wire \DLX_IDinst__n0445<42>/FROM ;
  wire \DLX_IDinst__n0445<42>/GROM ;
  wire \CHOICE3554/FROM ;
  wire \CHOICE3554/GROM ;
  wire \N100440/FROM ;
  wire \N100440/GROM ;
  wire \CHOICE3556/FROM ;
  wire \CHOICE3556/GROM ;
  wire \DLX_IDinst__n0445<43>/FROM ;
  wire \DLX_IDinst__n0445<43>/GROM ;
  wire \CHOICE3112/FROM ;
  wire \CHOICE3112/GROM ;
  wire \DLX_EXlc_md_wint18/FROM ;
  wire \DLX_EXlc_md_wint18/GROM ;
  wire \DLX_IDinst__n0445<44>/FROM ;
  wire \DLX_IDinst__n0445<44>/GROM ;
  wire \CHOICE3728/FROM ;
  wire \CHOICE3728/GROM ;
  wire \CHOICE3249/GROM ;
  wire \CHOICE3713/FROM ;
  wire \CHOICE3713/GROM ;
  wire \DLX_IDinst__n0445<45>/FROM ;
  wire \DLX_IDinst__n0445<45>/GROM ;
  wire \CHOICE4196/FROM ;
  wire \CHOICE4196/GROM ;
  wire \DLX_IDinst__n0445<46>/FROM ;
  wire \DLX_IDinst__n0445<46>/GROM ;
  wire \DLX_EXlc_md_wint30/FROM ;
  wire \DLX_EXlc_md_wint30/GROM ;
  wire \DLX_EXlc_md_wint17/FROM ;
  wire \DLX_EXlc_md_wint17/GROM ;
  wire \DLX_IDinst_branch_address<10>/FROM ;
  wire N105724;
  wire \N102270/FROM ;
  wire \N102270/GROM ;
  wire \N101725/FROM ;
  wire \N101725/GROM ;
  wire \DLX_EXinst_ALU_result<8>/FROM ;
  wire \DLX_EXinst_ALU_result<8>/GROM ;
  wire \CHOICE3725/FROM ;
  wire \CHOICE3725/GROM ;
  wire \CHOICE1976/FROM ;
  wire \CHOICE1976/GROM ;
  wire \CHOICE5746/FROM ;
  wire \CHOICE5746/GROM ;
  wire \DLX_RF_delay_inst_wint16/GROM ;
  wire \DLX_RF_delay_inst_wint24/FROM ;
  wire \DLX_RF_delay_inst_wint24/GROM ;
  wire \DM_delay_inst_wint4/GROM ;
  wire \DLX_MEMlc_md_wint8/FROM ;
  wire \DLX_MEMlc_md_wint8/GROM ;
  wire \DLX_RF_delay_inst_wint17/GROM ;
  wire \DM_delay_inst_wint5/GROM ;
  wire \vga_top_vga1_N73394/GROM ;
  wire \DLX_RF_delay_inst_wint18/GROM ;
  wire \DLX_RF_delay_inst_wint26/GROM ;
  wire \DM_delay_inst_wint6/GROM ;
  wire \DLX_IDinst_N70077/FROM ;
  wire \DLX_IDinst_N70077/GROM ;
  wire \DLX_RF_delay_inst_wint19/GROM ;
  wire \DLX_RF_delay_inst_wint27/GROM ;
  wire \DM_delay_inst_wint7/GROM ;
  wire \CHOICE5657/FROM ;
  wire \CHOICE5657/GROM ;
  wire \DLX_IDinst_IR_opcode_field<1>/FROM ;
  wire \DLX_RF_delay_inst_wint28/GROM ;
  wire \DM_delay_inst_wint8/GROM ;
  wire \CHOICE51/FROM ;
  wire \CHOICE51/GROM ;
  wire \DLX_RF_delay_inst_wint29/GROM ;
  wire \DM_delay_inst_wint9/GROM ;
  wire \CHOICE5411/FROM ;
  wire \CHOICE5411/GROM ;
  wire \N127139/FROM ;
  wire \N127139/GROM ;
  wire \CHOICE3525/FROM ;
  wire \CHOICE3525/GROM ;
  wire \vga_top_vga1_N73399/FROM ;
  wire \vga_top_vga1_N73399/GROM ;
  wire \CHOICE5020/FROM ;
  wire \CHOICE5020/GROM ;
  wire \N127378/FROM ;
  wire \N127378/GROM ;
  wire \DLX_IFlc_md_wint33/FROM ;
  wire \DLX_IFlc_md_wint33/GROM ;
  wire \DLX_IDinst__n0338/FROM ;
  wire \DLX_IDinst__n0338/GROM ;
  wire \DLX_IFlc_md_wint32/FROM ;
  wire \DLX_IFlc_md_wint32/GROM ;
  wire \N126847/FROM ;
  wire \N126847/GROM ;
  wire \CHOICE3317/FROM ;
  wire \CHOICE3317/GROM ;
  wire \DLX_IFinst_PC<9>/FFY/RST ;
  wire \DLX_IFlc_md_wint29/FROM ;
  wire \DLX_IFlc_md_wint29/GROM ;
  wire \DLX_IFlc_md_wint28/FROM ;
  wire \DLX_IFlc_md_wint28/GROM ;
  wire \N126580/FROM ;
  wire \N126580/GROM ;
  wire \DLX_EXinst_N63129/FROM ;
  wire \DLX_EXinst_N63129/GROM ;
  wire \DLX_IDinst_Imm_31_1/FROM ;
  wire \DLX_IDinst_Imm_31_1/GROM ;
  wire \N93383/FROM ;
  wire \N93383/GROM ;
  wire \DLX_IDinst__n0250/FROM ;
  wire \DLX_IDinst__n0250/GROM ;
  wire \DLX_EXinst_N63484/FROM ;
  wire \DLX_EXinst_N63484/GROM ;
  wire \DLX_IDinst_branch_sig/FROM ;
  wire \DLX_IDinst_branch_sig/GROM ;
  wire \DLX_IFlc_md_wint25/FROM ;
  wire \DLX_IFlc_md_wint25/GROM ;
  wire \DLX_IFlc_md_wint24/FROM ;
  wire \DLX_IFlc_md_wint24/GROM ;
  wire \DLX_EXinst__n0017<9>/FROM ;
  wire \DLX_EXinst__n0017<9>/GROM ;
  wire \CHOICE292/FROM ;
  wire \CHOICE292/GROM ;
  wire \DLX_EXinst_N62806/FROM ;
  wire \DLX_EXinst_N62806/GROM ;
  wire \CHOICE4396/FROM ;
  wire \CHOICE4396/GROM ;
  wire \DLX_IFlc_md_wint30/FROM ;
  wire \DLX_IFlc_md_wint30/GROM ;
  wire \DLX_IFlc_md_wint19/FROM ;
  wire \DLX_IFlc_md_wint19/GROM ;
  wire \DLX_IFlc_md_wint23/FROM ;
  wire \DLX_IFlc_md_wint23/GROM ;
  wire \DLX_EXinst_N62811/FROM ;
  wire \DLX_EXinst_N62811/GROM ;
  wire \DLX_EXinst_N66485/FROM ;
  wire \DLX_EXinst_N66485/GROM ;
  wire \DLX_EXinst_N63026/FROM ;
  wire \DLX_EXinst_N63026/GROM ;
  wire \CHOICE1324/FROM ;
  wire \CHOICE1324/GROM ;
  wire \DLX_EXinst_N63011/FROM ;
  wire \DLX_EXinst_N63011/GROM ;
  wire \N125959/FROM ;
  wire \N125959/GROM ;
  wire \PIPEEMPTY_OBUF/GROM ;
  wire \DLX_IFlc_md_wint18/FROM ;
  wire \DLX_IFlc_md_wint18/GROM ;
  wire \DLX_EXinst_Mshift__n0024_Sh<25>/FROM ;
  wire \DLX_EXinst_Mshift__n0024_Sh<25>/GROM ;
  wire \DLX_EXinst_ALU_result<24>/FROM ;
  wire N112254;
  wire \DLX_EXinst_N63036/FROM ;
  wire \DLX_EXinst_N63036/GROM ;
  wire \DLX_EXinst__n0017<10>/FROM ;
  wire \DLX_EXinst__n0017<10>/GROM ;
  wire \DLX_IDinst_IR_opcode_field<3>/FROM ;
  wire \DLX_EXinst_Mshift__n0024_Sh<27>/FROM ;
  wire \DLX_EXinst_Mshift__n0024_Sh<27>/GROM ;
  wire \DLX_EXinst_N63046/FROM ;
  wire \DLX_EXinst_N63046/GROM ;
  wire \DLX_EXinst__n0017<13>/FROM ;
  wire \DLX_EXinst__n0017<13>/GROM ;
  wire \DLX_IFlc_md_wint9/FROM ;
  wire \DLX_IFlc_md_wint9/GROM ;
  wire \DLX_IFlc_md_wint17/FROM ;
  wire \DLX_IFlc_md_wint17/GROM ;
  wire \DLX_EXinst_N63056/FROM ;
  wire \DLX_EXinst_N63056/GROM ;
  wire \CHOICE4990/FROM ;
  wire \CHOICE4990/GROM ;
  wire \DLX_EXinst_N63339/FROM ;
  wire \DLX_EXinst_N63339/GROM ;
  wire \DLX_EXinst__n0017<15>/FROM ;
  wire \DLX_EXinst__n0017<15>/GROM ;
  wire \DLX_EXinst_N63041/FROM ;
  wire \DLX_EXinst_N63041/GROM ;
  wire \CHOICE3917/FROM ;
  wire \CHOICE3917/GROM ;
  wire \vga_top_vga1_helpcounter<0>/BXMUXNOT ;
  wire \DLX_EXinst_N63066/FROM ;
  wire \DLX_EXinst_N63066/GROM ;
  wire \N127404/FROM ;
  wire \N127404/GROM ;
  wire \DLX_EXinst_N63404/FROM ;
  wire \DLX_EXinst_N63404/GROM ;
  wire \DLX_EXinst_N63157/GROM ;
  wire \DLX_EXinst_N63061/FROM ;
  wire \DLX_EXinst_N63061/GROM ;
  wire \DLX_EXinst_N63279/FROM ;
  wire \DLX_EXinst_N63279/GROM ;
  wire \N127322/FROM ;
  wire \N127322/GROM ;
  wire \DLX_IDinst__n0442/FROM ;
  wire \DLX_IDinst__n0442/GROM ;
  wire \DLX_EXinst_N63414/FROM ;
  wire \DLX_EXinst_N63414/GROM ;
  wire \DLX_EXinst_N62946/FROM ;
  wire \DLX_EXinst_N62946/GROM ;
  wire \N127126/FROM ;
  wire \N127126/GROM ;
  wire \DLX_IDinst_N70885/FROM ;
  wire \DLX_IDinst_N70885/GROM ;
  wire \DM_delay_inst_wint10/GROM ;
  wire \DLX_IDinst_regB_eff<1>/FROM ;
  wire \DLX_IDinst_regB_eff<1>/GROM ;
  wire \DLX_IFlc_md_wint34/FROM ;
  wire \DLX_IFlc_md_wint34/GROM ;
  wire \DLX_IFlc_md_wint26/FROM ;
  wire \DLX_IFlc_md_wint26/GROM ;
  wire \CHOICE2099/FROM ;
  wire \CHOICE2099/GROM ;
  wire \DM_delay_inst_wint11/GROM ;
  wire \DLX_EXinst_N63424/FROM ;
  wire \DLX_EXinst_N63424/GROM ;
  wire \DLX_EXinst_N64560/FROM ;
  wire \DLX_EXinst_N64560/GROM ;
  wire \DLX_EXinst_N63504/FROM ;
  wire \DLX_EXinst_N63504/GROM ;
  wire \DM_delay_inst_wint12/GROM ;
  wire \DM_delay_inst_wint20/FROM ;
  wire \DM_delay_inst_wint20/GROM ;
  wire \DLX_EXlc_slave_ctrlEX_l/GROM ;
  wire \DLX_IDinst_regB_eff<2>/FROM ;
  wire \DLX_IDinst_regB_eff<2>/GROM ;
  wire \N126811/FROM ;
  wire \N126811/GROM ;
  wire \CHOICE1321/FROM ;
  wire \CHOICE1321/GROM ;
  wire \DLX_EXinst_N63081/FROM ;
  wire \DLX_EXinst_N63081/GROM ;
  wire \DLX_EXinst_N63409/FROM ;
  wire \DLX_EXinst_N63409/GROM ;
  wire \DLX_EXinst_N63329/FROM ;
  wire \DLX_EXinst_N63329/GROM ;
  wire \CHOICE3736/FROM ;
  wire \CHOICE3736/GROM ;
  wire \DM_delay_inst_wint13/GROM ;
  wire \CHOICE1184/FROM ;
  wire \CHOICE1184/GROM ;
  wire \DLX_EXinst_N63780/FROM ;
  wire \DLX_EXinst_N63780/GROM ;
  wire \DLX_EXinst_N64314/FROM ;
  wire \DLX_EXinst_N64314/GROM ;
  wire \DLX_EXinst_N63514/FROM ;
  wire \DLX_EXinst_N63514/GROM ;
  wire \DM_delay_inst_wint14/GROM ;
  wire \DM_read/OFF/RST ;
  wire \DM_delay_inst_wint22/GROM ;
  wire \DM_delay_inst_wint30/GROM ;
  wire \DLX_IDinst_regB_eff<3>/FROM ;
  wire \DLX_IDinst_regB_eff<3>/GROM ;
  wire \DLX_IDinst_regB_eff<4>/FROM ;
  wire \DLX_IDinst_regB_eff<4>/GROM ;
  wire \DLX_EXinst_N63419/FROM ;
  wire \DLX_EXinst_N63419/GROM ;
  wire \CHOICE5244/FROM ;
  wire \CHOICE5244/GROM ;
  wire \CHOICE5333/FROM ;
  wire \CHOICE5333/GROM ;
  wire \DM_delay_inst_wint15/GROM ;
  wire \DM_delay_inst_wint23/GROM ;
  wire \DM_delay_inst_wint31/GROM ;
  wire \DLX_EXinst_N62976/FROM ;
  wire \DLX_EXinst_N62976/GROM ;
  wire \DLX_EXinst_N63364/FROM ;
  wire \DLX_EXinst_N63364/GROM ;
  wire \DLX_EXinst_N64324/FROM ;
  wire \DLX_EXinst_N64324/GROM ;
  wire \N127396/FROM ;
  wire \N127396/GROM ;
  wire \DLX_clk_IF/FROM ;
  wire \DLX_clk_IF/GROM ;
  wire \DM_delay_inst_wint16/GROM ;
  wire \DM_delay_inst_wint24/GROM ;
  wire \DM_delay_inst_wint32/GROM ;
  wire \DM_delay_inst_wint40/GROM ;
  wire \DLX_IDinst_regB_eff<5>/FROM ;
  wire \DLX_IDinst_regB_eff<5>/GROM ;
  wire \DLX_IDinst_regB_eff<6>/FROM ;
  wire \DLX_IDinst_regB_eff<6>/GROM ;
  wire \DLX_EXinst_N62733/FROM ;
  wire \DLX_EXinst_N62733/GROM ;
  wire \DLX_EXinst_N62709/FROM ;
  wire \DLX_EXinst_N62709/GROM ;
  wire \DLX_EXinst_N63269/FROM ;
  wire \DLX_EXinst_N63269/GROM ;
  wire \DLX_EXinst_N63429/FROM ;
  wire \DLX_EXinst_N63429/GROM ;
  wire \DLX_EXinst_N63509/FROM ;
  wire \DLX_EXinst_N63509/GROM ;
  wire \N126263/FROM ;
  wire \N126263/GROM ;
  wire \CHOICE4610/FROM ;
  wire \CHOICE4610/GROM ;
  wire \NPC_eff<10>/OFF/RST ;
  wire \DM_delay_inst_wint17/GROM ;
  wire \DM_delay_inst_wint25/GROM ;
  wire \DM_delay_inst_wint33/GROM ;
  wire \DLX_IDinst_rt_addr<0>/FROM ;
  wire \DLX_EXinst_N63374/FROM ;
  wire \DLX_EXinst_N63374/GROM ;
  wire \DLX_IDinst_IR_opcode_field<4>/FROM ;
  wire \DLX_EXinst_N63294/FROM ;
  wire \DLX_EXinst_N63294/GROM ;
  wire \NPC_eff<11>/OFF/RST ;
  wire \DLX_EXinst_N64334/FROM ;
  wire \DLX_EXinst_N64334/GROM ;
  wire \DLX_EXinst_N63454/FROM ;
  wire \DLX_EXinst_N63454/GROM ;
  wire \DLX_EXinst_N64094/FROM ;
  wire \DLX_EXinst_N64094/GROM ;
  wire \N127314/FROM ;
  wire \N127314/GROM ;
  wire \DM_delay_inst_wint18/GROM ;
  wire \DM_delay_inst_wint26/FROM ;
  wire \DM_delay_inst_wint26/GROM ;
  wire \DM_delay_inst_wint34/FROM ;
  wire \DM_delay_inst_wint34/GROM ;
  wire \CHOICE5864/FROM ;
  wire \CHOICE5864/GROM ;
  wire \DLX_IDinst_regB_eff<7>/FROM ;
  wire \DLX_IDinst_regB_eff<7>/GROM ;
  wire \DLX_IDinst_regB_eff<8>/FROM ;
  wire \DLX_IDinst_regB_eff<8>/GROM ;
  wire \DLX_IDinst_regB_eff<9>/FROM ;
  wire \DLX_IDinst_regB_eff<9>/GROM ;
  wire \DLX_IFlc_md_wint8/FROM ;
  wire \DLX_IFlc_md_wint8/GROM ;
  wire \DLX_EXinst_N62631/FROM ;
  wire \DLX_EXinst_N62631/GROM ;
  wire \N94155/FROM ;
  wire \N94155/GROM ;
  wire \DLX_EXinst_N63359/FROM ;
  wire \DLX_EXinst_N63359/GROM ;
  wire \DLX_EXinst_N63474/FROM ;
  wire \DLX_EXinst_N63474/GROM ;
  wire \DLX_EXinst_N64319/FROM ;
  wire \DLX_EXinst_N64319/GROM ;
  wire \NPC_eff<12>/OFF/RST ;
  wire \N94305/FROM ;
  wire \N94305/GROM ;
  wire \DLX_EXinst_N63439/FROM ;
  wire \DLX_EXinst_N63439/GROM ;
  wire \N57312/FROM ;
  wire \N57312/GROM ;
  wire \DLX_IFlc_md_wint7/FROM ;
  wire \DLX_IFlc_md_wint7/GROM ;
  wire \DM_delay_inst_wint19/GROM ;
  wire \DLX_EXinst_N66112/FROM ;
  wire \DLX_EXinst_N66112/GROM ;
  wire \DLX_EXinst_N63384/FROM ;
  wire \DLX_EXinst_N63384/GROM ;
  wire \DLX_EXinst_N63464/FROM ;
  wire \DLX_EXinst_N63464/GROM ;
  wire \DM_delay_inst_wint28/GROM ;
  wire \DM_delay_inst_wint36/GROM ;
  wire \reset_IBUF_1/FROM ;
  wire \reset_IBUF_1/GROM ;
  wire \DLX_IDinst_regB_eff<16>/FROM ;
  wire \DLX_IDinst_regB_eff<16>/GROM ;
  wire \DLX_IDinst_regB_eff<17>/FROM ;
  wire \DLX_IDinst_regB_eff<17>/GROM ;
  wire \DLX_IDinst_regB_eff<18>/FROM ;
  wire \DLX_IDinst_regB_eff<18>/GROM ;
  wire \DLX_EXinst_N63369/FROM ;
  wire \DLX_EXinst_N63369/GROM ;
  wire \DLX_EXinst_N66105/FROM ;
  wire \DLX_EXinst_N66105/GROM ;
  wire \DLX_EXinst_N62721/FROM ;
  wire \DLX_EXinst_N62721/GROM ;
  wire \NPC_eff<13>/OFF/RST ;
  wire \DLX_EXinst_N63449/FROM ;
  wire \DLX_EXinst_N63449/GROM ;
  wire \DLX_EXinst_N64329/FROM ;
  wire \DLX_EXinst_N64329/GROM ;
  wire \reset_IBUF_2/GROM ;
  wire \CHOICE5408/FROM ;
  wire \CHOICE5408/GROM ;
  wire \CHOICE4675/FROM ;
  wire \CHOICE4675/GROM ;
  wire \DM_delay_inst_wint29/GROM ;
  wire \DM_delay_inst_wint37/GROM ;
  wire \reset_IBUF_3/GROM ;
  wire \DLX_EXinst_N66202/FROM ;
  wire \DLX_EXinst_N66202/GROM ;
  wire \reset_IBUF_4/GROM ;
  wire \DM_delay_inst_wint38/GROM ;
  wire \reset_IBUF_5/GROM ;
  wire \DLX_IDinst_regB_eff<19>/FROM ;
  wire \DLX_IDinst_regB_eff<19>/GROM ;
  wire \DLX_IFlc_md_wint6/FROM ;
  wire \DLX_IFlc_md_wint6/GROM ;
  wire \DLX_EXinst_N63379/FROM ;
  wire \DLX_EXinst_N63379/GROM ;
  wire \CHOICE3836/FROM ;
  wire \CHOICE3836/GROM ;
  wire \DLX_EXinst_N63459/FROM ;
  wire \DLX_EXinst_N63459/GROM ;
  wire \NPC_eff<14>/OFF/RST ;
  wire \CHOICE3818/FROM ;
  wire \CHOICE3818/GROM ;
  wire \DLX_IFlc_md_wint5/FROM ;
  wire \DLX_IFlc_md_wint5/GROM ;
  wire \DM_delay_inst_wint39/GROM ;
  wire \DLX_EXinst_N62740/FROM ;
  wire \DLX_EXinst_N62740/GROM ;
  wire \CHOICE3692/FROM ;
  wire \CHOICE3692/GROM ;
  wire \DLX_IDinst_regB_eff<26>/FROM ;
  wire \DLX_IDinst_regB_eff<26>/GROM ;
  wire \DLX_EXinst_N62821/FROM ;
  wire \DLX_EXinst_N62821/GROM ;
  wire \CHOICE1294/FROM ;
  wire \CHOICE1294/GROM ;
  wire \DLX_EXinst_N63469/FROM ;
  wire \DLX_EXinst_N63469/GROM ;
  wire \DLX_EXinst_N63389/FROM ;
  wire \DLX_EXinst_N63389/GROM ;
  wire \CHOICE5256/FROM ;
  wire \CHOICE5256/GROM ;
  wire \DLX_EXinst_N62766/FROM ;
  wire \DLX_EXinst_N62766/GROM ;
  wire \DLX_EXinst_N63494/FROM ;
  wire \DLX_EXinst_N63494/GROM ;
  wire \DLX_IFlc_md_wint38/FROM ;
  wire \DLX_IFlc_md_wint38/GROM ;
  wire \DLX_EXinst_N64587/FROM ;
  wire \DLX_EXinst_N64587/GROM ;
  wire \CHOICE4438/FROM ;
  wire \CHOICE4438/GROM ;
  wire \DLX_EXinst_N64550/FROM ;
  wire \DLX_EXinst_N64550/GROM ;
  wire \DLX_EXinst_N62856/FROM ;
  wire \DLX_EXinst_N62856/GROM ;
  wire \DLX_EXinst_N62921/FROM ;
  wire \DLX_EXinst_N62921/GROM ;
  wire \N94255/FROM ;
  wire \N94255/GROM ;
  wire \DLX_IDinst_regB_eff<28>/FROM ;
  wire \DLX_IDinst_regB_eff<28>/GROM ;
  wire \N95468/FROM ;
  wire \N95468/GROM ;
  wire \CHOICE1446/FROM ;
  wire \CHOICE1446/GROM ;
  wire \DLX_IDlc_md_wint4/FROM ;
  wire \DLX_IDlc_md_wint4/GROM ;
  wire \DLX_IDinst_reg_out_A<10>/FROM ;
  wire N103352;
  wire \CHOICE2446/FROM ;
  wire \CHOICE2446/GROM ;
  wire \CHOICE2924/FROM ;
  wire \CHOICE2924/GROM ;
  wire \DLX_EXinst_Mshift__n0027_Sh<6>/FROM ;
  wire \DLX_EXinst_Mshift__n0027_Sh<6>/GROM ;
  wire \DLX_EXinst_Mshift__n0024_Sh<61>/FROM ;
  wire \DLX_EXinst_Mshift__n0024_Sh<61>/GROM ;
  wire \DLX_EXinst_Mshift__n0024_Sh<29>/FROM ;
  wire \DLX_EXinst_Mshift__n0024_Sh<29>/GROM ;
  wire \DLX_IDlc_md_wint2/GROM ;
  wire \DLX_EXinst_Mshift__n0028_Sh<50>/FROM ;
  wire \DLX_EXinst_Mshift__n0028_Sh<50>/GROM ;
  wire \DLX_EXinst_Mshift__n0028_Sh<18>/FROM ;
  wire \DLX_EXinst_Mshift__n0028_Sh<18>/GROM ;
  wire \DLX_IDinst_reg_out_A<11>/FROM ;
  wire N103488;
  wire \CHOICE2326/FROM ;
  wire \CHOICE2326/GROM ;
  wire \N127257/FROM ;
  wire \N127257/GROM ;
  wire \N107780/FROM ;
  wire \N107780/GROM ;
  wire \DLX_IDlc_md_wint3/GROM ;
  wire \DLX_EXinst_Mshift__n0024_Sh<80>/GROM ;
  wire \DLX_IDinst_reg_out_A<12>/FROM ;
  wire N103420;
  wire \DLX_IDinst_reg_out_A<20>/FROM ;
  wire N104032;
  wire \CHOICE3406/FROM ;
  wire \CHOICE3406/GROM ;
  wire \CHOICE1424/FROM ;
  wire \CHOICE1424/GROM ;
  wire \CHOICE2494/FROM ;
  wire \CHOICE2494/GROM ;
  wire \DLX_IFlc_pd_wint1/FROM ;
  wire \DLX_IFlc_pd_wint1/GROM ;
  wire \N126205/FROM ;
  wire \N126205/GROM ;
  wire \N93587/FROM ;
  wire \N93587/GROM ;
  wire \DLX_IDinst_reg_out_A<21>/FROM ;
  wire N104168;
  wire \DLX_IDinst_reg_out_A<13>/FROM ;
  wire N103556;
  wire \CHOICE2170/FROM ;
  wire \CHOICE2170/GROM ;
  wire \N126816/FROM ;
  wire \N126816/GROM ;
  wire \DLX_IDinst_reg_out_A<22>/FROM ;
  wire N104100;
  wire \DLX_IDinst_reg_out_A<14>/FROM ;
  wire N103624;
  wire \DLX_IDinst_reg_out_A<30>/FROM ;
  wire N104712;
  wire \DLX_EXinst_N62966/FROM ;
  wire \DLX_EXinst_N62966/GROM ;
  wire \DLX_EXinst_N63489/FROM ;
  wire \DLX_EXinst_N63489/GROM ;
  wire \DLX_EXinst_N62866/FROM ;
  wire \DLX_EXinst_N62866/GROM ;
  wire \DLX_EXinst_N62786/FROM ;
  wire \DLX_EXinst_N62786/GROM ;
  wire \CHOICE1018/FROM ;
  wire \CHOICE1018/GROM ;
  wire \DLX_EXinst_N64914/FROM ;
  wire \DLX_EXinst_N64914/GROM ;
  wire \NPC_eff<15>/OFF/RST ;
  wire \DLX_EXinst_N66130/FROM ;
  wire \DLX_EXinst_N66130/GROM ;
  wire \DLX_IDinst_Mmux__n0148__net123/GROM ;
  wire \N126134/FROM ;
  wire \N126134/GROM ;
  wire \DLX_IFlc_md_wint39/FROM ;
  wire \DLX_IFlc_md_wint39/GROM ;
  wire \DLX_EXinst_N62851/FROM ;
  wire \DLX_EXinst_N62851/GROM ;
  wire \DLX_EXinst_N63785/FROM ;
  wire \DLX_EXinst_N63785/GROM ;
  wire \DLX_EXinst_N63499/FROM ;
  wire \DLX_EXinst_N63499/GROM ;
  wire \CHOICE4554/FROM ;
  wire \CHOICE4554/GROM ;
  wire \CHOICE3978/FROM ;
  wire \CHOICE3978/GROM ;
  wire \vga_top_vga1__n0010/FROM ;
  wire \vga_top_vga1__n0010/GROM ;
  wire \DLX_EXinst_N62876/FROM ;
  wire \DLX_EXinst_N62876/GROM ;
  wire \DLX_EXinst_N62796/FROM ;
  wire \DLX_EXinst_N62796/GROM ;
  wire \CHOICE1364/FROM ;
  wire \CHOICE1364/GROM ;
  wire \CHOICE4567/FROM ;
  wire \CHOICE4567/GROM ;
  wire \DLX_EXinst__n0017<12>/FROM ;
  wire \DLX_EXinst__n0017<12>/GROM ;
  wire \DLX_IDinst_WB_data_eff<29>/FROM ;
  wire \DLX_IDinst_WB_data_eff<29>/GROM ;
  wire \DLX_EXinst_N62861/FROM ;
  wire \DLX_EXinst_N62861/GROM ;
  wire \N127334/FROM ;
  wire \N127334/GROM ;
  wire \CHOICE5216/FROM ;
  wire \CHOICE5216/GROM ;
  wire \DLX_EXinst_N64565/FROM ;
  wire \DLX_EXinst_N64565/GROM ;
  wire \DM_write_data<0>/OFF/RST ;
  wire \CHOICE1060/FROM ;
  wire \CHOICE1060/GROM ;
  wire \DLX_EXinst_N62886/FROM ;
  wire \DLX_EXinst_N62886/GROM ;
  wire \DLX_EXinst_N64067/FROM ;
  wire \DLX_EXinst_N64067/GROM ;
  wire \DLX_EXinst_N66078/FROM ;
  wire \DLX_EXinst_N66078/GROM ;
  wire \N127107/FROM ;
  wire \N127107/GROM ;
  wire \DLX_EXinst_N64864/FROM ;
  wire \DLX_EXinst_N64864/GROM ;
  wire \DLX_EXinst_N62951/FROM ;
  wire \DLX_EXinst_N62951/GROM ;
  wire \DLX_EXinst_N62871/FROM ;
  wire \DLX_EXinst_N62871/GROM ;
  wire \DLX_EXinst_N62791/FROM ;
  wire \DLX_EXinst_N62791/GROM ;
  wire \DLX_EXinst_N66087/FROM ;
  wire \DLX_EXinst_N66087/GROM ;
  wire \DLX_EXinst_N64904/FROM ;
  wire \DLX_EXinst_N64904/GROM ;
  wire \DLX_EXinst_N62891/FROM ;
  wire \DLX_EXinst_N62891/GROM ;
  wire \DLX_EXinst_N66096/FROM ;
  wire \DLX_EXinst_N66096/GROM ;
  wire \CHOICE1359/FROM ;
  wire \CHOICE1359/GROM ;
  wire \DLX_EXinst_N63915/FROM ;
  wire \DLX_EXinst_N63915/GROM ;
  wire \CHOICE4504/FROM ;
  wire \CHOICE4504/GROM ;
  wire \DLX_EXinst_N62881/FROM ;
  wire \DLX_EXinst_N62881/GROM ;
  wire \DLX_EXinst_N62801/FROM ;
  wire \DLX_EXinst_N62801/GROM ;
  wire \CHOICE1084/FROM ;
  wire \CHOICE1084/GROM ;
  wire \DLX_EXinst_N62986/FROM ;
  wire \DLX_EXinst_N62986/GROM ;
  wire \CHOICE3992/FROM ;
  wire \CHOICE3992/GROM ;
  wire \N127306/FROM ;
  wire \N127306/GROM ;
  wire \CHOICE3674/FROM ;
  wire \CHOICE3674/GROM ;
  wire \N95300/FROM ;
  wire \N95300/GROM ;
  wire \DLX_EXinst_N62971/FROM ;
  wire \DLX_EXinst_N62971/GROM ;
  wire \N89980/FROM ;
  wire \N89980/GROM ;
  wire \DLX_EXinst_Mshift__n0025_Sh<4>/FROM ;
  wire \DLX_EXinst_Mshift__n0025_Sh<4>/GROM ;
  wire \CHOICE4429/FROM ;
  wire \CHOICE4429/GROM ;
  wire \DLX_EXinst_N62996/FROM ;
  wire \DLX_EXinst_N62996/GROM ;
  wire \DLX_EXinst_ALU_result<21>/FROM ;
  wire N114850;
  wire \DLX_IDinst_zflag/FROM ;
  wire \DLX_IDinst_zflag/GROM ;
  wire \DLX_EXinst__n0082/FROM ;
  wire \DLX_EXinst__n0082/GROM ;
  wire \DLX_EXinst_N62981/FROM ;
  wire \DLX_EXinst_N62981/GROM ;
  wire \DLX_EXinst_N66421/FROM ;
  wire \DLX_EXinst_N66421/GROM ;
  wire \DLX_EXinst_N66525/FROM ;
  wire \DLX_EXinst_N66525/GROM ;
  wire \DLX_EXinst_N66437/FROM ;
  wire \DLX_EXinst_N66437/GROM ;
  wire \CHOICE1012/FROM ;
  wire \CHOICE1012/GROM ;
  wire \CHOICE3802/FROM ;
  wire \CHOICE3802/GROM ;
  wire \N90461/FROM ;
  wire \N90461/GROM ;
  wire \DLX_EXinst_N63790/FROM ;
  wire \DLX_EXinst_N63790/GROM ;
  wire \DLX_EXinst_reg_out_B_EX<15>/FROM ;
  wire \CHOICE1072/FROM ;
  wire \CHOICE1072/GROM ;
  wire \N90557/FROM ;
  wire \N90557/GROM ;
  wire \DLX_EXinst_N62991/FROM ;
  wire \DLX_EXinst_N62991/GROM ;
  wire \DLX_EXinst_N66535/FROM ;
  wire \DLX_EXinst_N66535/GROM ;
  wire \DLX_EXinst_reg_out_B_EX<31>/FROM ;
  wire \CHOICE5223/FROM ;
  wire \CHOICE5223/GROM ;
  wire \DLX_EXinst_Mshift__n0025_Sh<5>/GROM ;
  wire \DLX_EXinst__n0061/FROM ;
  wire \DLX_EXinst__n0061/GROM ;
  wire \CHOICE3812/FROM ;
  wire \CHOICE3812/GROM ;
  wire \CHOICE4361/FROM ;
  wire \CHOICE4361/GROM ;
  wire \DLX_EXinst__n0114/FROM ;
  wire \DLX_EXinst__n0114/GROM ;
  wire \DLX_EXinst_N66392/FROM ;
  wire \DLX_EXinst_N66392/GROM ;
  wire \DLX_EXinst_N63001/FROM ;
  wire \DLX_EXinst_N63001/GROM ;
  wire \CHOICE1300/FROM ;
  wire \CHOICE1300/GROM ;
  wire \CHOICE3610/FROM ;
  wire \CHOICE3610/GROM ;
  wire \CHOICE4492/FROM ;
  wire \CHOICE4492/GROM ;
  wire \CHOICE2075/FROM ;
  wire \CHOICE2075/GROM ;
  wire \DLX_EXinst_Mshift__n0025_Sh<6>/GROM ;
  wire \CHOICE3809/FROM ;
  wire \CHOICE3809/GROM ;
  wire \CHOICE4599/FROM ;
  wire \CHOICE4599/GROM ;
  wire \DLX_EXinst__n0046/FROM ;
  wire \DLX_EXinst__n0046/GROM ;
  wire \CHOICE4119/FROM ;
  wire \CHOICE4119/GROM ;
  wire \N127412/FROM ;
  wire \N127412/GROM ;
  wire \DLX_EXinst__n0048/FROM ;
  wire \DLX_EXinst__n0048/GROM ;
  wire \N90344/FROM ;
  wire \N90344/GROM ;
  wire \DLX_EXinst__n0049/FROM ;
  wire \DLX_EXinst__n0049/GROM ;
  wire \DLX_EXinst__n0081/FROM ;
  wire \DLX_EXinst__n0081/GROM ;
  wire \vga_top_vga1_helpme/LOGIC_ZERO ;
  wire \CHOICE3691/FROM ;
  wire \CHOICE3691/GROM ;
  wire \DLX_IFinst_PC<13>/FFY/RST ;
  wire \DLX_IFinst_PC<23>/FFY/RST ;
  wire \DLX_IFinst_PC<15>/FFY/RST ;
  wire \CHOICE2558/FROM ;
  wire \CHOICE2558/GROM ;
  wire \CHOICE3603/FROM ;
  wire \CHOICE3603/GROM ;
  wire \CHOICE4560/FROM ;
  wire \CHOICE4560/GROM ;
  wire \DLX_IFinst_PC<17>/FFY/RST ;
  wire \CHOICE3876/FROM ;
  wire \CHOICE3876/GROM ;
  wire \DLX_IDinst_slot_num_FFd2/FROM ;
  wire \DLX_IDinst_slot_num_FFd2-In ;
  wire \DLX_EXinst__n0077/FROM ;
  wire \DLX_EXinst__n0077/GROM ;
  wire \DLX_IFinst_PC<19>/FFY/RST ;
  wire \CHOICE2635/FROM ;
  wire \CHOICE2635/GROM ;
  wire \CHOICE2877/FROM ;
  wire \CHOICE2877/GROM ;
  wire \DLX_EXinst__n0017<24>/FROM ;
  wire \DLX_EXinst__n0017<24>/GROM ;
  wire \DLX_IDinst__n0331/FROM ;
  wire \DLX_IDinst__n0331/GROM ;
  wire \DLX_EXinst__n0078/FROM ;
  wire \DLX_EXinst__n0078/GROM ;
  wire \DLX_IDinst__n0443/FROM ;
  wire \DLX_IDinst__n0443/GROM ;
  wire \CHOICE283/FROM ;
  wire \CHOICE283/GROM ;
  wire \DLX_IDinst__n0440/FROM ;
  wire \DLX_IDinst__n0440/GROM ;
  wire \DLX_EXinst__n0079/FROM ;
  wire \DLX_EXinst__n0079/GROM ;
  wire \CHOICE2712/FROM ;
  wire \CHOICE2712/GROM ;
  wire \CHOICE2756/FROM ;
  wire \CHOICE2756/GROM ;
  wire \DLX_EXinst__n0017<22>/FROM ;
  wire \DLX_EXinst__n0017<22>/GROM ;
  wire \N95654/FROM ;
  wire \N95654/GROM ;
  wire \N95611/FROM ;
  wire \N95611/GROM ;
  wire \CHOICE4954/FROM ;
  wire \CHOICE4954/GROM ;
  wire \CHOICE2811/FROM ;
  wire \CHOICE2811/GROM ;
  wire \CHOICE2657/FROM ;
  wire \CHOICE2657/GROM ;
  wire \DLX_EXinst__n0017<17>/FROM ;
  wire \DLX_EXinst__n0017<17>/GROM ;
  wire \CHOICE4508/FROM ;
  wire \CHOICE4508/GROM ;
  wire \blue_2_OBUF/FROM ;
  wire \blue_2_OBUF/GROM ;
  wire \CHOICE2569/FROM ;
  wire \CHOICE2569/GROM ;
  wire \DLX_EXinst__n0017<18>/FROM ;
  wire \DLX_EXinst__n0017<18>/GROM ;
  wire \DLX_EXinst__n0017<28>/FROM ;
  wire \DLX_EXinst__n0017<28>/GROM ;
  wire \DLX_EXinst_Mshift__n0025_Sh<1>/FROM ;
  wire \DLX_EXinst_Mshift__n0025_Sh<1>/GROM ;
  wire \DLX_IDinst_branch_address<0>/FROM ;
  wire N105098;
  wire \CHOICE2591/FROM ;
  wire \CHOICE2591/GROM ;
  wire \CHOICE2888/FROM ;
  wire \CHOICE2888/GROM ;
  wire \DLX_EXinst_ALU_result<17>/FROM ;
  wire N123529;
  wire \DLX_EXinst_ALU_result<25>/FROM ;
  wire N118327;
  wire \blue_1_OBUF/FROM ;
  wire \blue_1_OBUF/GROM ;
  wire \DLX_reqout_EX/GROM ;
  wire \CHOICE2580/FROM ;
  wire \CHOICE2580/GROM ;
  wire \CHOICE2899/FROM ;
  wire \CHOICE2899/GROM ;
  wire \DLX_EXinst__n0017<27>/FROM ;
  wire \DLX_EXinst__n0017<27>/GROM ;
  wire \CHOICE3412/FROM ;
  wire \CHOICE3412/GROM ;
  wire \DLX_IDinst_branch_address<1>/FROM ;
  wire N105224;
  wire \CHOICE2602/FROM ;
  wire \CHOICE2602/GROM ;
  wire \CHOICE2613/FROM ;
  wire \CHOICE2613/GROM ;
  wire \DLX_EXinst__n0017<29>/FROM ;
  wire \DLX_EXinst__n0017<29>/GROM ;
  wire \N125999/FROM ;
  wire \N125999/GROM ;
  wire \DLX_IDinst_branch_address<2>/FROM ;
  wire N105161;
  wire \CHOICE1410/FROM ;
  wire \CHOICE1410/GROM ;
  wire \N126597/FROM ;
  wire \N126597/GROM ;
  wire \CHOICE2881/FROM ;
  wire \CHOICE2881/GROM ;
  wire \N98420/FROM ;
  wire \N98420/GROM ;
  wire \DLX_IDinst_N70333/GROM ;
  wire \DLX_IDinst_branch_address<3>/FROM ;
  wire N105287;
  wire \DLX_IDinst_N70328/FROM ;
  wire \DLX_IDinst_N70328/GROM ;
  wire \DLX_IDinst_branch_address<4>/FROM ;
  wire N105350;
  wire \N100688/FROM ;
  wire \N100688/GROM ;
  wire \DLX_IDinst_branch_address<5>/FROM ;
  wire N105413;
  wire \DLX_IDinst_N70623/FROM ;
  wire \DLX_IDinst_N70623/GROM ;
  wire \DLX_IDinst_branch_address<6>/FROM ;
  wire N105535;
  wire \DLX_IDinst_branch_address<7>/FROM ;
  wire N105474;
  wire \DLX_IDinst__n0252/FROM ;
  wire \DLX_IDinst__n0252/GROM ;
  wire \DLX_IDinst_N70716/FROM ;
  wire \DLX_IDinst_N70716/GROM ;
  wire \N127366/FROM ;
  wire \N127366/GROM ;
  wire \N127362/FROM ;
  wire \N127362/GROM ;
  wire \N90497/FROM ;
  wire \N90497/GROM ;
  wire \CHOICE1479/FROM ;
  wire \CHOICE1479/GROM ;
  wire \CHOICE1757/FROM ;
  wire \CHOICE1757/GROM ;
  wire \DLX_IDinst_regA_eff<0>/FROM ;
  wire \DLX_IDinst_regA_eff<0>/GROM ;
  wire \DLX_IDinst_regA_eff<1>/FROM ;
  wire \DLX_IDinst_regA_eff<1>/GROM ;
  wire \DLX_IDinst_N70673/FROM ;
  wire \DLX_IDinst_N70673/GROM ;
  wire \DLX_IDinst_branch_address<8>/FROM ;
  wire N105598;
  wire \DLX_IDinst_N70570/FROM ;
  wire \DLX_IDinst_N70570/GROM ;
  wire \CHOICE4498/FROM ;
  wire \CHOICE4498/GROM ;
  wire \DLX_IDinst_regA_eff<2>/FROM ;
  wire \DLX_IDinst_regA_eff<2>/GROM ;
  wire \CHOICE4248/FROM ;
  wire \CHOICE4248/GROM ;
  wire \DLX_IDinst_regA_eff<3>/FROM ;
  wire \DLX_IDinst_regA_eff<3>/GROM ;
  wire \DLX_IDinst_branch_address<9>/FROM ;
  wire N105661;
  wire \DLX_IDinst_rd_addr<0>/FROM ;
  wire \CHOICE3928/FROM ;
  wire \CHOICE3928/GROM ;
  wire \DLX_IDinst_regA_eff<4>/FROM ;
  wire \DLX_IDinst_regA_eff<4>/GROM ;
  wire \DLX_EXinst_Mshift__n0023_Sh<127>/FROM ;
  wire \DLX_EXinst_Mshift__n0023_Sh<127>/GROM ;
  wire \CHOICE5047/FROM ;
  wire \CHOICE5047/GROM ;
  wire \CHOICE4185/FROM ;
  wire \CHOICE4185/GROM ;
  wire \DLX_IDinst_regA_eff<5>/FROM ;
  wire \DLX_IDinst_regA_eff<5>/GROM ;
  wire \N90656/FROM ;
  wire \N90656/GROM ;
  wire \N109741/FROM ;
  wire \N109741/GROM ;
  wire \DLX_IDinst_N70786/FROM ;
  wire \DLX_IDinst_N70786/GROM ;
  wire \CHOICE1444/FROM ;
  wire \CHOICE1444/GROM ;
  wire \CHOICE4234/FROM ;
  wire \CHOICE4234/GROM ;
  wire \N126419/FROM ;
  wire \N126419/GROM ;
  wire \CHOICE4621/FROM ;
  wire \CHOICE4621/GROM ;
  wire \DLX_IDinst_regA_eff<6>/FROM ;
  wire \DLX_IDinst_regA_eff<6>/GROM ;
  wire \DLX_EXinst__n0063/FROM ;
  wire \DLX_EXinst__n0063/GROM ;
  wire \N126239/FROM ;
  wire \N126239/GROM ;
  wire \CHOICE4611/FROM ;
  wire \CHOICE4611/GROM ;
  wire \N127354/FROM ;
  wire \N127354/GROM ;
  wire \CHOICE3877/FROM ;
  wire \CHOICE3877/GROM ;
  wire \CHOICE4676/FROM ;
  wire \CHOICE4676/GROM ;
  wire \CHOICE3755/FROM ;
  wire \CHOICE3755/GROM ;
  wire \DLX_IDinst_regA_eff<7>/FROM ;
  wire \DLX_IDinst_regA_eff<7>/GROM ;
  wire \DLX_IDinst_delay_slot/FROM ;
  wire N109531;
  wire \CHOICE4242/FROM ;
  wire \CHOICE4242/GROM ;
  wire \N100282/FROM ;
  wire \N100282/GROM ;
  wire \CHOICE4741/FROM ;
  wire \CHOICE4741/GROM ;
  wire \CHOICE4884/FROM ;
  wire \CHOICE4884/GROM ;
  wire \DLX_IDinst_regA_eff<8>/FROM ;
  wire \DLX_IDinst_regA_eff<8>/GROM ;
  wire \CHOICE4173/FROM ;
  wire \CHOICE4173/GROM ;
  wire \CHOICE4241/FROM ;
  wire \CHOICE4241/GROM ;
  wire \CHOICE5421/FROM ;
  wire \CHOICE5421/GROM ;
  wire \DLX_IDinst_regA_eff<9>/FROM ;
  wire \DLX_IDinst_regA_eff<9>/GROM ;
  wire \DLX_IDinst_N70985/FROM ;
  wire \DLX_IDinst_N70985/GROM ;
  wire \CHOICE4309/FROM ;
  wire \CHOICE4309/GROM ;
  wire \CHOICE4686/FROM ;
  wire \CHOICE4686/GROM ;
  wire \CHOICE4811/FROM ;
  wire \CHOICE4811/GROM ;
  wire \CHOICE4107/FROM ;
  wire \CHOICE4107/GROM ;
  wire \CHOICE5341/FROM ;
  wire \CHOICE5341/GROM ;
  wire \CHOICE4249/FROM ;
  wire \CHOICE4249/GROM ;
  wire \CHOICE19/FROM ;
  wire \CHOICE19/GROM ;
  wire \DLX_EXlc_md_wint33/FROM ;
  wire \DLX_EXlc_md_wint33/GROM ;
  wire \CHOICE4021/FROM ;
  wire \CHOICE4021/GROM ;
  wire \CHOICE4817/FROM ;
  wire \CHOICE4817/GROM ;
  wire \DLX_IDinst_N70991/FROM ;
  wire \DLX_IDinst_N70991/GROM ;
  wire \N126482/FROM ;
  wire \N126482/GROM ;
  wire \CHOICE5617/FROM ;
  wire \CHOICE5617/GROM ;
  wire \CHOICE4041/FROM ;
  wire \CHOICE4041/GROM ;
  wire \N126054/FROM ;
  wire \N126054/GROM ;
  wire \CHOICE2548/FROM ;
  wire \CHOICE2548/GROM ;
  wire \CHOICE3743/FROM ;
  wire \CHOICE3743/GROM ;
  wire \DLX_EXlc_ridp3/FROM ;
  wire \DLX_EXlc_ridp3/GROM ;
  wire \CHOICE5875/FROM ;
  wire \CHOICE5875/GROM ;
  wire \CHOICE5276/FROM ;
  wire \CHOICE5276/GROM ;
  wire \CHOICE3085/FROM ;
  wire \CHOICE3085/GROM ;
  wire \DLX_IDinst__n03641_1/FROM ;
  wire \DLX_IDinst__n03641_1/GROM ;
  wire \DLX_IDinst_Imm<11>/FROM ;
  wire DLX_IDinst__n0094;
  wire \CHOICE5917/FROM ;
  wire \CHOICE5917/GROM ;
  wire \CHOICE3068/FROM ;
  wire \CHOICE3068/GROM ;
  wire \CHOICE5046/FROM ;
  wire \CHOICE5046/GROM ;
  wire \CHOICE4751/FROM ;
  wire \CHOICE4751/GROM ;
  wire \CHOICE2060/FROM ;
  wire \CHOICE2060/GROM ;
  wire \CHOICE5587/FROM ;
  wire \CHOICE5587/GROM ;
  wire \DLX_IDinst_Imm<12>/FROM ;
  wire DLX_IDinst__n0093;
  wire \DLX_IDinst_Imm<5>/FROM ;
  wire DLX_IDinst__n0100;
  wire \CHOICE1138/FROM ;
  wire \CHOICE1138/GROM ;
  wire \DLX_MEMlc_pd_wint1/FROM ;
  wire \DLX_MEMlc_pd_wint1/GROM ;
  wire \CHOICE4980/FROM ;
  wire \CHOICE4980/GROM ;
  wire \CHOICE1868/FROM ;
  wire \CHOICE1868/GROM ;
  wire \DLX_EXlc_md_wint32/FROM ;
  wire \DLX_EXlc_md_wint32/GROM ;
  wire \CHOICE5953/FROM ;
  wire \CHOICE5953/GROM ;
  wire \CHOICE1957/FROM ;
  wire \CHOICE1957/GROM ;
  wire \DLX_IDinst_Imm<13>/FROM ;
  wire DLX_IDinst__n0092;
  wire \CHOICE5704/FROM ;
  wire \CHOICE5704/GROM ;
  wire \CHOICE4123/FROM ;
  wire \CHOICE4123/GROM ;
  wire \CHOICE4758/FROM ;
  wire \CHOICE4758/GROM ;
  wire \CHOICE5914/FROM ;
  wire \CHOICE5914/GROM ;
  wire \CHOICE1825/FROM ;
  wire \CHOICE1825/GROM ;
  wire \DLX_IDinst_Imm<14>/FROM ;
  wire DLX_IDinst__n0091;
  wire \CHOICE5517/FROM ;
  wire \CHOICE5517/GROM ;
  wire \N101641/FROM ;
  wire \N101641/GROM ;
  wire \CHOICE2046/FROM ;
  wire \CHOICE2046/GROM ;
  wire \DLX_EXinst_Mshift__n0023_Sh<25>/FROM ;
  wire \DLX_EXinst_Mshift__n0023_Sh<25>/GROM ;
  wire \DLX_EXlc_md_wint29/FROM ;
  wire \DLX_EXlc_md_wint29/GROM ;
  wire \DLX_EXinst_Mshift__n0026_Sh<24>/FROM ;
  wire \DLX_EXinst_Mshift__n0026_Sh<24>/GROM ;
  wire \CHOICE5686/FROM ;
  wire \CHOICE5686/GROM ;
  wire \DLX_EXinst_Mshift__n0023_Sh<29>/FROM ;
  wire \DLX_EXinst_Mshift__n0023_Sh<29>/GROM ;
  wire \CHOICE5943/FROM ;
  wire \CHOICE5943/GROM ;
  wire \DLX_IDinst_Imm<15>/FROM ;
  wire DLX_IDinst__n0090;
  wire \CHOICE1962/FROM ;
  wire \CHOICE1962/GROM ;
  wire \CHOICE5724/FROM ;
  wire \CHOICE5724/GROM ;
  wire \CHOICE1036/FROM ;
  wire \CHOICE1036/GROM ;
  wire \CHOICE4693/FROM ;
  wire \CHOICE4693/GROM ;
  wire \CHOICE4763/FROM ;
  wire \CHOICE4763/GROM ;
  wire \CHOICE1144/FROM ;
  wire \CHOICE1144/GROM ;
  wire \DLX_EXinst_Mshift__n0026_Sh<50>/FROM ;
  wire \DLX_EXinst_Mshift__n0026_Sh<50>/GROM ;
  wire \CHOICE5730/FROM ;
  wire \CHOICE5730/GROM ;
  wire \N127346/FROM ;
  wire \N127346/GROM ;
  wire \CHOICE1911/FROM ;
  wire \CHOICE1911/GROM ;
  wire \CHOICE1972/FROM ;
  wire \CHOICE1972/GROM ;
  wire \DLX_EXinst_Mshift__n0023_Sh<26>/FROM ;
  wire \DLX_EXinst_Mshift__n0023_Sh<26>/GROM ;
  wire \CHOICE5714/FROM ;
  wire \CHOICE5714/GROM ;
  wire \CHOICE1276/FROM ;
  wire \CHOICE1276/GROM ;
  wire \CHOICE4520/FROM ;
  wire \CHOICE4520/GROM ;
  wire \DLX_EXlc_md_wint28/FROM ;
  wire \DLX_EXlc_md_wint28/GROM ;
  wire \CHOICE3032/FROM ;
  wire \CHOICE3032/GROM ;
  wire \N98808/FROM ;
  wire \N98808/GROM ;
  wire \DLX_EXinst_ALU_result<0>/FROM ;
  wire \DLX_EXinst_ALU_result<0>/GROM ;
  wire \N125971/FROM ;
  wire \N125971/GROM ;
  wire \CHOICE5982/FROM ;
  wire \CHOICE5982/GROM ;
  wire \DLX_EXinst_ALU_result<1>/FROM ;
  wire \DLX_EXinst_ALU_result<1>/GROM ;
  wire \CHOICE4453/FROM ;
  wire \CHOICE4453/GROM ;
  wire \CHOICE4698/FROM ;
  wire \CHOICE4698/GROM ;
  wire \vga_top_vga1_videoon/LOGIC_ONE ;
  wire \CHOICE1379/FROM ;
  wire \CHOICE1379/GROM ;
  wire \CHOICE1150/FROM ;
  wire \CHOICE1150/GROM ;
  wire \CHOICE2069/FROM ;
  wire \CHOICE2069/GROM ;
  wire \DLX_EXlc_md_wint25/FROM ;
  wire \DLX_EXlc_md_wint25/GROM ;
  wire \CHOICE5542/FROM ;
  wire \CHOICE5542/GROM ;
  wire \CHOICE4130/FROM ;
  wire \CHOICE4130/GROM ;
  wire \CHOICE4385/FROM ;
  wire \CHOICE4385/GROM ;
  wire \CHOICE5520/FROM ;
  wire \CHOICE5520/GROM ;
  wire \CHOICE5988/FROM ;
  wire \CHOICE5988/GROM ;
  wire \CHOICE2980/FROM ;
  wire \CHOICE2980/GROM ;
  wire \CHOICE5558/FROM ;
  wire \CHOICE5558/GROM ;
  wire \N94205/FROM ;
  wire \N94205/GROM ;
  wire \DLX_EXinst_Mshift__n0026_Sh<30>/FROM ;
  wire \DLX_EXinst_Mshift__n0026_Sh<30>/GROM ;
  wire \CHOICE3069/FROM ;
  wire \CHOICE3069/GROM ;
  wire \DLX_EXlc_md_wint24/FROM ;
  wire \DLX_EXlc_md_wint24/GROM ;
  wire \DLX_EXinst_Mshift__n0026_Sh<6>/FROM ;
  wire \DLX_EXinst_Mshift__n0026_Sh<6>/GROM ;
  wire \CHOICE4537/FROM ;
  wire \CHOICE4537/GROM ;
  wire \CHOICE5548/FROM ;
  wire \CHOICE5548/GROM ;
  wire \CHOICE5300/FROM ;
  wire \CHOICE5300/GROM ;
  wire \CHOICE1349/FROM ;
  wire \CHOICE1349/GROM ;
  wire \CHOICE1102/FROM ;
  wire \CHOICE1102/GROM ;
  wire \DLX_EXinst_Mshift__n0026_Sh<21>/FROM ;
  wire \DLX_EXinst_Mshift__n0026_Sh<21>/GROM ;
  wire \DLX_EXlc_md_wint23/FROM ;
  wire \DLX_EXlc_md_wint23/GROM ;
  wire \CHOICE5201/FROM ;
  wire \CHOICE5201/GROM ;
  wire \CHOICE5049/FROM ;
  wire \CHOICE5049/GROM ;
  wire \N126006/FROM ;
  wire \N126006/GROM ;
  wire \CHOICE5086/FROM ;
  wire \CHOICE5086/GROM ;
  wire \DLX_EXinst_Mshift__n0026_Sh<22>/FROM ;
  wire \DLX_EXinst_Mshift__n0026_Sh<22>/GROM ;
  wire \N100191/FROM ;
  wire \N100191/GROM ;
  wire \CHOICE1337/FROM ;
  wire \CHOICE1337/GROM ;
  wire \N107444/FROM ;
  wire \N107444/GROM ;
  wire \DLX_EXinst_N66072/FROM ;
  wire \DLX_EXinst_N66072/GROM ;
  wire \N127350/FROM ;
  wire \N127350/GROM ;
  wire \DLX_EXlc_md_wint22/FROM ;
  wire \DLX_EXlc_md_wint22/GROM ;
  wire \CHOICE5353/FROM ;
  wire \CHOICE5353/GROM ;
  wire \DLX_EXinst_ALU_result<3>/FROM ;
  wire \DLX_EXinst_ALU_result<3>/GROM ;
  wire \CHOICE3214/FROM ;
  wire \CHOICE3214/GROM ;
  wire \CHOICE5056/FROM ;
  wire \CHOICE5056/GROM ;
  wire \N109350/FROM ;
  wire \N109350/GROM ;
  wire \DLX_EXinst_Mshift__n0026_Sh<16>/FROM ;
  wire \DLX_EXinst_Mshift__n0026_Sh<16>/GROM ;
  wire \CHOICE4003/FROM ;
  wire \CHOICE4003/GROM ;
  wire \DLX_EXinst_Mshift__n0028_Sh<57>/FROM ;
  wire \DLX_EXinst_Mshift__n0028_Sh<57>/GROM ;
  wire \CHOICE1180/FROM ;
  wire \CHOICE1180/GROM ;
  wire \DLX_IDinst_reg_out_B<0>/FROM ;
  wire \N94921/FROM ;
  wire \N94921/GROM ;
  wire \CHOICE4464/FROM ;
  wire \CHOICE4464/GROM ;
  wire \CHOICE3844/FROM ;
  wire \CHOICE3844/GROM ;
  wire \CHOICE5613/FROM ;
  wire \CHOICE5613/GROM ;
  wire \CHOICE1288/FROM ;
  wire \CHOICE1288/GROM ;
  wire \CHOICE3564/FROM ;
  wire \CHOICE3564/GROM ;
  wire \CHOICE1048/FROM ;
  wire \CHOICE1048/GROM ;
  wire \DLX_EXinst_ALU_result<4>/FROM ;
  wire \DLX_EXinst_ALU_result<4>/GROM ;
  wire \CHOICE4017/FROM ;
  wire \CHOICE4017/GROM ;
  wire \CHOICE5236/FROM ;
  wire \CHOICE5236/GROM ;
  wire \DLX_IDinst_WB_data_eff<30>/FROM ;
  wire \DLX_IDinst_WB_data_eff<30>/GROM ;
  wire \CHOICE3415/FROM ;
  wire \CHOICE3415/GROM ;
  wire \N94107/FROM ;
  wire \N94107/GROM ;
  wire \DLX_IDinst_WB_data_eff<28>/FROM ;
  wire \DLX_IDinst_WB_data_eff<28>/GROM ;
  wire \CHOICE4064/FROM ;
  wire \CHOICE4064/GROM ;
  wire \N97892/FROM ;
  wire \N97892/GROM ;
  wire \CHOICE4446/FROM ;
  wire \CHOICE4446/GROM ;
  wire \DLX_IDinst_WB_data_eff<27>/FROM ;
  wire \DLX_IDinst_WB_data_eff<27>/GROM ;
  wire \CHOICE3547/FROM ;
  wire \CHOICE3547/GROM ;
  wire \DLX_IDinst_WB_data_eff<26>/FROM ;
  wire \DLX_IDinst_WB_data_eff<26>/GROM ;
  wire \CHOICE4475/FROM ;
  wire \CHOICE4475/GROM ;
  wire \DLX_EXinst_ALU_result<5>/FROM ;
  wire \DLX_EXinst_ALU_result<5>/GROM ;
  wire \DLX_IDinst_WB_data_eff<25>/FROM ;
  wire \DLX_IDinst_WB_data_eff<25>/GROM ;
  wire \DLX_IDinst_WB_data_eff<19>/FROM ;
  wire \DLX_IDinst_WB_data_eff<19>/GROM ;
  wire \CHOICE3551/FROM ;
  wire \CHOICE3551/GROM ;
  wire \CHOICE3024/FROM ;
  wire \CHOICE3024/GROM ;
  wire \N127338/FROM ;
  wire \N127338/GROM ;
  wire \N127342/FROM ;
  wire \N127342/GROM ;
  wire \DLX_IDinst_N69781/FROM ;
  wire \DLX_IDinst_N69781/GROM ;
  wire \CHOICE4596/FROM ;
  wire \CHOICE4596/GROM ;
  wire \CHOICE5801/FROM ;
  wire \CHOICE5801/GROM ;
  wire \CHOICE1096/FROM ;
  wire \CHOICE1096/GROM ;
  wire \DLX_IDinst_WB_data_eff<18>/FROM ;
  wire \DLX_IDinst_WB_data_eff<18>/GROM ;
  wire \N126571/FROM ;
  wire \N126571/GROM ;
  wire \N94857/FROM ;
  wire \N94857/GROM ;
  wire \CHOICE4378/FROM ;
  wire \CHOICE4378/GROM ;
  wire \CHOICE4478/FROM ;
  wire \CHOICE4478/GROM ;
  wire \CHOICE4397/FROM ;
  wire \CHOICE4397/GROM ;
  wire \CHOICE1417/FROM ;
  wire \CHOICE1417/GROM ;
  wire \DLX_EXinst_Mshift__n0026_Sh<49>/FROM ;
  wire \DLX_EXinst_Mshift__n0026_Sh<49>/GROM ;
  wire \CHOICE1216/FROM ;
  wire \CHOICE1216/GROM ;
  wire \CHOICE3377/FROM ;
  wire \CHOICE3377/GROM ;
  wire \DLX_EXinst_ALU_result<22>/FROM ;
  wire N114452;
  wire \DLX_EXinst_ALU_result<6>/FROM ;
  wire \DLX_EXinst_ALU_result<6>/GROM ;
  wire \CHOICE4407/FROM ;
  wire \CHOICE4407/GROM ;
  wire \CHOICE1108/FROM ;
  wire \CHOICE1108/GROM ;
  wire \CHOICE5383/FROM ;
  wire \CHOICE5383/GROM ;
  wire \DLX_EXlc_md_wint21/FROM ;
  wire \DLX_EXlc_md_wint21/GROM ;
  wire \CHOICE1926/FROM ;
  wire \CHOICE1926/GROM ;
  wire \CHOICE4410/FROM ;
  wire \CHOICE4410/GROM ;
  wire \CHOICE3826/FROM ;
  wire \CHOICE3826/GROM ;
  wire \CHOICE2815/FROM ;
  wire \CHOICE2815/GROM ;
  wire \CHOICE3045/FROM ;
  wire \CHOICE3045/GROM ;
  wire \CHOICE4576/FROM ;
  wire \CHOICE4576/GROM ;
  wire \DLX_IFlc_master_ctrlIF_nro/FROM ;
  wire \DLX_IFlc_master_ctrlIF_nro/GROM ;
  wire \CHOICE3491/FROM ;
  wire \CHOICE3491/GROM ;
  wire \DLX_IDinst_branch_address<11>/FROM ;
  wire N105787;
  wire \DLX_IDinst_mem_to_reg/FROM ;
  wire DLX_IDinst__n0110;
  wire \DLX_EXlc_md_wint36/FROM ;
  wire \DLX_EXlc_md_wint36/GROM ;
  wire \DLX_EXinst_Mshift__n0027_Sh<0>/FROM ;
  wire \DLX_EXinst_Mshift__n0027_Sh<0>/GROM ;
  wire \DLX_EXinst_Mshift__n0027_Sh<41>/FROM ;
  wire \DLX_EXinst_Mshift__n0027_Sh<41>/GROM ;
  wire \CHOICE4588/FROM ;
  wire \CHOICE4588/GROM ;
  wire \DLX_EXinst_ALU_result<18>/FROM ;
  wire N122511;
  wire \DLX_EXinst_ALU_result<26>/FROM ;
  wire N117936;
  wire \CHOICE3295/FROM ;
  wire \CHOICE3295/GROM ;
  wire \CHOICE994/FROM ;
  wire \CHOICE994/GROM ;
  wire \DLX_RF_delay_inst_wint4/GROM ;
  wire \CHOICE2551/FROM ;
  wire \CHOICE2551/GROM ;
  wire \DLX_IDinst_CLI/FROM ;
  wire \DLX_IDinst_CLI/GROM ;
  wire \DLX_IDinst__n0135/FROM ;
  wire \DLX_IDinst__n0135/GROM ;
  wire \DLX_RF_delay_inst_wint5/GROM ;
  wire \CHOICE4602/FROM ;
  wire \CHOICE4602/GROM ;
  wire \DLX_IDinst__n0145/FROM ;
  wire \DLX_IDinst__n0145/GROM ;
  wire \DLX_IDinst__n0144/FROM ;
  wire \DLX_IDinst__n0144/GROM ;
  wire \DLX_IDinst_branch_address<12>/FROM ;
  wire N105850;
  wire \DLX_EXlc_md_wint37/FROM ;
  wire \DLX_EXlc_md_wint37/GROM ;
  wire \DLX_IDinst_branch_address<20>/FROM ;
  wire N106354;
  wire \DLX_EXinst_ALU_result<9>/FROM ;
  wire \DLX_EXinst_ALU_result<9>/GROM ;
  wire \DLX_RF_delay_inst_wint6/GROM ;
  wire \DLX_IDinst_Ker709161_1/FROM ;
  wire \DLX_IDinst_Ker709161_1/GROM ;
  wire \DLX_RF_delay_inst_wint7/GROM ;
  wire \DLX_RF_delay_inst_wint8/GROM ;
  wire \DLX_IDinst__n0147/FROM ;
  wire \DLX_IDinst__n0147/GROM ;
  wire \N90255/FROM ;
  wire \N90255/GROM ;
  wire \DLX_RF_delay_inst_wint9/GROM ;
  wire \DLX_IDinst_branch_address<21>/FROM ;
  wire N106480;
  wire \DLX_IDinst_branch_address<13>/FROM ;
  wire N105913;
  wire \DLX_IDlc_md_wint33/FROM ;
  wire \DLX_IDlc_md_wint33/GROM ;
  wire \CHOICE1168/FROM ;
  wire \CHOICE1168/GROM ;
  wire \CHOICE1436/FROM ;
  wire \CHOICE1436/GROM ;
  wire \DLX_IDinst__n0173/FROM ;
  wire \DLX_IDinst__n0173/GROM ;
  wire \CHOICE2760/FROM ;
  wire \CHOICE2760/GROM ;
  wire \DLX_EXinst_noop/FROM ;
  wire N101911;
  wire \DLX_IDinst__n0350/FROM ;
  wire \DLX_IDinst__n0350/GROM ;
  wire \DLX_IDinst__n0441/FROM ;
  wire \DLX_IDinst__n0441/GROM ;
  wire \N126388/FROM ;
  wire \N126388/GROM ;
  wire \DLX_IDinst_branch_address<14>/FROM ;
  wire N105976;
  wire \DLX_IDinst_branch_address<22>/FROM ;
  wire N106606;
  wire \DLX_IDinst_branch_address<30>/FROM ;
  wire N106417;
  wire \DLX_IDinst__n0344/FROM ;
  wire \DLX_IDinst__n0344/GROM ;
  wire \DLX_EXlc_md_wint34/FROM ;
  wire \DLX_EXlc_md_wint34/GROM ;
  wire \DLX_EXlc_md_wint26/FROM ;
  wire \DLX_EXlc_md_wint26/GROM ;
  wire \DLX_IDinst_branch_address<31>/FROM ;
  wire N107102;
  wire \CHOICE2182/FROM ;
  wire \CHOICE2182/GROM ;
  wire \CHOICE2727/GROM ;
  wire \DLX_EXinst_Mshift__n0027_Sh<7>/FROM ;
  wire \DLX_EXinst_Mshift__n0027_Sh<7>/GROM ;
  wire \CHOICE3466/FROM ;
  wire \CHOICE3466/GROM ;
  wire \DLX_IFlc_ridp3/GROM ;
  wire \DLX_IDinst_branch_address<23>/FROM ;
  wire N106543;
  wire \DLX_IDinst_branch_address<15>/FROM ;
  wire N106039;
  wire \DLX_IDinst__n0348/FROM ;
  wire \DLX_IDinst__n0348/GROM ;
  wire \DLX_IDinst__n0364/FROM ;
  wire \DLX_IDinst__n0364/GROM ;
  wire \DLX_EXinst_Mshift__n0027_Sh<9>/FROM ;
  wire \DLX_EXinst_Mshift__n0027_Sh<9>/GROM ;
  wire \DLX_IDinst_branch_address<16>/FROM ;
  wire N106102;
  wire \DLX_IDinst_branch_address<24>/FROM ;
  wire N106669;
  wire \CHOICE1786/FROM ;
  wire \CHOICE1786/GROM ;
  wire \DLX_EXlc_pd_wint2/GROM ;
  wire \DLX_EXinst__n0030_1/FROM ;
  wire \DLX_EXinst__n0030_1/GROM ;
  wire \N127555/FROM ;
  wire \N127555/GROM ;
  wire \DLX_EXlc_pd_wint3/GROM ;
  wire \DLX_EXlc_pd_wint4/GROM ;
  wire \DLX_IDinst_stall/FROM ;
  wire \DLX_IDinst_stall/GROM ;
  wire \DLX_EXlc_pd_wint5/FROM ;
  wire \DLX_EXlc_pd_wint5/GROM ;
  wire \DLX_IDinst_branch_address<17>/FROM ;
  wire N106165;
  wire \DLX_IDinst_branch_address<25>/FROM ;
  wire N106789;
  wire \DLX_EXinst_N62715/FROM ;
  wire \DLX_EXinst_N62715/GROM ;
  wire \DLX_IFinst_NPC<10>/FROM ;
  wire \DLX_IFinst_NPC<10>/GROM ;
  wire \DLX_IDinst_branch_address<26>/FROM ;
  wire N106852;
  wire \DLX_IDinst_branch_address<18>/FROM ;
  wire N106291;
  wire \CHOICE5/FROM ;
  wire \CHOICE5/GROM ;
  wire \DLX_EXlc_md_wint38/GROM ;
  wire \DLX_EXinst_N62727/FROM ;
  wire \DLX_EXinst_N62727/GROM ;
  wire \DLX_EXinst_N64181/FROM ;
  wire \DLX_EXinst_N64181/GROM ;
  wire \DLX_IDinst_branch_address<27>/FROM ;
  wire N106915;
  wire \DLX_IDinst_branch_address<19>/FROM ;
  wire N106228;
  wire \DLX_EXlc_md_wint39/GROM ;
  wire \DLX_EXinst_N64448/FROM ;
  wire \DLX_EXinst_N64448/GROM ;
  wire \N126428/FROM ;
  wire \N126428/GROM ;
  wire \CHOICE1790/FROM ;
  wire \CHOICE1790/GROM ;
  wire \DLX_IDinst_branch_address<28>/FROM ;
  wire N106978;
  wire \N126169/FROM ;
  wire \N126169/GROM ;
  wire \DLX_EXinst_ALU_result<14>/FROM ;
  wire \DLX_EXinst_ALU_result<14>/GROM ;
  wire \DLX_EXinst__n0030/FROM ;
  wire \DLX_EXinst__n0030/GROM ;
  wire \DLX_IDinst_branch_address<29>/FROM ;
  wire N107041;
  wire \DLX_EXinst_N66519/FROM ;
  wire \DLX_EXinst_N66519/GROM ;
  wire \DLX_EXinst_N64919/FROM ;
  wire \DLX_EXinst_N64919/GROM ;
  wire \N126490/FROM ;
  wire \N126490/GROM ;
  wire \DLX_IFinst_NPC<11>/FROM ;
  wire \DLX_IFinst_NPC<11>/GROM ;
  wire \DLX_EXinst__n0128/FROM ;
  wire \DLX_EXinst__n0128/GROM ;
  wire \DLX_IDlc_md_wint32/FROM ;
  wire \DLX_IDlc_md_wint32/GROM ;
  wire \DLX_IDlc_md_wint29/FROM ;
  wire \DLX_IDlc_md_wint29/GROM ;
  wire \CHOICE4217/FROM ;
  wire \CHOICE4217/GROM ;
  wire \DLX_IFinst_NPC<20>/FROM ;
  wire \DLX_IFinst_NPC<12>/FROM ;
  wire \DLX_IFinst_NPC<12>/GROM ;
  wire \DLX_IDlc_md_wint28/FROM ;
  wire \DLX_IDlc_md_wint28/GROM ;
  wire \DLX_IDlc_md_wint25/FROM ;
  wire \DLX_IDlc_md_wint25/GROM ;
  wire \clk_DM_OBUF/GROM ;
  wire \DLX_IFinst_NPC<0>/FROM ;
  wire \DLX_IFinst_NPC<0>/GROM ;
  wire \DLX_IDlc_md_wint24/FROM ;
  wire \DLX_IDlc_md_wint24/GROM ;
  wire \DLX_IDlc_md_wint23/FROM ;
  wire \DLX_IDlc_md_wint23/GROM ;
  wire \N126048/FROM ;
  wire \N126048/GROM ;
  wire \CHOICE2646/GROM ;
  wire \DLX_IDinst_regA_eff<10>/FROM ;
  wire \DLX_IDinst_regA_eff<10>/GROM ;
  wire \DLX_IDlc_md_wint30/FROM ;
  wire \DLX_IDlc_md_wint30/GROM ;
  wire \DLX_IDlc_md_wint19/FROM ;
  wire \DLX_IDlc_md_wint19/GROM ;
  wire \DLX_IDlc_md_wint18/FROM ;
  wire \DLX_IDlc_md_wint18/GROM ;
  wire \CHOICE32/FROM ;
  wire \CHOICE32/GROM ;
  wire \CHOICE3328/FROM ;
  wire \CHOICE3328/GROM ;
  wire \DLX_IDinst_regA_eff<11>/FROM ;
  wire \DLX_IDinst_regA_eff<11>/GROM ;
  wire \N95327/FROM ;
  wire \N95327/GROM ;
  wire \DLX_IDinst_regA_eff<12>/FROM ;
  wire \DLX_IDinst_regA_eff<12>/GROM ;
  wire \DLX_IDinst_regA_eff<20>/FROM ;
  wire \DLX_IDinst_regA_eff<20>/GROM ;
  wire \DLX_IDlc_md_wint17/FROM ;
  wire \DLX_IDlc_md_wint17/GROM ;
  wire \DLX_EXinst_Mshift__n0027_Sh<10>/FROM ;
  wire \DLX_EXinst_Mshift__n0027_Sh<10>/GROM ;
  wire \DLX_EXinst_Mshift__n0023_Sh<30>/FROM ;
  wire \DLX_EXinst_Mshift__n0023_Sh<30>/GROM ;
  wire \DLX_MEMinst_noop/CKMUXNOT ;
  wire \DLX_IDinst_regA_eff<13>/FROM ;
  wire \DLX_IDinst_regA_eff<13>/GROM ;
  wire \DLX_IDinst_regA_eff<21>/FROM ;
  wire \DLX_IDinst_regA_eff<21>/GROM ;
  wire \DLX_IFinst_NPC<13>/FROM ;
  wire \DLX_IFinst_NPC<13>/GROM ;
  wire \DLX_IFinst_NPC<21>/FROM ;
  wire \DLX_IDinst_regA_eff<14>/FROM ;
  wire \DLX_IDinst_regA_eff<14>/GROM ;
  wire \DLX_IDinst_regA_eff<22>/FROM ;
  wire \DLX_IDinst_regA_eff<22>/GROM ;
  wire \CHOICE3343/FROM ;
  wire \CHOICE3343/GROM ;
  wire \DLX_IDlc_md_wint9/FROM ;
  wire \DLX_IDlc_md_wint9/GROM ;
  wire \DLX_EXinst_Mshift__n0027_Sh<12>/FROM ;
  wire \DLX_EXinst_Mshift__n0027_Sh<12>/GROM ;
  wire \DLX_IDinst_regA_eff<15>/FROM ;
  wire \DLX_IDinst_regA_eff<15>/GROM ;
  wire \DLX_IDinst_regA_eff<23>/FROM ;
  wire \DLX_IDinst_regA_eff<23>/GROM ;
  wire \DLX_IDinst_regA_eff<31>/FROM ;
  wire \DLX_IDinst_regA_eff<31>/GROM ;
  wire \DLX_EXinst_Mshift__n0027_Sh<13>/FROM ;
  wire \DLX_EXinst_Mshift__n0027_Sh<13>/GROM ;
  wire \DLX_IFinst_NPC<1>/FROM ;
  wire \DLX_IFinst_NPC<1>/GROM ;
  wire \DLX_IDinst_regA_eff<16>/FROM ;
  wire \DLX_IDinst_regA_eff<16>/GROM ;
  wire \DLX_IDinst_regA_eff<24>/FROM ;
  wire \DLX_IDinst_regA_eff<24>/GROM ;
  wire \DLX_EXinst_Mshift__n0027_Sh<14>/FROM ;
  wire \DLX_EXinst_Mshift__n0027_Sh<14>/GROM ;
  wire \CHOICE4514/FROM ;
  wire \CHOICE4514/GROM ;
  wire \DLX_IDinst_regA_eff<17>/FROM ;
  wire \DLX_IDinst_regA_eff<17>/GROM ;
  wire \DLX_IDinst_regA_eff<25>/FROM ;
  wire \DLX_IDinst_regA_eff<25>/GROM ;
  wire \DLX_IDinst_regA_eff<18>/FROM ;
  wire \DLX_IDinst_regA_eff<18>/GROM ;
  wire \DLX_IDinst_regA_eff<26>/FROM ;
  wire \DLX_IDinst_regA_eff<26>/GROM ;
  wire \DLX_IDlc_md_wint34/FROM ;
  wire \DLX_IDlc_md_wint34/GROM ;
  wire \DLX_IDlc_md_wint26/FROM ;
  wire \DLX_IDlc_md_wint26/GROM ;
  wire \CHOICE4540/FROM ;
  wire \CHOICE4540/GROM ;
  wire \DLX_IDinst_regA_eff<19>/FROM ;
  wire \DLX_IDinst_regA_eff<19>/GROM ;
  wire \DLX_IDinst_regA_eff<27>/FROM ;
  wire \DLX_IDinst_regA_eff<27>/GROM ;
  wire \DLX_EXinst_Mshift__n0023_Sh<61>/FROM ;
  wire \DLX_EXinst_Mshift__n0023_Sh<61>/GROM ;
  wire \CHOICE4532/FROM ;
  wire \CHOICE4532/GROM ;
  wire \DLX_IDinst_regA_eff<28>/FROM ;
  wire \DLX_IDinst_regA_eff<28>/GROM ;
  wire \N126564/FROM ;
  wire \N126564/GROM ;
  wire \DLX_EXinst_ALU_result<10>/FROM ;
  wire \DLX_EXinst_ALU_result<10>/GROM ;
  wire \CHOICE3944/FROM ;
  wire \CHOICE3944/GROM ;
  wire \DLX_IDinst_regA_eff<29>/FROM ;
  wire \DLX_IDinst_regA_eff<29>/GROM ;
  wire \DLX_IFinst_NPC<30>/FROM ;
  wire \DLX_IFinst_NPC<14>/FROM ;
  wire \DLX_IFinst_NPC<14>/GROM ;
  wire \DLX_IFinst_NPC<22>/FROM ;
  wire \CHOICE3966/FROM ;
  wire \CHOICE3966/GROM ;
  wire \DLX_IDinst_reg_dst/FROM ;
  wire N110380;
  wire \DLX_EXinst__n0093/FROM ;
  wire \DLX_EXinst__n0093/GROM ;
  wire \CHOICE4643/FROM ;
  wire \CHOICE4643/GROM ;
  wire \DLX_IDlc_md_wint8/FROM ;
  wire \DLX_IDlc_md_wint8/GROM ;
  wire \CHOICE5451/FROM ;
  wire \CHOICE5451/GROM ;
  wire \DLX_EXinst_ALU_result<11>/FROM ;
  wire \DLX_EXinst_ALU_result<11>/GROM ;
  wire \DLX_IFinst_NPC<2>/FROM ;
  wire \DLX_IFinst_NPC<2>/GROM ;
  wire \CHOICE3963/FROM ;
  wire \CHOICE3963/GROM ;
  wire \DLX_IDlc_md_wint7/FROM ;
  wire \DLX_IDlc_md_wint7/GROM ;
  wire \CHOICE5321/FROM ;
  wire \CHOICE5321/GROM ;
  wire \DLX_EXinst_ALU_result<20>/FROM ;
  wire N119151;
  wire \CHOICE1000/FROM ;
  wire \CHOICE1000/GROM ;
  wire \CHOICE5447/FROM ;
  wire \CHOICE5447/GROM ;
  wire \CHOICE2521/FROM ;
  wire \CHOICE2521/GROM ;
  wire \CHOICE4928/FROM ;
  wire \CHOICE4928/GROM ;
  wire \CHOICE3908/FROM ;
  wire \CHOICE3908/GROM ;
  wire \CHOICE1120/FROM ;
  wire \CHOICE1120/GROM ;
  wire \CHOICE4925/FROM ;
  wire \CHOICE4925/GROM ;
  wire \DLX_IDlc_md_wint6/FROM ;
  wire \DLX_IDlc_md_wint6/GROM ;
  wire \CHOICE4145/FROM ;
  wire \CHOICE4145/GROM ;
  wire \CHOICE4057/FROM ;
  wire \CHOICE4057/GROM ;
  wire \CHOICE3895/FROM ;
  wire \CHOICE3895/GROM ;
  wire \vga_select_6<0>/FROM ;
  wire \vga_select_6<0>/GROM ;
  wire \CHOICE4256/FROM ;
  wire \CHOICE4256/GROM ;
  wire \CHOICE3903/FROM ;
  wire \CHOICE3903/GROM ;
  wire \CHOICE4913/FROM ;
  wire \CHOICE4913/GROM ;
  wire \vga_select_6<5>/FROM ;
  wire \vga_select_6<5>/GROM ;
  wire \DLX_EXinst_Mshift__n0027_Sh<4>/FROM ;
  wire \DLX_EXinst_Mshift__n0027_Sh<4>/GROM ;
  wire \DLX_IDlc_md_wint5/FROM ;
  wire \DLX_IDlc_md_wint5/GROM ;
  wire \DLX_EXinst_ALU_result<23>/FROM ;
  wire N114054;
  wire \CHOICE4999/FROM ;
  wire \CHOICE4999/GROM ;
  wire \DLX_IFinst_NPC<15>/FROM ;
  wire \DLX_IFinst_NPC<15>/GROM ;
  wire \DLX_IFinst_NPC<31>/FROM ;
  wire \DLX_IFinst_NPC<23>/FROM ;
  wire \CHOICE4219/FROM ;
  wire \CHOICE4219/GROM ;
  wire \CHOICE1024/FROM ;
  wire \CHOICE1024/GROM ;
  wire \CHOICE4708/FROM ;
  wire \CHOICE4708/GROM ;
  wire \DLX_EXlc_master_ctrlEX_nro/FROM ;
  wire \DLX_EXlc_master_ctrlEX_nro/GROM ;
  wire \CHOICE4342/FROM ;
  wire \CHOICE4342/GROM ;
  wire \CHOICE4205/FROM ;
  wire \CHOICE4205/GROM ;
  wire \CHOICE4337/FROM ;
  wire \CHOICE4337/GROM ;
  wire \CHOICE4327/FROM ;
  wire \CHOICE4327/GROM ;
  wire \vga_select_6<4>/FROM ;
  wire \vga_select_6<4>/GROM ;
  wire \DLX_IFinst_NPC<3>/FROM ;
  wire \DLX_IFinst_NPC<3>/GROM ;
  wire \CHOICE4154/FROM ;
  wire \CHOICE4154/GROM ;
  wire \CHOICE4151/FROM ;
  wire \CHOICE4151/GROM ;
  wire \DLX_IDinst_slot_num_FFd3/FROM ;
  wire \DLX_IDinst_slot_num_FFd3-In ;
  wire \N127567/FROM ;
  wire \N127567/GROM ;
  wire \CHOICE4282/FROM ;
  wire \CHOICE4282/GROM ;
  wire \CHOICE4139/FROM ;
  wire \CHOICE4139/GROM ;
  wire \CHOICE4277/FROM ;
  wire \CHOICE4277/GROM ;
  wire \CHOICE4267/FROM ;
  wire \CHOICE4267/GROM ;
  wire \CHOICE5247/FROM ;
  wire \CHOICE5247/GROM ;
  wire \CHOICE4831/GROM ;
  wire \CHOICE5784/FROM ;
  wire \CHOICE5784/GROM ;
  wire \CHOICE5315/FROM ;
  wire \CHOICE5315/GROM ;
  wire \CHOICE4860/FROM ;
  wire \CHOICE4860/GROM ;
  wire \CHOICE5169/FROM ;
  wire \CHOICE5169/GROM ;
  wire \CHOICE4085/FROM ;
  wire \CHOICE4085/GROM ;
  wire \DLX_IFinst_NPC<24>/FROM ;
  wire \DLX_IFinst_NPC<16>/FROM ;
  wire \DLX_EXinst_ALU_result<30>/FROM ;
  wire N121549;
  wire \N127563/FROM ;
  wire \N127563/GROM ;
  wire \CHOICE3766/FROM ;
  wire \CHOICE3766/GROM ;
  wire \CHOICE4865/FROM ;
  wire \CHOICE4865/GROM ;
  wire \CHOICE4073/FROM ;
  wire \CHOICE4073/GROM ;
  wire \CHOICE5440/FROM ;
  wire \CHOICE5440/GROM ;
  wire \CHOICE5785/FROM ;
  wire \CHOICE5785/GROM ;
  wire \DLX_IFinst_NPC<4>/FROM ;
  wire \DLX_IFinst_NPC<4>/GROM ;
  wire \DLX_EXinst_ALU_result<27>/FROM ;
  wire N117545;
  wire \DLX_EXinst_ALU_result<15>/FROM ;
  wire N118737;
  wire \DLX_MEMinst_reg_dst_out<1>/CKMUXNOT ;
  wire \CHOICE5818/FROM ;
  wire \CHOICE5818/GROM ;
  wire \DLX_EXinst_ALU_result<31>/FROM ;
  wire N124731;
  wire \CHOICE5128/GROM ;
  wire \DLX_MEMinst_reg_dst_out<3>/CKMUXNOT ;
  wire \CHOICE3789/FROM ;
  wire \CHOICE3789/GROM ;
  wire \CHOICE5145/FROM ;
  wire \CHOICE5145/GROM ;
  wire \DLX_MEMinst_reg_dst_out<4>/CKMUXNOT ;
  wire \DLX_reqout_MEM/FROM ;
  wire \DLX_reqout_MEM/GROM ;
  wire \DLX_MEMlc_md_wint10/FROM ;
  wire \DLX_MEMlc_md_wint10/GROM ;
  wire \CHOICE5824/FROM ;
  wire \CHOICE5824/GROM ;
  wire \CHOICE5168/GROM ;
  wire \N126344/FROM ;
  wire \N126344/GROM ;
  wire \CHOICE3773/FROM ;
  wire \CHOICE3773/GROM ;
  wire \CHOICE5603/FROM ;
  wire \CHOICE5603/GROM ;
  wire \N127423/GROM ;
  wire \DLX_IFinst_NPC<17>/FROM ;
  wire \N90373/FROM ;
  wire \N90373/GROM ;
  wire \CHOICE5642/FROM ;
  wire \CHOICE5642/GROM ;
  wire \DLX_IFinst_NPC<25>/FROM ;
  wire \CHOICE3783/FROM ;
  wire \CHOICE3783/GROM ;
  wire \DLX_EXinst_ALU_result<16>/FROM ;
  wire N120627;
  wire \CHOICE4790/FROM ;
  wire \CHOICE4790/GROM ;
  wire \vga_select_6<1>/GROM ;
  wire \CHOICE5625/FROM ;
  wire \CHOICE5625/GROM ;
  wire \CHOICE4701/FROM ;
  wire \CHOICE4701/GROM ;
  wire \vga_select_6<2>/FROM ;
  wire \vga_select_6<2>/GROM ;
  wire \CHOICE4773/GROM ;
  wire \CHOICE5646/FROM ;
  wire \CHOICE5646/GROM ;
  wire \DLX_IFinst_NPC<5>/FROM ;
  wire \DLX_IFinst_NPC<5>/GROM ;
  wire \CHOICE4782/FROM ;
  wire \CHOICE4782/GROM ;
  wire \vga_select_6<3>/FROM ;
  wire \vga_select_6<3>/GROM ;
  wire \CHOICE2937/FROM ;
  wire \CHOICE2937/GROM ;
  wire \CHOICE5437/FROM ;
  wire \CHOICE5437/GROM ;
  wire \CHOICE5476/FROM ;
  wire \CHOICE5476/GROM ;
  wire \CHOICE4725/FROM ;
  wire \CHOICE4725/GROM ;
  wire \CHOICE4731/FROM ;
  wire \CHOICE4731/GROM ;
  wire \DLX_MEMlc_md_wint14/FROM ;
  wire \DLX_MEMlc_md_wint14/GROM ;
  wire \CHOICE5459/FROM ;
  wire \CHOICE5459/GROM ;
  wire \CHOICE4715/FROM ;
  wire \CHOICE4715/GROM ;
  wire \DLX_reqout_ID/FROM ;
  wire \DLX_reqout_ID/GROM ;
  wire \red_1_OBUF/FROM ;
  wire \red_1_OBUF/GROM ;
  wire \CHOICE5480/FROM ;
  wire \CHOICE5480/GROM ;
  wire \N107291/FROM ;
  wire \N107291/GROM ;
  wire \DLX_EXinst_Mshift__n0025_Sh<7>/FROM ;
  wire \DLX_EXinst_Mshift__n0025_Sh<7>/GROM ;
  wire \N126542/FROM ;
  wire \N126542/GROM ;
  wire \DLX_EXinst__n0095/FROM ;
  wire \DLX_EXinst__n0095/GROM ;
  wire \DLX_IFinst_NPC<26>/FROM ;
  wire \N126432/FROM ;
  wire \N126432/GROM ;
  wire \DLX_IFinst_NPC<18>/FROM ;
  wire \CHOICE4660/FROM ;
  wire \CHOICE4660/GROM ;
  wire \CHOICE4666/FROM ;
  wire \CHOICE4666/GROM ;
  wire \DLX_MEMlc_md_wint18/FROM ;
  wire \DLX_MEMlc_md_wint18/GROM ;
  wire \CHOICE4650/FROM ;
  wire \CHOICE4650/GROM ;
  wire \CHOICE5008/GROM ;
  wire \N108101/FROM ;
  wire \N108101/GROM ;
  wire \DLX_MEMlc_md_wint19/FROM ;
  wire \DLX_MEMlc_md_wint19/GROM ;
  wire \DLX_IFinst_NPC<6>/FROM ;
  wire \DLX_IFinst_NPC<6>/GROM ;
  wire \DLX_IDinst_reg_write/FROM ;
  wire N110803;
  wire \DLX_IDlc_pd_wint1/FROM ;
  wire \DLX_IDlc_pd_wint1/GROM ;
  wire \DLX_IDinst_counter<0>/FROM ;
  wire N107173;
  wire \DLX_EXinst_Mshift__n0024_Sh<127>/FROM ;
  wire \DLX_EXinst_Mshift__n0024_Sh<127>/GROM ;
  wire \CHOICE5384/FROM ;
  wire \CHOICE5384/GROM ;
  wire \CHOICE5238/FROM ;
  wire \CHOICE5238/GROM ;
  wire \DLX_EXinst_ALU_result<28>/FROM ;
  wire N121082;
  wire \N126551/FROM ;
  wire \N126551/GROM ;
  wire \DLX_IFinst_NPC<19>/FROM ;
  wire \DLX_IFinst_NPC<27>/FROM ;
  wire \N108266/FROM ;
  wire \N108266/GROM ;
  wire \DLX_IDinst_N69568/FROM ;
  wire \DLX_IDinst_N69568/GROM ;
  wire \CHOICE1114/FROM ;
  wire \CHOICE1114/GROM ;
  wire \CHOICE5398/GROM ;
  wire \CHOICE2100/FROM ;
  wire \CHOICE2100/GROM ;
  wire \DLX_IFinst_NPC<7>/FROM ;
  wire \DLX_IFinst_NPC<7>/GROM ;
  wire \N94733/FROM ;
  wire \N94733/GROM ;
  wire \CHOICE5392/FROM ;
  wire \CHOICE5392/GROM ;
  wire \DLX_IDlc_master_ctrlID_nro/GROM ;
  wire \DLX_EXinst_ALU_result<29>/FROM ;
  wire N122016;
  wire \N126207/FROM ;
  wire \N126207/GROM ;
  wire \N126379/FROM ;
  wire \N126379/GROM ;
  wire \DLX_IFinst_NPC<28>/FROM ;
  wire \CHOICE1880/FROM ;
  wire \CHOICE1880/GROM ;
  wire \DM_read_data<25>/FROM ;
  wire \DM_read_data<25>/GROM ;
  wire \DLX_IFinst_NPC<8>/FROM ;
  wire \DLX_IFinst_NPC<8>/GROM ;
  wire \N94673/FROM ;
  wire \N94673/GROM ;
  wire \DM_read_data<26>/FROM ;
  wire \DM_read_data<26>/GROM ;
  wire \DLX_EXinst_Mshift__n0028_Sh<30>/FROM ;
  wire \DLX_EXinst_Mshift__n0028_Sh<30>/GROM ;
  wire \N126620/FROM ;
  wire \N126620/GROM ;
  wire \DM_read_data<27>/FROM ;
  wire \DM_read_data<27>/GROM ;
  wire \DM_read_data<28>/FROM ;
  wire \DM_read_data<28>/GROM ;
  wire \DLX_EXinst_Mshift__n0024_Sh<26>/FROM ;
  wire \DLX_EXinst_Mshift__n0024_Sh<26>/GROM ;
  wire \N126776/GROM ;
  wire \DM_read_data<29>/FROM ;
  wire \DM_read_data<29>/GROM ;
  wire \DM_read_data<31>/FROM ;
  wire \DM_read_data<31>/GROM ;
  wire \red_0_OBUF/GROM ;
  wire \DM_read_data<1>/FROM ;
  wire \DM_read_data<1>/GROM ;
  wire \DM_read_data<2>/FROM ;
  wire \DM_read_data<2>/GROM ;
  wire \N102532/FROM ;
  wire \N102532/GROM ;
  wire \CHOICE2112/GROM ;
  wire \N126473/FROM ;
  wire \N126473/GROM ;
  wire \DM_read_data<3>/FROM ;
  wire \DM_read_data<3>/GROM ;
  wire \DM_read_data<4>/FROM ;
  wire \DM_read_data<4>/GROM ;
  wire \CHOICE3225/FROM ;
  wire \CHOICE3225/GROM ;
  wire \DLX_EXinst_Mshift__n0024_Sh<30>/FROM ;
  wire \DLX_EXinst_Mshift__n0024_Sh<30>/GROM ;
  wire \CHOICE1132/FROM ;
  wire \CHOICE1132/GROM ;
  wire \DLX_IFinst_NPC<29>/FROM ;
  wire \CHOICE3427/GROM ;
  wire \DM_read_data<5>/FROM ;
  wire \DM_read_data<5>/GROM ;
  wire \DM_read_data<6>/FROM ;
  wire \DM_read_data<6>/GROM ;
  wire \N90291/FROM ;
  wire \N90291/GROM ;
  wire \DM_read_data<7>/FROM ;
  wire \DM_read_data<7>/GROM ;
  wire \DLX_MEMinst_reg_write_MEM/CKMUXNOT ;
  wire \CHOICE25/FROM ;
  wire \CHOICE25/GROM ;
  wire \DLX_EXinst_Mshift__n0028_Sh<21>/FROM ;
  wire \DLX_EXinst_Mshift__n0028_Sh<21>/GROM ;
  wire \DM_read_data<8>/FROM ;
  wire \DM_read_data<8>/GROM ;
  wire \DLX_IFinst_NPC<9>/FROM ;
  wire \DLX_IFinst_NPC<9>/GROM ;
  wire \DLX_EXinst_Mshift__n0028_Sh<22>/FROM ;
  wire \DLX_EXinst_Mshift__n0028_Sh<22>/GROM ;
  wire \DM_read_data<9>/FROM ;
  wire \DM_read_data<9>/GROM ;
  wire \N126362/GROM ;
  wire \CHOICE2470/FROM ;
  wire \CHOICE2470/GROM ;
  wire \CHOICE2158/FROM ;
  wire \CHOICE2158/GROM ;
  wire \CHOICE2122/FROM ;
  wire \CHOICE2122/GROM ;
  wire \DLX_EXinst_Mshift__n0028_Sh<49>/FROM ;
  wire \DLX_EXinst_Mshift__n0028_Sh<49>/GROM ;
  wire \CHOICE2362/FROM ;
  wire \CHOICE2362/GROM ;
  wire \DLX_IDinst_reg_out_A<23>/FROM ;
  wire N104236;
  wire \DLX_IDinst_reg_out_A<31>/FROM ;
  wire N102604;
  wire \DLX_IDinst_reg_out_A<15>/FROM ;
  wire N103692;
  wire \DLX_IDinst_reg_out_A<0>/FROM ;
  wire N102740;
  wire \CHOICE2350/FROM ;
  wire \CHOICE2350/GROM ;
  wire \CHOICE2458/FROM ;
  wire \CHOICE2458/GROM ;
  wire \DLX_IDinst_reg_out_A<24>/FROM ;
  wire N104372;
  wire \DLX_IDinst_reg_out_A<16>/FROM ;
  wire N103828;
  wire \CHOICE1459/FROM ;
  wire \CHOICE1459/GROM ;
  wire \DLX_IDinst_reg_out_A<1>/FROM ;
  wire N102672;
  wire \N93641/FROM ;
  wire \N93641/GROM ;
  wire \DLX_IDinst_reg_out_A<17>/FROM ;
  wire N103760;
  wire \DLX_IDinst_reg_out_A<25>/FROM ;
  wire N104304;
  wire \DLX_IDinst_reg_out_A<2>/FROM ;
  wire N102808;
  wire \CHOICE1481/FROM ;
  wire \CHOICE1481/GROM ;
  wire \CHOICE1471/GROM ;
  wire \DLX_IDinst_reg_out_A<26>/FROM ;
  wire N104440;
  wire \DLX_IDinst_reg_out_A<18>/FROM ;
  wire N103896;
  wire \DLX_IDinst_reg_out_A<3>/FROM ;
  wire N102944;
  wire \DLX_IDinst_reg_out_A<27>/FROM ;
  wire N104576;
  wire \DLX_IDinst_reg_out_A<19>/FROM ;
  wire N103964;
  wire \DLX_IDinst_reg_out_A<4>/FROM ;
  wire N102876;
  wire \N90186/FROM ;
  wire \N90186/GROM ;
  wire \DLX_IFinst_IR_latched<10>/FFX/RST ;
  wire \DLX_IFinst_IR_latched<11>/FFX/RST ;
  wire \DLX_IFinst_IR_latched<12>/FFX/RST ;
  wire \DLX_IFinst_IR_latched<20>/FFX/RST ;
  wire \DLX_IFinst_IR_latched<13>/FFX/RST ;
  wire \DLX_IFinst_IR_latched<21>/FFX/RST ;
  wire \DLX_IFinst_IR_latched<14>/FFX/RST ;
  wire \DLX_MEMinst_RF_data_in<11>/FFX/RST ;
  wire \DLX_MEMinst_RF_data_in<21>/FFX/RST ;
  wire \DLX_MEMinst_RF_data_in<13>/FFX/RST ;
  wire \DLX_MEMinst_RF_data_in<31>/FFX/RST ;
  wire \DLX_MEMinst_RF_data_in<23>/FFX/RST ;
  wire \DLX_EXinst_reg_dst_out<4>/FFY/RST ;
  wire \DLX_IDinst_reg_out_B<11>/FFX/RST ;
  wire \DLX_IDinst_reg_out_B<21>/FFX/RST ;
  wire \DLX_IDinst_reg_out_B<13>/FFY/RST ;
  wire \DLX_IDinst_reg_out_B<13>/FFX/RST ;
  wire \DLX_IDinst_reg_out_B<31>/FFY/RST ;
  wire \DLX_IDinst_reg_out_B<31>/FFX/RST ;
  wire \DLX_IDinst_reg_out_B<23>/FFY/RST ;
  wire \DLX_IDinst_reg_out_B<23>/FFX/RST ;
  wire \DLX_IDinst_reg_out_B<15>/FFY/RST ;
  wire \DLX_IFinst_IR_latched<0>/FFX/RST ;
  wire \DLX_IFinst_IR_latched<1>/FFX/RST ;
  wire \DLX_IFinst_IR_latched<2>/FFX/RST ;
  wire \DLX_IFinst_IR_latched<3>/FFX/RST ;
  wire \DLX_IFinst_IR_latched<4>/FFX/RST ;
  wire \DLX_IFinst_IR_latched<5>/FFX/RST ;
  wire \DLX_IFinst_IR_latched<6>/FFX/RST ;
  wire \DLX_IFinst_IR_latched<30>/FFX/RST ;
  wire \DLX_IFinst_IR_latched<22>/FFX/RST ;
  wire \DLX_IFinst_IR_latched<23>/FFX/RST ;
  wire \DLX_IFinst_IR_latched<31>/FFX/RST ;
  wire \DLX_IFinst_IR_latched<15>/FFX/RST ;
  wire \DLX_IFinst_IR_latched<16>/FFX/RST ;
  wire \DLX_IFinst_IR_latched<24>/FFX/RST ;
  wire \DLX_IFinst_IR_latched<25>/FFX/RST ;
  wire \DLX_IFinst_IR_latched<17>/FFX/RST ;
  wire \DLX_IFinst_IR_latched<26>/FFX/RST ;
  wire \DLX_IFinst_IR_latched<18>/FFX/RST ;
  wire \DLX_IFinst_IR_latched<27>/FFX/RST ;
  wire \DLX_IFinst_IR_latched<19>/FFX/RST ;
  wire \DLX_IFinst_IR_latched<28>/FFX/RST ;
  wire \DLX_IFinst_IR_latched<29>/FFX/RST ;
  wire \DLX_IFinst_IR_latched<7>/FFX/RST ;
  wire \DLX_IFinst_IR_latched<8>/FFX/RST ;
  wire \DLX_IFinst_IR_latched<9>/FFX/RST ;
  wire \DLX_IFinst_PC<1>/FFY/RST ;
  wire \DLX_EXinst_ALU_result<19>/FFY/RST ;
  wire \DLX_IDinst_reg_out_A<8>/FFY/RST ;
  wire \DLX_IDinst_reg_out_A<9>/FFY/RST ;
  wire \DLX_IDinst_IR_opcode_field<1>/FFY/RST ;
  wire \DLX_IDinst_Imm<11>/FFY/RST ;
  wire \DLX_IDinst_delay_slot/FFY/RST ;
  wire \DLX_EXinst_reg_out_B_EX<30>/FFY/RST ;
  wire \DLX_MEMinst_RF_data_in<15>/FFX/RST ;
  wire \DLX_MEMinst_RF_data_in<25>/FFX/RST ;
  wire \DLX_MEMinst_RF_data_in<17>/FFX/RST ;
  wire \DLX_MEMinst_RF_data_in<27>/FFX/RST ;
  wire \DLX_EXinst_mem_to_reg_EX/FFX/RST ;
  wire \DLX_IDinst_EPC<9>/FFX/RST ;
  wire \DLX_IDinst_reg_out_B_2_1/FFY/RST ;
  wire \DLX_IDinst_reg_out_B<3>/FFY/RST ;
  wire \DLX_EXinst_ALU_result<13>/FFY/RST ;
  wire \DLX_IDinst_reg_out_B<3>/FFX/RST ;
  wire \DLX_EXinst_ALU_result<13>/FFX/RST ;
  wire \DLX_IDinst_current_IR<7>/FFX/RST ;
  wire \DLX_IDinst_EPC<1>/FFY/RST ;
  wire \DLX_IDinst_current_IR<9>/FFX/RST ;
  wire \DLX_IDinst_EPC<1>/FFX/RST ;
  wire \DLX_IDinst_EPC<3>/FFY/RST ;
  wire \DLX_IDinst_EPC<3>/FFX/RST ;
  wire \DLX_IDinst_EPC<5>/FFY/RST ;
  wire \DLX_IDinst_EPC<5>/FFX/RST ;
  wire \DLX_IDinst_EPC<7>/FFY/RST ;
  wire \DLX_IDinst_EPC<7>/FFX/RST ;
  wire \DLX_IDinst_EPC<9>/FFY/RST ;
  wire \DLX_IDinst_current_IR<1>/FFY/RST ;
  wire \DLX_IDinst_current_IR<3>/FFY/RST ;
  wire \DLX_IDinst_current_IR<1>/FFX/RST ;
  wire \DLX_IDinst_current_IR<5>/FFY/RST ;
  wire \DLX_IDinst_current_IR<3>/FFX/RST ;
  wire \DLX_IDinst_current_IR<7>/FFY/RST ;
  wire \DLX_IDinst_current_IR<5>/FFX/RST ;
  wire \DLX_IDinst_current_IR<9>/FFY/RST ;
  wire \DLX_IDinst_slot_num_FFd1/FFY/RST ;
  wire \DLX_IDinst_Cause_Reg<1>/FFY/RST ;
  wire \DLX_EXinst_reg_write_EX/FFY/RST ;
  wire \DLX_IDinst_Cause_Reg<3>/FFY/RST ;
  wire \DLX_EXinst_reg_write_EX/FFX/RST ;
  wire \DLX_IDinst_Cause_Reg<1>/FFX/RST ;
  wire \DLX_IDinst_Cause_Reg<3>/FFX/RST ;
  wire \DLX_IDinst_Cause_Reg<5>/FFY/RST ;
  wire \DLX_IDinst_Cause_Reg<5>/FFX/RST ;
  wire \DLX_IDinst_Cause_Reg<7>/FFY/RST ;
  wire \DLX_IDinst_EPC<11>/FFX/RST ;
  wire \DLX_IDinst_EPC<13>/FFX/RST ;
  wire \DLX_IDinst_EPC<21>/FFY/RST ;
  wire \DLX_IDinst_EPC<21>/FFX/RST ;
  wire \DLX_IDinst_EPC<15>/FFY/RST ;
  wire \DLX_IDinst_EPC<15>/FFX/RST ;
  wire \DLX_IDinst_EPC<23>/FFY/RST ;
  wire \DLX_IDinst_EPC<23>/FFX/RST ;
  wire \DLX_IDinst_EPC<25>/FFY/RST ;
  wire \DLX_IDinst_EPC<31>/FFY/RST ;
  wire \DLX_IDinst_EPC<31>/FFX/RST ;
  wire \DLX_IDinst_EPC<17>/FFY/RST ;
  wire \DLX_MEMinst_RF_data_in<19>/FFX/RST ;
  wire \DLX_MEMinst_RF_data_in<29>/FFX/RST ;
  wire \DLX_IDinst_current_IR<20>/FFY/RST ;
  wire \DLX_IDinst_current_IR<11>/FFX/RST ;
  wire \DLX_IDinst_current_IR<15>/FFY/RST ;
  wire \DLX_IDinst_current_IR<13>/FFY/RST ;
  wire \DLX_IDinst_current_IR<13>/FFX/RST ;
  wire \DLX_IDinst_current_IR<21>/FFX/RST ;
  wire \DLX_IDinst_current_IR<17>/FFX/RST ;
  wire \DLX_IDinst_current_IR<26>/FFX/RST ;
  wire \DLX_IDinst_current_IR<19>/FFY/RST ;
  wire \DLX_IDinst_current_IR<19>/FFX/RST ;
  wire \DLX_IDinst_current_IR<27>/FFX/RST ;
  wire \DLX_IDinst_current_IR<28>/FFX/RST ;
  wire \DLX_IDinst_current_IR<29>/FFX/RST ;
  wire \DLX_IDinst_EPC<11>/FFY/RST ;
  wire \DLX_IDinst_EPC<13>/FFY/RST ;
  wire \DLX_IDinst_current_IR<23>/FFY/RST ;
  wire \DLX_IDinst_current_IR<15>/FFX/RST ;
  wire \DLX_IDinst_current_IR<23>/FFX/RST ;
  wire \DLX_IDinst_current_IR<30>/FFX/RST ;
  wire \DLX_IDinst_current_IR<31>/FFX/RST ;
  wire \DLX_IDinst_current_IR<24>/FFX/RST ;
  wire \DLX_IDinst_current_IR<17>/FFY/RST ;
  wire \DLX_IDinst_current_IR<25>/FFY/RST ;
  wire \DLX_IDinst_Cause_Reg<7>/FFX/RST ;
  wire \DLX_IDinst_Cause_Reg<9>/FFY/RST ;
  wire \DLX_IDinst_Cause_Reg<9>/FFX/RST ;
  wire \DLX_EXinst_reg_out_B_EX<11>/FFY/RST ;
  wire \DLX_EXinst_reg_out_B_EX<11>/FFX/RST ;
  wire \DLX_IDinst_IR_function_field<0>/FFY/RST ;
  wire \DLX_EXinst_reg_out_B_EX<13>/FFY/RST ;
  wire \DLX_EXinst_reg_out_B_EX<13>/FFX/RST ;
  wire \DLX_IDinst_IR_function_field<0>/FFX/RST ;
  wire \DLX_EXinst_reg_out_B_EX<21>/FFY/RST ;
  wire \DLX_EXinst_reg_out_B_EX<23>/FFY/RST ;
  wire \DLX_EXinst_reg_out_B_EX<21>/FFX/RST ;
  wire \DLX_IDinst_EPC<17>/FFX/RST ;
  wire \DLX_IDinst_EPC<25>/FFX/RST ;
  wire \DLX_IDinst_EPC<19>/FFY/RST ;
  wire \DLX_IDinst_EPC<19>/FFX/RST ;
  wire \DLX_IDinst_EPC<27>/FFY/RST ;
  wire \DLX_IDinst_EPC<27>/FFX/RST ;
  wire \DLX_IDinst_EPC<29>/FFY/RST ;
  wire \DLX_IDinst_EPC<29>/FFX/RST ;
  wire \DLX_IDinst_counter<1>/FFY/RST ;
  wire \DLX_EXinst_reg_out_B_EX<19>/FFX/RST ;
  wire \DLX_EXinst_reg_out_B_EX<27>/FFY/RST ;
  wire \DLX_EXinst_reg_out_B_EX<27>/FFX/RST ;
  wire \DLX_IDinst_IR_function_field<2>/FFY/RST ;
  wire \DLX_EXinst_reg_out_B_EX<29>/FFY/RST ;
  wire \DLX_EXinst_reg_out_B_EX<29>/FFX/RST ;
  wire \DLX_IDinst_IR_function_field<2>/FFX/RST ;
  wire \DLX_IDinst_IR_function_field<3>/FFY/RST ;
  wire \DLX_IDinst_reg_out_B<21>/FFY/RST ;
  wire \DLX_IDinst_reg_out_B<11>/FFY/RST ;
  wire \DLX_IDinst_IR_function_field<3>/FFX/RST ;
  wire \DLX_EXinst_reg_out_B_EX<23>/FFX/RST ;
  wire \DLX_EXinst_reg_out_B_EX<14>/FFY/RST ;
  wire \DLX_EXinst_reg_out_B_EX<25>/FFX/RST ;
  wire \DLX_IDinst_IR_function_field<1>/FFY/RST ;
  wire \DLX_EXinst_reg_out_B_EX<25>/FFY/RST ;
  wire \DLX_IDinst_IR_function_field<1>/FFX/RST ;
  wire \DLX_EXinst_reg_out_B_EX<17>/FFY/RST ;
  wire \DLX_EXinst_reg_out_B_EX<17>/FFX/RST ;
  wire \DLX_EXinst_reg_out_B_EX<19>/FFY/RST ;
  wire \DLX_IDinst_reg_out_B<29>/FFX/RST ;
  wire \DLX_IDinst_Imm<8>/FFY/RST ;
  wire \DLX_EXinst_ALU_result<2>/FFY/RST ;
  wire \DLX_IDinst_IR_opcode_field<2>/FFY/RST ;
  wire \DLX_IDinst_IR_opcode_field<2>/FFX/RST ;
  wire \DLX_RF_data_in<1>/FFX/RST ;
  wire \DLX_IDinst_Imm<8>/FFX/RST ;
  wire \DLX_RF_data_in<3>/FFY/RST ;
  wire \DLX_RF_data_in<1>/FFY/RST ;
  wire \DLX_IDinst_Imm<10>/FFY/RST ;
  wire \DLX_IDinst_reg_out_B<15>/FFX/RST ;
  wire \DLX_IDinst_reg_out_B<25>/FFY/RST ;
  wire \DLX_IDinst_reg_out_B<25>/FFX/RST ;
  wire \DLX_IDinst_reg_out_B<17>/FFY/RST ;
  wire \DLX_IDinst_reg_out_B<17>/FFX/RST ;
  wire \DLX_IDinst_reg_out_B<27>/FFY/RST ;
  wire \DLX_IDinst_reg_out_B<27>/FFX/RST ;
  wire \DLX_IDinst_reg_out_B<19>/FFY/RST ;
  wire \DLX_IDinst_reg_out_B<29>/FFY/RST ;
  wire \DLX_IDinst_reg_out_B<19>/FFX/RST ;
  wire \DLX_IDinst_Imm<10>/FFX/RST ;
  wire \DLX_RF_data_in<3>/FFX/RST ;
  wire \DLX_RF_data_in<5>/FFY/RST ;
  wire \DLX_RF_data_in<5>/FFX/RST ;
  wire \DLX_RF_data_in<7>/FFY/RST ;
  wire \DLX_RF_data_in<7>/FFX/RST ;
  wire \DLX_MEMinst_RF_data_in<9>/FFY/RST ;
  wire \DLX_MEMinst_RF_data_in<9>/FFX/RST ;
  wire \DLX_EXinst_word/FFY/RST ;
  wire \DLX_IDinst_reg_out_B<5>/FFX/RST ;
  wire \DLX_IDinst_reg_out_B<7>/FFY/RST ;
  wire \DLX_IDinst_reg_out_B<7>/FFX/RST ;
  wire \DLX_IDinst_reg_out_B<9>/FFY/RST ;
  wire \DLX_IDinst_reg_out_B<9>/FFX/RST ;
  wire \DLX_IDinst_rt_addr<1>/FFY/RST ;
  wire \DLX_IDinst_rt_addr<3>/FFX/RST ;
  wire \DLX_IDinst_rt_addr<3>/FFY/RST ;
  wire \DLX_IDinst_mem_read/FFY/RST ;
  wire \DLX_IDinst_IR_opcode_field<5>/FFX/RST ;
  wire \DLX_EXinst_word/FFX/RST ;
  wire \DLX_IFinst_stalled/FFY/RST ;
  wire \DLX_IDinst_rd_addr<3>/FFX/RST ;
  wire \DLX_IDinst_rd_addr<4>/FFY/RST ;
  wire \DLX_IDinst_rd_addr<4>/FFX/RST ;
  wire \DLX_IDinst_rd_addr<3>/FFY/RST ;
  wire \DLX_IDinst_reg_out_B<5>/FFY/RST ;
  wire \DLX_IDinst_reg_out_B<1>/FFY/RST ;
  wire \DLX_IDinst_Cause_Reg<11>/FFY/RST ;
  wire \DLX_IDinst_Cause_Reg<11>/FFX/RST ;
  wire \DLX_IDinst_Cause_Reg<13>/FFY/RST ;
  wire \DLX_IDinst_Cause_Reg<13>/FFX/RST ;
  wire \DLX_IDinst_Cause_Reg<21>/FFY/RST ;
  wire \DLX_IDinst_Cause_Reg<21>/FFX/RST ;
  wire \DLX_IDinst_mem_write/FFY/RST ;
  wire \DLX_IDinst_Cause_Reg<15>/FFY/RST ;
  wire \DLX_IDinst_Cause_Reg<15>/FFX/RST ;
  wire \DLX_IDinst_Cause_Reg<23>/FFY/RST ;
  wire \DLX_IDinst_Cause_Reg<23>/FFX/RST ;
  wire \DLX_IDinst_Cause_Reg<31>/FFY/RST ;
  wire \DLX_IDinst_Cause_Reg<31>/FFX/RST ;
  wire \DLX_IDinst_Cause_Reg<17>/FFY/RST ;
  wire \DLX_IDinst_Cause_Reg<17>/FFX/RST ;
  wire \DLX_IDinst_Cause_Reg<25>/FFY/RST ;
  wire \DLX_IDinst_Cause_Reg<25>/FFX/RST ;
  wire \DLX_IDinst_Cause_Reg<19>/FFY/RST ;
  wire \DLX_IDinst_Cause_Reg<19>/FFX/RST ;
  wire \DLX_IDinst_Cause_Reg<27>/FFY/RST ;
  wire \DLX_IDinst_Cause_Reg<27>/FFX/RST ;
  wire \DLX_IDinst_Cause_Reg<29>/FFY/RST ;
  wire \DLX_EXinst_reg_out_B_EX<5>/FFX/RST ;
  wire \DLX_EXinst_reg_out_B_EX<3>/FFY/RST ;
  wire \DLX_IDinst_Cause_Reg<29>/FFX/RST ;
  wire \DLX_EXinst_reg_out_B_EX<1>/FFY/RST ;
  wire \DLX_EXinst_reg_out_B_EX<1>/FFX/RST ;
  wire \DLX_EXinst_reg_out_B_EX<3>/FFX/RST ;
  wire \DLX_EXinst_reg_out_B_EX<5>/FFY/RST ;
  wire \DLX_EXinst_reg_out_B_EX<7>/FFX/RST ;
  wire \DLX_EXinst_reg_out_B_EX<7>/FFY/RST ;
  wire \DLX_EXinst_reg_out_B_EX<9>/FFY/RST ;
  wire \DLX_EXinst_reg_dst_out<1>/FFY/RST ;
  wire \DLX_IDinst_reg_out_A<29>/FFY/RST ;
  wire \DLX_EXinst_reg_out_B_EX<9>/FFX/RST ;
  wire \DLX_EXinst_reg_dst_out<1>/FFX/RST ;
  wire \DLX_EXinst_reg_dst_out<3>/FFX/RST ;
  wire \DLX_IDinst_IR_function_field<5>/FFX/RST ;
  wire \DLX_IDinst_reg_out_A<28>/FFY/RST ;
  wire \DLX_IDinst_reg_out_A<5>/FFY/RST ;
  wire \DLX_IDinst_reg_out_A<7>/FFY/RST ;
  wire \DLX_IDinst_IR_opcode_field<3>/FFY/RST ;
  wire \DLX_IFinst_PC<3>/FFY/RST ;
  wire \DLX_IFinst_PC<1>/FFX/RST ;
  wire \DLX_IFinst_PC<5>/FFY/RST ;
  wire \DLX_IFinst_PC<3>/FFX/RST ;
  wire \DLX_IFinst_PC<7>/FFY/RST ;
  wire \DLX_IFinst_PC<5>/FFX/RST ;
  wire \DLX_IFinst_PC<7>/FFX/RST ;
  wire \DLX_IFinst_PC<9>/FFX/RST ;
  wire \DLX_IDinst_Imm_31_1/FFY/RST ;
  wire \DLX_IDinst_Imm_31_1/FFX/RST ;
  wire \DLX_IDinst_branch_sig/FFY/RST ;
  wire \DLX_EXinst_ALU_result<24>/FFY/RST ;
  wire \DLX_EXinst_ALU_result<21>/FFY/RST ;
  wire \DLX_MEMinst_noop/FFY/SET ;
  wire \DLX_IFinst_NPC<13>/FFY/RST ;
  wire \DLX_IFinst_NPC<21>/FFY/RST ;
  wire \DLX_IDinst_rt_addr<0>/FFY/RST ;
  wire \DLX_IDinst_IR_opcode_field<4>/FFY/RST ;
  wire \DLX_EXinst_ALU_result<0>/FFY/RST ;
  wire \DLX_EXinst_ALU_result<1>/FFY/RST ;
  wire \DLX_EXinst_reg_out_B_EX<15>/FFY/RST ;
  wire \DLX_EXinst_reg_out_B_EX<31>/FFY/RST ;
  wire \DLX_IFinst_PC<11>/FFY/RST ;
  wire \DLX_IDinst_branch_address<0>/FFY/RST ;
  wire \DLX_EXinst_ALU_result<17>/FFY/RST ;
  wire \DLX_EXinst_ALU_result<25>/FFY/RST ;
  wire \DLX_IFinst_PC<11>/FFX/RST ;
  wire \DLX_IFinst_PC<21>/FFY/RST ;
  wire \DLX_IFinst_PC<21>/FFX/RST ;
  wire \DLX_IFinst_PC<13>/FFX/RST ;
  wire \DLX_IFinst_PC<31>/FFX/RST ;
  wire \DLX_IFinst_PC<31>/FFY/RST ;
  wire \DLX_IFinst_PC<23>/FFX/RST ;
  wire \DLX_IFinst_PC<15>/FFX/RST ;
  wire \DLX_IFinst_PC<25>/FFY/RST ;
  wire \DLX_IFinst_PC<25>/FFX/RST ;
  wire \DLX_IDinst_slot_num_FFd2/FFY/RST ;
  wire \DLX_IFinst_PC<17>/FFX/RST ;
  wire \DLX_IFinst_PC<27>/FFY/RST ;
  wire \DLX_IFinst_PC<27>/FFX/RST ;
  wire \DLX_IFinst_PC<19>/FFX/RST ;
  wire \DLX_IFinst_PC<29>/FFY/RST ;
  wire \DLX_IFinst_PC<29>/FFX/RST ;
  wire \DLX_IDinst_branch_address<1>/FFY/RST ;
  wire \DLX_IDinst_branch_address<2>/FFY/RST ;
  wire \DLX_IDinst_branch_address<3>/FFY/RST ;
  wire \DLX_IDinst_branch_address<4>/FFY/RST ;
  wire \DLX_IDinst_branch_address<5>/FFY/RST ;
  wire \DLX_IDinst_branch_address<6>/FFY/RST ;
  wire \DLX_IDinst_branch_address<7>/FFY/RST ;
  wire \DLX_IDinst_branch_address<8>/FFY/RST ;
  wire \DLX_IDinst_rd_addr<0>/FFY/RST ;
  wire \DLX_IDinst_branch_address<9>/FFY/RST ;
  wire \DLX_IDinst_Imm<12>/FFY/RST ;
  wire \DLX_IDinst_Imm<5>/FFY/RST ;
  wire \DLX_IDinst_Imm<13>/FFY/RST ;
  wire \DLX_IDinst_Imm<14>/FFY/RST ;
  wire \DLX_IDinst_Imm<15>/FFY/RST ;
  wire \DLX_EXinst_ALU_result<3>/FFY/RST ;
  wire \DLX_IDinst_reg_out_B<0>/FFY/RST ;
  wire \DLX_EXinst_ALU_result<4>/FFY/RST ;
  wire \DLX_EXinst_ALU_result<5>/FFY/RST ;
  wire \DLX_EXinst_ALU_result<22>/FFY/RST ;
  wire \DLX_EXinst_ALU_result<6>/FFY/RST ;
  wire \DLX_EXinst_ALU_result<7>/FFY/RST ;
  wire \DLX_IDinst_branch_address<11>/FFY/RST ;
  wire \DLX_IDinst_mem_to_reg/FFY/RST ;
  wire \DLX_IDinst_branch_address<10>/FFY/RST ;
  wire \DLX_EXinst_ALU_result<8>/FFY/RST ;
  wire \DLX_IDinst_branch_address<12>/FFY/RST ;
  wire \DLX_IDinst_branch_address<20>/FFY/RST ;
  wire \DLX_EXinst_ALU_result<9>/FFY/RST ;
  wire \DLX_EXinst_ALU_result<18>/FFY/RST ;
  wire \DLX_EXinst_ALU_result<26>/FFY/RST ;
  wire \DLX_IDinst_CLI/FFY/RST ;
  wire \DLX_EXinst_noop/FFY/SET ;
  wire \DLX_IDinst_branch_address<14>/FFY/RST ;
  wire \DLX_IDinst_branch_address<30>/FFY/RST ;
  wire \DLX_IDinst_branch_address<22>/FFY/RST ;
  wire \DLX_IDinst_branch_address<21>/FFY/RST ;
  wire \DLX_IDinst_branch_address<13>/FFY/RST ;
  wire \DLX_IDinst_stall/FFY/RST ;
  wire \DLX_IDinst_branch_address<17>/FFY/RST ;
  wire \DLX_IDinst_branch_address<25>/FFY/RST ;
  wire \DLX_IFinst_NPC<10>/FFY/RST ;
  wire \DLX_IDinst_branch_address<31>/FFY/RST ;
  wire \DLX_IFinst_NPC<20>/FFY/RST ;
  wire \DLX_IFinst_NPC<12>/FFY/RST ;
  wire \DLX_IFinst_NPC<0>/FFY/RST ;
  wire \DLX_IDinst_branch_address<23>/FFY/RST ;
  wire \DLX_IDinst_branch_address<15>/FFY/RST ;
  wire \DLX_IDinst_branch_address<16>/FFY/RST ;
  wire \DLX_IDinst_branch_address<24>/FFY/RST ;
  wire \DLX_IDinst_branch_address<26>/FFY/RST ;
  wire \DLX_IDinst_branch_address<18>/FFY/RST ;
  wire \DLX_IDinst_branch_address<27>/FFY/RST ;
  wire \DLX_IDinst_branch_address<19>/FFY/RST ;
  wire \DLX_IDinst_branch_address<28>/FFY/RST ;
  wire \DLX_EXinst_ALU_result<14>/FFY/RST ;
  wire \DLX_IDinst_branch_address<29>/FFY/RST ;
  wire \DLX_IFinst_NPC<11>/FFY/RST ;
  wire \DLX_IFinst_NPC<1>/FFY/RST ;
  wire \DLX_IFinst_NPC<4>/FFY/RST ;
  wire \DLX_EXinst_ALU_result<27>/FFY/RST ;
  wire \DLX_EXinst_ALU_result<15>/FFY/RST ;
  wire \DLX_MEMinst_reg_dst_out<1>/FFY/RST ;
  wire \DLX_MEMinst_reg_dst_out<1>/FFX/RST ;
  wire \DLX_EXinst_ALU_result<31>/FFY/RST ;
  wire \DLX_EXinst_ALU_result<10>/FFY/RST ;
  wire \DLX_IFinst_NPC<30>/FFY/RST ;
  wire \DLX_IFinst_NPC<14>/FFY/RST ;
  wire \DLX_IFinst_NPC<22>/FFY/RST ;
  wire \DLX_IDinst_reg_dst/FFY/RST ;
  wire \DLX_EXinst_ALU_result<11>/FFY/RST ;
  wire \DLX_IFinst_NPC<2>/FFY/RST ;
  wire \DLX_EXinst_ALU_result<20>/FFY/RST ;
  wire \DLX_EXinst_ALU_result<23>/FFY/RST ;
  wire \DLX_IFinst_NPC<15>/FFY/RST ;
  wire \DLX_IFinst_NPC<31>/FFY/RST ;
  wire \DLX_IFinst_NPC<23>/FFY/RST ;
  wire \DLX_IFinst_NPC<3>/FFY/RST ;
  wire \DLX_MEMinst_reg_dst_out<3>/FFY/RST ;
  wire \DLX_MEMinst_reg_dst_out<3>/FFX/RST ;
  wire \DLX_MEMinst_reg_dst_out<4>/FFY/RST ;
  wire \DLX_IDinst_slot_num_FFd3/FFY/SET ;
  wire \DLX_IDinst_reg_out_B<2>/FFY/RST ;
  wire \DLX_IFinst_NPC<24>/FFY/RST ;
  wire \DLX_IFinst_NPC<16>/FFY/RST ;
  wire \DLX_EXinst_ALU_result<30>/FFY/RST ;
  wire \DLX_IFinst_NPC<26>/FFY/RST ;
  wire \DLX_IFinst_NPC<18>/FFY/RST ;
  wire \DLX_IFinst_NPC<17>/FFY/RST ;
  wire \DLX_IFinst_NPC<25>/FFY/RST ;
  wire \DLX_EXinst_ALU_result<16>/FFY/RST ;
  wire \DLX_IDinst_reg_out_A<21>/FFY/RST ;
  wire \DLX_IDinst_reg_out_A<13>/FFY/RST ;
  wire \DLX_IFinst_NPC<5>/FFY/RST ;
  wire \DLX_IFinst_NPC<6>/FFY/RST ;
  wire \DLX_IDinst_reg_write/FFY/RST ;
  wire \DLX_IDinst_counter<0>/FFY/RST ;
  wire \DLX_EXinst_ALU_result<28>/FFY/RST ;
  wire \DLX_IFinst_NPC<19>/FFY/RST ;
  wire \DLX_IFinst_NPC<27>/FFY/RST ;
  wire \DLX_IFinst_NPC<7>/FFY/RST ;
  wire \DLX_EXinst_ALU_result<29>/FFY/RST ;
  wire \DLX_IFinst_NPC<28>/FFY/RST ;
  wire \DLX_IFinst_NPC<8>/FFY/RST ;
  wire \DLX_IFinst_NPC<29>/FFY/RST ;
  wire \DLX_IDinst_reg_out_A<11>/FFY/RST ;
  wire \DLX_IDinst_reg_out_A<12>/FFY/RST ;
  wire \DLX_IDinst_reg_out_A<20>/FFY/RST ;
  wire \DLX_MEMinst_reg_write_MEM/FFY/RST ;
  wire \DLX_IFinst_NPC<9>/FFY/RST ;
  wire \DLX_IDinst_reg_out_A<10>/FFY/RST ;
  wire \DLX_IDinst_reg_out_A<14>/FFY/RST ;
  wire \DLX_IDinst_reg_out_A<22>/FFY/RST ;
  wire \DLX_IDinst_reg_out_A<30>/FFY/RST ;
  wire \DLX_IDinst_reg_out_A<23>/FFY/RST ;
  wire \DLX_IDinst_reg_out_A<31>/FFY/RST ;
  wire \DLX_IDinst_reg_out_A<15>/FFY/RST ;
  wire \DLX_IDinst_reg_out_A<0>/FFY/RST ;
  wire \DLX_IDinst_reg_out_A<24>/FFY/RST ;
  wire \DLX_IDinst_reg_out_A<16>/FFY/RST ;
  wire \DLX_IDinst_reg_out_A<1>/FFY/RST ;
  wire \DLX_IDinst_reg_out_A<17>/FFY/RST ;
  wire \DLX_IDinst_reg_out_A<25>/FFY/RST ;
  wire \DLX_IDinst_reg_out_A<2>/FFY/RST ;
  wire \DLX_IDinst_reg_out_A<26>/FFY/RST ;
  wire \DLX_IDinst_reg_out_A<18>/FFY/RST ;
  wire \DLX_IDinst_reg_out_A<3>/FFY/RST ;
  wire \DLX_IDinst_reg_out_A<27>/FFY/RST ;
  wire \DLX_IDinst_reg_out_A<19>/FFY/RST ;
  wire \DLX_IDinst_reg_out_A<4>/FFY/RST ;
  wire \DLX_clkbuf2/CE ;
  wire \DLX_clkbuf3/CE ;
  wire \clkbuf2/CE ;
  wire \clkbuf3/CE ;
  wire \PWR_VCC_0/FROM ;
  wire \PWR_VCC_0/GROM ;
  wire \PWR_VCC_1/FROM ;
  wire \PWR_VCC_1/GROM ;
  wire \PWR_VCC_2/FROM ;
  wire \PWR_VCC_2/GROM ;
  wire \PWR_VCC_3/FROM ;
  wire \PWR_VCC_3/GROM ;
  wire \PWR_VCC_4/FROM ;
  wire \PWR_VCC_4/GROM ;
  wire \PWR_GND_0/GROM ;
  wire \PWR_GND_1/GROM ;
  wire \PWR_GND_2/GROM ;
  wire \PWR_GND_3/GROM ;
  wire \PWR_GND_4/GROM ;
  wire \PWR_GND_5/GROM ;
  wire \PWR_GND_6/GROM ;
  wire VCC;
  wire GND;
  wire \NLW_Mmux__COND_2_inst_mux_f6_0.F51_IA_UNCONNECTED ;
  wire [0 : 0] DM_write_data;
  wire [31 : 0] DLX_IFinst__n0001;
  wire [31 : 0] DLX_EXinst__n0007;
  wire [4 : 0] DLX_IDinst_regA_index;
  wire [4 : 0] DLX_MEMinst_reg_dst_out;
  wire [7 : 0] DLX_RF_data_in;
  wire [31 : 8] DLX_IDinst_WB_data_eff;
  wire [31 : 0] DLX_IDinst_reg_out_A_RF;
  wire [4 : 0] DLX_IDinst_regB_index;
  wire [31 : 0] DLX_IDinst_reg_out_B_RF;
  wire [31 : 0] DLX_EXinst_ALU_result;
  wire [31 : 0] DLX_IFinst_NPC;
  wire [31 : 0] DLX_EXinst_reg_out_B_EX;
  wire [31 : 0] RAM_read_data;
  wire [23 : 0] IR;
  wire [5 : 0] vga_select_6;
  wire [14 : 6] vga_address;
  wire [8 : 0] vga_top_vga1_gridhcounter;
  wire [4 : 0] vram_out_cpu;
  wire [4 : 0] vram_out_vga;
  wire [31 : 0] DLX_IDinst_reg_out_B;
  wire [31 : 0] DLX_IDinst_reg_out_A;
  wire [31 : 26] DLX_IDinst_IR_latched;
  wire [5 : 0] DLX_IDinst_IR_function_field;
  wire [31 : 0] DLX_IFinst_IR_previous;
  wire [31 : 0] DLX_IFinst_IR_curr;
  wire [31 : 0] DLX_IFinst_IR_latched;
  wire [8 : 0] vga_top_vga1_gridvcounter;
  wire [4 : 0] DLX_reg_dst_of_EX;
  wire [4 : 0] DLX_IDinst_rt_addr;
  wire [4 : 0] DLX_IDinst_rd_addr;
  wire [4 : 0] DLX_reg_dst_of_MEM;
  wire [5 : 0] DLX_IDinst_IR_opcode_field;
  wire [4 : 0] DLX_EXinst_reg_dst_out;
  wire [15 : 0] DLX_IDinst_jtarget;
  wire [31 : 1] DLX_IDinst__n0129;
  wire [31 : 0] DLX_IDinst_current_IR;
  wire [9 : 0] vga_top_vga1_vcounter;
  wire [15 : 0] vga_top_vga1_hcounter;
  wire [31 : 0] DLX_EXinst__n0017;
  wire [31 : 0] DLX_EXinst__n0016;
  wire [31 : 3] DLX_IFinst__n0015;
  wire [31 : 0] DLX_IDinst__n0128;
  wire [1 : 0] DLX_IDinst_counter;
  wire [31 : 0] DLX_IDinst_EPC;
  wire [2 : 0] vga_top_vga1_helpcounter;
  wire [31 : 0] DLX_IDinst_regB_eff;
  wire [31 : 0] DLX_IDinst__n0118;
  wire [31 : 0] DM_read_data;
  wire [31 : 8] DLX_MEMinst_RF_data_in;
  wire [31 : 0] DLX_IDinst_Cause_Reg;
  wire [4 : 0] DLX_IDinst__n0023;
  wire [1 : 1] DLX_IDinst__n0448;
  wire [5 : 5] DLX_IDinst__n0030;
  wire [31 : 0] DLX_IDinst_regA_eff;
  wire [5 : 0] DLX_opcode_of_MEM;
  wire [5 : 0] DLX_opcode_of_WB;
  wire [31 : 0] DLX_IFinst_PC;
  wire [31 : 0] DLX_IDinst_branch_address;
  wire [47 : 40] DLX_IDinst__n0445;
  wire [31 : 0] DLX_IFinst__n0003;
  wire [4 : 0] DLX_EXinst__n0008;
  wire [4 : 0] DLX_IDinst__n0106;
  wire [9 : 1] vga_top_vga1_vcounter__n0000;
  wire [15 : 1] vga_top_vga1_hcounter__n0000;
  wire [8 : 1] vga_top_vga1_gridvcounter__n0000;
  wire [8 : 1] vga_top_vga1_gridhcounter__n0000;
  wire [31 : 0] DLX_IDinst__n0123;
  wire [2 : 1] vga_top_vga1_helpcounter__n0000;
  wire [31 : 0] DLX_MEMinst__n0000;
  wire [1 : 1] DLX_IDinst__n0116;
  wire [31 : 0] DLX_IDinst__n0127;
  wire [5 : 0] DLX_IDinst__n0113;
  wire [4 : 0] DLX_IDinst__n0107;
  wire [5 : 5] DLX_IDinst__n0114;
  assign
    DM_write_data_0 = DM_write_data[0];
  initial $sdf_annotate("DLX_top_timesim.sdf");
  X_OPAD \mask<1>/PAD  (
    .PAD(mask[1])
  );
  X_TRI mask_1_OBUF_0 (
    .I(\mask<1>/OUTMUX ),
    .CTL(\mask<1>/ENABLE ),
    .O(mask[1])
  );
  X_INV \mask<1>/ENABLEINV  (
    .I(\mask<1>/TORGTS ),
    .O(\mask<1>/ENABLE )
  );
  X_BUF \mask<1>/GTS_OR  (
    .I(GTS),
    .O(\mask<1>/TORGTS )
  );
  X_BUF \mask<1>/OUTMUX_1  (
    .I(mask_1_OBUF),
    .O(\mask<1>/OUTMUX )
  );
  X_OR2 \DM_write/OFF/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DM_write/OFF/RST )
  );
  defparam DLX_EXinst_mem_write_EX_1_2.INIT = 1'b0;
  X_FF DLX_EXinst_mem_write_EX_1_2 (
    .I(\DM_write/OD ),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DM_write/OFF/RST ),
    .O(DLX_EXinst_mem_write_EX_1)
  );
  X_OPAD \DM_write/PAD  (
    .PAD(DM_write)
  );
  X_TRI DM_write_OBUF (
    .I(\DM_write/OUTMUX ),
    .CTL(\DM_write/ENABLE ),
    .O(DM_write)
  );
  X_INV \DM_write/ENABLEINV  (
    .I(\DM_write/TORGTS ),
    .O(\DM_write/ENABLE )
  );
  X_BUF \DM_write/GTS_OR  (
    .I(GTS),
    .O(\DM_write/TORGTS )
  );
  X_BUF \DM_write/OUTMUX_3  (
    .I(DLX_EXinst_mem_write_EX_1),
    .O(\DM_write/OUTMUX )
  );
  X_BUF \DM_write/OMUX  (
    .I(DLX_EXinst__n0012),
    .O(\DM_write/OD )
  );
  X_OPAD \mask<2>/PAD  (
    .PAD(mask[2])
  );
  X_TRI mask_2_OBUF_4 (
    .I(\mask<2>/OUTMUX ),
    .CTL(\mask<2>/ENABLE ),
    .O(mask[2])
  );
  X_INV \mask<2>/ENABLEINV  (
    .I(\mask<2>/TORGTS ),
    .O(\mask<2>/ENABLE )
  );
  X_BUF \mask<2>/GTS_OR  (
    .I(GTS),
    .O(\mask<2>/TORGTS )
  );
  X_BUF \mask<2>/OUTMUX_5  (
    .I(mask_2_OBUF),
    .O(\mask<2>/OUTMUX )
  );
  X_OPAD \PIPEEMPTY/PAD  (
    .PAD(PIPEEMPTY)
  );
  X_TRI PIPEEMPTY_OBUF_6 (
    .I(\PIPEEMPTY/OUTMUX ),
    .CTL(\PIPEEMPTY/ENABLE ),
    .O(PIPEEMPTY)
  );
  X_INV \PIPEEMPTY/ENABLEINV  (
    .I(\PIPEEMPTY/TORGTS ),
    .O(\PIPEEMPTY/ENABLE )
  );
  X_BUF \PIPEEMPTY/GTS_OR  (
    .I(GTS),
    .O(\PIPEEMPTY/TORGTS )
  );
  X_BUF \PIPEEMPTY/OUTMUX_7  (
    .I(PIPEEMPTY_OBUF),
    .O(\PIPEEMPTY/OUTMUX )
  );
  X_OPAD \clk_IF_del/PAD  (
    .PAD(clk_IF_del)
  );
  X_TRI clk_IF_del_OBUF (
    .I(\clk_IF_del/OUTMUX ),
    .CTL(\clk_IF_del/ENABLE ),
    .O(clk_IF_del)
  );
  X_INV \clk_IF_del/ENABLEINV  (
    .I(\clk_IF_del/TORGTS ),
    .O(\clk_IF_del/ENABLE )
  );
  X_BUF \clk_IF_del/GTS_OR  (
    .I(GTS),
    .O(\clk_IF_del/TORGTS )
  );
  X_BUF \clk_IF_del/OUTMUX_8  (
    .I(DLX_clk_IF_del),
    .O(\clk_IF_del/OUTMUX )
  );
  X_OR2 \DM_addr_eff<10>/OFF/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DM_addr_eff<10>/OFF/RST )
  );
  defparam DLX_EXinst_ALU_result_10_1_9.INIT = 1'b0;
  X_FF DLX_EXinst_ALU_result_10_1_9 (
    .I(\DM_addr_eff<10>/OD ),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DM_addr_eff<10>/OFF/RST ),
    .O(DLX_EXinst_ALU_result_10_1)
  );
  X_OPAD \DM_addr_eff<10>/PAD  (
    .PAD(DM_addr_eff[10])
  );
  X_TRI DM_addr_eff_10_OBUF (
    .I(\DM_addr_eff<10>/OUTMUX ),
    .CTL(\DM_addr_eff<10>/ENABLE ),
    .O(DM_addr_eff[10])
  );
  X_INV \DM_addr_eff<10>/ENABLEINV  (
    .I(\DM_addr_eff<10>/TORGTS ),
    .O(\DM_addr_eff<10>/ENABLE )
  );
  X_BUF \DM_addr_eff<10>/GTS_OR  (
    .I(GTS),
    .O(\DM_addr_eff<10>/TORGTS )
  );
  X_BUF \DM_addr_eff<10>/OUTMUX_10  (
    .I(DLX_EXinst_ALU_result_10_1),
    .O(\DM_addr_eff<10>/OUTMUX )
  );
  X_BUF \DM_addr_eff<10>/OMUX  (
    .I(N116776),
    .O(\DM_addr_eff<10>/OD )
  );
  X_OR2 \DM_addr_eff<11>/OFF/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DM_addr_eff<11>/OFF/RST )
  );
  defparam DLX_EXinst_ALU_result_11_1_11.INIT = 1'b0;
  X_FF DLX_EXinst_ALU_result_11_1_11 (
    .I(\DM_addr_eff<11>/OD ),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DM_addr_eff<11>/OFF/RST ),
    .O(DLX_EXinst_ALU_result_11_1)
  );
  X_OPAD \DM_addr_eff<11>/PAD  (
    .PAD(DM_addr_eff[11])
  );
  X_TRI DM_addr_eff_11_OBUF (
    .I(\DM_addr_eff<11>/OUTMUX ),
    .CTL(\DM_addr_eff<11>/ENABLE ),
    .O(DM_addr_eff[11])
  );
  X_INV \DM_addr_eff<11>/ENABLEINV  (
    .I(\DM_addr_eff<11>/TORGTS ),
    .O(\DM_addr_eff<11>/ENABLE )
  );
  X_BUF \DM_addr_eff<11>/GTS_OR  (
    .I(GTS),
    .O(\DM_addr_eff<11>/TORGTS )
  );
  X_BUF \DM_addr_eff<11>/OUTMUX_12  (
    .I(DLX_EXinst_ALU_result_11_1),
    .O(\DM_addr_eff<11>/OUTMUX )
  );
  X_BUF \DM_addr_eff<11>/OMUX  (
    .I(N113314),
    .O(\DM_addr_eff<11>/OD )
  );
  X_OR2 \DM_addr_eff<12>/OFF/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DM_addr_eff<12>/OFF/RST )
  );
  defparam DLX_EXinst_ALU_result_12_1_13.INIT = 1'b0;
  X_FF DLX_EXinst_ALU_result_12_1_13 (
    .I(\DM_addr_eff<12>/OD ),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DM_addr_eff<12>/OFF/RST ),
    .O(DLX_EXinst_ALU_result_12_1)
  );
  X_OPAD \DM_addr_eff<12>/PAD  (
    .PAD(DM_addr_eff[12])
  );
  X_TRI DM_addr_eff_12_OBUF (
    .I(\DM_addr_eff<12>/OUTMUX ),
    .CTL(\DM_addr_eff<12>/ENABLE ),
    .O(DM_addr_eff[12])
  );
  X_INV \DM_addr_eff<12>/ENABLEINV  (
    .I(\DM_addr_eff<12>/TORGTS ),
    .O(\DM_addr_eff<12>/ENABLE )
  );
  X_BUF \DM_addr_eff<12>/GTS_OR  (
    .I(GTS),
    .O(\DM_addr_eff<12>/TORGTS )
  );
  X_BUF \DM_addr_eff<12>/OUTMUX_14  (
    .I(DLX_EXinst_ALU_result_12_1),
    .O(\DM_addr_eff<12>/OUTMUX )
  );
  X_BUF \DM_addr_eff<12>/OMUX  (
    .I(N112968),
    .O(\DM_addr_eff<12>/OD )
  );
  X_OPAD \DM_addr_eff<13>/PAD  (
    .PAD(DM_addr_eff[13])
  );
  X_TRI DM_addr_eff_13_OBUF (
    .I(\DM_addr_eff<13>/OUTMUX ),
    .CTL(\DM_addr_eff<13>/ENABLE ),
    .O(DM_addr_eff[13])
  );
  X_INV \DM_addr_eff<13>/ENABLEINV  (
    .I(\DM_addr_eff<13>/TORGTS ),
    .O(\DM_addr_eff<13>/ENABLE )
  );
  X_BUF \DM_addr_eff<13>/GTS_OR  (
    .I(GTS),
    .O(\DM_addr_eff<13>/TORGTS )
  );
  X_BUF \DM_addr_eff<13>/OUTMUX_15  (
    .I(DLX_EXinst_ALU_result_13_1),
    .O(\DM_addr_eff<13>/OUTMUX )
  );
  X_BUF \DM_addr_eff<13>/OMUX  (
    .I(N115578),
    .O(\DM_addr_eff<13>/OD )
  );
  X_OPAD \DM_addr_eff<14>/PAD  (
    .PAD(DM_addr_eff[14])
  );
  X_TRI DM_addr_eff_14_OBUF (
    .I(\DM_addr_eff<14>/OUTMUX ),
    .CTL(\DM_addr_eff<14>/ENABLE ),
    .O(DM_addr_eff[14])
  );
  X_INV \DM_addr_eff<14>/ENABLEINV  (
    .I(\DM_addr_eff<14>/TORGTS ),
    .O(\DM_addr_eff<14>/ENABLE )
  );
  X_BUF \DM_addr_eff<14>/GTS_OR  (
    .I(GTS),
    .O(\DM_addr_eff<14>/TORGTS )
  );
  X_BUF \DM_addr_eff<14>/OUTMUX_16  (
    .I(DLX_EXinst_ALU_result_14_1),
    .O(\DM_addr_eff<14>/OUTMUX )
  );
  X_BUF \DM_addr_eff<14>/OMUX  (
    .I(N115216),
    .O(\DM_addr_eff<14>/OD )
  );
  X_OPAD \branch_sig/PAD  (
    .PAD(branch_sig)
  );
  X_TRI branch_sig_OBUF (
    .I(\branch_sig/OUTMUX ),
    .CTL(\branch_sig/ENABLE ),
    .O(branch_sig)
  );
  X_INV \branch_sig/ENABLEINV  (
    .I(\branch_sig/TORGTS ),
    .O(\branch_sig/ENABLE )
  );
  X_BUF \branch_sig/GTS_OR  (
    .I(GTS),
    .O(\branch_sig/TORGTS )
  );
  X_BUF \branch_sig/OUTMUX_17  (
    .I(DLX_IDinst_branch_sig_1),
    .O(\branch_sig/OUTMUX )
  );
  X_BUF \branch_sig/OMUX  (
    .I(N110516),
    .O(\branch_sig/OD )
  );
  X_OPAD \clk_DM/PAD  (
    .PAD(clk_DM)
  );
  X_TRI clk_DM_OBUF_18 (
    .I(\clk_DM/OUTMUX ),
    .CTL(\clk_DM/ENABLE ),
    .O(clk_DM)
  );
  X_INV \clk_DM/ENABLEINV  (
    .I(\clk_DM/TORGTS ),
    .O(\clk_DM/ENABLE )
  );
  X_BUF \clk_DM/GTS_OR  (
    .I(GTS),
    .O(\clk_DM/TORGTS )
  );
  X_BUF \clk_DM/OUTMUX_19  (
    .I(clk_DM_OBUF),
    .O(\clk_DM/OUTMUX )
  );
  X_OPAD \clk_ID/PAD  (
    .PAD(clk_ID)
  );
  X_TRI clk_ID_OBUF (
    .I(\clk_ID/OUTMUX ),
    .CTL(\clk_ID/ENABLE ),
    .O(clk_ID)
  );
  X_INV \clk_ID/ENABLEINV  (
    .I(\clk_ID/TORGTS ),
    .O(\clk_ID/ENABLE )
  );
  X_BUF \clk_ID/GTS_OR  (
    .I(GTS),
    .O(\clk_ID/TORGTS )
  );
  X_BUF \clk_ID/OUTMUX_20  (
    .I(DLX_clk_ID),
    .O(\clk_ID/OUTMUX )
  );
  X_OPAD \clk_IF/PAD  (
    .PAD(clk_IF)
  );
  X_TRI clk_IF_OBUF (
    .I(\clk_IF/OUTMUX ),
    .CTL(\clk_IF/ENABLE ),
    .O(clk_IF)
  );
  X_INV \clk_IF/ENABLEINV  (
    .I(\clk_IF/TORGTS ),
    .O(\clk_IF/ENABLE )
  );
  X_BUF \clk_IF/GTS_OR  (
    .I(GTS),
    .O(\clk_IF/TORGTS )
  );
  X_BUF \clk_IF/OUTMUX_21  (
    .I(DLX_clk_IF),
    .O(\clk_IF/OUTMUX )
  );
  X_OPAD \clk_EX/PAD  (
    .PAD(clk_EX)
  );
  X_TRI clk_EX_OBUF (
    .I(\clk_EX/OUTMUX ),
    .CTL(\clk_EX/ENABLE ),
    .O(clk_EX)
  );
  X_INV \clk_EX/ENABLEINV  (
    .I(\clk_EX/TORGTS ),
    .O(\clk_EX/ENABLE )
  );
  X_BUF \clk_EX/GTS_OR  (
    .I(GTS),
    .O(\clk_EX/TORGTS )
  );
  X_BUF \clk_EX/OUTMUX_22  (
    .I(DLX_clk_EX),
    .O(\clk_EX/OUTMUX )
  );
  X_ZERO \hsync/LOGIC_ZERO_23  (
    .O(\hsync/LOGIC_ZERO )
  );
  X_OPAD \hsync/PAD  (
    .PAD(hsync)
  );
  X_TRI hsync_OBUF (
    .I(\hsync/OUTMUX ),
    .CTL(\hsync/ENABLE ),
    .O(hsync)
  );
  X_INV \hsync/ENABLEINV  (
    .I(\hsync/TORGTS ),
    .O(\hsync/ENABLE )
  );
  X_BUF \hsync/GTS_OR  (
    .I(GTS),
    .O(\hsync/TORGTS )
  );
  X_BUF \hsync/OUTMUX_24  (
    .I(vga_top_vga1_hsyncout),
    .O(\hsync/OUTMUX )
  );
  X_OPAD \green<0>/PAD  (
    .PAD(green[0])
  );
  X_TRI green_0_OBUF_25 (
    .I(\green<0>/OUTMUX ),
    .CTL(\green<0>/ENABLE ),
    .O(green[0])
  );
  X_INV \green<0>/ENABLEINV  (
    .I(\green<0>/TORGTS ),
    .O(\green<0>/ENABLE )
  );
  X_BUF \green<0>/GTS_OR  (
    .I(GTS),
    .O(\green<0>/TORGTS )
  );
  X_BUF \green<0>/OUTMUX_26  (
    .I(green_0_OBUF),
    .O(\green<0>/OUTMUX )
  );
  X_OPAD \green<1>/PAD  (
    .PAD(green[1])
  );
  X_TRI green_1_OBUF_27 (
    .I(\green<1>/OUTMUX ),
    .CTL(\green<1>/ENABLE ),
    .O(green[1])
  );
  X_INV \green<1>/ENABLEINV  (
    .I(\green<1>/TORGTS ),
    .O(\green<1>/ENABLE )
  );
  X_BUF \green<1>/GTS_OR  (
    .I(GTS),
    .O(\green<1>/TORGTS )
  );
  X_BUF \green<1>/OUTMUX_28  (
    .I(green_1_OBUF),
    .O(\green<1>/OUTMUX )
  );
  X_OPAD \green<2>/PAD  (
    .PAD(green[2])
  );
  X_TRI green_2_OBUF_29 (
    .I(\green<2>/OUTMUX ),
    .CTL(\green<2>/ENABLE ),
    .O(green[2])
  );
  X_INV \green<2>/ENABLEINV  (
    .I(\green<2>/TORGTS ),
    .O(\green<2>/ENABLE )
  );
  X_BUF \green<2>/GTS_OR  (
    .I(GTS),
    .O(\green<2>/TORGTS )
  );
  X_BUF \green<2>/OUTMUX_30  (
    .I(green_2_OBUF),
    .O(\green<2>/OUTMUX )
  );
  X_IPAD \reset/PAD  (
    .PAD(reset)
  );
  X_BUF \reset/IMUX  (
    .I(\reset/IBUF ),
    .O(reset_IBUF)
  );
  X_BUF reset_IBUF_31 (
    .I(reset),
    .O(\reset/IBUF )
  );
  X_OPAD \red<0>/PAD  (
    .PAD(red[0])
  );
  X_TRI red_0_OBUF_32 (
    .I(\red<0>/OUTMUX ),
    .CTL(\red<0>/ENABLE ),
    .O(red[0])
  );
  X_INV \red<0>/ENABLEINV  (
    .I(\red<0>/TORGTS ),
    .O(\red<0>/ENABLE )
  );
  X_BUF \red<0>/GTS_OR  (
    .I(GTS),
    .O(\red<0>/TORGTS )
  );
  X_BUF \red<0>/OUTMUX_33  (
    .I(red_0_OBUF),
    .O(\red<0>/OUTMUX )
  );
  X_OPAD \red<1>/PAD  (
    .PAD(red[1])
  );
  X_TRI red_1_OBUF_34 (
    .I(\red<1>/OUTMUX ),
    .CTL(\red<1>/ENABLE ),
    .O(red[1])
  );
  X_INV \red<1>/ENABLEINV  (
    .I(\red<1>/TORGTS ),
    .O(\red<1>/ENABLE )
  );
  X_BUF \red<1>/GTS_OR  (
    .I(GTS),
    .O(\red<1>/TORGTS )
  );
  X_BUF \red<1>/OUTMUX_35  (
    .I(red_1_OBUF),
    .O(\red<1>/OUTMUX )
  );
  X_OPAD \NPC_eff<0>/PAD  (
    .PAD(NPC_eff[0])
  );
  X_TRI NPC_eff_0_OBUF (
    .I(\NPC_eff<0>/OUTMUX ),
    .CTL(\NPC_eff<0>/ENABLE ),
    .O(NPC_eff[0])
  );
  X_INV \NPC_eff<0>/ENABLEINV  (
    .I(\NPC_eff<0>/TORGTS ),
    .O(\NPC_eff<0>/ENABLE )
  );
  X_BUF \NPC_eff<0>/GTS_OR  (
    .I(GTS),
    .O(\NPC_eff<0>/TORGTS )
  );
  X_BUF \NPC_eff<0>/OUTMUX_36  (
    .I(DLX_IFinst_NPC_0_1),
    .O(\NPC_eff<0>/OUTMUX )
  );
  X_BUF \NPC_eff<0>/OMUX  (
    .I(DLX_IFinst__n0001[0]),
    .O(\NPC_eff<0>/OD )
  );
  defparam DLX_EXinst_ALU_result_13_1_37.INIT = 1'b0;
  X_FF DLX_EXinst_ALU_result_13_1_37 (
    .I(\DM_addr_eff<13>/OD ),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DM_addr_eff<13>/OFF/RST ),
    .O(DLX_EXinst_ALU_result_13_1)
  );
  X_OR2 \DM_addr_eff<13>/OFF/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DM_addr_eff<13>/OFF/RST )
  );
  X_OPAD \NPC_eff<1>/PAD  (
    .PAD(NPC_eff[1])
  );
  X_TRI NPC_eff_1_OBUF (
    .I(\NPC_eff<1>/OUTMUX ),
    .CTL(\NPC_eff<1>/ENABLE ),
    .O(NPC_eff[1])
  );
  X_INV \NPC_eff<1>/ENABLEINV  (
    .I(\NPC_eff<1>/TORGTS ),
    .O(\NPC_eff<1>/ENABLE )
  );
  X_BUF \NPC_eff<1>/GTS_OR  (
    .I(GTS),
    .O(\NPC_eff<1>/TORGTS )
  );
  X_BUF \NPC_eff<1>/OUTMUX_38  (
    .I(DLX_IFinst_NPC_1_1),
    .O(\NPC_eff<1>/OUTMUX )
  );
  X_BUF \NPC_eff<1>/OMUX  (
    .I(DLX_IFinst__n0001[1]),
    .O(\NPC_eff<1>/OD )
  );
  X_OPAD \NPC_eff<2>/PAD  (
    .PAD(NPC_eff[2])
  );
  X_TRI NPC_eff_2_OBUF (
    .I(\NPC_eff<2>/OUTMUX ),
    .CTL(\NPC_eff<2>/ENABLE ),
    .O(NPC_eff[2])
  );
  X_INV \NPC_eff<2>/ENABLEINV  (
    .I(\NPC_eff<2>/TORGTS ),
    .O(\NPC_eff<2>/ENABLE )
  );
  X_BUF \NPC_eff<2>/GTS_OR  (
    .I(GTS),
    .O(\NPC_eff<2>/TORGTS )
  );
  X_BUF \NPC_eff<2>/OUTMUX_39  (
    .I(DLX_IFinst_NPC_2_1),
    .O(\NPC_eff<2>/OUTMUX )
  );
  X_BUF \NPC_eff<2>/OMUX  (
    .I(DLX_IFinst__n0001[2]),
    .O(\NPC_eff<2>/OD )
  );
  X_OPAD \NPC_eff<3>/PAD  (
    .PAD(NPC_eff[3])
  );
  X_TRI NPC_eff_3_OBUF (
    .I(\NPC_eff<3>/OUTMUX ),
    .CTL(\NPC_eff<3>/ENABLE ),
    .O(NPC_eff[3])
  );
  X_INV \NPC_eff<3>/ENABLEINV  (
    .I(\NPC_eff<3>/TORGTS ),
    .O(\NPC_eff<3>/ENABLE )
  );
  X_BUF \NPC_eff<3>/GTS_OR  (
    .I(GTS),
    .O(\NPC_eff<3>/TORGTS )
  );
  X_BUF \NPC_eff<3>/OUTMUX_40  (
    .I(DLX_IFinst_NPC_3_1),
    .O(\NPC_eff<3>/OUTMUX )
  );
  X_BUF \NPC_eff<3>/OMUX  (
    .I(DLX_IFinst__n0001[3]),
    .O(\NPC_eff<3>/OD )
  );
  X_OPAD \NPC_eff<4>/PAD  (
    .PAD(NPC_eff[4])
  );
  X_TRI NPC_eff_4_OBUF (
    .I(\NPC_eff<4>/OUTMUX ),
    .CTL(\NPC_eff<4>/ENABLE ),
    .O(NPC_eff[4])
  );
  X_INV \NPC_eff<4>/ENABLEINV  (
    .I(\NPC_eff<4>/TORGTS ),
    .O(\NPC_eff<4>/ENABLE )
  );
  X_BUF \NPC_eff<4>/GTS_OR  (
    .I(GTS),
    .O(\NPC_eff<4>/TORGTS )
  );
  X_BUF \NPC_eff<4>/OUTMUX_41  (
    .I(DLX_IFinst_NPC_4_1),
    .O(\NPC_eff<4>/OUTMUX )
  );
  X_BUF \NPC_eff<4>/OMUX  (
    .I(DLX_IFinst__n0001[4]),
    .O(\NPC_eff<4>/OD )
  );
  X_OPAD \NPC_eff<5>/PAD  (
    .PAD(NPC_eff[5])
  );
  X_TRI NPC_eff_5_OBUF (
    .I(\NPC_eff<5>/OUTMUX ),
    .CTL(\NPC_eff<5>/ENABLE ),
    .O(NPC_eff[5])
  );
  X_INV \NPC_eff<5>/ENABLEINV  (
    .I(\NPC_eff<5>/TORGTS ),
    .O(\NPC_eff<5>/ENABLE )
  );
  X_BUF \NPC_eff<5>/GTS_OR  (
    .I(GTS),
    .O(\NPC_eff<5>/TORGTS )
  );
  X_BUF \NPC_eff<5>/OUTMUX_42  (
    .I(DLX_IFinst_NPC_5_1),
    .O(\NPC_eff<5>/OUTMUX )
  );
  X_BUF \NPC_eff<5>/OMUX  (
    .I(DLX_IFinst__n0001[5]),
    .O(\NPC_eff<5>/OD )
  );
  X_OPAD \NPC_eff<6>/PAD  (
    .PAD(NPC_eff[6])
  );
  X_TRI NPC_eff_6_OBUF (
    .I(\NPC_eff<6>/OUTMUX ),
    .CTL(\NPC_eff<6>/ENABLE ),
    .O(NPC_eff[6])
  );
  X_INV \NPC_eff<6>/ENABLEINV  (
    .I(\NPC_eff<6>/TORGTS ),
    .O(\NPC_eff<6>/ENABLE )
  );
  X_BUF \NPC_eff<6>/GTS_OR  (
    .I(GTS),
    .O(\NPC_eff<6>/TORGTS )
  );
  X_BUF \NPC_eff<6>/OUTMUX_43  (
    .I(DLX_IFinst_NPC_6_1),
    .O(\NPC_eff<6>/OUTMUX )
  );
  X_BUF \NPC_eff<6>/OMUX  (
    .I(DLX_IFinst__n0001[6]),
    .O(\NPC_eff<6>/OD )
  );
  X_OPAD \NPC_eff<7>/PAD  (
    .PAD(NPC_eff[7])
  );
  X_TRI NPC_eff_7_OBUF (
    .I(\NPC_eff<7>/OUTMUX ),
    .CTL(\NPC_eff<7>/ENABLE ),
    .O(NPC_eff[7])
  );
  X_INV \NPC_eff<7>/ENABLEINV  (
    .I(\NPC_eff<7>/TORGTS ),
    .O(\NPC_eff<7>/ENABLE )
  );
  X_BUF \NPC_eff<7>/GTS_OR  (
    .I(GTS),
    .O(\NPC_eff<7>/TORGTS )
  );
  X_BUF \NPC_eff<7>/OUTMUX_44  (
    .I(DLX_IFinst_NPC_7_1),
    .O(\NPC_eff<7>/OUTMUX )
  );
  X_BUF \NPC_eff<7>/OMUX  (
    .I(DLX_IFinst__n0001[7]),
    .O(\NPC_eff<7>/OD )
  );
  X_OPAD \NPC_eff<8>/PAD  (
    .PAD(NPC_eff[8])
  );
  X_TRI NPC_eff_8_OBUF (
    .I(\NPC_eff<8>/OUTMUX ),
    .CTL(\NPC_eff<8>/ENABLE ),
    .O(NPC_eff[8])
  );
  X_INV \NPC_eff<8>/ENABLEINV  (
    .I(\NPC_eff<8>/TORGTS ),
    .O(\NPC_eff<8>/ENABLE )
  );
  X_BUF \NPC_eff<8>/GTS_OR  (
    .I(GTS),
    .O(\NPC_eff<8>/TORGTS )
  );
  X_BUF \NPC_eff<8>/OUTMUX_45  (
    .I(DLX_IFinst_NPC_8_1),
    .O(\NPC_eff<8>/OUTMUX )
  );
  X_BUF \NPC_eff<8>/OMUX  (
    .I(DLX_IFinst__n0001[8]),
    .O(\NPC_eff<8>/OD )
  );
  X_OPAD \NPC_eff<9>/PAD  (
    .PAD(NPC_eff[9])
  );
  X_TRI NPC_eff_9_OBUF (
    .I(\NPC_eff<9>/OUTMUX ),
    .CTL(\NPC_eff<9>/ENABLE ),
    .O(NPC_eff[9])
  );
  X_INV \NPC_eff<9>/ENABLEINV  (
    .I(\NPC_eff<9>/TORGTS ),
    .O(\NPC_eff<9>/ENABLE )
  );
  X_BUF \NPC_eff<9>/GTS_OR  (
    .I(GTS),
    .O(\NPC_eff<9>/TORGTS )
  );
  X_BUF \NPC_eff<9>/OUTMUX_46  (
    .I(DLX_IFinst_NPC_9_1),
    .O(\NPC_eff<9>/OUTMUX )
  );
  X_BUF \NPC_eff<9>/OMUX  (
    .I(DLX_IFinst__n0001[9]),
    .O(\NPC_eff<9>/OD )
  );
  X_OPAD \stall/PAD  (
    .PAD(stall)
  );
  X_TRI stall_OBUF (
    .I(\stall/OUTMUX ),
    .CTL(\stall/ENABLE ),
    .O(stall)
  );
  X_INV \stall/ENABLEINV  (
    .I(\stall/TORGTS ),
    .O(\stall/ENABLE )
  );
  X_BUF \stall/GTS_OR  (
    .I(GTS),
    .O(\stall/TORGTS )
  );
  X_BUF \stall/OUTMUX_47  (
    .I(DLX_IDinst_stall_1),
    .O(\stall/OUTMUX )
  );
  X_BUF \stall/OMUX  (
    .I(N110648),
    .O(\stall/OD )
  );
  X_OPAD \CLI/PAD  (
    .PAD(CLI)
  );
  X_TRI CLI_OBUF (
    .I(\CLI/OUTMUX ),
    .CTL(\CLI/ENABLE ),
    .O(CLI)
  );
  X_INV \CLI/ENABLEINV  (
    .I(\CLI/TORGTS ),
    .O(\CLI/ENABLE )
  );
  X_BUF \CLI/GTS_OR  (
    .I(GTS),
    .O(\CLI/TORGTS )
  );
  X_BUF \CLI/OUTMUX_48  (
    .I(DLX_IDinst_CLI_1),
    .O(\CLI/OUTMUX )
  );
  X_BUF \CLI/OMUX  (
    .I(DLX_IDinst__n0124),
    .O(\CLI/OD )
  );
  X_IPAD \INT/PAD  (
    .PAD(INT)
  );
  X_BUF \INT/IMUX  (
    .I(\INT/IBUF ),
    .O(INT_IBUF)
  );
  X_BUF INT_IBUF_49 (
    .I(INT),
    .O(\INT/IBUF )
  );
  X_OPAD \DM_addr_eff<0>/PAD  (
    .PAD(DM_addr_eff[0])
  );
  X_TRI DM_addr_eff_0_OBUF (
    .I(\DM_addr_eff<0>/OUTMUX ),
    .CTL(\DM_addr_eff<0>/ENABLE ),
    .O(DM_addr_eff[0])
  );
  X_INV \DM_addr_eff<0>/ENABLEINV  (
    .I(\DM_addr_eff<0>/TORGTS ),
    .O(\DM_addr_eff<0>/ENABLE )
  );
  X_BUF \DM_addr_eff<0>/GTS_OR  (
    .I(GTS),
    .O(\DM_addr_eff<0>/TORGTS )
  );
  X_BUF \DM_addr_eff<0>/OUTMUX_50  (
    .I(DLX_EXinst_ALU_result_0_1),
    .O(\DM_addr_eff<0>/OUTMUX )
  );
  X_BUF \DM_addr_eff<0>/OMUX  (
    .I(N125635),
    .O(\DM_addr_eff<0>/OD )
  );
  X_OPAD \DM_addr_eff<1>/PAD  (
    .PAD(DM_addr_eff[1])
  );
  X_TRI DM_addr_eff_1_OBUF (
    .I(\DM_addr_eff<1>/OUTMUX ),
    .CTL(\DM_addr_eff<1>/ENABLE ),
    .O(DM_addr_eff[1])
  );
  X_INV \DM_addr_eff<1>/ENABLEINV  (
    .I(\DM_addr_eff<1>/TORGTS ),
    .O(\DM_addr_eff<1>/ENABLE )
  );
  X_BUF \DM_addr_eff<1>/GTS_OR  (
    .I(GTS),
    .O(\DM_addr_eff<1>/TORGTS )
  );
  X_BUF \DM_addr_eff<1>/OUTMUX_51  (
    .I(DLX_EXinst_ALU_result_1_1),
    .O(\DM_addr_eff<1>/OUTMUX )
  );
  X_BUF \DM_addr_eff<1>/OMUX  (
    .I(N124056),
    .O(\DM_addr_eff<1>/OD )
  );
  X_OPAD \DM_addr_eff<2>/PAD  (
    .PAD(DM_addr_eff[2])
  );
  X_TRI DM_addr_eff_2_OBUF (
    .I(\DM_addr_eff<2>/OUTMUX ),
    .CTL(\DM_addr_eff<2>/ENABLE ),
    .O(DM_addr_eff[2])
  );
  X_INV \DM_addr_eff<2>/ENABLEINV  (
    .I(\DM_addr_eff<2>/TORGTS ),
    .O(\DM_addr_eff<2>/ENABLE )
  );
  X_BUF \DM_addr_eff<2>/GTS_OR  (
    .I(GTS),
    .O(\DM_addr_eff<2>/TORGTS )
  );
  X_BUF \DM_addr_eff<2>/OUTMUX_52  (
    .I(DLX_EXinst_ALU_result_2_1),
    .O(\DM_addr_eff<2>/OUTMUX )
  );
  X_BUF \DM_addr_eff<2>/OMUX  (
    .I(N123038),
    .O(\DM_addr_eff<2>/OD )
  );
  X_OPAD \DM_addr_eff<3>/PAD  (
    .PAD(DM_addr_eff[3])
  );
  X_TRI DM_addr_eff_3_OBUF (
    .I(\DM_addr_eff<3>/OUTMUX ),
    .CTL(\DM_addr_eff<3>/ENABLE ),
    .O(DM_addr_eff[3])
  );
  X_INV \DM_addr_eff<3>/ENABLEINV  (
    .I(\DM_addr_eff<3>/TORGTS ),
    .O(\DM_addr_eff<3>/ENABLE )
  );
  X_BUF \DM_addr_eff<3>/GTS_OR  (
    .I(GTS),
    .O(\DM_addr_eff<3>/TORGTS )
  );
  X_BUF \DM_addr_eff<3>/OUTMUX_53  (
    .I(DLX_EXinst_ALU_result_3_1),
    .O(\DM_addr_eff<3>/OUTMUX )
  );
  X_BUF \DM_addr_eff<3>/OMUX  (
    .I(N120114),
    .O(\DM_addr_eff<3>/OD )
  );
  X_OPAD \DM_addr_eff<4>/PAD  (
    .PAD(DM_addr_eff[4])
  );
  X_TRI DM_addr_eff_4_OBUF (
    .I(\DM_addr_eff<4>/OUTMUX ),
    .CTL(\DM_addr_eff<4>/ENABLE ),
    .O(DM_addr_eff[4])
  );
  X_INV \DM_addr_eff<4>/ENABLEINV  (
    .I(\DM_addr_eff<4>/TORGTS ),
    .O(\DM_addr_eff<4>/ENABLE )
  );
  X_BUF \DM_addr_eff<4>/GTS_OR  (
    .I(GTS),
    .O(\DM_addr_eff<4>/TORGTS )
  );
  X_BUF \DM_addr_eff<4>/OUTMUX_54  (
    .I(DLX_EXinst_ALU_result_4_1),
    .O(\DM_addr_eff<4>/OUTMUX )
  );
  X_BUF \DM_addr_eff<4>/OMUX  (
    .I(N113660),
    .O(\DM_addr_eff<4>/OD )
  );
  defparam DLX_EXinst_ALU_result_14_1_55.INIT = 1'b0;
  X_FF DLX_EXinst_ALU_result_14_1_55 (
    .I(\DM_addr_eff<14>/OD ),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DM_addr_eff<14>/OFF/RST ),
    .O(DLX_EXinst_ALU_result_14_1)
  );
  X_OR2 \DM_addr_eff<14>/OFF/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DM_addr_eff<14>/OFF/RST )
  );
  X_OPAD \DM_addr_eff<5>/PAD  (
    .PAD(DM_addr_eff[5])
  );
  X_TRI DM_addr_eff_5_OBUF (
    .I(\DM_addr_eff<5>/OUTMUX ),
    .CTL(\DM_addr_eff<5>/ENABLE ),
    .O(DM_addr_eff[5])
  );
  X_INV \DM_addr_eff<5>/ENABLEINV  (
    .I(\DM_addr_eff<5>/TORGTS ),
    .O(\DM_addr_eff<5>/ENABLE )
  );
  X_BUF \DM_addr_eff<5>/GTS_OR  (
    .I(GTS),
    .O(\DM_addr_eff<5>/TORGTS )
  );
  X_BUF \DM_addr_eff<5>/OUTMUX_56  (
    .I(DLX_EXinst_ALU_result_5_1),
    .O(\DM_addr_eff<5>/OUTMUX )
  );
  X_BUF \DM_addr_eff<5>/OMUX  (
    .I(N116396),
    .O(\DM_addr_eff<5>/OD )
  );
  X_OPAD \DM_addr_eff<6>/PAD  (
    .PAD(DM_addr_eff[6])
  );
  X_TRI DM_addr_eff_6_OBUF (
    .I(\DM_addr_eff<6>/OUTMUX ),
    .CTL(\DM_addr_eff<6>/ENABLE ),
    .O(DM_addr_eff[6])
  );
  X_INV \DM_addr_eff<6>/ENABLEINV  (
    .I(\DM_addr_eff<6>/TORGTS ),
    .O(\DM_addr_eff<6>/ENABLE )
  );
  X_BUF \DM_addr_eff<6>/GTS_OR  (
    .I(GTS),
    .O(\DM_addr_eff<6>/TORGTS )
  );
  X_BUF \DM_addr_eff<6>/OUTMUX_57  (
    .I(DLX_EXinst_ALU_result_6_1),
    .O(\DM_addr_eff<6>/OUTMUX )
  );
  X_BUF \DM_addr_eff<6>/OMUX  (
    .I(N115984),
    .O(\DM_addr_eff<6>/OD )
  );
  X_OPAD \DM_addr_eff<7>/PAD  (
    .PAD(DM_addr_eff[7])
  );
  X_TRI DM_addr_eff_7_OBUF (
    .I(\DM_addr_eff<7>/OUTMUX ),
    .CTL(\DM_addr_eff<7>/ENABLE ),
    .O(DM_addr_eff[7])
  );
  X_INV \DM_addr_eff<7>/ENABLEINV  (
    .I(\DM_addr_eff<7>/TORGTS ),
    .O(\DM_addr_eff<7>/ENABLE )
  );
  X_BUF \DM_addr_eff<7>/GTS_OR  (
    .I(GTS),
    .O(\DM_addr_eff<7>/TORGTS )
  );
  X_BUF \DM_addr_eff<7>/OUTMUX_58  (
    .I(DLX_EXinst_ALU_result_7_1),
    .O(\DM_addr_eff<7>/OUTMUX )
  );
  X_BUF \DM_addr_eff<7>/OMUX  (
    .I(N112616),
    .O(\DM_addr_eff<7>/OD )
  );
  X_OPAD \DM_addr_eff<8>/PAD  (
    .PAD(DM_addr_eff[8])
  );
  X_TRI DM_addr_eff_8_OBUF (
    .I(\DM_addr_eff<8>/OUTMUX ),
    .CTL(\DM_addr_eff<8>/ENABLE ),
    .O(DM_addr_eff[8])
  );
  X_INV \DM_addr_eff<8>/ENABLEINV  (
    .I(\DM_addr_eff<8>/TORGTS ),
    .O(\DM_addr_eff<8>/ENABLE )
  );
  X_BUF \DM_addr_eff<8>/GTS_OR  (
    .I(GTS),
    .O(\DM_addr_eff<8>/TORGTS )
  );
  X_BUF \DM_addr_eff<8>/OUTMUX_59  (
    .I(DLX_EXinst_ALU_result_8_1),
    .O(\DM_addr_eff<8>/OUTMUX )
  );
  X_BUF \DM_addr_eff<8>/OMUX  (
    .I(N111878),
    .O(\DM_addr_eff<8>/OD )
  );
  X_OPAD \DM_addr_eff<9>/PAD  (
    .PAD(DM_addr_eff[9])
  );
  X_TRI DM_addr_eff_9_OBUF (
    .I(\DM_addr_eff<9>/OUTMUX ),
    .CTL(\DM_addr_eff<9>/ENABLE ),
    .O(DM_addr_eff[9])
  );
  X_INV \DM_addr_eff<9>/ENABLEINV  (
    .I(\DM_addr_eff<9>/TORGTS ),
    .O(\DM_addr_eff<9>/ENABLE )
  );
  X_BUF \DM_addr_eff<9>/GTS_OR  (
    .I(GTS),
    .O(\DM_addr_eff<9>/TORGTS )
  );
  X_BUF \DM_addr_eff<9>/OUTMUX_60  (
    .I(DLX_EXinst_ALU_result_9_1),
    .O(\DM_addr_eff<9>/OUTMUX )
  );
  X_BUF \DM_addr_eff<9>/OMUX  (
    .I(N117154),
    .O(\DM_addr_eff<9>/OD )
  );
  X_ZERO \vsync/LOGIC_ZERO_61  (
    .O(\vsync/LOGIC_ZERO )
  );
  X_OPAD \vsync/PAD  (
    .PAD(vsync)
  );
  X_TRI vsync_OBUF (
    .I(\vsync/OUTMUX ),
    .CTL(\vsync/ENABLE ),
    .O(vsync)
  );
  X_INV \vsync/ENABLEINV  (
    .I(\vsync/TORGTS ),
    .O(\vsync/ENABLE )
  );
  X_BUF \vsync/GTS_OR  (
    .I(GTS),
    .O(\vsync/TORGTS )
  );
  X_BUF \vsync/OUTMUX_62  (
    .I(vga_top_vga1_vsyncout),
    .O(\vsync/OUTMUX )
  );
  X_IPAD \FREEZE/PAD  (
    .PAD(FREEZE)
  );
  X_BUF \FREEZE/IMUX  (
    .I(\FREEZE/IBUF ),
    .O(FREEZE_IBUF)
  );
  X_BUF FREEZE_IBUF_63 (
    .I(FREEZE),
    .O(\FREEZE/IBUF )
  );
  X_OPAD \IR_MSB<0>/PAD  (
    .PAD(IR_MSB[0])
  );
  X_TRI IR_MSB_0_OBUF_64 (
    .I(\IR_MSB<0>/OUTMUX ),
    .CTL(\IR_MSB<0>/ENABLE ),
    .O(IR_MSB[0])
  );
  X_INV \IR_MSB<0>/ENABLEINV  (
    .I(\IR_MSB<0>/TORGTS ),
    .O(\IR_MSB<0>/ENABLE )
  );
  X_BUF \IR_MSB<0>/GTS_OR  (
    .I(GTS),
    .O(\IR_MSB<0>/TORGTS )
  );
  X_BUF \IR_MSB<0>/OUTMUX_65  (
    .I(IR_MSB_0_OBUF),
    .O(\IR_MSB<0>/OUTMUX )
  );
  X_OPAD \IR_MSB<1>/PAD  (
    .PAD(IR_MSB[1])
  );
  X_TRI IR_MSB_1_OBUF_66 (
    .I(\IR_MSB<1>/OUTMUX ),
    .CTL(\IR_MSB<1>/ENABLE ),
    .O(IR_MSB[1])
  );
  X_INV \IR_MSB<1>/ENABLEINV  (
    .I(\IR_MSB<1>/TORGTS ),
    .O(\IR_MSB<1>/ENABLE )
  );
  X_BUF \IR_MSB<1>/GTS_OR  (
    .I(GTS),
    .O(\IR_MSB<1>/TORGTS )
  );
  X_BUF \IR_MSB<1>/OUTMUX_67  (
    .I(IR_MSB_1_OBUF),
    .O(\IR_MSB<1>/OUTMUX )
  );
  X_OPAD \IR_MSB<2>/PAD  (
    .PAD(IR_MSB[2])
  );
  X_TRI IR_MSB_2_OBUF_68 (
    .I(\IR_MSB<2>/OUTMUX ),
    .CTL(\IR_MSB<2>/ENABLE ),
    .O(IR_MSB[2])
  );
  X_INV \IR_MSB<2>/ENABLEINV  (
    .I(\IR_MSB<2>/TORGTS ),
    .O(\IR_MSB<2>/ENABLE )
  );
  X_BUF \IR_MSB<2>/GTS_OR  (
    .I(GTS),
    .O(\IR_MSB<2>/TORGTS )
  );
  X_BUF \IR_MSB<2>/OUTMUX_69  (
    .I(IR_MSB_2_OBUF),
    .O(\IR_MSB<2>/OUTMUX )
  );
  X_OPAD \IR_MSB<3>/PAD  (
    .PAD(IR_MSB[3])
  );
  X_TRI IR_MSB_3_OBUF_70 (
    .I(\IR_MSB<3>/OUTMUX ),
    .CTL(\IR_MSB<3>/ENABLE ),
    .O(IR_MSB[3])
  );
  X_INV \IR_MSB<3>/ENABLEINV  (
    .I(\IR_MSB<3>/TORGTS ),
    .O(\IR_MSB<3>/ENABLE )
  );
  X_BUF \IR_MSB<3>/GTS_OR  (
    .I(GTS),
    .O(\IR_MSB<3>/TORGTS )
  );
  X_BUF \IR_MSB<3>/OUTMUX_71  (
    .I(IR_MSB_3_OBUF),
    .O(\IR_MSB<3>/OUTMUX )
  );
  X_OPAD \IR_MSB<4>/PAD  (
    .PAD(IR_MSB[4])
  );
  X_TRI IR_MSB_4_OBUF_72 (
    .I(\IR_MSB<4>/OUTMUX ),
    .CTL(\IR_MSB<4>/ENABLE ),
    .O(IR_MSB[4])
  );
  X_INV \IR_MSB<4>/ENABLEINV  (
    .I(\IR_MSB<4>/TORGTS ),
    .O(\IR_MSB<4>/ENABLE )
  );
  X_BUF \IR_MSB<4>/GTS_OR  (
    .I(GTS),
    .O(\IR_MSB<4>/TORGTS )
  );
  X_BUF \IR_MSB<4>/OUTMUX_73  (
    .I(IR_MSB_4_OBUF),
    .O(\IR_MSB<4>/OUTMUX )
  );
  X_OPAD \IR_MSB<5>/PAD  (
    .PAD(IR_MSB[5])
  );
  X_TRI IR_MSB_5_OBUF_74 (
    .I(\IR_MSB<5>/OUTMUX ),
    .CTL(\IR_MSB<5>/ENABLE ),
    .O(IR_MSB[5])
  );
  X_INV \IR_MSB<5>/ENABLEINV  (
    .I(\IR_MSB<5>/TORGTS ),
    .O(\IR_MSB<5>/ENABLE )
  );
  X_BUF \IR_MSB<5>/GTS_OR  (
    .I(GTS),
    .O(\IR_MSB<5>/TORGTS )
  );
  X_BUF \IR_MSB<5>/OUTMUX_75  (
    .I(IR_MSB_5_OBUF),
    .O(\IR_MSB<5>/OUTMUX )
  );
  X_OPAD \IR_MSB<6>/PAD  (
    .PAD(IR_MSB[6])
  );
  X_TRI IR_MSB_6_OBUF_76 (
    .I(\IR_MSB<6>/OUTMUX ),
    .CTL(\IR_MSB<6>/ENABLE ),
    .O(IR_MSB[6])
  );
  X_INV \IR_MSB<6>/ENABLEINV  (
    .I(\IR_MSB<6>/TORGTS ),
    .O(\IR_MSB<6>/ENABLE )
  );
  X_BUF \IR_MSB<6>/GTS_OR  (
    .I(GTS),
    .O(\IR_MSB<6>/TORGTS )
  );
  X_BUF \IR_MSB<6>/OUTMUX_77  (
    .I(IR_MSB_6_OBUF),
    .O(\IR_MSB<6>/OUTMUX )
  );
  X_OPAD \IR_MSB<7>/PAD  (
    .PAD(IR_MSB[7])
  );
  X_TRI IR_MSB_7_OBUF_78 (
    .I(\IR_MSB<7>/OUTMUX ),
    .CTL(\IR_MSB<7>/ENABLE ),
    .O(IR_MSB[7])
  );
  X_INV \IR_MSB<7>/ENABLEINV  (
    .I(\IR_MSB<7>/TORGTS ),
    .O(\IR_MSB<7>/ENABLE )
  );
  X_BUF \IR_MSB<7>/GTS_OR  (
    .I(GTS),
    .O(\IR_MSB<7>/TORGTS )
  );
  X_BUF \IR_MSB<7>/OUTMUX_79  (
    .I(IR_MSB_7_OBUF),
    .O(\IR_MSB<7>/OUTMUX )
  );
  X_IPAD \delay_selectDM<0>/PAD  (
    .PAD(delay_selectDM[0])
  );
  X_BUF \delay_selectDM<0>/IMUX  (
    .I(\delay_selectDM<0>/IBUF ),
    .O(delay_selectDM_0_IBUF)
  );
  X_BUF delay_selectDM_0_IBUF_80 (
    .I(delay_selectDM[0]),
    .O(\delay_selectDM<0>/IBUF )
  );
  X_IPAD \delay_selectDM<1>/PAD  (
    .PAD(delay_selectDM[1])
  );
  X_BUF \delay_selectDM<1>/IMUX  (
    .I(\delay_selectDM<1>/IBUF ),
    .O(delay_selectDM_1_IBUF)
  );
  X_BUF delay_selectDM_1_IBUF_81 (
    .I(delay_selectDM[1]),
    .O(\delay_selectDM<1>/IBUF )
  );
  defparam DLX_IDinst_branch_sig_1_82.INIT = 1'b0;
  X_FF DLX_IDinst_branch_sig_1_82 (
    .I(\branch_sig/OD ),
    .CE(DLX_IDinst__n0422),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\branch_sig/OFF/RST ),
    .O(DLX_IDinst_branch_sig_1)
  );
  X_OR2 \branch_sig/OFF/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\branch_sig/OFF/RST )
  );
  X_IPAD \delay_selectID<0>/PAD  (
    .PAD(delay_selectID[0])
  );
  X_BUF \delay_selectID<0>/IMUX  (
    .I(\delay_selectID<0>/IBUF ),
    .O(delay_selectID_0_IBUF)
  );
  X_BUF delay_selectID_0_IBUF_83 (
    .I(delay_selectID[0]),
    .O(\delay_selectID<0>/IBUF )
  );
  X_IPAD \delay_selectID<1>/PAD  (
    .PAD(delay_selectID[1])
  );
  X_BUF \delay_selectID<1>/IMUX  (
    .I(\delay_selectID<1>/IBUF ),
    .O(delay_selectID_1_IBUF)
  );
  X_BUF delay_selectID_1_IBUF_84 (
    .I(delay_selectID[1]),
    .O(\delay_selectID<1>/IBUF )
  );
  X_OPAD \clk_MEM/PAD  (
    .PAD(clk_MEM)
  );
  X_TRI clk_MEM_OBUF (
    .I(\clk_MEM/OUTMUX ),
    .CTL(\clk_MEM/ENABLE ),
    .O(clk_MEM)
  );
  X_INV \clk_MEM/ENABLEINV  (
    .I(\clk_MEM/TORGTS ),
    .O(\clk_MEM/ENABLE )
  );
  X_BUF \clk_MEM/GTS_OR  (
    .I(GTS),
    .O(\clk_MEM/TORGTS )
  );
  X_BUF \clk_MEM/OUTMUX_85  (
    .I(\clk_MEM/ODNOT ),
    .O(\clk_MEM/OUTMUX )
  );
  X_INV \clk_MEM/OMUX  (
    .I(DLX_MEMlc_master_ctrlMEM_l),
    .O(\clk_MEM/ODNOT )
  );
  X_IPAD \delay_selectIF<0>/PAD  (
    .PAD(delay_selectIF[0])
  );
  X_BUF \delay_selectIF<0>/IMUX  (
    .I(\delay_selectIF<0>/IBUF ),
    .O(delay_selectIF_0_IBUF)
  );
  X_BUF delay_selectIF_0_IBUF_86 (
    .I(delay_selectIF[0]),
    .O(\delay_selectIF<0>/IBUF )
  );
  X_IPAD \delay_selectIF<1>/PAD  (
    .PAD(delay_selectIF[1])
  );
  X_BUF \delay_selectIF<1>/IMUX  (
    .I(\delay_selectIF<1>/IBUF ),
    .O(delay_selectIF_1_IBUF)
  );
  X_BUF delay_selectIF_1_IBUF_87 (
    .I(delay_selectIF[1]),
    .O(\delay_selectIF<1>/IBUF )
  );
  X_IPAD \delay_selectMEM<0>/PAD  (
    .PAD(delay_selectMEM[0])
  );
  X_BUF \delay_selectMEM<0>/IMUX  (
    .I(\delay_selectMEM<0>/IBUF ),
    .O(delay_selectMEM_0_IBUF)
  );
  X_BUF delay_selectMEM_0_IBUF_88 (
    .I(delay_selectMEM[0]),
    .O(\delay_selectMEM<0>/IBUF )
  );
  X_IPAD \delay_selectMEM<1>/PAD  (
    .PAD(delay_selectMEM[1])
  );
  X_BUF \delay_selectMEM<1>/IMUX  (
    .I(\delay_selectMEM<1>/IBUF ),
    .O(delay_selectMEM_1_IBUF)
  );
  X_BUF delay_selectMEM_1_IBUF_89 (
    .I(delay_selectMEM[1]),
    .O(\delay_selectMEM<1>/IBUF )
  );
  X_OPAD \blue<0>/PAD  (
    .PAD(blue[0])
  );
  X_TRI blue_0_OBUF_90 (
    .I(\blue<0>/OUTMUX ),
    .CTL(\blue<0>/ENABLE ),
    .O(blue[0])
  );
  X_INV \blue<0>/ENABLEINV  (
    .I(\blue<0>/TORGTS ),
    .O(\blue<0>/ENABLE )
  );
  X_BUF \blue<0>/GTS_OR  (
    .I(GTS),
    .O(\blue<0>/TORGTS )
  );
  X_BUF \blue<0>/OUTMUX_91  (
    .I(blue_0_OBUF),
    .O(\blue<0>/OUTMUX )
  );
  X_OPAD \blue<1>/PAD  (
    .PAD(blue[1])
  );
  X_TRI blue_1_OBUF_92 (
    .I(\blue<1>/OUTMUX ),
    .CTL(\blue<1>/ENABLE ),
    .O(blue[1])
  );
  X_INV \blue<1>/ENABLEINV  (
    .I(\blue<1>/TORGTS ),
    .O(\blue<1>/ENABLE )
  );
  X_BUF \blue<1>/GTS_OR  (
    .I(GTS),
    .O(\blue<1>/TORGTS )
  );
  X_BUF \blue<1>/OUTMUX_93  (
    .I(blue_1_OBUF),
    .O(\blue<1>/OUTMUX )
  );
  X_OPAD \blue<2>/PAD  (
    .PAD(blue[2])
  );
  X_TRI blue_2_OBUF_94 (
    .I(\blue<2>/OUTMUX ),
    .CTL(\blue<2>/ENABLE ),
    .O(blue[2])
  );
  X_INV \blue<2>/ENABLEINV  (
    .I(\blue<2>/TORGTS ),
    .O(\blue<2>/ENABLE )
  );
  X_BUF \blue<2>/GTS_OR  (
    .I(GTS),
    .O(\blue<2>/TORGTS )
  );
  X_BUF \blue<2>/OUTMUX_95  (
    .I(blue_2_OBUF),
    .O(\blue<2>/OUTMUX )
  );
  X_IPAD \STOP_fetch/PAD  (
    .PAD(STOP_fetch)
  );
  X_BUF \STOP_fetch/IMUX  (
    .I(\STOP_fetch/IBUF ),
    .O(STOP_fetch_IBUF)
  );
  X_BUF STOP_fetch_IBUF_96 (
    .I(STOP_fetch),
    .O(\STOP_fetch/IBUF )
  );
  X_IPAD \delay_selectEX<0>/PAD  (
    .PAD(delay_selectEX[0])
  );
  X_BUF \delay_selectEX<0>/IMUX  (
    .I(\delay_selectEX<0>/IBUF ),
    .O(delay_selectEX_0_IBUF)
  );
  X_BUF delay_selectEX_0_IBUF_97 (
    .I(delay_selectEX[0]),
    .O(\delay_selectEX<0>/IBUF )
  );
  X_IPAD \delay_selectEX<1>/PAD  (
    .PAD(delay_selectEX[1])
  );
  X_BUF \delay_selectEX<1>/IMUX  (
    .I(\delay_selectEX<1>/IBUF ),
    .O(delay_selectEX_1_IBUF)
  );
  X_BUF delay_selectEX_1_IBUF_98 (
    .I(delay_selectEX[1]),
    .O(\delay_selectEX<1>/IBUF )
  );
  X_OPAD \mask<0>/PAD  (
    .PAD(mask[0])
  );
  X_TRI mask_0_OBUF_99 (
    .I(\mask<0>/OUTMUX ),
    .CTL(\mask<0>/ENABLE ),
    .O(mask[0])
  );
  X_INV \mask<0>/ENABLEINV  (
    .I(\mask<0>/TORGTS ),
    .O(\mask<0>/ENABLE )
  );
  X_BUF \mask<0>/GTS_OR  (
    .I(GTS),
    .O(\mask<0>/TORGTS )
  );
  X_BUF \mask<0>/OUTMUX_100  (
    .I(mask_0_OBUF),
    .O(\mask<0>/OUTMUX )
  );
  X_IPAD \delay_selectRF<0>/PAD  (
    .PAD(delay_selectRF[0])
  );
  X_BUF \delay_selectRF<0>/IMUX  (
    .I(\delay_selectRF<0>/IBUF ),
    .O(delay_selectRF_0_IBUF)
  );
  X_BUF delay_selectRF_0_IBUF_101 (
    .I(delay_selectRF[0]),
    .O(\delay_selectRF<0>/IBUF )
  );
  X_IPAD \delay_selectRF<1>/PAD  (
    .PAD(delay_selectRF[1])
  );
  X_BUF \delay_selectRF<1>/IMUX  (
    .I(\delay_selectRF<1>/IBUF ),
    .O(delay_selectRF_1_IBUF)
  );
  X_BUF delay_selectRF_1_IBUF_102 (
    .I(delay_selectRF[1]),
    .O(\delay_selectRF<1>/IBUF )
  );
  X_OPAD \DM_read/PAD  (
    .PAD(DM_read)
  );
  X_TRI DM_read_OBUF (
    .I(\DM_read/OUTMUX ),
    .CTL(\DM_read/ENABLE ),
    .O(DM_read)
  );
  X_INV \DM_read/ENABLEINV  (
    .I(\DM_read/TORGTS ),
    .O(\DM_read/ENABLE )
  );
  X_BUF \DM_read/GTS_OR  (
    .I(GTS),
    .O(\DM_read/TORGTS )
  );
  X_BUF \DM_read/OUTMUX_103  (
    .I(DLX_EXinst_mem_read_EX_1),
    .O(\DM_read/OUTMUX )
  );
  X_BUF \DM_read/OMUX  (
    .I(DLX_EXinst__n0011),
    .O(\DM_read/OD )
  );
  X_OPAD \mask<3>/PAD  (
    .PAD(mask[3])
  );
  X_TRI mask_3_OBUF_104 (
    .I(\mask<3>/OUTMUX ),
    .CTL(\mask<3>/ENABLE ),
    .O(mask[3])
  );
  X_INV \mask<3>/ENABLEINV  (
    .I(\mask<3>/TORGTS ),
    .O(\mask<3>/ENABLE )
  );
  X_BUF \mask<3>/GTS_OR  (
    .I(GTS),
    .O(\mask<3>/TORGTS )
  );
  X_BUF \mask<3>/OUTMUX_105  (
    .I(mask_3_OBUF),
    .O(\mask<3>/OUTMUX )
  );
  X_OPAD \NPC_eff<10>/PAD  (
    .PAD(NPC_eff[10])
  );
  X_TRI NPC_eff_10_OBUF (
    .I(\NPC_eff<10>/OUTMUX ),
    .CTL(\NPC_eff<10>/ENABLE ),
    .O(NPC_eff[10])
  );
  X_INV \NPC_eff<10>/ENABLEINV  (
    .I(\NPC_eff<10>/TORGTS ),
    .O(\NPC_eff<10>/ENABLE )
  );
  X_BUF \NPC_eff<10>/GTS_OR  (
    .I(GTS),
    .O(\NPC_eff<10>/TORGTS )
  );
  X_BUF \NPC_eff<10>/OUTMUX_106  (
    .I(DLX_IFinst_NPC_10_1),
    .O(\NPC_eff<10>/OUTMUX )
  );
  X_BUF \NPC_eff<10>/OMUX  (
    .I(DLX_IFinst__n0001[10]),
    .O(\NPC_eff<10>/OD )
  );
  X_OPAD \NPC_eff<11>/PAD  (
    .PAD(NPC_eff[11])
  );
  X_TRI NPC_eff_11_OBUF (
    .I(\NPC_eff<11>/OUTMUX ),
    .CTL(\NPC_eff<11>/ENABLE ),
    .O(NPC_eff[11])
  );
  X_INV \NPC_eff<11>/ENABLEINV  (
    .I(\NPC_eff<11>/TORGTS ),
    .O(\NPC_eff<11>/ENABLE )
  );
  X_BUF \NPC_eff<11>/GTS_OR  (
    .I(GTS),
    .O(\NPC_eff<11>/TORGTS )
  );
  X_BUF \NPC_eff<11>/OUTMUX_107  (
    .I(DLX_IFinst_NPC_11_1),
    .O(\NPC_eff<11>/OUTMUX )
  );
  X_BUF \NPC_eff<11>/OMUX  (
    .I(DLX_IFinst__n0001[11]),
    .O(\NPC_eff<11>/OD )
  );
  X_OPAD \NPC_eff<12>/PAD  (
    .PAD(NPC_eff[12])
  );
  X_TRI NPC_eff_12_OBUF (
    .I(\NPC_eff<12>/OUTMUX ),
    .CTL(\NPC_eff<12>/ENABLE ),
    .O(NPC_eff[12])
  );
  X_INV \NPC_eff<12>/ENABLEINV  (
    .I(\NPC_eff<12>/TORGTS ),
    .O(\NPC_eff<12>/ENABLE )
  );
  X_BUF \NPC_eff<12>/GTS_OR  (
    .I(GTS),
    .O(\NPC_eff<12>/TORGTS )
  );
  X_BUF \NPC_eff<12>/OUTMUX_108  (
    .I(DLX_IFinst_NPC_12_1),
    .O(\NPC_eff<12>/OUTMUX )
  );
  X_BUF \NPC_eff<12>/OMUX  (
    .I(DLX_IFinst__n0001[12]),
    .O(\NPC_eff<12>/OD )
  );
  X_OPAD \NPC_eff<13>/PAD  (
    .PAD(NPC_eff[13])
  );
  X_TRI NPC_eff_13_OBUF (
    .I(\NPC_eff<13>/OUTMUX ),
    .CTL(\NPC_eff<13>/ENABLE ),
    .O(NPC_eff[13])
  );
  X_INV \NPC_eff<13>/ENABLEINV  (
    .I(\NPC_eff<13>/TORGTS ),
    .O(\NPC_eff<13>/ENABLE )
  );
  X_BUF \NPC_eff<13>/GTS_OR  (
    .I(GTS),
    .O(\NPC_eff<13>/TORGTS )
  );
  X_BUF \NPC_eff<13>/OUTMUX_109  (
    .I(DLX_IFinst_NPC_13_1),
    .O(\NPC_eff<13>/OUTMUX )
  );
  X_BUF \NPC_eff<13>/OMUX  (
    .I(DLX_IFinst__n0001[13]),
    .O(\NPC_eff<13>/OD )
  );
  X_OPAD \NPC_eff<14>/PAD  (
    .PAD(NPC_eff[14])
  );
  X_TRI NPC_eff_14_OBUF (
    .I(\NPC_eff<14>/OUTMUX ),
    .CTL(\NPC_eff<14>/ENABLE ),
    .O(NPC_eff[14])
  );
  X_INV \NPC_eff<14>/ENABLEINV  (
    .I(\NPC_eff<14>/TORGTS ),
    .O(\NPC_eff<14>/ENABLE )
  );
  X_BUF \NPC_eff<14>/GTS_OR  (
    .I(GTS),
    .O(\NPC_eff<14>/TORGTS )
  );
  X_BUF \NPC_eff<14>/OUTMUX_110  (
    .I(DLX_IFinst_NPC_14_1),
    .O(\NPC_eff<14>/OUTMUX )
  );
  X_BUF \NPC_eff<14>/OMUX  (
    .I(DLX_IFinst__n0001[14]),
    .O(\NPC_eff<14>/OD )
  );
  X_OPAD \NPC_eff<15>/PAD  (
    .PAD(NPC_eff[15])
  );
  X_TRI NPC_eff_15_OBUF (
    .I(\NPC_eff<15>/OUTMUX ),
    .CTL(\NPC_eff<15>/ENABLE ),
    .O(NPC_eff[15])
  );
  X_INV \NPC_eff<15>/ENABLEINV  (
    .I(\NPC_eff<15>/TORGTS ),
    .O(\NPC_eff<15>/ENABLE )
  );
  X_BUF \NPC_eff<15>/GTS_OR  (
    .I(GTS),
    .O(\NPC_eff<15>/TORGTS )
  );
  X_BUF \NPC_eff<15>/OUTMUX_111  (
    .I(DLX_IFinst_NPC_15_1),
    .O(\NPC_eff<15>/OUTMUX )
  );
  X_BUF \NPC_eff<15>/OMUX  (
    .I(DLX_IFinst__n0001[15]),
    .O(\NPC_eff<15>/OD )
  );
  X_OPAD \DM_write_data<0>/PAD  (
    .PAD(DM_write_data[0])
  );
  X_TRI DM_write_data_0_OBUF (
    .I(\DM_write_data<0>/OUTMUX ),
    .CTL(\DM_write_data<0>/ENABLE ),
    .O(DM_write_data[0])
  );
  X_INV \DM_write_data<0>/ENABLEINV  (
    .I(\DM_write_data<0>/TORGTS ),
    .O(\DM_write_data<0>/ENABLE )
  );
  X_BUF \DM_write_data<0>/GTS_OR  (
    .I(GTS),
    .O(\DM_write_data<0>/TORGTS )
  );
  X_BUF \DM_write_data<0>/OUTMUX_112  (
    .I(DLX_EXinst_reg_out_B_EX_0_1),
    .O(\DM_write_data<0>/OUTMUX )
  );
  X_BUF \DM_write_data<0>/OMUX  (
    .I(DLX_EXinst__n0007[0]),
    .O(\DM_write_data<0>/OD )
  );
  X_ZERO \clkdivider/LOGIC_ZERO_113  (
    .O(\clkdivider/LOGIC_ZERO )
  );
  defparam clkdivider.CLKDV_DIVIDE = 2.0;
  defparam clkdivider.DUTY_CYCLE_CORRECTION = "TRUE";
  defparam clkdivider.MAXPERCLKIN = 40000;
  X_CLKDLLE clkdivider (
    .CLKIN(clkbuf),
    .CLKFB(clk0buf),
    .RST(\clkdivider/LOGIC_ZERO ),
    .CLK0(clk0),
    .CLK90(\clkdivider/CLK90 ),
    .CLK180(\clkdivider/CLK180 ),
    .CLK270(\clkdivider/CLK270 ),
    .CLK2X(\clkdivider/CLK2X ),
    .CLK2X180(\clkdivider/CLK2X180 ),
    .CLKDV(clkdivub),
    .LOCKED(\clkdivider/LOCKED )
  );
  X_ZERO \DLX_IDinst_RF_block0s0/LOGIC_ZERO_114  (
    .O(\DLX_IDinst_RF_block0s0/LOGIC_ZERO )
  );
  defparam DLX_IDinst_RF_block0s0.INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block0s0.INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block0s0.INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block0s0.INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block0s0.INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block0s0.INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block0s0.INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block0s0.INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block0s0.INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block0s0.INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block0s0.INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block0s0.INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block0s0.INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block0s0.INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block0s0.INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block0s0.INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block0s0.SETUP_ALL = 2701;
  X_RAMB4_S16_S16 DLX_IDinst_RF_block0s0 (
    .CLKA(DLX_clk_IF_del),
    .CLKB(DLX_clk_ID),
    .ENA(DLX_IDinst__n0000),
    .ENB(DLX_IDinst__n0410),
    .RSTA(DLX_IDinst__n0002),
    .RSTB(\DLX_IDinst_RF_block0s0/LOGIC_ZERO ),
    .WEA(\DLX_IDinst_RF_block0s0/LOGIC_ZERO ),
    .WEB(DLX_MEMinst_reg_write_MEM),
    .GSR(GSR),
    .ADDRA({GLOBAL_LOGIC0, GLOBAL_LOGIC0_2, GLOBAL_LOGIC0_1, DLX_IDinst_regA_index[4], DLX_IDinst_regA_index[3], DLX_IDinst_regA_index[2], 
DLX_IDinst_regA_index[1], DLX_IDinst_regA_index[0]}),
    .ADDRB({GLOBAL_LOGIC0_1, GLOBAL_LOGIC0_2, GLOBAL_LOGIC0_1, DLX_MEMinst_reg_dst_out[4], DLX_MEMinst_reg_dst_out[3], DLX_MEMinst_reg_dst_out[2], 
DLX_MEMinst_reg_dst_out[1], DLX_MEMinst_reg_dst_out[0]}),
    .DIA({\DLX_IDinst_RF_block0s0/DIA15 , \DLX_IDinst_RF_block0s0/DIA14 , \DLX_IDinst_RF_block0s0/DIA13 , \DLX_IDinst_RF_block0s0/DIA12 , 
\DLX_IDinst_RF_block0s0/DIA11 , \DLX_IDinst_RF_block0s0/DIA10 , \DLX_IDinst_RF_block0s0/DIA9 , \DLX_IDinst_RF_block0s0/DIA8 , 
\DLX_IDinst_RF_block0s0/DIA7 , \DLX_IDinst_RF_block0s0/DIA6 , \DLX_IDinst_RF_block0s0/DIA5 , \DLX_IDinst_RF_block0s0/DIA4 , 
\DLX_IDinst_RF_block0s0/DIA3 , \DLX_IDinst_RF_block0s0/DIA2 , \DLX_IDinst_RF_block0s0/DIA1 , \DLX_IDinst_RF_block0s0/DIA0 }),
    .DIB({DLX_IDinst_WB_data_eff[15], DLX_IDinst_WB_data_eff[14], DLX_IDinst_WB_data_eff[13], DLX_IDinst_WB_data_eff[12], DLX_IDinst_WB_data_eff[11], 
DLX_IDinst_WB_data_eff[10], DLX_IDinst_WB_data_eff[9], DLX_IDinst_WB_data_eff[8], DLX_RF_data_in[7], DLX_RF_data_in[6], DLX_RF_data_in[5], 
DLX_RF_data_in[4], DLX_RF_data_in[3], DLX_RF_data_in[2], DLX_RF_data_in[1], DLX_RF_data_in[0]}),
    .DOA({DLX_IDinst_reg_out_A_RF[15], DLX_IDinst_reg_out_A_RF[14], DLX_IDinst_reg_out_A_RF[13], DLX_IDinst_reg_out_A_RF[12], 
DLX_IDinst_reg_out_A_RF[11], DLX_IDinst_reg_out_A_RF[10], DLX_IDinst_reg_out_A_RF[9], DLX_IDinst_reg_out_A_RF[8], DLX_IDinst_reg_out_A_RF[7], 
DLX_IDinst_reg_out_A_RF[6], DLX_IDinst_reg_out_A_RF[5], DLX_IDinst_reg_out_A_RF[4], DLX_IDinst_reg_out_A_RF[3], DLX_IDinst_reg_out_A_RF[2], 
DLX_IDinst_reg_out_A_RF[1], DLX_IDinst_reg_out_A_RF[0]}),
    .DOB({\DLX_IDinst_RF_block0s0/DOB15 , \DLX_IDinst_RF_block0s0/DOB14 , \DLX_IDinst_RF_block0s0/DOB13 , \DLX_IDinst_RF_block0s0/DOB12 , 
\DLX_IDinst_RF_block0s0/DOB11 , \DLX_IDinst_RF_block0s0/DOB10 , \DLX_IDinst_RF_block0s0/DOB9 , \DLX_IDinst_RF_block0s0/DOB8 , 
\DLX_IDinst_RF_block0s0/DOB7 , \DLX_IDinst_RF_block0s0/DOB6 , \DLX_IDinst_RF_block0s0/DOB5 , \DLX_IDinst_RF_block0s0/DOB4 , 
\DLX_IDinst_RF_block0s0/DOB3 , \DLX_IDinst_RF_block0s0/DOB2 , \DLX_IDinst_RF_block0s0/DOB1 , \DLX_IDinst_RF_block0s0/DOB0 })
  );
  X_ZERO \DLX_IDinst_RF_block0s1/LOGIC_ZERO_115  (
    .O(\DLX_IDinst_RF_block0s1/LOGIC_ZERO )
  );
  defparam DLX_IDinst_RF_block0s1.INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block0s1.INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block0s1.INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block0s1.INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block0s1.INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block0s1.INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block0s1.INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block0s1.INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block0s1.INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block0s1.INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block0s1.INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block0s1.INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block0s1.INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block0s1.INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block0s1.INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block0s1.INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block0s1.SETUP_ALL = 2701;
  X_RAMB4_S16_S16 DLX_IDinst_RF_block0s1 (
    .CLKA(DLX_clk_IF_del),
    .CLKB(DLX_clk_ID),
    .ENA(DLX_IDinst__n0003),
    .ENB(DLX_IDinst__n0410),
    .RSTA(DLX_IDinst__n0004),
    .RSTB(\DLX_IDinst_RF_block0s1/LOGIC_ZERO ),
    .WEA(\DLX_IDinst_RF_block0s1/LOGIC_ZERO ),
    .WEB(DLX_MEMinst_reg_write_MEM),
    .GSR(GSR),
    .ADDRA({GLOBAL_LOGIC0_3, GLOBAL_LOGIC0_3, GLOBAL_LOGIC0_3, DLX_IDinst_regB_index[4], DLX_IDinst_regB_index[3], DLX_IDinst_regB_index[2], 
DLX_IDinst_regB_index[1], DLX_IDinst_regB_index[0]}),
    .ADDRB({GLOBAL_LOGIC0_3, GLOBAL_LOGIC0_3, GLOBAL_LOGIC0_3, DLX_MEMinst_reg_dst_out[4], DLX_MEMinst_reg_dst_out[3], DLX_MEMinst_reg_dst_out[2], 
DLX_MEMinst_reg_dst_out[1], DLX_MEMinst_reg_dst_out[0]}),
    .DIA({\DLX_IDinst_RF_block0s1/DIA15 , \DLX_IDinst_RF_block0s1/DIA14 , \DLX_IDinst_RF_block0s1/DIA13 , \DLX_IDinst_RF_block0s1/DIA12 , 
\DLX_IDinst_RF_block0s1/DIA11 , \DLX_IDinst_RF_block0s1/DIA10 , \DLX_IDinst_RF_block0s1/DIA9 , \DLX_IDinst_RF_block0s1/DIA8 , 
\DLX_IDinst_RF_block0s1/DIA7 , \DLX_IDinst_RF_block0s1/DIA6 , \DLX_IDinst_RF_block0s1/DIA5 , \DLX_IDinst_RF_block0s1/DIA4 , 
\DLX_IDinst_RF_block0s1/DIA3 , \DLX_IDinst_RF_block0s1/DIA2 , \DLX_IDinst_RF_block0s1/DIA1 , \DLX_IDinst_RF_block0s1/DIA0 }),
    .DIB({DLX_IDinst_WB_data_eff[15], DLX_IDinst_WB_data_eff[14], DLX_IDinst_WB_data_eff[13], DLX_IDinst_WB_data_eff[12], DLX_IDinst_WB_data_eff[11], 
DLX_IDinst_WB_data_eff[10], DLX_IDinst_WB_data_eff[9], DLX_IDinst_WB_data_eff[8], DLX_RF_data_in[7], DLX_RF_data_in[6], DLX_RF_data_in[5], 
DLX_RF_data_in[4], DLX_RF_data_in[3], DLX_RF_data_in[2], DLX_RF_data_in[1], DLX_RF_data_in[0]}),
    .DOA({DLX_IDinst_reg_out_B_RF[15], DLX_IDinst_reg_out_B_RF[14], DLX_IDinst_reg_out_B_RF[13], DLX_IDinst_reg_out_B_RF[12], 
DLX_IDinst_reg_out_B_RF[11], DLX_IDinst_reg_out_B_RF[10], DLX_IDinst_reg_out_B_RF[9], DLX_IDinst_reg_out_B_RF[8], DLX_IDinst_reg_out_B_RF[7], 
DLX_IDinst_reg_out_B_RF[6], DLX_IDinst_reg_out_B_RF[5], DLX_IDinst_reg_out_B_RF[4], DLX_IDinst_reg_out_B_RF[3], DLX_IDinst_reg_out_B_RF[2], 
DLX_IDinst_reg_out_B_RF[1], DLX_IDinst_reg_out_B_RF[0]}),
    .DOB({\DLX_IDinst_RF_block0s1/DOB15 , \DLX_IDinst_RF_block0s1/DOB14 , \DLX_IDinst_RF_block0s1/DOB13 , \DLX_IDinst_RF_block0s1/DOB12 , 
\DLX_IDinst_RF_block0s1/DOB11 , \DLX_IDinst_RF_block0s1/DOB10 , \DLX_IDinst_RF_block0s1/DOB9 , \DLX_IDinst_RF_block0s1/DOB8 , 
\DLX_IDinst_RF_block0s1/DOB7 , \DLX_IDinst_RF_block0s1/DOB6 , \DLX_IDinst_RF_block0s1/DOB5 , \DLX_IDinst_RF_block0s1/DOB4 , 
\DLX_IDinst_RF_block0s1/DOB3 , \DLX_IDinst_RF_block0s1/DOB2 , \DLX_IDinst_RF_block0s1/DOB1 , \DLX_IDinst_RF_block0s1/DOB0 })
  );
  X_ZERO \DLX_IDinst_RF_block1s0/LOGIC_ZERO_116  (
    .O(\DLX_IDinst_RF_block1s0/LOGIC_ZERO )
  );
  defparam DLX_IDinst_RF_block1s0.INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block1s0.INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block1s0.INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block1s0.INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block1s0.INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block1s0.INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block1s0.INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block1s0.INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block1s0.INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block1s0.INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block1s0.INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block1s0.INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block1s0.INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block1s0.INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block1s0.INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block1s0.INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block1s0.SETUP_ALL = 2701;
  X_RAMB4_S16_S16 DLX_IDinst_RF_block1s0 (
    .CLKA(DLX_clk_IF_del),
    .CLKB(DLX_clk_ID),
    .ENA(DLX_IDinst__n0000),
    .ENB(DLX_IDinst__n0410),
    .RSTA(DLX_IDinst__n0002),
    .RSTB(\DLX_IDinst_RF_block1s0/LOGIC_ZERO ),
    .WEA(\DLX_IDinst_RF_block1s0/LOGIC_ZERO ),
    .WEB(DLX_MEMinst_reg_write_MEM),
    .GSR(GSR),
    .ADDRA({GLOBAL_LOGIC0_0, GLOBAL_LOGIC0_0, GLOBAL_LOGIC0_0, DLX_IDinst_regA_index[4], DLX_IDinst_regA_index[3], DLX_IDinst_regA_index[2], 
DLX_IDinst_regA_index[1], DLX_IDinst_regA_index[0]}),
    .ADDRB({GLOBAL_LOGIC0_0, GLOBAL_LOGIC0_0, GLOBAL_LOGIC0_0, DLX_MEMinst_reg_dst_out[4], DLX_MEMinst_reg_dst_out[3], DLX_MEMinst_reg_dst_out[2], 
DLX_MEMinst_reg_dst_out[1], DLX_MEMinst_reg_dst_out[0]}),
    .DIA({\DLX_IDinst_RF_block1s0/DIA15 , \DLX_IDinst_RF_block1s0/DIA14 , \DLX_IDinst_RF_block1s0/DIA13 , \DLX_IDinst_RF_block1s0/DIA12 , 
\DLX_IDinst_RF_block1s0/DIA11 , \DLX_IDinst_RF_block1s0/DIA10 , \DLX_IDinst_RF_block1s0/DIA9 , \DLX_IDinst_RF_block1s0/DIA8 , 
\DLX_IDinst_RF_block1s0/DIA7 , \DLX_IDinst_RF_block1s0/DIA6 , \DLX_IDinst_RF_block1s0/DIA5 , \DLX_IDinst_RF_block1s0/DIA4 , 
\DLX_IDinst_RF_block1s0/DIA3 , \DLX_IDinst_RF_block1s0/DIA2 , \DLX_IDinst_RF_block1s0/DIA1 , \DLX_IDinst_RF_block1s0/DIA0 }),
    .DIB({DLX_IDinst_WB_data_eff[31], DLX_IDinst_WB_data_eff[30], DLX_IDinst_WB_data_eff[29], DLX_IDinst_WB_data_eff[28], DLX_IDinst_WB_data_eff[27], 
DLX_IDinst_WB_data_eff[26], DLX_IDinst_WB_data_eff[25], DLX_IDinst_WB_data_eff[24], DLX_IDinst_WB_data_eff[23], DLX_IDinst_WB_data_eff[22], 
DLX_IDinst_WB_data_eff[21], DLX_IDinst_WB_data_eff[20], DLX_IDinst_WB_data_eff[19], DLX_IDinst_WB_data_eff[18], DLX_IDinst_WB_data_eff[17], 
DLX_IDinst_WB_data_eff[16]}),
    .DOA({DLX_IDinst_reg_out_A_RF[31], DLX_IDinst_reg_out_A_RF[30], DLX_IDinst_reg_out_A_RF[29], DLX_IDinst_reg_out_A_RF[28], 
DLX_IDinst_reg_out_A_RF[27], DLX_IDinst_reg_out_A_RF[26], DLX_IDinst_reg_out_A_RF[25], DLX_IDinst_reg_out_A_RF[24], DLX_IDinst_reg_out_A_RF[23], 
DLX_IDinst_reg_out_A_RF[22], DLX_IDinst_reg_out_A_RF[21], DLX_IDinst_reg_out_A_RF[20], DLX_IDinst_reg_out_A_RF[19], DLX_IDinst_reg_out_A_RF[18], 
DLX_IDinst_reg_out_A_RF[17], DLX_IDinst_reg_out_A_RF[16]}),
    .DOB({\DLX_IDinst_RF_block1s0/DOB15 , \DLX_IDinst_RF_block1s0/DOB14 , \DLX_IDinst_RF_block1s0/DOB13 , \DLX_IDinst_RF_block1s0/DOB12 , 
\DLX_IDinst_RF_block1s0/DOB11 , \DLX_IDinst_RF_block1s0/DOB10 , \DLX_IDinst_RF_block1s0/DOB9 , \DLX_IDinst_RF_block1s0/DOB8 , 
\DLX_IDinst_RF_block1s0/DOB7 , \DLX_IDinst_RF_block1s0/DOB6 , \DLX_IDinst_RF_block1s0/DOB5 , \DLX_IDinst_RF_block1s0/DOB4 , 
\DLX_IDinst_RF_block1s0/DOB3 , \DLX_IDinst_RF_block1s0/DOB2 , \DLX_IDinst_RF_block1s0/DOB1 , \DLX_IDinst_RF_block1s0/DOB0 })
  );
  X_ZERO \DLX_IDinst_RF_block1s1/LOGIC_ZERO_117  (
    .O(\DLX_IDinst_RF_block1s1/LOGIC_ZERO )
  );
  defparam DLX_IDinst_RF_block1s1.INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block1s1.INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block1s1.INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block1s1.INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block1s1.INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block1s1.INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block1s1.INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block1s1.INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block1s1.INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block1s1.INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block1s1.INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block1s1.INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block1s1.INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block1s1.INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block1s1.INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block1s1.INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam DLX_IDinst_RF_block1s1.SETUP_ALL = 2701;
  X_RAMB4_S16_S16 DLX_IDinst_RF_block1s1 (
    .CLKA(DLX_clk_IF_del),
    .CLKB(DLX_clk_ID),
    .ENA(DLX_IDinst__n0003),
    .ENB(DLX_IDinst__n0410),
    .RSTA(DLX_IDinst__n0004),
    .RSTB(\DLX_IDinst_RF_block1s1/LOGIC_ZERO ),
    .WEA(\DLX_IDinst_RF_block1s1/LOGIC_ZERO ),
    .WEB(DLX_MEMinst_reg_write_MEM),
    .GSR(GSR),
    .ADDRA({GLOBAL_LOGIC0_4, GLOBAL_LOGIC0_4, GLOBAL_LOGIC0_4, DLX_IDinst_regB_index[4], DLX_IDinst_regB_index[3], DLX_IDinst_regB_index[2], 
DLX_IDinst_regB_index[1], DLX_IDinst_regB_index[0]}),
    .ADDRB({GLOBAL_LOGIC0_4, GLOBAL_LOGIC0_4, GLOBAL_LOGIC0_4, DLX_MEMinst_reg_dst_out[4], DLX_MEMinst_reg_dst_out[3], DLX_MEMinst_reg_dst_out[2], 
DLX_MEMinst_reg_dst_out[1], DLX_MEMinst_reg_dst_out[0]}),
    .DIA({\DLX_IDinst_RF_block1s1/DIA15 , \DLX_IDinst_RF_block1s1/DIA14 , \DLX_IDinst_RF_block1s1/DIA13 , \DLX_IDinst_RF_block1s1/DIA12 , 
\DLX_IDinst_RF_block1s1/DIA11 , \DLX_IDinst_RF_block1s1/DIA10 , \DLX_IDinst_RF_block1s1/DIA9 , \DLX_IDinst_RF_block1s1/DIA8 , 
\DLX_IDinst_RF_block1s1/DIA7 , \DLX_IDinst_RF_block1s1/DIA6 , \DLX_IDinst_RF_block1s1/DIA5 , \DLX_IDinst_RF_block1s1/DIA4 , 
\DLX_IDinst_RF_block1s1/DIA3 , \DLX_IDinst_RF_block1s1/DIA2 , \DLX_IDinst_RF_block1s1/DIA1 , \DLX_IDinst_RF_block1s1/DIA0 }),
    .DIB({DLX_IDinst_WB_data_eff[31], DLX_IDinst_WB_data_eff[30], DLX_IDinst_WB_data_eff[29], DLX_IDinst_WB_data_eff[28], DLX_IDinst_WB_data_eff[27], 
DLX_IDinst_WB_data_eff[26], DLX_IDinst_WB_data_eff[25], DLX_IDinst_WB_data_eff[24], DLX_IDinst_WB_data_eff[23], DLX_IDinst_WB_data_eff[22], 
DLX_IDinst_WB_data_eff[21], DLX_IDinst_WB_data_eff[20], DLX_IDinst_WB_data_eff[19], DLX_IDinst_WB_data_eff[18], DLX_IDinst_WB_data_eff[17], 
DLX_IDinst_WB_data_eff[16]}),
    .DOA({DLX_IDinst_reg_out_B_RF[31], DLX_IDinst_reg_out_B_RF[30], DLX_IDinst_reg_out_B_RF[29], DLX_IDinst_reg_out_B_RF[28], 
DLX_IDinst_reg_out_B_RF[27], DLX_IDinst_reg_out_B_RF[26], DLX_IDinst_reg_out_B_RF[25], DLX_IDinst_reg_out_B_RF[24], DLX_IDinst_reg_out_B_RF[23], 
DLX_IDinst_reg_out_B_RF[22], DLX_IDinst_reg_out_B_RF[21], DLX_IDinst_reg_out_B_RF[20], DLX_IDinst_reg_out_B_RF[19], DLX_IDinst_reg_out_B_RF[18], 
DLX_IDinst_reg_out_B_RF[17], DLX_IDinst_reg_out_B_RF[16]}),
    .DOB({\DLX_IDinst_RF_block1s1/DOB15 , \DLX_IDinst_RF_block1s1/DOB14 , \DLX_IDinst_RF_block1s1/DOB13 , \DLX_IDinst_RF_block1s1/DOB12 , 
\DLX_IDinst_RF_block1s1/DOB11 , \DLX_IDinst_RF_block1s1/DOB10 , \DLX_IDinst_RF_block1s1/DOB9 , \DLX_IDinst_RF_block1s1/DOB8 , 
\DLX_IDinst_RF_block1s1/DOB7 , \DLX_IDinst_RF_block1s1/DOB6 , \DLX_IDinst_RF_block1s1/DOB5 , \DLX_IDinst_RF_block1s1/DOB4 , 
\DLX_IDinst_RF_block1s1/DOB3 , \DLX_IDinst_RF_block1s1/DOB2 , \DLX_IDinst_RF_block1s1/DOB1 , \DLX_IDinst_RF_block1s1/DOB0 })
  );
  X_ONE \block0/LOGIC_ONE_118  (
    .O(\block0/LOGIC_ONE )
  );
  X_ZERO \block0/LOGIC_ZERO_119  (
    .O(\block0/LOGIC_ZERO )
  );
  defparam block0.INIT_00 = 256'h0000000000000000000000000000000000000000000000000000E80000000000;
  defparam block0.INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block0.INIT_02 = 256'hD0140001A000E8000001A00000280020203C00F4000000F00100200000E80000;
  defparam block0.INIT_03 = 256'h0205A02000003C001020280000244440A0000000C47801A000B4005CA0000000;
  defparam block0.INIT_04 = 256'h0028004C2020A0100C080400000000B401010021212101000820240006001F21;
  defparam block0.INIT_05 = 256'h008461FF603F9FA0A101002C0090202000002000C0010100250006001F200205;
  defparam block0.INIT_06 = 256'h019FA001002C009077002861605FA1A09F01010050019FC16061A09F01002C9F;
  defparam block0.INIT_07 = 256'hA0002C00905F606101019FA0A100B8FF6061773F01A0A1002C9F00EC5F60C19F;
  defparam block0.INIT_08 = 256'h0004A1A09F01019FA0A1002C013F9FA09F01A0A1002C9F00603F9F01A1A0019F;
  defparam block0.INIT_09 = 256'h0008000100080001000800010008000100080001000800010008000100080020;
  defparam block0.INIT_0A = 256'h0000000000EC0401001405200000010008202404010020010008200300200001;
  defparam block0.INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block0.INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block0.INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block0.INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block0.INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block0.SETUP_ALL = 2701;
  X_RAMB4_S8_S8 block0 (
    .CLKA(clk_DM_OBUF),
    .CLKB(DLX_clk_IF),
    .ENA(mask_0_OBUF),
    .ENB(\block0/LOGIC_ONE ),
    .RSTA(\block0/LOGIC_ZERO ),
    .RSTB(\block0/LOGIC_ZERO ),
    .WEA(DLX_EXinst_mem_write_EX),
    .WEB(\block0/LOGIC_ZERO ),
    .GSR(GSR),
    .ADDRA({DLX_EXinst_ALU_result[10], DLX_EXinst_ALU_result[9], DLX_EXinst_ALU_result[8], DLX_EXinst_ALU_result[7], DLX_EXinst_ALU_result[6], 
DLX_EXinst_ALU_result[5], DLX_EXinst_ALU_result[4], DLX_EXinst_ALU_result[3], DLX_EXinst_ALU_result[2]}),
    .ADDRB({DLX_IFinst_NPC[10], DLX_IFinst_NPC[9], DLX_IFinst_NPC[8], DLX_IFinst_NPC[7], DLX_IFinst_NPC[6], DLX_IFinst_NPC[5], DLX_IFinst_NPC[4], 
DLX_IFinst_NPC[3], DLX_IFinst_NPC[2]}),
    .DIA({DLX_EXinst_reg_out_B_EX[7], DLX_EXinst_reg_out_B_EX[6], DLX_EXinst_reg_out_B_EX[5], DLX_EXinst_reg_out_B_EX[4], DLX_EXinst_reg_out_B_EX[3], 
DLX_EXinst_reg_out_B_EX[2], DLX_EXinst_reg_out_B_EX[1], DLX_EXinst_reg_out_B_EX[0]}),
    .DIB({\block0/DIB7 , \block0/DIB6 , \block0/DIB5 , \block0/DIB4 , \block0/DIB3 , \block0/DIB2 , \block0/DIB1 , \block0/DIB0 }),
    .DOA({RAM_read_data[7], RAM_read_data[6], RAM_read_data[5], RAM_read_data[4], RAM_read_data[3], RAM_read_data[2], RAM_read_data[1], 
RAM_read_data[0]}),
    .DOB({IR[7], IR[6], IR[5], IR[4], IR[3], IR[2], IR[1], IR[0]})
  );
  X_ONE \block1/LOGIC_ONE_120  (
    .O(\block1/LOGIC_ONE )
  );
  X_ZERO \block1/LOGIC_ZERO_121  (
    .O(\block1/LOGIC_ZERO )
  );
  defparam block1.INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block1.INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block1.INIT_02 = 256'h00080000000000080000000001080088800800FF000000FF0000000000031000;
  defparam block1.INIT_03 = 256'h000000B80000080000C008000000080800080000FF0000000003000000080000;
  defparam block1.INIT_04 = 256'h000000006068000000000000000000FF000000A0A0A0000000A89800A08000B0;
  defparam block1.INIT_05 = 256'h00014A4A4A010000000000000000D0D00000F800FF000000B000B88000C80000;
  defparam block1.INIT_06 = 256'h00000000000000000000014A4A4A000000000000010000494A4A000000000000;
  defparam block1.INIT_07 = 256'h00000000004A4A4A000000000000004A4A4A000100000000000000004A4A4900;
  defparam block1.INIT_08 = 256'h0000000000000000000000000001000000000000000000000001000000000000;
  defparam block1.INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000040;
  defparam block1.INIT_0A = 256'h0000000000FF0000080800C8000000000008A000000000000000080000000000;
  defparam block1.INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block1.INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block1.INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block1.INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block1.INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block1.SETUP_ALL = 2701;
  X_RAMB4_S8_S8 block1 (
    .CLKA(clk_DM_OBUF),
    .CLKB(DLX_clk_IF),
    .ENA(mask_1_OBUF),
    .ENB(\block1/LOGIC_ONE ),
    .RSTA(\block1/LOGIC_ZERO ),
    .RSTB(\block1/LOGIC_ZERO ),
    .WEA(DLX_EXinst_mem_write_EX),
    .WEB(\block1/LOGIC_ZERO ),
    .GSR(GSR),
    .ADDRA({DLX_EXinst_ALU_result[10], DLX_EXinst_ALU_result[9], DLX_EXinst_ALU_result[8], DLX_EXinst_ALU_result[7], DLX_EXinst_ALU_result[6], 
DLX_EXinst_ALU_result[5], DLX_EXinst_ALU_result[4], DLX_EXinst_ALU_result[3], DLX_EXinst_ALU_result[2]}),
    .ADDRB({DLX_IFinst_NPC[10], DLX_IFinst_NPC[9], DLX_IFinst_NPC[8], DLX_IFinst_NPC[7], DLX_IFinst_NPC[6], DLX_IFinst_NPC[5], DLX_IFinst_NPC[4], 
DLX_IFinst_NPC[3], DLX_IFinst_NPC[2]}),
    .DIA({DLX_EXinst_reg_out_B_EX[15], DLX_EXinst_reg_out_B_EX[14], DLX_EXinst_reg_out_B_EX[13], DLX_EXinst_reg_out_B_EX[12], 
DLX_EXinst_reg_out_B_EX[11], DLX_EXinst_reg_out_B_EX[10], DLX_EXinst_reg_out_B_EX[9], DLX_EXinst_reg_out_B_EX[8]}),
    .DIB({\block1/DIB7 , \block1/DIB6 , \block1/DIB5 , \block1/DIB4 , \block1/DIB3 , \block1/DIB2 , \block1/DIB1 , \block1/DIB0 }),
    .DOA({RAM_read_data[15], RAM_read_data[14], RAM_read_data[13], RAM_read_data[12], RAM_read_data[11], RAM_read_data[10], RAM_read_data[9], 
RAM_read_data[8]}),
    .DOB({IR[15], IR[14], IR[13], IR[12], IR[11], IR[10], IR[9], IR[8]})
  );
  X_ONE \block2/LOGIC_ONE_122  (
    .O(\block2/LOGIC_ONE )
  );
  X_ZERO \block2/LOGIC_ZERO_123  (
    .O(\block2/LOGIC_ZERO )
  );
  defparam block2.INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block2.INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block2.INIT_02 = 256'h00EF0F31100000EF0F31100000EF0F00001F00FF000000FF2900000000096303;
  defparam block2.INIT_03 = 256'hD6F6120000E01F00000039190000181018391900A02531100000000018391900;
  defparam block2.INIT_04 = 256'h002000001F000EE0E0E0E0E000E0004052F795839817B500600074D39514F5D9;
  defparam block2.INIT_05 = 256'h0000575958545653525500A000204D7000E00C00C0CEAD36D736F817B82F39B9;
  defparam block2.INIT_06 = 256'h5957585500A000203900005758595253545556000052555758595354560020B9;
  defparam block2.INIT_07 = 256'h5800A000005253545556575859000052535455575658590020B9000052535456;
  defparam block2.INIT_08 = 256'h00005253545556575859000054575553545658590020B9000054565952535557;
  defparam block2.INIT_09 = 256'h00605B0800607B0800609B080060BB080060DB080060FB0800601B0800603B00;
  defparam block2.INIT_0A = 256'h000000E0000039183737180000E0010080009818140000010000000800C05608;
  defparam block2.INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block2.INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block2.INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block2.INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block2.INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block2.SETUP_ALL = 2701;
  X_RAMB4_S8_S8 block2 (
    .CLKA(clk_DM_OBUF),
    .CLKB(DLX_clk_IF),
    .ENA(mask_2_OBUF),
    .ENB(\block2/LOGIC_ONE ),
    .RSTA(\block2/LOGIC_ZERO ),
    .RSTB(\block2/LOGIC_ZERO ),
    .WEA(DLX_EXinst_mem_write_EX),
    .WEB(\block2/LOGIC_ZERO ),
    .GSR(GSR),
    .ADDRA({DLX_EXinst_ALU_result[10], DLX_EXinst_ALU_result[9], DLX_EXinst_ALU_result[8], DLX_EXinst_ALU_result[7], DLX_EXinst_ALU_result[6], 
DLX_EXinst_ALU_result[5], DLX_EXinst_ALU_result[4], DLX_EXinst_ALU_result[3], DLX_EXinst_ALU_result[2]}),
    .ADDRB({DLX_IFinst_NPC[10], DLX_IFinst_NPC[9], DLX_IFinst_NPC[8], DLX_IFinst_NPC[7], DLX_IFinst_NPC[6], DLX_IFinst_NPC[5], DLX_IFinst_NPC[4], 
DLX_IFinst_NPC[3], DLX_IFinst_NPC[2]}),
    .DIA({DLX_EXinst_reg_out_B_EX[23], DLX_EXinst_reg_out_B_EX[22], DLX_EXinst_reg_out_B_EX[21], DLX_EXinst_reg_out_B_EX[20], 
DLX_EXinst_reg_out_B_EX[19], DLX_EXinst_reg_out_B_EX[18], DLX_EXinst_reg_out_B_EX[17], DLX_EXinst_reg_out_B_EX[16]}),
    .DIB({\block2/DIB7 , \block2/DIB6 , \block2/DIB5 , \block2/DIB4 , \block2/DIB3 , \block2/DIB2 , \block2/DIB1 , \block2/DIB0 }),
    .DOA({RAM_read_data[23], RAM_read_data[22], RAM_read_data[21], RAM_read_data[20], RAM_read_data[19], RAM_read_data[18], RAM_read_data[17], 
RAM_read_data[16]}),
    .DOB({IR[23], IR[22], IR[21], IR[20], IR[19], IR[18], IR[17], IR[16]})
  );
  X_ONE \block3/LOGIC_ONE_124  (
    .O(\block3/LOGIC_ONE )
  );
  X_ZERO \block3/LOGIC_ZERO_125  (
    .O(\block3/LOGIC_ZERO )
  );
  defparam block3.INIT_00 = 256'h0000000000000000000000000000000000000000000000000054085454545454;
  defparam block3.INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block3.INIT_02 = 256'h0C253C2622540C253C2622540C253C0000AC540B5454540F2D540C545420243C;
  defparam block3.INIT_03 = 256'h525A2000544B8C540C00273C540CACAC2E273C54142E2626540C540C2E273C54;
  defparam block3.INIT_04 = 256'h5410540C000020ADADADADAD544B54162E26A202020026541200028E023C3202;
  defparam block3.INIT_05 = 256'h54082727272727272727541554160300544B0054152D25AF028F023C31035359;
  defparam block3.INIT_06 = 256'h2F2F2F27541554172E5408272727272727272F5408272F27272727272F54172D;
  defparam block3.INIT_07 = 256'h2F541554082F2F2F272F2F2F2F54082F2F2F2F2F2F2F2F54172D54082F2F2F27;
  defparam block3.INIT_08 = 256'h5408272727272F2F2F2F5408272F2F27272F2F2F54172D540827272F2727272F;
  defparam block3.INIT_09 = 256'h5413822554138225541382255413822554138225541382255413832554138300;
  defparam block3.INIT_0A = 256'h0000544B5417272FAF8F2000544B2054120002696D5408245415002D54168325;
  defparam block3.INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block3.INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block3.INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block3.INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block3.INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block3.SETUP_ALL = 2701;
  X_RAMB4_S8_S8 block3 (
    .CLKA(clk_DM_OBUF),
    .CLKB(DLX_clk_IF),
    .ENA(mask_3_OBUF),
    .ENB(\block3/LOGIC_ONE ),
    .RSTA(\block3/LOGIC_ZERO ),
    .RSTB(\block3/LOGIC_ZERO ),
    .WEA(DLX_EXinst_mem_write_EX),
    .WEB(\block3/LOGIC_ZERO ),
    .GSR(GSR),
    .ADDRA({DLX_EXinst_ALU_result[10], DLX_EXinst_ALU_result[9], DLX_EXinst_ALU_result[8], DLX_EXinst_ALU_result[7], DLX_EXinst_ALU_result[6], 
DLX_EXinst_ALU_result[5], DLX_EXinst_ALU_result[4], DLX_EXinst_ALU_result[3], DLX_EXinst_ALU_result[2]}),
    .ADDRB({DLX_IFinst_NPC[10], DLX_IFinst_NPC[9], DLX_IFinst_NPC[8], DLX_IFinst_NPC[7], DLX_IFinst_NPC[6], DLX_IFinst_NPC[5], DLX_IFinst_NPC[4], 
DLX_IFinst_NPC[3], DLX_IFinst_NPC[2]}),
    .DIA({DLX_EXinst_reg_out_B_EX[31], DLX_EXinst_reg_out_B_EX[30], DLX_EXinst_reg_out_B_EX[29], DLX_EXinst_reg_out_B_EX[28], 
DLX_EXinst_reg_out_B_EX[27], DLX_EXinst_reg_out_B_EX[26], DLX_EXinst_reg_out_B_EX[25], DLX_EXinst_reg_out_B_EX[24]}),
    .DIB({\block3/DIB7 , \block3/DIB6 , \block3/DIB5 , \block3/DIB4 , \block3/DIB3 , \block3/DIB2 , \block3/DIB1 , \block3/DIB0 }),
    .DOA({RAM_read_data[31], RAM_read_data[30], RAM_read_data[29], RAM_read_data[28], RAM_read_data[27], RAM_read_data[26], RAM_read_data[25], 
RAM_read_data[24]}),
    .DOB({IR_MSB_7_OBUF, IR_MSB_6_OBUF, IR_MSB_5_OBUF, IR_MSB_4_OBUF, IR_MSB_3_OBUF, IR_MSB_2_OBUF, IR_MSB_1_OBUF, IR_MSB_0_OBUF})
  );
  X_ZERO \vga0/LOGIC_ZERO_126  (
    .O(\vga0/LOGIC_ZERO )
  );
  X_ONE \vga0/LOGIC_ONE_127  (
    .O(\vga0/LOGIC_ONE )
  );
  defparam vga0.INIT_00 = 256'h000000000000000000001CE080F000008003FF00000000000000000000007F00;
  defparam vga0.INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga0.INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga0.INIT_03 = 256'h0000000000000000000000000000000000000000000000000000007000000000;
  defparam vga0.INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga0.INIT_05 = 256'h0000000000000000000000380000000000000000000000000000000000000070;
  defparam vga0.INIT_06 = 256'h0000E06000000000000000000000000000000000000000300000000000000000;
  defparam vga0.INIT_07 = 256'h00000000000001C000000000186060600000000000000000000001C000000000;
  defparam vga0.INIT_08 = 256'h00000000000080208000000000000000000000C0000000000000C02000000000;
  defparam vga0.INIT_09 = 256'h8000000000000000000000C000000000000080208000000000000000000000C0;
  defparam vga0.INIT_0A = 256'h000000C000000000000080208000000000000000000000800000000000008000;
  defparam vga0.INIT_0B = 256'h0000800080000000000000000000008000000000000080008000000000000000;
  defparam vga0.INIT_0C = 256'h0000000000000080000000000000800000000000000000000000008000000000;
  defparam vga0.INIT_0D = 256'h00000000000080008000000000000000000000C0000000000000802080000000;
  defparam vga0.INIT_0E = 256'h0000000000000008000000400000300000000000800000000000000000000080;
  defparam vga0.INIT_0F = 256'h0000003000001800000000000000000000000004000000600000300000000000;
  defparam vga0.SETUP_ALL = 2701;
  X_RAMB4_S1_S1 vga0 (
    .CLKA(clk_DM_OBUF),
    .CLKB(clkdiv_vga),
    .ENA(vga_select_6[1]),
    .ENB(\vga0/LOGIC_ONE ),
    .RSTA(reset_IBUF_1),
    .RSTB(reset_IBUF_1),
    .WEA(DLX_EXinst_mem_write_EX),
    .WEB(\vga0/LOGIC_ZERO ),
    .GSR(GSR),
    .ADDRA({DLX_EXinst_ALU_result[11], DLX_EXinst_ALU_result[10], DLX_EXinst_ALU_result[9], DLX_EXinst_ALU_result[8], DLX_EXinst_ALU_result[7], 
DLX_EXinst_ALU_result[6], DLX_EXinst_ALU_result[5], DLX_EXinst_ALU_result[4], DLX_EXinst_ALU_result[3], DLX_EXinst_ALU_result[2], 
DLX_EXinst_ALU_result[1], DLX_EXinst_ALU_result[0]}),
    .ADDRB({vga_address[11], vga_address[10], vga_address[9], vga_address[8], vga_address[7], vga_address[6], 
vga_top_vga1_Madd_addressout_inst_lut2_331, vga_top_vga1_gridhcounter[4], vga_top_vga1_gridhcounter[3], vga_top_vga1_gridhcounter[2], 
vga_top_vga1_gridhcounter[1], vga_top_vga1_gridhcounter[0]}),
    .DIA({DLX_EXinst_reg_out_B_EX[0]}),
    .DIB({\vga0/DIB0 }),
    .DOA({vram_out_cpu[0]}),
    .DOB({vram_out_vga[0]})
  );
  X_ZERO \vga1/LOGIC_ZERO_128  (
    .O(\vga1/LOGIC_ZERO )
  );
  X_ONE \vga1/LOGIC_ONE_129  (
    .O(\vga1/LOGIC_ONE )
  );
  defparam vga1.INIT_00 = 256'h000000010000000001400000000000300000180000000000000000000180001C;
  defparam vga1.INIT_01 = 256'h0000000000000018000010000000000100000000010000000000001800401000;
  defparam vga1.INIT_02 = 256'h0040100000000011000000000000000000000018004010000000000100000000;
  defparam vga1.INIT_03 = 256'h0000000000000000000000180040000000000001000000000000000000000008;
  defparam vga1.INIT_04 = 256'h0000000800000000000000000000000000000000000000180040000000000000;
  defparam vga1.INIT_05 = 256'h00000000C0000000C00000000000001000000000000000000000000000000000;
  defparam vga1.INIT_06 = 256'h00000000000000100000000000000000C0000000000000000000001000000000;
  defparam vga1.INIT_07 = 256'h0000000000000000C000000000000000000000000000000000000000C0000000;
  defparam vga1.INIT_08 = 256'h0000000000000000038000000000000000000000C00000000000000000000000;
  defparam vga1.INIT_09 = 256'h0380000000000000000000000000000000000000038000000000000000000000;
  defparam vga1.INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga1.INIT_0B = 256'h00000000C000000000000000000000000000000000000000C000000000000000;
  defparam vga1.INIT_0C = 256'h00000000000000000000000000000000C0000000000000000000000000000000;
  defparam vga1.INIT_0D = 256'h00000000000000000000000000000000000000000000000000000000C0000000;
  defparam vga1.INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga1.INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga1.SETUP_ALL = 2701;
  X_RAMB4_S1_S1 vga1 (
    .CLKA(clk_DM_OBUF),
    .CLKB(clkdiv_vga),
    .ENA(vga_select_6[2]),
    .ENB(\vga1/LOGIC_ONE ),
    .RSTA(reset_IBUF_1),
    .RSTB(reset_IBUF_1),
    .WEA(DLX_EXinst_mem_write_EX),
    .WEB(\vga1/LOGIC_ZERO ),
    .GSR(GSR),
    .ADDRA({DLX_EXinst_ALU_result[11], DLX_EXinst_ALU_result[10], DLX_EXinst_ALU_result[9], DLX_EXinst_ALU_result[8], DLX_EXinst_ALU_result[7], 
DLX_EXinst_ALU_result[6], DLX_EXinst_ALU_result[5], DLX_EXinst_ALU_result[4], DLX_EXinst_ALU_result[3], DLX_EXinst_ALU_result[2], 
DLX_EXinst_ALU_result[1], DLX_EXinst_ALU_result[0]}),
    .ADDRB({vga_address[11], vga_address[10], vga_address[9], vga_address[8], vga_address[7], vga_address[6], 
vga_top_vga1_Madd_addressout_inst_lut2_331, vga_top_vga1_gridhcounter[4], vga_top_vga1_gridhcounter[3], vga_top_vga1_gridhcounter[2], 
vga_top_vga1_gridhcounter[1], vga_top_vga1_gridhcounter[0]}),
    .DIA({DLX_EXinst_reg_out_B_EX[0]}),
    .DIB({\vga1/DIB0 }),
    .DOA({vram_out_cpu[1]}),
    .DOB({vram_out_vga[1]})
  );
  X_ZERO \vga2/LOGIC_ZERO_130  (
    .O(\vga2/LOGIC_ZERO )
  );
  X_ONE \vga2/LOGIC_ONE_131  (
    .O(\vga2/LOGIC_ONE )
  );
  defparam vga2.INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga2.INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga2.INIT_02 = 256'h0000000000000000000000000000001C00000000800000008000000000000000;
  defparam vga2.INIT_03 = 256'h000000000000001C000000000000000000000000000000000000001C00000000;
  defparam vga2.INIT_04 = 256'h0000000080000000800000000000000000000000000000000000000000000000;
  defparam vga2.INIT_05 = 256'h8000000000000000000000000000000080000000800000000000000000000000;
  defparam vga2.INIT_06 = 256'h0000000000000000800000008000000000000000000000000000000080000000;
  defparam vga2.INIT_07 = 256'h0000000000000000000000000000000000000000800000000000000000000000;
  defparam vga2.INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga2.INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga2.INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga2.INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga2.INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga2.INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga2.INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga2.INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga2.SETUP_ALL = 2701;
  X_RAMB4_S1_S1 vga2 (
    .CLKA(clk_DM_OBUF),
    .CLKB(clkdiv_vga),
    .ENA(vga_select_6[3]),
    .ENB(\vga2/LOGIC_ONE ),
    .RSTA(reset_IBUF_1),
    .RSTB(reset_IBUF_1),
    .WEA(DLX_EXinst_mem_write_EX),
    .WEB(\vga2/LOGIC_ZERO ),
    .GSR(GSR),
    .ADDRA({DLX_EXinst_ALU_result[11], DLX_EXinst_ALU_result[10], DLX_EXinst_ALU_result[9], DLX_EXinst_ALU_result[8], DLX_EXinst_ALU_result[7], 
DLX_EXinst_ALU_result[6], DLX_EXinst_ALU_result[5], DLX_EXinst_ALU_result[4], DLX_EXinst_ALU_result[3], DLX_EXinst_ALU_result[2], 
DLX_EXinst_ALU_result[1], DLX_EXinst_ALU_result[0]}),
    .ADDRB({vga_address[11], vga_address[10], vga_address[9], vga_address[8], vga_address[7], vga_address[6], 
vga_top_vga1_Madd_addressout_inst_lut2_331, vga_top_vga1_gridhcounter[4], vga_top_vga1_gridhcounter[3], vga_top_vga1_gridhcounter[2], 
vga_top_vga1_gridhcounter[1], vga_top_vga1_gridhcounter[0]}),
    .DIA({DLX_EXinst_reg_out_B_EX[0]}),
    .DIB({\vga2/DIB0 }),
    .DOA({vram_out_cpu[2]}),
    .DOB({vram_out_vga[2]})
  );
  X_ZERO \vga3/LOGIC_ZERO_132  (
    .O(\vga3/LOGIC_ZERO )
  );
  X_ONE \vga3/LOGIC_ONE_133  (
    .O(\vga3/LOGIC_ONE )
  );
  defparam vga3.INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga3.INIT_01 = 256'h0000000000000000000000000000000000000400000000000000000000000000;
  defparam vga3.INIT_02 = 256'h0000000000000000000012000000000000000000000000000000000000000C00;
  defparam vga3.INIT_03 = 256'h0000000000000000000000000000000000001800000000000000000000000000;
  defparam vga3.INIT_04 = 256'h0000000000000000000008000000000000003FF0000000000000000000000800;
  defparam vga3.INIT_05 = 256'h0000038000000000000000000000000000000000000000000000000000000000;
  defparam vga3.INIT_06 = 256'h0000000000000000000000000000008000000000000000000000000000000000;
  defparam vga3.INIT_07 = 256'h01C000000000000000000000000000000000000000000000010000000003FF00;
  defparam vga3.INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga3.INIT_09 = 256'h0000E00000000000000000000000000000000000000080000000000000000000;
  defparam vga3.INIT_0A = 256'h0000000000000000000000000000004000000000000000000000000000000000;
  defparam vga3.INIT_0B = 256'h00000000000001F000000000000000000000000000000000000000E000000000;
  defparam vga3.INIT_0C = 256'h00000000000000000000000000000000000003F8000000000000000000000000;
  defparam vga3.INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga3.INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga3.INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga3.SETUP_ALL = 2701;
  X_RAMB4_S1_S1 vga3 (
    .CLKA(clk_DM_OBUF),
    .CLKB(clkdiv_vga),
    .ENA(vga_select_6[4]),
    .ENB(\vga3/LOGIC_ONE ),
    .RSTA(reset_IBUF_1),
    .RSTB(reset_IBUF_1),
    .WEA(DLX_EXinst_mem_write_EX),
    .WEB(\vga3/LOGIC_ZERO ),
    .GSR(GSR),
    .ADDRA({DLX_EXinst_ALU_result[11], DLX_EXinst_ALU_result[10], DLX_EXinst_ALU_result[9], DLX_EXinst_ALU_result[8], DLX_EXinst_ALU_result[7], 
DLX_EXinst_ALU_result[6], DLX_EXinst_ALU_result[5], DLX_EXinst_ALU_result[4], DLX_EXinst_ALU_result[3], DLX_EXinst_ALU_result[2], 
DLX_EXinst_ALU_result[1], DLX_EXinst_ALU_result[0]}),
    .ADDRB({vga_address[11], vga_address[10], vga_address[9], vga_address[8], vga_address[7], vga_address[6], 
vga_top_vga1_Madd_addressout_inst_lut2_331, vga_top_vga1_gridhcounter[4], vga_top_vga1_gridhcounter[3], vga_top_vga1_gridhcounter[2], 
vga_top_vga1_gridhcounter[1], vga_top_vga1_gridhcounter[0]}),
    .DIA({DLX_EXinst_reg_out_B_EX[0]}),
    .DIB({\vga3/DIB0 }),
    .DOA({vram_out_cpu[3]}),
    .DOB({vram_out_vga[3]})
  );
  X_ZERO \vga4/LOGIC_ZERO_134  (
    .O(\vga4/LOGIC_ZERO )
  );
  X_ONE \vga4/LOGIC_ONE_135  (
    .O(\vga4/LOGIC_ONE )
  );
  defparam vga4.INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga4.INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga4.INIT_02 = 256'h00000000000000000003E000000000000000000000000000000000000003E000;
  defparam vga4.INIT_03 = 256'h0003E000000000000000000000000000000000000003E0000000000000000000;
  defparam vga4.INIT_04 = 256'h0000000000000000000000000003E00000000000000000000000000000000000;
  defparam vga4.INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga4.INIT_06 = 256'h0000000000000000006000000000000000700000000000000000000000C00000;
  defparam vga4.INIT_07 = 256'h000C00000000000000100000001E000000000000003000000000000000700000;
  defparam vga4.INIT_08 = 256'h0000000000000000000000000006000000000000000000000000000000000000;
  defparam vga4.INIT_09 = 256'h0000000000060000000000000000000000000000000000000006000000000000;
  defparam vga4.INIT_0A = 256'h00000000000000000000000000000000000600F0000000000000000000000000;
  defparam vga4.INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga4.INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga4.INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga4.INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga4.INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga4.SETUP_ALL = 2701;
  X_RAMB4_S1_S1 vga4 (
    .CLKA(clk_DM_OBUF),
    .CLKB(clkdiv_vga),
    .ENA(vga_select_6[5]),
    .ENB(\vga4/LOGIC_ONE ),
    .RSTA(reset_IBUF_1),
    .RSTB(reset_IBUF_1),
    .WEA(DLX_EXinst_mem_write_EX),
    .WEB(\vga4/LOGIC_ZERO ),
    .GSR(GSR),
    .ADDRA({DLX_EXinst_ALU_result[11], DLX_EXinst_ALU_result[10], DLX_EXinst_ALU_result[9], DLX_EXinst_ALU_result[8], DLX_EXinst_ALU_result[7], 
DLX_EXinst_ALU_result[6], DLX_EXinst_ALU_result[5], DLX_EXinst_ALU_result[4], DLX_EXinst_ALU_result[3], DLX_EXinst_ALU_result[2], 
DLX_EXinst_ALU_result[1], DLX_EXinst_ALU_result[0]}),
    .ADDRB({vga_address[11], vga_address[10], vga_address[9], vga_address[8], vga_address[7], vga_address[6], 
vga_top_vga1_Madd_addressout_inst_lut2_331, vga_top_vga1_gridhcounter[4], vga_top_vga1_gridhcounter[3], vga_top_vga1_gridhcounter[2], 
vga_top_vga1_gridhcounter[1], vga_top_vga1_gridhcounter[0]}),
    .DIA({DLX_EXinst_reg_out_B_EX[0]}),
    .DIB({\vga4/DIB0 }),
    .DOA({vram_out_cpu[4]}),
    .DOB({vram_out_vga[4]})
  );
  X_MUX2 DLX_EXinst_Ker64882106 (
    .IA(N127639),
    .IB(N127641),
    .SEL(DLX_IDinst_reg_out_B_3_1),
    .O(\N108593/F5MUX )
  );
  defparam DLX_EXinst_Ker64882106_G.INIT = 16'h00C0;
  X_LUT4 DLX_EXinst_Ker64882106_G (
    .ADR0(VCC),
    .ADR1(N111221),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(DLX_IDinst_reg_out_B[5]),
    .O(N127641)
  );
  defparam DLX_EXinst_Ker64882106_F.INIT = 16'hFFA8;
  X_LUT4 DLX_EXinst_Ker64882106_F (
    .ADR0(N111221),
    .ADR1(CHOICE3145),
    .ADR2(CHOICE3139),
    .ADR3(CHOICE3152),
    .O(N127639)
  );
  X_BUF \N108593/XUSED  (
    .I(\N108593/F5MUX ),
    .O(N108593)
  );
  X_MUX2 DLX_EXinst_Ker64867103 (
    .IA(N127699),
    .IB(N127701),
    .SEL(DLX_IDinst_reg_out_B_2_1),
    .O(\CHOICE3132/F5MUX )
  );
  defparam DLX_EXinst_Ker64867103_G.INIT = 16'h4440;
  X_LUT4 DLX_EXinst_Ker64867103_G (
    .ADR0(DLX_IDinst_reg_out_B_3_1),
    .ADR1(DLX_EXinst_N66494),
    .ADR2(CHOICE1306),
    .ADR3(CHOICE1312),
    .O(N127701)
  );
  defparam DLX_EXinst_Ker64867103_F.INIT = 16'h8C80;
  X_LUT4 DLX_EXinst_Ker64867103_F (
    .ADR0(\DLX_EXinst_Mshift__n0026_Sh[29] ),
    .ADR1(DLX_EXinst_N66494),
    .ADR2(DLX_IDinst_reg_out_B_3_1),
    .ADR3(\DLX_EXinst_Mshift__n0026_Sh[21] ),
    .O(N127699)
  );
  X_BUF \CHOICE3132/XUSED  (
    .I(\CHOICE3132/F5MUX ),
    .O(CHOICE3132)
  );
  X_MUX2 DLX_EXinst_Ker64887102 (
    .IA(N127684),
    .IB(N127686),
    .SEL(DLX_IDinst_reg_out_B_3_1),
    .O(\N107934/F5MUX )
  );
  defparam DLX_EXinst_Ker64887102_G.INIT = 16'h0808;
  X_LUT4 DLX_EXinst_Ker64887102_G (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(N111221),
    .ADR2(DLX_IDinst_reg_out_B[5]),
    .ADR3(VCC),
    .O(N127686)
  );
  defparam DLX_EXinst_Ker64887102_F.INIT = 16'hFCF8;
  X_LUT4 DLX_EXinst_Ker64887102_F (
    .ADR0(CHOICE3032),
    .ADR1(N111221),
    .ADR2(CHOICE3045),
    .ADR3(CHOICE3038),
    .O(N127684)
  );
  X_BUF \N107934/XUSED  (
    .I(\N107934/F5MUX ),
    .O(N107934)
  );
  X_MUX2 DLX_IDinst__n012269 (
    .IA(N127924),
    .IB(N127926),
    .SEL(DLX_IDinst_IR_latched[28]),
    .O(\CHOICE3311/F5MUX )
  );
  defparam DLX_IDinst__n012269_G.INIT = 16'h3000;
  X_LUT4 DLX_IDinst__n012269_G (
    .ADR0(VCC),
    .ADR1(N126675),
    .ADR2(DLX_IDinst__n0377),
    .ADR3(DLX_IDinst_N70909),
    .O(N127926)
  );
  defparam DLX_IDinst__n012269_F.INIT = 16'hB000;
  X_LUT4 DLX_IDinst__n012269_F (
    .ADR0(DLX_IDinst_N70985),
    .ADR1(DLX_IDinst_IR_latched[30]),
    .ADR2(DLX_IDinst_IR_latched[27]),
    .ADR3(DLX_IDinst_N70909),
    .O(N127924)
  );
  X_BUF \CHOICE3311/XUSED  (
    .I(\CHOICE3311/F5MUX ),
    .O(CHOICE3311)
  );
  X_MUX2 \DLX_EXinst__n0006<28>99_SW0  (
    .IA(N128064),
    .IB(N128066),
    .SEL(DLX_IDinst_IR_function_field[4]),
    .O(\N126636/F5MUX )
  );
  defparam \DLX_EXinst__n0006<28>99_SW0_G .INIT = 16'hC8C8;
  X_LUT4 \DLX_EXinst__n0006<28>99_SW0_G  (
    .ADR0(CHOICE1042),
    .ADR1(DLX_EXinst_N66202),
    .ADR2(CHOICE1048),
    .ADR3(VCC),
    .O(N128066)
  );
  defparam \DLX_EXinst__n0006<28>99_SW0_F .INIT = 16'hA0C0;
  X_LUT4 \DLX_EXinst__n0006<28>99_SW0_F  (
    .ADR0(N97960),
    .ADR1(CHOICE5189),
    .ADR2(DLX_EXinst_N66202),
    .ADR3(DLX_IDinst_IR_function_field[2]),
    .O(N128064)
  );
  X_BUF \N126636/XUSED  (
    .I(\N126636/F5MUX ),
    .O(N126636)
  );
  X_MUX2 DLX_IDinst__n033958 (
    .IA(N128094),
    .IB(N128096),
    .SEL(DLX_IDinst_IR_latched[30]),
    .O(\CHOICE1402/F5MUX )
  );
  defparam DLX_IDinst__n033958_G.INIT = 16'h7A7E;
  X_LUT4 DLX_IDinst__n033958_G (
    .ADR0(DLX_IDinst_IR_latched[29]),
    .ADR1(DLX_IDinst_IR_latched[28]),
    .ADR2(DLX_IDinst_IR_latched[27]),
    .ADR3(DLX_IDinst_IR_latched[26]),
    .O(N128096)
  );
  defparam DLX_IDinst__n033958_F.INIT = 16'h7F00;
  X_LUT4 DLX_IDinst__n033958_F (
    .ADR0(DLX_IDinst_IR_latched[26]),
    .ADR1(DLX_IDinst_IR_latched[28]),
    .ADR2(DLX_IDinst_IR_latched[27]),
    .ADR3(DLX_IDinst_IR_latched[29]),
    .O(N128094)
  );
  X_BUF \CHOICE1402/XUSED  (
    .I(\CHOICE1402/F5MUX ),
    .O(CHOICE1402)
  );
  X_MUX2 DLX_IFlc_md_Mmux_outp2_inst_mux_f5_3111 (
    .IA(N127944),
    .IB(N127946),
    .SEL(delay_selectIF_0_IBUF),
    .O(\DLX_IFlc_md_outp2/F5MUX )
  );
  defparam DLX_IFlc_md_Mmux_outp2_inst_mux_f5_3111_G.INIT = 16'hFA0A;
  X_LUT4 DLX_IFlc_md_Mmux_outp2_inst_mux_f5_3111_G (
    .ADR0(DLX_IFlc_md_wint30),
    .ADR1(VCC),
    .ADR2(delay_selectIF_1_IBUF),
    .ADR3(DLX_IFlc_md_wint40),
    .O(N127946)
  );
  defparam DLX_IFlc_md_Mmux_outp2_inst_mux_f5_3111_F.INIT = 16'hF3C0;
  X_LUT4 DLX_IFlc_md_Mmux_outp2_inst_mux_f5_3111_F (
    .ADR0(VCC),
    .ADR1(delay_selectIF_1_IBUF),
    .ADR2(DLX_IFlc_md_wint34),
    .ADR3(DLX_IFlc_md_wint26),
    .O(N127944)
  );
  X_BUF \DLX_IFlc_md_outp2/XUSED  (
    .I(\DLX_IFlc_md_outp2/F5MUX ),
    .O(DLX_IFlc_md_outp2)
  );
  X_MUX2 DLX_IDlc_md_Mmux_outp2_inst_mux_f5_4111 (
    .IA(N127939),
    .IB(N127941),
    .SEL(delay_selectID_0_IBUF),
    .O(\DLX_IDlc_md_outp2/F5MUX )
  );
  defparam DLX_IDlc_md_Mmux_outp2_inst_mux_f5_4111_G.INIT = 16'hFA50;
  X_LUT4 DLX_IDlc_md_Mmux_outp2_inst_mux_f5_4111_G (
    .ADR0(delay_selectID_1_IBUF),
    .ADR1(VCC),
    .ADR2(DLX_IDlc_md_wint30),
    .ADR3(DLX_IDlc_md_wint40),
    .O(N127941)
  );
  defparam DLX_IDlc_md_Mmux_outp2_inst_mux_f5_4111_F.INIT = 16'hFA50;
  X_LUT4 DLX_IDlc_md_Mmux_outp2_inst_mux_f5_4111_F (
    .ADR0(delay_selectID_1_IBUF),
    .ADR1(VCC),
    .ADR2(DLX_IDlc_md_wint26),
    .ADR3(DLX_IDlc_md_wint34),
    .O(N127939)
  );
  X_BUF \DLX_IDlc_md_outp2/XUSED  (
    .I(\DLX_IDlc_md_outp2/F5MUX ),
    .O(DLX_IDlc_md_outp2)
  );
  X_MUX2 DLX_EXlc_md_Mmux_outp2_inst_mux_f5_5111 (
    .IA(N127934),
    .IB(N127936),
    .SEL(delay_selectEX_0_IBUF),
    .O(\DLX_EXlc_md_outp2/F5MUX )
  );
  defparam DLX_EXlc_md_Mmux_outp2_inst_mux_f5_5111_G.INIT = 16'hBB88;
  X_LUT4 DLX_EXlc_md_Mmux_outp2_inst_mux_f5_5111_G (
    .ADR0(DLX_EXlc_md_wint40),
    .ADR1(delay_selectEX_1_IBUF),
    .ADR2(VCC),
    .ADR3(DLX_EXlc_md_wint30),
    .O(N127936)
  );
  defparam DLX_EXlc_md_Mmux_outp2_inst_mux_f5_5111_F.INIT = 16'hBB88;
  X_LUT4 DLX_EXlc_md_Mmux_outp2_inst_mux_f5_5111_F (
    .ADR0(DLX_EXlc_md_wint34),
    .ADR1(delay_selectEX_1_IBUF),
    .ADR2(VCC),
    .ADR3(DLX_EXlc_md_wint26),
    .O(N127934)
  );
  X_BUF \DLX_EXlc_md_outp2/XUSED  (
    .I(\DLX_EXlc_md_outp2/F5MUX ),
    .O(DLX_EXlc_md_outp2)
  );
  X_MUX2 \DLX_EXinst__n0006<2>71  (
    .IA(N127879),
    .IB(N127881),
    .SEL(DLX_IDinst_IR_function_field[3]),
    .O(\CHOICE5509/F5MUX )
  );
  defparam \DLX_EXinst__n0006<2>71_G .INIT = 16'h5140;
  X_LUT4 \DLX_EXinst__n0006<2>71_G  (
    .ADR0(DLX_IDinst_IR_function_field[2]),
    .ADR1(DLX_IDinst_IR_function_field[0]),
    .ADR2(DLX_EXinst_N62986),
    .ADR3(DLX_EXinst_N63489),
    .O(N127881)
  );
  defparam \DLX_EXinst__n0006<2>71_F .INIT = 16'h0A0C;
  X_LUT4 \DLX_EXinst__n0006<2>71_F  (
    .ADR0(DLX_EXinst_N65165),
    .ADR1(DLX_EXinst_N64474),
    .ADR2(DLX_IDinst_IR_function_field[2]),
    .ADR3(DLX_IDinst_IR_function_field[0]),
    .O(N127879)
  );
  X_BUF \CHOICE5509/XUSED  (
    .I(\CHOICE5509/F5MUX ),
    .O(CHOICE5509)
  );
  X_MUX2 DLX_MEMlc_md_Mmux_outp2_inst_mux_f5_6111 (
    .IA(N127929),
    .IB(N127931),
    .SEL(delay_selectMEM_0_IBUF),
    .O(\DLX_MEMlc_md_outp2/F5MUX )
  );
  defparam DLX_MEMlc_md_Mmux_outp2_inst_mux_f5_6111_G.INIT = 16'hF0AA;
  X_LUT4 DLX_MEMlc_md_Mmux_outp2_inst_mux_f5_6111_G (
    .ADR0(DLX_MEMlc_md_wint10),
    .ADR1(VCC),
    .ADR2(DLX_MEMlc_md_wint20),
    .ADR3(delay_selectMEM_1_IBUF),
    .O(N127931)
  );
  defparam DLX_MEMlc_md_Mmux_outp2_inst_mux_f5_6111_F.INIT = 16'hCCF0;
  X_LUT4 DLX_MEMlc_md_Mmux_outp2_inst_mux_f5_6111_F (
    .ADR0(VCC),
    .ADR1(DLX_MEMlc_md_wint14),
    .ADR2(DLX_MEMlc_md_wint8),
    .ADR3(delay_selectMEM_1_IBUF),
    .O(N127929)
  );
  X_BUF \DLX_MEMlc_md_outp2/XUSED  (
    .I(\DLX_MEMlc_md_outp2/F5MUX ),
    .O(DLX_MEMlc_md_outp2)
  );
  X_MUX2 \DLX_EXinst__n0006<29>99_SW0  (
    .IA(N127779),
    .IB(N127781),
    .SEL(DLX_IDinst_IR_function_field[4]),
    .O(\N126486/F5MUX )
  );
  defparam \DLX_EXinst__n0006<29>99_SW0_G .INIT = 16'hA808;
  X_LUT4 \DLX_EXinst__n0006<29>99_SW0_G  (
    .ADR0(DLX_EXinst_N66202),
    .ADR1(N93279),
    .ADR2(DLX_IDinst_IR_function_field[3]),
    .ADR3(DLX_EXinst_N62821),
    .O(N127781)
  );
  defparam \DLX_EXinst__n0006<29>99_SW0_F .INIT = 16'hA280;
  X_LUT4 \DLX_EXinst__n0006<29>99_SW0_F  (
    .ADR0(DLX_EXinst_N66202),
    .ADR1(DLX_IDinst_IR_function_field[2]),
    .ADR2(N97665),
    .ADR3(CHOICE5341),
    .O(N127779)
  );
  X_BUF \N126486/XUSED  (
    .I(\N126486/F5MUX ),
    .O(N126486)
  );
  X_MUX2 DLX_IDinst_Ker69961 (
    .IA(N127884),
    .IB(N127886),
    .SEL(DLX_IDinst__n0135),
    .O(\DLX_IDinst_N69963/F5MUX )
  );
  defparam DLX_IDinst_Ker69961_G.INIT = 16'h0333;
  X_LUT4 DLX_IDinst_Ker69961_G (
    .ADR0(VCC),
    .ADR1(N98613),
    .ADR2(DLX_IDinst_N70647),
    .ADR3(N98420),
    .O(N127886)
  );
  defparam DLX_IDinst_Ker69961_F.INIT = 16'h550C;
  X_LUT4 DLX_IDinst_Ker69961_F (
    .ADR0(DLX_IDinst__n0344),
    .ADR1(DLX_IDinst__n0345),
    .ADR2(DLX_IDinst__n0347),
    .ADR3(DLX_IDinst__n0136),
    .O(N127884)
  );
  X_BUF \DLX_IDinst_N69963/XUSED  (
    .I(\DLX_IDinst_N69963/F5MUX ),
    .O(DLX_IDinst_N69963)
  );
  X_MUX2 DM_delay_inst_Mmux_outp_inst_mux_f5_1111 (
    .IA(N127999),
    .IB(N128001),
    .SEL(delay_selectDM_0_IBUF),
    .O(\clk_EX_del/F5MUX )
  );
  defparam DM_delay_inst_Mmux_outp_inst_mux_f5_1111_G.INIT = 16'hF5A0;
  X_LUT4 DM_delay_inst_Mmux_outp_inst_mux_f5_1111_G (
    .ADR0(delay_selectDM_1_IBUF),
    .ADR1(VCC),
    .ADR2(DM_delay_inst_wint40),
    .ADR3(DM_delay_inst_wint26),
    .O(N128001)
  );
  defparam DM_delay_inst_Mmux_outp_inst_mux_f5_1111_F.INIT = 16'hB8B8;
  X_LUT4 DM_delay_inst_Mmux_outp_inst_mux_f5_1111_F (
    .ADR0(DM_delay_inst_wint34),
    .ADR1(delay_selectDM_1_IBUF),
    .ADR2(DM_delay_inst_wint20),
    .ADR3(VCC),
    .O(N127999)
  );
  X_BUF \clk_EX_del/XUSED  (
    .I(\clk_EX_del/F5MUX ),
    .O(clk_EX_del)
  );
  X_MUX2 \DLX_IFinst__n0003<10>  (
    .IA(N127694),
    .IB(N127696),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[10])
  );
  defparam \DLX_IFinst__n0003<10>_G .INIT = 16'hFC30;
  X_LUT4 \DLX_IFinst__n0003<10>_G  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(DLX_IFinst_IR_previous[10]),
    .ADR3(IR[10]),
    .O(N127696)
  );
  defparam \DLX_IFinst__n0003<10>_F .INIT = 16'hF2D0;
  X_LUT4 \DLX_IFinst__n0003<10>_F  (
    .ADR0(DLX_IFinst_stalled),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(IR[10]),
    .ADR3(DLX_IFinst_IR_curr[10]),
    .O(N127694)
  );
  X_MUX2 \DLX_IFinst__n0003<11>  (
    .IA(N127784),
    .IB(N127786),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[11])
  );
  defparam \DLX_IFinst__n0003<11>_G .INIT = 16'hBB88;
  X_LUT4 \DLX_IFinst__n0003<11>_G  (
    .ADR0(IR[11]),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(VCC),
    .ADR3(DLX_IFinst_IR_previous[11]),
    .O(N127786)
  );
  defparam \DLX_IFinst__n0003<11>_F .INIT = 16'hBA8A;
  X_LUT4 \DLX_IFinst__n0003<11>_F  (
    .ADR0(IR[11]),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(DLX_IFinst_stalled),
    .ADR3(DLX_IFinst_IR_curr[11]),
    .O(N127784)
  );
  X_MUX2 \DLX_IFinst__n0003<12>  (
    .IA(N127904),
    .IB(N127906),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[12])
  );
  defparam \DLX_IFinst__n0003<12>_G .INIT = 16'hF0AA;
  X_LUT4 \DLX_IFinst__n0003<12>_G  (
    .ADR0(DLX_IFinst_IR_previous[12]),
    .ADR1(VCC),
    .ADR2(IR[12]),
    .ADR3(DLX_IDinst_branch_sig),
    .O(N127906)
  );
  defparam \DLX_IFinst__n0003<12>_F .INIT = 16'hF2D0;
  X_LUT4 \DLX_IFinst__n0003<12>_F  (
    .ADR0(DLX_IFinst_stalled),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(IR[12]),
    .ADR3(DLX_IFinst_IR_curr[12]),
    .O(N127904)
  );
  X_MUX2 \DLX_IFinst__n0003<20>  (
    .IA(N127674),
    .IB(N127676),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[20])
  );
  defparam \DLX_IFinst__n0003<20>_G .INIT = 16'hE2E2;
  X_LUT4 \DLX_IFinst__n0003<20>_G  (
    .ADR0(DLX_IFinst_IR_previous[20]),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(IR[20]),
    .ADR3(VCC),
    .O(N127676)
  );
  defparam \DLX_IFinst__n0003<20>_F .INIT = 16'hAEA2;
  X_LUT4 \DLX_IFinst__n0003<20>_F  (
    .ADR0(IR[20]),
    .ADR1(DLX_IFinst_stalled),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(DLX_IFinst_IR_curr[20]),
    .O(N127674)
  );
  defparam vga_top_vga1_hsyncout_136.INIT = 1'b1;
  X_SFF vga_top_vga1_hsyncout_136 (
    .I(\hsync/LOGIC_ZERO ),
    .CE(VCC),
    .CLK(clkdiv_vga),
    .SET(GSR),
    .RST(GND),
    .SSET(vga_top_vga1__n0010),
    .SRST(GND),
    .O(vga_top_vga1_hsyncout)
  );
  X_MUX2 DLX_RF_delay_inst_Mmux_outp_inst_mux_f5_2111 (
    .IA(N127994),
    .IB(N127996),
    .SEL(delay_selectRF_0_IBUF),
    .O(\DLX_clk_IF_del/F5MUX )
  );
  defparam DLX_RF_delay_inst_Mmux_outp_inst_mux_f5_2111_G.INIT = 16'hFC30;
  X_LUT4 DLX_RF_delay_inst_Mmux_outp_inst_mux_f5_2111_G (
    .ADR0(VCC),
    .ADR1(delay_selectRF_1_IBUF),
    .ADR2(DLX_RF_delay_inst_wint20),
    .ADR3(DLX_RF_delay_inst_wint30),
    .O(N127996)
  );
  defparam DLX_RF_delay_inst_Mmux_outp_inst_mux_f5_2111_F.INIT = 16'hFA0A;
  X_LUT4 DLX_RF_delay_inst_Mmux_outp_inst_mux_f5_2111_F (
    .ADR0(DLX_RF_delay_inst_wint14),
    .ADR1(VCC),
    .ADR2(delay_selectRF_1_IBUF),
    .ADR3(DLX_RF_delay_inst_wint24),
    .O(N127994)
  );
  X_BUF \DLX_clk_IF_del/XUSED  (
    .I(\DLX_clk_IF_del/F5MUX ),
    .O(DLX_clk_IF_del)
  );
  X_MUX2 \DLX_IFinst__n0003<13>  (
    .IA(N127754),
    .IB(N127756),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[13])
  );
  defparam \DLX_IFinst__n0003<13>_G .INIT = 16'hEE22;
  X_LUT4 \DLX_IFinst__n0003<13>_G  (
    .ADR0(DLX_IFinst_IR_previous[13]),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(VCC),
    .ADR3(IR[13]),
    .O(N127756)
  );
  defparam \DLX_IFinst__n0003<13>_F .INIT = 16'hB8AA;
  X_LUT4 \DLX_IFinst__n0003<13>_F  (
    .ADR0(IR[13]),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(DLX_IFinst_IR_curr[13]),
    .ADR3(DLX_IFinst_stalled),
    .O(N127754)
  );
  X_MUX2 \DLX_IFinst__n0003<21>  (
    .IA(N127664),
    .IB(N127666),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[21])
  );
  defparam \DLX_IFinst__n0003<21>_G .INIT = 16'hCFC0;
  X_LUT4 \DLX_IFinst__n0003<21>_G  (
    .ADR0(VCC),
    .ADR1(IR[21]),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(DLX_IFinst_IR_previous[21]),
    .O(N127666)
  );
  defparam \DLX_IFinst__n0003<21>_F .INIT = 16'hCCAC;
  X_LUT4 \DLX_IFinst__n0003<21>_F  (
    .ADR0(DLX_IFinst_IR_curr[21]),
    .ADR1(IR[21]),
    .ADR2(DLX_IFinst_stalled),
    .ADR3(DLX_IDinst_branch_sig),
    .O(N127664)
  );
  X_MUX2 \DLX_IFinst__n0003<14>  (
    .IA(N128099),
    .IB(N128101),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[14])
  );
  defparam \DLX_IFinst__n0003<14>_G .INIT = 16'hEE22;
  X_LUT4 \DLX_IFinst__n0003<14>_G  (
    .ADR0(DLX_IFinst_IR_previous[14]),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(VCC),
    .ADR3(IR[14]),
    .O(N128101)
  );
  defparam \DLX_IFinst__n0003<14>_F .INIT = 16'hEF20;
  X_LUT4 \DLX_IFinst__n0003<14>_F  (
    .ADR0(DLX_IFinst_IR_curr[14]),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(DLX_IFinst_stalled),
    .ADR3(IR[14]),
    .O(N128099)
  );
  X_MUX2 \DLX_IFinst__n0003<30>  (
    .IA(N127839),
    .IB(N127841),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[30])
  );
  defparam \DLX_IFinst__n0003<30>_G .INIT = 16'hF5A0;
  X_LUT4 \DLX_IFinst__n0003<30>_G  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(VCC),
    .ADR2(IR_MSB_6_OBUF),
    .ADR3(DLX_IFinst_IR_previous[30]),
    .O(N127841)
  );
  defparam \DLX_IFinst__n0003<30>_F .INIT = 16'hE4F0;
  X_LUT4 \DLX_IFinst__n0003<30>_F  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(DLX_IFinst_IR_curr[30]),
    .ADR2(IR_MSB_6_OBUF),
    .ADR3(DLX_IFinst_stalled),
    .O(N127839)
  );
  X_MUX2 \DLX_IFinst__n0003<22>  (
    .IA(N127704),
    .IB(N127706),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[22])
  );
  defparam \DLX_IFinst__n0003<22>_G .INIT = 16'hFA0A;
  X_LUT4 \DLX_IFinst__n0003<22>_G  (
    .ADR0(DLX_IFinst_IR_previous[22]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(IR[22]),
    .O(N127706)
  );
  defparam \DLX_IFinst__n0003<22>_F .INIT = 16'hF0D8;
  X_LUT4 \DLX_IFinst__n0003<22>_F  (
    .ADR0(DLX_IFinst_stalled),
    .ADR1(DLX_IFinst_IR_curr[22]),
    .ADR2(IR[22]),
    .ADR3(DLX_IDinst_branch_sig),
    .O(N127704)
  );
  X_MUX2 \DLX_IFinst__n0003<23>  (
    .IA(N127859),
    .IB(N127861),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[23])
  );
  defparam \DLX_IFinst__n0003<23>_G .INIT = 16'hDD88;
  X_LUT4 \DLX_IFinst__n0003<23>_G  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(IR[23]),
    .ADR2(VCC),
    .ADR3(DLX_IFinst_IR_previous[23]),
    .O(N127861)
  );
  defparam \DLX_IFinst__n0003<23>_F .INIT = 16'hCACC;
  X_LUT4 \DLX_IFinst__n0003<23>_F  (
    .ADR0(DLX_IFinst_IR_curr[23]),
    .ADR1(IR[23]),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(DLX_IFinst_stalled),
    .O(N127859)
  );
  X_MUX2 \DLX_IFinst__n0003<31>  (
    .IA(N127849),
    .IB(N127851),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[31])
  );
  defparam \DLX_IFinst__n0003<31>_G .INIT = 16'hCCAA;
  X_LUT4 \DLX_IFinst__n0003<31>_G  (
    .ADR0(DLX_IFinst_IR_previous[31]),
    .ADR1(IR_MSB_7_OBUF),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_branch_sig),
    .O(N127851)
  );
  defparam \DLX_IFinst__n0003<31>_F .INIT = 16'hCCAC;
  X_LUT4 \DLX_IFinst__n0003<31>_F  (
    .ADR0(DLX_IFinst_IR_curr[31]),
    .ADR1(IR_MSB_7_OBUF),
    .ADR2(DLX_IFinst_stalled),
    .ADR3(DLX_IDinst_branch_sig),
    .O(N127849)
  );
  X_MUX2 \DLX_IFinst__n0003<15>  (
    .IA(N127749),
    .IB(N127751),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[15])
  );
  defparam \DLX_IFinst__n0003<15>_G .INIT = 16'hBB88;
  X_LUT4 \DLX_IFinst__n0003<15>_G  (
    .ADR0(IR[15]),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(VCC),
    .ADR3(DLX_IFinst_IR_previous[15]),
    .O(N127751)
  );
  defparam \DLX_IFinst__n0003<15>_F .INIT = 16'hE2F0;
  X_LUT4 \DLX_IFinst__n0003<15>_F  (
    .ADR0(DLX_IFinst_IR_curr[15]),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(IR[15]),
    .ADR3(DLX_IFinst_stalled),
    .O(N127749)
  );
  X_MUX2 \DLX_EXinst_Mshift__n0025_Sh<40>  (
    .IA(N127919),
    .IB(N127921),
    .SEL(DLX_IDinst_reg_out_B_3_1),
    .O(\DLX_EXinst_Mshift__n0025_Sh<40>/F5MUX )
  );
  defparam \DLX_EXinst_Mshift__n0025_Sh<40>_G .INIT = 16'h0010;
  X_LUT4 \DLX_EXinst_Mshift__n0025_Sh<40>_G  (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(DLX_IDinst_reg_out_B[0]),
    .ADR2(DLX_IDinst_reg_out_A[0]),
    .ADR3(DLX_IDinst_reg_out_B_2_1),
    .O(N127921)
  );
  defparam \DLX_EXinst_Mshift__n0025_Sh<40>_F .INIT = 16'hFCAA;
  X_LUT4 \DLX_EXinst_Mshift__n0025_Sh<40>_F  (
    .ADR0(\DLX_EXinst_Mshift__n0025_Sh[8] ),
    .ADR1(CHOICE1084),
    .ADR2(CHOICE1078),
    .ADR3(DLX_IDinst_reg_out_B_2_1),
    .O(N127919)
  );
  X_BUF \DLX_EXinst_Mshift__n0025_Sh<40>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0025_Sh<40>/F5MUX ),
    .O(\DLX_EXinst_Mshift__n0025_Sh[40] )
  );
  X_MUX2 \DLX_IFinst__n0003<16>  (
    .IA(N128059),
    .IB(N128061),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[16])
  );
  defparam \DLX_IFinst__n0003<16>_G .INIT = 16'hE2E2;
  X_LUT4 \DLX_IFinst__n0003<16>_G  (
    .ADR0(DLX_IFinst_IR_previous[16]),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(IR[16]),
    .ADR3(VCC),
    .O(N128061)
  );
  defparam \DLX_IFinst__n0003<16>_F .INIT = 16'hF4B0;
  X_LUT4 \DLX_IFinst__n0003<16>_F  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(DLX_IFinst_stalled),
    .ADR2(IR[16]),
    .ADR3(DLX_IFinst_IR_curr[16]),
    .O(N128059)
  );
  X_MUX2 \DLX_IFinst__n0003<24>  (
    .IA(N127739),
    .IB(N127741),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[24])
  );
  defparam \DLX_IFinst__n0003<24>_G .INIT = 16'hFC30;
  X_LUT4 \DLX_IFinst__n0003<24>_G  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(DLX_IFinst_IR_previous[24]),
    .ADR3(IR_MSB_0_OBUF),
    .O(N127741)
  );
  defparam \DLX_IFinst__n0003<24>_F .INIT = 16'hD8CC;
  X_LUT4 \DLX_IFinst__n0003<24>_F  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(IR_MSB_0_OBUF),
    .ADR2(DLX_IFinst_IR_curr[24]),
    .ADR3(DLX_IFinst_stalled),
    .O(N127739)
  );
  X_MUX2 \DLX_IFinst__n0003<25>  (
    .IA(N127969),
    .IB(N127971),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[25])
  );
  defparam \DLX_IFinst__n0003<25>_G .INIT = 16'hCFC0;
  X_LUT4 \DLX_IFinst__n0003<25>_G  (
    .ADR0(VCC),
    .ADR1(IR_MSB_1_OBUF),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(DLX_IFinst_IR_previous[25]),
    .O(N127971)
  );
  defparam \DLX_IFinst__n0003<25>_F .INIT = 16'hCACC;
  X_LUT4 \DLX_IFinst__n0003<25>_F  (
    .ADR0(DLX_IFinst_IR_curr[25]),
    .ADR1(IR_MSB_1_OBUF),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(DLX_IFinst_stalled),
    .O(N127969)
  );
  X_MUX2 \DLX_IFinst__n0003<17>  (
    .IA(N127629),
    .IB(N127631),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[17])
  );
  defparam \DLX_IFinst__n0003<17>_G .INIT = 16'hBB88;
  X_LUT4 \DLX_IFinst__n0003<17>_G  (
    .ADR0(IR[17]),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(VCC),
    .ADR3(DLX_IFinst_IR_previous[17]),
    .O(N127631)
  );
  defparam \DLX_IFinst__n0003<17>_F .INIT = 16'hFD08;
  X_LUT4 \DLX_IFinst__n0003<17>_F  (
    .ADR0(DLX_IFinst_stalled),
    .ADR1(DLX_IFinst_IR_curr[17]),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(IR[17]),
    .O(N127629)
  );
  X_MUX2 \DLX_IFinst__n0003<26>  (
    .IA(N127734),
    .IB(N127736),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[26])
  );
  defparam \DLX_IFinst__n0003<26>_G .INIT = 16'hE2E2;
  X_LUT4 \DLX_IFinst__n0003<26>_G  (
    .ADR0(DLX_IFinst_IR_previous[26]),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(IR_MSB_2_OBUF),
    .ADR3(VCC),
    .O(N127736)
  );
  defparam \DLX_IFinst__n0003<26>_F .INIT = 16'hDC8C;
  X_LUT4 \DLX_IFinst__n0003<26>_F  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(IR_MSB_2_OBUF),
    .ADR2(DLX_IFinst_stalled),
    .ADR3(DLX_IFinst_IR_curr[26]),
    .O(N127734)
  );
  X_MUX2 \DLX_IFinst__n0003<18>  (
    .IA(N127609),
    .IB(N127611),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[18])
  );
  defparam \DLX_IFinst__n0003<18>_G .INIT = 16'hBB88;
  X_LUT4 \DLX_IFinst__n0003<18>_G  (
    .ADR0(IR[18]),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(VCC),
    .ADR3(DLX_IFinst_IR_previous[18]),
    .O(N127611)
  );
  defparam \DLX_IFinst__n0003<18>_F .INIT = 16'hF0B8;
  X_LUT4 \DLX_IFinst__n0003<18>_F  (
    .ADR0(DLX_IFinst_IR_curr[18]),
    .ADR1(DLX_IFinst_stalled),
    .ADR2(IR[18]),
    .ADR3(DLX_IDinst_branch_sig),
    .O(N127609)
  );
  X_MUX2 \DLX_EXinst_Mshift__n0025_Sh<43>  (
    .IA(N127989),
    .IB(N127991),
    .SEL(DLX_IDinst_reg_out_B_2_1),
    .O(\DLX_EXinst_Mshift__n0025_Sh<43>/F5MUX )
  );
  defparam \DLX_EXinst_Mshift__n0025_Sh<43>_G .INIT = 16'h3120;
  X_LUT4 \DLX_EXinst_Mshift__n0025_Sh<43>_G  (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(DLX_IDinst_reg_out_B_3_1),
    .ADR2(N94305),
    .ADR3(DLX_EXinst_N62851),
    .O(N127991)
  );
  defparam \DLX_EXinst_Mshift__n0025_Sh<43>_F .INIT = 16'hFACA;
  X_LUT4 \DLX_EXinst_Mshift__n0025_Sh<43>_F  (
    .ADR0(\DLX_EXinst_Mshift__n0025_Sh[11] ),
    .ADR1(CHOICE1054),
    .ADR2(DLX_IDinst_reg_out_B_3_1),
    .ADR3(CHOICE1060),
    .O(N127989)
  );
  X_BUF \DLX_EXinst_Mshift__n0025_Sh<43>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0025_Sh<43>/F5MUX ),
    .O(\DLX_EXinst_Mshift__n0025_Sh[43] )
  );
  X_MUX2 \DLX_IFinst__n0003<27>  (
    .IA(N127809),
    .IB(N127811),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[27])
  );
  defparam \DLX_IFinst__n0003<27>_G .INIT = 16'hE2E2;
  X_LUT4 \DLX_IFinst__n0003<27>_G  (
    .ADR0(DLX_IFinst_IR_previous[27]),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(IR_MSB_3_OBUF),
    .ADR3(VCC),
    .O(N127811)
  );
  defparam \DLX_IFinst__n0003<27>_F .INIT = 16'hBA8A;
  X_LUT4 \DLX_IFinst__n0003<27>_F  (
    .ADR0(IR_MSB_3_OBUF),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(DLX_IFinst_stalled),
    .ADR3(DLX_IFinst_IR_curr[27]),
    .O(N127809)
  );
  X_MUX2 \DLX_IFinst__n0003<19>  (
    .IA(N127649),
    .IB(N127651),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[19])
  );
  defparam \DLX_IFinst__n0003<19>_G .INIT = 16'hFA0A;
  X_LUT4 \DLX_IFinst__n0003<19>_G  (
    .ADR0(DLX_IFinst_IR_previous[19]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(IR[19]),
    .O(N127651)
  );
  defparam \DLX_IFinst__n0003<19>_F .INIT = 16'hE2F0;
  X_LUT4 \DLX_IFinst__n0003<19>_F  (
    .ADR0(DLX_IFinst_IR_curr[19]),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(IR[19]),
    .ADR3(DLX_IFinst_stalled),
    .O(N127649)
  );
  X_MUX2 \DLX_IFinst__n0003<28>  (
    .IA(N127914),
    .IB(N127916),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[28])
  );
  defparam \DLX_IFinst__n0003<28>_G .INIT = 16'hEE44;
  X_LUT4 \DLX_IFinst__n0003<28>_G  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(DLX_IFinst_IR_previous[28]),
    .ADR2(VCC),
    .ADR3(IR_MSB_4_OBUF),
    .O(N127916)
  );
  defparam \DLX_IFinst__n0003<28>_F .INIT = 16'hF2D0;
  X_LUT4 \DLX_IFinst__n0003<28>_F  (
    .ADR0(DLX_IFinst_stalled),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(IR_MSB_4_OBUF),
    .ADR3(DLX_IFinst_IR_curr[28]),
    .O(N127914)
  );
  X_MUX2 \DLX_IFinst__n0003<29>  (
    .IA(N127834),
    .IB(N127836),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[29])
  );
  defparam \DLX_IFinst__n0003<29>_G .INIT = 16'hCCF0;
  X_LUT4 \DLX_IFinst__n0003<29>_G  (
    .ADR0(VCC),
    .ADR1(IR_MSB_5_OBUF),
    .ADR2(DLX_IFinst_IR_previous[29]),
    .ADR3(DLX_IDinst_branch_sig),
    .O(N127836)
  );
  defparam \DLX_IFinst__n0003<29>_F .INIT = 16'hCACC;
  X_LUT4 \DLX_IFinst__n0003<29>_F  (
    .ADR0(DLX_IFinst_IR_curr[29]),
    .ADR1(IR_MSB_5_OBUF),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(DLX_IFinst_stalled),
    .O(N127834)
  );
  X_MUX2 \DLX_EXinst__n0006<30>99_SW0  (
    .IA(N128084),
    .IB(N128086),
    .SEL(DLX_IDinst_IR_function_field[4]),
    .O(\N126560/F5MUX )
  );
  defparam \DLX_EXinst__n0006<30>99_SW0_G .INIT = 16'h88C0;
  X_LUT4 \DLX_EXinst__n0006<30>99_SW0_G  (
    .ADR0(DLX_EXinst_N62826),
    .ADR1(DLX_EXinst_N66202),
    .ADR2(N93331),
    .ADR3(DLX_IDinst_IR_function_field[3]),
    .O(N128086)
  );
  defparam \DLX_EXinst__n0006<30>99_SW0_F .INIT = 16'hB080;
  X_LUT4 \DLX_EXinst__n0006<30>99_SW0_F  (
    .ADR0(N98032),
    .ADR1(DLX_IDinst_IR_function_field[2]),
    .ADR2(DLX_EXinst_N66202),
    .ADR3(CHOICE5264),
    .O(N128084)
  );
  X_BUF \N126560/XUSED  (
    .I(\N126560/F5MUX ),
    .O(N126560)
  );
  X_MUX2 \DLX_EXinst__n0006<0>119  (
    .IA(N127789),
    .IB(N127791),
    .SEL(DLX_IDinst_reg_out_B[4]),
    .O(\CHOICE5871/F5MUX )
  );
  defparam \DLX_EXinst__n0006<0>119_G .INIT = 16'hC480;
  X_LUT4 \DLX_EXinst__n0006<0>119_G  (
    .ADR0(DLX_IDinst_reg_out_B[2]),
    .ADR1(DLX_EXinst_N62631),
    .ADR2(DLX_EXinst_N62727),
    .ADR3(DLX_EXinst_N64319),
    .O(N127791)
  );
  defparam \DLX_EXinst__n0006<0>119_F .INIT = 16'hE0C0;
  X_LUT4 \DLX_EXinst__n0006<0>119_F  (
    .ADR0(N96153),
    .ADR1(CHOICE5866),
    .ADR2(DLX_EXinst_N62631),
    .ADR3(DLX_IDinst_reg_out_B[2]),
    .O(N127789)
  );
  X_BUF \CHOICE5871/XUSED  (
    .I(\CHOICE5871/F5MUX ),
    .O(CHOICE5871)
  );
  X_MUX2 \DLX_EXinst__n0006<16>16  (
    .IA(N128044),
    .IB(N128046),
    .SEL(DLX_IDinst_IR_function_field[4]),
    .O(\CHOICE5100/F5MUX )
  );
  defparam \DLX_EXinst__n0006<16>16_G .INIT = 16'h3000;
  X_LUT4 \DLX_EXinst__n0006<16>16_G  (
    .ADR0(VCC),
    .ADR1(\DLX_IDinst_Imm[5] ),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(N110065),
    .O(N128046)
  );
  defparam \DLX_EXinst__n0006<16>16_F .INIT = 16'hA808;
  X_LUT4 \DLX_EXinst__n0006<16>16_F  (
    .ADR0(DLX_EXinst_N63185),
    .ADR1(DLX_EXinst_N64565),
    .ADR2(DLX_IDinst_IR_function_field[2]),
    .ADR3(DLX_EXinst_N62715),
    .O(N128044)
  );
  X_BUF \CHOICE5100/XUSED  (
    .I(\CHOICE5100/F5MUX ),
    .O(CHOICE5100)
  );
  X_MUX2 \DLX_EXinst__n0006<16>90  (
    .IA(N127719),
    .IB(N127721),
    .SEL(DLX_IDinst_IR_function_field[2]),
    .O(\CHOICE5125/F5MUX )
  );
  defparam \DLX_EXinst__n0006<16>90_G .INIT = 16'h0D08;
  X_LUT4 \DLX_EXinst__n0006<16>90_G  (
    .ADR0(DLX_IDinst_IR_function_field[3]),
    .ADR1(\DLX_EXinst_Mshift__n0027_Sh[4] ),
    .ADR2(DLX_IDinst_IR_function_field[4]),
    .ADR3(\DLX_EXinst_Mshift__n0027_Sh[12] ),
    .O(N127721)
  );
  defparam \DLX_EXinst__n0006<16>90_F .INIT = 16'h3120;
  X_LUT4 \DLX_EXinst__n0006<16>90_F  (
    .ADR0(DLX_IDinst_IR_function_field[3]),
    .ADR1(DLX_IDinst_IR_function_field[4]),
    .ADR2(\DLX_EXinst_Mshift__n0027_Sh[8] ),
    .ADR3(N93179),
    .O(N127719)
  );
  X_BUF \CHOICE5125/XUSED  (
    .I(\CHOICE5125/F5MUX ),
    .O(CHOICE5125)
  );
  X_MUX2 \DLX_EXinst__n0006<17>74  (
    .IA(N127864),
    .IB(N127866),
    .SEL(DLX_IDinst_IR_function_field[3]),
    .O(\CHOICE5598/F5MUX )
  );
  defparam \DLX_EXinst__n0006<17>74_G .INIT = 16'hCA00;
  X_LUT4 \DLX_EXinst__n0006<17>74_G  (
    .ADR0(\DLX_EXinst_Mshift__n0027_Sh[9] ),
    .ADR1(\DLX_EXinst_Mshift__n0027_Sh[5] ),
    .ADR2(DLX_IDinst_IR_function_field[2]),
    .ADR3(DLX_EXinst__n0081),
    .O(N127866)
  );
  defparam \DLX_EXinst__n0006<17>74_F .INIT = 16'h88C0;
  X_LUT4 \DLX_EXinst__n0006<17>74_F  (
    .ADR0(\DLX_EXinst_Mshift__n0027_Sh[13] ),
    .ADR1(DLX_EXinst__n0081),
    .ADR2(N93127),
    .ADR3(DLX_IDinst_IR_function_field[2]),
    .O(N127864)
  );
  X_BUF \CHOICE5598/XUSED  (
    .I(\CHOICE5598/F5MUX ),
    .O(CHOICE5598)
  );
  X_MUX2 \DLX_EXinst__n0006<0>619  (
    .IA(N127894),
    .IB(N127896),
    .SEL(DLX_IDinst_IR_function_field[2]),
    .O(\CHOICE5973/F5MUX )
  );
  defparam \DLX_EXinst__n0006<0>619_G .INIT = 16'hEE00;
  X_LUT4 \DLX_EXinst__n0006<0>619_G  (
    .ADR0(CHOICE1276),
    .ADR1(CHOICE1270),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N63185),
    .O(N127896)
  );
  defparam \DLX_EXinst__n0006<0>619_F .INIT = 16'hA888;
  X_LUT4 \DLX_EXinst__n0006<0>619_F  (
    .ADR0(DLX_EXinst_N63185),
    .ADR1(CHOICE5969),
    .ADR2(\DLX_EXinst_Mshift__n0028_Sh[8] ),
    .ADR3(DLX_IDinst_IR_function_field[3]),
    .O(N127894)
  );
  X_BUF \CHOICE5973/XUSED  (
    .I(\CHOICE5973/F5MUX ),
    .O(CHOICE5973)
  );
  X_MUX2 DLX_EXinst_Ker6505418 (
    .IA(N127654),
    .IB(N127656),
    .SEL(DLX_EXinst__n0030_1),
    .O(\CHOICE1771/F5MUX )
  );
  defparam DLX_EXinst_Ker6505418_G.INIT = 16'h0808;
  X_LUT4 DLX_EXinst_Ker6505418_G (
    .ADR0(N111221),
    .ADR1(DLX_IDinst_reg_out_B[4]),
    .ADR2(DLX_IDinst_reg_out_B[5]),
    .ADR3(VCC),
    .O(N127656)
  );
  defparam DLX_EXinst_Ker6505418_F.INIT = 16'h3000;
  X_LUT4 DLX_EXinst_Ker6505418_F (
    .ADR0(VCC),
    .ADR1(\DLX_IDinst_Imm[5] ),
    .ADR2(N110065),
    .ADR3(DLX_IDinst_IR_function_field[4]),
    .O(N127654)
  );
  X_BUF \CHOICE1771/XUSED  (
    .I(\CHOICE1771/F5MUX ),
    .O(CHOICE1771)
  );
  X_MUX2 \DLX_EXinst__n0006<1>254  (
    .IA(N127764),
    .IB(N127766),
    .SEL(DLX_IDinst_reg_out_B[4]),
    .O(\CHOICE5709/F5MUX )
  );
  defparam \DLX_EXinst__n0006<1>254_G .INIT = 16'hCC80;
  X_LUT4 \DLX_EXinst__n0006<1>254_G  (
    .ADR0(DLX_IDinst_reg_out_B[5]),
    .ADR1(N111221),
    .ADR2(CHOICE1919),
    .ADR3(CHOICE1926),
    .O(N127766)
  );
  defparam \DLX_EXinst__n0006<1>254_F .INIT = 16'hE0E0;
  X_LUT4 \DLX_EXinst__n0006<1>254_F  (
    .ADR0(CHOICE5706),
    .ADR1(CHOICE5696),
    .ADR2(DLX_EXinst_N62631),
    .ADR3(VCC),
    .O(N127764)
  );
  X_BUF \CHOICE5709/XUSED  (
    .I(\CHOICE5709/F5MUX ),
    .O(CHOICE5709)
  );
  X_MUX2 \DLX_EXinst__n0006<18>74  (
    .IA(N127824),
    .IB(N127826),
    .SEL(DLX_IDinst_IR_function_field[3]),
    .O(\CHOICE5432/F5MUX )
  );
  defparam \DLX_EXinst__n0006<18>74_G .INIT = 16'hC808;
  X_LUT4 \DLX_EXinst__n0006<18>74_G  (
    .ADR0(\DLX_EXinst_Mshift__n0027_Sh[10] ),
    .ADR1(DLX_EXinst__n0081),
    .ADR2(DLX_IDinst_IR_function_field[2]),
    .ADR3(\DLX_EXinst_Mshift__n0027_Sh[6] ),
    .O(N127826)
  );
  defparam \DLX_EXinst__n0006<18>74_F .INIT = 16'hA808;
  X_LUT4 \DLX_EXinst__n0006<18>74_F  (
    .ADR0(DLX_EXinst__n0081),
    .ADR1(N93229),
    .ADR2(DLX_IDinst_IR_function_field[2]),
    .ADR3(\DLX_EXinst_Mshift__n0027_Sh[14] ),
    .O(N127824)
  );
  X_BUF \CHOICE5432/XUSED  (
    .I(\CHOICE5432/F5MUX ),
    .O(CHOICE5432)
  );
  X_MUX2 \DLX_EXinst__n0006<2>217  (
    .IA(N128009),
    .IB(N128011),
    .SEL(DLX_IDinst_reg_out_B[0]),
    .O(\CHOICE5540/F5MUX )
  );
  defparam \DLX_EXinst__n0006<2>217_G .INIT = 16'h2320;
  X_LUT4 \DLX_EXinst__n0006<2>217_G  (
    .ADR0(DLX_EXinst_N63036),
    .ADR1(DLX_IDinst_reg_out_B[2]),
    .ADR2(DLX_IDinst_reg_out_B[3]),
    .ADR3(DLX_EXinst_N64904),
    .O(N128011)
  );
  defparam \DLX_EXinst__n0006<2>217_F .INIT = 16'h3022;
  X_LUT4 \DLX_EXinst__n0006<2>217_F  (
    .ADR0(DLX_EXinst_N64255),
    .ADR1(DLX_IDinst_reg_out_B[2]),
    .ADR2(DLX_EXinst_N63329),
    .ADR3(DLX_IDinst_reg_out_B[3]),
    .O(N128009)
  );
  X_BUF \CHOICE5540/XUSED  (
    .I(\CHOICE5540/F5MUX ),
    .O(CHOICE5540)
  );
  X_MUX2 \DLX_EXinst__n0006<19>74  (
    .IA(N128069),
    .IB(N128071),
    .SEL(DLX_IDinst_IR_function_field[3]),
    .O(\CHOICE4965/F5MUX )
  );
  defparam \DLX_EXinst__n0006<19>74_G .INIT = 16'hE020;
  X_LUT4 \DLX_EXinst__n0006<19>74_G  (
    .ADR0(\DLX_EXinst_Mshift__n0027_Sh[11] ),
    .ADR1(DLX_IDinst_IR_function_field[2]),
    .ADR2(DLX_EXinst__n0081),
    .ADR3(\DLX_EXinst_Mshift__n0027_Sh[7] ),
    .O(N128071)
  );
  defparam \DLX_EXinst__n0006<19>74_F .INIT = 16'hC0A0;
  X_LUT4 \DLX_EXinst__n0006<19>74_F  (
    .ADR0(\DLX_EXinst_Mshift__n0027_Sh[19] ),
    .ADR1(\DLX_EXinst_Mshift__n0027_Sh[15] ),
    .ADR2(DLX_EXinst__n0081),
    .ADR3(DLX_IDinst_IR_function_field[2]),
    .O(N128069)
  );
  X_BUF \CHOICE4965/XUSED  (
    .I(\CHOICE4965/F5MUX ),
    .O(CHOICE4965)
  );
  X_MUX2 DLX_EXinst_Ker6512856 (
    .IA(N128019),
    .IB(N128021),
    .SEL(\DLX_IDinst_Imm[5] ),
    .O(\N101537/F5MUX )
  );
  defparam DLX_EXinst_Ker6512856_G.INIT = 16'h70F0;
  X_LUT4 DLX_EXinst_Ker6512856_G (
    .ADR0(DLX_EXinst_N63129),
    .ADR1(DLX_IDinst_IR_function_field_2_1),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(DLX_IDinst_IR_function_field_3_1),
    .O(N128021)
  );
  defparam DLX_EXinst_Ker6512856_F.INIT = 16'hFFC0;
  X_LUT4 DLX_EXinst_Ker6512856_F (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N66421),
    .ADR2(DLX_IDinst_IR_function_field_2_1),
    .ADR3(N125971),
    .O(N128019)
  );
  X_BUF \N101537/XUSED  (
    .I(\N101537/F5MUX ),
    .O(N101537)
  );
  X_MUX2 DLX_EXinst_Ker6508317 (
    .IA(N127724),
    .IB(N127726),
    .SEL(DLX_IDinst_reg_out_B[5]),
    .O(\N95810/F5MUX )
  );
  defparam DLX_EXinst_Ker6508317_G.INIT = 16'h0030;
  X_LUT4 DLX_EXinst_Ker6508317_G (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_B_2_1),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(DLX_IDinst_reg_out_B_3_1),
    .O(N127726)
  );
  defparam DLX_EXinst_Ker6508317_F.INIT = 16'hFAAA;
  X_LUT4 DLX_EXinst_Ker6508317_F (
    .ADR0(\DLX_EXinst_Mshift__n0026_Sh[60] ),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(DLX_EXinst_N62740),
    .O(N127724)
  );
  X_BUF \N95810/XUSED  (
    .I(\N95810/F5MUX ),
    .O(N95810)
  );
  X_MUX2 DLX_EXinst_Ker6513856 (
    .IA(N128034),
    .IB(N128036),
    .SEL(DLX_IDinst_reg_out_B[5]),
    .O(\CHOICE2965/F5MUX )
  );
  defparam DLX_EXinst_Ker6513856_G.INIT = 16'h70F0;
  X_LUT4 DLX_EXinst_Ker6513856_G (
    .ADR0(DLX_IDinst_reg_out_B_2_1),
    .ADR1(DLX_IDinst_reg_out_B_3_1),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(DLX_EXinst_N63157),
    .O(N128036)
  );
  defparam DLX_EXinst_Ker6513856_F.INIT = 16'hECEC;
  X_LUT4 DLX_EXinst_Ker6513856_F (
    .ADR0(DLX_EXinst_N66431),
    .ADR1(N126006),
    .ADR2(DLX_IDinst_reg_out_B_2_1),
    .ADR3(VCC),
    .O(N128034)
  );
  X_BUF \CHOICE2965/XUSED  (
    .I(\CHOICE2965/F5MUX ),
    .O(CHOICE2965)
  );
  X_MUX2 DLX_EXinst_Ker6514860 (
    .IA(N127619),
    .IB(N127621),
    .SEL(\DLX_IDinst_Imm[5] ),
    .O(\CHOICE3097/F5MUX )
  );
  defparam DLX_EXinst_Ker6514860_G.INIT = 16'h30AA;
  X_LUT4 DLX_EXinst_Ker6514860_G (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(DLX_IDinst_IR_function_field_2_1),
    .ADR2(\DLX_EXinst_Mshift__n0024_Sh[61] ),
    .ADR3(DLX_IDinst_IR_function_field_3_1),
    .O(N127621)
  );
  defparam DLX_EXinst_Ker6514860_F.INIT = 16'hAAFA;
  X_LUT4 DLX_EXinst_Ker6514860_F (
    .ADR0(CHOICE3085),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N62936),
    .ADR3(DLX_IDinst_IR_function_field_2_1),
    .O(N127619)
  );
  X_BUF \CHOICE3097/XUSED  (
    .I(\CHOICE3097/F5MUX ),
    .O(CHOICE3097)
  );
  X_MUX2 DLX_EXinst_Ker6517328 (
    .IA(N128054),
    .IB(N128056),
    .SEL(DLX_IDinst_reg_out_B[0]),
    .O(\N97089/F5MUX )
  );
  defparam DLX_EXinst_Ker6517328_G.INIT = 16'hEEAA;
  X_LUT4 DLX_EXinst_Ker6517328_G (
    .ADR0(CHOICE1184),
    .ADR1(DLX_EXinst_N63374),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B_3_1),
    .O(N128056)
  );
  defparam DLX_EXinst_Ker6517328_F.INIT = 16'hF0CC;
  X_LUT4 DLX_EXinst_Ker6517328_F (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N62896),
    .ADR2(DLX_EXinst_N62876),
    .ADR3(DLX_IDinst_reg_out_B_3_1),
    .O(N128054)
  );
  X_BUF \N97089/XUSED  (
    .I(\N97089/F5MUX ),
    .O(N97089)
  );
  X_MUX2 DLX_EXinst_Ker6453328 (
    .IA(N127799),
    .IB(N127801),
    .SEL(DLX_IDinst_reg_out_B_3_1),
    .O(\N97449/F5MUX )
  );
  defparam DLX_EXinst_Ker6453328_G.INIT = 16'hAFA0;
  X_LUT4 DLX_EXinst_Ker6453328_G (
    .ADR0(DLX_EXinst_N63780),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[0]),
    .ADR3(DLX_EXinst_N63066),
    .O(N127801)
  );
  defparam DLX_EXinst_Ker6453328_F.INIT = 16'hFA50;
  X_LUT4 DLX_EXinst_Ker6453328_F (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N63046),
    .ADR3(DLX_EXinst_N63419),
    .O(N127799)
  );
  X_BUF \N97449/XUSED  (
    .I(\N97449/F5MUX ),
    .O(N97449)
  );
  X_MUX2 DLX_EXinst_Ker6435737 (
    .IA(N127614),
    .IB(N127616),
    .SEL(DLX_IDinst_reg_out_B[0]),
    .O(\N100843/F5MUX )
  );
  defparam DLX_EXinst_Ker6435737_G.INIT = 16'hBBB8;
  X_LUT4 DLX_EXinst_Ker6435737_G (
    .ADR0(DLX_EXinst_N63379),
    .ADR1(DLX_IDinst_reg_out_B_3_1),
    .ADR2(CHOICE1825),
    .ADR3(DLX_EXinst_N63274),
    .O(N127616)
  );
  defparam DLX_EXinst_Ker6435737_F.INIT = 16'hE4E4;
  X_LUT4 DLX_EXinst_Ker6435737_F (
    .ADR0(DLX_IDinst_reg_out_B_3_1),
    .ADR1(CHOICE1825),
    .ADR2(DLX_EXinst_N62881),
    .ADR3(VCC),
    .O(N127614)
  );
  X_BUF \N100843/XUSED  (
    .I(\N100843/F5MUX ),
    .O(N100843)
  );
  X_MUX2 \DLX_EXinst__n0006<3>262  (
    .IA(N127854),
    .IB(N127856),
    .SEL(DLX_IDinst_reg_out_B[2]),
    .O(\CHOICE5077/F5MUX )
  );
  defparam \DLX_EXinst__n0006<3>262_G .INIT = 16'hCCC0;
  X_LUT4 \DLX_EXinst__n0006<3>262_G  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N62631),
    .ADR2(CHOICE1168),
    .ADR3(CHOICE1162),
    .O(N127856)
  );
  defparam \DLX_EXinst__n0006<3>262_F .INIT = 16'hEC00;
  X_LUT4 \DLX_EXinst__n0006<3>262_F  (
    .ADR0(DLX_IDinst_reg_out_B[3]),
    .ADR1(CHOICE5073),
    .ADR2(\DLX_EXinst_Mshift__n0026_Sh[11] ),
    .ADR3(DLX_EXinst_N62631),
    .O(N127854)
  );
  X_BUF \CHOICE5077/XUSED  (
    .I(\CHOICE5077/F5MUX ),
    .O(CHOICE5077)
  );
  X_MUX2 DLX_EXinst_Ker6455328 (
    .IA(N127759),
    .IB(N127761),
    .SEL(DLX_IDinst_IR_function_field[3]),
    .O(\N97305/F5MUX )
  );
  defparam DLX_EXinst_Ker6455328_G.INIT = 16'hDD88;
  X_LUT4 DLX_EXinst_Ker6455328_G (
    .ADR0(DLX_IDinst_IR_function_field[0]),
    .ADR1(DLX_EXinst_N63279),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N63016),
    .O(N127761)
  );
  defparam DLX_EXinst_Ker6455328_F.INIT = 16'hBB88;
  X_LUT4 DLX_EXinst_Ker6455328_F (
    .ADR0(DLX_EXinst_N63504),
    .ADR1(DLX_IDinst_IR_function_field[0]),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N62996),
    .O(N127759)
  );
  X_BUF \N97305/XUSED  (
    .I(\N97305/F5MUX ),
    .O(N97305)
  );
  X_MUX2 Mmux__COND_2_inst_mux_f5_0 (
    .IA(Mmux__COND_2__net0),
    .IB(Mmux__COND_2__net1),
    .SEL(vga_address[13]),
    .O(\Mmux__COND_2__net2/F5MUX )
  );
  defparam Mmux__COND_2_inst_lut3_11.INIT = 16'hBB88;
  X_LUT4 Mmux__COND_2_inst_lut3_11 (
    .ADR0(vram_out_vga[3]),
    .ADR1(vga_address[12]),
    .ADR2(VCC),
    .ADR3(vram_out_vga[2]),
    .O(Mmux__COND_2__net1)
  );
  defparam Mmux__COND_2_inst_lut3_01.INIT = 16'hAACC;
  X_LUT4 Mmux__COND_2_inst_lut3_01 (
    .ADR0(vram_out_vga[1]),
    .ADR1(vram_out_vga[0]),
    .ADR2(VCC),
    .ADR3(vga_address[12]),
    .O(Mmux__COND_2__net0)
  );
  X_BUF \Mmux__COND_2__net2/F5USED  (
    .I(\Mmux__COND_2__net2/F5MUX ),
    .O(Mmux__COND_2__net2)
  );
  X_MUX2 DLX_EXinst_Ker6453828 (
    .IA(N128074),
    .IB(N128076),
    .SEL(DLX_IDinst_reg_out_B_3_1),
    .O(\N97375/F5MUX )
  );
  defparam DLX_EXinst_Ker6453828_G.INIT = 16'hCCAA;
  X_LUT4 DLX_EXinst_Ker6453828_G (
    .ADR0(DLX_EXinst_N63429),
    .ADR1(DLX_EXinst_N63061),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[0]),
    .O(N128076)
  );
  defparam DLX_EXinst_Ker6453828_F.INIT = 16'hDD88;
  X_LUT4 DLX_EXinst_Ker6453828_F (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(DLX_EXinst_N63041),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N63409),
    .O(N128074)
  );
  X_BUF \N97375/XUSED  (
    .I(\N97375/F5MUX ),
    .O(N97375)
  );
  X_MUX2 DLX_EXinst_Ker6517828 (
    .IA(N127794),
    .IB(N127796),
    .SEL(DLX_IDinst_reg_out_B[0]),
    .O(\N97161/F5MUX )
  );
  defparam DLX_EXinst_Ker6517828_G.INIT = 16'hE4E4;
  X_LUT4 DLX_EXinst_Ker6517828_G (
    .ADR0(DLX_IDinst_reg_out_B_3_1),
    .ADR1(DLX_EXinst_N62891),
    .ADR2(DLX_EXinst_N62871),
    .ADR3(VCC),
    .O(N127796)
  );
  defparam DLX_EXinst_Ker6517828_F.INIT = 16'hFCF0;
  X_LUT4 DLX_EXinst_Ker6517828_F (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N63374),
    .ADR2(CHOICE1184),
    .ADR3(DLX_IDinst_reg_out_B_3_1),
    .O(N127794)
  );
  X_BUF \N97161/XUSED  (
    .I(\N97161/F5MUX ),
    .O(N97161)
  );
  X_MUX2 DLX_EXinst_Ker6458037 (
    .IA(N127949),
    .IB(N127951),
    .SEL(DLX_IDinst_IR_function_field[3]),
    .O(\N100919/F5MUX )
  );
  defparam DLX_EXinst_Ker6458037_G.INIT = 16'hACAC;
  X_LUT4 DLX_EXinst_Ker6458037_G (
    .ADR0(DLX_EXinst_N63459),
    .ADR1(DLX_EXinst_N62796),
    .ADR2(DLX_IDinst_IR_function_field[0]),
    .ADR3(VCC),
    .O(N127951)
  );
  defparam DLX_EXinst_Ker6458037_F.INIT = 16'hFFC0;
  X_LUT4 DLX_EXinst_Ker6458037_F (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_IR_function_field[0]),
    .ADR2(DLX_EXinst_N63309),
    .ADR3(CHOICE1838),
    .O(N127949)
  );
  X_BUF \N100919/XUSED  (
    .I(\N100919/F5MUX ),
    .O(N100919)
  );
  X_MUX2 DLX_EXinst_Ker6483236 (
    .IA(N128029),
    .IB(N128031),
    .SEL(DLX_IDinst_reg_out_B[5]),
    .O(\N101009/F5MUX )
  );
  defparam DLX_EXinst_Ker6483236_G.INIT = 16'h2AAA;
  X_LUT4 DLX_EXinst_Ker6483236_G (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(DLX_IDinst_reg_out_B_2_1),
    .ADR2(DLX_IDinst_reg_out_B_3_1),
    .ADR3(DLX_IDinst_reg_out_B[1]),
    .O(N128031)
  );
  defparam DLX_EXinst_Ker6483236_F.INIT = 16'hFC0C;
  X_LUT4 DLX_EXinst_Ker6483236_F (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N64334),
    .ADR2(DLX_IDinst_reg_out_B_2_1),
    .ADR3(DLX_EXinst_N62971),
    .O(N128029)
  );
  X_BUF \N101009/XUSED  (
    .I(\N101009/F5MUX ),
    .O(N101009)
  );
  X_MUX2 DLX_EXinst_Ker6483746 (
    .IA(N127869),
    .IB(N127871),
    .SEL(\DLX_IDinst_Imm[5] ),
    .O(\N101253/F5MUX )
  );
  defparam DLX_EXinst_Ker6483746_G.INIT = 16'h1300;
  X_LUT4 DLX_EXinst_Ker6483746_G (
    .ADR0(DLX_EXinst_N63129),
    .ADR1(DLX_IDinst_IR_function_field_3_1),
    .ADR2(DLX_IDinst_IR_function_field_2_1),
    .ADR3(DLX_IDinst_reg_out_A[31]),
    .O(N127871)
  );
  defparam DLX_EXinst_Ker6483746_F.INIT = 16'hFE04;
  X_LUT4 DLX_EXinst_Ker6483746_F (
    .ADR0(DLX_IDinst_IR_function_field_3_1),
    .ADR1(\DLX_EXinst_Mshift__n0024_Sh[27] ),
    .ADR2(DLX_IDinst_IR_function_field_2_1),
    .ADR3(DLX_IDinst_reg_out_A[31]),
    .O(N127869)
  );
  X_BUF \N101253/XUSED  (
    .I(\N101253/F5MUX ),
    .O(N101253)
  );
  X_MUX2 DLX_EXinst_Ker6539928 (
    .IA(N127829),
    .IB(N127831),
    .SEL(DLX_IDinst_IR_function_field_3_1),
    .O(\N97521/F5MUX )
  );
  defparam DLX_EXinst_Ker6539928_G.INIT = 16'hFC0C;
  X_LUT4 DLX_EXinst_Ker6539928_G (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N63499),
    .ADR2(DLX_IDinst_IR_function_field[0]),
    .ADR3(DLX_EXinst_N62996),
    .O(N127831)
  );
  defparam DLX_EXinst_Ker6539928_F.INIT = 16'hFA0A;
  X_LUT4 DLX_EXinst_Ker6539928_F (
    .ADR0(DLX_EXinst_N63334),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_IR_function_field[0]),
    .ADR3(DLX_EXinst_N62921),
    .O(N127829)
  );
  X_BUF \N97521/XUSED  (
    .I(\N97521/F5MUX ),
    .O(N97521)
  );
  X_MUX2 DLX_EXinst_Ker6487265 (
    .IA(N127634),
    .IB(N127636),
    .SEL(DLX_IDinst_reg_out_B[5]),
    .O(\CHOICE3198/F5MUX )
  );
  defparam DLX_EXinst_Ker6487265_G.INIT = 16'h5070;
  X_LUT4 DLX_EXinst_Ker6487265_G (
    .ADR0(DLX_IDinst_reg_out_B_3_1),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(DLX_IDinst_reg_out_B_2_1),
    .O(N127636)
  );
  defparam DLX_EXinst_Ker6487265_F.INIT = 16'hF8F0;
  X_LUT4 DLX_EXinst_Ker6487265_F (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(DLX_IDinst_reg_out_B_2_1),
    .ADR2(CHOICE3196),
    .ADR3(DLX_IDinst_reg_out_B_3_1),
    .O(N127634)
  );
  X_BUF \CHOICE3198/XUSED  (
    .I(\CHOICE3198/F5MUX ),
    .O(CHOICE3198)
  );
  X_MUX2 DLX_EXinst_Ker6489244 (
    .IA(N127909),
    .IB(N127911),
    .SEL(DLX_IDinst_reg_out_B[5]),
    .O(\CHOICE2542/F5MUX )
  );
  defparam DLX_EXinst_Ker6489244_G.INIT = 16'h1300;
  X_LUT4 DLX_EXinst_Ker6489244_G (
    .ADR0(DLX_IDinst_reg_out_B_2_1),
    .ADR1(DLX_IDinst_reg_out_B_3_1),
    .ADR2(DLX_EXinst_N63157),
    .ADR3(DLX_IDinst_reg_out_A[31]),
    .O(N127911)
  );
  defparam DLX_EXinst_Ker6489244_F.INIT = 16'hCCF0;
  X_LUT4 DLX_EXinst_Ker6489244_F (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[31]),
    .ADR2(\DLX_EXinst_Mshift__n0023_Sh[27] ),
    .ADR3(DLX_EXinst_N62740),
    .O(N127909)
  );
  X_BUF \CHOICE2542/XUSED  (
    .I(\CHOICE2542/F5MUX ),
    .O(CHOICE2542)
  );
  X_MUX2 \DLX_EXinst_Mshift__n0027_Sh<40>  (
    .IA(N127624),
    .IB(N127626),
    .SEL(DLX_IDinst_IR_function_field_3_1),
    .O(\DLX_EXinst_Mshift__n0027_Sh<40>/F5MUX )
  );
  defparam \DLX_EXinst_Mshift__n0027_Sh<40>_G .INIT = 16'h0100;
  X_LUT4 \DLX_EXinst_Mshift__n0027_Sh<40>_G  (
    .ADR0(DLX_IDinst_IR_function_field_0_1),
    .ADR1(DLX_IDinst_IR_function_field_1_1),
    .ADR2(DLX_IDinst_IR_function_field_2_1),
    .ADR3(DLX_IDinst_reg_out_A[0]),
    .O(N127626)
  );
  defparam \DLX_EXinst_Mshift__n0027_Sh<40>_F .INIT = 16'hFDA8;
  X_LUT4 \DLX_EXinst_Mshift__n0027_Sh<40>_F  (
    .ADR0(DLX_IDinst_IR_function_field_2_1),
    .ADR1(CHOICE1006),
    .ADR2(CHOICE1012),
    .ADR3(\DLX_EXinst_Mshift__n0027_Sh[8] ),
    .O(N127624)
  );
  X_BUF \DLX_EXinst_Mshift__n0027_Sh<40>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0027_Sh<40>/F5MUX ),
    .O(\DLX_EXinst_Mshift__n0027_Sh[40] )
  );
  X_MUX2 DLX_EXinst_Ker6486759 (
    .IA(N127889),
    .IB(N127891),
    .SEL(DLX_IDinst_reg_out_B[5]),
    .O(\CHOICE3124/F5MUX )
  );
  defparam DLX_EXinst_Ker6486759_G.INIT = 16'h2F20;
  X_LUT4 DLX_EXinst_Ker6486759_G (
    .ADR0(\DLX_EXinst_Mshift__n0023_Sh[61] ),
    .ADR1(DLX_IDinst_reg_out_B_2_1),
    .ADR2(DLX_IDinst_reg_out_B_3_1),
    .ADR3(DLX_IDinst_reg_out_A[31]),
    .O(N127891)
  );
  defparam DLX_EXinst_Ker6486759_F.INIT = 16'hFF0C;
  X_LUT4 DLX_EXinst_Ker6486759_F (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N62966),
    .ADR2(DLX_IDinst_reg_out_B_2_1),
    .ADR3(CHOICE3112),
    .O(N127889)
  );
  X_BUF \CHOICE3124/XUSED  (
    .I(\CHOICE3124/F5MUX ),
    .O(CHOICE3124)
  );
  X_MUX2 \DLX_EXinst__n0006<9>155  (
    .IA(N127689),
    .IB(N127691),
    .SEL(DLX_IDinst_reg_out_B[3]),
    .O(\CHOICE4587/F5MUX )
  );
  defparam \DLX_EXinst__n0006<9>155_G .INIT = 16'hD800;
  X_LUT4 \DLX_EXinst__n0006<9>155_G  (
    .ADR0(DLX_IDinst_reg_out_B[2]),
    .ADR1(\DLX_EXinst_Mshift__n0026_Sh[21] ),
    .ADR2(\DLX_EXinst_Mshift__n0026_Sh[17] ),
    .ADR3(DLX_EXinst_N62631),
    .O(N127691)
  );
  defparam \DLX_EXinst__n0006<9>155_F .INIT = 16'hE200;
  X_LUT4 \DLX_EXinst__n0006<9>155_F  (
    .ADR0(\DLX_EXinst_Mshift__n0023_Sh[9] ),
    .ADR1(DLX_IDinst_reg_out_B[2]),
    .ADR2(\DLX_EXinst_Mshift__n0026_Sh[13] ),
    .ADR3(DLX_EXinst_N62631),
    .O(N127689)
  );
  X_BUF \CHOICE4587/XUSED  (
    .I(\CHOICE4587/F5MUX ),
    .O(CHOICE4587)
  );
  X_MUX2 \DLX_EXinst_Mshift__n0027_Sh<42>  (
    .IA(N127594),
    .IB(N127596),
    .SEL(DLX_IDinst_IR_function_field_2_1),
    .O(\DLX_EXinst_Mshift__n0027_Sh<42>/F5MUX )
  );
  defparam \DLX_EXinst_Mshift__n0027_Sh<42>_G .INIT = 16'h00AC;
  X_LUT4 \DLX_EXinst_Mshift__n0027_Sh<42>_G  (
    .ADR0(N94155),
    .ADR1(DLX_EXinst_N63479),
    .ADR2(DLX_IDinst_IR_function_field_0_1),
    .ADR3(DLX_IDinst_IR_function_field_3_1),
    .O(N127596)
  );
  defparam \DLX_EXinst_Mshift__n0027_Sh<42>_F .INIT = 16'hBB88;
  X_LUT4 \DLX_EXinst_Mshift__n0027_Sh<42>_F  (
    .ADR0(\DLX_EXinst_Mshift__n0027_Sh[2] ),
    .ADR1(DLX_IDinst_IR_function_field_3_1),
    .ADR2(VCC),
    .ADR3(\DLX_EXinst_Mshift__n0027_Sh[10] ),
    .O(N127594)
  );
  X_BUF \DLX_EXinst_Mshift__n0027_Sh<42>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0027_Sh<42>/F5MUX ),
    .O(\DLX_EXinst_Mshift__n0027_Sh[42] )
  );
  X_MUX2 \DLX_EXinst_Mshift__n0027_Sh<43>  (
    .IA(N127604),
    .IB(N127606),
    .SEL(DLX_IDinst_IR_function_field_2_1),
    .O(\DLX_EXinst_Mshift__n0027_Sh<43>/F5MUX )
  );
  defparam \DLX_EXinst_Mshift__n0027_Sh<43>_G .INIT = 16'h0C0A;
  X_LUT4 \DLX_EXinst_Mshift__n0027_Sh<43>_G  (
    .ADR0(DLX_EXinst_N62766),
    .ADR1(DLX_EXinst_N63479),
    .ADR2(DLX_IDinst_IR_function_field_3_1),
    .ADR3(DLX_IDinst_IR_function_field_0_1),
    .O(N127606)
  );
  defparam \DLX_EXinst_Mshift__n0027_Sh<43>_F .INIT = 16'hFACC;
  X_LUT4 \DLX_EXinst_Mshift__n0027_Sh<43>_F  (
    .ADR0(CHOICE994),
    .ADR1(\DLX_EXinst_Mshift__n0027_Sh[11] ),
    .ADR2(CHOICE1000),
    .ADR3(DLX_IDinst_IR_function_field_3_1),
    .O(N127604)
  );
  X_BUF \DLX_EXinst_Mshift__n0027_Sh<43>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0027_Sh<43>/F5MUX ),
    .O(\DLX_EXinst_Mshift__n0027_Sh[43] )
  );
  X_MUX2 DLX_EXinst_Ker64877107_SW0 (
    .IA(N127804),
    .IB(N127806),
    .SEL(DLX_IDinst_reg_out_B[5]),
    .O(\N126268/F5MUX )
  );
  defparam DLX_EXinst_Ker64877107_SW0_G.INIT = 16'h3070;
  X_LUT4 DLX_EXinst_Ker64877107_SW0_G (
    .ADR0(DLX_IDinst_reg_out_B_2_1),
    .ADR1(DLX_IDinst_reg_out_B_3_1),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(DLX_EXinst_N63157),
    .O(N127806)
  );
  defparam DLX_EXinst_Ker64877107_SW0_F.INIT = 16'hF5F0;
  X_LUT4 DLX_EXinst_Ker64877107_SW0_F (
    .ADR0(DLX_IDinst_reg_out_B_2_1),
    .ADR1(VCC),
    .ADR2(CHOICE2980),
    .ADR3(DLX_EXinst_N66431),
    .O(N127804)
  );
  X_BUF \N126268/XUSED  (
    .I(\N126268/F5MUX ),
    .O(N126268)
  );
  X_MUX2 DLX_EXinst_Ker65088 (
    .IA(N127814),
    .IB(N127816),
    .SEL(DLX_IDinst_reg_out_B[5]),
    .O(\DLX_EXinst_N65090/F5MUX )
  );
  defparam DLX_EXinst_Ker65088_G.INIT = 16'h1050;
  X_LUT4 DLX_EXinst_Ker65088_G (
    .ADR0(DLX_EXinst_N62740),
    .ADR1(DLX_IDinst_reg_out_B[0]),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(DLX_IDinst_reg_out_B[1]),
    .O(N127816)
  );
  defparam DLX_EXinst_Ker65088_F.INIT = 16'hCCCA;
  X_LUT4 DLX_EXinst_Ker65088_F (
    .ADR0(DLX_EXinst_N62721),
    .ADR1(DLX_IDinst_reg_out_A[31]),
    .ADR2(DLX_IDinst_reg_out_B[1]),
    .ADR3(DLX_EXinst_N62740),
    .O(N127814)
  );
  X_BUF \DLX_EXinst_N65090/XUSED  (
    .I(\DLX_EXinst_N65090/F5MUX ),
    .O(DLX_EXinst_N65090)
  );
  X_MUX2 DLX_EXinst_Ker64498 (
    .IA(N127769),
    .IB(N127771),
    .SEL(DLX_IDinst_reg_out_B_2_1),
    .O(\DLX_EXinst_N64500/F5MUX )
  );
  defparam DLX_EXinst_Ker64498_G.INIT = 16'h0AAC;
  X_LUT4 DLX_EXinst_Ker64498_G (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(\DLX_EXinst_Mshift__n0026_Sh[24] ),
    .ADR2(DLX_IDinst_reg_out_B[5]),
    .ADR3(DLX_IDinst_reg_out_B_3_1),
    .O(N127771)
  );
  defparam DLX_EXinst_Ker64498_F.INIT = 16'hCCF0;
  X_LUT4 DLX_EXinst_Ker64498_F (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[31]),
    .ADR2(DLX_EXinst_N62727),
    .ADR3(DLX_IDinst_reg_out_B[5]),
    .O(N127769)
  );
  X_BUF \DLX_EXinst_N64500/XUSED  (
    .I(\DLX_EXinst_N64500/F5MUX ),
    .O(DLX_EXinst_N64500)
  );
  X_MUX2 \DLX_IFinst__n0003<0>  (
    .IA(N128079),
    .IB(N128081),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[0])
  );
  defparam \DLX_IFinst__n0003<0>_G .INIT = 16'hBB88;
  X_LUT4 \DLX_IFinst__n0003<0>_G  (
    .ADR0(IR[0]),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(VCC),
    .ADR3(DLX_IFinst_IR_previous[0]),
    .O(N128081)
  );
  defparam \DLX_IFinst__n0003<0>_F .INIT = 16'hEF20;
  X_LUT4 \DLX_IFinst__n0003<0>_F  (
    .ADR0(DLX_IFinst_IR_curr[0]),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(DLX_IFinst_stalled),
    .ADR3(IR[0]),
    .O(N128079)
  );
  X_MUX2 \DLX_IFinst__n0003<1>  (
    .IA(N128004),
    .IB(N128006),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[1])
  );
  defparam \DLX_IFinst__n0003<1>_G .INIT = 16'hFA0A;
  X_LUT4 \DLX_IFinst__n0003<1>_G  (
    .ADR0(DLX_IFinst_IR_previous[1]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(IR[1]),
    .O(N128006)
  );
  defparam \DLX_IFinst__n0003<1>_F .INIT = 16'hEF40;
  X_LUT4 \DLX_IFinst__n0003<1>_F  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(DLX_IFinst_IR_curr[1]),
    .ADR2(DLX_IFinst_stalled),
    .ADR3(IR[1]),
    .O(N128004)
  );
  X_MUX2 \DLX_IFinst__n0003<2>  (
    .IA(N128039),
    .IB(N128041),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[2])
  );
  defparam \DLX_IFinst__n0003<2>_G .INIT = 16'hB8B8;
  X_LUT4 \DLX_IFinst__n0003<2>_G  (
    .ADR0(IR[2]),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(DLX_IFinst_IR_previous[2]),
    .ADR3(VCC),
    .O(N128041)
  );
  defparam \DLX_IFinst__n0003<2>_F .INIT = 16'hE2F0;
  X_LUT4 \DLX_IFinst__n0003<2>_F  (
    .ADR0(DLX_IFinst_IR_curr[2]),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(IR[2]),
    .ADR3(DLX_IFinst_stalled),
    .O(N128039)
  );
  X_MUX2 \DLX_IFinst__n0003<3>  (
    .IA(N127979),
    .IB(N127981),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[3])
  );
  defparam \DLX_IFinst__n0003<3>_G .INIT = 16'hBB88;
  X_LUT4 \DLX_IFinst__n0003<3>_G  (
    .ADR0(IR[3]),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(VCC),
    .ADR3(DLX_IFinst_IR_previous[3]),
    .O(N127981)
  );
  defparam \DLX_IFinst__n0003<3>_F .INIT = 16'hAEA2;
  X_LUT4 \DLX_IFinst__n0003<3>_F  (
    .ADR0(IR[3]),
    .ADR1(DLX_IFinst_stalled),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(DLX_IFinst_IR_curr[3]),
    .O(N127979)
  );
  X_MUX2 \DLX_IFinst__n0003<4>  (
    .IA(N127959),
    .IB(N127961),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[4])
  );
  defparam \DLX_IFinst__n0003<4>_G .INIT = 16'hD8D8;
  X_LUT4 \DLX_IFinst__n0003<4>_G  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(IR[4]),
    .ADR2(DLX_IFinst_IR_previous[4]),
    .ADR3(VCC),
    .O(N127961)
  );
  defparam \DLX_IFinst__n0003<4>_F .INIT = 16'hEF40;
  X_LUT4 \DLX_IFinst__n0003<4>_F  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(DLX_IFinst_IR_curr[4]),
    .ADR2(DLX_IFinst_stalled),
    .ADR3(IR[4]),
    .O(N127959)
  );
  X_MUX2 \DLX_IFinst__n0003<5>  (
    .IA(N127984),
    .IB(N127986),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[5])
  );
  defparam \DLX_IFinst__n0003<5>_G .INIT = 16'hCACA;
  X_LUT4 \DLX_IFinst__n0003<5>_G  (
    .ADR0(DLX_IFinst_IR_previous[5]),
    .ADR1(IR[5]),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(VCC),
    .O(N127986)
  );
  defparam \DLX_IFinst__n0003<5>_F .INIT = 16'hE4F0;
  X_LUT4 \DLX_IFinst__n0003<5>_F  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(DLX_IFinst_IR_curr[5]),
    .ADR2(IR[5]),
    .ADR3(DLX_IFinst_stalled),
    .O(N127984)
  );
  X_MUX2 \DLX_IFinst__n0003<6>  (
    .IA(N127874),
    .IB(N127876),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[6])
  );
  defparam \DLX_IFinst__n0003<6>_G .INIT = 16'hF0AA;
  X_LUT4 \DLX_IFinst__n0003<6>_G  (
    .ADR0(DLX_IFinst_IR_previous[6]),
    .ADR1(VCC),
    .ADR2(IR[6]),
    .ADR3(DLX_IDinst_branch_sig),
    .O(N127876)
  );
  defparam \DLX_IFinst__n0003<6>_F .INIT = 16'hF2D0;
  X_LUT4 \DLX_IFinst__n0003<6>_F  (
    .ADR0(DLX_IFinst_stalled),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(IR[6]),
    .ADR3(DLX_IFinst_IR_curr[6]),
    .O(N127874)
  );
  X_MUX2 \DLX_IFinst__n0003<7>  (
    .IA(N127964),
    .IB(N127966),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[7])
  );
  defparam \DLX_IFinst__n0003<7>_G .INIT = 16'hDD88;
  X_LUT4 \DLX_IFinst__n0003<7>_G  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(IR[7]),
    .ADR2(VCC),
    .ADR3(DLX_IFinst_IR_previous[7]),
    .O(N127966)
  );
  defparam \DLX_IFinst__n0003<7>_F .INIT = 16'hACAA;
  X_LUT4 \DLX_IFinst__n0003<7>_F  (
    .ADR0(IR[7]),
    .ADR1(DLX_IFinst_IR_curr[7]),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(DLX_IFinst_stalled),
    .O(N127964)
  );
  X_MUX2 \DLX_IFinst__n0003<8>  (
    .IA(N127744),
    .IB(N127746),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[8])
  );
  defparam \DLX_IFinst__n0003<8>_G .INIT = 16'hF0CC;
  X_LUT4 \DLX_IFinst__n0003<8>_G  (
    .ADR0(VCC),
    .ADR1(DLX_IFinst_IR_previous[8]),
    .ADR2(IR[8]),
    .ADR3(DLX_IDinst_branch_sig),
    .O(N127746)
  );
  defparam \DLX_IFinst__n0003<8>_F .INIT = 16'hF4B0;
  X_LUT4 \DLX_IFinst__n0003<8>_F  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(DLX_IFinst_stalled),
    .ADR2(IR[8]),
    .ADR3(DLX_IFinst_IR_curr[8]),
    .O(N127744)
  );
  X_MUX2 \DLX_IFinst__n0003<9>  (
    .IA(N127774),
    .IB(N127776),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[9])
  );
  defparam \DLX_IFinst__n0003<9>_G .INIT = 16'hCACA;
  X_LUT4 \DLX_IFinst__n0003<9>_G  (
    .ADR0(DLX_IFinst_IR_previous[9]),
    .ADR1(IR[9]),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(VCC),
    .O(N127776)
  );
  defparam \DLX_IFinst__n0003<9>_F .INIT = 16'hAEA2;
  X_LUT4 \DLX_IFinst__n0003<9>_F  (
    .ADR0(IR[9]),
    .ADR1(DLX_IFinst_stalled),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(DLX_IFinst_IR_curr[9]),
    .O(N127774)
  );
  X_MUX2 \DLX_EXinst_Mshift__n0028_Sh<59>  (
    .IA(N128089),
    .IB(N128091),
    .SEL(DLX_IDinst_IR_function_field_2_1),
    .O(\DLX_EXinst_Mshift__n0028_Sh<59>/F5MUX )
  );
  defparam \DLX_EXinst_Mshift__n0028_Sh<59>_G .INIT = 16'h0100;
  X_LUT4 \DLX_EXinst_Mshift__n0028_Sh<59>_G  (
    .ADR0(DLX_IDinst_IR_function_field_3_1),
    .ADR1(DLX_IDinst_IR_function_field_1_1),
    .ADR2(DLX_IDinst_IR_function_field_0_1),
    .ADR3(DLX_IDinst_reg_out_A[31]),
    .O(N128091)
  );
  defparam \DLX_EXinst_Mshift__n0028_Sh<59>_F .INIT = 16'h3210;
  X_LUT4 \DLX_EXinst_Mshift__n0028_Sh<59>_F  (
    .ADR0(DLX_IDinst_IR_function_field_1_1),
    .ADR1(DLX_IDinst_IR_function_field_3_1),
    .ADR2(N93799),
    .ADR3(DLX_EXinst_N62709),
    .O(N128089)
  );
  X_BUF \DLX_EXinst_Mshift__n0028_Sh<59>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0028_Sh<59>/F5MUX ),
    .O(\DLX_EXinst_Mshift__n0028_Sh[59] )
  );
  X_MUX2 \DLX_EXinst__n0006<10>177  (
    .IA(N127709),
    .IB(N127711),
    .SEL(DLX_IDinst_reg_out_B[3]),
    .O(\CHOICE4531/F5MUX )
  );
  defparam \DLX_EXinst__n0006<10>177_G .INIT = 16'hE200;
  X_LUT4 \DLX_EXinst__n0006<10>177_G  (
    .ADR0(\DLX_EXinst_Mshift__n0026_Sh[18] ),
    .ADR1(DLX_IDinst_reg_out_B[2]),
    .ADR2(\DLX_EXinst_Mshift__n0026_Sh[22] ),
    .ADR3(DLX_EXinst_N62631),
    .O(N127711)
  );
  defparam \DLX_EXinst__n0006<10>177_F .INIT = 16'hE200;
  X_LUT4 \DLX_EXinst__n0006<10>177_F  (
    .ADR0(\DLX_EXinst_Mshift__n0026_Sh[10] ),
    .ADR1(DLX_IDinst_reg_out_B[2]),
    .ADR2(\DLX_EXinst_Mshift__n0026_Sh[14] ),
    .ADR3(DLX_EXinst_N62631),
    .O(N127709)
  );
  X_BUF \CHOICE4531/XUSED  (
    .I(\CHOICE4531/F5MUX ),
    .O(CHOICE4531)
  );
  X_MUX2 \DLX_EXinst__n0006<31>224_SW0  (
    .IA(N127669),
    .IB(N127671),
    .SEL(DLX_IDinst_reg_out_B[4]),
    .O(\N126500/F5MUX )
  );
  defparam \DLX_EXinst__n0006<31>224_SW0_G .INIT = 16'hC044;
  X_LUT4 \DLX_EXinst__n0006<31>224_SW0_G  (
    .ADR0(N93695),
    .ADR1(DLX_EXinst__n0048),
    .ADR2(DLX_EXinst_N62916),
    .ADR3(DLX_IDinst_reg_out_B[3]),
    .O(N127671)
  );
  defparam \DLX_EXinst__n0006<31>224_SW0_F .INIT = 16'hA088;
  X_LUT4 \DLX_EXinst__n0006<31>224_SW0_F  (
    .ADR0(DLX_EXinst__n0048),
    .ADR1(N126169),
    .ADR2(N100843),
    .ADR3(DLX_IDinst_reg_out_B[2]),
    .O(N127669)
  );
  X_BUF \N126500/XUSED  (
    .I(\N126500/F5MUX ),
    .O(N126500)
  );
  X_MUX2 \DLX_EXinst__n0006<30>202  (
    .IA(N127729),
    .IB(N127731),
    .SEL(DLX_IDinst_reg_out_B[4]),
    .O(\CHOICE5297/F5MUX )
  );
  defparam \DLX_EXinst__n0006<30>202_G .INIT = 16'h880A;
  X_LUT4 \DLX_EXinst__n0006<30>202_G  (
    .ADR0(DLX_EXinst__n0048),
    .ADR1(DLX_EXinst_N62911),
    .ADR2(N93747),
    .ADR3(DLX_IDinst_reg_out_B[3]),
    .O(N127731)
  );
  defparam \DLX_EXinst__n0006<30>202_F .INIT = 16'hC480;
  X_LUT4 \DLX_EXinst__n0006<30>202_F  (
    .ADR0(DLX_IDinst_reg_out_B[2]),
    .ADR1(DLX_EXinst__n0048),
    .ADR2(N97017),
    .ADR3(CHOICE5291),
    .O(N127729)
  );
  X_BUF \CHOICE5297/XUSED  (
    .I(\CHOICE5297/F5MUX ),
    .O(CHOICE5297)
  );
  X_MUX2 \DLX_EXinst__n0006<1>129_SW0_SW0  (
    .IA(N127954),
    .IB(N127956),
    .SEL(DLX_IDinst_IR_function_field[3]),
    .O(\N127444/F5MUX )
  );
  defparam \DLX_EXinst__n0006<1>129_SW0_SW0_G .INIT = 16'hB8B8;
  X_LUT4 \DLX_EXinst__n0006<1>129_SW0_SW0_G  (
    .ADR0(DLX_EXinst_N63489),
    .ADR1(DLX_IDinst_IR_function_field[0]),
    .ADR2(DLX_EXinst_N62981),
    .ADR3(VCC),
    .O(N127956)
  );
  defparam \DLX_EXinst__n0006<1>129_SW0_SW0_F .INIT = 16'hFC30;
  X_LUT4 \DLX_EXinst__n0006<1>129_SW0_SW0_F  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_IR_function_field[0]),
    .ADR2(DLX_EXinst_N65135),
    .ADR3(DLX_EXinst_N64474),
    .O(N127954)
  );
  X_BUF \N127444/XUSED  (
    .I(\N127444/F5MUX ),
    .O(N127444)
  );
  X_MUX2 \DLX_EXinst__n0006<31>426  (
    .IA(N127714),
    .IB(N127716),
    .SEL(DLX_IDinst_IR_function_field[4]),
    .O(\CHOICE5815/F5MUX )
  );
  defparam \DLX_EXinst__n0006<31>426_G .INIT = 16'hB080;
  X_LUT4 \DLX_EXinst__n0006<31>426_G  (
    .ADR0(DLX_EXinst_N62831),
    .ADR1(DLX_IDinst_IR_function_field[3]),
    .ADR2(DLX_EXinst__n0081),
    .ADR3(N93383),
    .O(N127716)
  );
  defparam \DLX_EXinst__n0006<31>426_F .INIT = 16'hA808;
  X_LUT4 \DLX_EXinst__n0006<31>426_F  (
    .ADR0(DLX_EXinst__n0081),
    .ADR1(N126154),
    .ADR2(DLX_IDinst_IR_function_field[2]),
    .ADR3(N100919),
    .O(N127714)
  );
  X_BUF \CHOICE5815/XUSED  (
    .I(\CHOICE5815/F5MUX ),
    .O(CHOICE5815)
  );
  X_MUX2 \DLX_EXinst__n0006<31>542  (
    .IA(N127819),
    .IB(N127821),
    .SEL(DLX_IDinst_reg_out_A[31]),
    .O(\CHOICE5842/F5MUX )
  );
  defparam \DLX_EXinst__n0006<31>542_G .INIT = 16'hFEFC;
  X_LUT4 \DLX_EXinst__n0006<31>542_G  (
    .ADR0(DLX_EXinst__n0078),
    .ADR1(DLX_EXinst__n0079),
    .ADR2(CHOICE5839),
    .ADR3(\DLX_IDinst_Imm[31] ),
    .O(N127821)
  );
  defparam \DLX_EXinst__n0006<31>542_F .INIT = 16'hEE00;
  X_LUT4 \DLX_EXinst__n0006<31>542_F  (
    .ADR0(DLX_EXinst__n0079),
    .ADR1(DLX_EXinst__n0080),
    .ADR2(VCC),
    .ADR3(\DLX_IDinst_Imm[31] ),
    .O(N127819)
  );
  X_BUF \CHOICE5842/XUSED  (
    .I(\CHOICE5842/F5MUX ),
    .O(CHOICE5842)
  );
  X_MUX2 \DLX_EXinst__n0006<16>280  (
    .IA(N128014),
    .IB(N128016),
    .SEL(DLX_IDinst_reg_out_B[4]),
    .O(\CHOICE5166/F5MUX )
  );
  defparam \DLX_EXinst__n0006<16>280_G .INIT = 16'h0002;
  X_LUT4 \DLX_EXinst__n0006<16>280_G  (
    .ADR0(DLX_IDinst_reg_out_A[0]),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(DLX_IDinst_reg_out_B[0]),
    .ADR3(DLX_EXinst_N62740),
    .O(N128016)
  );
  defparam \DLX_EXinst__n0006<16>280_F .INIT = 16'hFF0A;
  X_LUT4 \DLX_EXinst__n0006<16>280_F  (
    .ADR0(DLX_EXinst_N64914),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[2]),
    .ADR3(CHOICE5162),
    .O(N128014)
  );
  X_BUF \CHOICE5166/XUSED  (
    .I(\CHOICE5166/F5MUX ),
    .O(CHOICE5166)
  );
  X_MUX2 \DLX_EXinst__n0006<16>196  (
    .IA(N127899),
    .IB(N127901),
    .SEL(DLX_IDinst_reg_out_B[4]),
    .O(\CHOICE5140/F5MUX )
  );
  defparam \DLX_EXinst__n0006<16>196_G .INIT = 16'h2200;
  X_LUT4 \DLX_EXinst__n0006<16>196_G  (
    .ADR0(N111221),
    .ADR1(DLX_IDinst_reg_out_B[5]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[31]),
    .O(N127901)
  );
  defparam \DLX_EXinst__n0006<16>196_F .INIT = 16'hD080;
  X_LUT4 \DLX_EXinst__n0006<16>196_F  (
    .ADR0(DLX_IDinst_reg_out_B[2]),
    .ADR1(DLX_EXinst_N62727),
    .ADR2(DLX_EXinst_N62631),
    .ADR3(DLX_EXinst_N64319),
    .O(N127899)
  );
  X_BUF \CHOICE5140/XUSED  (
    .I(\CHOICE5140/F5MUX ),
    .O(CHOICE5140)
  );
  X_MUX2 \DLX_EXinst__n0006<17>267  (
    .IA(N128024),
    .IB(N128026),
    .SEL(DLX_IDinst_reg_out_B[3]),
    .O(\CHOICE5637/F5MUX )
  );
  defparam \DLX_EXinst__n0006<17>267_G .INIT = 16'hC808;
  X_LUT4 \DLX_EXinst__n0006<17>267_G  (
    .ADR0(\DLX_EXinst_Mshift__n0025_Sh[9] ),
    .ADR1(DLX_EXinst__n0048),
    .ADR2(DLX_IDinst_reg_out_B[2]),
    .ADR3(\DLX_EXinst_Mshift__n0025_Sh[5] ),
    .O(N128026)
  );
  defparam \DLX_EXinst__n0006<17>267_F .INIT = 16'hC840;
  X_LUT4 \DLX_EXinst__n0006<17>267_F  (
    .ADR0(DLX_IDinst_reg_out_B[2]),
    .ADR1(DLX_EXinst__n0048),
    .ADR2(N93487),
    .ADR3(\DLX_EXinst_Mshift__n0025_Sh[13] ),
    .O(N128024)
  );
  X_BUF \CHOICE5637/XUSED  (
    .I(\CHOICE5637/F5MUX ),
    .O(CHOICE5637)
  );
  X_MUX2 \DLX_EXinst__n0006<18>267  (
    .IA(N127844),
    .IB(N127846),
    .SEL(DLX_IDinst_reg_out_B[3]),
    .O(\CHOICE5471/F5MUX )
  );
  defparam \DLX_EXinst__n0006<18>267_G .INIT = 16'hAC00;
  X_LUT4 \DLX_EXinst__n0006<18>267_G  (
    .ADR0(\DLX_EXinst_Mshift__n0025_Sh[6] ),
    .ADR1(\DLX_EXinst_Mshift__n0025_Sh[10] ),
    .ADR2(DLX_IDinst_reg_out_B[2]),
    .ADR3(DLX_EXinst__n0048),
    .O(N127846)
  );
  defparam \DLX_EXinst__n0006<18>267_F .INIT = 16'h8C80;
  X_LUT4 \DLX_EXinst__n0006<18>267_F  (
    .ADR0(\DLX_EXinst_Mshift__n0025_Sh[14] ),
    .ADR1(DLX_EXinst__n0048),
    .ADR2(DLX_IDinst_reg_out_B[2]),
    .ADR3(N93537),
    .O(N127844)
  );
  X_BUF \CHOICE5471/XUSED  (
    .I(\CHOICE5471/F5MUX ),
    .O(CHOICE5471)
  );
  X_MUX2 \DLX_EXinst__n0006<19>243  (
    .IA(N127644),
    .IB(N127646),
    .SEL(DLX_IDinst_reg_out_B[4]),
    .O(\CHOICE4994/F5MUX )
  );
  defparam \DLX_EXinst__n0006<19>243_G .INIT = 16'h0032;
  X_LUT4 \DLX_EXinst__n0006<19>243_G  (
    .ADR0(CHOICE1054),
    .ADR1(DLX_IDinst_reg_out_B[2]),
    .ADR2(CHOICE1060),
    .ADR3(DLX_IDinst_reg_out_B[3]),
    .O(N127646)
  );
  defparam \DLX_EXinst__n0006<19>243_F .INIT = 16'hF4F4;
  X_LUT4 \DLX_EXinst__n0006<19>243_F  (
    .ADR0(DLX_IDinst_reg_out_B[2]),
    .ADR1(DLX_EXinst_N63920),
    .ADR2(CHOICE4990),
    .ADR3(VCC),
    .O(N127644)
  );
  X_BUF \CHOICE4994/XUSED  (
    .I(\CHOICE4994/F5MUX ),
    .O(CHOICE4994)
  );
  X_MUX2 \DLX_EXinst__n0006<28>202  (
    .IA(N127599),
    .IB(N127601),
    .SEL(DLX_IDinst_reg_out_B[4]),
    .O(\CHOICE5222/F5MUX )
  );
  defparam \DLX_EXinst__n0006<28>202_G .INIT = 16'h80B0;
  X_LUT4 \DLX_EXinst__n0006<28>202_G  (
    .ADR0(DLX_EXinst_N62901),
    .ADR1(DLX_IDinst_reg_out_B[3]),
    .ADR2(DLX_EXinst__n0048),
    .ADR3(N93587),
    .O(N127601)
  );
  defparam \DLX_EXinst__n0006<28>202_F .INIT = 16'h8C80;
  X_LUT4 \DLX_EXinst__n0006<28>202_F  (
    .ADR0(N97161),
    .ADR1(DLX_EXinst__n0048),
    .ADR2(DLX_IDinst_reg_out_B[2]),
    .ADR3(CHOICE5216),
    .O(N127599)
  );
  X_BUF \CHOICE5222/XUSED  (
    .I(\CHOICE5222/F5MUX ),
    .O(CHOICE5222)
  );
  X_MUX2 \DLX_EXinst__n0006<29>202  (
    .IA(N127679),
    .IB(N127681),
    .SEL(DLX_IDinst_reg_out_B[4]),
    .O(\CHOICE5374/F5MUX )
  );
  defparam \DLX_EXinst__n0006<29>202_G .INIT = 16'hC404;
  X_LUT4 \DLX_EXinst__n0006<29>202_G  (
    .ADR0(N93641),
    .ADR1(DLX_EXinst__n0048),
    .ADR2(DLX_IDinst_reg_out_B[3]),
    .ADR3(DLX_EXinst_N62906),
    .O(N127681)
  );
  defparam \DLX_EXinst__n0006<29>202_F .INIT = 16'h8A80;
  X_LUT4 \DLX_EXinst__n0006<29>202_F  (
    .ADR0(DLX_EXinst__n0048),
    .ADR1(N97089),
    .ADR2(DLX_IDinst_reg_out_B[2]),
    .ADR3(CHOICE5368),
    .O(N127679)
  );
  X_BUF \CHOICE5374/XUSED  (
    .I(\CHOICE5374/F5MUX ),
    .O(CHOICE5374)
  );
  X_MUX2 \DLX_EXinst__n0006<3>129_SW0_SW0  (
    .IA(N127659),
    .IB(N127661),
    .SEL(DLX_IDinst_IR_function_field[3]),
    .O(\N127440/F5MUX )
  );
  defparam \DLX_EXinst__n0006<3>129_SW0_SW0_G .INIT = 16'hAFA0;
  X_LUT4 \DLX_EXinst__n0006<3>129_SW0_SW0_G  (
    .ADR0(DLX_EXinst_N63494),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_IR_function_field[0]),
    .ADR3(DLX_EXinst_N62986),
    .O(N127661)
  );
  defparam \DLX_EXinst__n0006<3>129_SW0_SW0_F .INIT = 16'hDD88;
  X_LUT4 \DLX_EXinst__n0006<3>129_SW0_SW0_F  (
    .ADR0(DLX_IDinst_IR_function_field[0]),
    .ADR1(DLX_EXinst_N64909),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N65165),
    .O(N127659)
  );
  X_BUF \N127440/XUSED  (
    .I(\N127440/F5MUX ),
    .O(N127440)
  );
  defparam DLX_IFinst_NPC_0_1_137.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_0_1_137 (
    .I(\NPC_eff<0>/OD ),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\NPC_eff<0>/OFF/RST ),
    .O(DLX_IFinst_NPC_0_1)
  );
  X_OR2 \NPC_eff<0>/OFF/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\NPC_eff<0>/OFF/RST )
  );
  X_MUX2 DLX_EXinst_Ker65384107_SW0 (
    .IA(N127974),
    .IB(N127976),
    .SEL(\DLX_IDinst_Imm[5] ),
    .O(\N126272/F5MUX )
  );
  defparam DLX_EXinst_Ker65384107_SW0_G.INIT = 16'h02AA;
  X_LUT4 DLX_EXinst_Ker65384107_SW0_G (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(DLX_IDinst_IR_function_field_2_1),
    .ADR2(DLX_EXinst_N63129),
    .ADR3(DLX_IDinst_IR_function_field_3_1),
    .O(N127976)
  );
  defparam DLX_EXinst_Ker65384107_SW0_F.INIT = 16'hF0FC;
  X_LUT4 DLX_EXinst_Ker65384107_SW0_F (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N66421),
    .ADR2(CHOICE3007),
    .ADR3(DLX_IDinst_IR_function_field_2_1),
    .O(N127974)
  );
  X_BUF \N126272/XUSED  (
    .I(\N126272/F5MUX ),
    .O(N126272)
  );
  X_ONE \vram_out_vga_eff/LOGIC_ONE_138  (
    .O(\vram_out_vga_eff/LOGIC_ONE )
  );
  X_MUX2 \Mmux__COND_2_inst_mux_f6_0.F51_139  (
    .IA(\NLW_Mmux__COND_2_inst_mux_f6_0.F51_IA_UNCONNECTED ),
    .IB(\vram_out_vga<4>_rt ),
    .SEL(\vram_out_vga_eff/LOGIC_ONE ),
    .O(\Mmux__COND_2_inst_mux_f6_0.F51 )
  );
  defparam \vram_out_vga<4>_rt_140 .INIT = 16'hCCCC;
  X_LUT4 \vram_out_vga<4>_rt_140  (
    .ADR0(VCC),
    .ADR1(vram_out_vga[4]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\vram_out_vga<4>_rt )
  );
  X_BUF \vram_out_vga_eff/YUSED  (
    .I(\vram_out_vga_eff/F6MUX ),
    .O(vram_out_vga_eff)
  );
  X_MUX2 Mmux__COND_2_inst_mux_f6_0 (
    .IA(Mmux__COND_2__net2),
    .IB(\Mmux__COND_2_inst_mux_f6_0.F51 ),
    .SEL(vga_address[14]),
    .O(\vram_out_vga_eff/F6MUX )
  );
  X_MUX2 \DLX_EXinst_Mshift__n0023_Sh<27>  (
    .IA(N128049),
    .IB(N128051),
    .SEL(DLX_IDinst_reg_out_B[1]),
    .O(\DLX_EXinst_Mshift__n0023_Sh<27>/F5MUX )
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<27>_G .INIT = 16'hF0CC;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<27>_G  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[29]),
    .ADR2(DLX_IDinst_reg_out_A[30]),
    .ADR3(DLX_IDinst_reg_out_B[0]),
    .O(N128051)
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<27>_F .INIT = 16'hFC0C;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<27>_F  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[27]),
    .ADR2(DLX_IDinst_reg_out_B[0]),
    .ADR3(DLX_IDinst_reg_out_A[28]),
    .O(N128049)
  );
  X_BUF \DLX_EXinst_Mshift__n0023_Sh<27>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0023_Sh<27>/F5MUX ),
    .O(\DLX_EXinst_Mshift__n0023_Sh[27] )
  );
  X_ZERO \vga_top_vga1_Madd_addressout_inst_lut2_331/LOGIC_ZERO_141  (
    .O(\vga_top_vga1_Madd_addressout_inst_lut2_331/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_Madd_addressout_inst_cy_465_142 (
    .IA(vga_top_vga1_gridhcounter[5]),
    .IB(\vga_top_vga1_Madd_addressout_inst_lut2_331/LOGIC_ZERO ),
    .SEL(\vga_top_vga1_Madd_addressout_inst_lut2_331/FROM ),
    .O(vga_top_vga1_Madd_addressout_inst_cy_465)
  );
  defparam vga_top_vga1_Madd_addressout_inst_lut2_3311.INIT = 16'h5A5A;
  X_LUT4 vga_top_vga1_Madd_addressout_inst_lut2_3311 (
    .ADR0(vga_top_vga1_gridhcounter[5]),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_gridvcounter[0]),
    .ADR3(VCC),
    .O(\vga_top_vga1_Madd_addressout_inst_lut2_331/FROM )
  );
  defparam vga_top_vga1_Madd_addressout_inst_lut2_3321.INIT = 16'h6666;
  X_LUT4 vga_top_vga1_Madd_addressout_inst_lut2_3321 (
    .ADR0(vga_top_vga1_gridhcounter[6]),
    .ADR1(vga_top_vga1_gridvcounter[1]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(vga_top_vga1_Madd_addressout_inst_lut2_332)
  );
  X_BUF \vga_top_vga1_Madd_addressout_inst_lut2_331/COUTUSED  (
    .I(\vga_top_vga1_Madd_addressout_inst_lut2_331/CYMUXG ),
    .O(vga_top_vga1_Madd_addressout_inst_cy_466)
  );
  X_BUF \vga_top_vga1_Madd_addressout_inst_lut2_331/XUSED  (
    .I(\vga_top_vga1_Madd_addressout_inst_lut2_331/FROM ),
    .O(vga_top_vga1_Madd_addressout_inst_lut2_331)
  );
  X_BUF \vga_top_vga1_Madd_addressout_inst_lut2_331/YUSED  (
    .I(\vga_top_vga1_Madd_addressout_inst_lut2_331/XORG ),
    .O(vga_address[6])
  );
  X_MUX2 vga_top_vga1_Madd_addressout_inst_cy_466_143 (
    .IA(vga_top_vga1_gridhcounter[6]),
    .IB(vga_top_vga1_Madd_addressout_inst_cy_465),
    .SEL(vga_top_vga1_Madd_addressout_inst_lut2_332),
    .O(\vga_top_vga1_Madd_addressout_inst_lut2_331/CYMUXG )
  );
  X_XOR2 vga_top_vga1_Madd_addressout_inst_sum_254 (
    .I0(vga_top_vga1_Madd_addressout_inst_cy_465),
    .I1(vga_top_vga1_Madd_addressout_inst_lut2_332),
    .O(\vga_top_vga1_Madd_addressout_inst_lut2_331/XORG )
  );
  X_MUX2 vga_top_vga1_Madd_addressout_inst_cy_467_144 (
    .IA(vga_top_vga1_gridhcounter[7]),
    .IB(\vga_address<7>/CYINIT ),
    .SEL(vga_top_vga1_Madd_addressout_inst_lut2_333),
    .O(vga_top_vga1_Madd_addressout_inst_cy_467)
  );
  X_XOR2 vga_top_vga1_Madd_addressout_inst_sum_255 (
    .I0(\vga_address<7>/CYINIT ),
    .I1(vga_top_vga1_Madd_addressout_inst_lut2_333),
    .O(\vga_address<7>/XORF )
  );
  defparam vga_top_vga1_Madd_addressout_inst_lut2_3331.INIT = 16'h9966;
  X_LUT4 vga_top_vga1_Madd_addressout_inst_lut2_3331 (
    .ADR0(vga_top_vga1_gridhcounter[7]),
    .ADR1(vga_top_vga1_gridvcounter[2]),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_gridvcounter[0]),
    .O(vga_top_vga1_Madd_addressout_inst_lut2_333)
  );
  defparam vga_top_vga1_Madd_addressout_inst_lut2_3341.INIT = 16'h6666;
  X_LUT4 vga_top_vga1_Madd_addressout_inst_lut2_3341 (
    .ADR0(vga_top_vga1_gridhcounter[8]),
    .ADR1(vga_top_vga1_Mmult__n0043_inst_lut2_317),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(vga_top_vga1_Madd_addressout_inst_lut2_334)
  );
  X_BUF \vga_address<7>/COUTUSED  (
    .I(\vga_address<7>/CYMUXG ),
    .O(vga_top_vga1_Madd_addressout_inst_cy_468)
  );
  X_BUF \vga_address<7>/XUSED  (
    .I(\vga_address<7>/XORF ),
    .O(vga_address[7])
  );
  X_BUF \vga_address<7>/YUSED  (
    .I(\vga_address<7>/XORG ),
    .O(vga_address[8])
  );
  X_MUX2 vga_top_vga1_Madd_addressout_inst_cy_468_145 (
    .IA(vga_top_vga1_gridhcounter[8]),
    .IB(vga_top_vga1_Madd_addressout_inst_cy_467),
    .SEL(vga_top_vga1_Madd_addressout_inst_lut2_334),
    .O(\vga_address<7>/CYMUXG )
  );
  X_XOR2 vga_top_vga1_Madd_addressout_inst_sum_256 (
    .I0(vga_top_vga1_Madd_addressout_inst_cy_467),
    .I1(vga_top_vga1_Madd_addressout_inst_lut2_334),
    .O(\vga_address<7>/XORG )
  );
  X_BUF \vga_address<7>/CYINIT_146  (
    .I(vga_top_vga1_Madd_addressout_inst_cy_466),
    .O(\vga_address<7>/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0061_inst_cy_212_147 (
    .IA(DLX_IDinst_reg_out_A[14]),
    .IB(\DLX_EXinst_Mcompar__n0061_inst_cy_213/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0061_inst_lut2_148),
    .O(DLX_EXinst_Mcompar__n0061_inst_cy_212)
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_lut2_1481.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_lut2_1481 (
    .ADR0(DLX_IDinst_reg_out_A[14]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[14]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0061_inst_lut2_148)
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_lut2_1491.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_lut2_1491 (
    .ADR0(DLX_IDinst_reg_out_A[15]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[15]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0061_inst_lut2_149)
  );
  X_BUF \DLX_EXinst_Mcompar__n0061_inst_cy_213/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0061_inst_cy_213/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0061_inst_cy_213)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0061_inst_cy_213_148 (
    .IA(DLX_IDinst_reg_out_A[15]),
    .IB(DLX_EXinst_Mcompar__n0061_inst_cy_212),
    .SEL(DLX_EXinst_Mcompar__n0061_inst_lut2_149),
    .O(\DLX_EXinst_Mcompar__n0061_inst_cy_213/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0061_inst_cy_213/CYINIT_149  (
    .I(DLX_EXinst_Mcompar__n0061_inst_cy_211),
    .O(\DLX_EXinst_Mcompar__n0061_inst_cy_213/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0061_inst_cy_214_150 (
    .IA(DLX_IDinst_reg_out_A[16]),
    .IB(\DLX_EXinst_Mcompar__n0061_inst_cy_215/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0061_inst_lut2_150),
    .O(DLX_EXinst_Mcompar__n0061_inst_cy_214)
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_lut2_1501.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_lut2_1501 (
    .ADR0(DLX_IDinst_reg_out_A[16]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[16]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0061_inst_lut2_150)
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_lut2_1511.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_lut2_1511 (
    .ADR0(DLX_IDinst_reg_out_A[17]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[17]),
    .O(DLX_EXinst_Mcompar__n0061_inst_lut2_151)
  );
  X_BUF \DLX_EXinst_Mcompar__n0061_inst_cy_215/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0061_inst_cy_215/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0061_inst_cy_215)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0061_inst_cy_215_151 (
    .IA(DLX_IDinst_reg_out_A[17]),
    .IB(DLX_EXinst_Mcompar__n0061_inst_cy_214),
    .SEL(DLX_EXinst_Mcompar__n0061_inst_lut2_151),
    .O(\DLX_EXinst_Mcompar__n0061_inst_cy_215/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0061_inst_cy_215/CYINIT_152  (
    .I(DLX_EXinst_Mcompar__n0061_inst_cy_213),
    .O(\DLX_EXinst_Mcompar__n0061_inst_cy_215/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0061_inst_cy_216_153 (
    .IA(DLX_IDinst_reg_out_A[18]),
    .IB(\DLX_EXinst_Mcompar__n0061_inst_cy_217/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0061_inst_lut2_152),
    .O(DLX_EXinst_Mcompar__n0061_inst_cy_216)
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_lut2_1521.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_lut2_1521 (
    .ADR0(DLX_IDinst_reg_out_A[18]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[18]),
    .O(DLX_EXinst_Mcompar__n0061_inst_lut2_152)
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_lut2_1531.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_lut2_1531 (
    .ADR0(DLX_IDinst_reg_out_A[19]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[19]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0061_inst_lut2_153)
  );
  X_BUF \DLX_EXinst_Mcompar__n0061_inst_cy_217/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0061_inst_cy_217/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0061_inst_cy_217)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0061_inst_cy_217_154 (
    .IA(DLX_IDinst_reg_out_A[19]),
    .IB(DLX_EXinst_Mcompar__n0061_inst_cy_216),
    .SEL(DLX_EXinst_Mcompar__n0061_inst_lut2_153),
    .O(\DLX_EXinst_Mcompar__n0061_inst_cy_217/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0061_inst_cy_217/CYINIT_155  (
    .I(DLX_EXinst_Mcompar__n0061_inst_cy_215),
    .O(\DLX_EXinst_Mcompar__n0061_inst_cy_217/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0061_inst_cy_218_156 (
    .IA(DLX_IDinst_reg_out_A[20]),
    .IB(\DLX_EXinst_Mcompar__n0061_inst_cy_219/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0061_inst_lut2_154),
    .O(DLX_EXinst_Mcompar__n0061_inst_cy_218)
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_lut2_1541.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_lut2_1541 (
    .ADR0(DLX_IDinst_reg_out_A[20]),
    .ADR1(DLX_IDinst_reg_out_B[20]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0061_inst_lut2_154)
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_lut2_1551.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_lut2_1551 (
    .ADR0(DLX_IDinst_reg_out_A[21]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[21]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0061_inst_lut2_155)
  );
  X_BUF \DLX_EXinst_Mcompar__n0061_inst_cy_219/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0061_inst_cy_219/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0061_inst_cy_219)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0061_inst_cy_219_157 (
    .IA(DLX_IDinst_reg_out_A[21]),
    .IB(DLX_EXinst_Mcompar__n0061_inst_cy_218),
    .SEL(DLX_EXinst_Mcompar__n0061_inst_lut2_155),
    .O(\DLX_EXinst_Mcompar__n0061_inst_cy_219/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0061_inst_cy_219/CYINIT_158  (
    .I(DLX_EXinst_Mcompar__n0061_inst_cy_217),
    .O(\DLX_EXinst_Mcompar__n0061_inst_cy_219/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0061_inst_cy_220_159 (
    .IA(DLX_IDinst_reg_out_A[22]),
    .IB(\DLX_EXinst_Mcompar__n0061_inst_cy_221/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0061_inst_lut2_156),
    .O(DLX_EXinst_Mcompar__n0061_inst_cy_220)
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_lut2_1561.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_lut2_1561 (
    .ADR0(DLX_IDinst_reg_out_A[22]),
    .ADR1(DLX_IDinst_reg_out_B[22]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0061_inst_lut2_156)
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_lut2_1571.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_lut2_1571 (
    .ADR0(DLX_IDinst_reg_out_A[23]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[23]),
    .O(DLX_EXinst_Mcompar__n0061_inst_lut2_157)
  );
  X_BUF \DLX_EXinst_Mcompar__n0061_inst_cy_221/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0061_inst_cy_221/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0061_inst_cy_221)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0061_inst_cy_221_160 (
    .IA(DLX_IDinst_reg_out_A[23]),
    .IB(DLX_EXinst_Mcompar__n0061_inst_cy_220),
    .SEL(DLX_EXinst_Mcompar__n0061_inst_lut2_157),
    .O(\DLX_EXinst_Mcompar__n0061_inst_cy_221/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0061_inst_cy_221/CYINIT_161  (
    .I(DLX_EXinst_Mcompar__n0061_inst_cy_219),
    .O(\DLX_EXinst_Mcompar__n0061_inst_cy_221/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0061_inst_cy_222_162 (
    .IA(DLX_IDinst_reg_out_A[24]),
    .IB(\DLX_EXinst_Mcompar__n0061_inst_cy_223/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0061_inst_lut2_158),
    .O(DLX_EXinst_Mcompar__n0061_inst_cy_222)
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_lut2_1581.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_lut2_1581 (
    .ADR0(DLX_IDinst_reg_out_A[24]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[24]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0061_inst_lut2_158)
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_lut2_1591.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_lut2_1591 (
    .ADR0(DLX_IDinst_reg_out_A[25]),
    .ADR1(DLX_IDinst_reg_out_B[25]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0061_inst_lut2_159)
  );
  X_BUF \DLX_EXinst_Mcompar__n0061_inst_cy_223/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0061_inst_cy_223/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0061_inst_cy_223)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0061_inst_cy_223_163 (
    .IA(DLX_IDinst_reg_out_A[25]),
    .IB(DLX_EXinst_Mcompar__n0061_inst_cy_222),
    .SEL(DLX_EXinst_Mcompar__n0061_inst_lut2_159),
    .O(\DLX_EXinst_Mcompar__n0061_inst_cy_223/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0061_inst_cy_223/CYINIT_164  (
    .I(DLX_EXinst_Mcompar__n0061_inst_cy_221),
    .O(\DLX_EXinst_Mcompar__n0061_inst_cy_223/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0061_inst_cy_224_165 (
    .IA(DLX_IDinst_reg_out_A[26]),
    .IB(\DLX_EXinst_Mcompar__n0061_inst_cy_225/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0061_inst_lut2_160),
    .O(DLX_EXinst_Mcompar__n0061_inst_cy_224)
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_lut2_1601.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_lut2_1601 (
    .ADR0(DLX_IDinst_reg_out_A[26]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[26]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0061_inst_lut2_160)
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_lut2_1611.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_lut2_1611 (
    .ADR0(DLX_IDinst_reg_out_A[27]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[27]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0061_inst_lut2_161)
  );
  X_BUF \DLX_EXinst_Mcompar__n0061_inst_cy_225/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0061_inst_cy_225/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0061_inst_cy_225)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0061_inst_cy_225_166 (
    .IA(DLX_IDinst_reg_out_A[27]),
    .IB(DLX_EXinst_Mcompar__n0061_inst_cy_224),
    .SEL(DLX_EXinst_Mcompar__n0061_inst_lut2_161),
    .O(\DLX_EXinst_Mcompar__n0061_inst_cy_225/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0061_inst_cy_225/CYINIT_167  (
    .I(DLX_EXinst_Mcompar__n0061_inst_cy_223),
    .O(\DLX_EXinst_Mcompar__n0061_inst_cy_225/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0061_inst_cy_226_168 (
    .IA(DLX_IDinst_reg_out_A[28]),
    .IB(\DLX_EXinst_Mcompar__n0061_inst_cy_227/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0061_inst_lut2_162),
    .O(DLX_EXinst_Mcompar__n0061_inst_cy_226)
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_lut2_1621.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_lut2_1621 (
    .ADR0(DLX_IDinst_reg_out_A[28]),
    .ADR1(DLX_IDinst_reg_out_B[28]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0061_inst_lut2_162)
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_lut2_1631.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_lut2_1631 (
    .ADR0(DLX_IDinst_reg_out_A[29]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[29]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0061_inst_lut2_163)
  );
  X_BUF \DLX_EXinst_Mcompar__n0061_inst_cy_227/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0061_inst_cy_227/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0061_inst_cy_227)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0061_inst_cy_227_169 (
    .IA(DLX_IDinst_reg_out_A[29]),
    .IB(DLX_EXinst_Mcompar__n0061_inst_cy_226),
    .SEL(DLX_EXinst_Mcompar__n0061_inst_lut2_163),
    .O(\DLX_EXinst_Mcompar__n0061_inst_cy_227/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0061_inst_cy_227/CYINIT_170  (
    .I(DLX_EXinst_Mcompar__n0061_inst_cy_225),
    .O(\DLX_EXinst_Mcompar__n0061_inst_cy_227/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0061_inst_cy_228_171 (
    .IA(DLX_IDinst_reg_out_A[30]),
    .IB(\DLX_EXinst_reg_out_B_EX<30>/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0061_inst_lut2_164),
    .O(\DLX_EXinst_reg_out_B_EX<30>/CYMUXF )
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_lut2_1641.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_lut2_1641 (
    .ADR0(DLX_IDinst_reg_out_A[30]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[30]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0061_inst_lut2_164)
  );
  defparam \DLX_EXinst__n0007<30>1 .INIT = 16'hA0A0;
  X_LUT4 \DLX_EXinst__n0007<30>1  (
    .ADR0(DLX_IDinst_reg_out_B[30]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N66271),
    .ADR3(VCC),
    .O(DLX_EXinst__n0007[30])
  );
  X_BUF \DLX_EXinst_reg_out_B_EX<30>/XBUSED  (
    .I(\DLX_EXinst_reg_out_B_EX<30>/CYMUXF ),
    .O(DLX_EXinst_Mcompar__n0061_inst_cy_228)
  );
  X_BUF \DLX_EXinst_reg_out_B_EX<30>/CYINIT_172  (
    .I(DLX_EXinst_Mcompar__n0061_inst_cy_227),
    .O(\DLX_EXinst_reg_out_B_EX<30>/CYINIT )
  );
  X_ONE \vga_top_vga1_Mcompar__n0029_inst_cy_374/LOGIC_ONE_173  (
    .O(\vga_top_vga1_Mcompar__n0029_inst_cy_374/LOGIC_ONE )
  );
  X_ZERO \vga_top_vga1_Mcompar__n0029_inst_cy_374/LOGIC_ZERO_174  (
    .O(\vga_top_vga1_Mcompar__n0029_inst_cy_374/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0029_inst_cy_373_175 (
    .IA(\vga_top_vga1_Mcompar__n0029_inst_cy_374/LOGIC_ZERO ),
    .IB(\vga_top_vga1_Mcompar__n0029_inst_cy_374/LOGIC_ONE ),
    .SEL(vga_top_vga1_Mcompar__n0029_inst_lut1_22),
    .O(vga_top_vga1_Mcompar__n0029_inst_cy_373)
  );
  defparam vga_top_vga1_Mcompar__n0029_inst_lut1_221.INIT = 16'h00FF;
  X_LUT4 vga_top_vga1_Mcompar__n0029_inst_lut1_221 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[4]),
    .O(vga_top_vga1_Mcompar__n0029_inst_lut1_22)
  );
  defparam vga_top_vga1_Mcompar__n0029_inst_lut1_231.INIT = 16'h3333;
  X_LUT4 vga_top_vga1_Mcompar__n0029_inst_lut1_231 (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_hcounter[4]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(vga_top_vga1_Mcompar__n0029_inst_lut1_23)
  );
  X_BUF \vga_top_vga1_Mcompar__n0029_inst_cy_374/COUTUSED  (
    .I(\vga_top_vga1_Mcompar__n0029_inst_cy_374/CYMUXG ),
    .O(vga_top_vga1_Mcompar__n0029_inst_cy_374)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0029_inst_cy_374_176 (
    .IA(\vga_top_vga1_Mcompar__n0029_inst_cy_374/LOGIC_ZERO ),
    .IB(vga_top_vga1_Mcompar__n0029_inst_cy_373),
    .SEL(vga_top_vga1_Mcompar__n0029_inst_lut1_23),
    .O(\vga_top_vga1_Mcompar__n0029_inst_cy_374/CYMUXG )
  );
  X_ONE \vga_top_vga1_Mcompar__n0029_inst_cy_376/LOGIC_ONE_177  (
    .O(\vga_top_vga1_Mcompar__n0029_inst_cy_376/LOGIC_ONE )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0029_inst_cy_375_178 (
    .IA(\vga_top_vga1_Mcompar__n0029_inst_cy_376/LOGIC_ONE ),
    .IB(\vga_top_vga1_Mcompar__n0029_inst_cy_376/CYINIT ),
    .SEL(\$SIG_13 ),
    .O(vga_top_vga1_Mcompar__n0029_inst_cy_375)
  );
  defparam \$BEL_13 .INIT = 16'hAAAA;
  X_LUT4 \$BEL_13  (
    .ADR0(vga_top_vga1_hcounter[5]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\$SIG_13 )
  );
  defparam \$BEL_14 .INIT = 16'hFF00;
  X_LUT4 \$BEL_14  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[5]),
    .O(\$SIG_14 )
  );
  X_BUF \vga_top_vga1_Mcompar__n0029_inst_cy_376/COUTUSED  (
    .I(\vga_top_vga1_Mcompar__n0029_inst_cy_376/CYMUXG ),
    .O(vga_top_vga1_Mcompar__n0029_inst_cy_376)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0029_inst_cy_376_179 (
    .IA(\vga_top_vga1_Mcompar__n0029_inst_cy_376/LOGIC_ONE ),
    .IB(vga_top_vga1_Mcompar__n0029_inst_cy_375),
    .SEL(\$SIG_14 ),
    .O(\vga_top_vga1_Mcompar__n0029_inst_cy_376/CYMUXG )
  );
  X_BUF \vga_top_vga1_Mcompar__n0029_inst_cy_376/CYINIT_180  (
    .I(vga_top_vga1_Mcompar__n0029_inst_cy_374),
    .O(\vga_top_vga1_Mcompar__n0029_inst_cy_376/CYINIT )
  );
  X_ZERO \vga_top_vga1_Mcompar__n0029_inst_cy_378/LOGIC_ZERO_181  (
    .O(\vga_top_vga1_Mcompar__n0029_inst_cy_378/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0029_inst_cy_377_182 (
    .IA(\vga_top_vga1_Mcompar__n0029_inst_cy_378/LOGIC_ZERO ),
    .IB(\vga_top_vga1_Mcompar__n0029_inst_cy_378/CYINIT ),
    .SEL(vga_top_vga1_Mcompar__n0029_inst_lut4_51),
    .O(vga_top_vga1_Mcompar__n0029_inst_cy_377)
  );
  defparam vga_top_vga1_Mcompar__n0029_inst_lut4_511.INIT = 16'h0001;
  X_LUT4 vga_top_vga1_Mcompar__n0029_inst_lut4_511 (
    .ADR0(vga_top_vga1_hcounter[8]),
    .ADR1(vga_top_vga1_hcounter[6]),
    .ADR2(vga_top_vga1_hcounter[9]),
    .ADR3(vga_top_vga1_hcounter[7]),
    .O(vga_top_vga1_Mcompar__n0029_inst_lut4_51)
  );
  defparam vga_top_vga1_Mcompar__n0029_inst_lut4_521.INIT = 16'h0001;
  X_LUT4 vga_top_vga1_Mcompar__n0029_inst_lut4_521 (
    .ADR0(vga_top_vga1_hcounter[7]),
    .ADR1(vga_top_vga1_hcounter[6]),
    .ADR2(vga_top_vga1_hcounter[8]),
    .ADR3(vga_top_vga1_hcounter[9]),
    .O(vga_top_vga1_Mcompar__n0029_inst_lut4_52)
  );
  X_BUF \vga_top_vga1_Mcompar__n0029_inst_cy_378/COUTUSED  (
    .I(\vga_top_vga1_Mcompar__n0029_inst_cy_378/CYMUXG ),
    .O(vga_top_vga1_Mcompar__n0029_inst_cy_378)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0029_inst_cy_378_183 (
    .IA(\vga_top_vga1_Mcompar__n0029_inst_cy_378/LOGIC_ZERO ),
    .IB(vga_top_vga1_Mcompar__n0029_inst_cy_377),
    .SEL(vga_top_vga1_Mcompar__n0029_inst_lut4_52),
    .O(\vga_top_vga1_Mcompar__n0029_inst_cy_378/CYMUXG )
  );
  X_BUF \vga_top_vga1_Mcompar__n0029_inst_cy_378/CYINIT_184  (
    .I(vga_top_vga1_Mcompar__n0029_inst_cy_376),
    .O(\vga_top_vga1_Mcompar__n0029_inst_cy_378/CYINIT )
  );
  defparam DLX_EXinst_ALU_result_4_1_185.INIT = 1'b0;
  X_FF DLX_EXinst_ALU_result_4_1_185 (
    .I(\DM_addr_eff<4>/OD ),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DM_addr_eff<4>/OFF/RST ),
    .O(DLX_EXinst_ALU_result_4_1)
  );
  X_OR2 \DM_addr_eff<4>/OFF/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DM_addr_eff<4>/OFF/RST )
  );
  X_ZERO \vga_top_vga1__n0029/LOGIC_ZERO_186  (
    .O(\vga_top_vga1__n0029/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0029_inst_cy_379_187 (
    .IA(\vga_top_vga1__n0029/LOGIC_ZERO ),
    .IB(\vga_top_vga1__n0029/CYINIT ),
    .SEL(vga_top_vga1_Mcompar__n0029_inst_lut4_53),
    .O(vga_top_vga1_Mcompar__n0029_inst_cy_379)
  );
  defparam vga_top_vga1_Mcompar__n0029_inst_lut4_531.INIT = 16'h0001;
  X_LUT4 vga_top_vga1_Mcompar__n0029_inst_lut4_531 (
    .ADR0(vga_top_vga1_hcounter[11]),
    .ADR1(vga_top_vga1_hcounter[10]),
    .ADR2(vga_top_vga1_hcounter[12]),
    .ADR3(vga_top_vga1_hcounter[13]),
    .O(vga_top_vga1_Mcompar__n0029_inst_lut4_53)
  );
  defparam vga_top_vga1_Mcompar__n0029_inst_lut2_2751.INIT = 16'h0505;
  X_LUT4 vga_top_vga1_Mcompar__n0029_inst_lut2_2751 (
    .ADR0(vga_top_vga1_hcounter[14]),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_hcounter[15]),
    .ADR3(VCC),
    .O(vga_top_vga1_Mcompar__n0029_inst_lut2_275)
  );
  X_BUF \vga_top_vga1__n0029/COUTUSED  (
    .I(\vga_top_vga1__n0029/CYMUXG ),
    .O(vga_top_vga1__n0029)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0029_inst_cy_380 (
    .IA(\vga_top_vga1__n0029/LOGIC_ZERO ),
    .IB(vga_top_vga1_Mcompar__n0029_inst_cy_379),
    .SEL(vga_top_vga1_Mcompar__n0029_inst_lut2_275),
    .O(\vga_top_vga1__n0029/CYMUXG )
  );
  X_BUF \vga_top_vga1__n0029/CYINIT_188  (
    .I(vga_top_vga1_Mcompar__n0029_inst_cy_378),
    .O(\vga_top_vga1__n0029/CYINIT )
  );
  X_ONE \vga_top_vga1_Mcompar__n0037_inst_cy_475/LOGIC_ONE_189  (
    .O(\vga_top_vga1_Mcompar__n0037_inst_cy_475/LOGIC_ONE )
  );
  X_ZERO \vga_top_vga1_Mcompar__n0037_inst_cy_475/LOGIC_ZERO_190  (
    .O(\vga_top_vga1_Mcompar__n0037_inst_cy_475/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0037_inst_cy_474_191 (
    .IA(\vga_top_vga1_Mcompar__n0037_inst_cy_475/LOGIC_ZERO ),
    .IB(\vga_top_vga1_Mcompar__n0037_inst_cy_475/LOGIC_ONE ),
    .SEL(vga_top_vga1_Mcompar__n0037_inst_lut2_341),
    .O(vga_top_vga1_Mcompar__n0037_inst_cy_474)
  );
  defparam vga_top_vga1_Mcompar__n0037_inst_lut2_3411.INIT = 16'hAA00;
  X_LUT4 vga_top_vga1_Mcompar__n0037_inst_lut2_3411 (
    .ADR0(vga_top_vga1_hcounter[4]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[5]),
    .O(vga_top_vga1_Mcompar__n0037_inst_lut2_341)
  );
  defparam vga_top_vga1_Mcompar__n0037_inst_lut2_3421.INIT = 16'hF000;
  X_LUT4 vga_top_vga1_Mcompar__n0037_inst_lut2_3421 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_hcounter[5]),
    .ADR3(vga_top_vga1_hcounter[4]),
    .O(vga_top_vga1_Mcompar__n0037_inst_lut2_342)
  );
  X_BUF \vga_top_vga1_Mcompar__n0037_inst_cy_475/COUTUSED  (
    .I(\vga_top_vga1_Mcompar__n0037_inst_cy_475/CYMUXG ),
    .O(vga_top_vga1_Mcompar__n0037_inst_cy_475)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0037_inst_cy_475_192 (
    .IA(\vga_top_vga1_Mcompar__n0037_inst_cy_475/LOGIC_ZERO ),
    .IB(vga_top_vga1_Mcompar__n0037_inst_cy_474),
    .SEL(vga_top_vga1_Mcompar__n0037_inst_lut2_342),
    .O(\vga_top_vga1_Mcompar__n0037_inst_cy_475/CYMUXG )
  );
  X_ONE \vga_top_vga1_Mcompar__n0037_inst_cy_477/LOGIC_ONE_193  (
    .O(\vga_top_vga1_Mcompar__n0037_inst_cy_477/LOGIC_ONE )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0037_inst_cy_476_194 (
    .IA(\vga_top_vga1_Mcompar__n0037_inst_cy_477/LOGIC_ONE ),
    .IB(\vga_top_vga1_Mcompar__n0037_inst_cy_477/CYINIT ),
    .SEL(vga_top_vga1_Mcompar__n0037_inst_lut4_86),
    .O(vga_top_vga1_Mcompar__n0037_inst_cy_476)
  );
  defparam vga_top_vga1_Mcompar__n0037_inst_lut4_861.INIT = 16'h0001;
  X_LUT4 vga_top_vga1_Mcompar__n0037_inst_lut4_861 (
    .ADR0(vga_top_vga1_hcounter[9]),
    .ADR1(vga_top_vga1_hcounter[8]),
    .ADR2(vga_top_vga1_hcounter[7]),
    .ADR3(vga_top_vga1_hcounter[6]),
    .O(vga_top_vga1_Mcompar__n0037_inst_lut4_86)
  );
  defparam vga_top_vga1_Mcompar__n0037_inst_lut4_871.INIT = 16'h0001;
  X_LUT4 vga_top_vga1_Mcompar__n0037_inst_lut4_871 (
    .ADR0(vga_top_vga1_hcounter[8]),
    .ADR1(vga_top_vga1_hcounter[6]),
    .ADR2(vga_top_vga1_hcounter[9]),
    .ADR3(vga_top_vga1_hcounter[7]),
    .O(vga_top_vga1_Mcompar__n0037_inst_lut4_87)
  );
  X_BUF \vga_top_vga1_Mcompar__n0037_inst_cy_477/COUTUSED  (
    .I(\vga_top_vga1_Mcompar__n0037_inst_cy_477/CYMUXG ),
    .O(vga_top_vga1_Mcompar__n0037_inst_cy_477)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0037_inst_cy_477_195 (
    .IA(\vga_top_vga1_Mcompar__n0037_inst_cy_477/LOGIC_ONE ),
    .IB(vga_top_vga1_Mcompar__n0037_inst_cy_476),
    .SEL(vga_top_vga1_Mcompar__n0037_inst_lut4_87),
    .O(\vga_top_vga1_Mcompar__n0037_inst_cy_477/CYMUXG )
  );
  X_BUF \vga_top_vga1_Mcompar__n0037_inst_cy_477/CYINIT_196  (
    .I(vga_top_vga1_Mcompar__n0037_inst_cy_475),
    .O(\vga_top_vga1_Mcompar__n0037_inst_cy_477/CYINIT )
  );
  X_ONE \vga_top_vga1__n0037/LOGIC_ONE_197  (
    .O(\vga_top_vga1__n0037/LOGIC_ONE )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0037_inst_cy_478_198 (
    .IA(\vga_top_vga1__n0037/LOGIC_ONE ),
    .IB(\vga_top_vga1__n0037/CYINIT ),
    .SEL(vga_top_vga1_Mcompar__n0037_inst_lut4_88),
    .O(vga_top_vga1_Mcompar__n0037_inst_cy_478)
  );
  defparam vga_top_vga1_Mcompar__n0037_inst_lut4_881.INIT = 16'h0001;
  X_LUT4 vga_top_vga1_Mcompar__n0037_inst_lut4_881 (
    .ADR0(vga_top_vga1_hcounter[10]),
    .ADR1(vga_top_vga1_hcounter[11]),
    .ADR2(vga_top_vga1_hcounter[12]),
    .ADR3(vga_top_vga1_hcounter[13]),
    .O(vga_top_vga1_Mcompar__n0037_inst_lut4_88)
  );
  defparam vga_top_vga1_Mcompar__n0037_inst_lut2_3431.INIT = 16'h000F;
  X_LUT4 vga_top_vga1_Mcompar__n0037_inst_lut2_3431 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_hcounter[14]),
    .ADR3(vga_top_vga1_hcounter[15]),
    .O(vga_top_vga1_Mcompar__n0037_inst_lut2_343)
  );
  X_BUF \vga_top_vga1__n0037/COUTUSED  (
    .I(\vga_top_vga1__n0037/CYMUXG ),
    .O(vga_top_vga1__n0037)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0037_inst_cy_479 (
    .IA(\vga_top_vga1__n0037/LOGIC_ONE ),
    .IB(vga_top_vga1_Mcompar__n0037_inst_cy_478),
    .SEL(vga_top_vga1_Mcompar__n0037_inst_lut2_343),
    .O(\vga_top_vga1__n0037/CYMUXG )
  );
  X_BUF \vga_top_vga1__n0037/CYINIT_199  (
    .I(vga_top_vga1_Mcompar__n0037_inst_cy_477),
    .O(\vga_top_vga1__n0037/CYINIT )
  );
  X_ZERO \DLX_EXinst_Mcompar__n0055_inst_cy_119/LOGIC_ZERO_200  (
    .O(\DLX_EXinst_Mcompar__n0055_inst_cy_119/LOGIC_ZERO )
  );
  X_ONE \DLX_EXinst_Mcompar__n0055_inst_cy_119/LOGIC_ONE_201  (
    .O(\DLX_EXinst_Mcompar__n0055_inst_cy_119/LOGIC_ONE )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0055_inst_cy_118_202 (
    .IA(\DLX_EXinst_Mcompar__n0055_inst_cy_119/LOGIC_ONE ),
    .IB(\DLX_EXinst_Mcompar__n0055_inst_cy_119/LOGIC_ZERO ),
    .SEL(DLX_EXinst_Mcompar__n0055_inst_lut4_16),
    .O(DLX_EXinst_Mcompar__n0055_inst_cy_118)
  );
  defparam DLX_EXinst_Mcompar__n0055_inst_lut4_161.INIT = 16'h8421;
  X_LUT4 DLX_EXinst_Mcompar__n0055_inst_lut4_161 (
    .ADR0(DLX_IDinst_reg_out_A[1]),
    .ADR1(DLX_IDinst_reg_out_A[0]),
    .ADR2(DLX_IDinst_reg_out_B[1]),
    .ADR3(DLX_IDinst_reg_out_B[0]),
    .O(DLX_EXinst_Mcompar__n0055_inst_lut4_16)
  );
  defparam DLX_EXinst_Mcompar__n0055_inst_lut4_171.INIT = 16'h9009;
  X_LUT4 DLX_EXinst_Mcompar__n0055_inst_lut4_171 (
    .ADR0(DLX_IDinst_reg_out_A[2]),
    .ADR1(DLX_IDinst_reg_out_B_2_1),
    .ADR2(DLX_IDinst_reg_out_B_3_1),
    .ADR3(DLX_IDinst_reg_out_A[3]),
    .O(DLX_EXinst_Mcompar__n0055_inst_lut4_17)
  );
  X_BUF \DLX_EXinst_Mcompar__n0055_inst_cy_119/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0055_inst_cy_119/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0055_inst_cy_119)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0055_inst_cy_119_203 (
    .IA(\DLX_EXinst_Mcompar__n0055_inst_cy_119/LOGIC_ONE ),
    .IB(DLX_EXinst_Mcompar__n0055_inst_cy_118),
    .SEL(DLX_EXinst_Mcompar__n0055_inst_lut4_17),
    .O(\DLX_EXinst_Mcompar__n0055_inst_cy_119/CYMUXG )
  );
  X_ONE \DLX_EXinst_Mcompar__n0055_inst_cy_121/LOGIC_ONE_204  (
    .O(\DLX_EXinst_Mcompar__n0055_inst_cy_121/LOGIC_ONE )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0055_inst_cy_120_205 (
    .IA(\DLX_EXinst_Mcompar__n0055_inst_cy_121/LOGIC_ONE ),
    .IB(\DLX_EXinst_Mcompar__n0055_inst_cy_121/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0055_inst_lut4_18),
    .O(DLX_EXinst_Mcompar__n0055_inst_cy_120)
  );
  defparam DLX_EXinst_Mcompar__n0055_inst_lut4_181.INIT = 16'h8421;
  X_LUT4 DLX_EXinst_Mcompar__n0055_inst_lut4_181 (
    .ADR0(DLX_IDinst_reg_out_A[4]),
    .ADR1(DLX_IDinst_reg_out_A[5]),
    .ADR2(DLX_IDinst_reg_out_B[4]),
    .ADR3(DLX_IDinst_reg_out_B[5]),
    .O(DLX_EXinst_Mcompar__n0055_inst_lut4_18)
  );
  defparam DLX_EXinst_Mcompar__n0055_inst_lut4_191.INIT = 16'h8241;
  X_LUT4 DLX_EXinst_Mcompar__n0055_inst_lut4_191 (
    .ADR0(DLX_IDinst_reg_out_B[6]),
    .ADR1(DLX_IDinst_reg_out_A[7]),
    .ADR2(DLX_IDinst_reg_out_B[7]),
    .ADR3(DLX_IDinst_reg_out_A[6]),
    .O(DLX_EXinst_Mcompar__n0055_inst_lut4_19)
  );
  X_BUF \DLX_EXinst_Mcompar__n0055_inst_cy_121/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0055_inst_cy_121/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0055_inst_cy_121)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0055_inst_cy_121_206 (
    .IA(\DLX_EXinst_Mcompar__n0055_inst_cy_121/LOGIC_ONE ),
    .IB(DLX_EXinst_Mcompar__n0055_inst_cy_120),
    .SEL(DLX_EXinst_Mcompar__n0055_inst_lut4_19),
    .O(\DLX_EXinst_Mcompar__n0055_inst_cy_121/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0055_inst_cy_121/CYINIT_207  (
    .I(DLX_EXinst_Mcompar__n0055_inst_cy_119),
    .O(\DLX_EXinst_Mcompar__n0055_inst_cy_121/CYINIT )
  );
  X_ONE \DLX_EXinst_Mcompar__n0055_inst_cy_123/LOGIC_ONE_208  (
    .O(\DLX_EXinst_Mcompar__n0055_inst_cy_123/LOGIC_ONE )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0055_inst_cy_122_209 (
    .IA(\DLX_EXinst_Mcompar__n0055_inst_cy_123/LOGIC_ONE ),
    .IB(\DLX_EXinst_Mcompar__n0055_inst_cy_123/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0055_inst_lut4_20),
    .O(DLX_EXinst_Mcompar__n0055_inst_cy_122)
  );
  defparam DLX_EXinst_Mcompar__n0055_inst_lut4_201.INIT = 16'h8241;
  X_LUT4 DLX_EXinst_Mcompar__n0055_inst_lut4_201 (
    .ADR0(DLX_IDinst_reg_out_B[9]),
    .ADR1(DLX_IDinst_reg_out_A[8]),
    .ADR2(DLX_IDinst_reg_out_B[8]),
    .ADR3(DLX_IDinst_reg_out_A[9]),
    .O(DLX_EXinst_Mcompar__n0055_inst_lut4_20)
  );
  defparam DLX_EXinst_Mcompar__n0055_inst_lut4_211.INIT = 16'h8421;
  X_LUT4 DLX_EXinst_Mcompar__n0055_inst_lut4_211 (
    .ADR0(DLX_IDinst_reg_out_B[10]),
    .ADR1(DLX_IDinst_reg_out_B[11]),
    .ADR2(DLX_IDinst_reg_out_A[10]),
    .ADR3(DLX_IDinst_reg_out_A[11]),
    .O(DLX_EXinst_Mcompar__n0055_inst_lut4_21)
  );
  X_BUF \DLX_EXinst_Mcompar__n0055_inst_cy_123/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0055_inst_cy_123/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0055_inst_cy_123)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0055_inst_cy_123_210 (
    .IA(\DLX_EXinst_Mcompar__n0055_inst_cy_123/LOGIC_ONE ),
    .IB(DLX_EXinst_Mcompar__n0055_inst_cy_122),
    .SEL(DLX_EXinst_Mcompar__n0055_inst_lut4_21),
    .O(\DLX_EXinst_Mcompar__n0055_inst_cy_123/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0055_inst_cy_123/CYINIT_211  (
    .I(DLX_EXinst_Mcompar__n0055_inst_cy_121),
    .O(\DLX_EXinst_Mcompar__n0055_inst_cy_123/CYINIT )
  );
  X_ONE \DLX_EXinst_Mcompar__n0055_inst_cy_125/LOGIC_ONE_212  (
    .O(\DLX_EXinst_Mcompar__n0055_inst_cy_125/LOGIC_ONE )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0055_inst_cy_124_213 (
    .IA(\DLX_EXinst_Mcompar__n0055_inst_cy_125/LOGIC_ONE ),
    .IB(\DLX_EXinst_Mcompar__n0055_inst_cy_125/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0055_inst_lut4_22),
    .O(DLX_EXinst_Mcompar__n0055_inst_cy_124)
  );
  defparam DLX_EXinst_Mcompar__n0055_inst_lut4_221.INIT = 16'h8241;
  X_LUT4 DLX_EXinst_Mcompar__n0055_inst_lut4_221 (
    .ADR0(DLX_IDinst_reg_out_B[12]),
    .ADR1(DLX_IDinst_reg_out_A[13]),
    .ADR2(DLX_IDinst_reg_out_B[13]),
    .ADR3(DLX_IDinst_reg_out_A[12]),
    .O(DLX_EXinst_Mcompar__n0055_inst_lut4_22)
  );
  defparam DLX_EXinst_Mcompar__n0055_inst_lut4_231.INIT = 16'h8241;
  X_LUT4 DLX_EXinst_Mcompar__n0055_inst_lut4_231 (
    .ADR0(DLX_IDinst_reg_out_A[15]),
    .ADR1(DLX_IDinst_reg_out_A[14]),
    .ADR2(DLX_IDinst_reg_out_B[14]),
    .ADR3(DLX_IDinst_reg_out_B[15]),
    .O(DLX_EXinst_Mcompar__n0055_inst_lut4_23)
  );
  X_BUF \DLX_EXinst_Mcompar__n0055_inst_cy_125/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0055_inst_cy_125/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0055_inst_cy_125)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0055_inst_cy_125_214 (
    .IA(\DLX_EXinst_Mcompar__n0055_inst_cy_125/LOGIC_ONE ),
    .IB(DLX_EXinst_Mcompar__n0055_inst_cy_124),
    .SEL(DLX_EXinst_Mcompar__n0055_inst_lut4_23),
    .O(\DLX_EXinst_Mcompar__n0055_inst_cy_125/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0055_inst_cy_125/CYINIT_215  (
    .I(DLX_EXinst_Mcompar__n0055_inst_cy_123),
    .O(\DLX_EXinst_Mcompar__n0055_inst_cy_125/CYINIT )
  );
  X_ONE \DLX_EXinst_Mcompar__n0055_inst_cy_127/LOGIC_ONE_216  (
    .O(\DLX_EXinst_Mcompar__n0055_inst_cy_127/LOGIC_ONE )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0055_inst_cy_126_217 (
    .IA(\DLX_EXinst_Mcompar__n0055_inst_cy_127/LOGIC_ONE ),
    .IB(\DLX_EXinst_Mcompar__n0055_inst_cy_127/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0055_inst_lut4_24),
    .O(DLX_EXinst_Mcompar__n0055_inst_cy_126)
  );
  defparam DLX_EXinst_Mcompar__n0055_inst_lut4_241.INIT = 16'h8241;
  X_LUT4 DLX_EXinst_Mcompar__n0055_inst_lut4_241 (
    .ADR0(DLX_IDinst_reg_out_B[17]),
    .ADR1(DLX_IDinst_reg_out_A[16]),
    .ADR2(DLX_IDinst_reg_out_B[16]),
    .ADR3(DLX_IDinst_reg_out_A[17]),
    .O(DLX_EXinst_Mcompar__n0055_inst_lut4_24)
  );
  defparam DLX_EXinst_Mcompar__n0055_inst_lut4_251.INIT = 16'h8241;
  X_LUT4 DLX_EXinst_Mcompar__n0055_inst_lut4_251 (
    .ADR0(DLX_IDinst_reg_out_B[18]),
    .ADR1(DLX_IDinst_reg_out_B[19]),
    .ADR2(DLX_IDinst_reg_out_A[19]),
    .ADR3(DLX_IDinst_reg_out_A[18]),
    .O(DLX_EXinst_Mcompar__n0055_inst_lut4_25)
  );
  X_BUF \DLX_EXinst_Mcompar__n0055_inst_cy_127/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0055_inst_cy_127/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0055_inst_cy_127)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0055_inst_cy_127_218 (
    .IA(\DLX_EXinst_Mcompar__n0055_inst_cy_127/LOGIC_ONE ),
    .IB(DLX_EXinst_Mcompar__n0055_inst_cy_126),
    .SEL(DLX_EXinst_Mcompar__n0055_inst_lut4_25),
    .O(\DLX_EXinst_Mcompar__n0055_inst_cy_127/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0055_inst_cy_127/CYINIT_219  (
    .I(DLX_EXinst_Mcompar__n0055_inst_cy_125),
    .O(\DLX_EXinst_Mcompar__n0055_inst_cy_127/CYINIT )
  );
  X_ONE \DLX_EXinst_Mcompar__n0055_inst_cy_129/LOGIC_ONE_220  (
    .O(\DLX_EXinst_Mcompar__n0055_inst_cy_129/LOGIC_ONE )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0055_inst_cy_128_221 (
    .IA(\DLX_EXinst_Mcompar__n0055_inst_cy_129/LOGIC_ONE ),
    .IB(\DLX_EXinst_Mcompar__n0055_inst_cy_129/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0055_inst_lut4_26),
    .O(DLX_EXinst_Mcompar__n0055_inst_cy_128)
  );
  defparam DLX_EXinst_Mcompar__n0055_inst_lut4_261.INIT = 16'h8241;
  X_LUT4 DLX_EXinst_Mcompar__n0055_inst_lut4_261 (
    .ADR0(DLX_IDinst_reg_out_B[21]),
    .ADR1(DLX_IDinst_reg_out_A[20]),
    .ADR2(DLX_IDinst_reg_out_B[20]),
    .ADR3(DLX_IDinst_reg_out_A[21]),
    .O(DLX_EXinst_Mcompar__n0055_inst_lut4_26)
  );
  defparam DLX_EXinst_Mcompar__n0055_inst_lut4_271.INIT = 16'h8421;
  X_LUT4 DLX_EXinst_Mcompar__n0055_inst_lut4_271 (
    .ADR0(DLX_IDinst_reg_out_A[22]),
    .ADR1(DLX_IDinst_reg_out_A[23]),
    .ADR2(DLX_IDinst_reg_out_B[22]),
    .ADR3(DLX_IDinst_reg_out_B[23]),
    .O(DLX_EXinst_Mcompar__n0055_inst_lut4_27)
  );
  X_BUF \DLX_EXinst_Mcompar__n0055_inst_cy_129/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0055_inst_cy_129/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0055_inst_cy_129)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0055_inst_cy_129_222 (
    .IA(\DLX_EXinst_Mcompar__n0055_inst_cy_129/LOGIC_ONE ),
    .IB(DLX_EXinst_Mcompar__n0055_inst_cy_128),
    .SEL(DLX_EXinst_Mcompar__n0055_inst_lut4_27),
    .O(\DLX_EXinst_Mcompar__n0055_inst_cy_129/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0055_inst_cy_129/CYINIT_223  (
    .I(DLX_EXinst_Mcompar__n0055_inst_cy_127),
    .O(\DLX_EXinst_Mcompar__n0055_inst_cy_129/CYINIT )
  );
  X_ONE \DLX_EXinst_Mcompar__n0055_inst_cy_131/LOGIC_ONE_224  (
    .O(\DLX_EXinst_Mcompar__n0055_inst_cy_131/LOGIC_ONE )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0055_inst_cy_130_225 (
    .IA(\DLX_EXinst_Mcompar__n0055_inst_cy_131/LOGIC_ONE ),
    .IB(\DLX_EXinst_Mcompar__n0055_inst_cy_131/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0055_inst_lut4_28),
    .O(DLX_EXinst_Mcompar__n0055_inst_cy_130)
  );
  defparam DLX_EXinst_Mcompar__n0055_inst_lut4_281.INIT = 16'h8241;
  X_LUT4 DLX_EXinst_Mcompar__n0055_inst_lut4_281 (
    .ADR0(DLX_IDinst_reg_out_B[25]),
    .ADR1(DLX_IDinst_reg_out_B[24]),
    .ADR2(DLX_IDinst_reg_out_A[24]),
    .ADR3(DLX_IDinst_reg_out_A[25]),
    .O(DLX_EXinst_Mcompar__n0055_inst_lut4_28)
  );
  defparam DLX_EXinst_Mcompar__n0055_inst_lut4_291.INIT = 16'h8241;
  X_LUT4 DLX_EXinst_Mcompar__n0055_inst_lut4_291 (
    .ADR0(DLX_IDinst_reg_out_A[26]),
    .ADR1(DLX_IDinst_reg_out_B[27]),
    .ADR2(DLX_IDinst_reg_out_A[27]),
    .ADR3(DLX_IDinst_reg_out_B[26]),
    .O(DLX_EXinst_Mcompar__n0055_inst_lut4_29)
  );
  X_BUF \DLX_EXinst_Mcompar__n0055_inst_cy_131/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0055_inst_cy_131/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0055_inst_cy_131)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0055_inst_cy_131_226 (
    .IA(\DLX_EXinst_Mcompar__n0055_inst_cy_131/LOGIC_ONE ),
    .IB(DLX_EXinst_Mcompar__n0055_inst_cy_130),
    .SEL(DLX_EXinst_Mcompar__n0055_inst_lut4_29),
    .O(\DLX_EXinst_Mcompar__n0055_inst_cy_131/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0055_inst_cy_131/CYINIT_227  (
    .I(DLX_EXinst_Mcompar__n0055_inst_cy_129),
    .O(\DLX_EXinst_Mcompar__n0055_inst_cy_131/CYINIT )
  );
  X_ONE \DLX_EXinst__n0055/LOGIC_ONE_228  (
    .O(\DLX_EXinst__n0055/LOGIC_ONE )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0055_inst_cy_132_229 (
    .IA(\DLX_EXinst__n0055/LOGIC_ONE ),
    .IB(\DLX_EXinst__n0055/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0055_inst_lut4_30),
    .O(DLX_EXinst_Mcompar__n0055_inst_cy_132)
  );
  defparam DLX_EXinst_Mcompar__n0055_inst_lut4_301.INIT = 16'h8241;
  X_LUT4 DLX_EXinst_Mcompar__n0055_inst_lut4_301 (
    .ADR0(DLX_IDinst_reg_out_A[29]),
    .ADR1(DLX_IDinst_reg_out_A[28]),
    .ADR2(DLX_IDinst_reg_out_B[28]),
    .ADR3(DLX_IDinst_reg_out_B[29]),
    .O(DLX_EXinst_Mcompar__n0055_inst_lut4_30)
  );
  defparam DLX_EXinst_Mcompar__n0055_inst_lut4_311.INIT = 16'h9009;
  X_LUT4 DLX_EXinst_Mcompar__n0055_inst_lut4_311 (
    .ADR0(DLX_IDinst_reg_out_A[30]),
    .ADR1(DLX_IDinst_reg_out_B[30]),
    .ADR2(DLX_IDinst_reg_out_B[31]),
    .ADR3(DLX_IDinst_reg_out_A[31]),
    .O(DLX_EXinst_Mcompar__n0055_inst_lut4_31)
  );
  X_BUF \DLX_EXinst__n0055/COUTUSED  (
    .I(\DLX_EXinst__n0055/CYMUXG ),
    .O(DLX_EXinst__n0055)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0055_inst_cy_133 (
    .IA(\DLX_EXinst__n0055/LOGIC_ONE ),
    .IB(DLX_EXinst_Mcompar__n0055_inst_cy_132),
    .SEL(DLX_EXinst_Mcompar__n0055_inst_lut4_31),
    .O(\DLX_EXinst__n0055/CYMUXG )
  );
  X_BUF \DLX_EXinst__n0055/CYINIT_230  (
    .I(DLX_EXinst_Mcompar__n0055_inst_cy_131),
    .O(\DLX_EXinst__n0055/CYINIT )
  );
  X_ZERO \DLX_EXinst_Mcompar__n0063_inst_cy_231/LOGIC_ZERO_231  (
    .O(\DLX_EXinst_Mcompar__n0063_inst_cy_231/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_230_232 (
    .IA(DLX_IDinst_reg_out_B[0]),
    .IB(\DLX_EXinst_Mcompar__n0063_inst_cy_231/LOGIC_ZERO ),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_166),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_230)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_1661.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_1661 (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[0]),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_166)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_1671.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_1671 (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(DLX_IDinst_reg_out_A[1]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_167)
  );
  X_BUF \DLX_EXinst_Mcompar__n0063_inst_cy_231/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0063_inst_cy_231/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_231)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_231_233 (
    .IA(DLX_IDinst_reg_out_B[1]),
    .IB(DLX_EXinst_Mcompar__n0063_inst_cy_230),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_167),
    .O(\DLX_EXinst_Mcompar__n0063_inst_cy_231/CYMUXG )
  );
  X_ZERO \vga_address<9>/LOGIC_ZERO_234  (
    .O(\vga_address<9>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_Madd_addressout_inst_cy_469_235 (
    .IA(\vga_address<9>/LOGIC_ZERO ),
    .IB(\vga_address<9>/CYINIT ),
    .SEL(\vga_address<9>/FROM ),
    .O(vga_top_vga1_Madd_addressout_inst_cy_469)
  );
  X_XOR2 vga_top_vga1_Madd_addressout_inst_sum_257 (
    .I0(\vga_address<9>/CYINIT ),
    .I1(\vga_address<9>/FROM ),
    .O(\vga_address<9>/XORF )
  );
  defparam \vga_address<9>/F .INIT = 16'hCCCC;
  X_LUT4 \vga_address<9>/F  (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_Mmult__n0043_inst_lut2_318),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\vga_address<9>/FROM )
  );
  defparam \vga_address<9>/G .INIT = 16'hAAAA;
  X_LUT4 \vga_address<9>/G  (
    .ADR0(vga_top_vga1_Mmult__n0043_inst_lut2_319),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\vga_address<9>/GROM )
  );
  X_BUF \vga_address<9>/COUTUSED  (
    .I(\vga_address<9>/CYMUXG ),
    .O(vga_top_vga1_Madd_addressout_inst_cy_470)
  );
  X_BUF \vga_address<9>/XUSED  (
    .I(\vga_address<9>/XORF ),
    .O(vga_address[9])
  );
  X_BUF \vga_address<9>/YUSED  (
    .I(\vga_address<9>/XORG ),
    .O(vga_address[10])
  );
  X_MUX2 vga_top_vga1_Madd_addressout_inst_cy_470_236 (
    .IA(\vga_address<9>/LOGIC_ZERO ),
    .IB(vga_top_vga1_Madd_addressout_inst_cy_469),
    .SEL(\vga_address<9>/GROM ),
    .O(\vga_address<9>/CYMUXG )
  );
  X_XOR2 vga_top_vga1_Madd_addressout_inst_sum_258 (
    .I0(vga_top_vga1_Madd_addressout_inst_cy_469),
    .I1(\vga_address<9>/GROM ),
    .O(\vga_address<9>/XORG )
  );
  X_BUF \vga_address<9>/CYINIT_237  (
    .I(vga_top_vga1_Madd_addressout_inst_cy_468),
    .O(\vga_address<9>/CYINIT )
  );
  X_ZERO \vga_address<11>/LOGIC_ZERO_238  (
    .O(\vga_address<11>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_Madd_addressout_inst_cy_471_239 (
    .IA(\vga_address<11>/LOGIC_ZERO ),
    .IB(\vga_address<11>/CYINIT ),
    .SEL(\vga_address<11>/FROM ),
    .O(vga_top_vga1_Madd_addressout_inst_cy_471)
  );
  X_XOR2 vga_top_vga1_Madd_addressout_inst_sum_259 (
    .I0(\vga_address<11>/CYINIT ),
    .I1(\vga_address<11>/FROM ),
    .O(\vga_address<11>/XORF )
  );
  defparam \vga_address<11>/F .INIT = 16'hCCCC;
  X_LUT4 \vga_address<11>/F  (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_Mmult__n0043_inst_lut2_320),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\vga_address<11>/FROM )
  );
  defparam \vga_address<11>/G .INIT = 16'hAAAA;
  X_LUT4 \vga_address<11>/G  (
    .ADR0(vga_top_vga1_Mmult__n0043_inst_lut2_321),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\vga_address<11>/GROM )
  );
  X_BUF \vga_address<11>/COUTUSED  (
    .I(\vga_address<11>/CYMUXG ),
    .O(vga_top_vga1_Madd_addressout_inst_cy_472)
  );
  X_BUF \vga_address<11>/XUSED  (
    .I(\vga_address<11>/XORF ),
    .O(vga_address[11])
  );
  X_BUF \vga_address<11>/YUSED  (
    .I(\vga_address<11>/XORG ),
    .O(vga_address[12])
  );
  X_MUX2 vga_top_vga1_Madd_addressout_inst_cy_472_240 (
    .IA(\vga_address<11>/LOGIC_ZERO ),
    .IB(vga_top_vga1_Madd_addressout_inst_cy_471),
    .SEL(\vga_address<11>/GROM ),
    .O(\vga_address<11>/CYMUXG )
  );
  X_XOR2 vga_top_vga1_Madd_addressout_inst_sum_260 (
    .I0(vga_top_vga1_Madd_addressout_inst_cy_471),
    .I1(\vga_address<11>/GROM ),
    .O(\vga_address<11>/XORG )
  );
  X_BUF \vga_address<11>/CYINIT_241  (
    .I(vga_top_vga1_Madd_addressout_inst_cy_470),
    .O(\vga_address<11>/CYINIT )
  );
  defparam DLX_IFinst_NPC_1_1_242.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_1_1_242 (
    .I(\NPC_eff<1>/OD ),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\NPC_eff<1>/OFF/RST ),
    .O(DLX_IFinst_NPC_1_1)
  );
  X_OR2 \NPC_eff<1>/OFF/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\NPC_eff<1>/OFF/RST )
  );
  X_ZERO \vga_address<13>/LOGIC_ZERO_243  (
    .O(\vga_address<13>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_Madd_addressout_inst_cy_473_244 (
    .IA(\vga_address<13>/LOGIC_ZERO ),
    .IB(\vga_address<13>/CYINIT ),
    .SEL(\vga_address<13>/FROM ),
    .O(vga_top_vga1_Madd_addressout_inst_cy_473)
  );
  X_XOR2 vga_top_vga1_Madd_addressout_inst_sum_261 (
    .I0(\vga_address<13>/CYINIT ),
    .I1(\vga_address<13>/FROM ),
    .O(\vga_address<13>/XORF )
  );
  defparam \vga_address<13>/F .INIT = 16'hCCCC;
  X_LUT4 \vga_address<13>/F  (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_Mmult__n0043_inst_lut2_322),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\vga_address<13>/FROM )
  );
  defparam vga_top_vga1_Mmult__n0043_inst_lut2_323_rt_245.INIT = 16'hAAAA;
  X_LUT4 vga_top_vga1_Mmult__n0043_inst_lut2_323_rt_245 (
    .ADR0(vga_top_vga1_Mmult__n0043_inst_lut2_323),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(vga_top_vga1_Mmult__n0043_inst_lut2_323_rt)
  );
  X_BUF \vga_address<13>/XUSED  (
    .I(\vga_address<13>/XORF ),
    .O(vga_address[13])
  );
  X_BUF \vga_address<13>/YUSED  (
    .I(\vga_address<13>/XORG ),
    .O(vga_address[14])
  );
  X_XOR2 vga_top_vga1_Madd_addressout_inst_sum_262 (
    .I0(vga_top_vga1_Madd_addressout_inst_cy_473),
    .I1(vga_top_vga1_Mmult__n0043_inst_lut2_323_rt),
    .O(\vga_address<13>/XORG )
  );
  X_BUF \vga_address<13>/CYINIT_246  (
    .I(vga_top_vga1_Madd_addressout_inst_cy_472),
    .O(\vga_address<13>/CYINIT )
  );
  X_ZERO \DLX_EXinst_Mcompar__n0057_inst_cy_135/LOGIC_ZERO_247  (
    .O(\DLX_EXinst_Mcompar__n0057_inst_cy_135/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0057_inst_cy_134_248 (
    .IA(DLX_IDinst_reg_out_B[0]),
    .IB(\DLX_EXinst_Mcompar__n0057_inst_cy_135/LOGIC_ZERO ),
    .SEL(DLX_EXinst_Mcompar__n0057_inst_lut2_70),
    .O(DLX_EXinst_Mcompar__n0057_inst_cy_134)
  );
  defparam DLX_EXinst_Mcompar__n0057_inst_lut2_701.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0057_inst_lut2_701 (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(DLX_IDinst_reg_out_A[0]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0057_inst_lut2_70)
  );
  defparam DLX_EXinst_Mcompar__n0057_inst_lut2_711.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0057_inst_lut2_711 (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[1]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0057_inst_lut2_71)
  );
  X_BUF \DLX_EXinst_Mcompar__n0057_inst_cy_135/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0057_inst_cy_135/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0057_inst_cy_135)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0057_inst_cy_135_249 (
    .IA(DLX_IDinst_reg_out_B[1]),
    .IB(DLX_EXinst_Mcompar__n0057_inst_cy_134),
    .SEL(DLX_EXinst_Mcompar__n0057_inst_lut2_71),
    .O(\DLX_EXinst_Mcompar__n0057_inst_cy_135/CYMUXG )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0057_inst_cy_136_250 (
    .IA(DLX_IDinst_reg_out_B_2_1),
    .IB(\DLX_EXinst_Mcompar__n0057_inst_cy_137/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0057_inst_lut2_72),
    .O(DLX_EXinst_Mcompar__n0057_inst_cy_136)
  );
  defparam DLX_EXinst_Mcompar__n0057_inst_lut2_721.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0057_inst_lut2_721 (
    .ADR0(DLX_IDinst_reg_out_B_2_1),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[2]),
    .O(DLX_EXinst_Mcompar__n0057_inst_lut2_72)
  );
  defparam DLX_EXinst_Mcompar__n0057_inst_lut2_731.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0057_inst_lut2_731 (
    .ADR0(DLX_IDinst_reg_out_B_3_1),
    .ADR1(DLX_IDinst_reg_out_A[3]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0057_inst_lut2_73)
  );
  X_BUF \DLX_EXinst_Mcompar__n0057_inst_cy_137/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0057_inst_cy_137/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0057_inst_cy_137)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0057_inst_cy_137_251 (
    .IA(DLX_IDinst_reg_out_B_3_1),
    .IB(DLX_EXinst_Mcompar__n0057_inst_cy_136),
    .SEL(DLX_EXinst_Mcompar__n0057_inst_lut2_73),
    .O(\DLX_EXinst_Mcompar__n0057_inst_cy_137/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0057_inst_cy_137/CYINIT_252  (
    .I(DLX_EXinst_Mcompar__n0057_inst_cy_135),
    .O(\DLX_EXinst_Mcompar__n0057_inst_cy_137/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0057_inst_cy_138_253 (
    .IA(DLX_IDinst_reg_out_B[4]),
    .IB(\DLX_EXinst_Mcompar__n0057_inst_cy_139/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0057_inst_lut2_74),
    .O(DLX_EXinst_Mcompar__n0057_inst_cy_138)
  );
  defparam DLX_EXinst_Mcompar__n0057_inst_lut2_741.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0057_inst_lut2_741 (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(DLX_IDinst_reg_out_A[4]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0057_inst_lut2_74)
  );
  defparam DLX_EXinst_Mcompar__n0057_inst_lut2_751.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0057_inst_lut2_751 (
    .ADR0(DLX_IDinst_reg_out_B[5]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[5]),
    .O(DLX_EXinst_Mcompar__n0057_inst_lut2_75)
  );
  X_BUF \DLX_EXinst_Mcompar__n0057_inst_cy_139/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0057_inst_cy_139/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0057_inst_cy_139)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0057_inst_cy_139_254 (
    .IA(DLX_IDinst_reg_out_B[5]),
    .IB(DLX_EXinst_Mcompar__n0057_inst_cy_138),
    .SEL(DLX_EXinst_Mcompar__n0057_inst_lut2_75),
    .O(\DLX_EXinst_Mcompar__n0057_inst_cy_139/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0057_inst_cy_139/CYINIT_255  (
    .I(DLX_EXinst_Mcompar__n0057_inst_cy_137),
    .O(\DLX_EXinst_Mcompar__n0057_inst_cy_139/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0057_inst_cy_140_256 (
    .IA(DLX_IDinst_reg_out_B[6]),
    .IB(\DLX_EXinst_Mcompar__n0057_inst_cy_141/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0057_inst_lut2_76),
    .O(DLX_EXinst_Mcompar__n0057_inst_cy_140)
  );
  defparam DLX_EXinst_Mcompar__n0057_inst_lut2_761.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0057_inst_lut2_761 (
    .ADR0(DLX_IDinst_reg_out_B[6]),
    .ADR1(DLX_IDinst_reg_out_A[6]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0057_inst_lut2_76)
  );
  defparam DLX_EXinst_Mcompar__n0057_inst_lut2_771.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0057_inst_lut2_771 (
    .ADR0(DLX_IDinst_reg_out_B[7]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[7]),
    .O(DLX_EXinst_Mcompar__n0057_inst_lut2_77)
  );
  X_BUF \DLX_EXinst_Mcompar__n0057_inst_cy_141/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0057_inst_cy_141/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0057_inst_cy_141)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0057_inst_cy_141_257 (
    .IA(DLX_IDinst_reg_out_B[7]),
    .IB(DLX_EXinst_Mcompar__n0057_inst_cy_140),
    .SEL(DLX_EXinst_Mcompar__n0057_inst_lut2_77),
    .O(\DLX_EXinst_Mcompar__n0057_inst_cy_141/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0057_inst_cy_141/CYINIT_258  (
    .I(DLX_EXinst_Mcompar__n0057_inst_cy_139),
    .O(\DLX_EXinst_Mcompar__n0057_inst_cy_141/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0057_inst_cy_142_259 (
    .IA(DLX_IDinst_reg_out_B[8]),
    .IB(\DLX_EXinst_Mcompar__n0057_inst_cy_143/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0057_inst_lut2_78),
    .O(DLX_EXinst_Mcompar__n0057_inst_cy_142)
  );
  defparam DLX_EXinst_Mcompar__n0057_inst_lut2_781.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0057_inst_lut2_781 (
    .ADR0(DLX_IDinst_reg_out_B[8]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[8]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0057_inst_lut2_78)
  );
  defparam DLX_EXinst_Mcompar__n0057_inst_lut2_791.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0057_inst_lut2_791 (
    .ADR0(DLX_IDinst_reg_out_B[9]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[9]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0057_inst_lut2_79)
  );
  X_BUF \DLX_EXinst_Mcompar__n0057_inst_cy_143/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0057_inst_cy_143/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0057_inst_cy_143)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0057_inst_cy_143_260 (
    .IA(DLX_IDinst_reg_out_B[9]),
    .IB(DLX_EXinst_Mcompar__n0057_inst_cy_142),
    .SEL(DLX_EXinst_Mcompar__n0057_inst_lut2_79),
    .O(\DLX_EXinst_Mcompar__n0057_inst_cy_143/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0057_inst_cy_143/CYINIT_261  (
    .I(DLX_EXinst_Mcompar__n0057_inst_cy_141),
    .O(\DLX_EXinst_Mcompar__n0057_inst_cy_143/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0057_inst_cy_144_262 (
    .IA(DLX_IDinst_reg_out_B[10]),
    .IB(\DLX_EXinst_Mcompar__n0057_inst_cy_145/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0057_inst_lut2_80),
    .O(DLX_EXinst_Mcompar__n0057_inst_cy_144)
  );
  defparam DLX_EXinst_Mcompar__n0057_inst_lut2_801.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0057_inst_lut2_801 (
    .ADR0(DLX_IDinst_reg_out_B[10]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[10]),
    .O(DLX_EXinst_Mcompar__n0057_inst_lut2_80)
  );
  defparam DLX_EXinst_Mcompar__n0057_inst_lut2_811.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0057_inst_lut2_811 (
    .ADR0(DLX_IDinst_reg_out_B[11]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[11]),
    .O(DLX_EXinst_Mcompar__n0057_inst_lut2_81)
  );
  X_BUF \DLX_EXinst_Mcompar__n0057_inst_cy_145/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0057_inst_cy_145/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0057_inst_cy_145)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0057_inst_cy_145_263 (
    .IA(DLX_IDinst_reg_out_B[11]),
    .IB(DLX_EXinst_Mcompar__n0057_inst_cy_144),
    .SEL(DLX_EXinst_Mcompar__n0057_inst_lut2_81),
    .O(\DLX_EXinst_Mcompar__n0057_inst_cy_145/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0057_inst_cy_145/CYINIT_264  (
    .I(DLX_EXinst_Mcompar__n0057_inst_cy_143),
    .O(\DLX_EXinst_Mcompar__n0057_inst_cy_145/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0057_inst_cy_146_265 (
    .IA(DLX_IDinst_reg_out_B[12]),
    .IB(\DLX_EXinst_Mcompar__n0057_inst_cy_147/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0057_inst_lut2_82),
    .O(DLX_EXinst_Mcompar__n0057_inst_cy_146)
  );
  defparam DLX_EXinst_Mcompar__n0057_inst_lut2_821.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0057_inst_lut2_821 (
    .ADR0(DLX_IDinst_reg_out_B[12]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[12]),
    .O(DLX_EXinst_Mcompar__n0057_inst_lut2_82)
  );
  defparam DLX_EXinst_Mcompar__n0057_inst_lut2_831.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0057_inst_lut2_831 (
    .ADR0(DLX_IDinst_reg_out_B[13]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[13]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0057_inst_lut2_83)
  );
  X_BUF \DLX_EXinst_Mcompar__n0057_inst_cy_147/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0057_inst_cy_147/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0057_inst_cy_147)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0057_inst_cy_147_266 (
    .IA(DLX_IDinst_reg_out_B[13]),
    .IB(DLX_EXinst_Mcompar__n0057_inst_cy_146),
    .SEL(DLX_EXinst_Mcompar__n0057_inst_lut2_83),
    .O(\DLX_EXinst_Mcompar__n0057_inst_cy_147/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0057_inst_cy_147/CYINIT_267  (
    .I(DLX_EXinst_Mcompar__n0057_inst_cy_145),
    .O(\DLX_EXinst_Mcompar__n0057_inst_cy_147/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0057_inst_cy_148_268 (
    .IA(DLX_IDinst_reg_out_B[14]),
    .IB(\DLX_EXinst_Mcompar__n0057_inst_cy_149/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0057_inst_lut2_84),
    .O(DLX_EXinst_Mcompar__n0057_inst_cy_148)
  );
  defparam DLX_EXinst_Mcompar__n0057_inst_lut2_841.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0057_inst_lut2_841 (
    .ADR0(DLX_IDinst_reg_out_B[14]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[14]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0057_inst_lut2_84)
  );
  defparam DLX_EXinst_Mcompar__n0057_inst_lut2_851.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0057_inst_lut2_851 (
    .ADR0(DLX_IDinst_reg_out_B[15]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[15]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0057_inst_lut2_85)
  );
  X_BUF \DLX_EXinst_Mcompar__n0057_inst_cy_149/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0057_inst_cy_149/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0057_inst_cy_149)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0057_inst_cy_149_269 (
    .IA(DLX_IDinst_reg_out_B[15]),
    .IB(DLX_EXinst_Mcompar__n0057_inst_cy_148),
    .SEL(DLX_EXinst_Mcompar__n0057_inst_lut2_85),
    .O(\DLX_EXinst_Mcompar__n0057_inst_cy_149/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0057_inst_cy_149/CYINIT_270  (
    .I(DLX_EXinst_Mcompar__n0057_inst_cy_147),
    .O(\DLX_EXinst_Mcompar__n0057_inst_cy_149/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0057_inst_cy_150_271 (
    .IA(DLX_IDinst_reg_out_B[16]),
    .IB(\DLX_EXinst_Mcompar__n0057_inst_cy_151/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0057_inst_lut2_86),
    .O(DLX_EXinst_Mcompar__n0057_inst_cy_150)
  );
  defparam DLX_EXinst_Mcompar__n0057_inst_lut2_861.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0057_inst_lut2_861 (
    .ADR0(DLX_IDinst_reg_out_B[16]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[16]),
    .O(DLX_EXinst_Mcompar__n0057_inst_lut2_86)
  );
  defparam DLX_EXinst_Mcompar__n0057_inst_lut2_871.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0057_inst_lut2_871 (
    .ADR0(DLX_IDinst_reg_out_B[17]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[17]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0057_inst_lut2_87)
  );
  X_BUF \DLX_EXinst_Mcompar__n0057_inst_cy_151/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0057_inst_cy_151/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0057_inst_cy_151)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0057_inst_cy_151_272 (
    .IA(DLX_IDinst_reg_out_B[17]),
    .IB(DLX_EXinst_Mcompar__n0057_inst_cy_150),
    .SEL(DLX_EXinst_Mcompar__n0057_inst_lut2_87),
    .O(\DLX_EXinst_Mcompar__n0057_inst_cy_151/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0057_inst_cy_151/CYINIT_273  (
    .I(DLX_EXinst_Mcompar__n0057_inst_cy_149),
    .O(\DLX_EXinst_Mcompar__n0057_inst_cy_151/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0057_inst_cy_152_274 (
    .IA(DLX_IDinst_reg_out_B[18]),
    .IB(\DLX_EXinst_Mcompar__n0057_inst_cy_153/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0057_inst_lut2_88),
    .O(DLX_EXinst_Mcompar__n0057_inst_cy_152)
  );
  defparam DLX_EXinst_Mcompar__n0057_inst_lut2_881.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0057_inst_lut2_881 (
    .ADR0(DLX_IDinst_reg_out_B[18]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[18]),
    .O(DLX_EXinst_Mcompar__n0057_inst_lut2_88)
  );
  defparam DLX_EXinst_Mcompar__n0057_inst_lut2_891.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0057_inst_lut2_891 (
    .ADR0(DLX_IDinst_reg_out_B[19]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[19]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0057_inst_lut2_89)
  );
  X_BUF \DLX_EXinst_Mcompar__n0057_inst_cy_153/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0057_inst_cy_153/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0057_inst_cy_153)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0057_inst_cy_153_275 (
    .IA(DLX_IDinst_reg_out_B[19]),
    .IB(DLX_EXinst_Mcompar__n0057_inst_cy_152),
    .SEL(DLX_EXinst_Mcompar__n0057_inst_lut2_89),
    .O(\DLX_EXinst_Mcompar__n0057_inst_cy_153/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0057_inst_cy_153/CYINIT_276  (
    .I(DLX_EXinst_Mcompar__n0057_inst_cy_151),
    .O(\DLX_EXinst_Mcompar__n0057_inst_cy_153/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0057_inst_cy_154_277 (
    .IA(DLX_IDinst_reg_out_B[20]),
    .IB(\DLX_EXinst_Mcompar__n0057_inst_cy_155/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0057_inst_lut2_90),
    .O(DLX_EXinst_Mcompar__n0057_inst_cy_154)
  );
  defparam DLX_EXinst_Mcompar__n0057_inst_lut2_901.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0057_inst_lut2_901 (
    .ADR0(DLX_IDinst_reg_out_B[20]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[20]),
    .O(DLX_EXinst_Mcompar__n0057_inst_lut2_90)
  );
  defparam DLX_EXinst_Mcompar__n0057_inst_lut2_911.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0057_inst_lut2_911 (
    .ADR0(DLX_IDinst_reg_out_B[21]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[21]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0057_inst_lut2_91)
  );
  X_BUF \DLX_EXinst_Mcompar__n0057_inst_cy_155/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0057_inst_cy_155/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0057_inst_cy_155)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0057_inst_cy_155_278 (
    .IA(DLX_IDinst_reg_out_B[21]),
    .IB(DLX_EXinst_Mcompar__n0057_inst_cy_154),
    .SEL(DLX_EXinst_Mcompar__n0057_inst_lut2_91),
    .O(\DLX_EXinst_Mcompar__n0057_inst_cy_155/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0057_inst_cy_155/CYINIT_279  (
    .I(DLX_EXinst_Mcompar__n0057_inst_cy_153),
    .O(\DLX_EXinst_Mcompar__n0057_inst_cy_155/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0057_inst_cy_156_280 (
    .IA(DLX_IDinst_reg_out_B[22]),
    .IB(\DLX_EXinst_Mcompar__n0057_inst_cy_157/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0057_inst_lut2_92),
    .O(DLX_EXinst_Mcompar__n0057_inst_cy_156)
  );
  defparam DLX_EXinst_Mcompar__n0057_inst_lut2_921.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0057_inst_lut2_921 (
    .ADR0(DLX_IDinst_reg_out_B[22]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[22]),
    .O(DLX_EXinst_Mcompar__n0057_inst_lut2_92)
  );
  defparam DLX_EXinst_Mcompar__n0057_inst_lut2_931.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0057_inst_lut2_931 (
    .ADR0(DLX_IDinst_reg_out_B[23]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[23]),
    .O(DLX_EXinst_Mcompar__n0057_inst_lut2_93)
  );
  X_BUF \DLX_EXinst_Mcompar__n0057_inst_cy_157/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0057_inst_cy_157/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0057_inst_cy_157)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0057_inst_cy_157_281 (
    .IA(DLX_IDinst_reg_out_B[23]),
    .IB(DLX_EXinst_Mcompar__n0057_inst_cy_156),
    .SEL(DLX_EXinst_Mcompar__n0057_inst_lut2_93),
    .O(\DLX_EXinst_Mcompar__n0057_inst_cy_157/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0057_inst_cy_157/CYINIT_282  (
    .I(DLX_EXinst_Mcompar__n0057_inst_cy_155),
    .O(\DLX_EXinst_Mcompar__n0057_inst_cy_157/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0057_inst_cy_158_283 (
    .IA(DLX_IDinst_reg_out_B[24]),
    .IB(\DLX_EXinst_Mcompar__n0057_inst_cy_159/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0057_inst_lut2_94),
    .O(DLX_EXinst_Mcompar__n0057_inst_cy_158)
  );
  defparam DLX_EXinst_Mcompar__n0057_inst_lut2_941.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0057_inst_lut2_941 (
    .ADR0(DLX_IDinst_reg_out_B[24]),
    .ADR1(DLX_IDinst_reg_out_A[24]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0057_inst_lut2_94)
  );
  defparam DLX_EXinst_Mcompar__n0057_inst_lut2_951.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0057_inst_lut2_951 (
    .ADR0(DLX_IDinst_reg_out_B[25]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[25]),
    .O(DLX_EXinst_Mcompar__n0057_inst_lut2_95)
  );
  X_BUF \DLX_EXinst_Mcompar__n0057_inst_cy_159/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0057_inst_cy_159/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0057_inst_cy_159)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0057_inst_cy_159_284 (
    .IA(DLX_IDinst_reg_out_B[25]),
    .IB(DLX_EXinst_Mcompar__n0057_inst_cy_158),
    .SEL(DLX_EXinst_Mcompar__n0057_inst_lut2_95),
    .O(\DLX_EXinst_Mcompar__n0057_inst_cy_159/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0057_inst_cy_159/CYINIT_285  (
    .I(DLX_EXinst_Mcompar__n0057_inst_cy_157),
    .O(\DLX_EXinst_Mcompar__n0057_inst_cy_159/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0057_inst_cy_160_286 (
    .IA(DLX_IDinst_reg_out_B[26]),
    .IB(\DLX_EXinst_Mcompar__n0057_inst_cy_161/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0057_inst_lut2_96),
    .O(DLX_EXinst_Mcompar__n0057_inst_cy_160)
  );
  defparam DLX_EXinst_Mcompar__n0057_inst_lut2_961.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0057_inst_lut2_961 (
    .ADR0(DLX_IDinst_reg_out_B[26]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[26]),
    .O(DLX_EXinst_Mcompar__n0057_inst_lut2_96)
  );
  defparam DLX_EXinst_Mcompar__n0057_inst_lut2_971.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0057_inst_lut2_971 (
    .ADR0(DLX_IDinst_reg_out_B[27]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[27]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0057_inst_lut2_97)
  );
  X_BUF \DLX_EXinst_Mcompar__n0057_inst_cy_161/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0057_inst_cy_161/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0057_inst_cy_161)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0057_inst_cy_161_287 (
    .IA(DLX_IDinst_reg_out_B[27]),
    .IB(DLX_EXinst_Mcompar__n0057_inst_cy_160),
    .SEL(DLX_EXinst_Mcompar__n0057_inst_lut2_97),
    .O(\DLX_EXinst_Mcompar__n0057_inst_cy_161/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0057_inst_cy_161/CYINIT_288  (
    .I(DLX_EXinst_Mcompar__n0057_inst_cy_159),
    .O(\DLX_EXinst_Mcompar__n0057_inst_cy_161/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0057_inst_cy_162_289 (
    .IA(DLX_IDinst_reg_out_B[28]),
    .IB(\DLX_EXinst_Mcompar__n0057_inst_cy_163/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0057_inst_lut2_98),
    .O(DLX_EXinst_Mcompar__n0057_inst_cy_162)
  );
  defparam DLX_EXinst_Mcompar__n0057_inst_lut2_981.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0057_inst_lut2_981 (
    .ADR0(DLX_IDinst_reg_out_B[28]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[28]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0057_inst_lut2_98)
  );
  defparam DLX_EXinst_Mcompar__n0057_inst_lut2_991.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0057_inst_lut2_991 (
    .ADR0(DLX_IDinst_reg_out_B[29]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[29]),
    .O(DLX_EXinst_Mcompar__n0057_inst_lut2_99)
  );
  X_BUF \DLX_EXinst_Mcompar__n0057_inst_cy_163/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0057_inst_cy_163/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0057_inst_cy_163)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0057_inst_cy_163_290 (
    .IA(DLX_IDinst_reg_out_B[29]),
    .IB(DLX_EXinst_Mcompar__n0057_inst_cy_162),
    .SEL(DLX_EXinst_Mcompar__n0057_inst_lut2_99),
    .O(\DLX_EXinst_Mcompar__n0057_inst_cy_163/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0057_inst_cy_163/CYINIT_291  (
    .I(DLX_EXinst_Mcompar__n0057_inst_cy_161),
    .O(\DLX_EXinst_Mcompar__n0057_inst_cy_163/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0057_inst_cy_164_292 (
    .IA(DLX_IDinst_reg_out_B[30]),
    .IB(\CHOICE5306/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0057_inst_lut2_100),
    .O(\CHOICE5306/CYMUXF )
  );
  defparam DLX_EXinst_Mcompar__n0057_inst_lut2_1001.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0057_inst_lut2_1001 (
    .ADR0(DLX_IDinst_reg_out_B[30]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[30]),
    .O(DLX_EXinst_Mcompar__n0057_inst_lut2_100)
  );
  defparam \DLX_EXinst__n0006<30>253 .INIT = 16'h88A8;
  X_LUT4 \DLX_EXinst__n0006<30>253  (
    .ADR0(DLX_IDinst_reg_out_B[30]),
    .ADR1(DLX_EXinst__n0046),
    .ADR2(DLX_EXinst__n0047),
    .ADR3(DLX_IDinst_reg_out_A[30]),
    .O(\CHOICE5306/GROM )
  );
  X_BUF \CHOICE5306/XBUSED  (
    .I(\CHOICE5306/CYMUXF ),
    .O(DLX_EXinst_Mcompar__n0057_inst_cy_164)
  );
  X_BUF \CHOICE5306/YUSED  (
    .I(\CHOICE5306/GROM ),
    .O(CHOICE5306)
  );
  X_BUF \CHOICE5306/CYINIT_293  (
    .I(DLX_EXinst_Mcompar__n0057_inst_cy_163),
    .O(\CHOICE5306/CYINIT )
  );
  defparam DLX_IFinst_NPC_2_1_294.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_2_1_294 (
    .I(\NPC_eff<2>/OD ),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\NPC_eff<2>/OFF/RST ),
    .O(DLX_IFinst_NPC_2_1)
  );
  X_OR2 \NPC_eff<2>/OFF/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\NPC_eff<2>/OFF/RST )
  );
  X_ZERO \DLX_IDinst_Mcompar__n0000_inst_cy_266/LOGIC_ZERO_295  (
    .O(\DLX_IDinst_Mcompar__n0000_inst_cy_266/LOGIC_ZERO )
  );
  X_ONE \DLX_IDinst_Mcompar__n0000_inst_cy_266/LOGIC_ONE_296  (
    .O(\DLX_IDinst_Mcompar__n0000_inst_cy_266/LOGIC_ONE )
  );
  X_MUX2 DLX_IDinst_Mcompar__n0000_inst_cy_265_297 (
    .IA(\DLX_IDinst_Mcompar__n0000_inst_cy_266/LOGIC_ONE ),
    .IB(\DLX_IDinst_Mcompar__n0000_inst_cy_266/LOGIC_ZERO ),
    .SEL(DLX_IDinst_Mcompar__n0000_inst_lut4_43),
    .O(DLX_IDinst_Mcompar__n0000_inst_cy_265)
  );
  defparam DLX_IDinst_Mcompar__n0000_inst_lut4_431.INIT = 16'h8241;
  X_LUT4 DLX_IDinst_Mcompar__n0000_inst_lut4_431 (
    .ADR0(DLX_IDinst_regA_index[0]),
    .ADR1(DLX_MEMinst_reg_dst_out[1]),
    .ADR2(DLX_IDinst_regA_index[1]),
    .ADR3(DLX_MEMinst_reg_dst_out[0]),
    .O(DLX_IDinst_Mcompar__n0000_inst_lut4_43)
  );
  defparam DLX_IDinst_Mcompar__n0000_inst_lut4_441.INIT = 16'h8421;
  X_LUT4 DLX_IDinst_Mcompar__n0000_inst_lut4_441 (
    .ADR0(DLX_IDinst_regA_index[3]),
    .ADR1(DLX_MEMinst_reg_dst_out[2]),
    .ADR2(DLX_MEMinst_reg_dst_out[3]),
    .ADR3(DLX_IDinst_regA_index[2]),
    .O(DLX_IDinst_Mcompar__n0000_inst_lut4_44)
  );
  X_BUF \DLX_IDinst_Mcompar__n0000_inst_cy_266/COUTUSED  (
    .I(\DLX_IDinst_Mcompar__n0000_inst_cy_266/CYMUXG ),
    .O(DLX_IDinst_Mcompar__n0000_inst_cy_266)
  );
  X_MUX2 DLX_IDinst_Mcompar__n0000_inst_cy_266_298 (
    .IA(\DLX_IDinst_Mcompar__n0000_inst_cy_266/LOGIC_ONE ),
    .IB(DLX_IDinst_Mcompar__n0000_inst_cy_265),
    .SEL(DLX_IDinst_Mcompar__n0000_inst_lut4_44),
    .O(\DLX_IDinst_Mcompar__n0000_inst_cy_266/CYMUXG )
  );
  X_ONE \DLX_IDinst__n0000/LOGIC_ONE_299  (
    .O(\DLX_IDinst__n0000/LOGIC_ONE )
  );
  X_MUX2 DLX_IDinst_Mcompar__n0000_inst_cy_267 (
    .IA(\DLX_IDinst__n0000/LOGIC_ONE ),
    .IB(\DLX_IDinst__n0000/CYINIT ),
    .SEL(DLX_IDinst_Mcompar__n0000_inst_lut4_45),
    .O(\DLX_IDinst__n0000/CYMUXF )
  );
  defparam DLX_IDinst_Mcompar__n0000_inst_lut4_451.INIT = 16'hAA55;
  X_LUT4 DLX_IDinst_Mcompar__n0000_inst_lut4_451 (
    .ADR0(DLX_IDinst_regA_index[4]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_MEMinst_reg_dst_out[4]),
    .O(DLX_IDinst_Mcompar__n0000_inst_lut4_45)
  );
  X_BUF \DLX_IDinst__n0000/XBUSED  (
    .I(\DLX_IDinst__n0000/CYMUXF ),
    .O(DLX_IDinst__n0000)
  );
  X_BUF \DLX_IDinst__n0000/CYINIT_300  (
    .I(DLX_IDinst_Mcompar__n0000_inst_cy_266),
    .O(\DLX_IDinst__n0000/CYINIT )
  );
  X_ONE \DLX_IDinst_Mcompar__n0073_inst_cy_263/LOGIC_ONE_301  (
    .O(\DLX_IDinst_Mcompar__n0073_inst_cy_263/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mcompar__n0073_inst_cy_263/LOGIC_ZERO_302  (
    .O(\DLX_IDinst_Mcompar__n0073_inst_cy_263/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mcompar__n0073_inst_cy_262_303 (
    .IA(\DLX_IDinst_Mcompar__n0073_inst_cy_263/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mcompar__n0073_inst_cy_263/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mcompar__n0073_inst_lut4_40),
    .O(DLX_IDinst_Mcompar__n0073_inst_cy_262)
  );
  defparam DLX_IDinst_Mcompar__n0073_inst_lut4_401.INIT = 16'h8241;
  X_LUT4 DLX_IDinst_Mcompar__n0073_inst_lut4_401 (
    .ADR0(DLX_reg_dst_of_EX[1]),
    .ADR1(DLX_IDinst_regA_index[0]),
    .ADR2(DLX_reg_dst_of_EX[0]),
    .ADR3(DLX_IDinst_regA_index[1]),
    .O(DLX_IDinst_Mcompar__n0073_inst_lut4_40)
  );
  defparam DLX_IDinst_Mcompar__n0073_inst_lut4_411.INIT = 16'h8421;
  X_LUT4 DLX_IDinst_Mcompar__n0073_inst_lut4_411 (
    .ADR0(DLX_IDinst_regA_index[3]),
    .ADR1(DLX_IDinst_regA_index[2]),
    .ADR2(DLX_reg_dst_of_EX[3]),
    .ADR3(DLX_reg_dst_of_EX[2]),
    .O(DLX_IDinst_Mcompar__n0073_inst_lut4_41)
  );
  X_BUF \DLX_IDinst_Mcompar__n0073_inst_cy_263/COUTUSED  (
    .I(\DLX_IDinst_Mcompar__n0073_inst_cy_263/CYMUXG ),
    .O(DLX_IDinst_Mcompar__n0073_inst_cy_263)
  );
  X_MUX2 DLX_IDinst_Mcompar__n0073_inst_cy_263_304 (
    .IA(\DLX_IDinst_Mcompar__n0073_inst_cy_263/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mcompar__n0073_inst_cy_262),
    .SEL(DLX_IDinst_Mcompar__n0073_inst_lut4_41),
    .O(\DLX_IDinst_Mcompar__n0073_inst_cy_263/CYMUXG )
  );
  X_ZERO \DLX_reg_dst_of_MEM<4>/LOGIC_ZERO_305  (
    .O(\DLX_reg_dst_of_MEM<4>/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mcompar__n0073_inst_cy_264 (
    .IA(\DLX_reg_dst_of_MEM<4>/LOGIC_ZERO ),
    .IB(\DLX_reg_dst_of_MEM<4>/CYINIT ),
    .SEL(DLX_IDinst_Mcompar__n0073_inst_lut4_42),
    .O(\DLX_reg_dst_of_MEM<4>/CYMUXF )
  );
  defparam DLX_IDinst_Mcompar__n0073_inst_lut4_421.INIT = 16'hA5C3;
  X_LUT4 DLX_IDinst_Mcompar__n0073_inst_lut4_421 (
    .ADR0(DLX_IDinst_rd_addr[4]),
    .ADR1(DLX_IDinst_rt_addr[4]),
    .ADR2(DLX_IDinst_regA_index[4]),
    .ADR3(DLX_IDinst_reg_dst),
    .O(DLX_IDinst_Mcompar__n0073_inst_lut4_42)
  );
  defparam \DLX_Mmux_reg_dst_of_EX_Result<4>1 .INIT = 16'hFA50;
  X_LUT4 \DLX_Mmux_reg_dst_of_EX_Result<4>1  (
    .ADR0(DLX_IDinst_reg_dst),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_rt_addr[4]),
    .ADR3(DLX_IDinst_rd_addr[4]),
    .O(DLX_reg_dst_of_EX[4])
  );
  X_BUF \DLX_reg_dst_of_MEM<4>/XBUSED  (
    .I(\DLX_reg_dst_of_MEM<4>/CYMUXF ),
    .O(DLX_IDinst__n0073)
  );
  X_BUF \DLX_reg_dst_of_MEM<4>/CYINIT_306  (
    .I(DLX_IDinst_Mcompar__n0073_inst_cy_263),
    .O(\DLX_reg_dst_of_MEM<4>/CYINIT )
  );
  X_ONE \DLX_IDinst_Mcompar__n0314_inst_cy_263/LOGIC_ONE_307  (
    .O(\DLX_IDinst_Mcompar__n0314_inst_cy_263/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mcompar__n0314_inst_cy_263/LOGIC_ZERO_308  (
    .O(\DLX_IDinst_Mcompar__n0314_inst_cy_263/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mcompar__n0314_inst_cy_262_309 (
    .IA(\DLX_IDinst_Mcompar__n0314_inst_cy_263/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mcompar__n0314_inst_cy_263/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mcompar__n0314_inst_lut4_40),
    .O(DLX_IDinst_Mcompar__n0314_inst_cy_262)
  );
  defparam DLX_IDinst_Mcompar__n0314_inst_lut4_401.INIT = 16'h8421;
  X_LUT4 DLX_IDinst_Mcompar__n0314_inst_lut4_401 (
    .ADR0(DLX_MEMinst_reg_dst_out[0]),
    .ADR1(DLX_IDinst_regA_index[1]),
    .ADR2(DLX_IDinst_regA_index[0]),
    .ADR3(DLX_MEMinst_reg_dst_out[1]),
    .O(DLX_IDinst_Mcompar__n0314_inst_lut4_40)
  );
  defparam DLX_IDinst_Mcompar__n0314_inst_lut4_411.INIT = 16'h8421;
  X_LUT4 DLX_IDinst_Mcompar__n0314_inst_lut4_411 (
    .ADR0(DLX_MEMinst_reg_dst_out[3]),
    .ADR1(DLX_IDinst_regA_index[2]),
    .ADR2(DLX_IDinst_regA_index[3]),
    .ADR3(DLX_MEMinst_reg_dst_out[2]),
    .O(DLX_IDinst_Mcompar__n0314_inst_lut4_41)
  );
  X_BUF \DLX_IDinst_Mcompar__n0314_inst_cy_263/COUTUSED  (
    .I(\DLX_IDinst_Mcompar__n0314_inst_cy_263/CYMUXG ),
    .O(DLX_IDinst_Mcompar__n0314_inst_cy_263)
  );
  X_MUX2 DLX_IDinst_Mcompar__n0314_inst_cy_263_310 (
    .IA(\DLX_IDinst_Mcompar__n0314_inst_cy_263/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mcompar__n0314_inst_cy_262),
    .SEL(DLX_IDinst_Mcompar__n0314_inst_lut4_41),
    .O(\DLX_IDinst_Mcompar__n0314_inst_cy_263/CYMUXG )
  );
  X_ZERO \vga_top_vga1_Mmult__n0043_inst_lut2_317/LOGIC_ZERO_311  (
    .O(\vga_top_vga1_Mmult__n0043_inst_lut2_317/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_Mmult__n0043_inst_cy_439_312 (
    .IA(vga_top_vga1_gridvcounter[2]),
    .IB(\vga_top_vga1_Mmult__n0043_inst_lut2_317/LOGIC_ZERO ),
    .SEL(vga_top_vga1_Mmult__n0043_inst_lut2_303),
    .O(vga_top_vga1_Mmult__n0043_inst_cy_439)
  );
  defparam vga_top_vga1_Mmult__n0043_inst_lut2_3031.INIT = 16'h55AA;
  X_LUT4 vga_top_vga1_Mmult__n0043_inst_lut2_3031 (
    .ADR0(vga_top_vga1_gridvcounter[2]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_gridvcounter[0]),
    .O(vga_top_vga1_Mmult__n0043_inst_lut2_303)
  );
  defparam vga_top_vga1_Mmult__n0043_inst_lut2_3041.INIT = 16'h6666;
  X_LUT4 vga_top_vga1_Mmult__n0043_inst_lut2_3041 (
    .ADR0(vga_top_vga1_gridvcounter[3]),
    .ADR1(vga_top_vga1_gridvcounter[1]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(vga_top_vga1_Mmult__n0043_inst_lut2_304)
  );
  X_BUF \vga_top_vga1_Mmult__n0043_inst_lut2_317/COUTUSED  (
    .I(\vga_top_vga1_Mmult__n0043_inst_lut2_317/CYMUXG ),
    .O(vga_top_vga1_Mmult__n0043_inst_cy_440)
  );
  X_BUF \vga_top_vga1_Mmult__n0043_inst_lut2_317/YUSED  (
    .I(\vga_top_vga1_Mmult__n0043_inst_lut2_317/XORG ),
    .O(vga_top_vga1_Mmult__n0043_inst_lut2_317)
  );
  X_MUX2 vga_top_vga1_Mmult__n0043_inst_cy_440_313 (
    .IA(vga_top_vga1_gridvcounter[3]),
    .IB(vga_top_vga1_Mmult__n0043_inst_cy_439),
    .SEL(vga_top_vga1_Mmult__n0043_inst_lut2_304),
    .O(\vga_top_vga1_Mmult__n0043_inst_lut2_317/CYMUXG )
  );
  X_XOR2 vga_top_vga1_Mmult__n0043_inst_sum_226 (
    .I0(vga_top_vga1_Mmult__n0043_inst_cy_439),
    .I1(vga_top_vga1_Mmult__n0043_inst_lut2_304),
    .O(\vga_top_vga1_Mmult__n0043_inst_lut2_317/XORG )
  );
  X_MUX2 vga_top_vga1_Mmult__n0043_inst_cy_441_314 (
    .IA(vga_top_vga1_gridvcounter[4]),
    .IB(\vga_top_vga1_Mmult__n0043_inst_lut2_318/CYINIT ),
    .SEL(vga_top_vga1_Mmult__n0043_inst_lut2_305),
    .O(vga_top_vga1_Mmult__n0043_inst_cy_441)
  );
  X_XOR2 vga_top_vga1_Mmult__n0043_inst_sum_227 (
    .I0(\vga_top_vga1_Mmult__n0043_inst_lut2_318/CYINIT ),
    .I1(vga_top_vga1_Mmult__n0043_inst_lut2_305),
    .O(\vga_top_vga1_Mmult__n0043_inst_lut2_318/XORF )
  );
  defparam vga_top_vga1_Mmult__n0043_inst_lut2_3051.INIT = 16'h55AA;
  X_LUT4 vga_top_vga1_Mmult__n0043_inst_lut2_3051 (
    .ADR0(vga_top_vga1_gridvcounter[4]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_gridvcounter[2]),
    .O(vga_top_vga1_Mmult__n0043_inst_lut2_305)
  );
  defparam vga_top_vga1_Mmult__n0043_inst_lut2_3061.INIT = 16'h55AA;
  X_LUT4 vga_top_vga1_Mmult__n0043_inst_lut2_3061 (
    .ADR0(vga_top_vga1_gridvcounter[5]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_gridvcounter[3]),
    .O(vga_top_vga1_Mmult__n0043_inst_lut2_306)
  );
  X_BUF \vga_top_vga1_Mmult__n0043_inst_lut2_318/COUTUSED  (
    .I(\vga_top_vga1_Mmult__n0043_inst_lut2_318/CYMUXG ),
    .O(vga_top_vga1_Mmult__n0043_inst_cy_442)
  );
  X_BUF \vga_top_vga1_Mmult__n0043_inst_lut2_318/XUSED  (
    .I(\vga_top_vga1_Mmult__n0043_inst_lut2_318/XORF ),
    .O(vga_top_vga1_Mmult__n0043_inst_lut2_318)
  );
  X_BUF \vga_top_vga1_Mmult__n0043_inst_lut2_318/YUSED  (
    .I(\vga_top_vga1_Mmult__n0043_inst_lut2_318/XORG ),
    .O(vga_top_vga1_Mmult__n0043_inst_lut2_319)
  );
  X_MUX2 vga_top_vga1_Mmult__n0043_inst_cy_442_315 (
    .IA(vga_top_vga1_gridvcounter[5]),
    .IB(vga_top_vga1_Mmult__n0043_inst_cy_441),
    .SEL(vga_top_vga1_Mmult__n0043_inst_lut2_306),
    .O(\vga_top_vga1_Mmult__n0043_inst_lut2_318/CYMUXG )
  );
  X_XOR2 vga_top_vga1_Mmult__n0043_inst_sum_228 (
    .I0(vga_top_vga1_Mmult__n0043_inst_cy_441),
    .I1(vga_top_vga1_Mmult__n0043_inst_lut2_306),
    .O(\vga_top_vga1_Mmult__n0043_inst_lut2_318/XORG )
  );
  X_BUF \vga_top_vga1_Mmult__n0043_inst_lut2_318/CYINIT_316  (
    .I(vga_top_vga1_Mmult__n0043_inst_cy_440),
    .O(\vga_top_vga1_Mmult__n0043_inst_lut2_318/CYINIT )
  );
  X_MUX2 vga_top_vga1_Mmult__n0043_inst_cy_443_317 (
    .IA(vga_top_vga1_gridvcounter[6]),
    .IB(\vga_top_vga1_Mmult__n0043_inst_lut2_320/CYINIT ),
    .SEL(vga_top_vga1_Mmult__n0043_inst_lut2_307),
    .O(vga_top_vga1_Mmult__n0043_inst_cy_443)
  );
  X_XOR2 vga_top_vga1_Mmult__n0043_inst_sum_229 (
    .I0(\vga_top_vga1_Mmult__n0043_inst_lut2_320/CYINIT ),
    .I1(vga_top_vga1_Mmult__n0043_inst_lut2_307),
    .O(\vga_top_vga1_Mmult__n0043_inst_lut2_320/XORF )
  );
  defparam vga_top_vga1_Mmult__n0043_inst_lut2_3071.INIT = 16'h5A5A;
  X_LUT4 vga_top_vga1_Mmult__n0043_inst_lut2_3071 (
    .ADR0(vga_top_vga1_gridvcounter[6]),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_gridvcounter[4]),
    .ADR3(VCC),
    .O(vga_top_vga1_Mmult__n0043_inst_lut2_307)
  );
  defparam vga_top_vga1_Mmult__n0043_inst_lut2_3081.INIT = 16'h55AA;
  X_LUT4 vga_top_vga1_Mmult__n0043_inst_lut2_3081 (
    .ADR0(vga_top_vga1_gridvcounter[7]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_gridvcounter[5]),
    .O(vga_top_vga1_Mmult__n0043_inst_lut2_308)
  );
  X_BUF \vga_top_vga1_Mmult__n0043_inst_lut2_320/COUTUSED  (
    .I(\vga_top_vga1_Mmult__n0043_inst_lut2_320/CYMUXG ),
    .O(vga_top_vga1_Mmult__n0043_inst_cy_444)
  );
  X_BUF \vga_top_vga1_Mmult__n0043_inst_lut2_320/XUSED  (
    .I(\vga_top_vga1_Mmult__n0043_inst_lut2_320/XORF ),
    .O(vga_top_vga1_Mmult__n0043_inst_lut2_320)
  );
  X_BUF \vga_top_vga1_Mmult__n0043_inst_lut2_320/YUSED  (
    .I(\vga_top_vga1_Mmult__n0043_inst_lut2_320/XORG ),
    .O(vga_top_vga1_Mmult__n0043_inst_lut2_321)
  );
  X_MUX2 vga_top_vga1_Mmult__n0043_inst_cy_444_318 (
    .IA(vga_top_vga1_gridvcounter[7]),
    .IB(vga_top_vga1_Mmult__n0043_inst_cy_443),
    .SEL(vga_top_vga1_Mmult__n0043_inst_lut2_308),
    .O(\vga_top_vga1_Mmult__n0043_inst_lut2_320/CYMUXG )
  );
  X_XOR2 vga_top_vga1_Mmult__n0043_inst_sum_230 (
    .I0(vga_top_vga1_Mmult__n0043_inst_cy_443),
    .I1(vga_top_vga1_Mmult__n0043_inst_lut2_308),
    .O(\vga_top_vga1_Mmult__n0043_inst_lut2_320/XORG )
  );
  X_BUF \vga_top_vga1_Mmult__n0043_inst_lut2_320/CYINIT_319  (
    .I(vga_top_vga1_Mmult__n0043_inst_cy_442),
    .O(\vga_top_vga1_Mmult__n0043_inst_lut2_320/CYINIT )
  );
  X_MUX2 vga_top_vga1_Mmult__n0043_inst_cy_445_320 (
    .IA(vga_top_vga1_gridvcounter[8]),
    .IB(\vga_top_vga1_Mmult__n0043_inst_lut2_322/CYINIT ),
    .SEL(vga_top_vga1_Mmult__n0043_inst_lut2_309),
    .O(vga_top_vga1_Mmult__n0043_inst_cy_445)
  );
  X_XOR2 vga_top_vga1_Mmult__n0043_inst_sum_231 (
    .I0(\vga_top_vga1_Mmult__n0043_inst_lut2_322/CYINIT ),
    .I1(vga_top_vga1_Mmult__n0043_inst_lut2_309),
    .O(\vga_top_vga1_Mmult__n0043_inst_lut2_322/XORF )
  );
  defparam vga_top_vga1_Mmult__n0043_inst_lut2_3091.INIT = 16'h5A5A;
  X_LUT4 vga_top_vga1_Mmult__n0043_inst_lut2_3091 (
    .ADR0(vga_top_vga1_gridvcounter[8]),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_gridvcounter[6]),
    .ADR3(VCC),
    .O(vga_top_vga1_Mmult__n0043_inst_lut2_309)
  );
  defparam \vga_top_vga1_gridvcounter<7>_rt_321 .INIT = 16'hAAAA;
  X_LUT4 \vga_top_vga1_gridvcounter<7>_rt_321  (
    .ADR0(vga_top_vga1_gridvcounter[7]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\vga_top_vga1_gridvcounter<7>_rt )
  );
  X_BUF \vga_top_vga1_Mmult__n0043_inst_lut2_322/XUSED  (
    .I(\vga_top_vga1_Mmult__n0043_inst_lut2_322/XORF ),
    .O(vga_top_vga1_Mmult__n0043_inst_lut2_322)
  );
  X_BUF \vga_top_vga1_Mmult__n0043_inst_lut2_322/YUSED  (
    .I(\vga_top_vga1_Mmult__n0043_inst_lut2_322/XORG ),
    .O(vga_top_vga1_Mmult__n0043_inst_lut2_323)
  );
  X_XOR2 vga_top_vga1_Mmult__n0043_inst_sum_232 (
    .I0(vga_top_vga1_Mmult__n0043_inst_cy_445),
    .I1(\vga_top_vga1_gridvcounter<7>_rt ),
    .O(\vga_top_vga1_Mmult__n0043_inst_lut2_322/XORG )
  );
  X_BUF \vga_top_vga1_Mmult__n0043_inst_lut2_322/CYINIT_322  (
    .I(vga_top_vga1_Mmult__n0043_inst_cy_444),
    .O(\vga_top_vga1_Mmult__n0043_inst_lut2_322/CYINIT )
  );
  X_ZERO \DLX_EXinst_Mcompar__n0091_inst_cy_167/LOGIC_ZERO_323  (
    .O(\DLX_EXinst_Mcompar__n0091_inst_cy_167/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_166_324 (
    .IA(DLX_IDinst_reg_out_A[0]),
    .IB(\DLX_EXinst_Mcompar__n0091_inst_cy_167/LOGIC_ZERO ),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_102),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_166)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1021.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1021 (
    .ADR0(DLX_IDinst_reg_out_A[0]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_IR_function_field_0_1),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_102)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1031.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1031 (
    .ADR0(DLX_IDinst_reg_out_A[1]),
    .ADR1(DLX_IDinst_IR_function_field_1_1),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_103)
  );
  X_BUF \DLX_EXinst_Mcompar__n0091_inst_cy_167/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0091_inst_cy_167/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_167)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_167_325 (
    .IA(DLX_IDinst_reg_out_A[1]),
    .IB(DLX_EXinst_Mcompar__n0091_inst_cy_166),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_103),
    .O(\DLX_EXinst_Mcompar__n0091_inst_cy_167/CYMUXG )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_168_326 (
    .IA(DLX_IDinst_reg_out_A[2]),
    .IB(\DLX_EXinst_Mcompar__n0091_inst_cy_169/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_104),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_168)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1041.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1041 (
    .ADR0(DLX_IDinst_reg_out_A[2]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_IR_function_field_2_1),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_104)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1051.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1051 (
    .ADR0(DLX_IDinst_reg_out_A[3]),
    .ADR1(DLX_IDinst_IR_function_field_3_1),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_105)
  );
  X_BUF \DLX_EXinst_Mcompar__n0091_inst_cy_169/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0091_inst_cy_169/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_169)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_169_327 (
    .IA(DLX_IDinst_reg_out_A[3]),
    .IB(DLX_EXinst_Mcompar__n0091_inst_cy_168),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_105),
    .O(\DLX_EXinst_Mcompar__n0091_inst_cy_169/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0091_inst_cy_169/CYINIT_328  (
    .I(DLX_EXinst_Mcompar__n0091_inst_cy_167),
    .O(\DLX_EXinst_Mcompar__n0091_inst_cy_169/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_170_329 (
    .IA(DLX_IDinst_reg_out_A[4]),
    .IB(\DLX_EXinst_Mcompar__n0091_inst_cy_171/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_106),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_170)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1061.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1061 (
    .ADR0(DLX_IDinst_reg_out_A[4]),
    .ADR1(DLX_IDinst_IR_function_field[4]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_106)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1071.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1071 (
    .ADR0(DLX_IDinst_reg_out_A[5]),
    .ADR1(\DLX_IDinst_Imm[5] ),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_107)
  );
  X_BUF \DLX_EXinst_Mcompar__n0091_inst_cy_171/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0091_inst_cy_171/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_171)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_171_330 (
    .IA(DLX_IDinst_reg_out_A[5]),
    .IB(DLX_EXinst_Mcompar__n0091_inst_cy_170),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_107),
    .O(\DLX_EXinst_Mcompar__n0091_inst_cy_171/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0091_inst_cy_171/CYINIT_331  (
    .I(DLX_EXinst_Mcompar__n0091_inst_cy_169),
    .O(\DLX_EXinst_Mcompar__n0091_inst_cy_171/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_172_332 (
    .IA(DLX_IDinst_reg_out_A[6]),
    .IB(\DLX_EXinst_Mcompar__n0091_inst_cy_173/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_108),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_172)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1081.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1081 (
    .ADR0(DLX_IDinst_reg_out_A[6]),
    .ADR1(\DLX_IDinst_Imm[6] ),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_108)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1091.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1091 (
    .ADR0(DLX_IDinst_reg_out_A[7]),
    .ADR1(VCC),
    .ADR2(\DLX_IDinst_Imm[7] ),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_109)
  );
  X_BUF \DLX_EXinst_Mcompar__n0091_inst_cy_173/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0091_inst_cy_173/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_173)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_173_333 (
    .IA(DLX_IDinst_reg_out_A[7]),
    .IB(DLX_EXinst_Mcompar__n0091_inst_cy_172),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_109),
    .O(\DLX_EXinst_Mcompar__n0091_inst_cy_173/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0091_inst_cy_173/CYINIT_334  (
    .I(DLX_EXinst_Mcompar__n0091_inst_cy_171),
    .O(\DLX_EXinst_Mcompar__n0091_inst_cy_173/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_174_335 (
    .IA(DLX_IDinst_reg_out_A[8]),
    .IB(\DLX_EXinst_Mcompar__n0091_inst_cy_175/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_110),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_174)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1101.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1101 (
    .ADR0(DLX_IDinst_reg_out_A[8]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(\DLX_IDinst_Imm[8] ),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_110)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1111.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1111 (
    .ADR0(DLX_IDinst_reg_out_A[9]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(\DLX_IDinst_Imm[9] ),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_111)
  );
  X_BUF \DLX_EXinst_Mcompar__n0091_inst_cy_175/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0091_inst_cy_175/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_175)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_175_336 (
    .IA(DLX_IDinst_reg_out_A[9]),
    .IB(DLX_EXinst_Mcompar__n0091_inst_cy_174),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_111),
    .O(\DLX_EXinst_Mcompar__n0091_inst_cy_175/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0091_inst_cy_175/CYINIT_337  (
    .I(DLX_EXinst_Mcompar__n0091_inst_cy_173),
    .O(\DLX_EXinst_Mcompar__n0091_inst_cy_175/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_176_338 (
    .IA(DLX_IDinst_reg_out_A[10]),
    .IB(\DLX_EXinst_Mcompar__n0091_inst_cy_177/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_112),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_176)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1121.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1121 (
    .ADR0(DLX_IDinst_reg_out_A[10]),
    .ADR1(VCC),
    .ADR2(\DLX_IDinst_Imm[10] ),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_112)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1131.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1131 (
    .ADR0(DLX_IDinst_reg_out_A[11]),
    .ADR1(VCC),
    .ADR2(\DLX_IDinst_Imm[11] ),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_113)
  );
  X_BUF \DLX_EXinst_Mcompar__n0091_inst_cy_177/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0091_inst_cy_177/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_177)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_177_339 (
    .IA(DLX_IDinst_reg_out_A[11]),
    .IB(DLX_EXinst_Mcompar__n0091_inst_cy_176),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_113),
    .O(\DLX_EXinst_Mcompar__n0091_inst_cy_177/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0091_inst_cy_177/CYINIT_340  (
    .I(DLX_EXinst_Mcompar__n0091_inst_cy_175),
    .O(\DLX_EXinst_Mcompar__n0091_inst_cy_177/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_178_341 (
    .IA(DLX_IDinst_reg_out_A[12]),
    .IB(\DLX_EXinst_Mcompar__n0091_inst_cy_179/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_114),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_178)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1141.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1141 (
    .ADR0(DLX_IDinst_reg_out_A[12]),
    .ADR1(VCC),
    .ADR2(\DLX_IDinst_Imm[12] ),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_114)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1151.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1151 (
    .ADR0(DLX_IDinst_reg_out_A[13]),
    .ADR1(VCC),
    .ADR2(\DLX_IDinst_Imm[13] ),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_115)
  );
  X_BUF \DLX_EXinst_Mcompar__n0091_inst_cy_179/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0091_inst_cy_179/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_179)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_179_342 (
    .IA(DLX_IDinst_reg_out_A[13]),
    .IB(DLX_EXinst_Mcompar__n0091_inst_cy_178),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_115),
    .O(\DLX_EXinst_Mcompar__n0091_inst_cy_179/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0091_inst_cy_179/CYINIT_343  (
    .I(DLX_EXinst_Mcompar__n0091_inst_cy_177),
    .O(\DLX_EXinst_Mcompar__n0091_inst_cy_179/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_180_344 (
    .IA(DLX_IDinst_reg_out_A[14]),
    .IB(\DLX_EXinst_Mcompar__n0091_inst_cy_181/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_116),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_180)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1161.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1161 (
    .ADR0(DLX_IDinst_reg_out_A[14]),
    .ADR1(\DLX_IDinst_Imm[14] ),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_116)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1171.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1171 (
    .ADR0(DLX_IDinst_reg_out_A[15]),
    .ADR1(\DLX_IDinst_Imm[15] ),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_117)
  );
  X_BUF \DLX_EXinst_Mcompar__n0091_inst_cy_181/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0091_inst_cy_181/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_181)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_181_345 (
    .IA(DLX_IDinst_reg_out_A[15]),
    .IB(DLX_EXinst_Mcompar__n0091_inst_cy_180),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_117),
    .O(\DLX_EXinst_Mcompar__n0091_inst_cy_181/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0091_inst_cy_181/CYINIT_346  (
    .I(DLX_EXinst_Mcompar__n0091_inst_cy_179),
    .O(\DLX_EXinst_Mcompar__n0091_inst_cy_181/CYINIT )
  );
  defparam DLX_IFinst_NPC_3_1_347.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_3_1_347 (
    .I(\NPC_eff<3>/OD ),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\NPC_eff<3>/OFF/RST ),
    .O(DLX_IFinst_NPC_3_1)
  );
  X_OR2 \NPC_eff<3>/OFF/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\NPC_eff<3>/OFF/RST )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_182_348 (
    .IA(DLX_IDinst_reg_out_A[16]),
    .IB(\DLX_EXinst_Mcompar__n0091_inst_cy_183/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_118),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_182)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1181.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1181 (
    .ADR0(DLX_IDinst_reg_out_A[16]),
    .ADR1(DLX_IDinst_Imm_31_1),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_118)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1191.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1191 (
    .ADR0(DLX_IDinst_reg_out_A[17]),
    .ADR1(DLX_IDinst_Imm_31_1),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_119)
  );
  X_BUF \DLX_EXinst_Mcompar__n0091_inst_cy_183/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0091_inst_cy_183/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_183)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_183_349 (
    .IA(DLX_IDinst_reg_out_A[17]),
    .IB(DLX_EXinst_Mcompar__n0091_inst_cy_182),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_119),
    .O(\DLX_EXinst_Mcompar__n0091_inst_cy_183/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0091_inst_cy_183/CYINIT_350  (
    .I(DLX_EXinst_Mcompar__n0091_inst_cy_181),
    .O(\DLX_EXinst_Mcompar__n0091_inst_cy_183/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_184_351 (
    .IA(DLX_IDinst_reg_out_A[18]),
    .IB(\DLX_EXinst_Mcompar__n0091_inst_cy_185/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_120),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_184)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1201.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1201 (
    .ADR0(DLX_IDinst_reg_out_A[18]),
    .ADR1(DLX_IDinst_Imm_31_1),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_120)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1211.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1211 (
    .ADR0(DLX_IDinst_reg_out_A[19]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_Imm_31_1),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_121)
  );
  X_BUF \DLX_EXinst_Mcompar__n0091_inst_cy_185/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0091_inst_cy_185/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_185)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_185_352 (
    .IA(DLX_IDinst_reg_out_A[19]),
    .IB(DLX_EXinst_Mcompar__n0091_inst_cy_184),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_121),
    .O(\DLX_EXinst_Mcompar__n0091_inst_cy_185/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0091_inst_cy_185/CYINIT_353  (
    .I(DLX_EXinst_Mcompar__n0091_inst_cy_183),
    .O(\DLX_EXinst_Mcompar__n0091_inst_cy_185/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_186_354 (
    .IA(DLX_IDinst_reg_out_A[20]),
    .IB(\DLX_EXinst_Mcompar__n0091_inst_cy_187/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_122),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_186)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1221.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1221 (
    .ADR0(DLX_IDinst_reg_out_A[20]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_Imm_31_1),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_122)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1231.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1231 (
    .ADR0(DLX_IDinst_reg_out_A[21]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_Imm_31_1),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_123)
  );
  X_BUF \DLX_EXinst_Mcompar__n0091_inst_cy_187/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0091_inst_cy_187/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_187)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_187_355 (
    .IA(DLX_IDinst_reg_out_A[21]),
    .IB(DLX_EXinst_Mcompar__n0091_inst_cy_186),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_123),
    .O(\DLX_EXinst_Mcompar__n0091_inst_cy_187/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0091_inst_cy_187/CYINIT_356  (
    .I(DLX_EXinst_Mcompar__n0091_inst_cy_185),
    .O(\DLX_EXinst_Mcompar__n0091_inst_cy_187/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_188_357 (
    .IA(DLX_IDinst_reg_out_A[22]),
    .IB(\DLX_EXinst_Mcompar__n0091_inst_cy_189/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_124),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_188)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1241.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1241 (
    .ADR0(DLX_IDinst_reg_out_A[22]),
    .ADR1(DLX_IDinst_Imm_31_1),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_124)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1251.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1251 (
    .ADR0(DLX_IDinst_reg_out_A[23]),
    .ADR1(DLX_IDinst_Imm_31_1),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_125)
  );
  X_BUF \DLX_EXinst_Mcompar__n0091_inst_cy_189/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0091_inst_cy_189/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_189)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_189_358 (
    .IA(DLX_IDinst_reg_out_A[23]),
    .IB(DLX_EXinst_Mcompar__n0091_inst_cy_188),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_125),
    .O(\DLX_EXinst_Mcompar__n0091_inst_cy_189/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0091_inst_cy_189/CYINIT_359  (
    .I(DLX_EXinst_Mcompar__n0091_inst_cy_187),
    .O(\DLX_EXinst_Mcompar__n0091_inst_cy_189/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_190_360 (
    .IA(DLX_IDinst_reg_out_A[24]),
    .IB(\DLX_EXinst_Mcompar__n0091_inst_cy_191/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_126),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_190)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1261.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1261 (
    .ADR0(DLX_IDinst_reg_out_A[24]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_Imm_31_1),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_126)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1271.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1271 (
    .ADR0(DLX_IDinst_reg_out_A[25]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_Imm_31_1),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_127)
  );
  X_BUF \DLX_EXinst_Mcompar__n0091_inst_cy_191/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0091_inst_cy_191/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_191)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_191_361 (
    .IA(DLX_IDinst_reg_out_A[25]),
    .IB(DLX_EXinst_Mcompar__n0091_inst_cy_190),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_127),
    .O(\DLX_EXinst_Mcompar__n0091_inst_cy_191/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0091_inst_cy_191/CYINIT_362  (
    .I(DLX_EXinst_Mcompar__n0091_inst_cy_189),
    .O(\DLX_EXinst_Mcompar__n0091_inst_cy_191/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_192_363 (
    .IA(DLX_IDinst_reg_out_A[26]),
    .IB(\DLX_EXinst_Mcompar__n0091_inst_cy_193/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_128),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_192)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1281.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1281 (
    .ADR0(DLX_IDinst_reg_out_A[26]),
    .ADR1(DLX_IDinst_Imm_31_1),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_128)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1291.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1291 (
    .ADR0(DLX_IDinst_reg_out_A[27]),
    .ADR1(DLX_IDinst_Imm_31_1),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_129)
  );
  X_BUF \DLX_EXinst_Mcompar__n0091_inst_cy_193/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0091_inst_cy_193/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_193)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_193_364 (
    .IA(DLX_IDinst_reg_out_A[27]),
    .IB(DLX_EXinst_Mcompar__n0091_inst_cy_192),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_129),
    .O(\DLX_EXinst_Mcompar__n0091_inst_cy_193/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0091_inst_cy_193/CYINIT_365  (
    .I(DLX_EXinst_Mcompar__n0091_inst_cy_191),
    .O(\DLX_EXinst_Mcompar__n0091_inst_cy_193/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_194_366 (
    .IA(DLX_IDinst_reg_out_A[28]),
    .IB(\DLX_EXinst_Mcompar__n0091_inst_cy_195/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_130),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_194)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1301.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1301 (
    .ADR0(DLX_IDinst_reg_out_A[28]),
    .ADR1(DLX_IDinst_Imm_31_1),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_130)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1311.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1311 (
    .ADR0(DLX_IDinst_reg_out_A[29]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_Imm_31_1),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_131)
  );
  X_BUF \DLX_EXinst_Mcompar__n0091_inst_cy_195/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0091_inst_cy_195/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_195)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_195_367 (
    .IA(DLX_IDinst_reg_out_A[29]),
    .IB(DLX_EXinst_Mcompar__n0091_inst_cy_194),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_131),
    .O(\DLX_EXinst_Mcompar__n0091_inst_cy_195/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0091_inst_cy_195/CYINIT_368  (
    .I(DLX_EXinst_Mcompar__n0091_inst_cy_193),
    .O(\DLX_EXinst_Mcompar__n0091_inst_cy_195/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_196_369 (
    .IA(DLX_IDinst_reg_out_A[30]),
    .IB(\N127408/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_132),
    .O(\N127408/CYMUXF )
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1321.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1321 (
    .ADR0(DLX_IDinst_reg_out_A[30]),
    .ADR1(DLX_IDinst_Imm_31_1),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_132)
  );
  defparam \DLX_EXinst__n0006<30>88_SW0 .INIT = 16'h0505;
  X_LUT4 \DLX_EXinst__n0006<30>88_SW0  (
    .ADR0(DLX_IDinst_IR_opcode_field[0]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[30]),
    .ADR3(VCC),
    .O(\N127408/GROM )
  );
  X_BUF \N127408/XBUSED  (
    .I(\N127408/CYMUXF ),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_196)
  );
  X_BUF \N127408/YUSED  (
    .I(\N127408/GROM ),
    .O(N127408)
  );
  X_BUF \N127408/CYINIT_370  (
    .I(DLX_EXinst_Mcompar__n0091_inst_cy_195),
    .O(\N127408/CYINIT )
  );
  X_ZERO \DLX_EXinst_Mcompar__n0059_inst_cy_167/LOGIC_ZERO_371  (
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_167/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0059_inst_cy_166_372 (
    .IA(DLX_IDinst_reg_out_A[0]),
    .IB(\DLX_EXinst_Mcompar__n0059_inst_cy_167/LOGIC_ZERO ),
    .SEL(DLX_EXinst_Mcompar__n0059_inst_lut2_102),
    .O(DLX_EXinst_Mcompar__n0059_inst_cy_166)
  );
  defparam DLX_EXinst_Mcompar__n0059_inst_lut2_1021.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0059_inst_lut2_1021 (
    .ADR0(DLX_IDinst_reg_out_A[0]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[0]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0059_inst_lut2_102)
  );
  defparam DLX_EXinst_Mcompar__n0059_inst_lut2_1031.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0059_inst_lut2_1031 (
    .ADR0(DLX_IDinst_reg_out_A[1]),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0059_inst_lut2_103)
  );
  X_BUF \DLX_EXinst_Mcompar__n0059_inst_cy_167/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0059_inst_cy_167/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0059_inst_cy_167)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0059_inst_cy_167_373 (
    .IA(DLX_IDinst_reg_out_A[1]),
    .IB(DLX_EXinst_Mcompar__n0059_inst_cy_166),
    .SEL(DLX_EXinst_Mcompar__n0059_inst_lut2_103),
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_167/CYMUXG )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0059_inst_cy_168_374 (
    .IA(DLX_IDinst_reg_out_A[2]),
    .IB(\DLX_EXinst_Mcompar__n0059_inst_cy_169/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0059_inst_lut2_104),
    .O(DLX_EXinst_Mcompar__n0059_inst_cy_168)
  );
  defparam DLX_EXinst_Mcompar__n0059_inst_lut2_1041.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0059_inst_lut2_1041 (
    .ADR0(DLX_IDinst_reg_out_A[2]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B_2_1),
    .O(DLX_EXinst_Mcompar__n0059_inst_lut2_104)
  );
  defparam DLX_EXinst_Mcompar__n0059_inst_lut2_1051.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0059_inst_lut2_1051 (
    .ADR0(DLX_IDinst_reg_out_A[3]),
    .ADR1(DLX_IDinst_reg_out_B_3_1),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0059_inst_lut2_105)
  );
  X_BUF \DLX_EXinst_Mcompar__n0059_inst_cy_169/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0059_inst_cy_169/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0059_inst_cy_169)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0059_inst_cy_169_375 (
    .IA(DLX_IDinst_reg_out_A[3]),
    .IB(DLX_EXinst_Mcompar__n0059_inst_cy_168),
    .SEL(DLX_EXinst_Mcompar__n0059_inst_lut2_105),
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_169/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0059_inst_cy_169/CYINIT_376  (
    .I(DLX_EXinst_Mcompar__n0059_inst_cy_167),
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_169/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0059_inst_cy_170_377 (
    .IA(DLX_IDinst_reg_out_A[4]),
    .IB(\DLX_EXinst_Mcompar__n0059_inst_cy_171/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0059_inst_lut2_106),
    .O(DLX_EXinst_Mcompar__n0059_inst_cy_170)
  );
  defparam DLX_EXinst_Mcompar__n0059_inst_lut2_1061.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0059_inst_lut2_1061 (
    .ADR0(DLX_IDinst_reg_out_A[4]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[4]),
    .O(DLX_EXinst_Mcompar__n0059_inst_lut2_106)
  );
  defparam DLX_EXinst_Mcompar__n0059_inst_lut2_1071.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0059_inst_lut2_1071 (
    .ADR0(DLX_IDinst_reg_out_A[5]),
    .ADR1(DLX_IDinst_reg_out_B[5]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0059_inst_lut2_107)
  );
  X_BUF \DLX_EXinst_Mcompar__n0059_inst_cy_171/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0059_inst_cy_171/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0059_inst_cy_171)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0059_inst_cy_171_378 (
    .IA(DLX_IDinst_reg_out_A[5]),
    .IB(DLX_EXinst_Mcompar__n0059_inst_cy_170),
    .SEL(DLX_EXinst_Mcompar__n0059_inst_lut2_107),
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_171/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0059_inst_cy_171/CYINIT_379  (
    .I(DLX_EXinst_Mcompar__n0059_inst_cy_169),
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_171/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0059_inst_cy_172_380 (
    .IA(DLX_IDinst_reg_out_A[6]),
    .IB(\DLX_EXinst_Mcompar__n0059_inst_cy_173/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0059_inst_lut2_108),
    .O(DLX_EXinst_Mcompar__n0059_inst_cy_172)
  );
  defparam DLX_EXinst_Mcompar__n0059_inst_lut2_1081.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0059_inst_lut2_1081 (
    .ADR0(DLX_IDinst_reg_out_A[6]),
    .ADR1(DLX_IDinst_reg_out_B[6]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0059_inst_lut2_108)
  );
  defparam DLX_EXinst_Mcompar__n0059_inst_lut2_1091.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0059_inst_lut2_1091 (
    .ADR0(DLX_IDinst_reg_out_A[7]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[7]),
    .O(DLX_EXinst_Mcompar__n0059_inst_lut2_109)
  );
  X_BUF \DLX_EXinst_Mcompar__n0059_inst_cy_173/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0059_inst_cy_173/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0059_inst_cy_173)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0059_inst_cy_173_381 (
    .IA(DLX_IDinst_reg_out_A[7]),
    .IB(DLX_EXinst_Mcompar__n0059_inst_cy_172),
    .SEL(DLX_EXinst_Mcompar__n0059_inst_lut2_109),
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_173/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0059_inst_cy_173/CYINIT_382  (
    .I(DLX_EXinst_Mcompar__n0059_inst_cy_171),
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_173/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0059_inst_cy_174_383 (
    .IA(DLX_IDinst_reg_out_A[8]),
    .IB(\DLX_EXinst_Mcompar__n0059_inst_cy_175/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0059_inst_lut2_110),
    .O(DLX_EXinst_Mcompar__n0059_inst_cy_174)
  );
  defparam DLX_EXinst_Mcompar__n0059_inst_lut2_1101.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0059_inst_lut2_1101 (
    .ADR0(DLX_IDinst_reg_out_A[8]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[8]),
    .O(DLX_EXinst_Mcompar__n0059_inst_lut2_110)
  );
  defparam DLX_EXinst_Mcompar__n0059_inst_lut2_1111.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0059_inst_lut2_1111 (
    .ADR0(DLX_IDinst_reg_out_A[9]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[9]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0059_inst_lut2_111)
  );
  X_BUF \DLX_EXinst_Mcompar__n0059_inst_cy_175/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0059_inst_cy_175/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0059_inst_cy_175)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0059_inst_cy_175_384 (
    .IA(DLX_IDinst_reg_out_A[9]),
    .IB(DLX_EXinst_Mcompar__n0059_inst_cy_174),
    .SEL(DLX_EXinst_Mcompar__n0059_inst_lut2_111),
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_175/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0059_inst_cy_175/CYINIT_385  (
    .I(DLX_EXinst_Mcompar__n0059_inst_cy_173),
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_175/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0059_inst_cy_176_386 (
    .IA(DLX_IDinst_reg_out_A[10]),
    .IB(\DLX_EXinst_Mcompar__n0059_inst_cy_177/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0059_inst_lut2_112),
    .O(DLX_EXinst_Mcompar__n0059_inst_cy_176)
  );
  defparam DLX_EXinst_Mcompar__n0059_inst_lut2_1121.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0059_inst_lut2_1121 (
    .ADR0(DLX_IDinst_reg_out_A[10]),
    .ADR1(DLX_IDinst_reg_out_B[10]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0059_inst_lut2_112)
  );
  defparam DLX_EXinst_Mcompar__n0059_inst_lut2_1131.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0059_inst_lut2_1131 (
    .ADR0(DLX_IDinst_reg_out_A[11]),
    .ADR1(DLX_IDinst_reg_out_B[11]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0059_inst_lut2_113)
  );
  X_BUF \DLX_EXinst_Mcompar__n0059_inst_cy_177/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0059_inst_cy_177/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0059_inst_cy_177)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0059_inst_cy_177_387 (
    .IA(DLX_IDinst_reg_out_A[11]),
    .IB(DLX_EXinst_Mcompar__n0059_inst_cy_176),
    .SEL(DLX_EXinst_Mcompar__n0059_inst_lut2_113),
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_177/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0059_inst_cy_177/CYINIT_388  (
    .I(DLX_EXinst_Mcompar__n0059_inst_cy_175),
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_177/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0059_inst_cy_178_389 (
    .IA(DLX_IDinst_reg_out_A[12]),
    .IB(\DLX_EXinst_Mcompar__n0059_inst_cy_179/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0059_inst_lut2_114),
    .O(DLX_EXinst_Mcompar__n0059_inst_cy_178)
  );
  defparam DLX_EXinst_Mcompar__n0059_inst_lut2_1141.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0059_inst_lut2_1141 (
    .ADR0(DLX_IDinst_reg_out_A[12]),
    .ADR1(DLX_IDinst_reg_out_B[12]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0059_inst_lut2_114)
  );
  defparam DLX_EXinst_Mcompar__n0059_inst_lut2_1151.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0059_inst_lut2_1151 (
    .ADR0(DLX_IDinst_reg_out_A[13]),
    .ADR1(DLX_IDinst_reg_out_B[13]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0059_inst_lut2_115)
  );
  X_BUF \DLX_EXinst_Mcompar__n0059_inst_cy_179/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0059_inst_cy_179/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0059_inst_cy_179)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0059_inst_cy_179_390 (
    .IA(DLX_IDinst_reg_out_A[13]),
    .IB(DLX_EXinst_Mcompar__n0059_inst_cy_178),
    .SEL(DLX_EXinst_Mcompar__n0059_inst_lut2_115),
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_179/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0059_inst_cy_179/CYINIT_391  (
    .I(DLX_EXinst_Mcompar__n0059_inst_cy_177),
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_179/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0059_inst_cy_180_392 (
    .IA(DLX_IDinst_reg_out_A[14]),
    .IB(\DLX_EXinst_Mcompar__n0059_inst_cy_181/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0059_inst_lut2_116),
    .O(DLX_EXinst_Mcompar__n0059_inst_cy_180)
  );
  defparam DLX_EXinst_Mcompar__n0059_inst_lut2_1161.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0059_inst_lut2_1161 (
    .ADR0(DLX_IDinst_reg_out_A[14]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[14]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0059_inst_lut2_116)
  );
  defparam DLX_EXinst_Mcompar__n0059_inst_lut2_1171.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0059_inst_lut2_1171 (
    .ADR0(DLX_IDinst_reg_out_A[15]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[15]),
    .O(DLX_EXinst_Mcompar__n0059_inst_lut2_117)
  );
  X_BUF \DLX_EXinst_Mcompar__n0059_inst_cy_181/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0059_inst_cy_181/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0059_inst_cy_181)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0059_inst_cy_181_393 (
    .IA(DLX_IDinst_reg_out_A[15]),
    .IB(DLX_EXinst_Mcompar__n0059_inst_cy_180),
    .SEL(DLX_EXinst_Mcompar__n0059_inst_lut2_117),
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_181/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0059_inst_cy_181/CYINIT_394  (
    .I(DLX_EXinst_Mcompar__n0059_inst_cy_179),
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_181/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0059_inst_cy_182_395 (
    .IA(DLX_IDinst_reg_out_A[16]),
    .IB(\DLX_EXinst_Mcompar__n0059_inst_cy_183/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0059_inst_lut2_118),
    .O(DLX_EXinst_Mcompar__n0059_inst_cy_182)
  );
  defparam DLX_EXinst_Mcompar__n0059_inst_lut2_1181.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0059_inst_lut2_1181 (
    .ADR0(DLX_IDinst_reg_out_A[16]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[16]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0059_inst_lut2_118)
  );
  defparam DLX_EXinst_Mcompar__n0059_inst_lut2_1191.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0059_inst_lut2_1191 (
    .ADR0(DLX_IDinst_reg_out_A[17]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[17]),
    .O(DLX_EXinst_Mcompar__n0059_inst_lut2_119)
  );
  X_BUF \DLX_EXinst_Mcompar__n0059_inst_cy_183/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0059_inst_cy_183/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0059_inst_cy_183)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0059_inst_cy_183_396 (
    .IA(DLX_IDinst_reg_out_A[17]),
    .IB(DLX_EXinst_Mcompar__n0059_inst_cy_182),
    .SEL(DLX_EXinst_Mcompar__n0059_inst_lut2_119),
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_183/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0059_inst_cy_183/CYINIT_397  (
    .I(DLX_EXinst_Mcompar__n0059_inst_cy_181),
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_183/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0059_inst_cy_184_398 (
    .IA(DLX_IDinst_reg_out_A[18]),
    .IB(\DLX_EXinst_Mcompar__n0059_inst_cy_185/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0059_inst_lut2_120),
    .O(DLX_EXinst_Mcompar__n0059_inst_cy_184)
  );
  defparam DLX_EXinst_Mcompar__n0059_inst_lut2_1201.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0059_inst_lut2_1201 (
    .ADR0(DLX_IDinst_reg_out_A[18]),
    .ADR1(DLX_IDinst_reg_out_B[18]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0059_inst_lut2_120)
  );
  defparam DLX_EXinst_Mcompar__n0059_inst_lut2_1211.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0059_inst_lut2_1211 (
    .ADR0(DLX_IDinst_reg_out_A[19]),
    .ADR1(DLX_IDinst_reg_out_B[19]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0059_inst_lut2_121)
  );
  X_BUF \DLX_EXinst_Mcompar__n0059_inst_cy_185/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0059_inst_cy_185/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0059_inst_cy_185)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0059_inst_cy_185_399 (
    .IA(DLX_IDinst_reg_out_A[19]),
    .IB(DLX_EXinst_Mcompar__n0059_inst_cy_184),
    .SEL(DLX_EXinst_Mcompar__n0059_inst_lut2_121),
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_185/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0059_inst_cy_185/CYINIT_400  (
    .I(DLX_EXinst_Mcompar__n0059_inst_cy_183),
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_185/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0059_inst_cy_186_401 (
    .IA(DLX_IDinst_reg_out_A[20]),
    .IB(\DLX_EXinst_Mcompar__n0059_inst_cy_187/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0059_inst_lut2_122),
    .O(DLX_EXinst_Mcompar__n0059_inst_cy_186)
  );
  defparam DLX_EXinst_Mcompar__n0059_inst_lut2_1221.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0059_inst_lut2_1221 (
    .ADR0(DLX_IDinst_reg_out_A[20]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[20]),
    .O(DLX_EXinst_Mcompar__n0059_inst_lut2_122)
  );
  defparam DLX_EXinst_Mcompar__n0059_inst_lut2_1231.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0059_inst_lut2_1231 (
    .ADR0(DLX_IDinst_reg_out_A[21]),
    .ADR1(DLX_IDinst_reg_out_B[21]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0059_inst_lut2_123)
  );
  X_BUF \DLX_EXinst_Mcompar__n0059_inst_cy_187/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0059_inst_cy_187/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0059_inst_cy_187)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0059_inst_cy_187_402 (
    .IA(DLX_IDinst_reg_out_A[21]),
    .IB(DLX_EXinst_Mcompar__n0059_inst_cy_186),
    .SEL(DLX_EXinst_Mcompar__n0059_inst_lut2_123),
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_187/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0059_inst_cy_187/CYINIT_403  (
    .I(DLX_EXinst_Mcompar__n0059_inst_cy_185),
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_187/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0059_inst_cy_188_404 (
    .IA(DLX_IDinst_reg_out_A[22]),
    .IB(\DLX_EXinst_Mcompar__n0059_inst_cy_189/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0059_inst_lut2_124),
    .O(DLX_EXinst_Mcompar__n0059_inst_cy_188)
  );
  defparam DLX_EXinst_Mcompar__n0059_inst_lut2_1241.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0059_inst_lut2_1241 (
    .ADR0(DLX_IDinst_reg_out_A[22]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[22]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0059_inst_lut2_124)
  );
  defparam DLX_EXinst_Mcompar__n0059_inst_lut2_1251.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0059_inst_lut2_1251 (
    .ADR0(DLX_IDinst_reg_out_A[23]),
    .ADR1(DLX_IDinst_reg_out_B[23]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0059_inst_lut2_125)
  );
  X_BUF \DLX_EXinst_Mcompar__n0059_inst_cy_189/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0059_inst_cy_189/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0059_inst_cy_189)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0059_inst_cy_189_405 (
    .IA(DLX_IDinst_reg_out_A[23]),
    .IB(DLX_EXinst_Mcompar__n0059_inst_cy_188),
    .SEL(DLX_EXinst_Mcompar__n0059_inst_lut2_125),
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_189/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0059_inst_cy_189/CYINIT_406  (
    .I(DLX_EXinst_Mcompar__n0059_inst_cy_187),
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_189/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0059_inst_cy_190_407 (
    .IA(DLX_IDinst_reg_out_A[24]),
    .IB(\DLX_EXinst_Mcompar__n0059_inst_cy_191/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0059_inst_lut2_126),
    .O(DLX_EXinst_Mcompar__n0059_inst_cy_190)
  );
  defparam DLX_EXinst_Mcompar__n0059_inst_lut2_1261.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0059_inst_lut2_1261 (
    .ADR0(DLX_IDinst_reg_out_A[24]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[24]),
    .O(DLX_EXinst_Mcompar__n0059_inst_lut2_126)
  );
  defparam DLX_EXinst_Mcompar__n0059_inst_lut2_1271.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0059_inst_lut2_1271 (
    .ADR0(DLX_IDinst_reg_out_A[25]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[25]),
    .O(DLX_EXinst_Mcompar__n0059_inst_lut2_127)
  );
  X_BUF \DLX_EXinst_Mcompar__n0059_inst_cy_191/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0059_inst_cy_191/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0059_inst_cy_191)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0059_inst_cy_191_408 (
    .IA(DLX_IDinst_reg_out_A[25]),
    .IB(DLX_EXinst_Mcompar__n0059_inst_cy_190),
    .SEL(DLX_EXinst_Mcompar__n0059_inst_lut2_127),
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_191/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0059_inst_cy_191/CYINIT_409  (
    .I(DLX_EXinst_Mcompar__n0059_inst_cy_189),
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_191/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0059_inst_cy_192_410 (
    .IA(DLX_IDinst_reg_out_A[26]),
    .IB(\DLX_EXinst_Mcompar__n0059_inst_cy_193/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0059_inst_lut2_128),
    .O(DLX_EXinst_Mcompar__n0059_inst_cy_192)
  );
  defparam DLX_EXinst_Mcompar__n0059_inst_lut2_1281.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0059_inst_lut2_1281 (
    .ADR0(DLX_IDinst_reg_out_A[26]),
    .ADR1(DLX_IDinst_reg_out_B[26]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0059_inst_lut2_128)
  );
  defparam DLX_EXinst_Mcompar__n0059_inst_lut2_1291.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0059_inst_lut2_1291 (
    .ADR0(DLX_IDinst_reg_out_A[27]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[27]),
    .O(DLX_EXinst_Mcompar__n0059_inst_lut2_129)
  );
  X_BUF \DLX_EXinst_Mcompar__n0059_inst_cy_193/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0059_inst_cy_193/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0059_inst_cy_193)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0059_inst_cy_193_411 (
    .IA(DLX_IDinst_reg_out_A[27]),
    .IB(DLX_EXinst_Mcompar__n0059_inst_cy_192),
    .SEL(DLX_EXinst_Mcompar__n0059_inst_lut2_129),
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_193/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0059_inst_cy_193/CYINIT_412  (
    .I(DLX_EXinst_Mcompar__n0059_inst_cy_191),
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_193/CYINIT )
  );
  defparam DLX_IFinst_NPC_4_1_413.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_4_1_413 (
    .I(\NPC_eff<4>/OD ),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\NPC_eff<4>/OFF/RST ),
    .O(DLX_IFinst_NPC_4_1)
  );
  X_OR2 \NPC_eff<4>/OFF/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\NPC_eff<4>/OFF/RST )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0059_inst_cy_194_414 (
    .IA(DLX_IDinst_reg_out_A[28]),
    .IB(\DLX_EXinst_Mcompar__n0059_inst_cy_195/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0059_inst_lut2_130),
    .O(DLX_EXinst_Mcompar__n0059_inst_cy_194)
  );
  defparam DLX_EXinst_Mcompar__n0059_inst_lut2_1301.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0059_inst_lut2_1301 (
    .ADR0(DLX_IDinst_reg_out_A[28]),
    .ADR1(DLX_IDinst_reg_out_B[28]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0059_inst_lut2_130)
  );
  defparam DLX_EXinst_Mcompar__n0059_inst_lut2_1311.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0059_inst_lut2_1311 (
    .ADR0(DLX_IDinst_reg_out_A[29]),
    .ADR1(DLX_IDinst_reg_out_B[29]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0059_inst_lut2_131)
  );
  X_BUF \DLX_EXinst_Mcompar__n0059_inst_cy_195/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0059_inst_cy_195/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0059_inst_cy_195)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0059_inst_cy_195_415 (
    .IA(DLX_IDinst_reg_out_A[29]),
    .IB(DLX_EXinst_Mcompar__n0059_inst_cy_194),
    .SEL(DLX_EXinst_Mcompar__n0059_inst_lut2_131),
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_195/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0059_inst_cy_195/CYINIT_416  (
    .I(DLX_EXinst_Mcompar__n0059_inst_cy_193),
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_195/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0059_inst_cy_196_417 (
    .IA(DLX_IDinst_reg_out_A[30]),
    .IB(\CHOICE5313/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0059_inst_lut2_132),
    .O(\CHOICE5313/CYMUXF )
  );
  defparam DLX_EXinst_Mcompar__n0059_inst_lut2_1321.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0059_inst_lut2_1321 (
    .ADR0(DLX_IDinst_reg_out_A[30]),
    .ADR1(DLX_IDinst_reg_out_B[30]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0059_inst_lut2_132)
  );
  defparam \DLX_EXinst__n0006<30>275 .INIT = 16'hECEC;
  X_LUT4 \DLX_EXinst__n0006<30>275  (
    .ADR0(DLX_EXinst__n0045),
    .ADR1(DLX_EXinst_N64448),
    .ADR2(DLX_IDinst_reg_out_B[30]),
    .ADR3(VCC),
    .O(\CHOICE5313/GROM )
  );
  X_BUF \CHOICE5313/XBUSED  (
    .I(\CHOICE5313/CYMUXF ),
    .O(DLX_EXinst_Mcompar__n0059_inst_cy_196)
  );
  X_BUF \CHOICE5313/YUSED  (
    .I(\CHOICE5313/GROM ),
    .O(CHOICE5313)
  );
  X_BUF \CHOICE5313/CYINIT_418  (
    .I(DLX_EXinst_Mcompar__n0059_inst_cy_195),
    .O(\CHOICE5313/CYINIT )
  );
  X_ONE \DLX_IDinst_Mcompar__n0075_inst_cy_263/LOGIC_ONE_419  (
    .O(\DLX_IDinst_Mcompar__n0075_inst_cy_263/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mcompar__n0075_inst_cy_263/LOGIC_ZERO_420  (
    .O(\DLX_IDinst_Mcompar__n0075_inst_cy_263/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mcompar__n0075_inst_cy_262_421 (
    .IA(\DLX_IDinst_Mcompar__n0075_inst_cy_263/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mcompar__n0075_inst_cy_263/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mcompar__n0075_inst_lut4_40),
    .O(DLX_IDinst_Mcompar__n0075_inst_cy_262)
  );
  defparam DLX_IDinst_Mcompar__n0075_inst_lut4_401.INIT = 16'h9009;
  X_LUT4 DLX_IDinst_Mcompar__n0075_inst_lut4_401 (
    .ADR0(DLX_reg_dst_of_EX[1]),
    .ADR1(DLX_IDinst_regB_index[1]),
    .ADR2(DLX_reg_dst_of_EX[0]),
    .ADR3(DLX_IDinst_regB_index[0]),
    .O(DLX_IDinst_Mcompar__n0075_inst_lut4_40)
  );
  defparam DLX_IDinst_Mcompar__n0075_inst_lut4_411.INIT = 16'h9009;
  X_LUT4 DLX_IDinst_Mcompar__n0075_inst_lut4_411 (
    .ADR0(DLX_reg_dst_of_EX[3]),
    .ADR1(DLX_IDinst_regB_index[3]),
    .ADR2(DLX_IDinst_regB_index[2]),
    .ADR3(DLX_reg_dst_of_EX[2]),
    .O(DLX_IDinst_Mcompar__n0075_inst_lut4_41)
  );
  X_BUF \DLX_IDinst_Mcompar__n0075_inst_cy_263/COUTUSED  (
    .I(\DLX_IDinst_Mcompar__n0075_inst_cy_263/CYMUXG ),
    .O(DLX_IDinst_Mcompar__n0075_inst_cy_263)
  );
  X_MUX2 DLX_IDinst_Mcompar__n0075_inst_cy_263_422 (
    .IA(\DLX_IDinst_Mcompar__n0075_inst_cy_263/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mcompar__n0075_inst_cy_262),
    .SEL(DLX_IDinst_Mcompar__n0075_inst_lut4_41),
    .O(\DLX_IDinst_Mcompar__n0075_inst_cy_263/CYMUXG )
  );
  X_ZERO \DLX_EXinst_reg_dst_out<4>/LOGIC_ZERO_423  (
    .O(\DLX_EXinst_reg_dst_out<4>/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mcompar__n0075_inst_cy_264 (
    .IA(\DLX_EXinst_reg_dst_out<4>/LOGIC_ZERO ),
    .IB(\DLX_EXinst_reg_dst_out<4>/CYINIT ),
    .SEL(DLX_IDinst_Mcompar__n0075_inst_lut4_42),
    .O(\DLX_EXinst_reg_dst_out<4>/CYMUXF )
  );
  defparam DLX_IDinst_Mcompar__n0075_inst_lut4_421.INIT = 16'hC399;
  X_LUT4 DLX_IDinst_Mcompar__n0075_inst_lut4_421 (
    .ADR0(DLX_IDinst_rt_addr[4]),
    .ADR1(DLX_IDinst_regB_index[4]),
    .ADR2(DLX_IDinst_rd_addr[4]),
    .ADR3(DLX_IDinst_reg_dst),
    .O(DLX_IDinst_Mcompar__n0075_inst_lut4_42)
  );
  defparam \DLX_EXinst__n0008<4>1 .INIT = 16'hA280;
  X_LUT4 \DLX_EXinst__n0008<4>1  (
    .ADR0(DLX_EXinst__n0149),
    .ADR1(DLX_IDinst_reg_dst),
    .ADR2(DLX_IDinst_rd_addr[4]),
    .ADR3(DLX_IDinst_rt_addr[4]),
    .O(DLX_EXinst__n0008[4])
  );
  X_BUF \DLX_EXinst_reg_dst_out<4>/XBUSED  (
    .I(\DLX_EXinst_reg_dst_out<4>/CYMUXF ),
    .O(DLX_IDinst__n0075)
  );
  X_BUF \DLX_EXinst_reg_dst_out<4>/CYINIT_424  (
    .I(DLX_IDinst_Mcompar__n0075_inst_cy_263),
    .O(\DLX_EXinst_reg_dst_out<4>/CYINIT )
  );
  X_ONE \DLX_IDinst_Mcompar__n0315_inst_cy_263/LOGIC_ONE_425  (
    .O(\DLX_IDinst_Mcompar__n0315_inst_cy_263/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mcompar__n0315_inst_cy_263/LOGIC_ZERO_426  (
    .O(\DLX_IDinst_Mcompar__n0315_inst_cy_263/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mcompar__n0315_inst_cy_262_427 (
    .IA(\DLX_IDinst_Mcompar__n0315_inst_cy_263/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mcompar__n0315_inst_cy_263/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mcompar__n0315_inst_lut4_40),
    .O(DLX_IDinst_Mcompar__n0315_inst_cy_262)
  );
  defparam DLX_IDinst_Mcompar__n0315_inst_lut4_401.INIT = 16'h8421;
  X_LUT4 DLX_IDinst_Mcompar__n0315_inst_lut4_401 (
    .ADR0(DLX_MEMinst_reg_dst_out[1]),
    .ADR1(DLX_MEMinst_reg_dst_out[0]),
    .ADR2(DLX_IDinst_regB_index[1]),
    .ADR3(DLX_IDinst_regB_index[0]),
    .O(DLX_IDinst_Mcompar__n0315_inst_lut4_40)
  );
  defparam DLX_IDinst_Mcompar__n0315_inst_lut4_411.INIT = 16'h8241;
  X_LUT4 DLX_IDinst_Mcompar__n0315_inst_lut4_411 (
    .ADR0(DLX_IDinst_regB_index[2]),
    .ADR1(DLX_IDinst_regB_index[3]),
    .ADR2(DLX_MEMinst_reg_dst_out[3]),
    .ADR3(DLX_MEMinst_reg_dst_out[2]),
    .O(DLX_IDinst_Mcompar__n0315_inst_lut4_41)
  );
  X_BUF \DLX_IDinst_Mcompar__n0315_inst_cy_263/COUTUSED  (
    .I(\DLX_IDinst_Mcompar__n0315_inst_cy_263/CYMUXG ),
    .O(DLX_IDinst_Mcompar__n0315_inst_cy_263)
  );
  X_MUX2 DLX_IDinst_Mcompar__n0315_inst_cy_263_428 (
    .IA(\DLX_IDinst_Mcompar__n0315_inst_cy_263/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mcompar__n0315_inst_cy_262),
    .SEL(DLX_IDinst_Mcompar__n0315_inst_lut4_41),
    .O(\DLX_IDinst_Mcompar__n0315_inst_cy_263/CYMUXG )
  );
  X_ZERO \DLX_IDinst_Madd__n0129_inst_lut2_198/LOGIC_ZERO_429  (
    .O(\DLX_IDinst_Madd__n0129_inst_lut2_198/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Madd__n0129_inst_cy_268_430 (
    .IA(DLX_IFinst_NPC[0]),
    .IB(\DLX_IDinst_Madd__n0129_inst_lut2_198/LOGIC_ZERO ),
    .SEL(\DLX_IDinst_Madd__n0129_inst_lut2_198/FROM ),
    .O(DLX_IDinst_Madd__n0129_inst_cy_268)
  );
  defparam DLX_IDinst_Madd__n0129_inst_lut2_1981.INIT = 16'h55AA;
  X_LUT4 DLX_IDinst_Madd__n0129_inst_lut2_1981 (
    .ADR0(DLX_IFinst_NPC[0]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_jtarget[0]),
    .O(\DLX_IDinst_Madd__n0129_inst_lut2_198/FROM )
  );
  defparam DLX_IDinst_Madd__n0129_inst_lut2_1991.INIT = 16'h6666;
  X_LUT4 DLX_IDinst_Madd__n0129_inst_lut2_1991 (
    .ADR0(DLX_IFinst_NPC[1]),
    .ADR1(DLX_IDinst_jtarget[1]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Madd__n0129_inst_lut2_199)
  );
  X_BUF \DLX_IDinst_Madd__n0129_inst_lut2_198/COUTUSED  (
    .I(\DLX_IDinst_Madd__n0129_inst_lut2_198/CYMUXG ),
    .O(DLX_IDinst_Madd__n0129_inst_cy_269)
  );
  X_BUF \DLX_IDinst_Madd__n0129_inst_lut2_198/XUSED  (
    .I(\DLX_IDinst_Madd__n0129_inst_lut2_198/FROM ),
    .O(DLX_IDinst_Madd__n0129_inst_lut2_198)
  );
  X_BUF \DLX_IDinst_Madd__n0129_inst_lut2_198/YUSED  (
    .I(\DLX_IDinst_Madd__n0129_inst_lut2_198/XORG ),
    .O(DLX_IDinst__n0129[1])
  );
  X_MUX2 DLX_IDinst_Madd__n0129_inst_cy_269_431 (
    .IA(DLX_IFinst_NPC[1]),
    .IB(DLX_IDinst_Madd__n0129_inst_cy_268),
    .SEL(DLX_IDinst_Madd__n0129_inst_lut2_199),
    .O(\DLX_IDinst_Madd__n0129_inst_lut2_198/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Madd__n0129_inst_sum_103 (
    .I0(DLX_IDinst_Madd__n0129_inst_cy_268),
    .I1(DLX_IDinst_Madd__n0129_inst_lut2_199),
    .O(\DLX_IDinst_Madd__n0129_inst_lut2_198/XORG )
  );
  X_MUX2 DLX_IDinst_Madd__n0129_inst_cy_270_432 (
    .IA(DLX_IFinst_NPC[2]),
    .IB(\DLX_IDinst__n0129<2>/CYINIT ),
    .SEL(DLX_IDinst_Madd__n0129_inst_lut2_200),
    .O(DLX_IDinst_Madd__n0129_inst_cy_270)
  );
  X_XOR2 DLX_IDinst_Madd__n0129_inst_sum_104 (
    .I0(\DLX_IDinst__n0129<2>/CYINIT ),
    .I1(DLX_IDinst_Madd__n0129_inst_lut2_200),
    .O(\DLX_IDinst__n0129<2>/XORF )
  );
  defparam DLX_IDinst_Madd__n0129_inst_lut2_2001.INIT = 16'h5A5A;
  X_LUT4 DLX_IDinst_Madd__n0129_inst_lut2_2001 (
    .ADR0(DLX_IFinst_NPC[2]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_jtarget[2]),
    .ADR3(VCC),
    .O(DLX_IDinst_Madd__n0129_inst_lut2_200)
  );
  defparam DLX_IDinst_Madd__n0129_inst_lut2_2011.INIT = 16'h665A;
  X_LUT4 DLX_IDinst_Madd__n0129_inst_lut2_2011 (
    .ADR0(DLX_IFinst_NPC[3]),
    .ADR1(DLX_IFinst_IR_latched[3]),
    .ADR2(DLX_IDinst_current_IR[3]),
    .ADR3(DLX_EXinst__n0149),
    .O(DLX_IDinst_Madd__n0129_inst_lut2_201)
  );
  X_BUF \DLX_IDinst__n0129<2>/COUTUSED  (
    .I(\DLX_IDinst__n0129<2>/CYMUXG ),
    .O(DLX_IDinst_Madd__n0129_inst_cy_271)
  );
  X_BUF \DLX_IDinst__n0129<2>/XUSED  (
    .I(\DLX_IDinst__n0129<2>/XORF ),
    .O(DLX_IDinst__n0129[2])
  );
  X_BUF \DLX_IDinst__n0129<2>/YUSED  (
    .I(\DLX_IDinst__n0129<2>/XORG ),
    .O(DLX_IDinst__n0129[3])
  );
  X_MUX2 DLX_IDinst_Madd__n0129_inst_cy_271_433 (
    .IA(DLX_IFinst_NPC[3]),
    .IB(DLX_IDinst_Madd__n0129_inst_cy_270),
    .SEL(DLX_IDinst_Madd__n0129_inst_lut2_201),
    .O(\DLX_IDinst__n0129<2>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Madd__n0129_inst_sum_105 (
    .I0(DLX_IDinst_Madd__n0129_inst_cy_270),
    .I1(DLX_IDinst_Madd__n0129_inst_lut2_201),
    .O(\DLX_IDinst__n0129<2>/XORG )
  );
  X_BUF \DLX_IDinst__n0129<2>/CYINIT_434  (
    .I(DLX_IDinst_Madd__n0129_inst_cy_269),
    .O(\DLX_IDinst__n0129<2>/CYINIT )
  );
  X_MUX2 DLX_IDinst_Madd__n0129_inst_cy_272_435 (
    .IA(DLX_IFinst_NPC[4]),
    .IB(\DLX_IDinst__n0129<4>/CYINIT ),
    .SEL(DLX_IDinst_Madd__n0129_inst_lut2_202),
    .O(DLX_IDinst_Madd__n0129_inst_cy_272)
  );
  X_XOR2 DLX_IDinst_Madd__n0129_inst_sum_106 (
    .I0(\DLX_IDinst__n0129<4>/CYINIT ),
    .I1(DLX_IDinst_Madd__n0129_inst_lut2_202),
    .O(\DLX_IDinst__n0129<4>/XORF )
  );
  defparam DLX_IDinst_Madd__n0129_inst_lut2_2021.INIT = 16'h656A;
  X_LUT4 DLX_IDinst_Madd__n0129_inst_lut2_2021 (
    .ADR0(DLX_IFinst_NPC[4]),
    .ADR1(DLX_IFinst_IR_latched[4]),
    .ADR2(DLX_EXinst__n0149),
    .ADR3(DLX_IDinst_current_IR[4]),
    .O(DLX_IDinst_Madd__n0129_inst_lut2_202)
  );
  defparam DLX_IDinst_Madd__n0129_inst_lut2_2031.INIT = 16'h56A6;
  X_LUT4 DLX_IDinst_Madd__n0129_inst_lut2_2031 (
    .ADR0(DLX_IFinst_NPC[5]),
    .ADR1(DLX_IDinst_current_IR[5]),
    .ADR2(DLX_EXinst__n0149),
    .ADR3(DLX_IFinst_IR_latched[5]),
    .O(DLX_IDinst_Madd__n0129_inst_lut2_203)
  );
  X_BUF \DLX_IDinst__n0129<4>/COUTUSED  (
    .I(\DLX_IDinst__n0129<4>/CYMUXG ),
    .O(DLX_IDinst_Madd__n0129_inst_cy_273)
  );
  X_BUF \DLX_IDinst__n0129<4>/XUSED  (
    .I(\DLX_IDinst__n0129<4>/XORF ),
    .O(DLX_IDinst__n0129[4])
  );
  X_BUF \DLX_IDinst__n0129<4>/YUSED  (
    .I(\DLX_IDinst__n0129<4>/XORG ),
    .O(DLX_IDinst__n0129[5])
  );
  X_MUX2 DLX_IDinst_Madd__n0129_inst_cy_273_436 (
    .IA(DLX_IFinst_NPC[5]),
    .IB(DLX_IDinst_Madd__n0129_inst_cy_272),
    .SEL(DLX_IDinst_Madd__n0129_inst_lut2_203),
    .O(\DLX_IDinst__n0129<4>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Madd__n0129_inst_sum_107 (
    .I0(DLX_IDinst_Madd__n0129_inst_cy_272),
    .I1(DLX_IDinst_Madd__n0129_inst_lut2_203),
    .O(\DLX_IDinst__n0129<4>/XORG )
  );
  X_BUF \DLX_IDinst__n0129<4>/CYINIT_437  (
    .I(DLX_IDinst_Madd__n0129_inst_cy_271),
    .O(\DLX_IDinst__n0129<4>/CYINIT )
  );
  X_MUX2 DLX_IDinst_Madd__n0129_inst_cy_274_438 (
    .IA(DLX_IFinst_NPC[6]),
    .IB(\DLX_IDinst__n0129<6>/CYINIT ),
    .SEL(DLX_IDinst_Madd__n0129_inst_lut2_204),
    .O(DLX_IDinst_Madd__n0129_inst_cy_274)
  );
  X_XOR2 DLX_IDinst_Madd__n0129_inst_sum_108 (
    .I0(\DLX_IDinst__n0129<6>/CYINIT ),
    .I1(DLX_IDinst_Madd__n0129_inst_lut2_204),
    .O(\DLX_IDinst__n0129<6>/XORF )
  );
  defparam DLX_IDinst_Madd__n0129_inst_lut2_2041.INIT = 16'h596A;
  X_LUT4 DLX_IDinst_Madd__n0129_inst_lut2_2041 (
    .ADR0(DLX_IFinst_NPC[6]),
    .ADR1(DLX_EXinst__n0149),
    .ADR2(DLX_IFinst_IR_latched[6]),
    .ADR3(DLX_IDinst_current_IR[6]),
    .O(DLX_IDinst_Madd__n0129_inst_lut2_204)
  );
  defparam DLX_IDinst_Madd__n0129_inst_lut2_2051.INIT = 16'h596A;
  X_LUT4 DLX_IDinst_Madd__n0129_inst_lut2_2051 (
    .ADR0(DLX_IFinst_NPC[7]),
    .ADR1(DLX_EXinst__n0149),
    .ADR2(DLX_IFinst_IR_latched[7]),
    .ADR3(DLX_IDinst_current_IR[7]),
    .O(DLX_IDinst_Madd__n0129_inst_lut2_205)
  );
  X_BUF \DLX_IDinst__n0129<6>/COUTUSED  (
    .I(\DLX_IDinst__n0129<6>/CYMUXG ),
    .O(DLX_IDinst_Madd__n0129_inst_cy_275)
  );
  X_BUF \DLX_IDinst__n0129<6>/XUSED  (
    .I(\DLX_IDinst__n0129<6>/XORF ),
    .O(DLX_IDinst__n0129[6])
  );
  X_BUF \DLX_IDinst__n0129<6>/YUSED  (
    .I(\DLX_IDinst__n0129<6>/XORG ),
    .O(DLX_IDinst__n0129[7])
  );
  X_MUX2 DLX_IDinst_Madd__n0129_inst_cy_275_439 (
    .IA(DLX_IFinst_NPC[7]),
    .IB(DLX_IDinst_Madd__n0129_inst_cy_274),
    .SEL(DLX_IDinst_Madd__n0129_inst_lut2_205),
    .O(\DLX_IDinst__n0129<6>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Madd__n0129_inst_sum_109 (
    .I0(DLX_IDinst_Madd__n0129_inst_cy_274),
    .I1(DLX_IDinst_Madd__n0129_inst_lut2_205),
    .O(\DLX_IDinst__n0129<6>/XORG )
  );
  X_BUF \DLX_IDinst__n0129<6>/CYINIT_440  (
    .I(DLX_IDinst_Madd__n0129_inst_cy_273),
    .O(\DLX_IDinst__n0129<6>/CYINIT )
  );
  X_MUX2 DLX_IDinst_Madd__n0129_inst_cy_276_441 (
    .IA(DLX_IFinst_NPC[8]),
    .IB(\DLX_IDinst__n0129<8>/CYINIT ),
    .SEL(DLX_IDinst_Madd__n0129_inst_lut2_206),
    .O(DLX_IDinst_Madd__n0129_inst_cy_276)
  );
  X_XOR2 DLX_IDinst_Madd__n0129_inst_sum_110 (
    .I0(\DLX_IDinst__n0129<8>/CYINIT ),
    .I1(DLX_IDinst_Madd__n0129_inst_lut2_206),
    .O(\DLX_IDinst__n0129<8>/XORF )
  );
  defparam DLX_IDinst_Madd__n0129_inst_lut2_2061.INIT = 16'h656A;
  X_LUT4 DLX_IDinst_Madd__n0129_inst_lut2_2061 (
    .ADR0(DLX_IFinst_NPC[8]),
    .ADR1(DLX_IFinst_IR_latched[8]),
    .ADR2(DLX_EXinst__n0149),
    .ADR3(DLX_IDinst_current_IR[8]),
    .O(DLX_IDinst_Madd__n0129_inst_lut2_206)
  );
  defparam DLX_IDinst_Madd__n0129_inst_lut2_2071.INIT = 16'h665A;
  X_LUT4 DLX_IDinst_Madd__n0129_inst_lut2_2071 (
    .ADR0(DLX_IFinst_NPC[9]),
    .ADR1(DLX_IFinst_IR_latched[9]),
    .ADR2(DLX_IDinst_current_IR[9]),
    .ADR3(DLX_EXinst__n0149),
    .O(DLX_IDinst_Madd__n0129_inst_lut2_207)
  );
  X_BUF \DLX_IDinst__n0129<8>/COUTUSED  (
    .I(\DLX_IDinst__n0129<8>/CYMUXG ),
    .O(DLX_IDinst_Madd__n0129_inst_cy_277)
  );
  X_BUF \DLX_IDinst__n0129<8>/XUSED  (
    .I(\DLX_IDinst__n0129<8>/XORF ),
    .O(DLX_IDinst__n0129[8])
  );
  X_BUF \DLX_IDinst__n0129<8>/YUSED  (
    .I(\DLX_IDinst__n0129<8>/XORG ),
    .O(DLX_IDinst__n0129[9])
  );
  X_MUX2 DLX_IDinst_Madd__n0129_inst_cy_277_442 (
    .IA(DLX_IFinst_NPC[9]),
    .IB(DLX_IDinst_Madd__n0129_inst_cy_276),
    .SEL(DLX_IDinst_Madd__n0129_inst_lut2_207),
    .O(\DLX_IDinst__n0129<8>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Madd__n0129_inst_sum_111 (
    .I0(DLX_IDinst_Madd__n0129_inst_cy_276),
    .I1(DLX_IDinst_Madd__n0129_inst_lut2_207),
    .O(\DLX_IDinst__n0129<8>/XORG )
  );
  X_BUF \DLX_IDinst__n0129<8>/CYINIT_443  (
    .I(DLX_IDinst_Madd__n0129_inst_cy_275),
    .O(\DLX_IDinst__n0129<8>/CYINIT )
  );
  X_MUX2 DLX_IDinst_Madd__n0129_inst_cy_278_444 (
    .IA(DLX_IFinst_NPC[10]),
    .IB(\DLX_IDinst__n0129<10>/CYINIT ),
    .SEL(DLX_IDinst_Madd__n0129_inst_lut2_208),
    .O(DLX_IDinst_Madd__n0129_inst_cy_278)
  );
  X_XOR2 DLX_IDinst_Madd__n0129_inst_sum_112 (
    .I0(\DLX_IDinst__n0129<10>/CYINIT ),
    .I1(DLX_IDinst_Madd__n0129_inst_lut2_208),
    .O(\DLX_IDinst__n0129<10>/XORF )
  );
  defparam DLX_IDinst_Madd__n0129_inst_lut2_2081.INIT = 16'h569A;
  X_LUT4 DLX_IDinst_Madd__n0129_inst_lut2_2081 (
    .ADR0(DLX_IFinst_NPC[10]),
    .ADR1(DLX_EXinst__n0149),
    .ADR2(DLX_IDinst_current_IR[10]),
    .ADR3(DLX_IFinst_IR_latched[10]),
    .O(DLX_IDinst_Madd__n0129_inst_lut2_208)
  );
  defparam DLX_IDinst_Madd__n0129_inst_lut2_2091.INIT = 16'h656A;
  X_LUT4 DLX_IDinst_Madd__n0129_inst_lut2_2091 (
    .ADR0(DLX_IFinst_NPC[11]),
    .ADR1(DLX_IFinst_IR_latched[11]),
    .ADR2(DLX_EXinst__n0149),
    .ADR3(DLX_IDinst_current_IR[11]),
    .O(DLX_IDinst_Madd__n0129_inst_lut2_209)
  );
  X_BUF \DLX_IDinst__n0129<10>/COUTUSED  (
    .I(\DLX_IDinst__n0129<10>/CYMUXG ),
    .O(DLX_IDinst_Madd__n0129_inst_cy_279)
  );
  X_BUF \DLX_IDinst__n0129<10>/XUSED  (
    .I(\DLX_IDinst__n0129<10>/XORF ),
    .O(DLX_IDinst__n0129[10])
  );
  X_BUF \DLX_IDinst__n0129<10>/YUSED  (
    .I(\DLX_IDinst__n0129<10>/XORG ),
    .O(DLX_IDinst__n0129[11])
  );
  X_MUX2 DLX_IDinst_Madd__n0129_inst_cy_279_445 (
    .IA(DLX_IFinst_NPC[11]),
    .IB(DLX_IDinst_Madd__n0129_inst_cy_278),
    .SEL(DLX_IDinst_Madd__n0129_inst_lut2_209),
    .O(\DLX_IDinst__n0129<10>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Madd__n0129_inst_sum_113 (
    .I0(DLX_IDinst_Madd__n0129_inst_cy_278),
    .I1(DLX_IDinst_Madd__n0129_inst_lut2_209),
    .O(\DLX_IDinst__n0129<10>/XORG )
  );
  X_BUF \DLX_IDinst__n0129<10>/CYINIT_446  (
    .I(DLX_IDinst_Madd__n0129_inst_cy_277),
    .O(\DLX_IDinst__n0129<10>/CYINIT )
  );
  X_MUX2 DLX_IDinst_Madd__n0129_inst_cy_280_447 (
    .IA(DLX_IFinst_NPC[12]),
    .IB(\DLX_IDinst__n0129<12>/CYINIT ),
    .SEL(DLX_IDinst_Madd__n0129_inst_lut2_210),
    .O(DLX_IDinst_Madd__n0129_inst_cy_280)
  );
  X_XOR2 DLX_IDinst_Madd__n0129_inst_sum_114 (
    .I0(\DLX_IDinst__n0129<12>/CYINIT ),
    .I1(DLX_IDinst_Madd__n0129_inst_lut2_210),
    .O(\DLX_IDinst__n0129<12>/XORF )
  );
  defparam DLX_IDinst_Madd__n0129_inst_lut2_2101.INIT = 16'h656A;
  X_LUT4 DLX_IDinst_Madd__n0129_inst_lut2_2101 (
    .ADR0(DLX_IFinst_NPC[12]),
    .ADR1(DLX_IFinst_IR_latched[12]),
    .ADR2(DLX_EXinst__n0149),
    .ADR3(DLX_IDinst_current_IR[12]),
    .O(DLX_IDinst_Madd__n0129_inst_lut2_210)
  );
  defparam DLX_IDinst_Madd__n0129_inst_lut2_2111.INIT = 16'h5A66;
  X_LUT4 DLX_IDinst_Madd__n0129_inst_lut2_2111 (
    .ADR0(DLX_IFinst_NPC[13]),
    .ADR1(DLX_IDinst_current_IR[13]),
    .ADR2(DLX_IFinst_IR_latched[13]),
    .ADR3(DLX_EXinst__n0149),
    .O(DLX_IDinst_Madd__n0129_inst_lut2_211)
  );
  X_BUF \DLX_IDinst__n0129<12>/COUTUSED  (
    .I(\DLX_IDinst__n0129<12>/CYMUXG ),
    .O(DLX_IDinst_Madd__n0129_inst_cy_281)
  );
  X_BUF \DLX_IDinst__n0129<12>/XUSED  (
    .I(\DLX_IDinst__n0129<12>/XORF ),
    .O(DLX_IDinst__n0129[12])
  );
  X_BUF \DLX_IDinst__n0129<12>/YUSED  (
    .I(\DLX_IDinst__n0129<12>/XORG ),
    .O(DLX_IDinst__n0129[13])
  );
  X_MUX2 DLX_IDinst_Madd__n0129_inst_cy_281_448 (
    .IA(DLX_IFinst_NPC[13]),
    .IB(DLX_IDinst_Madd__n0129_inst_cy_280),
    .SEL(DLX_IDinst_Madd__n0129_inst_lut2_211),
    .O(\DLX_IDinst__n0129<12>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Madd__n0129_inst_sum_115 (
    .I0(DLX_IDinst_Madd__n0129_inst_cy_280),
    .I1(DLX_IDinst_Madd__n0129_inst_lut2_211),
    .O(\DLX_IDinst__n0129<12>/XORG )
  );
  X_BUF \DLX_IDinst__n0129<12>/CYINIT_449  (
    .I(DLX_IDinst_Madd__n0129_inst_cy_279),
    .O(\DLX_IDinst__n0129<12>/CYINIT )
  );
  defparam DLX_IFinst_NPC_5_1_450.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_5_1_450 (
    .I(\NPC_eff<5>/OD ),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\NPC_eff<5>/OFF/RST ),
    .O(DLX_IFinst_NPC_5_1)
  );
  X_OR2 \NPC_eff<5>/OFF/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\NPC_eff<5>/OFF/RST )
  );
  X_MUX2 DLX_IDinst_Madd__n0129_inst_cy_282_451 (
    .IA(DLX_IFinst_NPC[14]),
    .IB(\DLX_IDinst__n0129<14>/CYINIT ),
    .SEL(DLX_IDinst_Madd__n0129_inst_lut2_212),
    .O(DLX_IDinst_Madd__n0129_inst_cy_282)
  );
  X_XOR2 DLX_IDinst_Madd__n0129_inst_sum_116 (
    .I0(\DLX_IDinst__n0129<14>/CYINIT ),
    .I1(DLX_IDinst_Madd__n0129_inst_lut2_212),
    .O(\DLX_IDinst__n0129<14>/XORF )
  );
  defparam DLX_IDinst_Madd__n0129_inst_lut2_2121.INIT = 16'h665A;
  X_LUT4 DLX_IDinst_Madd__n0129_inst_lut2_2121 (
    .ADR0(DLX_IFinst_NPC[14]),
    .ADR1(DLX_IFinst_IR_latched[14]),
    .ADR2(DLX_IDinst_current_IR[14]),
    .ADR3(DLX_EXinst__n0149),
    .O(DLX_IDinst_Madd__n0129_inst_lut2_212)
  );
  defparam DLX_IDinst_Madd__n0129_inst_lut2_2131.INIT = 16'h656A;
  X_LUT4 DLX_IDinst_Madd__n0129_inst_lut2_2131 (
    .ADR0(DLX_IFinst_NPC[15]),
    .ADR1(DLX_IFinst_IR_latched[15]),
    .ADR2(DLX_EXinst__n0149),
    .ADR3(DLX_IDinst_current_IR[15]),
    .O(DLX_IDinst_Madd__n0129_inst_lut2_213)
  );
  X_BUF \DLX_IDinst__n0129<14>/COUTUSED  (
    .I(\DLX_IDinst__n0129<14>/CYMUXG ),
    .O(DLX_IDinst_Madd__n0129_inst_cy_283)
  );
  X_BUF \DLX_IDinst__n0129<14>/XUSED  (
    .I(\DLX_IDinst__n0129<14>/XORF ),
    .O(DLX_IDinst__n0129[14])
  );
  X_BUF \DLX_IDinst__n0129<14>/YUSED  (
    .I(\DLX_IDinst__n0129<14>/XORG ),
    .O(DLX_IDinst__n0129[15])
  );
  X_MUX2 DLX_IDinst_Madd__n0129_inst_cy_283_452 (
    .IA(DLX_IFinst_NPC[15]),
    .IB(DLX_IDinst_Madd__n0129_inst_cy_282),
    .SEL(DLX_IDinst_Madd__n0129_inst_lut2_213),
    .O(\DLX_IDinst__n0129<14>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Madd__n0129_inst_sum_117 (
    .I0(DLX_IDinst_Madd__n0129_inst_cy_282),
    .I1(DLX_IDinst_Madd__n0129_inst_lut2_213),
    .O(\DLX_IDinst__n0129<14>/XORG )
  );
  X_BUF \DLX_IDinst__n0129<14>/CYINIT_453  (
    .I(DLX_IDinst_Madd__n0129_inst_cy_281),
    .O(\DLX_IDinst__n0129<14>/CYINIT )
  );
  X_MUX2 DLX_IDinst_Madd__n0129_inst_cy_284_454 (
    .IA(DLX_IFinst_NPC[16]),
    .IB(\DLX_IDinst__n0129<16>/CYINIT ),
    .SEL(DLX_IDinst_Madd__n0129_inst_lut2_214),
    .O(DLX_IDinst_Madd__n0129_inst_cy_284)
  );
  X_XOR2 DLX_IDinst_Madd__n0129_inst_sum_118 (
    .I0(\DLX_IDinst__n0129<16>/CYINIT ),
    .I1(DLX_IDinst_Madd__n0129_inst_lut2_214),
    .O(\DLX_IDinst__n0129<16>/XORF )
  );
  defparam DLX_IDinst_Madd__n0129_inst_lut2_2141.INIT = 16'h569A;
  X_LUT4 DLX_IDinst_Madd__n0129_inst_lut2_2141 (
    .ADR0(DLX_IFinst_NPC[16]),
    .ADR1(DLX_IDinst__n0456),
    .ADR2(DLX_IDinst_jtarget[15]),
    .ADR3(DLX_IDinst_regB_index[0]),
    .O(DLX_IDinst_Madd__n0129_inst_lut2_214)
  );
  defparam DLX_IDinst_Madd__n0129_inst_lut2_2151.INIT = 16'h656A;
  X_LUT4 DLX_IDinst_Madd__n0129_inst_lut2_2151 (
    .ADR0(DLX_IFinst_NPC[17]),
    .ADR1(DLX_IDinst_regB_index[1]),
    .ADR2(DLX_IDinst__n0456),
    .ADR3(DLX_IDinst_jtarget[15]),
    .O(DLX_IDinst_Madd__n0129_inst_lut2_215)
  );
  X_BUF \DLX_IDinst__n0129<16>/COUTUSED  (
    .I(\DLX_IDinst__n0129<16>/CYMUXG ),
    .O(DLX_IDinst_Madd__n0129_inst_cy_285)
  );
  X_BUF \DLX_IDinst__n0129<16>/XUSED  (
    .I(\DLX_IDinst__n0129<16>/XORF ),
    .O(DLX_IDinst__n0129[16])
  );
  X_BUF \DLX_IDinst__n0129<16>/YUSED  (
    .I(\DLX_IDinst__n0129<16>/XORG ),
    .O(DLX_IDinst__n0129[17])
  );
  X_MUX2 DLX_IDinst_Madd__n0129_inst_cy_285_455 (
    .IA(DLX_IFinst_NPC[17]),
    .IB(DLX_IDinst_Madd__n0129_inst_cy_284),
    .SEL(DLX_IDinst_Madd__n0129_inst_lut2_215),
    .O(\DLX_IDinst__n0129<16>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Madd__n0129_inst_sum_119 (
    .I0(DLX_IDinst_Madd__n0129_inst_cy_284),
    .I1(DLX_IDinst_Madd__n0129_inst_lut2_215),
    .O(\DLX_IDinst__n0129<16>/XORG )
  );
  X_BUF \DLX_IDinst__n0129<16>/CYINIT_456  (
    .I(DLX_IDinst_Madd__n0129_inst_cy_283),
    .O(\DLX_IDinst__n0129<16>/CYINIT )
  );
  X_MUX2 DLX_IDinst_Madd__n0129_inst_cy_286_457 (
    .IA(DLX_IFinst_NPC[18]),
    .IB(\DLX_IDinst__n0129<18>/CYINIT ),
    .SEL(DLX_IDinst_Madd__n0129_inst_lut2_216),
    .O(DLX_IDinst_Madd__n0129_inst_cy_286)
  );
  X_XOR2 DLX_IDinst_Madd__n0129_inst_sum_120 (
    .I0(\DLX_IDinst__n0129<18>/CYINIT ),
    .I1(DLX_IDinst_Madd__n0129_inst_lut2_216),
    .O(\DLX_IDinst__n0129<18>/XORF )
  );
  defparam DLX_IDinst_Madd__n0129_inst_lut2_2161.INIT = 16'h56A6;
  X_LUT4 DLX_IDinst_Madd__n0129_inst_lut2_2161 (
    .ADR0(DLX_IFinst_NPC[18]),
    .ADR1(DLX_IDinst_jtarget[15]),
    .ADR2(DLX_IDinst__n0456),
    .ADR3(DLX_IDinst_regB_index[2]),
    .O(DLX_IDinst_Madd__n0129_inst_lut2_216)
  );
  defparam DLX_IDinst_Madd__n0129_inst_lut2_2171.INIT = 16'h56A6;
  X_LUT4 DLX_IDinst_Madd__n0129_inst_lut2_2171 (
    .ADR0(DLX_IFinst_NPC[19]),
    .ADR1(DLX_IDinst_jtarget[15]),
    .ADR2(DLX_IDinst__n0456),
    .ADR3(DLX_IDinst_regB_index[3]),
    .O(DLX_IDinst_Madd__n0129_inst_lut2_217)
  );
  X_BUF \DLX_IDinst__n0129<18>/COUTUSED  (
    .I(\DLX_IDinst__n0129<18>/CYMUXG ),
    .O(DLX_IDinst_Madd__n0129_inst_cy_287)
  );
  X_BUF \DLX_IDinst__n0129<18>/XUSED  (
    .I(\DLX_IDinst__n0129<18>/XORF ),
    .O(DLX_IDinst__n0129[18])
  );
  X_BUF \DLX_IDinst__n0129<18>/YUSED  (
    .I(\DLX_IDinst__n0129<18>/XORG ),
    .O(DLX_IDinst__n0129[19])
  );
  X_MUX2 DLX_IDinst_Madd__n0129_inst_cy_287_458 (
    .IA(DLX_IFinst_NPC[19]),
    .IB(DLX_IDinst_Madd__n0129_inst_cy_286),
    .SEL(DLX_IDinst_Madd__n0129_inst_lut2_217),
    .O(\DLX_IDinst__n0129<18>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Madd__n0129_inst_sum_121 (
    .I0(DLX_IDinst_Madd__n0129_inst_cy_286),
    .I1(DLX_IDinst_Madd__n0129_inst_lut2_217),
    .O(\DLX_IDinst__n0129<18>/XORG )
  );
  X_BUF \DLX_IDinst__n0129<18>/CYINIT_459  (
    .I(DLX_IDinst_Madd__n0129_inst_cy_285),
    .O(\DLX_IDinst__n0129<18>/CYINIT )
  );
  X_MUX2 DLX_IDinst_Madd__n0129_inst_cy_288_460 (
    .IA(DLX_IFinst_NPC[20]),
    .IB(\DLX_IDinst__n0129<20>/CYINIT ),
    .SEL(DLX_IDinst_Madd__n0129_inst_lut2_218),
    .O(DLX_IDinst_Madd__n0129_inst_cy_288)
  );
  X_XOR2 DLX_IDinst_Madd__n0129_inst_sum_122 (
    .I0(\DLX_IDinst__n0129<20>/CYINIT ),
    .I1(DLX_IDinst_Madd__n0129_inst_lut2_218),
    .O(\DLX_IDinst__n0129<20>/XORF )
  );
  defparam DLX_IDinst_Madd__n0129_inst_lut2_2181.INIT = 16'h656A;
  X_LUT4 DLX_IDinst_Madd__n0129_inst_lut2_2181 (
    .ADR0(DLX_IFinst_NPC[20]),
    .ADR1(DLX_IDinst_regB_index[4]),
    .ADR2(DLX_IDinst__n0456),
    .ADR3(DLX_IDinst_jtarget[15]),
    .O(DLX_IDinst_Madd__n0129_inst_lut2_218)
  );
  defparam DLX_IDinst_Madd__n0129_inst_lut2_2191.INIT = 16'h656A;
  X_LUT4 DLX_IDinst_Madd__n0129_inst_lut2_2191 (
    .ADR0(DLX_IFinst_NPC[21]),
    .ADR1(DLX_IDinst_regA_index[0]),
    .ADR2(DLX_IDinst__n0456),
    .ADR3(DLX_IDinst_jtarget[15]),
    .O(DLX_IDinst_Madd__n0129_inst_lut2_219)
  );
  X_BUF \DLX_IDinst__n0129<20>/COUTUSED  (
    .I(\DLX_IDinst__n0129<20>/CYMUXG ),
    .O(DLX_IDinst_Madd__n0129_inst_cy_289)
  );
  X_BUF \DLX_IDinst__n0129<20>/XUSED  (
    .I(\DLX_IDinst__n0129<20>/XORF ),
    .O(DLX_IDinst__n0129[20])
  );
  X_BUF \DLX_IDinst__n0129<20>/YUSED  (
    .I(\DLX_IDinst__n0129<20>/XORG ),
    .O(DLX_IDinst__n0129[21])
  );
  X_MUX2 DLX_IDinst_Madd__n0129_inst_cy_289_461 (
    .IA(DLX_IFinst_NPC[21]),
    .IB(DLX_IDinst_Madd__n0129_inst_cy_288),
    .SEL(DLX_IDinst_Madd__n0129_inst_lut2_219),
    .O(\DLX_IDinst__n0129<20>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Madd__n0129_inst_sum_123 (
    .I0(DLX_IDinst_Madd__n0129_inst_cy_288),
    .I1(DLX_IDinst_Madd__n0129_inst_lut2_219),
    .O(\DLX_IDinst__n0129<20>/XORG )
  );
  X_BUF \DLX_IDinst__n0129<20>/CYINIT_462  (
    .I(DLX_IDinst_Madd__n0129_inst_cy_287),
    .O(\DLX_IDinst__n0129<20>/CYINIT )
  );
  X_MUX2 DLX_IDinst_Madd__n0129_inst_cy_290_463 (
    .IA(DLX_IFinst_NPC[22]),
    .IB(\DLX_IDinst__n0129<22>/CYINIT ),
    .SEL(DLX_IDinst_Madd__n0129_inst_lut2_220),
    .O(DLX_IDinst_Madd__n0129_inst_cy_290)
  );
  X_XOR2 DLX_IDinst_Madd__n0129_inst_sum_124 (
    .I0(\DLX_IDinst__n0129<22>/CYINIT ),
    .I1(DLX_IDinst_Madd__n0129_inst_lut2_220),
    .O(\DLX_IDinst__n0129<22>/XORF )
  );
  defparam DLX_IDinst_Madd__n0129_inst_lut2_2201.INIT = 16'h656A;
  X_LUT4 DLX_IDinst_Madd__n0129_inst_lut2_2201 (
    .ADR0(DLX_IFinst_NPC[22]),
    .ADR1(DLX_IDinst_regA_index[1]),
    .ADR2(DLX_IDinst__n0456),
    .ADR3(DLX_IDinst_jtarget[15]),
    .O(DLX_IDinst_Madd__n0129_inst_lut2_220)
  );
  defparam DLX_IDinst_Madd__n0129_inst_lut2_2211.INIT = 16'h656A;
  X_LUT4 DLX_IDinst_Madd__n0129_inst_lut2_2211 (
    .ADR0(DLX_IFinst_NPC[23]),
    .ADR1(DLX_IDinst_regA_index[2]),
    .ADR2(DLX_IDinst__n0456),
    .ADR3(DLX_IDinst_jtarget[15]),
    .O(DLX_IDinst_Madd__n0129_inst_lut2_221)
  );
  X_BUF \DLX_IDinst__n0129<22>/COUTUSED  (
    .I(\DLX_IDinst__n0129<22>/CYMUXG ),
    .O(DLX_IDinst_Madd__n0129_inst_cy_291)
  );
  X_BUF \DLX_IDinst__n0129<22>/XUSED  (
    .I(\DLX_IDinst__n0129<22>/XORF ),
    .O(DLX_IDinst__n0129[22])
  );
  X_BUF \DLX_IDinst__n0129<22>/YUSED  (
    .I(\DLX_IDinst__n0129<22>/XORG ),
    .O(DLX_IDinst__n0129[23])
  );
  X_MUX2 DLX_IDinst_Madd__n0129_inst_cy_291_464 (
    .IA(DLX_IFinst_NPC[23]),
    .IB(DLX_IDinst_Madd__n0129_inst_cy_290),
    .SEL(DLX_IDinst_Madd__n0129_inst_lut2_221),
    .O(\DLX_IDinst__n0129<22>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Madd__n0129_inst_sum_125 (
    .I0(DLX_IDinst_Madd__n0129_inst_cy_290),
    .I1(DLX_IDinst_Madd__n0129_inst_lut2_221),
    .O(\DLX_IDinst__n0129<22>/XORG )
  );
  X_BUF \DLX_IDinst__n0129<22>/CYINIT_465  (
    .I(DLX_IDinst_Madd__n0129_inst_cy_289),
    .O(\DLX_IDinst__n0129<22>/CYINIT )
  );
  X_MUX2 DLX_IDinst_Madd__n0129_inst_cy_292_466 (
    .IA(DLX_IFinst_NPC[24]),
    .IB(\DLX_IDinst__n0129<24>/CYINIT ),
    .SEL(DLX_IDinst_Madd__n0129_inst_lut2_222),
    .O(DLX_IDinst_Madd__n0129_inst_cy_292)
  );
  X_XOR2 DLX_IDinst_Madd__n0129_inst_sum_126 (
    .I0(\DLX_IDinst__n0129<24>/CYINIT ),
    .I1(DLX_IDinst_Madd__n0129_inst_lut2_222),
    .O(\DLX_IDinst__n0129<24>/XORF )
  );
  defparam DLX_IDinst_Madd__n0129_inst_lut2_2221.INIT = 16'h5A66;
  X_LUT4 DLX_IDinst_Madd__n0129_inst_lut2_2221 (
    .ADR0(DLX_IFinst_NPC[24]),
    .ADR1(DLX_IDinst_jtarget[15]),
    .ADR2(DLX_IDinst_regA_index[3]),
    .ADR3(DLX_IDinst__n0456),
    .O(DLX_IDinst_Madd__n0129_inst_lut2_222)
  );
  defparam DLX_IDinst_Madd__n0129_inst_lut2_2231.INIT = 16'h656A;
  X_LUT4 DLX_IDinst_Madd__n0129_inst_lut2_2231 (
    .ADR0(DLX_IFinst_NPC[25]),
    .ADR1(DLX_IDinst_regA_index[4]),
    .ADR2(DLX_IDinst__n0456),
    .ADR3(DLX_IDinst_jtarget[15]),
    .O(DLX_IDinst_Madd__n0129_inst_lut2_223)
  );
  X_BUF \DLX_IDinst__n0129<24>/COUTUSED  (
    .I(\DLX_IDinst__n0129<24>/CYMUXG ),
    .O(DLX_IDinst_Madd__n0129_inst_cy_293)
  );
  X_BUF \DLX_IDinst__n0129<24>/XUSED  (
    .I(\DLX_IDinst__n0129<24>/XORF ),
    .O(DLX_IDinst__n0129[24])
  );
  X_BUF \DLX_IDinst__n0129<24>/YUSED  (
    .I(\DLX_IDinst__n0129<24>/XORG ),
    .O(DLX_IDinst__n0129[25])
  );
  X_MUX2 DLX_IDinst_Madd__n0129_inst_cy_293_467 (
    .IA(DLX_IFinst_NPC[25]),
    .IB(DLX_IDinst_Madd__n0129_inst_cy_292),
    .SEL(DLX_IDinst_Madd__n0129_inst_lut2_223),
    .O(\DLX_IDinst__n0129<24>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Madd__n0129_inst_sum_127 (
    .I0(DLX_IDinst_Madd__n0129_inst_cy_292),
    .I1(DLX_IDinst_Madd__n0129_inst_lut2_223),
    .O(\DLX_IDinst__n0129<24>/XORG )
  );
  X_BUF \DLX_IDinst__n0129<24>/CYINIT_468  (
    .I(DLX_IDinst_Madd__n0129_inst_cy_291),
    .O(\DLX_IDinst__n0129<24>/CYINIT )
  );
  X_MUX2 DLX_IDinst_Madd__n0129_inst_cy_294_469 (
    .IA(DLX_IFinst_NPC[26]),
    .IB(\DLX_IDinst__n0129<26>/CYINIT ),
    .SEL(DLX_IDinst_Madd__n0129_inst_lut2_224),
    .O(DLX_IDinst_Madd__n0129_inst_cy_294)
  );
  X_XOR2 DLX_IDinst_Madd__n0129_inst_sum_128 (
    .I0(\DLX_IDinst__n0129<26>/CYINIT ),
    .I1(DLX_IDinst_Madd__n0129_inst_lut2_224),
    .O(\DLX_IDinst__n0129<26>/XORF )
  );
  defparam DLX_IDinst_Madd__n0129_inst_lut2_2241.INIT = 16'h596A;
  X_LUT4 DLX_IDinst_Madd__n0129_inst_lut2_2241 (
    .ADR0(DLX_IFinst_NPC[26]),
    .ADR1(DLX_IDinst__n0456),
    .ADR2(DLX_IDinst_regA_index[4]),
    .ADR3(DLX_IDinst_jtarget[15]),
    .O(DLX_IDinst_Madd__n0129_inst_lut2_224)
  );
  defparam DLX_IDinst_Madd__n0129_inst_lut2_2251.INIT = 16'h656A;
  X_LUT4 DLX_IDinst_Madd__n0129_inst_lut2_2251 (
    .ADR0(DLX_IFinst_NPC[27]),
    .ADR1(DLX_IDinst_regA_index[4]),
    .ADR2(DLX_IDinst__n0456),
    .ADR3(DLX_IDinst_jtarget[15]),
    .O(DLX_IDinst_Madd__n0129_inst_lut2_225)
  );
  X_BUF \DLX_IDinst__n0129<26>/COUTUSED  (
    .I(\DLX_IDinst__n0129<26>/CYMUXG ),
    .O(DLX_IDinst_Madd__n0129_inst_cy_295)
  );
  X_BUF \DLX_IDinst__n0129<26>/XUSED  (
    .I(\DLX_IDinst__n0129<26>/XORF ),
    .O(DLX_IDinst__n0129[26])
  );
  X_BUF \DLX_IDinst__n0129<26>/YUSED  (
    .I(\DLX_IDinst__n0129<26>/XORG ),
    .O(DLX_IDinst__n0129[27])
  );
  X_MUX2 DLX_IDinst_Madd__n0129_inst_cy_295_470 (
    .IA(DLX_IFinst_NPC[27]),
    .IB(DLX_IDinst_Madd__n0129_inst_cy_294),
    .SEL(DLX_IDinst_Madd__n0129_inst_lut2_225),
    .O(\DLX_IDinst__n0129<26>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Madd__n0129_inst_sum_129 (
    .I0(DLX_IDinst_Madd__n0129_inst_cy_294),
    .I1(DLX_IDinst_Madd__n0129_inst_lut2_225),
    .O(\DLX_IDinst__n0129<26>/XORG )
  );
  X_BUF \DLX_IDinst__n0129<26>/CYINIT_471  (
    .I(DLX_IDinst_Madd__n0129_inst_cy_293),
    .O(\DLX_IDinst__n0129<26>/CYINIT )
  );
  X_MUX2 DLX_IDinst_Madd__n0129_inst_cy_296_472 (
    .IA(DLX_IFinst_NPC[28]),
    .IB(\DLX_IDinst__n0129<28>/CYINIT ),
    .SEL(DLX_IDinst_Madd__n0129_inst_lut2_226),
    .O(DLX_IDinst_Madd__n0129_inst_cy_296)
  );
  X_XOR2 DLX_IDinst_Madd__n0129_inst_sum_130 (
    .I0(\DLX_IDinst__n0129<28>/CYINIT ),
    .I1(DLX_IDinst_Madd__n0129_inst_lut2_226),
    .O(\DLX_IDinst__n0129<28>/XORF )
  );
  defparam DLX_IDinst_Madd__n0129_inst_lut2_2261.INIT = 16'h656A;
  X_LUT4 DLX_IDinst_Madd__n0129_inst_lut2_2261 (
    .ADR0(DLX_IFinst_NPC[28]),
    .ADR1(DLX_IDinst_regA_index[4]),
    .ADR2(DLX_IDinst__n0456),
    .ADR3(DLX_IDinst_jtarget[15]),
    .O(DLX_IDinst_Madd__n0129_inst_lut2_226)
  );
  defparam DLX_IDinst_Madd__n0129_inst_lut2_2271.INIT = 16'h656A;
  X_LUT4 DLX_IDinst_Madd__n0129_inst_lut2_2271 (
    .ADR0(DLX_IFinst_NPC[29]),
    .ADR1(DLX_IDinst_regA_index[4]),
    .ADR2(DLX_IDinst__n0456),
    .ADR3(DLX_IDinst_jtarget[15]),
    .O(DLX_IDinst_Madd__n0129_inst_lut2_227)
  );
  X_BUF \DLX_IDinst__n0129<28>/COUTUSED  (
    .I(\DLX_IDinst__n0129<28>/CYMUXG ),
    .O(DLX_IDinst_Madd__n0129_inst_cy_297)
  );
  X_BUF \DLX_IDinst__n0129<28>/XUSED  (
    .I(\DLX_IDinst__n0129<28>/XORF ),
    .O(DLX_IDinst__n0129[28])
  );
  X_BUF \DLX_IDinst__n0129<28>/YUSED  (
    .I(\DLX_IDinst__n0129<28>/XORG ),
    .O(DLX_IDinst__n0129[29])
  );
  X_MUX2 DLX_IDinst_Madd__n0129_inst_cy_297_473 (
    .IA(DLX_IFinst_NPC[29]),
    .IB(DLX_IDinst_Madd__n0129_inst_cy_296),
    .SEL(DLX_IDinst_Madd__n0129_inst_lut2_227),
    .O(\DLX_IDinst__n0129<28>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Madd__n0129_inst_sum_131 (
    .I0(DLX_IDinst_Madd__n0129_inst_cy_296),
    .I1(DLX_IDinst_Madd__n0129_inst_lut2_227),
    .O(\DLX_IDinst__n0129<28>/XORG )
  );
  X_BUF \DLX_IDinst__n0129<28>/CYINIT_474  (
    .I(DLX_IDinst_Madd__n0129_inst_cy_295),
    .O(\DLX_IDinst__n0129<28>/CYINIT )
  );
  X_MUX2 DLX_IDinst_Madd__n0129_inst_cy_298_475 (
    .IA(DLX_IFinst_NPC[30]),
    .IB(\DLX_IDinst__n0129<30>/CYINIT ),
    .SEL(DLX_IDinst_Madd__n0129_inst_lut2_228),
    .O(DLX_IDinst_Madd__n0129_inst_cy_298)
  );
  X_XOR2 DLX_IDinst_Madd__n0129_inst_sum_132 (
    .I0(\DLX_IDinst__n0129<30>/CYINIT ),
    .I1(DLX_IDinst_Madd__n0129_inst_lut2_228),
    .O(\DLX_IDinst__n0129<30>/XORF )
  );
  defparam DLX_IDinst_Madd__n0129_inst_lut2_2281.INIT = 16'h569A;
  X_LUT4 DLX_IDinst_Madd__n0129_inst_lut2_2281 (
    .ADR0(DLX_IFinst_NPC[30]),
    .ADR1(DLX_IDinst__n0456),
    .ADR2(DLX_IDinst_jtarget[15]),
    .ADR3(DLX_IDinst_regA_index[4]),
    .O(DLX_IDinst_Madd__n0129_inst_lut2_228)
  );
  defparam DLX_IDinst_Madd__n0129_inst_lut2_2291.INIT = 16'h569A;
  X_LUT4 DLX_IDinst_Madd__n0129_inst_lut2_2291 (
    .ADR0(DLX_IFinst_NPC[31]),
    .ADR1(DLX_IDinst__n0456),
    .ADR2(DLX_IDinst_jtarget[15]),
    .ADR3(DLX_IDinst_regA_index[4]),
    .O(DLX_IDinst_Madd__n0129_inst_lut2_229)
  );
  X_BUF \DLX_IDinst__n0129<30>/XUSED  (
    .I(\DLX_IDinst__n0129<30>/XORF ),
    .O(DLX_IDinst__n0129[30])
  );
  X_BUF \DLX_IDinst__n0129<30>/YUSED  (
    .I(\DLX_IDinst__n0129<30>/XORG ),
    .O(DLX_IDinst__n0129[31])
  );
  X_XOR2 DLX_IDinst_Madd__n0129_inst_sum_133 (
    .I0(DLX_IDinst_Madd__n0129_inst_cy_298),
    .I1(DLX_IDinst_Madd__n0129_inst_lut2_229),
    .O(\DLX_IDinst__n0129<30>/XORG )
  );
  X_BUF \DLX_IDinst__n0129<30>/CYINIT_476  (
    .I(DLX_IDinst_Madd__n0129_inst_cy_297),
    .O(\DLX_IDinst__n0129<30>/CYINIT )
  );
  X_ZERO \DLX_IDinst_Mcompar__n0003_inst_cy_266/LOGIC_ZERO_477  (
    .O(\DLX_IDinst_Mcompar__n0003_inst_cy_266/LOGIC_ZERO )
  );
  X_ONE \DLX_IDinst_Mcompar__n0003_inst_cy_266/LOGIC_ONE_478  (
    .O(\DLX_IDinst_Mcompar__n0003_inst_cy_266/LOGIC_ONE )
  );
  X_MUX2 DLX_IDinst_Mcompar__n0003_inst_cy_265_479 (
    .IA(\DLX_IDinst_Mcompar__n0003_inst_cy_266/LOGIC_ONE ),
    .IB(\DLX_IDinst_Mcompar__n0003_inst_cy_266/LOGIC_ZERO ),
    .SEL(DLX_IDinst_Mcompar__n0003_inst_lut4_43),
    .O(DLX_IDinst_Mcompar__n0003_inst_cy_265)
  );
  defparam DLX_IDinst_Mcompar__n0003_inst_lut4_431.INIT = 16'h9009;
  X_LUT4 DLX_IDinst_Mcompar__n0003_inst_lut4_431 (
    .ADR0(DLX_MEMinst_reg_dst_out[0]),
    .ADR1(DLX_IDinst_regB_index[0]),
    .ADR2(DLX_MEMinst_reg_dst_out[1]),
    .ADR3(DLX_IDinst_regB_index[1]),
    .O(DLX_IDinst_Mcompar__n0003_inst_lut4_43)
  );
  defparam DLX_IDinst_Mcompar__n0003_inst_lut4_441.INIT = 16'h8421;
  X_LUT4 DLX_IDinst_Mcompar__n0003_inst_lut4_441 (
    .ADR0(DLX_IDinst_regB_index[2]),
    .ADR1(DLX_MEMinst_reg_dst_out[3]),
    .ADR2(DLX_MEMinst_reg_dst_out[2]),
    .ADR3(DLX_IDinst_regB_index[3]),
    .O(DLX_IDinst_Mcompar__n0003_inst_lut4_44)
  );
  X_BUF \DLX_IDinst_Mcompar__n0003_inst_cy_266/COUTUSED  (
    .I(\DLX_IDinst_Mcompar__n0003_inst_cy_266/CYMUXG ),
    .O(DLX_IDinst_Mcompar__n0003_inst_cy_266)
  );
  X_MUX2 DLX_IDinst_Mcompar__n0003_inst_cy_266_480 (
    .IA(\DLX_IDinst_Mcompar__n0003_inst_cy_266/LOGIC_ONE ),
    .IB(DLX_IDinst_Mcompar__n0003_inst_cy_265),
    .SEL(DLX_IDinst_Mcompar__n0003_inst_lut4_44),
    .O(\DLX_IDinst_Mcompar__n0003_inst_cy_266/CYMUXG )
  );
  X_OR2 \DLX_IDinst_rt_addr<4>/FFY/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IDinst_rt_addr<4>/FFY/RST )
  );
  defparam DLX_IDinst_rt_addr_4.INIT = 1'b0;
  X_FF DLX_IDinst_rt_addr_4 (
    .I(DLX_IDinst__n0106[4]),
    .CE(DLX_IDinst__n0422),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_rt_addr<4>/FFY/RST ),
    .O(DLX_IDinst_rt_addr[4])
  );
  X_ONE \DLX_IDinst_rt_addr<4>/LOGIC_ONE_481  (
    .O(\DLX_IDinst_rt_addr<4>/LOGIC_ONE )
  );
  X_MUX2 DLX_IDinst_Mcompar__n0003_inst_cy_267 (
    .IA(\DLX_IDinst_rt_addr<4>/LOGIC_ONE ),
    .IB(\DLX_IDinst_rt_addr<4>/CYINIT ),
    .SEL(DLX_IDinst_Mcompar__n0003_inst_lut4_45),
    .O(\DLX_IDinst_rt_addr<4>/CYMUXF )
  );
  defparam DLX_IDinst_Mcompar__n0003_inst_lut4_451.INIT = 16'h9999;
  X_LUT4 DLX_IDinst_Mcompar__n0003_inst_lut4_451 (
    .ADR0(DLX_IDinst_regB_index[4]),
    .ADR1(DLX_MEMinst_reg_dst_out[4]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Mcompar__n0003_inst_lut4_45)
  );
  defparam \DLX_IDinst__n0106<4> .INIT = 16'hE000;
  X_LUT4 \DLX_IDinst__n0106<4>  (
    .ADR0(N90703),
    .ADR1(DLX_IDinst__n0364),
    .ADR2(DLX_IDinst_regB_index[4]),
    .ADR3(DLX_IDinst_N70679),
    .O(DLX_IDinst__n0106[4])
  );
  X_BUF \DLX_IDinst_rt_addr<4>/XBUSED  (
    .I(\DLX_IDinst_rt_addr<4>/CYMUXF ),
    .O(DLX_IDinst__n0003)
  );
  X_BUF \DLX_IDinst_rt_addr<4>/CYINIT_482  (
    .I(DLX_IDinst_Mcompar__n0003_inst_cy_266),
    .O(\DLX_IDinst_rt_addr<4>/CYINIT )
  );
  defparam vga_top_vga1_vcounter_0.INIT = 1'b0;
  X_SFF vga_top_vga1_vcounter_0 (
    .I(vga_top_vga1_vcounter_Madd__n0000_inst_lut2_9),
    .CE(N108996),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0007),
    .O(vga_top_vga1_vcounter[0])
  );
  defparam vga_top_vga1_vcounter_1.INIT = 1'b0;
  X_SFF vga_top_vga1_vcounter_1 (
    .I(vga_top_vga1_vcounter__n0000[1]),
    .CE(N108996),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0007),
    .O(vga_top_vga1_vcounter[1])
  );
  X_ZERO \vga_top_vga1_vcounter<0>/LOGIC_ZERO_483  (
    .O(\vga_top_vga1_vcounter<0>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_vcounter_Madd__n0000_inst_cy_9_484 (
    .IA(GLOBAL_LOGIC1_3),
    .IB(\vga_top_vga1_vcounter<0>/LOGIC_ZERO ),
    .SEL(vga_top_vga1_vcounter_Madd__n0000_inst_lut2_9),
    .O(vga_top_vga1_vcounter_Madd__n0000_inst_cy_9)
  );
  defparam vga_top_vga1_vcounter_Madd__n0000_inst_lut2_91.INIT = 16'h00FF;
  X_LUT4 vga_top_vga1_vcounter_Madd__n0000_inst_lut2_91 (
    .ADR0(GLOBAL_LOGIC1_3),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_vcounter[0]),
    .O(vga_top_vga1_vcounter_Madd__n0000_inst_lut2_9)
  );
  defparam \vga_top_vga1_vcounter<0>/G .INIT = 16'hF0F0;
  X_LUT4 \vga_top_vga1_vcounter<0>/G  (
    .ADR0(GLOBAL_LOGIC0_5),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_vcounter[1]),
    .ADR3(VCC),
    .O(\vga_top_vga1_vcounter<0>/GROM )
  );
  X_BUF \vga_top_vga1_vcounter<0>/COUTUSED  (
    .I(\vga_top_vga1_vcounter<0>/CYMUXG ),
    .O(vga_top_vga1_vcounter_Madd__n0000_inst_cy_10)
  );
  X_MUX2 vga_top_vga1_vcounter_Madd__n0000_inst_cy_10_485 (
    .IA(GLOBAL_LOGIC0_5),
    .IB(vga_top_vga1_vcounter_Madd__n0000_inst_cy_9),
    .SEL(\vga_top_vga1_vcounter<0>/GROM ),
    .O(\vga_top_vga1_vcounter<0>/CYMUXG )
  );
  X_XOR2 vga_top_vga1_vcounter_Madd__n0000_inst_sum_10 (
    .I0(vga_top_vga1_vcounter_Madd__n0000_inst_cy_9),
    .I1(\vga_top_vga1_vcounter<0>/GROM ),
    .O(vga_top_vga1_vcounter__n0000[1])
  );
  defparam vga_top_vga1_vcounter_3.INIT = 1'b0;
  X_SFF vga_top_vga1_vcounter_3 (
    .I(vga_top_vga1_vcounter__n0000[3]),
    .CE(N108996),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0007),
    .O(vga_top_vga1_vcounter[3])
  );
  defparam vga_top_vga1_vcounter_2.INIT = 1'b0;
  X_SFF vga_top_vga1_vcounter_2 (
    .I(vga_top_vga1_vcounter__n0000[2]),
    .CE(N108996),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0007),
    .O(vga_top_vga1_vcounter[2])
  );
  X_ZERO \vga_top_vga1_vcounter<2>/LOGIC_ZERO_486  (
    .O(\vga_top_vga1_vcounter<2>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_vcounter_Madd__n0000_inst_cy_11_487 (
    .IA(\vga_top_vga1_vcounter<2>/LOGIC_ZERO ),
    .IB(\vga_top_vga1_vcounter<2>/CYINIT ),
    .SEL(\vga_top_vga1_vcounter<2>/FROM ),
    .O(vga_top_vga1_vcounter_Madd__n0000_inst_cy_11)
  );
  X_XOR2 vga_top_vga1_vcounter_Madd__n0000_inst_sum_11 (
    .I0(\vga_top_vga1_vcounter<2>/CYINIT ),
    .I1(\vga_top_vga1_vcounter<2>/FROM ),
    .O(vga_top_vga1_vcounter__n0000[2])
  );
  defparam \vga_top_vga1_vcounter<2>/F .INIT = 16'hFF00;
  X_LUT4 \vga_top_vga1_vcounter<2>/F  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_vcounter[2]),
    .O(\vga_top_vga1_vcounter<2>/FROM )
  );
  defparam \vga_top_vga1_vcounter<2>/G .INIT = 16'hAAAA;
  X_LUT4 \vga_top_vga1_vcounter<2>/G  (
    .ADR0(vga_top_vga1_vcounter[3]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\vga_top_vga1_vcounter<2>/GROM )
  );
  X_BUF \vga_top_vga1_vcounter<2>/COUTUSED  (
    .I(\vga_top_vga1_vcounter<2>/CYMUXG ),
    .O(vga_top_vga1_vcounter_Madd__n0000_inst_cy_12)
  );
  X_MUX2 vga_top_vga1_vcounter_Madd__n0000_inst_cy_12_488 (
    .IA(\vga_top_vga1_vcounter<2>/LOGIC_ZERO ),
    .IB(vga_top_vga1_vcounter_Madd__n0000_inst_cy_11),
    .SEL(\vga_top_vga1_vcounter<2>/GROM ),
    .O(\vga_top_vga1_vcounter<2>/CYMUXG )
  );
  X_XOR2 vga_top_vga1_vcounter_Madd__n0000_inst_sum_12 (
    .I0(vga_top_vga1_vcounter_Madd__n0000_inst_cy_11),
    .I1(\vga_top_vga1_vcounter<2>/GROM ),
    .O(vga_top_vga1_vcounter__n0000[3])
  );
  X_BUF \vga_top_vga1_vcounter<2>/CYINIT_489  (
    .I(vga_top_vga1_vcounter_Madd__n0000_inst_cy_10),
    .O(\vga_top_vga1_vcounter<2>/CYINIT )
  );
  defparam vga_top_vga1_vcounter_5.INIT = 1'b0;
  X_SFF vga_top_vga1_vcounter_5 (
    .I(vga_top_vga1_vcounter__n0000[5]),
    .CE(N108996),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0007),
    .O(vga_top_vga1_vcounter[5])
  );
  X_ZERO \vga_top_vga1_vcounter<4>/LOGIC_ZERO_490  (
    .O(\vga_top_vga1_vcounter<4>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_vcounter_Madd__n0000_inst_cy_13_491 (
    .IA(\vga_top_vga1_vcounter<4>/LOGIC_ZERO ),
    .IB(\vga_top_vga1_vcounter<4>/CYINIT ),
    .SEL(\vga_top_vga1_vcounter<4>/FROM ),
    .O(vga_top_vga1_vcounter_Madd__n0000_inst_cy_13)
  );
  X_XOR2 vga_top_vga1_vcounter_Madd__n0000_inst_sum_13 (
    .I0(\vga_top_vga1_vcounter<4>/CYINIT ),
    .I1(\vga_top_vga1_vcounter<4>/FROM ),
    .O(vga_top_vga1_vcounter__n0000[4])
  );
  defparam \vga_top_vga1_vcounter<4>/F .INIT = 16'hFF00;
  X_LUT4 \vga_top_vga1_vcounter<4>/F  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_vcounter[4]),
    .O(\vga_top_vga1_vcounter<4>/FROM )
  );
  defparam \vga_top_vga1_vcounter<4>/G .INIT = 16'hCCCC;
  X_LUT4 \vga_top_vga1_vcounter<4>/G  (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_vcounter[5]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\vga_top_vga1_vcounter<4>/GROM )
  );
  X_BUF \vga_top_vga1_vcounter<4>/COUTUSED  (
    .I(\vga_top_vga1_vcounter<4>/CYMUXG ),
    .O(vga_top_vga1_vcounter_Madd__n0000_inst_cy_14)
  );
  X_MUX2 vga_top_vga1_vcounter_Madd__n0000_inst_cy_14_492 (
    .IA(\vga_top_vga1_vcounter<4>/LOGIC_ZERO ),
    .IB(vga_top_vga1_vcounter_Madd__n0000_inst_cy_13),
    .SEL(\vga_top_vga1_vcounter<4>/GROM ),
    .O(\vga_top_vga1_vcounter<4>/CYMUXG )
  );
  X_XOR2 vga_top_vga1_vcounter_Madd__n0000_inst_sum_14 (
    .I0(vga_top_vga1_vcounter_Madd__n0000_inst_cy_13),
    .I1(\vga_top_vga1_vcounter<4>/GROM ),
    .O(vga_top_vga1_vcounter__n0000[5])
  );
  X_BUF \vga_top_vga1_vcounter<4>/CYINIT_493  (
    .I(vga_top_vga1_vcounter_Madd__n0000_inst_cy_12),
    .O(\vga_top_vga1_vcounter<4>/CYINIT )
  );
  defparam vga_top_vga1_vcounter_7.INIT = 1'b0;
  X_SFF vga_top_vga1_vcounter_7 (
    .I(vga_top_vga1_vcounter__n0000[7]),
    .CE(N108996),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0007),
    .O(vga_top_vga1_vcounter[7])
  );
  X_ZERO \vga_top_vga1_vcounter<6>/LOGIC_ZERO_494  (
    .O(\vga_top_vga1_vcounter<6>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_vcounter_Madd__n0000_inst_cy_15_495 (
    .IA(\vga_top_vga1_vcounter<6>/LOGIC_ZERO ),
    .IB(\vga_top_vga1_vcounter<6>/CYINIT ),
    .SEL(\vga_top_vga1_vcounter<6>/FROM ),
    .O(vga_top_vga1_vcounter_Madd__n0000_inst_cy_15)
  );
  X_XOR2 vga_top_vga1_vcounter_Madd__n0000_inst_sum_15 (
    .I0(\vga_top_vga1_vcounter<6>/CYINIT ),
    .I1(\vga_top_vga1_vcounter<6>/FROM ),
    .O(vga_top_vga1_vcounter__n0000[6])
  );
  defparam \vga_top_vga1_vcounter<6>/F .INIT = 16'hFF00;
  X_LUT4 \vga_top_vga1_vcounter<6>/F  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_vcounter[6]),
    .O(\vga_top_vga1_vcounter<6>/FROM )
  );
  defparam \vga_top_vga1_vcounter<6>/G .INIT = 16'hF0F0;
  X_LUT4 \vga_top_vga1_vcounter<6>/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_vcounter[7]),
    .ADR3(VCC),
    .O(\vga_top_vga1_vcounter<6>/GROM )
  );
  X_BUF \vga_top_vga1_vcounter<6>/COUTUSED  (
    .I(\vga_top_vga1_vcounter<6>/CYMUXG ),
    .O(vga_top_vga1_vcounter_Madd__n0000_inst_cy_16)
  );
  X_MUX2 vga_top_vga1_vcounter_Madd__n0000_inst_cy_16_496 (
    .IA(\vga_top_vga1_vcounter<6>/LOGIC_ZERO ),
    .IB(vga_top_vga1_vcounter_Madd__n0000_inst_cy_15),
    .SEL(\vga_top_vga1_vcounter<6>/GROM ),
    .O(\vga_top_vga1_vcounter<6>/CYMUXG )
  );
  X_XOR2 vga_top_vga1_vcounter_Madd__n0000_inst_sum_16 (
    .I0(vga_top_vga1_vcounter_Madd__n0000_inst_cy_15),
    .I1(\vga_top_vga1_vcounter<6>/GROM ),
    .O(vga_top_vga1_vcounter__n0000[7])
  );
  X_BUF \vga_top_vga1_vcounter<6>/CYINIT_497  (
    .I(vga_top_vga1_vcounter_Madd__n0000_inst_cy_14),
    .O(\vga_top_vga1_vcounter<6>/CYINIT )
  );
  X_ZERO \vga_top_vga1_vcounter<8>/LOGIC_ZERO_498  (
    .O(\vga_top_vga1_vcounter<8>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_vcounter_Madd__n0000_inst_cy_17_499 (
    .IA(\vga_top_vga1_vcounter<8>/LOGIC_ZERO ),
    .IB(\vga_top_vga1_vcounter<8>/CYINIT ),
    .SEL(\vga_top_vga1_vcounter<8>/FROM ),
    .O(vga_top_vga1_vcounter_Madd__n0000_inst_cy_17)
  );
  X_XOR2 vga_top_vga1_vcounter_Madd__n0000_inst_sum_17 (
    .I0(\vga_top_vga1_vcounter<8>/CYINIT ),
    .I1(\vga_top_vga1_vcounter<8>/FROM ),
    .O(vga_top_vga1_vcounter__n0000[8])
  );
  defparam \vga_top_vga1_vcounter<8>/F .INIT = 16'hFF00;
  X_LUT4 \vga_top_vga1_vcounter<8>/F  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_vcounter[8]),
    .O(\vga_top_vga1_vcounter<8>/FROM )
  );
  defparam \vga_top_vga1_vcounter<9>_rt_500 .INIT = 16'hFF00;
  X_LUT4 \vga_top_vga1_vcounter<9>_rt_500  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_vcounter[9]),
    .O(\vga_top_vga1_vcounter<9>_rt )
  );
  X_XOR2 vga_top_vga1_vcounter_Madd__n0000_inst_sum_18 (
    .I0(vga_top_vga1_vcounter_Madd__n0000_inst_cy_17),
    .I1(\vga_top_vga1_vcounter<9>_rt ),
    .O(vga_top_vga1_vcounter__n0000[9])
  );
  X_BUF \vga_top_vga1_vcounter<8>/CYINIT_501  (
    .I(vga_top_vga1_vcounter_Madd__n0000_inst_cy_16),
    .O(\vga_top_vga1_vcounter<8>/CYINIT )
  );
  X_ZERO \vga_top_vga1_hcounter<0>/LOGIC_ZERO_502  (
    .O(\vga_top_vga1_hcounter<0>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_hcounter_Madd__n0000_inst_cy_19_503 (
    .IA(GLOBAL_LOGIC1_2),
    .IB(\vga_top_vga1_hcounter<0>/LOGIC_ZERO ),
    .SEL(vga_top_vga1_hcounter_Madd__n0000_inst_lut2_19),
    .O(vga_top_vga1_hcounter_Madd__n0000_inst_cy_19)
  );
  defparam vga_top_vga1_hcounter_Madd__n0000_inst_lut2_191.INIT = 16'h0F0F;
  X_LUT4 vga_top_vga1_hcounter_Madd__n0000_inst_lut2_191 (
    .ADR0(GLOBAL_LOGIC1_2),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_hcounter[0]),
    .ADR3(VCC),
    .O(vga_top_vga1_hcounter_Madd__n0000_inst_lut2_19)
  );
  defparam \vga_top_vga1_hcounter<0>/G .INIT = 16'hFF00;
  X_LUT4 \vga_top_vga1_hcounter<0>/G  (
    .ADR0(GLOBAL_LOGIC0_6),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[1]),
    .O(\vga_top_vga1_hcounter<0>/GROM )
  );
  X_BUF \vga_top_vga1_hcounter<0>/COUTUSED  (
    .I(\vga_top_vga1_hcounter<0>/CYMUXG ),
    .O(vga_top_vga1_hcounter_Madd__n0000_inst_cy_20)
  );
  X_MUX2 vga_top_vga1_hcounter_Madd__n0000_inst_cy_20_504 (
    .IA(GLOBAL_LOGIC0_6),
    .IB(vga_top_vga1_hcounter_Madd__n0000_inst_cy_19),
    .SEL(\vga_top_vga1_hcounter<0>/GROM ),
    .O(\vga_top_vga1_hcounter<0>/CYMUXG )
  );
  X_XOR2 vga_top_vga1_hcounter_Madd__n0000_inst_sum_20 (
    .I0(vga_top_vga1_hcounter_Madd__n0000_inst_cy_19),
    .I1(\vga_top_vga1_hcounter<0>/GROM ),
    .O(vga_top_vga1_hcounter__n0000[1])
  );
  X_ZERO \vga_top_vga1_hcounter<2>/LOGIC_ZERO_505  (
    .O(\vga_top_vga1_hcounter<2>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_hcounter_Madd__n0000_inst_cy_21_506 (
    .IA(\vga_top_vga1_hcounter<2>/LOGIC_ZERO ),
    .IB(\vga_top_vga1_hcounter<2>/CYINIT ),
    .SEL(\vga_top_vga1_hcounter<2>/FROM ),
    .O(vga_top_vga1_hcounter_Madd__n0000_inst_cy_21)
  );
  X_XOR2 vga_top_vga1_hcounter_Madd__n0000_inst_sum_21 (
    .I0(\vga_top_vga1_hcounter<2>/CYINIT ),
    .I1(\vga_top_vga1_hcounter<2>/FROM ),
    .O(vga_top_vga1_hcounter__n0000[2])
  );
  defparam \vga_top_vga1_hcounter<2>/F .INIT = 16'hFF00;
  X_LUT4 \vga_top_vga1_hcounter<2>/F  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[2]),
    .O(\vga_top_vga1_hcounter<2>/FROM )
  );
  defparam \vga_top_vga1_hcounter<2>/G .INIT = 16'hCCCC;
  X_LUT4 \vga_top_vga1_hcounter<2>/G  (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_hcounter[3]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\vga_top_vga1_hcounter<2>/GROM )
  );
  X_BUF \vga_top_vga1_hcounter<2>/COUTUSED  (
    .I(\vga_top_vga1_hcounter<2>/CYMUXG ),
    .O(vga_top_vga1_hcounter_Madd__n0000_inst_cy_22)
  );
  X_MUX2 vga_top_vga1_hcounter_Madd__n0000_inst_cy_22_507 (
    .IA(\vga_top_vga1_hcounter<2>/LOGIC_ZERO ),
    .IB(vga_top_vga1_hcounter_Madd__n0000_inst_cy_21),
    .SEL(\vga_top_vga1_hcounter<2>/GROM ),
    .O(\vga_top_vga1_hcounter<2>/CYMUXG )
  );
  X_XOR2 vga_top_vga1_hcounter_Madd__n0000_inst_sum_22 (
    .I0(vga_top_vga1_hcounter_Madd__n0000_inst_cy_21),
    .I1(\vga_top_vga1_hcounter<2>/GROM ),
    .O(vga_top_vga1_hcounter__n0000[3])
  );
  X_BUF \vga_top_vga1_hcounter<2>/CYINIT_508  (
    .I(vga_top_vga1_hcounter_Madd__n0000_inst_cy_20),
    .O(\vga_top_vga1_hcounter<2>/CYINIT )
  );
  X_ZERO \vga_top_vga1_hcounter<4>/LOGIC_ZERO_509  (
    .O(\vga_top_vga1_hcounter<4>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_hcounter_Madd__n0000_inst_cy_23_510 (
    .IA(\vga_top_vga1_hcounter<4>/LOGIC_ZERO ),
    .IB(\vga_top_vga1_hcounter<4>/CYINIT ),
    .SEL(\vga_top_vga1_hcounter<4>/FROM ),
    .O(vga_top_vga1_hcounter_Madd__n0000_inst_cy_23)
  );
  X_XOR2 vga_top_vga1_hcounter_Madd__n0000_inst_sum_23 (
    .I0(\vga_top_vga1_hcounter<4>/CYINIT ),
    .I1(\vga_top_vga1_hcounter<4>/FROM ),
    .O(vga_top_vga1_hcounter__n0000[4])
  );
  defparam \vga_top_vga1_hcounter<4>/F .INIT = 16'hFF00;
  X_LUT4 \vga_top_vga1_hcounter<4>/F  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[4]),
    .O(\vga_top_vga1_hcounter<4>/FROM )
  );
  defparam \vga_top_vga1_hcounter<4>/G .INIT = 16'hF0F0;
  X_LUT4 \vga_top_vga1_hcounter<4>/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_hcounter[5]),
    .ADR3(VCC),
    .O(\vga_top_vga1_hcounter<4>/GROM )
  );
  X_BUF \vga_top_vga1_hcounter<4>/COUTUSED  (
    .I(\vga_top_vga1_hcounter<4>/CYMUXG ),
    .O(vga_top_vga1_hcounter_Madd__n0000_inst_cy_24)
  );
  X_MUX2 vga_top_vga1_hcounter_Madd__n0000_inst_cy_24_511 (
    .IA(\vga_top_vga1_hcounter<4>/LOGIC_ZERO ),
    .IB(vga_top_vga1_hcounter_Madd__n0000_inst_cy_23),
    .SEL(\vga_top_vga1_hcounter<4>/GROM ),
    .O(\vga_top_vga1_hcounter<4>/CYMUXG )
  );
  X_XOR2 vga_top_vga1_hcounter_Madd__n0000_inst_sum_24 (
    .I0(vga_top_vga1_hcounter_Madd__n0000_inst_cy_23),
    .I1(\vga_top_vga1_hcounter<4>/GROM ),
    .O(vga_top_vga1_hcounter__n0000[5])
  );
  X_BUF \vga_top_vga1_hcounter<4>/CYINIT_512  (
    .I(vga_top_vga1_hcounter_Madd__n0000_inst_cy_22),
    .O(\vga_top_vga1_hcounter<4>/CYINIT )
  );
  X_ZERO \vga_top_vga1_hcounter<6>/LOGIC_ZERO_513  (
    .O(\vga_top_vga1_hcounter<6>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_hcounter_Madd__n0000_inst_cy_25_514 (
    .IA(\vga_top_vga1_hcounter<6>/LOGIC_ZERO ),
    .IB(\vga_top_vga1_hcounter<6>/CYINIT ),
    .SEL(\vga_top_vga1_hcounter<6>/FROM ),
    .O(vga_top_vga1_hcounter_Madd__n0000_inst_cy_25)
  );
  X_XOR2 vga_top_vga1_hcounter_Madd__n0000_inst_sum_25 (
    .I0(\vga_top_vga1_hcounter<6>/CYINIT ),
    .I1(\vga_top_vga1_hcounter<6>/FROM ),
    .O(vga_top_vga1_hcounter__n0000[6])
  );
  defparam \vga_top_vga1_hcounter<6>/F .INIT = 16'hFF00;
  X_LUT4 \vga_top_vga1_hcounter<6>/F  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[6]),
    .O(\vga_top_vga1_hcounter<6>/FROM )
  );
  defparam \vga_top_vga1_hcounter<6>/G .INIT = 16'hFF00;
  X_LUT4 \vga_top_vga1_hcounter<6>/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[7]),
    .O(\vga_top_vga1_hcounter<6>/GROM )
  );
  X_BUF \vga_top_vga1_hcounter<6>/COUTUSED  (
    .I(\vga_top_vga1_hcounter<6>/CYMUXG ),
    .O(vga_top_vga1_hcounter_Madd__n0000_inst_cy_26)
  );
  X_MUX2 vga_top_vga1_hcounter_Madd__n0000_inst_cy_26_515 (
    .IA(\vga_top_vga1_hcounter<6>/LOGIC_ZERO ),
    .IB(vga_top_vga1_hcounter_Madd__n0000_inst_cy_25),
    .SEL(\vga_top_vga1_hcounter<6>/GROM ),
    .O(\vga_top_vga1_hcounter<6>/CYMUXG )
  );
  X_XOR2 vga_top_vga1_hcounter_Madd__n0000_inst_sum_26 (
    .I0(vga_top_vga1_hcounter_Madd__n0000_inst_cy_25),
    .I1(\vga_top_vga1_hcounter<6>/GROM ),
    .O(vga_top_vga1_hcounter__n0000[7])
  );
  X_BUF \vga_top_vga1_hcounter<6>/CYINIT_516  (
    .I(vga_top_vga1_hcounter_Madd__n0000_inst_cy_24),
    .O(\vga_top_vga1_hcounter<6>/CYINIT )
  );
  X_ZERO \vga_top_vga1_hcounter<8>/LOGIC_ZERO_517  (
    .O(\vga_top_vga1_hcounter<8>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_hcounter_Madd__n0000_inst_cy_27_518 (
    .IA(\vga_top_vga1_hcounter<8>/LOGIC_ZERO ),
    .IB(\vga_top_vga1_hcounter<8>/CYINIT ),
    .SEL(\vga_top_vga1_hcounter<8>/FROM ),
    .O(vga_top_vga1_hcounter_Madd__n0000_inst_cy_27)
  );
  X_XOR2 vga_top_vga1_hcounter_Madd__n0000_inst_sum_27 (
    .I0(\vga_top_vga1_hcounter<8>/CYINIT ),
    .I1(\vga_top_vga1_hcounter<8>/FROM ),
    .O(vga_top_vga1_hcounter__n0000[8])
  );
  defparam \vga_top_vga1_hcounter<8>/F .INIT = 16'hFF00;
  X_LUT4 \vga_top_vga1_hcounter<8>/F  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[8]),
    .O(\vga_top_vga1_hcounter<8>/FROM )
  );
  defparam \vga_top_vga1_hcounter<8>/G .INIT = 16'hFF00;
  X_LUT4 \vga_top_vga1_hcounter<8>/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[9]),
    .O(\vga_top_vga1_hcounter<8>/GROM )
  );
  X_BUF \vga_top_vga1_hcounter<8>/COUTUSED  (
    .I(\vga_top_vga1_hcounter<8>/CYMUXG ),
    .O(vga_top_vga1_hcounter_Madd__n0000_inst_cy_28)
  );
  X_MUX2 vga_top_vga1_hcounter_Madd__n0000_inst_cy_28_519 (
    .IA(\vga_top_vga1_hcounter<8>/LOGIC_ZERO ),
    .IB(vga_top_vga1_hcounter_Madd__n0000_inst_cy_27),
    .SEL(\vga_top_vga1_hcounter<8>/GROM ),
    .O(\vga_top_vga1_hcounter<8>/CYMUXG )
  );
  X_XOR2 vga_top_vga1_hcounter_Madd__n0000_inst_sum_28 (
    .I0(vga_top_vga1_hcounter_Madd__n0000_inst_cy_27),
    .I1(\vga_top_vga1_hcounter<8>/GROM ),
    .O(vga_top_vga1_hcounter__n0000[9])
  );
  X_BUF \vga_top_vga1_hcounter<8>/CYINIT_520  (
    .I(vga_top_vga1_hcounter_Madd__n0000_inst_cy_26),
    .O(\vga_top_vga1_hcounter<8>/CYINIT )
  );
  X_ZERO \vga_top_vga1_hcounter<10>/LOGIC_ZERO_521  (
    .O(\vga_top_vga1_hcounter<10>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_hcounter_Madd__n0000_inst_cy_29_522 (
    .IA(\vga_top_vga1_hcounter<10>/LOGIC_ZERO ),
    .IB(\vga_top_vga1_hcounter<10>/CYINIT ),
    .SEL(\vga_top_vga1_hcounter<10>/FROM ),
    .O(vga_top_vga1_hcounter_Madd__n0000_inst_cy_29)
  );
  X_XOR2 vga_top_vga1_hcounter_Madd__n0000_inst_sum_29 (
    .I0(\vga_top_vga1_hcounter<10>/CYINIT ),
    .I1(\vga_top_vga1_hcounter<10>/FROM ),
    .O(vga_top_vga1_hcounter__n0000[10])
  );
  defparam \vga_top_vga1_hcounter<10>/F .INIT = 16'hFF00;
  X_LUT4 \vga_top_vga1_hcounter<10>/F  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[10]),
    .O(\vga_top_vga1_hcounter<10>/FROM )
  );
  defparam \vga_top_vga1_hcounter<10>/G .INIT = 16'hFF00;
  X_LUT4 \vga_top_vga1_hcounter<10>/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[11]),
    .O(\vga_top_vga1_hcounter<10>/GROM )
  );
  X_BUF \vga_top_vga1_hcounter<10>/COUTUSED  (
    .I(\vga_top_vga1_hcounter<10>/CYMUXG ),
    .O(vga_top_vga1_hcounter_Madd__n0000_inst_cy_30)
  );
  X_MUX2 vga_top_vga1_hcounter_Madd__n0000_inst_cy_30_523 (
    .IA(\vga_top_vga1_hcounter<10>/LOGIC_ZERO ),
    .IB(vga_top_vga1_hcounter_Madd__n0000_inst_cy_29),
    .SEL(\vga_top_vga1_hcounter<10>/GROM ),
    .O(\vga_top_vga1_hcounter<10>/CYMUXG )
  );
  X_XOR2 vga_top_vga1_hcounter_Madd__n0000_inst_sum_30 (
    .I0(vga_top_vga1_hcounter_Madd__n0000_inst_cy_29),
    .I1(\vga_top_vga1_hcounter<10>/GROM ),
    .O(vga_top_vga1_hcounter__n0000[11])
  );
  X_BUF \vga_top_vga1_hcounter<10>/CYINIT_524  (
    .I(vga_top_vga1_hcounter_Madd__n0000_inst_cy_28),
    .O(\vga_top_vga1_hcounter<10>/CYINIT )
  );
  X_ZERO \vga_top_vga1_hcounter<12>/LOGIC_ZERO_525  (
    .O(\vga_top_vga1_hcounter<12>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_hcounter_Madd__n0000_inst_cy_31_526 (
    .IA(\vga_top_vga1_hcounter<12>/LOGIC_ZERO ),
    .IB(\vga_top_vga1_hcounter<12>/CYINIT ),
    .SEL(\vga_top_vga1_hcounter<12>/FROM ),
    .O(vga_top_vga1_hcounter_Madd__n0000_inst_cy_31)
  );
  X_XOR2 vga_top_vga1_hcounter_Madd__n0000_inst_sum_31 (
    .I0(\vga_top_vga1_hcounter<12>/CYINIT ),
    .I1(\vga_top_vga1_hcounter<12>/FROM ),
    .O(vga_top_vga1_hcounter__n0000[12])
  );
  defparam \vga_top_vga1_hcounter<12>/F .INIT = 16'hFF00;
  X_LUT4 \vga_top_vga1_hcounter<12>/F  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[12]),
    .O(\vga_top_vga1_hcounter<12>/FROM )
  );
  defparam \vga_top_vga1_hcounter<12>/G .INIT = 16'hFF00;
  X_LUT4 \vga_top_vga1_hcounter<12>/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[13]),
    .O(\vga_top_vga1_hcounter<12>/GROM )
  );
  X_BUF \vga_top_vga1_hcounter<12>/COUTUSED  (
    .I(\vga_top_vga1_hcounter<12>/CYMUXG ),
    .O(vga_top_vga1_hcounter_Madd__n0000_inst_cy_32)
  );
  X_MUX2 vga_top_vga1_hcounter_Madd__n0000_inst_cy_32_527 (
    .IA(\vga_top_vga1_hcounter<12>/LOGIC_ZERO ),
    .IB(vga_top_vga1_hcounter_Madd__n0000_inst_cy_31),
    .SEL(\vga_top_vga1_hcounter<12>/GROM ),
    .O(\vga_top_vga1_hcounter<12>/CYMUXG )
  );
  X_XOR2 vga_top_vga1_hcounter_Madd__n0000_inst_sum_32 (
    .I0(vga_top_vga1_hcounter_Madd__n0000_inst_cy_31),
    .I1(\vga_top_vga1_hcounter<12>/GROM ),
    .O(vga_top_vga1_hcounter__n0000[13])
  );
  X_BUF \vga_top_vga1_hcounter<12>/CYINIT_528  (
    .I(vga_top_vga1_hcounter_Madd__n0000_inst_cy_30),
    .O(\vga_top_vga1_hcounter<12>/CYINIT )
  );
  X_ZERO \vga_top_vga1_hcounter<14>/LOGIC_ZERO_529  (
    .O(\vga_top_vga1_hcounter<14>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_hcounter_Madd__n0000_inst_cy_33_530 (
    .IA(\vga_top_vga1_hcounter<14>/LOGIC_ZERO ),
    .IB(\vga_top_vga1_hcounter<14>/CYINIT ),
    .SEL(\vga_top_vga1_hcounter<14>/FROM ),
    .O(vga_top_vga1_hcounter_Madd__n0000_inst_cy_33)
  );
  X_XOR2 vga_top_vga1_hcounter_Madd__n0000_inst_sum_33 (
    .I0(\vga_top_vga1_hcounter<14>/CYINIT ),
    .I1(\vga_top_vga1_hcounter<14>/FROM ),
    .O(vga_top_vga1_hcounter__n0000[14])
  );
  defparam \vga_top_vga1_hcounter<14>/F .INIT = 16'hFF00;
  X_LUT4 \vga_top_vga1_hcounter<14>/F  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[14]),
    .O(\vga_top_vga1_hcounter<14>/FROM )
  );
  defparam \vga_top_vga1_hcounter<15>_rt_531 .INIT = 16'hFF00;
  X_LUT4 \vga_top_vga1_hcounter<15>_rt_531  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[15]),
    .O(\vga_top_vga1_hcounter<15>_rt )
  );
  X_XOR2 vga_top_vga1_hcounter_Madd__n0000_inst_sum_34 (
    .I0(vga_top_vga1_hcounter_Madd__n0000_inst_cy_33),
    .I1(\vga_top_vga1_hcounter<15>_rt ),
    .O(vga_top_vga1_hcounter__n0000[15])
  );
  X_BUF \vga_top_vga1_hcounter<14>/CYINIT_532  (
    .I(vga_top_vga1_hcounter_Madd__n0000_inst_cy_32),
    .O(\vga_top_vga1_hcounter<14>/CYINIT )
  );
  X_ONE \DLX_EXinst_Mcompar__n0085_inst_cy_103/LOGIC_ONE_533  (
    .O(\DLX_EXinst_Mcompar__n0085_inst_cy_103/LOGIC_ONE )
  );
  X_ZERO \DLX_EXinst_Mcompar__n0085_inst_cy_103/LOGIC_ZERO_534  (
    .O(\DLX_EXinst_Mcompar__n0085_inst_cy_103/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0085_inst_cy_102_535 (
    .IA(\DLX_EXinst_Mcompar__n0085_inst_cy_103/LOGIC_ZERO ),
    .IB(\DLX_EXinst_Mcompar__n0085_inst_cy_103/LOGIC_ONE ),
    .SEL(DLX_EXinst_Mcompar__n0085_inst_lut4_0),
    .O(DLX_EXinst_Mcompar__n0085_inst_cy_102)
  );
  defparam DLX_EXinst_Mcompar__n0085_inst_lut4_01.INIT = 16'h8241;
  X_LUT4 DLX_EXinst_Mcompar__n0085_inst_lut4_01 (
    .ADR0(DLX_IDinst_IR_function_field_0_1),
    .ADR1(DLX_IDinst_IR_function_field_1_1),
    .ADR2(DLX_IDinst_reg_out_A[1]),
    .ADR3(DLX_IDinst_reg_out_A[0]),
    .O(DLX_EXinst_Mcompar__n0085_inst_lut4_0)
  );
  defparam DLX_EXinst_Mcompar__n0085_inst_lut4_16.INIT = 16'h8241;
  X_LUT4 DLX_EXinst_Mcompar__n0085_inst_lut4_16 (
    .ADR0(DLX_IDinst_reg_out_A[3]),
    .ADR1(DLX_IDinst_reg_out_A[2]),
    .ADR2(DLX_IDinst_IR_function_field_2_1),
    .ADR3(DLX_IDinst_IR_function_field_3_1),
    .O(DLX_EXinst_Mcompar__n0085_inst_lut4_1)
  );
  X_BUF \DLX_EXinst_Mcompar__n0085_inst_cy_103/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0085_inst_cy_103/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0085_inst_cy_103)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0085_inst_cy_103_536 (
    .IA(\DLX_EXinst_Mcompar__n0085_inst_cy_103/LOGIC_ZERO ),
    .IB(DLX_EXinst_Mcompar__n0085_inst_cy_102),
    .SEL(DLX_EXinst_Mcompar__n0085_inst_lut4_1),
    .O(\DLX_EXinst_Mcompar__n0085_inst_cy_103/CYMUXG )
  );
  X_ZERO \DLX_EXinst_Mcompar__n0085_inst_cy_105/LOGIC_ZERO_537  (
    .O(\DLX_EXinst_Mcompar__n0085_inst_cy_105/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0085_inst_cy_104_538 (
    .IA(\DLX_EXinst_Mcompar__n0085_inst_cy_105/LOGIC_ZERO ),
    .IB(\DLX_EXinst_Mcompar__n0085_inst_cy_105/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0085_inst_lut4_2),
    .O(DLX_EXinst_Mcompar__n0085_inst_cy_104)
  );
  defparam DLX_EXinst_Mcompar__n0085_inst_lut4_21.INIT = 16'h8241;
  X_LUT4 DLX_EXinst_Mcompar__n0085_inst_lut4_21 (
    .ADR0(DLX_IDinst_IR_function_field[4]),
    .ADR1(\DLX_IDinst_Imm[5] ),
    .ADR2(DLX_IDinst_reg_out_A[5]),
    .ADR3(DLX_IDinst_reg_out_A[4]),
    .O(DLX_EXinst_Mcompar__n0085_inst_lut4_2)
  );
  defparam DLX_EXinst_Mcompar__n0085_inst_lut4_31.INIT = 16'h8241;
  X_LUT4 DLX_EXinst_Mcompar__n0085_inst_lut4_31 (
    .ADR0(\DLX_IDinst_Imm[7] ),
    .ADR1(\DLX_IDinst_Imm[6] ),
    .ADR2(DLX_IDinst_reg_out_A[6]),
    .ADR3(DLX_IDinst_reg_out_A[7]),
    .O(DLX_EXinst_Mcompar__n0085_inst_lut4_3)
  );
  X_BUF \DLX_EXinst_Mcompar__n0085_inst_cy_105/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0085_inst_cy_105/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0085_inst_cy_105)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0085_inst_cy_105_539 (
    .IA(\DLX_EXinst_Mcompar__n0085_inst_cy_105/LOGIC_ZERO ),
    .IB(DLX_EXinst_Mcompar__n0085_inst_cy_104),
    .SEL(DLX_EXinst_Mcompar__n0085_inst_lut4_3),
    .O(\DLX_EXinst_Mcompar__n0085_inst_cy_105/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0085_inst_cy_105/CYINIT_540  (
    .I(DLX_EXinst_Mcompar__n0085_inst_cy_103),
    .O(\DLX_EXinst_Mcompar__n0085_inst_cy_105/CYINIT )
  );
  X_ZERO \DLX_EXinst_Mcompar__n0085_inst_cy_107/LOGIC_ZERO_541  (
    .O(\DLX_EXinst_Mcompar__n0085_inst_cy_107/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0085_inst_cy_106_542 (
    .IA(\DLX_EXinst_Mcompar__n0085_inst_cy_107/LOGIC_ZERO ),
    .IB(\DLX_EXinst_Mcompar__n0085_inst_cy_107/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0085_inst_lut4_4),
    .O(DLX_EXinst_Mcompar__n0085_inst_cy_106)
  );
  defparam DLX_EXinst_Mcompar__n0085_inst_lut4_41.INIT = 16'h8241;
  X_LUT4 DLX_EXinst_Mcompar__n0085_inst_lut4_41 (
    .ADR0(\DLX_IDinst_Imm[9] ),
    .ADR1(DLX_IDinst_reg_out_A[8]),
    .ADR2(\DLX_IDinst_Imm[8] ),
    .ADR3(DLX_IDinst_reg_out_A[9]),
    .O(DLX_EXinst_Mcompar__n0085_inst_lut4_4)
  );
  defparam DLX_EXinst_Mcompar__n0085_inst_lut4_51.INIT = 16'h8241;
  X_LUT4 DLX_EXinst_Mcompar__n0085_inst_lut4_51 (
    .ADR0(DLX_IDinst_reg_out_A[10]),
    .ADR1(DLX_IDinst_reg_out_A[11]),
    .ADR2(\DLX_IDinst_Imm[11] ),
    .ADR3(\DLX_IDinst_Imm[10] ),
    .O(DLX_EXinst_Mcompar__n0085_inst_lut4_5)
  );
  X_BUF \DLX_EXinst_Mcompar__n0085_inst_cy_107/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0085_inst_cy_107/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0085_inst_cy_107)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0085_inst_cy_107_543 (
    .IA(\DLX_EXinst_Mcompar__n0085_inst_cy_107/LOGIC_ZERO ),
    .IB(DLX_EXinst_Mcompar__n0085_inst_cy_106),
    .SEL(DLX_EXinst_Mcompar__n0085_inst_lut4_5),
    .O(\DLX_EXinst_Mcompar__n0085_inst_cy_107/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0085_inst_cy_107/CYINIT_544  (
    .I(DLX_EXinst_Mcompar__n0085_inst_cy_105),
    .O(\DLX_EXinst_Mcompar__n0085_inst_cy_107/CYINIT )
  );
  defparam DLX_IFinst_NPC_6_1_545.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_6_1_545 (
    .I(\NPC_eff<6>/OD ),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\NPC_eff<6>/OFF/RST ),
    .O(DLX_IFinst_NPC_6_1)
  );
  X_OR2 \NPC_eff<6>/OFF/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\NPC_eff<6>/OFF/RST )
  );
  X_ZERO \DLX_EXinst_Mcompar__n0085_inst_cy_109/LOGIC_ZERO_546  (
    .O(\DLX_EXinst_Mcompar__n0085_inst_cy_109/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0085_inst_cy_108_547 (
    .IA(\DLX_EXinst_Mcompar__n0085_inst_cy_109/LOGIC_ZERO ),
    .IB(\DLX_EXinst_Mcompar__n0085_inst_cy_109/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0085_inst_lut4_6),
    .O(DLX_EXinst_Mcompar__n0085_inst_cy_108)
  );
  defparam DLX_EXinst_Mcompar__n0085_inst_lut4_61.INIT = 16'h8421;
  X_LUT4 DLX_EXinst_Mcompar__n0085_inst_lut4_61 (
    .ADR0(\DLX_IDinst_Imm[12] ),
    .ADR1(\DLX_IDinst_Imm[13] ),
    .ADR2(DLX_IDinst_reg_out_A[12]),
    .ADR3(DLX_IDinst_reg_out_A[13]),
    .O(DLX_EXinst_Mcompar__n0085_inst_lut4_6)
  );
  defparam DLX_EXinst_Mcompar__n0085_inst_lut4_71.INIT = 16'h8421;
  X_LUT4 DLX_EXinst_Mcompar__n0085_inst_lut4_71 (
    .ADR0(DLX_IDinst_reg_out_A[15]),
    .ADR1(DLX_IDinst_reg_out_A[14]),
    .ADR2(\DLX_IDinst_Imm[15] ),
    .ADR3(\DLX_IDinst_Imm[14] ),
    .O(DLX_EXinst_Mcompar__n0085_inst_lut4_7)
  );
  X_BUF \DLX_EXinst_Mcompar__n0085_inst_cy_109/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0085_inst_cy_109/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0085_inst_cy_109)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0085_inst_cy_109_548 (
    .IA(\DLX_EXinst_Mcompar__n0085_inst_cy_109/LOGIC_ZERO ),
    .IB(DLX_EXinst_Mcompar__n0085_inst_cy_108),
    .SEL(DLX_EXinst_Mcompar__n0085_inst_lut4_7),
    .O(\DLX_EXinst_Mcompar__n0085_inst_cy_109/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0085_inst_cy_109/CYINIT_549  (
    .I(DLX_EXinst_Mcompar__n0085_inst_cy_107),
    .O(\DLX_EXinst_Mcompar__n0085_inst_cy_109/CYINIT )
  );
  X_ZERO \DLX_EXinst_Mcompar__n0085_inst_cy_111/LOGIC_ZERO_550  (
    .O(\DLX_EXinst_Mcompar__n0085_inst_cy_111/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0085_inst_cy_110_551 (
    .IA(\DLX_EXinst_Mcompar__n0085_inst_cy_111/LOGIC_ZERO ),
    .IB(\DLX_EXinst_Mcompar__n0085_inst_cy_111/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0085_inst_lut4_8),
    .O(DLX_EXinst_Mcompar__n0085_inst_cy_110)
  );
  defparam DLX_EXinst_Mcompar__n0085_inst_lut4_81.INIT = 16'hC003;
  X_LUT4 DLX_EXinst_Mcompar__n0085_inst_lut4_81 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[17]),
    .ADR2(\DLX_IDinst_Imm[31] ),
    .ADR3(DLX_IDinst_reg_out_A[16]),
    .O(DLX_EXinst_Mcompar__n0085_inst_lut4_8)
  );
  defparam DLX_EXinst_Mcompar__n0085_inst_lut4_91.INIT = 16'h8181;
  X_LUT4 DLX_EXinst_Mcompar__n0085_inst_lut4_91 (
    .ADR0(DLX_IDinst_reg_out_A[18]),
    .ADR1(\DLX_IDinst_Imm[31] ),
    .ADR2(DLX_IDinst_reg_out_A[19]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0085_inst_lut4_9)
  );
  X_BUF \DLX_EXinst_Mcompar__n0085_inst_cy_111/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0085_inst_cy_111/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0085_inst_cy_111)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0085_inst_cy_111_552 (
    .IA(\DLX_EXinst_Mcompar__n0085_inst_cy_111/LOGIC_ZERO ),
    .IB(DLX_EXinst_Mcompar__n0085_inst_cy_110),
    .SEL(DLX_EXinst_Mcompar__n0085_inst_lut4_9),
    .O(\DLX_EXinst_Mcompar__n0085_inst_cy_111/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0085_inst_cy_111/CYINIT_553  (
    .I(DLX_EXinst_Mcompar__n0085_inst_cy_109),
    .O(\DLX_EXinst_Mcompar__n0085_inst_cy_111/CYINIT )
  );
  X_ZERO \DLX_EXinst_Mcompar__n0085_inst_cy_113/LOGIC_ZERO_554  (
    .O(\DLX_EXinst_Mcompar__n0085_inst_cy_113/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0085_inst_cy_112_555 (
    .IA(\DLX_EXinst_Mcompar__n0085_inst_cy_113/LOGIC_ZERO ),
    .IB(\DLX_EXinst_Mcompar__n0085_inst_cy_113/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0085_inst_lut4_10),
    .O(DLX_EXinst_Mcompar__n0085_inst_cy_112)
  );
  defparam DLX_EXinst_Mcompar__n0085_inst_lut4_101.INIT = 16'h8181;
  X_LUT4 DLX_EXinst_Mcompar__n0085_inst_lut4_101 (
    .ADR0(DLX_IDinst_reg_out_A[21]),
    .ADR1(\DLX_IDinst_Imm[31] ),
    .ADR2(DLX_IDinst_reg_out_A[20]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0085_inst_lut4_10)
  );
  defparam DLX_EXinst_Mcompar__n0085_inst_lut4_111.INIT = 16'h8811;
  X_LUT4 DLX_EXinst_Mcompar__n0085_inst_lut4_111 (
    .ADR0(DLX_IDinst_reg_out_A[22]),
    .ADR1(\DLX_IDinst_Imm[31] ),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[23]),
    .O(DLX_EXinst_Mcompar__n0085_inst_lut4_11)
  );
  X_BUF \DLX_EXinst_Mcompar__n0085_inst_cy_113/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0085_inst_cy_113/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0085_inst_cy_113)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0085_inst_cy_113_556 (
    .IA(\DLX_EXinst_Mcompar__n0085_inst_cy_113/LOGIC_ZERO ),
    .IB(DLX_EXinst_Mcompar__n0085_inst_cy_112),
    .SEL(DLX_EXinst_Mcompar__n0085_inst_lut4_11),
    .O(\DLX_EXinst_Mcompar__n0085_inst_cy_113/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0085_inst_cy_113/CYINIT_557  (
    .I(DLX_EXinst_Mcompar__n0085_inst_cy_111),
    .O(\DLX_EXinst_Mcompar__n0085_inst_cy_113/CYINIT )
  );
  X_ZERO \DLX_EXinst_Mcompar__n0085_inst_cy_115/LOGIC_ZERO_558  (
    .O(\DLX_EXinst_Mcompar__n0085_inst_cy_115/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0085_inst_cy_114_559 (
    .IA(\DLX_EXinst_Mcompar__n0085_inst_cy_115/LOGIC_ZERO ),
    .IB(\DLX_EXinst_Mcompar__n0085_inst_cy_115/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0085_inst_lut4_12),
    .O(DLX_EXinst_Mcompar__n0085_inst_cy_114)
  );
  defparam DLX_EXinst_Mcompar__n0085_inst_lut4_121.INIT = 16'h8181;
  X_LUT4 DLX_EXinst_Mcompar__n0085_inst_lut4_121 (
    .ADR0(\DLX_IDinst_Imm[31] ),
    .ADR1(DLX_IDinst_reg_out_A[25]),
    .ADR2(DLX_IDinst_reg_out_A[24]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0085_inst_lut4_12)
  );
  defparam DLX_EXinst_Mcompar__n0085_inst_lut4_131.INIT = 16'h8181;
  X_LUT4 DLX_EXinst_Mcompar__n0085_inst_lut4_131 (
    .ADR0(\DLX_IDinst_Imm[31] ),
    .ADR1(DLX_IDinst_reg_out_A[26]),
    .ADR2(DLX_IDinst_reg_out_A[27]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0085_inst_lut4_13)
  );
  X_BUF \DLX_EXinst_Mcompar__n0085_inst_cy_115/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0085_inst_cy_115/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0085_inst_cy_115)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0085_inst_cy_115_560 (
    .IA(\DLX_EXinst_Mcompar__n0085_inst_cy_115/LOGIC_ZERO ),
    .IB(DLX_EXinst_Mcompar__n0085_inst_cy_114),
    .SEL(DLX_EXinst_Mcompar__n0085_inst_lut4_13),
    .O(\DLX_EXinst_Mcompar__n0085_inst_cy_115/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0085_inst_cy_115/CYINIT_561  (
    .I(DLX_EXinst_Mcompar__n0085_inst_cy_113),
    .O(\DLX_EXinst_Mcompar__n0085_inst_cy_115/CYINIT )
  );
  X_ZERO \DLX_EXinst__n0085/LOGIC_ZERO_562  (
    .O(\DLX_EXinst__n0085/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0085_inst_cy_116_563 (
    .IA(\DLX_EXinst__n0085/LOGIC_ZERO ),
    .IB(\DLX_EXinst__n0085/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0085_inst_lut4_14),
    .O(DLX_EXinst_Mcompar__n0085_inst_cy_116)
  );
  defparam DLX_EXinst_Mcompar__n0085_inst_lut4_141.INIT = 16'hA005;
  X_LUT4 DLX_EXinst_Mcompar__n0085_inst_lut4_141 (
    .ADR0(DLX_IDinst_reg_out_A[29]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[28]),
    .ADR3(\DLX_IDinst_Imm[31] ),
    .O(DLX_EXinst_Mcompar__n0085_inst_lut4_14)
  );
  defparam DLX_EXinst_Mcompar__n0085_inst_lut4_151.INIT = 16'hA005;
  X_LUT4 DLX_EXinst_Mcompar__n0085_inst_lut4_151 (
    .ADR0(\DLX_IDinst_Imm[31] ),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(DLX_IDinst_reg_out_A[30]),
    .O(DLX_EXinst_Mcompar__n0085_inst_lut4_15)
  );
  X_BUF \DLX_EXinst__n0085/COUTUSED  (
    .I(\DLX_EXinst__n0085/CYMUXG ),
    .O(DLX_EXinst__n0085)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0085_inst_cy_117 (
    .IA(\DLX_EXinst__n0085/LOGIC_ZERO ),
    .IB(DLX_EXinst_Mcompar__n0085_inst_cy_116),
    .SEL(DLX_EXinst_Mcompar__n0085_inst_lut4_15),
    .O(\DLX_EXinst__n0085/CYMUXG )
  );
  X_BUF \DLX_EXinst__n0085/CYINIT_564  (
    .I(DLX_EXinst_Mcompar__n0085_inst_cy_115),
    .O(\DLX_EXinst__n0085/CYINIT )
  );
  X_ZERO \DLX_EXinst_Mcompar__n0093_inst_cy_199/LOGIC_ZERO_565  (
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_199/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_198_566 (
    .IA(DLX_IDinst_reg_out_A[0]),
    .IB(\DLX_EXinst_Mcompar__n0093_inst_cy_199/LOGIC_ZERO ),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_134),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_198)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1341.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1341 (
    .ADR0(DLX_IDinst_reg_out_A[0]),
    .ADR1(DLX_IDinst_IR_function_field_0_1),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_134)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1351.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1351 (
    .ADR0(DLX_IDinst_reg_out_A[1]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_IR_function_field_1_1),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_135)
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_199/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0093_inst_cy_199/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_199)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_199_567 (
    .IA(DLX_IDinst_reg_out_A[1]),
    .IB(DLX_EXinst_Mcompar__n0093_inst_cy_198),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_135),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_199/CYMUXG )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_200_568 (
    .IA(DLX_IDinst_reg_out_A[2]),
    .IB(\DLX_EXinst_Mcompar__n0093_inst_cy_201/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_136),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_200)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1361.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1361 (
    .ADR0(DLX_IDinst_reg_out_A[2]),
    .ADR1(DLX_IDinst_IR_function_field_2_1),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_136)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1371.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1371 (
    .ADR0(DLX_IDinst_reg_out_A[3]),
    .ADR1(DLX_IDinst_IR_function_field_3_1),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_137)
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_201/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0093_inst_cy_201/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_201)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_201_569 (
    .IA(DLX_IDinst_reg_out_A[3]),
    .IB(DLX_EXinst_Mcompar__n0093_inst_cy_200),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_137),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_201/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_201/CYINIT_570  (
    .I(DLX_EXinst_Mcompar__n0093_inst_cy_199),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_201/CYINIT )
  );
  defparam DLX_IFinst_NPC_7_1_571.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_7_1_571 (
    .I(\NPC_eff<7>/OD ),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\NPC_eff<7>/OFF/RST ),
    .O(DLX_IFinst_NPC_7_1)
  );
  X_OR2 \NPC_eff<7>/OFF/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\NPC_eff<7>/OFF/RST )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_202_572 (
    .IA(DLX_IDinst_reg_out_A[4]),
    .IB(\DLX_EXinst_Mcompar__n0093_inst_cy_203/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_138),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_202)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1381.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1381 (
    .ADR0(DLX_IDinst_reg_out_A[4]),
    .ADR1(DLX_IDinst_IR_function_field[4]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_138)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1391.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1391 (
    .ADR0(DLX_IDinst_reg_out_A[5]),
    .ADR1(\DLX_IDinst_Imm[5] ),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_139)
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_203/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0093_inst_cy_203/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_203)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_203_573 (
    .IA(DLX_IDinst_reg_out_A[5]),
    .IB(DLX_EXinst_Mcompar__n0093_inst_cy_202),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_139),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_203/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_203/CYINIT_574  (
    .I(DLX_EXinst_Mcompar__n0093_inst_cy_201),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_203/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_204_575 (
    .IA(DLX_IDinst_reg_out_A[6]),
    .IB(\DLX_EXinst_Mcompar__n0093_inst_cy_205/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_140),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_204)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1401.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1401 (
    .ADR0(DLX_IDinst_reg_out_A[6]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(\DLX_IDinst_Imm[6] ),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_140)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1411.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1411 (
    .ADR0(DLX_IDinst_reg_out_A[7]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(\DLX_IDinst_Imm[7] ),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_141)
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_205/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0093_inst_cy_205/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_205)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_205_576 (
    .IA(DLX_IDinst_reg_out_A[7]),
    .IB(DLX_EXinst_Mcompar__n0093_inst_cy_204),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_141),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_205/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_205/CYINIT_577  (
    .I(DLX_EXinst_Mcompar__n0093_inst_cy_203),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_205/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_206_578 (
    .IA(DLX_IDinst_reg_out_A[8]),
    .IB(\DLX_EXinst_Mcompar__n0093_inst_cy_207/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_142),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_206)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1421.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1421 (
    .ADR0(DLX_IDinst_reg_out_A[8]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(\DLX_IDinst_Imm[8] ),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_142)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1431.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1431 (
    .ADR0(DLX_IDinst_reg_out_A[9]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(\DLX_IDinst_Imm[9] ),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_143)
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_207/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0093_inst_cy_207/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_207)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_207_579 (
    .IA(DLX_IDinst_reg_out_A[9]),
    .IB(DLX_EXinst_Mcompar__n0093_inst_cy_206),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_143),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_207/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_207/CYINIT_580  (
    .I(DLX_EXinst_Mcompar__n0093_inst_cy_205),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_207/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_208_581 (
    .IA(DLX_IDinst_reg_out_A[10]),
    .IB(\DLX_EXinst_Mcompar__n0093_inst_cy_209/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_144),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_208)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1441.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1441 (
    .ADR0(DLX_IDinst_reg_out_A[10]),
    .ADR1(\DLX_IDinst_Imm[10] ),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_144)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1451.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1451 (
    .ADR0(DLX_IDinst_reg_out_A[11]),
    .ADR1(\DLX_IDinst_Imm[11] ),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_145)
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_209/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0093_inst_cy_209/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_209)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_209_582 (
    .IA(DLX_IDinst_reg_out_A[11]),
    .IB(DLX_EXinst_Mcompar__n0093_inst_cy_208),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_145),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_209/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_209/CYINIT_583  (
    .I(DLX_EXinst_Mcompar__n0093_inst_cy_207),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_209/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_210_584 (
    .IA(DLX_IDinst_reg_out_A[12]),
    .IB(\DLX_EXinst_Mcompar__n0093_inst_cy_211/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_146),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_210)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1461.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1461 (
    .ADR0(DLX_IDinst_reg_out_A[12]),
    .ADR1(VCC),
    .ADR2(\DLX_IDinst_Imm[12] ),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_146)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1471.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1471 (
    .ADR0(DLX_IDinst_reg_out_A[13]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(\DLX_IDinst_Imm[13] ),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_147)
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_211/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0093_inst_cy_211/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_211)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_211_585 (
    .IA(DLX_IDinst_reg_out_A[13]),
    .IB(DLX_EXinst_Mcompar__n0093_inst_cy_210),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_147),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_211/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_211/CYINIT_586  (
    .I(DLX_EXinst_Mcompar__n0093_inst_cy_209),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_211/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_212_587 (
    .IA(DLX_IDinst_reg_out_A[14]),
    .IB(\DLX_EXinst_Mcompar__n0093_inst_cy_213/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_148),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_212)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1481.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1481 (
    .ADR0(DLX_IDinst_reg_out_A[14]),
    .ADR1(VCC),
    .ADR2(\DLX_IDinst_Imm[14] ),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_148)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1491.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1491 (
    .ADR0(DLX_IDinst_reg_out_A[15]),
    .ADR1(\DLX_IDinst_Imm[15] ),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_149)
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_213/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0093_inst_cy_213/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_213)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_213_588 (
    .IA(DLX_IDinst_reg_out_A[15]),
    .IB(DLX_EXinst_Mcompar__n0093_inst_cy_212),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_149),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_213/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_213/CYINIT_589  (
    .I(DLX_EXinst_Mcompar__n0093_inst_cy_211),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_213/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_214_590 (
    .IA(DLX_IDinst_reg_out_A[16]),
    .IB(\DLX_EXinst_Mcompar__n0093_inst_cy_215/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_150),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_214)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1501.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1501 (
    .ADR0(DLX_IDinst_reg_out_A[16]),
    .ADR1(DLX_IDinst_Imm_31_1),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_150)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1511.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1511 (
    .ADR0(DLX_IDinst_reg_out_A[17]),
    .ADR1(DLX_IDinst_Imm_31_1),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_151)
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_215/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0093_inst_cy_215/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_215)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_215_591 (
    .IA(DLX_IDinst_reg_out_A[17]),
    .IB(DLX_EXinst_Mcompar__n0093_inst_cy_214),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_151),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_215/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_215/CYINIT_592  (
    .I(DLX_EXinst_Mcompar__n0093_inst_cy_213),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_215/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_216_593 (
    .IA(DLX_IDinst_reg_out_A[18]),
    .IB(\DLX_EXinst_Mcompar__n0093_inst_cy_217/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_152),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_216)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1521.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1521 (
    .ADR0(DLX_IDinst_reg_out_A[18]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_Imm_31_1),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_152)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1531.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1531 (
    .ADR0(DLX_IDinst_reg_out_A[19]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_Imm_31_1),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_153)
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_217/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0093_inst_cy_217/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_217)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_217_594 (
    .IA(DLX_IDinst_reg_out_A[19]),
    .IB(DLX_EXinst_Mcompar__n0093_inst_cy_216),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_153),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_217/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_217/CYINIT_595  (
    .I(DLX_EXinst_Mcompar__n0093_inst_cy_215),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_217/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_218_596 (
    .IA(DLX_IDinst_reg_out_A[20]),
    .IB(\DLX_EXinst_Mcompar__n0093_inst_cy_219/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_154),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_218)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1541.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1541 (
    .ADR0(DLX_IDinst_reg_out_A[20]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_Imm_31_1),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_154)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1551.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1551 (
    .ADR0(DLX_IDinst_reg_out_A[21]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_Imm_31_1),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_155)
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_219/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0093_inst_cy_219/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_219)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_219_597 (
    .IA(DLX_IDinst_reg_out_A[21]),
    .IB(DLX_EXinst_Mcompar__n0093_inst_cy_218),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_155),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_219/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_219/CYINIT_598  (
    .I(DLX_EXinst_Mcompar__n0093_inst_cy_217),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_219/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_220_599 (
    .IA(DLX_IDinst_reg_out_A[22]),
    .IB(\DLX_EXinst_Mcompar__n0093_inst_cy_221/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_156),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_220)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1561.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1561 (
    .ADR0(DLX_IDinst_reg_out_A[22]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_Imm_31_1),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_156)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1571.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1571 (
    .ADR0(DLX_IDinst_reg_out_A[23]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_Imm_31_1),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_157)
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_221/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0093_inst_cy_221/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_221)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_221_600 (
    .IA(DLX_IDinst_reg_out_A[23]),
    .IB(DLX_EXinst_Mcompar__n0093_inst_cy_220),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_157),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_221/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_221/CYINIT_601  (
    .I(DLX_EXinst_Mcompar__n0093_inst_cy_219),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_221/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_222_602 (
    .IA(DLX_IDinst_reg_out_A[24]),
    .IB(\DLX_EXinst_Mcompar__n0093_inst_cy_223/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_158),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_222)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1581.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1581 (
    .ADR0(DLX_IDinst_reg_out_A[24]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_Imm_31_1),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_158)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1591.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1591 (
    .ADR0(DLX_IDinst_reg_out_A[25]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_Imm_31_1),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_159)
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_223/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0093_inst_cy_223/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_223)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_223_603 (
    .IA(DLX_IDinst_reg_out_A[25]),
    .IB(DLX_EXinst_Mcompar__n0093_inst_cy_222),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_159),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_223/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_223/CYINIT_604  (
    .I(DLX_EXinst_Mcompar__n0093_inst_cy_221),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_223/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_224_605 (
    .IA(DLX_IDinst_reg_out_A[26]),
    .IB(\DLX_EXinst_Mcompar__n0093_inst_cy_225/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_160),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_224)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1601.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1601 (
    .ADR0(DLX_IDinst_reg_out_A[26]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_Imm_31_1),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_160)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1611.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1611 (
    .ADR0(DLX_IDinst_reg_out_A[27]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_Imm_31_1),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_161)
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_225/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0093_inst_cy_225/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_225)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_225_606 (
    .IA(DLX_IDinst_reg_out_A[27]),
    .IB(DLX_EXinst_Mcompar__n0093_inst_cy_224),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_161),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_225/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_225/CYINIT_607  (
    .I(DLX_EXinst_Mcompar__n0093_inst_cy_223),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_225/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_226_608 (
    .IA(DLX_IDinst_reg_out_A[28]),
    .IB(\DLX_EXinst_Mcompar__n0093_inst_cy_227/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_162),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_226)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1621.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1621 (
    .ADR0(DLX_IDinst_reg_out_A[28]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_Imm_31_1),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_162)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1631.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1631 (
    .ADR0(DLX_IDinst_reg_out_A[29]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_Imm_31_1),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_163)
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_227/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0093_inst_cy_227/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_227)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_227_609 (
    .IA(DLX_IDinst_reg_out_A[29]),
    .IB(DLX_EXinst_Mcompar__n0093_inst_cy_226),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_163),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_227/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_227/CYINIT_610  (
    .I(DLX_EXinst_Mcompar__n0093_inst_cy_225),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_227/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_228_611 (
    .IA(DLX_IDinst_reg_out_A[30]),
    .IB(\CHOICE1126/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_164),
    .O(\CHOICE1126/CYMUXF )
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1641.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1641 (
    .ADR0(DLX_IDinst_reg_out_A[30]),
    .ADR1(DLX_IDinst_Imm_31_1),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_164)
  );
  defparam \DLX_EXinst_Mshift__n0024_Sh<28>11 .INIT = 16'hA808;
  X_LUT4 \DLX_EXinst_Mshift__n0024_Sh<28>11  (
    .ADR0(DLX_IDinst_IR_function_field_1_1),
    .ADR1(DLX_IDinst_reg_out_A[30]),
    .ADR2(DLX_IDinst_IR_function_field_0_1),
    .ADR3(DLX_IDinst_reg_out_A[31]),
    .O(\CHOICE1126/GROM )
  );
  X_BUF \CHOICE1126/XBUSED  (
    .I(\CHOICE1126/CYMUXF ),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_228)
  );
  X_BUF \CHOICE1126/YUSED  (
    .I(\CHOICE1126/GROM ),
    .O(CHOICE1126)
  );
  X_BUF \CHOICE1126/CYINIT_612  (
    .I(DLX_EXinst_Mcompar__n0093_inst_cy_227),
    .O(\CHOICE1126/CYINIT )
  );
  X_ONE \DLX_IDinst_Mcompar__n0077_inst_cy_263/LOGIC_ONE_613  (
    .O(\DLX_IDinst_Mcompar__n0077_inst_cy_263/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mcompar__n0077_inst_cy_263/LOGIC_ZERO_614  (
    .O(\DLX_IDinst_Mcompar__n0077_inst_cy_263/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mcompar__n0077_inst_cy_262_615 (
    .IA(\DLX_IDinst_Mcompar__n0077_inst_cy_263/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mcompar__n0077_inst_cy_263/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mcompar__n0077_inst_lut4_40),
    .O(DLX_IDinst_Mcompar__n0077_inst_cy_262)
  );
  defparam DLX_IDinst_Mcompar__n0077_inst_lut4_401.INIT = 16'h8241;
  X_LUT4 DLX_IDinst_Mcompar__n0077_inst_lut4_401 (
    .ADR0(DLX_IDinst_regA_index[0]),
    .ADR1(DLX_reg_dst_of_MEM[1]),
    .ADR2(DLX_IDinst_regA_index[1]),
    .ADR3(DLX_reg_dst_of_MEM[0]),
    .O(DLX_IDinst_Mcompar__n0077_inst_lut4_40)
  );
  defparam DLX_IDinst_Mcompar__n0077_inst_lut4_411.INIT = 16'h8241;
  X_LUT4 DLX_IDinst_Mcompar__n0077_inst_lut4_411 (
    .ADR0(DLX_IDinst_regA_index[3]),
    .ADR1(DLX_IDinst_regA_index[2]),
    .ADR2(DLX_reg_dst_of_MEM[2]),
    .ADR3(DLX_reg_dst_of_MEM[3]),
    .O(DLX_IDinst_Mcompar__n0077_inst_lut4_41)
  );
  X_BUF \DLX_IDinst_Mcompar__n0077_inst_cy_263/COUTUSED  (
    .I(\DLX_IDinst_Mcompar__n0077_inst_cy_263/CYMUXG ),
    .O(DLX_IDinst_Mcompar__n0077_inst_cy_263)
  );
  X_MUX2 DLX_IDinst_Mcompar__n0077_inst_cy_263_616 (
    .IA(\DLX_IDinst_Mcompar__n0077_inst_cy_263/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mcompar__n0077_inst_cy_262),
    .SEL(DLX_IDinst_Mcompar__n0077_inst_lut4_41),
    .O(\DLX_IDinst_Mcompar__n0077_inst_cy_263/CYMUXG )
  );
  X_ZERO \DLX_IDinst__n0077/LOGIC_ZERO_617  (
    .O(\DLX_IDinst__n0077/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mcompar__n0077_inst_cy_264 (
    .IA(\DLX_IDinst__n0077/LOGIC_ZERO ),
    .IB(\DLX_IDinst__n0077/CYINIT ),
    .SEL(DLX_IDinst_Mcompar__n0077_inst_lut4_42),
    .O(\DLX_IDinst__n0077/CYMUXF )
  );
  defparam DLX_IDinst_Mcompar__n0077_inst_lut4_421.INIT = 16'hAA55;
  X_LUT4 DLX_IDinst_Mcompar__n0077_inst_lut4_421 (
    .ADR0(DLX_reg_dst_of_MEM[4]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_regA_index[4]),
    .O(DLX_IDinst_Mcompar__n0077_inst_lut4_42)
  );
  X_BUF \DLX_IDinst__n0077/XBUSED  (
    .I(\DLX_IDinst__n0077/CYMUXF ),
    .O(DLX_IDinst__n0077)
  );
  X_BUF \DLX_IDinst__n0077/CYINIT_618  (
    .I(DLX_IDinst_Mcompar__n0077_inst_cy_263),
    .O(\DLX_IDinst__n0077/CYINIT )
  );
  X_MUX2 DLX_EXinst_Maddsub__n0016_inst_cy_70_619 (
    .IA(DLX_IDinst_reg_out_A[0]),
    .IB(\DLX_EXinst__n0016<0>/CYINIT ),
    .SEL(DLX_EXinst_Maddsub__n0016_inst_lut3_6),
    .O(DLX_EXinst_Maddsub__n0016_inst_cy_70)
  );
  X_XOR2 DLX_EXinst_Maddsub__n0016_inst_sum_70 (
    .I0(\DLX_EXinst__n0016<0>/CYINIT ),
    .I1(DLX_EXinst_Maddsub__n0016_inst_lut3_6),
    .O(\DLX_EXinst__n0016<0>/XORF )
  );
  defparam DLX_EXinst_Maddsub__n0016_inst_lut3_61.INIT = 16'hA55A;
  X_LUT4 DLX_EXinst_Maddsub__n0016_inst_lut3_61 (
    .ADR0(DLX_IDinst_reg_out_A[0]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst__n0017[0]),
    .ADR3(N108704),
    .O(DLX_EXinst_Maddsub__n0016_inst_lut3_6)
  );
  defparam DLX_EXinst_Maddsub__n0016_inst_lut3_71.INIT = 16'hA55A;
  X_LUT4 DLX_EXinst_Maddsub__n0016_inst_lut3_71 (
    .ADR0(DLX_IDinst_reg_out_A[1]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst__n0017[1]),
    .ADR3(N108704),
    .O(DLX_EXinst_Maddsub__n0016_inst_lut3_7)
  );
  X_BUF \DLX_EXinst__n0016<0>/COUTUSED  (
    .I(\DLX_EXinst__n0016<0>/CYMUXG ),
    .O(DLX_EXinst_Maddsub__n0016_inst_cy_71)
  );
  X_BUF \DLX_EXinst__n0016<0>/XUSED  (
    .I(\DLX_EXinst__n0016<0>/XORF ),
    .O(DLX_EXinst__n0016[0])
  );
  X_BUF \DLX_EXinst__n0016<0>/YUSED  (
    .I(\DLX_EXinst__n0016<0>/XORG ),
    .O(DLX_EXinst__n0016[1])
  );
  X_MUX2 DLX_EXinst_Maddsub__n0016_inst_cy_71_620 (
    .IA(DLX_IDinst_reg_out_A[1]),
    .IB(DLX_EXinst_Maddsub__n0016_inst_cy_70),
    .SEL(DLX_EXinst_Maddsub__n0016_inst_lut3_7),
    .O(\DLX_EXinst__n0016<0>/CYMUXG )
  );
  X_XOR2 DLX_EXinst_Maddsub__n0016_inst_sum_71 (
    .I0(DLX_EXinst_Maddsub__n0016_inst_cy_70),
    .I1(DLX_EXinst_Maddsub__n0016_inst_lut3_7),
    .O(\DLX_EXinst__n0016<0>/XORG )
  );
  X_BUF \DLX_EXinst__n0016<0>/CYINIT_621  (
    .I(N108704),
    .O(\DLX_EXinst__n0016<0>/CYINIT )
  );
  X_MUX2 DLX_EXinst_Maddsub__n0016_inst_cy_72_622 (
    .IA(DLX_IDinst_reg_out_A[2]),
    .IB(\DLX_EXinst__n0016<2>/CYINIT ),
    .SEL(DLX_EXinst_Maddsub__n0016_inst_lut3_8),
    .O(DLX_EXinst_Maddsub__n0016_inst_cy_72)
  );
  X_XOR2 DLX_EXinst_Maddsub__n0016_inst_sum_72 (
    .I0(\DLX_EXinst__n0016<2>/CYINIT ),
    .I1(DLX_EXinst_Maddsub__n0016_inst_lut3_8),
    .O(\DLX_EXinst__n0016<2>/XORF )
  );
  defparam DLX_EXinst_Maddsub__n0016_inst_lut3_81.INIT = 16'h9696;
  X_LUT4 DLX_EXinst_Maddsub__n0016_inst_lut3_81 (
    .ADR0(DLX_IDinst_reg_out_A[2]),
    .ADR1(DLX_EXinst__n0017[2]),
    .ADR2(N108704),
    .ADR3(VCC),
    .O(DLX_EXinst_Maddsub__n0016_inst_lut3_8)
  );
  defparam DLX_EXinst_Maddsub__n0016_inst_lut3_91.INIT = 16'h9696;
  X_LUT4 DLX_EXinst_Maddsub__n0016_inst_lut3_91 (
    .ADR0(DLX_IDinst_reg_out_A[3]),
    .ADR1(N108704),
    .ADR2(DLX_EXinst__n0017[3]),
    .ADR3(VCC),
    .O(DLX_EXinst_Maddsub__n0016_inst_lut3_9)
  );
  X_BUF \DLX_EXinst__n0016<2>/COUTUSED  (
    .I(\DLX_EXinst__n0016<2>/CYMUXG ),
    .O(DLX_EXinst_Maddsub__n0016_inst_cy_73)
  );
  X_BUF \DLX_EXinst__n0016<2>/XUSED  (
    .I(\DLX_EXinst__n0016<2>/XORF ),
    .O(DLX_EXinst__n0016[2])
  );
  X_BUF \DLX_EXinst__n0016<2>/YUSED  (
    .I(\DLX_EXinst__n0016<2>/XORG ),
    .O(DLX_EXinst__n0016[3])
  );
  X_MUX2 DLX_EXinst_Maddsub__n0016_inst_cy_73_623 (
    .IA(DLX_IDinst_reg_out_A[3]),
    .IB(DLX_EXinst_Maddsub__n0016_inst_cy_72),
    .SEL(DLX_EXinst_Maddsub__n0016_inst_lut3_9),
    .O(\DLX_EXinst__n0016<2>/CYMUXG )
  );
  X_XOR2 DLX_EXinst_Maddsub__n0016_inst_sum_73 (
    .I0(DLX_EXinst_Maddsub__n0016_inst_cy_72),
    .I1(DLX_EXinst_Maddsub__n0016_inst_lut3_9),
    .O(\DLX_EXinst__n0016<2>/XORG )
  );
  X_BUF \DLX_EXinst__n0016<2>/CYINIT_624  (
    .I(DLX_EXinst_Maddsub__n0016_inst_cy_71),
    .O(\DLX_EXinst__n0016<2>/CYINIT )
  );
  X_MUX2 DLX_EXinst_Maddsub__n0016_inst_cy_74_625 (
    .IA(DLX_IDinst_reg_out_A[4]),
    .IB(\DLX_EXinst__n0016<4>/CYINIT ),
    .SEL(DLX_EXinst_Maddsub__n0016_inst_lut3_10),
    .O(DLX_EXinst_Maddsub__n0016_inst_cy_74)
  );
  X_XOR2 DLX_EXinst_Maddsub__n0016_inst_sum_74 (
    .I0(\DLX_EXinst__n0016<4>/CYINIT ),
    .I1(DLX_EXinst_Maddsub__n0016_inst_lut3_10),
    .O(\DLX_EXinst__n0016<4>/XORF )
  );
  defparam DLX_EXinst_Maddsub__n0016_inst_lut3_101.INIT = 16'h9966;
  X_LUT4 DLX_EXinst_Maddsub__n0016_inst_lut3_101 (
    .ADR0(DLX_IDinst_reg_out_A[4]),
    .ADR1(N108704),
    .ADR2(VCC),
    .ADR3(DLX_EXinst__n0017[4]),
    .O(DLX_EXinst_Maddsub__n0016_inst_lut3_10)
  );
  defparam DLX_EXinst_Maddsub__n0016_inst_lut3_111.INIT = 16'h9966;
  X_LUT4 DLX_EXinst_Maddsub__n0016_inst_lut3_111 (
    .ADR0(DLX_IDinst_reg_out_A[5]),
    .ADR1(N108704),
    .ADR2(VCC),
    .ADR3(DLX_EXinst__n0017[5]),
    .O(DLX_EXinst_Maddsub__n0016_inst_lut3_11)
  );
  X_BUF \DLX_EXinst__n0016<4>/COUTUSED  (
    .I(\DLX_EXinst__n0016<4>/CYMUXG ),
    .O(DLX_EXinst_Maddsub__n0016_inst_cy_75)
  );
  X_BUF \DLX_EXinst__n0016<4>/XUSED  (
    .I(\DLX_EXinst__n0016<4>/XORF ),
    .O(DLX_EXinst__n0016[4])
  );
  X_BUF \DLX_EXinst__n0016<4>/YUSED  (
    .I(\DLX_EXinst__n0016<4>/XORG ),
    .O(DLX_EXinst__n0016[5])
  );
  X_MUX2 DLX_EXinst_Maddsub__n0016_inst_cy_75_626 (
    .IA(DLX_IDinst_reg_out_A[5]),
    .IB(DLX_EXinst_Maddsub__n0016_inst_cy_74),
    .SEL(DLX_EXinst_Maddsub__n0016_inst_lut3_11),
    .O(\DLX_EXinst__n0016<4>/CYMUXG )
  );
  X_XOR2 DLX_EXinst_Maddsub__n0016_inst_sum_75 (
    .I0(DLX_EXinst_Maddsub__n0016_inst_cy_74),
    .I1(DLX_EXinst_Maddsub__n0016_inst_lut3_11),
    .O(\DLX_EXinst__n0016<4>/XORG )
  );
  X_BUF \DLX_EXinst__n0016<4>/CYINIT_627  (
    .I(DLX_EXinst_Maddsub__n0016_inst_cy_73),
    .O(\DLX_EXinst__n0016<4>/CYINIT )
  );
  X_MUX2 DLX_EXinst_Maddsub__n0016_inst_cy_76_628 (
    .IA(DLX_IDinst_reg_out_A[6]),
    .IB(\DLX_EXinst__n0016<6>/CYINIT ),
    .SEL(DLX_EXinst_Maddsub__n0016_inst_lut3_12),
    .O(DLX_EXinst_Maddsub__n0016_inst_cy_76)
  );
  X_XOR2 DLX_EXinst_Maddsub__n0016_inst_sum_76 (
    .I0(\DLX_EXinst__n0016<6>/CYINIT ),
    .I1(DLX_EXinst_Maddsub__n0016_inst_lut3_12),
    .O(\DLX_EXinst__n0016<6>/XORF )
  );
  defparam DLX_EXinst_Maddsub__n0016_inst_lut3_121.INIT = 16'h9696;
  X_LUT4 DLX_EXinst_Maddsub__n0016_inst_lut3_121 (
    .ADR0(DLX_IDinst_reg_out_A[6]),
    .ADR1(N108704),
    .ADR2(DLX_EXinst__n0017[6]),
    .ADR3(VCC),
    .O(DLX_EXinst_Maddsub__n0016_inst_lut3_12)
  );
  defparam DLX_EXinst_Maddsub__n0016_inst_lut3_131.INIT = 16'h9696;
  X_LUT4 DLX_EXinst_Maddsub__n0016_inst_lut3_131 (
    .ADR0(DLX_IDinst_reg_out_A[7]),
    .ADR1(N108704),
    .ADR2(DLX_EXinst__n0017[7]),
    .ADR3(VCC),
    .O(DLX_EXinst_Maddsub__n0016_inst_lut3_13)
  );
  X_BUF \DLX_EXinst__n0016<6>/COUTUSED  (
    .I(\DLX_EXinst__n0016<6>/CYMUXG ),
    .O(DLX_EXinst_Maddsub__n0016_inst_cy_77)
  );
  X_BUF \DLX_EXinst__n0016<6>/XUSED  (
    .I(\DLX_EXinst__n0016<6>/XORF ),
    .O(DLX_EXinst__n0016[6])
  );
  X_BUF \DLX_EXinst__n0016<6>/YUSED  (
    .I(\DLX_EXinst__n0016<6>/XORG ),
    .O(DLX_EXinst__n0016[7])
  );
  X_MUX2 DLX_EXinst_Maddsub__n0016_inst_cy_77_629 (
    .IA(DLX_IDinst_reg_out_A[7]),
    .IB(DLX_EXinst_Maddsub__n0016_inst_cy_76),
    .SEL(DLX_EXinst_Maddsub__n0016_inst_lut3_13),
    .O(\DLX_EXinst__n0016<6>/CYMUXG )
  );
  X_XOR2 DLX_EXinst_Maddsub__n0016_inst_sum_77 (
    .I0(DLX_EXinst_Maddsub__n0016_inst_cy_76),
    .I1(DLX_EXinst_Maddsub__n0016_inst_lut3_13),
    .O(\DLX_EXinst__n0016<6>/XORG )
  );
  X_BUF \DLX_EXinst__n0016<6>/CYINIT_630  (
    .I(DLX_EXinst_Maddsub__n0016_inst_cy_75),
    .O(\DLX_EXinst__n0016<6>/CYINIT )
  );
  X_MUX2 DLX_EXinst_Maddsub__n0016_inst_cy_78_631 (
    .IA(DLX_IDinst_reg_out_A[8]),
    .IB(\DLX_EXinst__n0016<8>/CYINIT ),
    .SEL(DLX_EXinst_Maddsub__n0016_inst_lut3_14),
    .O(DLX_EXinst_Maddsub__n0016_inst_cy_78)
  );
  X_XOR2 DLX_EXinst_Maddsub__n0016_inst_sum_78 (
    .I0(\DLX_EXinst__n0016<8>/CYINIT ),
    .I1(DLX_EXinst_Maddsub__n0016_inst_lut3_14),
    .O(\DLX_EXinst__n0016<8>/XORF )
  );
  defparam DLX_EXinst_Maddsub__n0016_inst_lut3_141.INIT = 16'hA55A;
  X_LUT4 DLX_EXinst_Maddsub__n0016_inst_lut3_141 (
    .ADR0(DLX_IDinst_reg_out_A[8]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst__n0017[8]),
    .ADR3(N108704),
    .O(DLX_EXinst_Maddsub__n0016_inst_lut3_14)
  );
  defparam DLX_EXinst_Maddsub__n0016_inst_lut3_151.INIT = 16'hA55A;
  X_LUT4 DLX_EXinst_Maddsub__n0016_inst_lut3_151 (
    .ADR0(DLX_IDinst_reg_out_A[9]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst__n0017[9]),
    .ADR3(N108704),
    .O(DLX_EXinst_Maddsub__n0016_inst_lut3_15)
  );
  X_BUF \DLX_EXinst__n0016<8>/COUTUSED  (
    .I(\DLX_EXinst__n0016<8>/CYMUXG ),
    .O(DLX_EXinst_Maddsub__n0016_inst_cy_79)
  );
  X_BUF \DLX_EXinst__n0016<8>/XUSED  (
    .I(\DLX_EXinst__n0016<8>/XORF ),
    .O(DLX_EXinst__n0016[8])
  );
  X_BUF \DLX_EXinst__n0016<8>/YUSED  (
    .I(\DLX_EXinst__n0016<8>/XORG ),
    .O(DLX_EXinst__n0016[9])
  );
  X_MUX2 DLX_EXinst_Maddsub__n0016_inst_cy_79_632 (
    .IA(DLX_IDinst_reg_out_A[9]),
    .IB(DLX_EXinst_Maddsub__n0016_inst_cy_78),
    .SEL(DLX_EXinst_Maddsub__n0016_inst_lut3_15),
    .O(\DLX_EXinst__n0016<8>/CYMUXG )
  );
  X_XOR2 DLX_EXinst_Maddsub__n0016_inst_sum_79 (
    .I0(DLX_EXinst_Maddsub__n0016_inst_cy_78),
    .I1(DLX_EXinst_Maddsub__n0016_inst_lut3_15),
    .O(\DLX_EXinst__n0016<8>/XORG )
  );
  X_BUF \DLX_EXinst__n0016<8>/CYINIT_633  (
    .I(DLX_EXinst_Maddsub__n0016_inst_cy_77),
    .O(\DLX_EXinst__n0016<8>/CYINIT )
  );
  X_MUX2 DLX_EXinst_Maddsub__n0016_inst_cy_80_634 (
    .IA(DLX_IDinst_reg_out_A[10]),
    .IB(\DLX_EXinst__n0016<10>/CYINIT ),
    .SEL(DLX_EXinst_Maddsub__n0016_inst_lut3_16),
    .O(DLX_EXinst_Maddsub__n0016_inst_cy_80)
  );
  X_XOR2 DLX_EXinst_Maddsub__n0016_inst_sum_80 (
    .I0(\DLX_EXinst__n0016<10>/CYINIT ),
    .I1(DLX_EXinst_Maddsub__n0016_inst_lut3_16),
    .O(\DLX_EXinst__n0016<10>/XORF )
  );
  defparam DLX_EXinst_Maddsub__n0016_inst_lut3_161.INIT = 16'h9966;
  X_LUT4 DLX_EXinst_Maddsub__n0016_inst_lut3_161 (
    .ADR0(DLX_IDinst_reg_out_A[10]),
    .ADR1(DLX_EXinst__n0017[10]),
    .ADR2(VCC),
    .ADR3(N108704),
    .O(DLX_EXinst_Maddsub__n0016_inst_lut3_16)
  );
  defparam DLX_EXinst_Maddsub__n0016_inst_lut3_171.INIT = 16'h9966;
  X_LUT4 DLX_EXinst_Maddsub__n0016_inst_lut3_171 (
    .ADR0(DLX_IDinst_reg_out_A[11]),
    .ADR1(DLX_EXinst__n0017[11]),
    .ADR2(VCC),
    .ADR3(N108704),
    .O(DLX_EXinst_Maddsub__n0016_inst_lut3_17)
  );
  X_BUF \DLX_EXinst__n0016<10>/COUTUSED  (
    .I(\DLX_EXinst__n0016<10>/CYMUXG ),
    .O(DLX_EXinst_Maddsub__n0016_inst_cy_81)
  );
  X_BUF \DLX_EXinst__n0016<10>/XUSED  (
    .I(\DLX_EXinst__n0016<10>/XORF ),
    .O(DLX_EXinst__n0016[10])
  );
  X_BUF \DLX_EXinst__n0016<10>/YUSED  (
    .I(\DLX_EXinst__n0016<10>/XORG ),
    .O(DLX_EXinst__n0016[11])
  );
  X_MUX2 DLX_EXinst_Maddsub__n0016_inst_cy_81_635 (
    .IA(DLX_IDinst_reg_out_A[11]),
    .IB(DLX_EXinst_Maddsub__n0016_inst_cy_80),
    .SEL(DLX_EXinst_Maddsub__n0016_inst_lut3_17),
    .O(\DLX_EXinst__n0016<10>/CYMUXG )
  );
  X_XOR2 DLX_EXinst_Maddsub__n0016_inst_sum_81 (
    .I0(DLX_EXinst_Maddsub__n0016_inst_cy_80),
    .I1(DLX_EXinst_Maddsub__n0016_inst_lut3_17),
    .O(\DLX_EXinst__n0016<10>/XORG )
  );
  X_BUF \DLX_EXinst__n0016<10>/CYINIT_636  (
    .I(DLX_EXinst_Maddsub__n0016_inst_cy_79),
    .O(\DLX_EXinst__n0016<10>/CYINIT )
  );
  defparam DLX_IFinst_NPC_8_1_637.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_8_1_637 (
    .I(\NPC_eff<8>/OD ),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\NPC_eff<8>/OFF/RST ),
    .O(DLX_IFinst_NPC_8_1)
  );
  X_OR2 \NPC_eff<8>/OFF/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\NPC_eff<8>/OFF/RST )
  );
  X_MUX2 DLX_EXinst_Maddsub__n0016_inst_cy_82_638 (
    .IA(DLX_IDinst_reg_out_A[12]),
    .IB(\DLX_EXinst__n0016<12>/CYINIT ),
    .SEL(DLX_EXinst_Maddsub__n0016_inst_lut3_18),
    .O(DLX_EXinst_Maddsub__n0016_inst_cy_82)
  );
  X_XOR2 DLX_EXinst_Maddsub__n0016_inst_sum_82 (
    .I0(\DLX_EXinst__n0016<12>/CYINIT ),
    .I1(DLX_EXinst_Maddsub__n0016_inst_lut3_18),
    .O(\DLX_EXinst__n0016<12>/XORF )
  );
  defparam DLX_EXinst_Maddsub__n0016_inst_lut3_181.INIT = 16'hA55A;
  X_LUT4 DLX_EXinst_Maddsub__n0016_inst_lut3_181 (
    .ADR0(DLX_IDinst_reg_out_A[12]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst__n0017[12]),
    .ADR3(N108704),
    .O(DLX_EXinst_Maddsub__n0016_inst_lut3_18)
  );
  defparam DLX_EXinst_Maddsub__n0016_inst_lut3_191.INIT = 16'h9966;
  X_LUT4 DLX_EXinst_Maddsub__n0016_inst_lut3_191 (
    .ADR0(DLX_IDinst_reg_out_A[13]),
    .ADR1(DLX_EXinst__n0017[13]),
    .ADR2(VCC),
    .ADR3(N108704),
    .O(DLX_EXinst_Maddsub__n0016_inst_lut3_19)
  );
  X_BUF \DLX_EXinst__n0016<12>/COUTUSED  (
    .I(\DLX_EXinst__n0016<12>/CYMUXG ),
    .O(DLX_EXinst_Maddsub__n0016_inst_cy_83)
  );
  X_BUF \DLX_EXinst__n0016<12>/XUSED  (
    .I(\DLX_EXinst__n0016<12>/XORF ),
    .O(DLX_EXinst__n0016[12])
  );
  X_BUF \DLX_EXinst__n0016<12>/YUSED  (
    .I(\DLX_EXinst__n0016<12>/XORG ),
    .O(DLX_EXinst__n0016[13])
  );
  X_MUX2 DLX_EXinst_Maddsub__n0016_inst_cy_83_639 (
    .IA(DLX_IDinst_reg_out_A[13]),
    .IB(DLX_EXinst_Maddsub__n0016_inst_cy_82),
    .SEL(DLX_EXinst_Maddsub__n0016_inst_lut3_19),
    .O(\DLX_EXinst__n0016<12>/CYMUXG )
  );
  X_XOR2 DLX_EXinst_Maddsub__n0016_inst_sum_83 (
    .I0(DLX_EXinst_Maddsub__n0016_inst_cy_82),
    .I1(DLX_EXinst_Maddsub__n0016_inst_lut3_19),
    .O(\DLX_EXinst__n0016<12>/XORG )
  );
  X_BUF \DLX_EXinst__n0016<12>/CYINIT_640  (
    .I(DLX_EXinst_Maddsub__n0016_inst_cy_81),
    .O(\DLX_EXinst__n0016<12>/CYINIT )
  );
  X_MUX2 DLX_EXinst_Maddsub__n0016_inst_cy_84_641 (
    .IA(DLX_IDinst_reg_out_A[14]),
    .IB(\DLX_EXinst__n0016<14>/CYINIT ),
    .SEL(DLX_EXinst_Maddsub__n0016_inst_lut3_20),
    .O(DLX_EXinst_Maddsub__n0016_inst_cy_84)
  );
  X_XOR2 DLX_EXinst_Maddsub__n0016_inst_sum_84 (
    .I0(\DLX_EXinst__n0016<14>/CYINIT ),
    .I1(DLX_EXinst_Maddsub__n0016_inst_lut3_20),
    .O(\DLX_EXinst__n0016<14>/XORF )
  );
  defparam DLX_EXinst_Maddsub__n0016_inst_lut3_201.INIT = 16'h9966;
  X_LUT4 DLX_EXinst_Maddsub__n0016_inst_lut3_201 (
    .ADR0(DLX_IDinst_reg_out_A[14]),
    .ADR1(N108704),
    .ADR2(VCC),
    .ADR3(DLX_EXinst__n0017[14]),
    .O(DLX_EXinst_Maddsub__n0016_inst_lut3_20)
  );
  defparam DLX_EXinst_Maddsub__n0016_inst_lut3_211.INIT = 16'h9966;
  X_LUT4 DLX_EXinst_Maddsub__n0016_inst_lut3_211 (
    .ADR0(DLX_IDinst_reg_out_A[15]),
    .ADR1(DLX_EXinst__n0017[15]),
    .ADR2(VCC),
    .ADR3(N108704),
    .O(DLX_EXinst_Maddsub__n0016_inst_lut3_21)
  );
  X_BUF \DLX_EXinst__n0016<14>/COUTUSED  (
    .I(\DLX_EXinst__n0016<14>/CYMUXG ),
    .O(DLX_EXinst_Maddsub__n0016_inst_cy_85)
  );
  X_BUF \DLX_EXinst__n0016<14>/XUSED  (
    .I(\DLX_EXinst__n0016<14>/XORF ),
    .O(DLX_EXinst__n0016[14])
  );
  X_BUF \DLX_EXinst__n0016<14>/YUSED  (
    .I(\DLX_EXinst__n0016<14>/XORG ),
    .O(DLX_EXinst__n0016[15])
  );
  X_MUX2 DLX_EXinst_Maddsub__n0016_inst_cy_85_642 (
    .IA(DLX_IDinst_reg_out_A[15]),
    .IB(DLX_EXinst_Maddsub__n0016_inst_cy_84),
    .SEL(DLX_EXinst_Maddsub__n0016_inst_lut3_21),
    .O(\DLX_EXinst__n0016<14>/CYMUXG )
  );
  X_XOR2 DLX_EXinst_Maddsub__n0016_inst_sum_85 (
    .I0(DLX_EXinst_Maddsub__n0016_inst_cy_84),
    .I1(DLX_EXinst_Maddsub__n0016_inst_lut3_21),
    .O(\DLX_EXinst__n0016<14>/XORG )
  );
  X_BUF \DLX_EXinst__n0016<14>/CYINIT_643  (
    .I(DLX_EXinst_Maddsub__n0016_inst_cy_83),
    .O(\DLX_EXinst__n0016<14>/CYINIT )
  );
  X_MUX2 DLX_EXinst_Maddsub__n0016_inst_cy_86_644 (
    .IA(DLX_IDinst_reg_out_A[16]),
    .IB(\DLX_EXinst__n0016<16>/CYINIT ),
    .SEL(DLX_EXinst_Maddsub__n0016_inst_lut3_22),
    .O(DLX_EXinst_Maddsub__n0016_inst_cy_86)
  );
  X_XOR2 DLX_EXinst_Maddsub__n0016_inst_sum_86 (
    .I0(\DLX_EXinst__n0016<16>/CYINIT ),
    .I1(DLX_EXinst_Maddsub__n0016_inst_lut3_22),
    .O(\DLX_EXinst__n0016<16>/XORF )
  );
  defparam DLX_EXinst_Maddsub__n0016_inst_lut3_221.INIT = 16'hA55A;
  X_LUT4 DLX_EXinst_Maddsub__n0016_inst_lut3_221 (
    .ADR0(DLX_IDinst_reg_out_A[16]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst__n0017[16]),
    .ADR3(N108704),
    .O(DLX_EXinst_Maddsub__n0016_inst_lut3_22)
  );
  defparam DLX_EXinst_Maddsub__n0016_inst_lut3_231.INIT = 16'h9696;
  X_LUT4 DLX_EXinst_Maddsub__n0016_inst_lut3_231 (
    .ADR0(DLX_IDinst_reg_out_A[17]),
    .ADR1(DLX_EXinst__n0017[17]),
    .ADR2(N108704),
    .ADR3(VCC),
    .O(DLX_EXinst_Maddsub__n0016_inst_lut3_23)
  );
  X_BUF \DLX_EXinst__n0016<16>/COUTUSED  (
    .I(\DLX_EXinst__n0016<16>/CYMUXG ),
    .O(DLX_EXinst_Maddsub__n0016_inst_cy_87)
  );
  X_BUF \DLX_EXinst__n0016<16>/XUSED  (
    .I(\DLX_EXinst__n0016<16>/XORF ),
    .O(DLX_EXinst__n0016[16])
  );
  X_BUF \DLX_EXinst__n0016<16>/YUSED  (
    .I(\DLX_EXinst__n0016<16>/XORG ),
    .O(DLX_EXinst__n0016[17])
  );
  X_MUX2 DLX_EXinst_Maddsub__n0016_inst_cy_87_645 (
    .IA(DLX_IDinst_reg_out_A[17]),
    .IB(DLX_EXinst_Maddsub__n0016_inst_cy_86),
    .SEL(DLX_EXinst_Maddsub__n0016_inst_lut3_23),
    .O(\DLX_EXinst__n0016<16>/CYMUXG )
  );
  X_XOR2 DLX_EXinst_Maddsub__n0016_inst_sum_87 (
    .I0(DLX_EXinst_Maddsub__n0016_inst_cy_86),
    .I1(DLX_EXinst_Maddsub__n0016_inst_lut3_23),
    .O(\DLX_EXinst__n0016<16>/XORG )
  );
  X_BUF \DLX_EXinst__n0016<16>/CYINIT_646  (
    .I(DLX_EXinst_Maddsub__n0016_inst_cy_85),
    .O(\DLX_EXinst__n0016<16>/CYINIT )
  );
  X_MUX2 DLX_EXinst_Maddsub__n0016_inst_cy_88_647 (
    .IA(DLX_IDinst_reg_out_A[18]),
    .IB(\DLX_EXinst__n0016<18>/CYINIT ),
    .SEL(DLX_EXinst_Maddsub__n0016_inst_lut3_24),
    .O(DLX_EXinst_Maddsub__n0016_inst_cy_88)
  );
  X_XOR2 DLX_EXinst_Maddsub__n0016_inst_sum_88 (
    .I0(\DLX_EXinst__n0016<18>/CYINIT ),
    .I1(DLX_EXinst_Maddsub__n0016_inst_lut3_24),
    .O(\DLX_EXinst__n0016<18>/XORF )
  );
  defparam DLX_EXinst_Maddsub__n0016_inst_lut3_241.INIT = 16'h9966;
  X_LUT4 DLX_EXinst_Maddsub__n0016_inst_lut3_241 (
    .ADR0(DLX_IDinst_reg_out_A[18]),
    .ADR1(DLX_EXinst__n0017[18]),
    .ADR2(VCC),
    .ADR3(N108704),
    .O(DLX_EXinst_Maddsub__n0016_inst_lut3_24)
  );
  defparam DLX_EXinst_Maddsub__n0016_inst_lut3_251.INIT = 16'hA55A;
  X_LUT4 DLX_EXinst_Maddsub__n0016_inst_lut3_251 (
    .ADR0(DLX_IDinst_reg_out_A[19]),
    .ADR1(VCC),
    .ADR2(N108704),
    .ADR3(DLX_EXinst__n0017[19]),
    .O(DLX_EXinst_Maddsub__n0016_inst_lut3_25)
  );
  X_BUF \DLX_EXinst__n0016<18>/COUTUSED  (
    .I(\DLX_EXinst__n0016<18>/CYMUXG ),
    .O(DLX_EXinst_Maddsub__n0016_inst_cy_89)
  );
  X_BUF \DLX_EXinst__n0016<18>/XUSED  (
    .I(\DLX_EXinst__n0016<18>/XORF ),
    .O(DLX_EXinst__n0016[18])
  );
  X_BUF \DLX_EXinst__n0016<18>/YUSED  (
    .I(\DLX_EXinst__n0016<18>/XORG ),
    .O(DLX_EXinst__n0016[19])
  );
  X_MUX2 DLX_EXinst_Maddsub__n0016_inst_cy_89_648 (
    .IA(DLX_IDinst_reg_out_A[19]),
    .IB(DLX_EXinst_Maddsub__n0016_inst_cy_88),
    .SEL(DLX_EXinst_Maddsub__n0016_inst_lut3_25),
    .O(\DLX_EXinst__n0016<18>/CYMUXG )
  );
  X_XOR2 DLX_EXinst_Maddsub__n0016_inst_sum_89 (
    .I0(DLX_EXinst_Maddsub__n0016_inst_cy_88),
    .I1(DLX_EXinst_Maddsub__n0016_inst_lut3_25),
    .O(\DLX_EXinst__n0016<18>/XORG )
  );
  X_BUF \DLX_EXinst__n0016<18>/CYINIT_649  (
    .I(DLX_EXinst_Maddsub__n0016_inst_cy_87),
    .O(\DLX_EXinst__n0016<18>/CYINIT )
  );
  X_MUX2 DLX_EXinst_Maddsub__n0016_inst_cy_90_650 (
    .IA(DLX_IDinst_reg_out_A[20]),
    .IB(\DLX_EXinst__n0016<20>/CYINIT ),
    .SEL(DLX_EXinst_Maddsub__n0016_inst_lut3_26),
    .O(DLX_EXinst_Maddsub__n0016_inst_cy_90)
  );
  X_XOR2 DLX_EXinst_Maddsub__n0016_inst_sum_90 (
    .I0(\DLX_EXinst__n0016<20>/CYINIT ),
    .I1(DLX_EXinst_Maddsub__n0016_inst_lut3_26),
    .O(\DLX_EXinst__n0016<20>/XORF )
  );
  defparam DLX_EXinst_Maddsub__n0016_inst_lut3_261.INIT = 16'h9696;
  X_LUT4 DLX_EXinst_Maddsub__n0016_inst_lut3_261 (
    .ADR0(DLX_IDinst_reg_out_A[20]),
    .ADR1(N108704),
    .ADR2(DLX_EXinst__n0017[20]),
    .ADR3(VCC),
    .O(DLX_EXinst_Maddsub__n0016_inst_lut3_26)
  );
  defparam DLX_EXinst_Maddsub__n0016_inst_lut3_271.INIT = 16'h9966;
  X_LUT4 DLX_EXinst_Maddsub__n0016_inst_lut3_271 (
    .ADR0(DLX_IDinst_reg_out_A[21]),
    .ADR1(DLX_EXinst__n0017[21]),
    .ADR2(VCC),
    .ADR3(N108704),
    .O(DLX_EXinst_Maddsub__n0016_inst_lut3_27)
  );
  X_BUF \DLX_EXinst__n0016<20>/COUTUSED  (
    .I(\DLX_EXinst__n0016<20>/CYMUXG ),
    .O(DLX_EXinst_Maddsub__n0016_inst_cy_91)
  );
  X_BUF \DLX_EXinst__n0016<20>/XUSED  (
    .I(\DLX_EXinst__n0016<20>/XORF ),
    .O(DLX_EXinst__n0016[20])
  );
  X_BUF \DLX_EXinst__n0016<20>/YUSED  (
    .I(\DLX_EXinst__n0016<20>/XORG ),
    .O(DLX_EXinst__n0016[21])
  );
  X_MUX2 DLX_EXinst_Maddsub__n0016_inst_cy_91_651 (
    .IA(DLX_IDinst_reg_out_A[21]),
    .IB(DLX_EXinst_Maddsub__n0016_inst_cy_90),
    .SEL(DLX_EXinst_Maddsub__n0016_inst_lut3_27),
    .O(\DLX_EXinst__n0016<20>/CYMUXG )
  );
  X_XOR2 DLX_EXinst_Maddsub__n0016_inst_sum_91 (
    .I0(DLX_EXinst_Maddsub__n0016_inst_cy_90),
    .I1(DLX_EXinst_Maddsub__n0016_inst_lut3_27),
    .O(\DLX_EXinst__n0016<20>/XORG )
  );
  X_BUF \DLX_EXinst__n0016<20>/CYINIT_652  (
    .I(DLX_EXinst_Maddsub__n0016_inst_cy_89),
    .O(\DLX_EXinst__n0016<20>/CYINIT )
  );
  X_MUX2 DLX_EXinst_Maddsub__n0016_inst_cy_92_653 (
    .IA(DLX_IDinst_reg_out_A[22]),
    .IB(\DLX_EXinst__n0016<22>/CYINIT ),
    .SEL(DLX_EXinst_Maddsub__n0016_inst_lut3_28),
    .O(DLX_EXinst_Maddsub__n0016_inst_cy_92)
  );
  X_XOR2 DLX_EXinst_Maddsub__n0016_inst_sum_92 (
    .I0(\DLX_EXinst__n0016<22>/CYINIT ),
    .I1(DLX_EXinst_Maddsub__n0016_inst_lut3_28),
    .O(\DLX_EXinst__n0016<22>/XORF )
  );
  defparam DLX_EXinst_Maddsub__n0016_inst_lut3_281.INIT = 16'h9696;
  X_LUT4 DLX_EXinst_Maddsub__n0016_inst_lut3_281 (
    .ADR0(DLX_IDinst_reg_out_A[22]),
    .ADR1(N108704),
    .ADR2(DLX_EXinst__n0017[22]),
    .ADR3(VCC),
    .O(DLX_EXinst_Maddsub__n0016_inst_lut3_28)
  );
  defparam DLX_EXinst_Maddsub__n0016_inst_lut3_291.INIT = 16'h9696;
  X_LUT4 DLX_EXinst_Maddsub__n0016_inst_lut3_291 (
    .ADR0(DLX_IDinst_reg_out_A[23]),
    .ADR1(N108704),
    .ADR2(DLX_EXinst__n0017[23]),
    .ADR3(VCC),
    .O(DLX_EXinst_Maddsub__n0016_inst_lut3_29)
  );
  X_BUF \DLX_EXinst__n0016<22>/COUTUSED  (
    .I(\DLX_EXinst__n0016<22>/CYMUXG ),
    .O(DLX_EXinst_Maddsub__n0016_inst_cy_93)
  );
  X_BUF \DLX_EXinst__n0016<22>/XUSED  (
    .I(\DLX_EXinst__n0016<22>/XORF ),
    .O(DLX_EXinst__n0016[22])
  );
  X_BUF \DLX_EXinst__n0016<22>/YUSED  (
    .I(\DLX_EXinst__n0016<22>/XORG ),
    .O(DLX_EXinst__n0016[23])
  );
  X_MUX2 DLX_EXinst_Maddsub__n0016_inst_cy_93_654 (
    .IA(DLX_IDinst_reg_out_A[23]),
    .IB(DLX_EXinst_Maddsub__n0016_inst_cy_92),
    .SEL(DLX_EXinst_Maddsub__n0016_inst_lut3_29),
    .O(\DLX_EXinst__n0016<22>/CYMUXG )
  );
  X_XOR2 DLX_EXinst_Maddsub__n0016_inst_sum_93 (
    .I0(DLX_EXinst_Maddsub__n0016_inst_cy_92),
    .I1(DLX_EXinst_Maddsub__n0016_inst_lut3_29),
    .O(\DLX_EXinst__n0016<22>/XORG )
  );
  X_BUF \DLX_EXinst__n0016<22>/CYINIT_655  (
    .I(DLX_EXinst_Maddsub__n0016_inst_cy_91),
    .O(\DLX_EXinst__n0016<22>/CYINIT )
  );
  X_MUX2 DLX_EXinst_Maddsub__n0016_inst_cy_94_656 (
    .IA(DLX_IDinst_reg_out_A[24]),
    .IB(\DLX_EXinst__n0016<24>/CYINIT ),
    .SEL(DLX_EXinst_Maddsub__n0016_inst_lut3_30),
    .O(DLX_EXinst_Maddsub__n0016_inst_cy_94)
  );
  X_XOR2 DLX_EXinst_Maddsub__n0016_inst_sum_94 (
    .I0(\DLX_EXinst__n0016<24>/CYINIT ),
    .I1(DLX_EXinst_Maddsub__n0016_inst_lut3_30),
    .O(\DLX_EXinst__n0016<24>/XORF )
  );
  defparam DLX_EXinst_Maddsub__n0016_inst_lut3_301.INIT = 16'h9696;
  X_LUT4 DLX_EXinst_Maddsub__n0016_inst_lut3_301 (
    .ADR0(DLX_IDinst_reg_out_A[24]),
    .ADR1(N108704),
    .ADR2(DLX_EXinst__n0017[24]),
    .ADR3(VCC),
    .O(DLX_EXinst_Maddsub__n0016_inst_lut3_30)
  );
  defparam DLX_EXinst_Maddsub__n0016_inst_lut3_311.INIT = 16'h9966;
  X_LUT4 DLX_EXinst_Maddsub__n0016_inst_lut3_311 (
    .ADR0(DLX_IDinst_reg_out_A[25]),
    .ADR1(N108704),
    .ADR2(VCC),
    .ADR3(DLX_EXinst__n0017[25]),
    .O(DLX_EXinst_Maddsub__n0016_inst_lut3_31)
  );
  X_BUF \DLX_EXinst__n0016<24>/COUTUSED  (
    .I(\DLX_EXinst__n0016<24>/CYMUXG ),
    .O(DLX_EXinst_Maddsub__n0016_inst_cy_95)
  );
  X_BUF \DLX_EXinst__n0016<24>/XUSED  (
    .I(\DLX_EXinst__n0016<24>/XORF ),
    .O(DLX_EXinst__n0016[24])
  );
  X_BUF \DLX_EXinst__n0016<24>/YUSED  (
    .I(\DLX_EXinst__n0016<24>/XORG ),
    .O(DLX_EXinst__n0016[25])
  );
  X_MUX2 DLX_EXinst_Maddsub__n0016_inst_cy_95_657 (
    .IA(DLX_IDinst_reg_out_A[25]),
    .IB(DLX_EXinst_Maddsub__n0016_inst_cy_94),
    .SEL(DLX_EXinst_Maddsub__n0016_inst_lut3_31),
    .O(\DLX_EXinst__n0016<24>/CYMUXG )
  );
  X_XOR2 DLX_EXinst_Maddsub__n0016_inst_sum_95 (
    .I0(DLX_EXinst_Maddsub__n0016_inst_cy_94),
    .I1(DLX_EXinst_Maddsub__n0016_inst_lut3_31),
    .O(\DLX_EXinst__n0016<24>/XORG )
  );
  X_BUF \DLX_EXinst__n0016<24>/CYINIT_658  (
    .I(DLX_EXinst_Maddsub__n0016_inst_cy_93),
    .O(\DLX_EXinst__n0016<24>/CYINIT )
  );
  X_MUX2 DLX_EXinst_Maddsub__n0016_inst_cy_96_659 (
    .IA(DLX_IDinst_reg_out_A[26]),
    .IB(\DLX_EXinst__n0016<26>/CYINIT ),
    .SEL(DLX_EXinst_Maddsub__n0016_inst_lut3_32),
    .O(DLX_EXinst_Maddsub__n0016_inst_cy_96)
  );
  X_XOR2 DLX_EXinst_Maddsub__n0016_inst_sum_96 (
    .I0(\DLX_EXinst__n0016<26>/CYINIT ),
    .I1(DLX_EXinst_Maddsub__n0016_inst_lut3_32),
    .O(\DLX_EXinst__n0016<26>/XORF )
  );
  defparam DLX_EXinst_Maddsub__n0016_inst_lut3_321.INIT = 16'h9696;
  X_LUT4 DLX_EXinst_Maddsub__n0016_inst_lut3_321 (
    .ADR0(DLX_IDinst_reg_out_A[26]),
    .ADR1(DLX_EXinst__n0017[26]),
    .ADR2(N108704),
    .ADR3(VCC),
    .O(DLX_EXinst_Maddsub__n0016_inst_lut3_32)
  );
  defparam DLX_EXinst_Maddsub__n0016_inst_lut3_331.INIT = 16'h9966;
  X_LUT4 DLX_EXinst_Maddsub__n0016_inst_lut3_331 (
    .ADR0(DLX_IDinst_reg_out_A[27]),
    .ADR1(N108704),
    .ADR2(VCC),
    .ADR3(DLX_EXinst__n0017[27]),
    .O(DLX_EXinst_Maddsub__n0016_inst_lut3_33)
  );
  X_BUF \DLX_EXinst__n0016<26>/COUTUSED  (
    .I(\DLX_EXinst__n0016<26>/CYMUXG ),
    .O(DLX_EXinst_Maddsub__n0016_inst_cy_97)
  );
  X_BUF \DLX_EXinst__n0016<26>/XUSED  (
    .I(\DLX_EXinst__n0016<26>/XORF ),
    .O(DLX_EXinst__n0016[26])
  );
  X_BUF \DLX_EXinst__n0016<26>/YUSED  (
    .I(\DLX_EXinst__n0016<26>/XORG ),
    .O(DLX_EXinst__n0016[27])
  );
  X_MUX2 DLX_EXinst_Maddsub__n0016_inst_cy_97_660 (
    .IA(DLX_IDinst_reg_out_A[27]),
    .IB(DLX_EXinst_Maddsub__n0016_inst_cy_96),
    .SEL(DLX_EXinst_Maddsub__n0016_inst_lut3_33),
    .O(\DLX_EXinst__n0016<26>/CYMUXG )
  );
  X_XOR2 DLX_EXinst_Maddsub__n0016_inst_sum_97 (
    .I0(DLX_EXinst_Maddsub__n0016_inst_cy_96),
    .I1(DLX_EXinst_Maddsub__n0016_inst_lut3_33),
    .O(\DLX_EXinst__n0016<26>/XORG )
  );
  X_BUF \DLX_EXinst__n0016<26>/CYINIT_661  (
    .I(DLX_EXinst_Maddsub__n0016_inst_cy_95),
    .O(\DLX_EXinst__n0016<26>/CYINIT )
  );
  X_MUX2 DLX_EXinst_Maddsub__n0016_inst_cy_98_662 (
    .IA(DLX_IDinst_reg_out_A[28]),
    .IB(\DLX_EXinst__n0016<28>/CYINIT ),
    .SEL(DLX_EXinst_Maddsub__n0016_inst_lut3_34),
    .O(DLX_EXinst_Maddsub__n0016_inst_cy_98)
  );
  X_XOR2 DLX_EXinst_Maddsub__n0016_inst_sum_98 (
    .I0(\DLX_EXinst__n0016<28>/CYINIT ),
    .I1(DLX_EXinst_Maddsub__n0016_inst_lut3_34),
    .O(\DLX_EXinst__n0016<28>/XORF )
  );
  defparam DLX_EXinst_Maddsub__n0016_inst_lut3_341.INIT = 16'h9696;
  X_LUT4 DLX_EXinst_Maddsub__n0016_inst_lut3_341 (
    .ADR0(DLX_IDinst_reg_out_A[28]),
    .ADR1(N108704),
    .ADR2(DLX_EXinst__n0017[28]),
    .ADR3(VCC),
    .O(DLX_EXinst_Maddsub__n0016_inst_lut3_34)
  );
  defparam DLX_EXinst_Maddsub__n0016_inst_lut3_351.INIT = 16'h9966;
  X_LUT4 DLX_EXinst_Maddsub__n0016_inst_lut3_351 (
    .ADR0(DLX_IDinst_reg_out_A[29]),
    .ADR1(N108704),
    .ADR2(VCC),
    .ADR3(DLX_EXinst__n0017[29]),
    .O(DLX_EXinst_Maddsub__n0016_inst_lut3_35)
  );
  X_BUF \DLX_EXinst__n0016<28>/COUTUSED  (
    .I(\DLX_EXinst__n0016<28>/CYMUXG ),
    .O(DLX_EXinst_Maddsub__n0016_inst_cy_99)
  );
  X_BUF \DLX_EXinst__n0016<28>/XUSED  (
    .I(\DLX_EXinst__n0016<28>/XORF ),
    .O(DLX_EXinst__n0016[28])
  );
  X_BUF \DLX_EXinst__n0016<28>/YUSED  (
    .I(\DLX_EXinst__n0016<28>/XORG ),
    .O(DLX_EXinst__n0016[29])
  );
  X_MUX2 DLX_EXinst_Maddsub__n0016_inst_cy_99_663 (
    .IA(DLX_IDinst_reg_out_A[29]),
    .IB(DLX_EXinst_Maddsub__n0016_inst_cy_98),
    .SEL(DLX_EXinst_Maddsub__n0016_inst_lut3_35),
    .O(\DLX_EXinst__n0016<28>/CYMUXG )
  );
  X_XOR2 DLX_EXinst_Maddsub__n0016_inst_sum_99 (
    .I0(DLX_EXinst_Maddsub__n0016_inst_cy_98),
    .I1(DLX_EXinst_Maddsub__n0016_inst_lut3_35),
    .O(\DLX_EXinst__n0016<28>/XORG )
  );
  X_BUF \DLX_EXinst__n0016<28>/CYINIT_664  (
    .I(DLX_EXinst_Maddsub__n0016_inst_cy_97),
    .O(\DLX_EXinst__n0016<28>/CYINIT )
  );
  X_MUX2 DLX_EXinst_Maddsub__n0016_inst_cy_100_665 (
    .IA(DLX_IDinst_reg_out_A[30]),
    .IB(\DLX_EXinst__n0016<30>/CYINIT ),
    .SEL(DLX_EXinst_Maddsub__n0016_inst_lut3_36),
    .O(DLX_EXinst_Maddsub__n0016_inst_cy_100)
  );
  X_XOR2 DLX_EXinst_Maddsub__n0016_inst_sum_100 (
    .I0(\DLX_EXinst__n0016<30>/CYINIT ),
    .I1(DLX_EXinst_Maddsub__n0016_inst_lut3_36),
    .O(\DLX_EXinst__n0016<30>/XORF )
  );
  defparam DLX_EXinst_Maddsub__n0016_inst_lut3_361.INIT = 16'h9696;
  X_LUT4 DLX_EXinst_Maddsub__n0016_inst_lut3_361 (
    .ADR0(DLX_IDinst_reg_out_A[30]),
    .ADR1(N108704),
    .ADR2(DLX_EXinst__n0017[30]),
    .ADR3(VCC),
    .O(DLX_EXinst_Maddsub__n0016_inst_lut3_36)
  );
  defparam DLX_EXinst_Maddsub__n0016_inst_lut3_371.INIT = 16'hA55A;
  X_LUT4 DLX_EXinst_Maddsub__n0016_inst_lut3_371 (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst__n0017[31]),
    .ADR3(N108704),
    .O(DLX_EXinst_Maddsub__n0016_inst_lut3_37)
  );
  X_BUF \DLX_EXinst__n0016<30>/XUSED  (
    .I(\DLX_EXinst__n0016<30>/XORF ),
    .O(DLX_EXinst__n0016[30])
  );
  X_BUF \DLX_EXinst__n0016<30>/YUSED  (
    .I(\DLX_EXinst__n0016<30>/XORG ),
    .O(DLX_EXinst__n0016[31])
  );
  X_XOR2 DLX_EXinst_Maddsub__n0016_inst_sum_101 (
    .I0(DLX_EXinst_Maddsub__n0016_inst_cy_100),
    .I1(DLX_EXinst_Maddsub__n0016_inst_lut3_37),
    .O(\DLX_EXinst__n0016<30>/XORG )
  );
  X_BUF \DLX_EXinst__n0016<30>/CYINIT_666  (
    .I(DLX_EXinst_Maddsub__n0016_inst_cy_99),
    .O(\DLX_EXinst__n0016<30>/CYINIT )
  );
  X_ONE \DLX_IDinst_Mcompar__n0078_inst_cy_263/LOGIC_ONE_667  (
    .O(\DLX_IDinst_Mcompar__n0078_inst_cy_263/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mcompar__n0078_inst_cy_263/LOGIC_ZERO_668  (
    .O(\DLX_IDinst_Mcompar__n0078_inst_cy_263/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mcompar__n0078_inst_cy_262_669 (
    .IA(\DLX_IDinst_Mcompar__n0078_inst_cy_263/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mcompar__n0078_inst_cy_263/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mcompar__n0078_inst_lut4_40),
    .O(DLX_IDinst_Mcompar__n0078_inst_cy_262)
  );
  defparam DLX_IDinst_Mcompar__n0078_inst_lut4_401.INIT = 16'h8421;
  X_LUT4 DLX_IDinst_Mcompar__n0078_inst_lut4_401 (
    .ADR0(DLX_reg_dst_of_MEM[0]),
    .ADR1(DLX_IDinst_regB_index[1]),
    .ADR2(DLX_IDinst_regB_index[0]),
    .ADR3(DLX_reg_dst_of_MEM[1]),
    .O(DLX_IDinst_Mcompar__n0078_inst_lut4_40)
  );
  defparam DLX_IDinst_Mcompar__n0078_inst_lut4_411.INIT = 16'h9009;
  X_LUT4 DLX_IDinst_Mcompar__n0078_inst_lut4_411 (
    .ADR0(DLX_IDinst_regB_index[2]),
    .ADR1(DLX_reg_dst_of_MEM[2]),
    .ADR2(DLX_reg_dst_of_MEM[3]),
    .ADR3(DLX_IDinst_regB_index[3]),
    .O(DLX_IDinst_Mcompar__n0078_inst_lut4_41)
  );
  X_BUF \DLX_IDinst_Mcompar__n0078_inst_cy_263/COUTUSED  (
    .I(\DLX_IDinst_Mcompar__n0078_inst_cy_263/CYMUXG ),
    .O(DLX_IDinst_Mcompar__n0078_inst_cy_263)
  );
  X_MUX2 DLX_IDinst_Mcompar__n0078_inst_cy_263_670 (
    .IA(\DLX_IDinst_Mcompar__n0078_inst_cy_263/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mcompar__n0078_inst_cy_262),
    .SEL(DLX_IDinst_Mcompar__n0078_inst_lut4_41),
    .O(\DLX_IDinst_Mcompar__n0078_inst_cy_263/CYMUXG )
  );
  X_ZERO \DLX_IDinst__n0078/LOGIC_ZERO_671  (
    .O(\DLX_IDinst__n0078/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mcompar__n0078_inst_cy_264 (
    .IA(\DLX_IDinst__n0078/LOGIC_ZERO ),
    .IB(\DLX_IDinst__n0078/CYINIT ),
    .SEL(DLX_IDinst_Mcompar__n0078_inst_lut4_42),
    .O(\DLX_IDinst__n0078/CYMUXF )
  );
  defparam DLX_IDinst_Mcompar__n0078_inst_lut4_421.INIT = 16'hAA55;
  X_LUT4 DLX_IDinst_Mcompar__n0078_inst_lut4_421 (
    .ADR0(DLX_reg_dst_of_MEM[4]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_regB_index[4]),
    .O(DLX_IDinst_Mcompar__n0078_inst_lut4_42)
  );
  X_BUF \DLX_IDinst__n0078/XBUSED  (
    .I(\DLX_IDinst__n0078/CYMUXF ),
    .O(DLX_IDinst__n0078)
  );
  X_BUF \DLX_IDinst__n0078/CYINIT_672  (
    .I(DLX_IDinst_Mcompar__n0078_inst_cy_263),
    .O(\DLX_IDinst__n0078/CYINIT )
  );
  defparam DLX_IFinst_NPC_9_1_673.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_9_1_673 (
    .I(\NPC_eff<9>/OD ),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\NPC_eff<9>/OFF/RST ),
    .O(DLX_IFinst_NPC_9_1)
  );
  X_OR2 \NPC_eff<9>/OFF/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\NPC_eff<9>/OFF/RST )
  );
  X_ZERO \DLX_EXinst_Mcompar__n0087_inst_cy_119/LOGIC_ZERO_674  (
    .O(\DLX_EXinst_Mcompar__n0087_inst_cy_119/LOGIC_ZERO )
  );
  X_ONE \DLX_EXinst_Mcompar__n0087_inst_cy_119/LOGIC_ONE_675  (
    .O(\DLX_EXinst_Mcompar__n0087_inst_cy_119/LOGIC_ONE )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0087_inst_cy_118_676 (
    .IA(\DLX_EXinst_Mcompar__n0087_inst_cy_119/LOGIC_ONE ),
    .IB(\DLX_EXinst_Mcompar__n0087_inst_cy_119/LOGIC_ZERO ),
    .SEL(DLX_EXinst_Mcompar__n0087_inst_lut4_16),
    .O(DLX_EXinst_Mcompar__n0087_inst_cy_118)
  );
  defparam DLX_EXinst_Mcompar__n0087_inst_lut4_161.INIT = 16'h8241;
  X_LUT4 DLX_EXinst_Mcompar__n0087_inst_lut4_161 (
    .ADR0(DLX_IDinst_IR_function_field_1_1),
    .ADR1(DLX_IDinst_reg_out_A[0]),
    .ADR2(DLX_IDinst_IR_function_field_0_1),
    .ADR3(DLX_IDinst_reg_out_A[1]),
    .O(DLX_EXinst_Mcompar__n0087_inst_lut4_16)
  );
  defparam DLX_EXinst_Mcompar__n0087_inst_lut4_171.INIT = 16'h8421;
  X_LUT4 DLX_EXinst_Mcompar__n0087_inst_lut4_171 (
    .ADR0(DLX_IDinst_IR_function_field_2_1),
    .ADR1(DLX_IDinst_IR_function_field_3_1),
    .ADR2(DLX_IDinst_reg_out_A[2]),
    .ADR3(DLX_IDinst_reg_out_A[3]),
    .O(DLX_EXinst_Mcompar__n0087_inst_lut4_17)
  );
  X_BUF \DLX_EXinst_Mcompar__n0087_inst_cy_119/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0087_inst_cy_119/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0087_inst_cy_119)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0087_inst_cy_119_677 (
    .IA(\DLX_EXinst_Mcompar__n0087_inst_cy_119/LOGIC_ONE ),
    .IB(DLX_EXinst_Mcompar__n0087_inst_cy_118),
    .SEL(DLX_EXinst_Mcompar__n0087_inst_lut4_17),
    .O(\DLX_EXinst_Mcompar__n0087_inst_cy_119/CYMUXG )
  );
  X_ONE \DLX_EXinst_Mcompar__n0087_inst_cy_121/LOGIC_ONE_678  (
    .O(\DLX_EXinst_Mcompar__n0087_inst_cy_121/LOGIC_ONE )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0087_inst_cy_120_679 (
    .IA(\DLX_EXinst_Mcompar__n0087_inst_cy_121/LOGIC_ONE ),
    .IB(\DLX_EXinst_Mcompar__n0087_inst_cy_121/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0087_inst_lut4_18),
    .O(DLX_EXinst_Mcompar__n0087_inst_cy_120)
  );
  defparam DLX_EXinst_Mcompar__n0087_inst_lut4_181.INIT = 16'h8421;
  X_LUT4 DLX_EXinst_Mcompar__n0087_inst_lut4_181 (
    .ADR0(DLX_IDinst_reg_out_A[5]),
    .ADR1(DLX_IDinst_reg_out_A[4]),
    .ADR2(\DLX_IDinst_Imm[5] ),
    .ADR3(DLX_IDinst_IR_function_field[4]),
    .O(DLX_EXinst_Mcompar__n0087_inst_lut4_18)
  );
  defparam DLX_EXinst_Mcompar__n0087_inst_lut4_191.INIT = 16'h8241;
  X_LUT4 DLX_EXinst_Mcompar__n0087_inst_lut4_191 (
    .ADR0(DLX_IDinst_reg_out_A[7]),
    .ADR1(\DLX_IDinst_Imm[6] ),
    .ADR2(DLX_IDinst_reg_out_A[6]),
    .ADR3(\DLX_IDinst_Imm[7] ),
    .O(DLX_EXinst_Mcompar__n0087_inst_lut4_19)
  );
  X_BUF \DLX_EXinst_Mcompar__n0087_inst_cy_121/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0087_inst_cy_121/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0087_inst_cy_121)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0087_inst_cy_121_680 (
    .IA(\DLX_EXinst_Mcompar__n0087_inst_cy_121/LOGIC_ONE ),
    .IB(DLX_EXinst_Mcompar__n0087_inst_cy_120),
    .SEL(DLX_EXinst_Mcompar__n0087_inst_lut4_19),
    .O(\DLX_EXinst_Mcompar__n0087_inst_cy_121/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0087_inst_cy_121/CYINIT_681  (
    .I(DLX_EXinst_Mcompar__n0087_inst_cy_119),
    .O(\DLX_EXinst_Mcompar__n0087_inst_cy_121/CYINIT )
  );
  X_ONE \DLX_EXinst_Mcompar__n0087_inst_cy_123/LOGIC_ONE_682  (
    .O(\DLX_EXinst_Mcompar__n0087_inst_cy_123/LOGIC_ONE )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0087_inst_cy_122_683 (
    .IA(\DLX_EXinst_Mcompar__n0087_inst_cy_123/LOGIC_ONE ),
    .IB(\DLX_EXinst_Mcompar__n0087_inst_cy_123/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0087_inst_lut4_20),
    .O(DLX_EXinst_Mcompar__n0087_inst_cy_122)
  );
  defparam DLX_EXinst_Mcompar__n0087_inst_lut4_201.INIT = 16'h8241;
  X_LUT4 DLX_EXinst_Mcompar__n0087_inst_lut4_201 (
    .ADR0(DLX_IDinst_reg_out_A[8]),
    .ADR1(DLX_IDinst_reg_out_A[9]),
    .ADR2(\DLX_IDinst_Imm[9] ),
    .ADR3(\DLX_IDinst_Imm[8] ),
    .O(DLX_EXinst_Mcompar__n0087_inst_lut4_20)
  );
  defparam DLX_EXinst_Mcompar__n0087_inst_lut4_211.INIT = 16'h8421;
  X_LUT4 DLX_EXinst_Mcompar__n0087_inst_lut4_211 (
    .ADR0(\DLX_IDinst_Imm[11] ),
    .ADR1(\DLX_IDinst_Imm[10] ),
    .ADR2(DLX_IDinst_reg_out_A[11]),
    .ADR3(DLX_IDinst_reg_out_A[10]),
    .O(DLX_EXinst_Mcompar__n0087_inst_lut4_21)
  );
  X_BUF \DLX_EXinst_Mcompar__n0087_inst_cy_123/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0087_inst_cy_123/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0087_inst_cy_123)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0087_inst_cy_123_684 (
    .IA(\DLX_EXinst_Mcompar__n0087_inst_cy_123/LOGIC_ONE ),
    .IB(DLX_EXinst_Mcompar__n0087_inst_cy_122),
    .SEL(DLX_EXinst_Mcompar__n0087_inst_lut4_21),
    .O(\DLX_EXinst_Mcompar__n0087_inst_cy_123/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0087_inst_cy_123/CYINIT_685  (
    .I(DLX_EXinst_Mcompar__n0087_inst_cy_121),
    .O(\DLX_EXinst_Mcompar__n0087_inst_cy_123/CYINIT )
  );
  X_ONE \DLX_EXinst_Mcompar__n0087_inst_cy_125/LOGIC_ONE_686  (
    .O(\DLX_EXinst_Mcompar__n0087_inst_cy_125/LOGIC_ONE )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0087_inst_cy_124_687 (
    .IA(\DLX_EXinst_Mcompar__n0087_inst_cy_125/LOGIC_ONE ),
    .IB(\DLX_EXinst_Mcompar__n0087_inst_cy_125/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0087_inst_lut4_22),
    .O(DLX_EXinst_Mcompar__n0087_inst_cy_124)
  );
  defparam DLX_EXinst_Mcompar__n0087_inst_lut4_221.INIT = 16'h8241;
  X_LUT4 DLX_EXinst_Mcompar__n0087_inst_lut4_221 (
    .ADR0(\DLX_IDinst_Imm[13] ),
    .ADR1(DLX_IDinst_reg_out_A[12]),
    .ADR2(\DLX_IDinst_Imm[12] ),
    .ADR3(DLX_IDinst_reg_out_A[13]),
    .O(DLX_EXinst_Mcompar__n0087_inst_lut4_22)
  );
  defparam DLX_EXinst_Mcompar__n0087_inst_lut4_231.INIT = 16'h8421;
  X_LUT4 DLX_EXinst_Mcompar__n0087_inst_lut4_231 (
    .ADR0(\DLX_IDinst_Imm[15] ),
    .ADR1(\DLX_IDinst_Imm[14] ),
    .ADR2(DLX_IDinst_reg_out_A[15]),
    .ADR3(DLX_IDinst_reg_out_A[14]),
    .O(DLX_EXinst_Mcompar__n0087_inst_lut4_23)
  );
  X_BUF \DLX_EXinst_Mcompar__n0087_inst_cy_125/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0087_inst_cy_125/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0087_inst_cy_125)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0087_inst_cy_125_688 (
    .IA(\DLX_EXinst_Mcompar__n0087_inst_cy_125/LOGIC_ONE ),
    .IB(DLX_EXinst_Mcompar__n0087_inst_cy_124),
    .SEL(DLX_EXinst_Mcompar__n0087_inst_lut4_23),
    .O(\DLX_EXinst_Mcompar__n0087_inst_cy_125/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0087_inst_cy_125/CYINIT_689  (
    .I(DLX_EXinst_Mcompar__n0087_inst_cy_123),
    .O(\DLX_EXinst_Mcompar__n0087_inst_cy_125/CYINIT )
  );
  X_ONE \DLX_EXinst_Mcompar__n0087_inst_cy_127/LOGIC_ONE_690  (
    .O(\DLX_EXinst_Mcompar__n0087_inst_cy_127/LOGIC_ONE )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0087_inst_cy_126_691 (
    .IA(\DLX_EXinst_Mcompar__n0087_inst_cy_127/LOGIC_ONE ),
    .IB(\DLX_EXinst_Mcompar__n0087_inst_cy_127/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0087_inst_lut4_24),
    .O(DLX_EXinst_Mcompar__n0087_inst_cy_126)
  );
  defparam DLX_EXinst_Mcompar__n0087_inst_lut4_241.INIT = 16'h8811;
  X_LUT4 DLX_EXinst_Mcompar__n0087_inst_lut4_241 (
    .ADR0(DLX_IDinst_reg_out_A[16]),
    .ADR1(DLX_IDinst_reg_out_A[17]),
    .ADR2(VCC),
    .ADR3(\DLX_IDinst_Imm[31] ),
    .O(DLX_EXinst_Mcompar__n0087_inst_lut4_24)
  );
  defparam DLX_EXinst_Mcompar__n0087_inst_lut4_251.INIT = 16'h8811;
  X_LUT4 DLX_EXinst_Mcompar__n0087_inst_lut4_251 (
    .ADR0(DLX_IDinst_reg_out_A[19]),
    .ADR1(DLX_IDinst_reg_out_A[18]),
    .ADR2(VCC),
    .ADR3(\DLX_IDinst_Imm[31] ),
    .O(DLX_EXinst_Mcompar__n0087_inst_lut4_25)
  );
  X_BUF \DLX_EXinst_Mcompar__n0087_inst_cy_127/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0087_inst_cy_127/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0087_inst_cy_127)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0087_inst_cy_127_692 (
    .IA(\DLX_EXinst_Mcompar__n0087_inst_cy_127/LOGIC_ONE ),
    .IB(DLX_EXinst_Mcompar__n0087_inst_cy_126),
    .SEL(DLX_EXinst_Mcompar__n0087_inst_lut4_25),
    .O(\DLX_EXinst_Mcompar__n0087_inst_cy_127/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0087_inst_cy_127/CYINIT_693  (
    .I(DLX_EXinst_Mcompar__n0087_inst_cy_125),
    .O(\DLX_EXinst_Mcompar__n0087_inst_cy_127/CYINIT )
  );
  X_ONE \DLX_EXinst_Mcompar__n0087_inst_cy_129/LOGIC_ONE_694  (
    .O(\DLX_EXinst_Mcompar__n0087_inst_cy_129/LOGIC_ONE )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0087_inst_cy_128_695 (
    .IA(\DLX_EXinst_Mcompar__n0087_inst_cy_129/LOGIC_ONE ),
    .IB(\DLX_EXinst_Mcompar__n0087_inst_cy_129/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0087_inst_lut4_26),
    .O(DLX_EXinst_Mcompar__n0087_inst_cy_128)
  );
  defparam DLX_EXinst_Mcompar__n0087_inst_lut4_261.INIT = 16'hC003;
  X_LUT4 DLX_EXinst_Mcompar__n0087_inst_lut4_261 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[20]),
    .ADR2(\DLX_IDinst_Imm[31] ),
    .ADR3(DLX_IDinst_reg_out_A[21]),
    .O(DLX_EXinst_Mcompar__n0087_inst_lut4_26)
  );
  defparam DLX_EXinst_Mcompar__n0087_inst_lut4_271.INIT = 16'hC003;
  X_LUT4 DLX_EXinst_Mcompar__n0087_inst_lut4_271 (
    .ADR0(VCC),
    .ADR1(\DLX_IDinst_Imm[31] ),
    .ADR2(DLX_IDinst_reg_out_A[22]),
    .ADR3(DLX_IDinst_reg_out_A[23]),
    .O(DLX_EXinst_Mcompar__n0087_inst_lut4_27)
  );
  X_BUF \DLX_EXinst_Mcompar__n0087_inst_cy_129/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0087_inst_cy_129/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0087_inst_cy_129)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0087_inst_cy_129_696 (
    .IA(\DLX_EXinst_Mcompar__n0087_inst_cy_129/LOGIC_ONE ),
    .IB(DLX_EXinst_Mcompar__n0087_inst_cy_128),
    .SEL(DLX_EXinst_Mcompar__n0087_inst_lut4_27),
    .O(\DLX_EXinst_Mcompar__n0087_inst_cy_129/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0087_inst_cy_129/CYINIT_697  (
    .I(DLX_EXinst_Mcompar__n0087_inst_cy_127),
    .O(\DLX_EXinst_Mcompar__n0087_inst_cy_129/CYINIT )
  );
  X_ONE \DLX_EXinst_Mcompar__n0087_inst_cy_131/LOGIC_ONE_698  (
    .O(\DLX_EXinst_Mcompar__n0087_inst_cy_131/LOGIC_ONE )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0087_inst_cy_130_699 (
    .IA(\DLX_EXinst_Mcompar__n0087_inst_cy_131/LOGIC_ONE ),
    .IB(\DLX_EXinst_Mcompar__n0087_inst_cy_131/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0087_inst_lut4_28),
    .O(DLX_EXinst_Mcompar__n0087_inst_cy_130)
  );
  defparam DLX_EXinst_Mcompar__n0087_inst_lut4_281.INIT = 16'hC003;
  X_LUT4 DLX_EXinst_Mcompar__n0087_inst_lut4_281 (
    .ADR0(VCC),
    .ADR1(\DLX_IDinst_Imm[31] ),
    .ADR2(DLX_IDinst_reg_out_A[25]),
    .ADR3(DLX_IDinst_reg_out_A[24]),
    .O(DLX_EXinst_Mcompar__n0087_inst_lut4_28)
  );
  defparam DLX_EXinst_Mcompar__n0087_inst_lut4_291.INIT = 16'h8811;
  X_LUT4 DLX_EXinst_Mcompar__n0087_inst_lut4_291 (
    .ADR0(DLX_IDinst_reg_out_A[26]),
    .ADR1(\DLX_IDinst_Imm[31] ),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[27]),
    .O(DLX_EXinst_Mcompar__n0087_inst_lut4_29)
  );
  X_BUF \DLX_EXinst_Mcompar__n0087_inst_cy_131/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0087_inst_cy_131/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0087_inst_cy_131)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0087_inst_cy_131_700 (
    .IA(\DLX_EXinst_Mcompar__n0087_inst_cy_131/LOGIC_ONE ),
    .IB(DLX_EXinst_Mcompar__n0087_inst_cy_130),
    .SEL(DLX_EXinst_Mcompar__n0087_inst_lut4_29),
    .O(\DLX_EXinst_Mcompar__n0087_inst_cy_131/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0087_inst_cy_131/CYINIT_701  (
    .I(DLX_EXinst_Mcompar__n0087_inst_cy_129),
    .O(\DLX_EXinst_Mcompar__n0087_inst_cy_131/CYINIT )
  );
  X_ONE \DLX_EXinst__n0087/LOGIC_ONE_702  (
    .O(\DLX_EXinst__n0087/LOGIC_ONE )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0087_inst_cy_132_703 (
    .IA(\DLX_EXinst__n0087/LOGIC_ONE ),
    .IB(\DLX_EXinst__n0087/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0087_inst_lut4_30),
    .O(DLX_EXinst_Mcompar__n0087_inst_cy_132)
  );
  defparam DLX_EXinst_Mcompar__n0087_inst_lut4_301.INIT = 16'h8181;
  X_LUT4 DLX_EXinst_Mcompar__n0087_inst_lut4_301 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(DLX_IDinst_reg_out_A[28]),
    .ADR2(DLX_IDinst_reg_out_A[29]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0087_inst_lut4_30)
  );
  defparam DLX_EXinst_Mcompar__n0087_inst_lut4_311.INIT = 16'h8811;
  X_LUT4 DLX_EXinst_Mcompar__n0087_inst_lut4_311 (
    .ADR0(DLX_IDinst_reg_out_A[30]),
    .ADR1(DLX_IDinst_Imm_31_1),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[31]),
    .O(DLX_EXinst_Mcompar__n0087_inst_lut4_31)
  );
  X_BUF \DLX_EXinst__n0087/COUTUSED  (
    .I(\DLX_EXinst__n0087/CYMUXG ),
    .O(DLX_EXinst__n0087)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0087_inst_cy_133 (
    .IA(\DLX_EXinst__n0087/LOGIC_ONE ),
    .IB(DLX_EXinst_Mcompar__n0087_inst_cy_132),
    .SEL(DLX_EXinst_Mcompar__n0087_inst_lut4_31),
    .O(\DLX_EXinst__n0087/CYMUXG )
  );
  X_BUF \DLX_EXinst__n0087/CYINIT_704  (
    .I(DLX_EXinst_Mcompar__n0087_inst_cy_131),
    .O(\DLX_EXinst__n0087/CYINIT )
  );
  X_ZERO \DLX_EXinst_Mcompar__n0095_inst_cy_231/LOGIC_ZERO_705  (
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_231/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_230_706 (
    .IA(DLX_IDinst_IR_function_field_0_1),
    .IB(\DLX_EXinst_Mcompar__n0095_inst_cy_231/LOGIC_ZERO ),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_166),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_230)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1661.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1661 (
    .ADR0(DLX_IDinst_IR_function_field_0_1),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[0]),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_166)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1671.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1671 (
    .ADR0(DLX_IDinst_IR_function_field_1_1),
    .ADR1(DLX_IDinst_reg_out_A[1]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_167)
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_231/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0095_inst_cy_231/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_231)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_231_707 (
    .IA(DLX_IDinst_IR_function_field_1_1),
    .IB(DLX_EXinst_Mcompar__n0095_inst_cy_230),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_167),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_231/CYMUXG )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_232_708 (
    .IA(DLX_IDinst_IR_function_field_2_1),
    .IB(\DLX_EXinst_Mcompar__n0095_inst_cy_233/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_168),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_232)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1681.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1681 (
    .ADR0(DLX_IDinst_IR_function_field_2_1),
    .ADR1(DLX_IDinst_reg_out_A[2]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_168)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1691.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1691 (
    .ADR0(DLX_IDinst_IR_function_field_3_1),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[3]),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_169)
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_233/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0095_inst_cy_233/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_233)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_233_709 (
    .IA(DLX_IDinst_IR_function_field_3_1),
    .IB(DLX_EXinst_Mcompar__n0095_inst_cy_232),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_169),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_233/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_233/CYINIT_710  (
    .I(DLX_EXinst_Mcompar__n0095_inst_cy_231),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_233/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_234_711 (
    .IA(DLX_IDinst_IR_function_field[4]),
    .IB(\DLX_EXinst_Mcompar__n0095_inst_cy_235/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_170),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_234)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1701.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1701 (
    .ADR0(DLX_IDinst_IR_function_field[4]),
    .ADR1(DLX_IDinst_reg_out_A[4]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_170)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1711.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1711 (
    .ADR0(\DLX_IDinst_Imm[5] ),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[5]),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_171)
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_235/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0095_inst_cy_235/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_235)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_235_712 (
    .IA(\DLX_IDinst_Imm[5] ),
    .IB(DLX_EXinst_Mcompar__n0095_inst_cy_234),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_171),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_235/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_235/CYINIT_713  (
    .I(DLX_EXinst_Mcompar__n0095_inst_cy_233),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_235/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_236_714 (
    .IA(\DLX_IDinst_Imm[6] ),
    .IB(\DLX_EXinst_Mcompar__n0095_inst_cy_237/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_172),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_236)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1721.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1721 (
    .ADR0(\DLX_IDinst_Imm[6] ),
    .ADR1(DLX_IDinst_reg_out_A[6]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_172)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1731.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1731 (
    .ADR0(\DLX_IDinst_Imm[7] ),
    .ADR1(DLX_IDinst_reg_out_A[7]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_173)
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_237/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0095_inst_cy_237/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_237)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_237_715 (
    .IA(\DLX_IDinst_Imm[7] ),
    .IB(DLX_EXinst_Mcompar__n0095_inst_cy_236),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_173),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_237/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_237/CYINIT_716  (
    .I(DLX_EXinst_Mcompar__n0095_inst_cy_235),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_237/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_238_717 (
    .IA(\DLX_IDinst_Imm[8] ),
    .IB(\DLX_EXinst_Mcompar__n0095_inst_cy_239/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_174),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_238)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1741.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1741 (
    .ADR0(\DLX_IDinst_Imm[8] ),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[8]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_174)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1751.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1751 (
    .ADR0(\DLX_IDinst_Imm[9] ),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[9]),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_175)
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_239/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0095_inst_cy_239/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_239)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_239_718 (
    .IA(\DLX_IDinst_Imm[9] ),
    .IB(DLX_EXinst_Mcompar__n0095_inst_cy_238),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_175),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_239/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_239/CYINIT_719  (
    .I(DLX_EXinst_Mcompar__n0095_inst_cy_237),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_239/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_240_720 (
    .IA(\DLX_IDinst_Imm[10] ),
    .IB(\DLX_EXinst_Mcompar__n0095_inst_cy_241/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_176),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_240)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1761.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1761 (
    .ADR0(\DLX_IDinst_Imm[10] ),
    .ADR1(DLX_IDinst_reg_out_A[10]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_176)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1771.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1771 (
    .ADR0(\DLX_IDinst_Imm[11] ),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[11]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_177)
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_241/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0095_inst_cy_241/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_241)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_241_721 (
    .IA(\DLX_IDinst_Imm[11] ),
    .IB(DLX_EXinst_Mcompar__n0095_inst_cy_240),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_177),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_241/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_241/CYINIT_722  (
    .I(DLX_EXinst_Mcompar__n0095_inst_cy_239),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_241/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_242_723 (
    .IA(\DLX_IDinst_Imm[12] ),
    .IB(\DLX_EXinst_Mcompar__n0095_inst_cy_243/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_178),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_242)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1781.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1781 (
    .ADR0(\DLX_IDinst_Imm[12] ),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[12]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_178)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1791.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1791 (
    .ADR0(\DLX_IDinst_Imm[13] ),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[13]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_179)
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_243/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0095_inst_cy_243/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_243)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_243_724 (
    .IA(\DLX_IDinst_Imm[13] ),
    .IB(DLX_EXinst_Mcompar__n0095_inst_cy_242),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_179),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_243/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_243/CYINIT_725  (
    .I(DLX_EXinst_Mcompar__n0095_inst_cy_241),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_243/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_244_726 (
    .IA(\DLX_IDinst_Imm[14] ),
    .IB(\DLX_EXinst_Mcompar__n0095_inst_cy_245/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_180),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_244)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1801.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1801 (
    .ADR0(\DLX_IDinst_Imm[14] ),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[14]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_180)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1811.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1811 (
    .ADR0(\DLX_IDinst_Imm[15] ),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[15]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_181)
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_245/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0095_inst_cy_245/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_245)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_245_727 (
    .IA(\DLX_IDinst_Imm[15] ),
    .IB(DLX_EXinst_Mcompar__n0095_inst_cy_244),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_181),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_245/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_245/CYINIT_728  (
    .I(DLX_EXinst_Mcompar__n0095_inst_cy_243),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_245/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_246_729 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(\DLX_EXinst_Mcompar__n0095_inst_cy_247/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_182),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_246)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1821.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1821 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[16]),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_182)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1831.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1831 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[17]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_183)
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_247/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0095_inst_cy_247/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_247)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_247_730 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(DLX_EXinst_Mcompar__n0095_inst_cy_246),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_183),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_247/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_247/CYINIT_731  (
    .I(DLX_EXinst_Mcompar__n0095_inst_cy_245),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_247/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_248_732 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(\DLX_EXinst_Mcompar__n0095_inst_cy_249/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_184),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_248)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1841.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1841 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[18]),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_184)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1851.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1851 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[19]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_185)
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_249/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0095_inst_cy_249/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_249)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_249_733 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(DLX_EXinst_Mcompar__n0095_inst_cy_248),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_185),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_249/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_249/CYINIT_734  (
    .I(DLX_EXinst_Mcompar__n0095_inst_cy_247),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_249/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_250_735 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(\DLX_EXinst_Mcompar__n0095_inst_cy_251/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_186),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_250)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1861.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1861 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[20]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_186)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1871.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1871 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[21]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_187)
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_251/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0095_inst_cy_251/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_251)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_251_736 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(DLX_EXinst_Mcompar__n0095_inst_cy_250),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_187),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_251/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_251/CYINIT_737  (
    .I(DLX_EXinst_Mcompar__n0095_inst_cy_249),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_251/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_252_738 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(\DLX_EXinst_Mcompar__n0095_inst_cy_253/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_188),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_252)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1881.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1881 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(DLX_IDinst_reg_out_A[22]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_188)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1891.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1891 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(DLX_IDinst_reg_out_A[23]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_189)
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_253/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0095_inst_cy_253/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_253)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_253_739 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(DLX_EXinst_Mcompar__n0095_inst_cy_252),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_189),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_253/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_253/CYINIT_740  (
    .I(DLX_EXinst_Mcompar__n0095_inst_cy_251),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_253/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_254_741 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(\DLX_EXinst_Mcompar__n0095_inst_cy_255/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_190),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_254)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1901.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1901 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[24]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_190)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1911.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1911 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(DLX_IDinst_reg_out_A[25]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_191)
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_255/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0095_inst_cy_255/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_255)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_255_742 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(DLX_EXinst_Mcompar__n0095_inst_cy_254),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_191),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_255/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_255/CYINIT_743  (
    .I(DLX_EXinst_Mcompar__n0095_inst_cy_253),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_255/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_256_744 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(\DLX_EXinst_Mcompar__n0095_inst_cy_257/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_192),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_256)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1921.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1921 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(DLX_IDinst_reg_out_A[26]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_192)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1931.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1931 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(DLX_IDinst_reg_out_A[27]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_193)
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_257/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0095_inst_cy_257/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_257)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_257_745 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(DLX_EXinst_Mcompar__n0095_inst_cy_256),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_193),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_257/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_257/CYINIT_746  (
    .I(DLX_EXinst_Mcompar__n0095_inst_cy_255),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_257/CYINIT )
  );
  defparam DLX_IDinst_stall_1_747.INIT = 1'b0;
  X_FF DLX_IDinst_stall_1_747 (
    .I(\stall/OD ),
    .CE(DLX_IDinst__n0441),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\stall/OFF/RST ),
    .O(DLX_IDinst_stall_1)
  );
  X_OR2 \stall/OFF/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\stall/OFF/RST )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_258_748 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(\DLX_EXinst_Mcompar__n0095_inst_cy_259/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_194),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_258)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1941.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1941 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[28]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_194)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1951.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1951 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[29]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_195)
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_259/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0095_inst_cy_259/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_259)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_259_749 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(DLX_EXinst_Mcompar__n0095_inst_cy_258),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_195),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_259/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_259/CYINIT_750  (
    .I(DLX_EXinst_Mcompar__n0095_inst_cy_257),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_259/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_260_751 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(\CHOICE5769/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_196),
    .O(\CHOICE5769/CYMUXF )
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1961.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1961 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[30]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_196)
  );
  defparam \DLX_EXinst__n0006<31>84 .INIT = 16'h88A0;
  X_LUT4 \DLX_EXinst__n0006<31>84  (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(DLX_IDinst_reg_out_A[28]),
    .ADR2(DLX_IDinst_reg_out_A[30]),
    .ADR3(DLX_IDinst_reg_out_B[1]),
    .O(\CHOICE5769/GROM )
  );
  X_BUF \CHOICE5769/XBUSED  (
    .I(\CHOICE5769/CYMUXF ),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_260)
  );
  X_BUF \CHOICE5769/YUSED  (
    .I(\CHOICE5769/GROM ),
    .O(CHOICE5769)
  );
  X_BUF \CHOICE5769/CYINIT_752  (
    .I(DLX_EXinst_Mcompar__n0095_inst_cy_259),
    .O(\CHOICE5769/CYINIT )
  );
  X_ONE \vga_top_vga1_Mcompar__n0030_inst_cy_358/LOGIC_ONE_753  (
    .O(\vga_top_vga1_Mcompar__n0030_inst_cy_358/LOGIC_ONE )
  );
  X_ZERO \vga_top_vga1_Mcompar__n0030_inst_cy_358/LOGIC_ZERO_754  (
    .O(\vga_top_vga1_Mcompar__n0030_inst_cy_358/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0030_inst_cy_357_755 (
    .IA(\vga_top_vga1_Mcompar__n0030_inst_cy_358/LOGIC_ZERO ),
    .IB(\vga_top_vga1_Mcompar__n0030_inst_cy_358/LOGIC_ONE ),
    .SEL(vga_top_vga1_Mcompar__n0030_inst_lut4_48),
    .O(vga_top_vga1_Mcompar__n0030_inst_cy_357)
  );
  defparam vga_top_vga1_Mcompar__n0030_inst_lut4_481.INIT = 16'h8000;
  X_LUT4 vga_top_vga1_Mcompar__n0030_inst_lut4_481 (
    .ADR0(vga_top_vga1_hcounter[1]),
    .ADR1(vga_top_vga1_hcounter[3]),
    .ADR2(vga_top_vga1_hcounter[0]),
    .ADR3(vga_top_vga1_hcounter[2]),
    .O(vga_top_vga1_Mcompar__n0030_inst_lut4_48)
  );
  defparam vga_top_vga1_Mcompar__n0030_inst_lut4_491.INIT = 16'h8000;
  X_LUT4 vga_top_vga1_Mcompar__n0030_inst_lut4_491 (
    .ADR0(vga_top_vga1_hcounter[0]),
    .ADR1(vga_top_vga1_hcounter[1]),
    .ADR2(vga_top_vga1_hcounter[2]),
    .ADR3(vga_top_vga1_hcounter[3]),
    .O(vga_top_vga1_Mcompar__n0030_inst_lut4_49)
  );
  X_BUF \vga_top_vga1_Mcompar__n0030_inst_cy_358/COUTUSED  (
    .I(\vga_top_vga1_Mcompar__n0030_inst_cy_358/CYMUXG ),
    .O(vga_top_vga1_Mcompar__n0030_inst_cy_358)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0030_inst_cy_358_756 (
    .IA(\vga_top_vga1_Mcompar__n0030_inst_cy_358/LOGIC_ZERO ),
    .IB(vga_top_vga1_Mcompar__n0030_inst_cy_357),
    .SEL(vga_top_vga1_Mcompar__n0030_inst_lut4_49),
    .O(\vga_top_vga1_Mcompar__n0030_inst_cy_358/CYMUXG )
  );
  X_ONE \vga_top_vga1_Mcompar__n0030_inst_cy_360/LOGIC_ONE_757  (
    .O(\vga_top_vga1_Mcompar__n0030_inst_cy_360/LOGIC_ONE )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0030_inst_cy_359_758 (
    .IA(\vga_top_vga1_Mcompar__n0030_inst_cy_360/LOGIC_ONE ),
    .IB(\vga_top_vga1_Mcompar__n0030_inst_cy_360/CYINIT ),
    .SEL(vga_top_vga1_Mcompar__n0030_inst_lut1_10),
    .O(vga_top_vga1_Mcompar__n0030_inst_cy_359)
  );
  defparam vga_top_vga1_Mcompar__n0030_inst_lut1_101.INIT = 16'h00FF;
  X_LUT4 vga_top_vga1_Mcompar__n0030_inst_lut1_101 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[4]),
    .O(vga_top_vga1_Mcompar__n0030_inst_lut1_10)
  );
  defparam vga_top_vga1_Mcompar__n0030_inst_lut1_111.INIT = 16'h0F0F;
  X_LUT4 vga_top_vga1_Mcompar__n0030_inst_lut1_111 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_hcounter[4]),
    .ADR3(VCC),
    .O(vga_top_vga1_Mcompar__n0030_inst_lut1_11)
  );
  X_BUF \vga_top_vga1_Mcompar__n0030_inst_cy_360/COUTUSED  (
    .I(\vga_top_vga1_Mcompar__n0030_inst_cy_360/CYMUXG ),
    .O(vga_top_vga1_Mcompar__n0030_inst_cy_360)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0030_inst_cy_360_759 (
    .IA(\vga_top_vga1_Mcompar__n0030_inst_cy_360/LOGIC_ONE ),
    .IB(vga_top_vga1_Mcompar__n0030_inst_cy_359),
    .SEL(vga_top_vga1_Mcompar__n0030_inst_lut1_11),
    .O(\vga_top_vga1_Mcompar__n0030_inst_cy_360/CYMUXG )
  );
  X_BUF \vga_top_vga1_Mcompar__n0030_inst_cy_360/CYINIT_760  (
    .I(vga_top_vga1_Mcompar__n0030_inst_cy_358),
    .O(\vga_top_vga1_Mcompar__n0030_inst_cy_360/CYINIT )
  );
  X_ZERO \vga_top_vga1_Mcompar__n0030_inst_cy_362/LOGIC_ZERO_761  (
    .O(\vga_top_vga1_Mcompar__n0030_inst_cy_362/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0030_inst_cy_361_762 (
    .IA(\vga_top_vga1_Mcompar__n0030_inst_cy_362/LOGIC_ZERO ),
    .IB(\vga_top_vga1_Mcompar__n0030_inst_cy_362/CYINIT ),
    .SEL(\$SIG_0 ),
    .O(vga_top_vga1_Mcompar__n0030_inst_cy_361)
  );
  defparam \$BEL_0 .INIT = 16'hCCCC;
  X_LUT4 \$BEL_0  (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_hcounter[5]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\$SIG_0 )
  );
  defparam \$BEL_1 .INIT = 16'hAAAA;
  X_LUT4 \$BEL_1  (
    .ADR0(vga_top_vga1_hcounter[5]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\$SIG_1 )
  );
  X_BUF \vga_top_vga1_Mcompar__n0030_inst_cy_362/COUTUSED  (
    .I(\vga_top_vga1_Mcompar__n0030_inst_cy_362/CYMUXG ),
    .O(vga_top_vga1_Mcompar__n0030_inst_cy_362)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0030_inst_cy_362_763 (
    .IA(\vga_top_vga1_Mcompar__n0030_inst_cy_362/LOGIC_ZERO ),
    .IB(vga_top_vga1_Mcompar__n0030_inst_cy_361),
    .SEL(\$SIG_1 ),
    .O(\vga_top_vga1_Mcompar__n0030_inst_cy_362/CYMUXG )
  );
  X_BUF \vga_top_vga1_Mcompar__n0030_inst_cy_362/CYINIT_764  (
    .I(vga_top_vga1_Mcompar__n0030_inst_cy_360),
    .O(\vga_top_vga1_Mcompar__n0030_inst_cy_362/CYINIT )
  );
  X_ONE \vga_top_vga1_Mcompar__n0030_inst_cy_364/LOGIC_ONE_765  (
    .O(\vga_top_vga1_Mcompar__n0030_inst_cy_364/LOGIC_ONE )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0030_inst_cy_363_766 (
    .IA(\vga_top_vga1_Mcompar__n0030_inst_cy_364/LOGIC_ONE ),
    .IB(\vga_top_vga1_Mcompar__n0030_inst_cy_364/CYINIT ),
    .SEL(vga_top_vga1_Mcompar__n0030_inst_lut1_14),
    .O(vga_top_vga1_Mcompar__n0030_inst_cy_363)
  );
  defparam vga_top_vga1_Mcompar__n0030_inst_lut1_141.INIT = 16'h5555;
  X_LUT4 vga_top_vga1_Mcompar__n0030_inst_lut1_141 (
    .ADR0(vga_top_vga1_hcounter[6]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(vga_top_vga1_Mcompar__n0030_inst_lut1_14)
  );
  defparam vga_top_vga1_Mcompar__n0030_inst_lut1_151.INIT = 16'h00FF;
  X_LUT4 vga_top_vga1_Mcompar__n0030_inst_lut1_151 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[6]),
    .O(vga_top_vga1_Mcompar__n0030_inst_lut1_15)
  );
  X_BUF \vga_top_vga1_Mcompar__n0030_inst_cy_364/COUTUSED  (
    .I(\vga_top_vga1_Mcompar__n0030_inst_cy_364/CYMUXG ),
    .O(vga_top_vga1_Mcompar__n0030_inst_cy_364)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0030_inst_cy_364_767 (
    .IA(\vga_top_vga1_Mcompar__n0030_inst_cy_364/LOGIC_ONE ),
    .IB(vga_top_vga1_Mcompar__n0030_inst_cy_363),
    .SEL(vga_top_vga1_Mcompar__n0030_inst_lut1_15),
    .O(\vga_top_vga1_Mcompar__n0030_inst_cy_364/CYMUXG )
  );
  X_BUF \vga_top_vga1_Mcompar__n0030_inst_cy_364/CYINIT_768  (
    .I(vga_top_vga1_Mcompar__n0030_inst_cy_362),
    .O(\vga_top_vga1_Mcompar__n0030_inst_cy_364/CYINIT )
  );
  X_ZERO \vga_top_vga1_Mcompar__n0030_inst_cy_366/LOGIC_ZERO_769  (
    .O(\vga_top_vga1_Mcompar__n0030_inst_cy_366/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0030_inst_cy_365_770 (
    .IA(\vga_top_vga1_Mcompar__n0030_inst_cy_366/LOGIC_ZERO ),
    .IB(\vga_top_vga1_Mcompar__n0030_inst_cy_366/CYINIT ),
    .SEL(\$SIG_2 ),
    .O(vga_top_vga1_Mcompar__n0030_inst_cy_365)
  );
  defparam \$BEL_2 .INIT = 16'hF0F0;
  X_LUT4 \$BEL_2  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_hcounter[7]),
    .ADR3(VCC),
    .O(\$SIG_2 )
  );
  defparam \$BEL_3 .INIT = 16'hF0F0;
  X_LUT4 \$BEL_3  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_hcounter[7]),
    .ADR3(VCC),
    .O(\$SIG_3 )
  );
  X_BUF \vga_top_vga1_Mcompar__n0030_inst_cy_366/COUTUSED  (
    .I(\vga_top_vga1_Mcompar__n0030_inst_cy_366/CYMUXG ),
    .O(vga_top_vga1_Mcompar__n0030_inst_cy_366)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0030_inst_cy_366_771 (
    .IA(\vga_top_vga1_Mcompar__n0030_inst_cy_366/LOGIC_ZERO ),
    .IB(vga_top_vga1_Mcompar__n0030_inst_cy_365),
    .SEL(\$SIG_3 ),
    .O(\vga_top_vga1_Mcompar__n0030_inst_cy_366/CYMUXG )
  );
  X_BUF \vga_top_vga1_Mcompar__n0030_inst_cy_366/CYINIT_772  (
    .I(vga_top_vga1_Mcompar__n0030_inst_cy_364),
    .O(\vga_top_vga1_Mcompar__n0030_inst_cy_366/CYINIT )
  );
  X_ONE \vga_top_vga1_Mcompar__n0030_inst_cy_368/LOGIC_ONE_773  (
    .O(\vga_top_vga1_Mcompar__n0030_inst_cy_368/LOGIC_ONE )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0030_inst_cy_367_774 (
    .IA(\vga_top_vga1_Mcompar__n0030_inst_cy_368/LOGIC_ONE ),
    .IB(\vga_top_vga1_Mcompar__n0030_inst_cy_368/CYINIT ),
    .SEL(vga_top_vga1_Mcompar__n0030_inst_lut1_18),
    .O(vga_top_vga1_Mcompar__n0030_inst_cy_367)
  );
  defparam vga_top_vga1_Mcompar__n0030_inst_lut1_181.INIT = 16'h0F0F;
  X_LUT4 vga_top_vga1_Mcompar__n0030_inst_lut1_181 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_hcounter[8]),
    .ADR3(VCC),
    .O(vga_top_vga1_Mcompar__n0030_inst_lut1_18)
  );
  defparam vga_top_vga1_Mcompar__n0030_inst_lut1_191.INIT = 16'h3333;
  X_LUT4 vga_top_vga1_Mcompar__n0030_inst_lut1_191 (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_hcounter[8]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(vga_top_vga1_Mcompar__n0030_inst_lut1_19)
  );
  X_BUF \vga_top_vga1_Mcompar__n0030_inst_cy_368/COUTUSED  (
    .I(\vga_top_vga1_Mcompar__n0030_inst_cy_368/CYMUXG ),
    .O(vga_top_vga1_Mcompar__n0030_inst_cy_368)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0030_inst_cy_368_775 (
    .IA(\vga_top_vga1_Mcompar__n0030_inst_cy_368/LOGIC_ONE ),
    .IB(vga_top_vga1_Mcompar__n0030_inst_cy_367),
    .SEL(vga_top_vga1_Mcompar__n0030_inst_lut1_19),
    .O(\vga_top_vga1_Mcompar__n0030_inst_cy_368/CYMUXG )
  );
  X_BUF \vga_top_vga1_Mcompar__n0030_inst_cy_368/CYINIT_776  (
    .I(vga_top_vga1_Mcompar__n0030_inst_cy_366),
    .O(\vga_top_vga1_Mcompar__n0030_inst_cy_368/CYINIT )
  );
  X_ZERO \vga_top_vga1_Mcompar__n0030_inst_cy_370/LOGIC_ZERO_777  (
    .O(\vga_top_vga1_Mcompar__n0030_inst_cy_370/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0030_inst_cy_369_778 (
    .IA(\vga_top_vga1_Mcompar__n0030_inst_cy_370/LOGIC_ZERO ),
    .IB(\vga_top_vga1_Mcompar__n0030_inst_cy_370/CYINIT ),
    .SEL(\$SIG_4 ),
    .O(vga_top_vga1_Mcompar__n0030_inst_cy_369)
  );
  defparam \$BEL_4 .INIT = 16'hF0F0;
  X_LUT4 \$BEL_4  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_hcounter[9]),
    .ADR3(VCC),
    .O(\$SIG_4 )
  );
  defparam \$BEL_5 .INIT = 16'hFF00;
  X_LUT4 \$BEL_5  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[9]),
    .O(\$SIG_5 )
  );
  X_BUF \vga_top_vga1_Mcompar__n0030_inst_cy_370/COUTUSED  (
    .I(\vga_top_vga1_Mcompar__n0030_inst_cy_370/CYMUXG ),
    .O(vga_top_vga1_Mcompar__n0030_inst_cy_370)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0030_inst_cy_370_779 (
    .IA(\vga_top_vga1_Mcompar__n0030_inst_cy_370/LOGIC_ZERO ),
    .IB(vga_top_vga1_Mcompar__n0030_inst_cy_369),
    .SEL(\$SIG_5 ),
    .O(\vga_top_vga1_Mcompar__n0030_inst_cy_370/CYMUXG )
  );
  X_BUF \vga_top_vga1_Mcompar__n0030_inst_cy_370/CYINIT_780  (
    .I(vga_top_vga1_Mcompar__n0030_inst_cy_368),
    .O(\vga_top_vga1_Mcompar__n0030_inst_cy_370/CYINIT )
  );
  X_ONE \vga_top_vga1__n0030/LOGIC_ONE_781  (
    .O(\vga_top_vga1__n0030/LOGIC_ONE )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0030_inst_cy_371_782 (
    .IA(\vga_top_vga1__n0030/LOGIC_ONE ),
    .IB(\vga_top_vga1__n0030/CYINIT ),
    .SEL(vga_top_vga1_Mcompar__n0030_inst_lut4_50),
    .O(vga_top_vga1_Mcompar__n0030_inst_cy_371)
  );
  defparam vga_top_vga1_Mcompar__n0030_inst_lut4_501.INIT = 16'h0001;
  X_LUT4 vga_top_vga1_Mcompar__n0030_inst_lut4_501 (
    .ADR0(vga_top_vga1_hcounter[10]),
    .ADR1(vga_top_vga1_hcounter[12]),
    .ADR2(vga_top_vga1_hcounter[11]),
    .ADR3(vga_top_vga1_hcounter[13]),
    .O(vga_top_vga1_Mcompar__n0030_inst_lut4_50)
  );
  defparam vga_top_vga1_Mcompar__n0030_inst_lut2_2741.INIT = 16'h0055;
  X_LUT4 vga_top_vga1_Mcompar__n0030_inst_lut2_2741 (
    .ADR0(vga_top_vga1_hcounter[14]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[15]),
    .O(vga_top_vga1_Mcompar__n0030_inst_lut2_274)
  );
  X_BUF \vga_top_vga1__n0030/COUTUSED  (
    .I(\vga_top_vga1__n0030/CYMUXG ),
    .O(vga_top_vga1__n0030)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0030_inst_cy_372 (
    .IA(\vga_top_vga1__n0030/LOGIC_ONE ),
    .IB(vga_top_vga1_Mcompar__n0030_inst_cy_371),
    .SEL(vga_top_vga1_Mcompar__n0030_inst_lut2_274),
    .O(\vga_top_vga1__n0030/CYMUXG )
  );
  X_BUF \vga_top_vga1__n0030/CYINIT_783  (
    .I(vga_top_vga1_Mcompar__n0030_inst_cy_370),
    .O(\vga_top_vga1__n0030/CYINIT )
  );
  X_ZERO \DLX_IFinst__n0015<3>/LOGIC_ZERO_784  (
    .O(\DLX_IFinst__n0015<3>/LOGIC_ZERO )
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_40_785 (
    .IA(GLOBAL_LOGIC1),
    .IB(\DLX_IFinst__n0015<3>/LOGIC_ZERO ),
    .SEL(DLX_IFinst_Madd__n0005_inst_lut2_40),
    .O(DLX_IFinst_Madd__n0005_inst_cy_40)
  );
  defparam DLX_IFinst_Madd__n0005_inst_lut2_401.INIT = 16'h3333;
  X_LUT4 DLX_IFinst_Madd__n0005_inst_lut2_401 (
    .ADR0(GLOBAL_LOGIC1),
    .ADR1(DLX_IFinst_NPC[2]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IFinst_Madd__n0005_inst_lut2_40)
  );
  defparam \DLX_IFinst__n0015<3>/G .INIT = 16'hFF00;
  X_LUT4 \DLX_IFinst__n0015<3>/G  (
    .ADR0(GLOBAL_LOGIC0_10),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IFinst_NPC[3]),
    .O(\DLX_IFinst__n0015<3>/GROM )
  );
  X_BUF \DLX_IFinst__n0015<3>/COUTUSED  (
    .I(\DLX_IFinst__n0015<3>/CYMUXG ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_41)
  );
  X_BUF \DLX_IFinst__n0015<3>/YUSED  (
    .I(\DLX_IFinst__n0015<3>/XORG ),
    .O(DLX_IFinst__n0015[3])
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_41_786 (
    .IA(GLOBAL_LOGIC0_10),
    .IB(DLX_IFinst_Madd__n0005_inst_cy_40),
    .SEL(\DLX_IFinst__n0015<3>/GROM ),
    .O(\DLX_IFinst__n0015<3>/CYMUXG )
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_41 (
    .I0(DLX_IFinst_Madd__n0005_inst_cy_40),
    .I1(\DLX_IFinst__n0015<3>/GROM ),
    .O(\DLX_IFinst__n0015<3>/XORG )
  );
  X_ZERO \DLX_IFinst__n0015<4>/LOGIC_ZERO_787  (
    .O(\DLX_IFinst__n0015<4>/LOGIC_ZERO )
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_42_788 (
    .IA(\DLX_IFinst__n0015<4>/LOGIC_ZERO ),
    .IB(\DLX_IFinst__n0015<4>/CYINIT ),
    .SEL(\DLX_IFinst__n0015<4>/FROM ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_42)
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_42 (
    .I0(\DLX_IFinst__n0015<4>/CYINIT ),
    .I1(\DLX_IFinst__n0015<4>/FROM ),
    .O(\DLX_IFinst__n0015<4>/XORF )
  );
  defparam \DLX_IFinst__n0015<4>/F .INIT = 16'hF0F0;
  X_LUT4 \DLX_IFinst__n0015<4>/F  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IFinst_NPC[4]),
    .ADR3(VCC),
    .O(\DLX_IFinst__n0015<4>/FROM )
  );
  defparam \DLX_IFinst__n0015<4>/G .INIT = 16'hAAAA;
  X_LUT4 \DLX_IFinst__n0015<4>/G  (
    .ADR0(DLX_IFinst_NPC[5]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IFinst__n0015<4>/GROM )
  );
  X_BUF \DLX_IFinst__n0015<4>/COUTUSED  (
    .I(\DLX_IFinst__n0015<4>/CYMUXG ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_43)
  );
  X_BUF \DLX_IFinst__n0015<4>/XUSED  (
    .I(\DLX_IFinst__n0015<4>/XORF ),
    .O(DLX_IFinst__n0015[4])
  );
  X_BUF \DLX_IFinst__n0015<4>/YUSED  (
    .I(\DLX_IFinst__n0015<4>/XORG ),
    .O(DLX_IFinst__n0015[5])
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_43_789 (
    .IA(\DLX_IFinst__n0015<4>/LOGIC_ZERO ),
    .IB(DLX_IFinst_Madd__n0005_inst_cy_42),
    .SEL(\DLX_IFinst__n0015<4>/GROM ),
    .O(\DLX_IFinst__n0015<4>/CYMUXG )
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_43 (
    .I0(DLX_IFinst_Madd__n0005_inst_cy_42),
    .I1(\DLX_IFinst__n0015<4>/GROM ),
    .O(\DLX_IFinst__n0015<4>/XORG )
  );
  X_BUF \DLX_IFinst__n0015<4>/CYINIT_790  (
    .I(DLX_IFinst_Madd__n0005_inst_cy_41),
    .O(\DLX_IFinst__n0015<4>/CYINIT )
  );
  X_ZERO \DLX_IFinst__n0015<6>/LOGIC_ZERO_791  (
    .O(\DLX_IFinst__n0015<6>/LOGIC_ZERO )
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_44_792 (
    .IA(\DLX_IFinst__n0015<6>/LOGIC_ZERO ),
    .IB(\DLX_IFinst__n0015<6>/CYINIT ),
    .SEL(\DLX_IFinst__n0015<6>/FROM ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_44)
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_44 (
    .I0(\DLX_IFinst__n0015<6>/CYINIT ),
    .I1(\DLX_IFinst__n0015<6>/FROM ),
    .O(\DLX_IFinst__n0015<6>/XORF )
  );
  defparam \DLX_IFinst__n0015<6>/F .INIT = 16'hFF00;
  X_LUT4 \DLX_IFinst__n0015<6>/F  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IFinst_NPC[6]),
    .O(\DLX_IFinst__n0015<6>/FROM )
  );
  defparam \DLX_IFinst__n0015<6>/G .INIT = 16'hF0F0;
  X_LUT4 \DLX_IFinst__n0015<6>/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IFinst_NPC[7]),
    .ADR3(VCC),
    .O(\DLX_IFinst__n0015<6>/GROM )
  );
  X_BUF \DLX_IFinst__n0015<6>/COUTUSED  (
    .I(\DLX_IFinst__n0015<6>/CYMUXG ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_45)
  );
  X_BUF \DLX_IFinst__n0015<6>/XUSED  (
    .I(\DLX_IFinst__n0015<6>/XORF ),
    .O(DLX_IFinst__n0015[6])
  );
  X_BUF \DLX_IFinst__n0015<6>/YUSED  (
    .I(\DLX_IFinst__n0015<6>/XORG ),
    .O(DLX_IFinst__n0015[7])
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_45_793 (
    .IA(\DLX_IFinst__n0015<6>/LOGIC_ZERO ),
    .IB(DLX_IFinst_Madd__n0005_inst_cy_44),
    .SEL(\DLX_IFinst__n0015<6>/GROM ),
    .O(\DLX_IFinst__n0015<6>/CYMUXG )
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_45 (
    .I0(DLX_IFinst_Madd__n0005_inst_cy_44),
    .I1(\DLX_IFinst__n0015<6>/GROM ),
    .O(\DLX_IFinst__n0015<6>/XORG )
  );
  X_BUF \DLX_IFinst__n0015<6>/CYINIT_794  (
    .I(DLX_IFinst_Madd__n0005_inst_cy_43),
    .O(\DLX_IFinst__n0015<6>/CYINIT )
  );
  X_ZERO \DLX_IFinst__n0015<8>/LOGIC_ZERO_795  (
    .O(\DLX_IFinst__n0015<8>/LOGIC_ZERO )
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_46_796 (
    .IA(\DLX_IFinst__n0015<8>/LOGIC_ZERO ),
    .IB(\DLX_IFinst__n0015<8>/CYINIT ),
    .SEL(\DLX_IFinst__n0015<8>/FROM ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_46)
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_46 (
    .I0(\DLX_IFinst__n0015<8>/CYINIT ),
    .I1(\DLX_IFinst__n0015<8>/FROM ),
    .O(\DLX_IFinst__n0015<8>/XORF )
  );
  defparam \DLX_IFinst__n0015<8>/F .INIT = 16'hFF00;
  X_LUT4 \DLX_IFinst__n0015<8>/F  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IFinst_NPC[8]),
    .O(\DLX_IFinst__n0015<8>/FROM )
  );
  defparam \DLX_IFinst__n0015<8>/G .INIT = 16'hFF00;
  X_LUT4 \DLX_IFinst__n0015<8>/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IFinst_NPC[9]),
    .O(\DLX_IFinst__n0015<8>/GROM )
  );
  X_BUF \DLX_IFinst__n0015<8>/COUTUSED  (
    .I(\DLX_IFinst__n0015<8>/CYMUXG ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_47)
  );
  X_BUF \DLX_IFinst__n0015<8>/XUSED  (
    .I(\DLX_IFinst__n0015<8>/XORF ),
    .O(DLX_IFinst__n0015[8])
  );
  X_BUF \DLX_IFinst__n0015<8>/YUSED  (
    .I(\DLX_IFinst__n0015<8>/XORG ),
    .O(DLX_IFinst__n0015[9])
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_47_797 (
    .IA(\DLX_IFinst__n0015<8>/LOGIC_ZERO ),
    .IB(DLX_IFinst_Madd__n0005_inst_cy_46),
    .SEL(\DLX_IFinst__n0015<8>/GROM ),
    .O(\DLX_IFinst__n0015<8>/CYMUXG )
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_47 (
    .I0(DLX_IFinst_Madd__n0005_inst_cy_46),
    .I1(\DLX_IFinst__n0015<8>/GROM ),
    .O(\DLX_IFinst__n0015<8>/XORG )
  );
  X_BUF \DLX_IFinst__n0015<8>/CYINIT_798  (
    .I(DLX_IFinst_Madd__n0005_inst_cy_45),
    .O(\DLX_IFinst__n0015<8>/CYINIT )
  );
  X_ZERO \DLX_IFinst__n0015<10>/LOGIC_ZERO_799  (
    .O(\DLX_IFinst__n0015<10>/LOGIC_ZERO )
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_48_800 (
    .IA(\DLX_IFinst__n0015<10>/LOGIC_ZERO ),
    .IB(\DLX_IFinst__n0015<10>/CYINIT ),
    .SEL(\DLX_IFinst__n0015<10>/FROM ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_48)
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_48 (
    .I0(\DLX_IFinst__n0015<10>/CYINIT ),
    .I1(\DLX_IFinst__n0015<10>/FROM ),
    .O(\DLX_IFinst__n0015<10>/XORF )
  );
  defparam \DLX_IFinst__n0015<10>/F .INIT = 16'hFF00;
  X_LUT4 \DLX_IFinst__n0015<10>/F  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IFinst_NPC[10]),
    .O(\DLX_IFinst__n0015<10>/FROM )
  );
  defparam \DLX_IFinst__n0015<10>/G .INIT = 16'hF0F0;
  X_LUT4 \DLX_IFinst__n0015<10>/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IFinst_NPC[11]),
    .ADR3(VCC),
    .O(\DLX_IFinst__n0015<10>/GROM )
  );
  X_BUF \DLX_IFinst__n0015<10>/COUTUSED  (
    .I(\DLX_IFinst__n0015<10>/CYMUXG ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_49)
  );
  X_BUF \DLX_IFinst__n0015<10>/XUSED  (
    .I(\DLX_IFinst__n0015<10>/XORF ),
    .O(DLX_IFinst__n0015[10])
  );
  X_BUF \DLX_IFinst__n0015<10>/YUSED  (
    .I(\DLX_IFinst__n0015<10>/XORG ),
    .O(DLX_IFinst__n0015[11])
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_49_801 (
    .IA(\DLX_IFinst__n0015<10>/LOGIC_ZERO ),
    .IB(DLX_IFinst_Madd__n0005_inst_cy_48),
    .SEL(\DLX_IFinst__n0015<10>/GROM ),
    .O(\DLX_IFinst__n0015<10>/CYMUXG )
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_49 (
    .I0(DLX_IFinst_Madd__n0005_inst_cy_48),
    .I1(\DLX_IFinst__n0015<10>/GROM ),
    .O(\DLX_IFinst__n0015<10>/XORG )
  );
  X_BUF \DLX_IFinst__n0015<10>/CYINIT_802  (
    .I(DLX_IFinst_Madd__n0005_inst_cy_47),
    .O(\DLX_IFinst__n0015<10>/CYINIT )
  );
  X_ZERO \DLX_IFinst__n0015<12>/LOGIC_ZERO_803  (
    .O(\DLX_IFinst__n0015<12>/LOGIC_ZERO )
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_50_804 (
    .IA(\DLX_IFinst__n0015<12>/LOGIC_ZERO ),
    .IB(\DLX_IFinst__n0015<12>/CYINIT ),
    .SEL(\DLX_IFinst__n0015<12>/FROM ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_50)
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_50 (
    .I0(\DLX_IFinst__n0015<12>/CYINIT ),
    .I1(\DLX_IFinst__n0015<12>/FROM ),
    .O(\DLX_IFinst__n0015<12>/XORF )
  );
  defparam \DLX_IFinst__n0015<12>/F .INIT = 16'hAAAA;
  X_LUT4 \DLX_IFinst__n0015<12>/F  (
    .ADR0(DLX_IFinst_NPC[12]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IFinst__n0015<12>/FROM )
  );
  defparam \DLX_IFinst__n0015<12>/G .INIT = 16'hCCCC;
  X_LUT4 \DLX_IFinst__n0015<12>/G  (
    .ADR0(VCC),
    .ADR1(DLX_IFinst_NPC[13]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IFinst__n0015<12>/GROM )
  );
  X_BUF \DLX_IFinst__n0015<12>/COUTUSED  (
    .I(\DLX_IFinst__n0015<12>/CYMUXG ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_51)
  );
  X_BUF \DLX_IFinst__n0015<12>/XUSED  (
    .I(\DLX_IFinst__n0015<12>/XORF ),
    .O(DLX_IFinst__n0015[12])
  );
  X_BUF \DLX_IFinst__n0015<12>/YUSED  (
    .I(\DLX_IFinst__n0015<12>/XORG ),
    .O(DLX_IFinst__n0015[13])
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_51_805 (
    .IA(\DLX_IFinst__n0015<12>/LOGIC_ZERO ),
    .IB(DLX_IFinst_Madd__n0005_inst_cy_50),
    .SEL(\DLX_IFinst__n0015<12>/GROM ),
    .O(\DLX_IFinst__n0015<12>/CYMUXG )
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_51 (
    .I0(DLX_IFinst_Madd__n0005_inst_cy_50),
    .I1(\DLX_IFinst__n0015<12>/GROM ),
    .O(\DLX_IFinst__n0015<12>/XORG )
  );
  X_BUF \DLX_IFinst__n0015<12>/CYINIT_806  (
    .I(DLX_IFinst_Madd__n0005_inst_cy_49),
    .O(\DLX_IFinst__n0015<12>/CYINIT )
  );
  X_ZERO \DLX_IFinst__n0015<14>/LOGIC_ZERO_807  (
    .O(\DLX_IFinst__n0015<14>/LOGIC_ZERO )
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_52_808 (
    .IA(\DLX_IFinst__n0015<14>/LOGIC_ZERO ),
    .IB(\DLX_IFinst__n0015<14>/CYINIT ),
    .SEL(\DLX_IFinst__n0015<14>/FROM ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_52)
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_52 (
    .I0(\DLX_IFinst__n0015<14>/CYINIT ),
    .I1(\DLX_IFinst__n0015<14>/FROM ),
    .O(\DLX_IFinst__n0015<14>/XORF )
  );
  defparam \DLX_IFinst__n0015<14>/F .INIT = 16'hCCCC;
  X_LUT4 \DLX_IFinst__n0015<14>/F  (
    .ADR0(VCC),
    .ADR1(DLX_IFinst_NPC[14]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IFinst__n0015<14>/FROM )
  );
  defparam \DLX_IFinst__n0015<14>/G .INIT = 16'hFF00;
  X_LUT4 \DLX_IFinst__n0015<14>/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IFinst_NPC[15]),
    .O(\DLX_IFinst__n0015<14>/GROM )
  );
  X_BUF \DLX_IFinst__n0015<14>/COUTUSED  (
    .I(\DLX_IFinst__n0015<14>/CYMUXG ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_53)
  );
  X_BUF \DLX_IFinst__n0015<14>/XUSED  (
    .I(\DLX_IFinst__n0015<14>/XORF ),
    .O(DLX_IFinst__n0015[14])
  );
  X_BUF \DLX_IFinst__n0015<14>/YUSED  (
    .I(\DLX_IFinst__n0015<14>/XORG ),
    .O(DLX_IFinst__n0015[15])
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_53_809 (
    .IA(\DLX_IFinst__n0015<14>/LOGIC_ZERO ),
    .IB(DLX_IFinst_Madd__n0005_inst_cy_52),
    .SEL(\DLX_IFinst__n0015<14>/GROM ),
    .O(\DLX_IFinst__n0015<14>/CYMUXG )
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_53 (
    .I0(DLX_IFinst_Madd__n0005_inst_cy_52),
    .I1(\DLX_IFinst__n0015<14>/GROM ),
    .O(\DLX_IFinst__n0015<14>/XORG )
  );
  X_BUF \DLX_IFinst__n0015<14>/CYINIT_810  (
    .I(DLX_IFinst_Madd__n0005_inst_cy_51),
    .O(\DLX_IFinst__n0015<14>/CYINIT )
  );
  X_ZERO \DLX_IFinst__n0015<16>/LOGIC_ZERO_811  (
    .O(\DLX_IFinst__n0015<16>/LOGIC_ZERO )
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_54_812 (
    .IA(\DLX_IFinst__n0015<16>/LOGIC_ZERO ),
    .IB(\DLX_IFinst__n0015<16>/CYINIT ),
    .SEL(\DLX_IFinst__n0015<16>/FROM ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_54)
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_54 (
    .I0(\DLX_IFinst__n0015<16>/CYINIT ),
    .I1(\DLX_IFinst__n0015<16>/FROM ),
    .O(\DLX_IFinst__n0015<16>/XORF )
  );
  defparam \DLX_IFinst__n0015<16>/F .INIT = 16'hF0F0;
  X_LUT4 \DLX_IFinst__n0015<16>/F  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IFinst_NPC[16]),
    .ADR3(VCC),
    .O(\DLX_IFinst__n0015<16>/FROM )
  );
  defparam \DLX_IFinst__n0015<16>/G .INIT = 16'hCCCC;
  X_LUT4 \DLX_IFinst__n0015<16>/G  (
    .ADR0(VCC),
    .ADR1(DLX_IFinst_NPC[17]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IFinst__n0015<16>/GROM )
  );
  X_BUF \DLX_IFinst__n0015<16>/COUTUSED  (
    .I(\DLX_IFinst__n0015<16>/CYMUXG ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_55)
  );
  X_BUF \DLX_IFinst__n0015<16>/XUSED  (
    .I(\DLX_IFinst__n0015<16>/XORF ),
    .O(DLX_IFinst__n0015[16])
  );
  X_BUF \DLX_IFinst__n0015<16>/YUSED  (
    .I(\DLX_IFinst__n0015<16>/XORG ),
    .O(DLX_IFinst__n0015[17])
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_55_813 (
    .IA(\DLX_IFinst__n0015<16>/LOGIC_ZERO ),
    .IB(DLX_IFinst_Madd__n0005_inst_cy_54),
    .SEL(\DLX_IFinst__n0015<16>/GROM ),
    .O(\DLX_IFinst__n0015<16>/CYMUXG )
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_55 (
    .I0(DLX_IFinst_Madd__n0005_inst_cy_54),
    .I1(\DLX_IFinst__n0015<16>/GROM ),
    .O(\DLX_IFinst__n0015<16>/XORG )
  );
  X_BUF \DLX_IFinst__n0015<16>/CYINIT_814  (
    .I(DLX_IFinst_Madd__n0005_inst_cy_53),
    .O(\DLX_IFinst__n0015<16>/CYINIT )
  );
  defparam DLX_IDinst_CLI_1_815.INIT = 1'b0;
  X_FF DLX_IDinst_CLI_1_815 (
    .I(\CLI/OD ),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\CLI/OFF/RST ),
    .O(DLX_IDinst_CLI_1)
  );
  X_OR2 \CLI/OFF/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\CLI/OFF/RST )
  );
  X_ZERO \DLX_IFinst__n0015<18>/LOGIC_ZERO_816  (
    .O(\DLX_IFinst__n0015<18>/LOGIC_ZERO )
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_56_817 (
    .IA(\DLX_IFinst__n0015<18>/LOGIC_ZERO ),
    .IB(\DLX_IFinst__n0015<18>/CYINIT ),
    .SEL(\DLX_IFinst__n0015<18>/FROM ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_56)
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_56 (
    .I0(\DLX_IFinst__n0015<18>/CYINIT ),
    .I1(\DLX_IFinst__n0015<18>/FROM ),
    .O(\DLX_IFinst__n0015<18>/XORF )
  );
  defparam \DLX_IFinst__n0015<18>/F .INIT = 16'hCCCC;
  X_LUT4 \DLX_IFinst__n0015<18>/F  (
    .ADR0(VCC),
    .ADR1(DLX_IFinst_NPC[18]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IFinst__n0015<18>/FROM )
  );
  defparam \DLX_IFinst__n0015<18>/G .INIT = 16'hFF00;
  X_LUT4 \DLX_IFinst__n0015<18>/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IFinst_NPC[19]),
    .O(\DLX_IFinst__n0015<18>/GROM )
  );
  X_BUF \DLX_IFinst__n0015<18>/COUTUSED  (
    .I(\DLX_IFinst__n0015<18>/CYMUXG ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_57)
  );
  X_BUF \DLX_IFinst__n0015<18>/XUSED  (
    .I(\DLX_IFinst__n0015<18>/XORF ),
    .O(DLX_IFinst__n0015[18])
  );
  X_BUF \DLX_IFinst__n0015<18>/YUSED  (
    .I(\DLX_IFinst__n0015<18>/XORG ),
    .O(DLX_IFinst__n0015[19])
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_57_818 (
    .IA(\DLX_IFinst__n0015<18>/LOGIC_ZERO ),
    .IB(DLX_IFinst_Madd__n0005_inst_cy_56),
    .SEL(\DLX_IFinst__n0015<18>/GROM ),
    .O(\DLX_IFinst__n0015<18>/CYMUXG )
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_57 (
    .I0(DLX_IFinst_Madd__n0005_inst_cy_56),
    .I1(\DLX_IFinst__n0015<18>/GROM ),
    .O(\DLX_IFinst__n0015<18>/XORG )
  );
  X_BUF \DLX_IFinst__n0015<18>/CYINIT_819  (
    .I(DLX_IFinst_Madd__n0005_inst_cy_55),
    .O(\DLX_IFinst__n0015<18>/CYINIT )
  );
  X_ZERO \DLX_IFinst__n0015<20>/LOGIC_ZERO_820  (
    .O(\DLX_IFinst__n0015<20>/LOGIC_ZERO )
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_58_821 (
    .IA(\DLX_IFinst__n0015<20>/LOGIC_ZERO ),
    .IB(\DLX_IFinst__n0015<20>/CYINIT ),
    .SEL(\DLX_IFinst__n0015<20>/FROM ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_58)
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_58 (
    .I0(\DLX_IFinst__n0015<20>/CYINIT ),
    .I1(\DLX_IFinst__n0015<20>/FROM ),
    .O(\DLX_IFinst__n0015<20>/XORF )
  );
  defparam \DLX_IFinst__n0015<20>/F .INIT = 16'hCCCC;
  X_LUT4 \DLX_IFinst__n0015<20>/F  (
    .ADR0(VCC),
    .ADR1(DLX_IFinst_NPC[20]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IFinst__n0015<20>/FROM )
  );
  defparam \DLX_IFinst__n0015<20>/G .INIT = 16'hAAAA;
  X_LUT4 \DLX_IFinst__n0015<20>/G  (
    .ADR0(DLX_IFinst_NPC[21]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IFinst__n0015<20>/GROM )
  );
  X_BUF \DLX_IFinst__n0015<20>/COUTUSED  (
    .I(\DLX_IFinst__n0015<20>/CYMUXG ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_59)
  );
  X_BUF \DLX_IFinst__n0015<20>/XUSED  (
    .I(\DLX_IFinst__n0015<20>/XORF ),
    .O(DLX_IFinst__n0015[20])
  );
  X_BUF \DLX_IFinst__n0015<20>/YUSED  (
    .I(\DLX_IFinst__n0015<20>/XORG ),
    .O(DLX_IFinst__n0015[21])
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_59_822 (
    .IA(\DLX_IFinst__n0015<20>/LOGIC_ZERO ),
    .IB(DLX_IFinst_Madd__n0005_inst_cy_58),
    .SEL(\DLX_IFinst__n0015<20>/GROM ),
    .O(\DLX_IFinst__n0015<20>/CYMUXG )
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_59 (
    .I0(DLX_IFinst_Madd__n0005_inst_cy_58),
    .I1(\DLX_IFinst__n0015<20>/GROM ),
    .O(\DLX_IFinst__n0015<20>/XORG )
  );
  X_BUF \DLX_IFinst__n0015<20>/CYINIT_823  (
    .I(DLX_IFinst_Madd__n0005_inst_cy_57),
    .O(\DLX_IFinst__n0015<20>/CYINIT )
  );
  X_ZERO \DLX_IFinst__n0015<22>/LOGIC_ZERO_824  (
    .O(\DLX_IFinst__n0015<22>/LOGIC_ZERO )
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_60_825 (
    .IA(\DLX_IFinst__n0015<22>/LOGIC_ZERO ),
    .IB(\DLX_IFinst__n0015<22>/CYINIT ),
    .SEL(\DLX_IFinst__n0015<22>/FROM ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_60)
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_60 (
    .I0(\DLX_IFinst__n0015<22>/CYINIT ),
    .I1(\DLX_IFinst__n0015<22>/FROM ),
    .O(\DLX_IFinst__n0015<22>/XORF )
  );
  defparam \DLX_IFinst__n0015<22>/F .INIT = 16'hF0F0;
  X_LUT4 \DLX_IFinst__n0015<22>/F  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IFinst_NPC[22]),
    .ADR3(VCC),
    .O(\DLX_IFinst__n0015<22>/FROM )
  );
  defparam \DLX_IFinst__n0015<22>/G .INIT = 16'hAAAA;
  X_LUT4 \DLX_IFinst__n0015<22>/G  (
    .ADR0(DLX_IFinst_NPC[23]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IFinst__n0015<22>/GROM )
  );
  X_BUF \DLX_IFinst__n0015<22>/COUTUSED  (
    .I(\DLX_IFinst__n0015<22>/CYMUXG ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_61)
  );
  X_BUF \DLX_IFinst__n0015<22>/XUSED  (
    .I(\DLX_IFinst__n0015<22>/XORF ),
    .O(DLX_IFinst__n0015[22])
  );
  X_BUF \DLX_IFinst__n0015<22>/YUSED  (
    .I(\DLX_IFinst__n0015<22>/XORG ),
    .O(DLX_IFinst__n0015[23])
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_61_826 (
    .IA(\DLX_IFinst__n0015<22>/LOGIC_ZERO ),
    .IB(DLX_IFinst_Madd__n0005_inst_cy_60),
    .SEL(\DLX_IFinst__n0015<22>/GROM ),
    .O(\DLX_IFinst__n0015<22>/CYMUXG )
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_61 (
    .I0(DLX_IFinst_Madd__n0005_inst_cy_60),
    .I1(\DLX_IFinst__n0015<22>/GROM ),
    .O(\DLX_IFinst__n0015<22>/XORG )
  );
  X_BUF \DLX_IFinst__n0015<22>/CYINIT_827  (
    .I(DLX_IFinst_Madd__n0005_inst_cy_59),
    .O(\DLX_IFinst__n0015<22>/CYINIT )
  );
  X_ZERO \DLX_IFinst__n0015<24>/LOGIC_ZERO_828  (
    .O(\DLX_IFinst__n0015<24>/LOGIC_ZERO )
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_62_829 (
    .IA(\DLX_IFinst__n0015<24>/LOGIC_ZERO ),
    .IB(\DLX_IFinst__n0015<24>/CYINIT ),
    .SEL(\DLX_IFinst__n0015<24>/FROM ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_62)
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_62 (
    .I0(\DLX_IFinst__n0015<24>/CYINIT ),
    .I1(\DLX_IFinst__n0015<24>/FROM ),
    .O(\DLX_IFinst__n0015<24>/XORF )
  );
  defparam \DLX_IFinst__n0015<24>/F .INIT = 16'hAAAA;
  X_LUT4 \DLX_IFinst__n0015<24>/F  (
    .ADR0(DLX_IFinst_NPC[24]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IFinst__n0015<24>/FROM )
  );
  defparam \DLX_IFinst__n0015<24>/G .INIT = 16'hFF00;
  X_LUT4 \DLX_IFinst__n0015<24>/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IFinst_NPC[25]),
    .O(\DLX_IFinst__n0015<24>/GROM )
  );
  X_BUF \DLX_IFinst__n0015<24>/COUTUSED  (
    .I(\DLX_IFinst__n0015<24>/CYMUXG ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_63)
  );
  X_BUF \DLX_IFinst__n0015<24>/XUSED  (
    .I(\DLX_IFinst__n0015<24>/XORF ),
    .O(DLX_IFinst__n0015[24])
  );
  X_BUF \DLX_IFinst__n0015<24>/YUSED  (
    .I(\DLX_IFinst__n0015<24>/XORG ),
    .O(DLX_IFinst__n0015[25])
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_63_830 (
    .IA(\DLX_IFinst__n0015<24>/LOGIC_ZERO ),
    .IB(DLX_IFinst_Madd__n0005_inst_cy_62),
    .SEL(\DLX_IFinst__n0015<24>/GROM ),
    .O(\DLX_IFinst__n0015<24>/CYMUXG )
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_63 (
    .I0(DLX_IFinst_Madd__n0005_inst_cy_62),
    .I1(\DLX_IFinst__n0015<24>/GROM ),
    .O(\DLX_IFinst__n0015<24>/XORG )
  );
  X_BUF \DLX_IFinst__n0015<24>/CYINIT_831  (
    .I(DLX_IFinst_Madd__n0005_inst_cy_61),
    .O(\DLX_IFinst__n0015<24>/CYINIT )
  );
  X_ZERO \DLX_IFinst__n0015<26>/LOGIC_ZERO_832  (
    .O(\DLX_IFinst__n0015<26>/LOGIC_ZERO )
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_64_833 (
    .IA(\DLX_IFinst__n0015<26>/LOGIC_ZERO ),
    .IB(\DLX_IFinst__n0015<26>/CYINIT ),
    .SEL(\DLX_IFinst__n0015<26>/FROM ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_64)
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_64 (
    .I0(\DLX_IFinst__n0015<26>/CYINIT ),
    .I1(\DLX_IFinst__n0015<26>/FROM ),
    .O(\DLX_IFinst__n0015<26>/XORF )
  );
  defparam \DLX_IFinst__n0015<26>/F .INIT = 16'hCCCC;
  X_LUT4 \DLX_IFinst__n0015<26>/F  (
    .ADR0(VCC),
    .ADR1(DLX_IFinst_NPC[26]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IFinst__n0015<26>/FROM )
  );
  defparam \DLX_IFinst__n0015<26>/G .INIT = 16'hFF00;
  X_LUT4 \DLX_IFinst__n0015<26>/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IFinst_NPC[27]),
    .O(\DLX_IFinst__n0015<26>/GROM )
  );
  X_BUF \DLX_IFinst__n0015<26>/COUTUSED  (
    .I(\DLX_IFinst__n0015<26>/CYMUXG ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_65)
  );
  X_BUF \DLX_IFinst__n0015<26>/XUSED  (
    .I(\DLX_IFinst__n0015<26>/XORF ),
    .O(DLX_IFinst__n0015[26])
  );
  X_BUF \DLX_IFinst__n0015<26>/YUSED  (
    .I(\DLX_IFinst__n0015<26>/XORG ),
    .O(DLX_IFinst__n0015[27])
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_65_834 (
    .IA(\DLX_IFinst__n0015<26>/LOGIC_ZERO ),
    .IB(DLX_IFinst_Madd__n0005_inst_cy_64),
    .SEL(\DLX_IFinst__n0015<26>/GROM ),
    .O(\DLX_IFinst__n0015<26>/CYMUXG )
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_65 (
    .I0(DLX_IFinst_Madd__n0005_inst_cy_64),
    .I1(\DLX_IFinst__n0015<26>/GROM ),
    .O(\DLX_IFinst__n0015<26>/XORG )
  );
  X_BUF \DLX_IFinst__n0015<26>/CYINIT_835  (
    .I(DLX_IFinst_Madd__n0005_inst_cy_63),
    .O(\DLX_IFinst__n0015<26>/CYINIT )
  );
  X_ZERO \DLX_IFinst__n0015<28>/LOGIC_ZERO_836  (
    .O(\DLX_IFinst__n0015<28>/LOGIC_ZERO )
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_66_837 (
    .IA(\DLX_IFinst__n0015<28>/LOGIC_ZERO ),
    .IB(\DLX_IFinst__n0015<28>/CYINIT ),
    .SEL(\DLX_IFinst__n0015<28>/FROM ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_66)
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_66 (
    .I0(\DLX_IFinst__n0015<28>/CYINIT ),
    .I1(\DLX_IFinst__n0015<28>/FROM ),
    .O(\DLX_IFinst__n0015<28>/XORF )
  );
  defparam \DLX_IFinst__n0015<28>/F .INIT = 16'hAAAA;
  X_LUT4 \DLX_IFinst__n0015<28>/F  (
    .ADR0(DLX_IFinst_NPC[28]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IFinst__n0015<28>/FROM )
  );
  defparam \DLX_IFinst__n0015<28>/G .INIT = 16'hAAAA;
  X_LUT4 \DLX_IFinst__n0015<28>/G  (
    .ADR0(DLX_IFinst_NPC[29]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IFinst__n0015<28>/GROM )
  );
  X_BUF \DLX_IFinst__n0015<28>/COUTUSED  (
    .I(\DLX_IFinst__n0015<28>/CYMUXG ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_67)
  );
  X_BUF \DLX_IFinst__n0015<28>/XUSED  (
    .I(\DLX_IFinst__n0015<28>/XORF ),
    .O(DLX_IFinst__n0015[28])
  );
  X_BUF \DLX_IFinst__n0015<28>/YUSED  (
    .I(\DLX_IFinst__n0015<28>/XORG ),
    .O(DLX_IFinst__n0015[29])
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_67_838 (
    .IA(\DLX_IFinst__n0015<28>/LOGIC_ZERO ),
    .IB(DLX_IFinst_Madd__n0005_inst_cy_66),
    .SEL(\DLX_IFinst__n0015<28>/GROM ),
    .O(\DLX_IFinst__n0015<28>/CYMUXG )
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_67 (
    .I0(DLX_IFinst_Madd__n0005_inst_cy_66),
    .I1(\DLX_IFinst__n0015<28>/GROM ),
    .O(\DLX_IFinst__n0015<28>/XORG )
  );
  X_BUF \DLX_IFinst__n0015<28>/CYINIT_839  (
    .I(DLX_IFinst_Madd__n0005_inst_cy_65),
    .O(\DLX_IFinst__n0015<28>/CYINIT )
  );
  X_ZERO \DLX_IFinst__n0015<30>/LOGIC_ZERO_840  (
    .O(\DLX_IFinst__n0015<30>/LOGIC_ZERO )
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_68_841 (
    .IA(\DLX_IFinst__n0015<30>/LOGIC_ZERO ),
    .IB(\DLX_IFinst__n0015<30>/CYINIT ),
    .SEL(\DLX_IFinst__n0015<30>/FROM ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_68)
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_68 (
    .I0(\DLX_IFinst__n0015<30>/CYINIT ),
    .I1(\DLX_IFinst__n0015<30>/FROM ),
    .O(\DLX_IFinst__n0015<30>/XORF )
  );
  defparam \DLX_IFinst__n0015<30>/F .INIT = 16'hCCCC;
  X_LUT4 \DLX_IFinst__n0015<30>/F  (
    .ADR0(VCC),
    .ADR1(DLX_IFinst_NPC[30]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IFinst__n0015<30>/FROM )
  );
  defparam \DLX_IFinst_NPC<31>_rt_842 .INIT = 16'hF0F0;
  X_LUT4 \DLX_IFinst_NPC<31>_rt_842  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IFinst_NPC[31]),
    .ADR3(VCC),
    .O(\DLX_IFinst_NPC<31>_rt )
  );
  X_BUF \DLX_IFinst__n0015<30>/XUSED  (
    .I(\DLX_IFinst__n0015<30>/XORF ),
    .O(DLX_IFinst__n0015[30])
  );
  X_BUF \DLX_IFinst__n0015<30>/YUSED  (
    .I(\DLX_IFinst__n0015<30>/XORG ),
    .O(DLX_IFinst__n0015[31])
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_69 (
    .I0(DLX_IFinst_Madd__n0005_inst_cy_68),
    .I1(\DLX_IFinst_NPC<31>_rt ),
    .O(\DLX_IFinst__n0015<30>/XORG )
  );
  X_BUF \DLX_IFinst__n0015<30>/CYINIT_843  (
    .I(DLX_IFinst_Madd__n0005_inst_cy_67),
    .O(\DLX_IFinst__n0015<30>/CYINIT )
  );
  X_ZERO \DLX_EXinst_Mcompar__n0089_inst_cy_135/LOGIC_ZERO_844  (
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_135/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_134_845 (
    .IA(DLX_IDinst_IR_function_field_0_1),
    .IB(\DLX_EXinst_Mcompar__n0089_inst_cy_135/LOGIC_ZERO ),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_70),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_134)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_701.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_701 (
    .ADR0(DLX_IDinst_IR_function_field_0_1),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[0]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_70)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_711.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_711 (
    .ADR0(DLX_IDinst_IR_function_field_1_1),
    .ADR1(DLX_IDinst_reg_out_A[1]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_71)
  );
  X_BUF \DLX_EXinst_Mcompar__n0089_inst_cy_135/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0089_inst_cy_135/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_135)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_135_846 (
    .IA(DLX_IDinst_IR_function_field_1_1),
    .IB(DLX_EXinst_Mcompar__n0089_inst_cy_134),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_71),
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_135/CYMUXG )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_136_847 (
    .IA(DLX_IDinst_IR_function_field_2_1),
    .IB(\DLX_EXinst_Mcompar__n0089_inst_cy_137/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_72),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_136)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_721.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_721 (
    .ADR0(DLX_IDinst_IR_function_field_2_1),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[2]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_72)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_731.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_731 (
    .ADR0(DLX_IDinst_IR_function_field_3_1),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[3]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_73)
  );
  X_BUF \DLX_EXinst_Mcompar__n0089_inst_cy_137/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0089_inst_cy_137/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_137)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_137_848 (
    .IA(DLX_IDinst_IR_function_field_3_1),
    .IB(DLX_EXinst_Mcompar__n0089_inst_cy_136),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_73),
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_137/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0089_inst_cy_137/CYINIT_849  (
    .I(DLX_EXinst_Mcompar__n0089_inst_cy_135),
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_137/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_138_850 (
    .IA(DLX_IDinst_IR_function_field[4]),
    .IB(\DLX_EXinst_Mcompar__n0089_inst_cy_139/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_74),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_138)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_741.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_741 (
    .ADR0(DLX_IDinst_IR_function_field[4]),
    .ADR1(DLX_IDinst_reg_out_A[4]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_74)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_751.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_751 (
    .ADR0(\DLX_IDinst_Imm[5] ),
    .ADR1(DLX_IDinst_reg_out_A[5]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_75)
  );
  X_BUF \DLX_EXinst_Mcompar__n0089_inst_cy_139/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0089_inst_cy_139/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_139)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_139_851 (
    .IA(\DLX_IDinst_Imm[5] ),
    .IB(DLX_EXinst_Mcompar__n0089_inst_cy_138),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_75),
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_139/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0089_inst_cy_139/CYINIT_852  (
    .I(DLX_EXinst_Mcompar__n0089_inst_cy_137),
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_139/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_140_853 (
    .IA(\DLX_IDinst_Imm[6] ),
    .IB(\DLX_EXinst_Mcompar__n0089_inst_cy_141/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_76),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_140)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_761.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_761 (
    .ADR0(\DLX_IDinst_Imm[6] ),
    .ADR1(DLX_IDinst_reg_out_A[6]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_76)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_771.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_771 (
    .ADR0(\DLX_IDinst_Imm[7] ),
    .ADR1(DLX_IDinst_reg_out_A[7]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_77)
  );
  X_BUF \DLX_EXinst_Mcompar__n0089_inst_cy_141/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0089_inst_cy_141/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_141)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_141_854 (
    .IA(\DLX_IDinst_Imm[7] ),
    .IB(DLX_EXinst_Mcompar__n0089_inst_cy_140),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_77),
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_141/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0089_inst_cy_141/CYINIT_855  (
    .I(DLX_EXinst_Mcompar__n0089_inst_cy_139),
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_141/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_142_856 (
    .IA(\DLX_IDinst_Imm[8] ),
    .IB(\DLX_EXinst_Mcompar__n0089_inst_cy_143/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_78),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_142)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_781.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_781 (
    .ADR0(\DLX_IDinst_Imm[8] ),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[8]),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_78)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_791.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_791 (
    .ADR0(\DLX_IDinst_Imm[9] ),
    .ADR1(DLX_IDinst_reg_out_A[9]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_79)
  );
  X_BUF \DLX_EXinst_Mcompar__n0089_inst_cy_143/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0089_inst_cy_143/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_143)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_143_857 (
    .IA(\DLX_IDinst_Imm[9] ),
    .IB(DLX_EXinst_Mcompar__n0089_inst_cy_142),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_79),
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_143/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0089_inst_cy_143/CYINIT_858  (
    .I(DLX_EXinst_Mcompar__n0089_inst_cy_141),
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_143/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_144_859 (
    .IA(\DLX_IDinst_Imm[10] ),
    .IB(\DLX_EXinst_Mcompar__n0089_inst_cy_145/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_80),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_144)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_801.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_801 (
    .ADR0(\DLX_IDinst_Imm[10] ),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[10]),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_80)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_811.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_811 (
    .ADR0(\DLX_IDinst_Imm[11] ),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[11]),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_81)
  );
  X_BUF \DLX_EXinst_Mcompar__n0089_inst_cy_145/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0089_inst_cy_145/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_145)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_145_860 (
    .IA(\DLX_IDinst_Imm[11] ),
    .IB(DLX_EXinst_Mcompar__n0089_inst_cy_144),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_81),
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_145/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0089_inst_cy_145/CYINIT_861  (
    .I(DLX_EXinst_Mcompar__n0089_inst_cy_143),
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_145/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_146_862 (
    .IA(\DLX_IDinst_Imm[12] ),
    .IB(\DLX_EXinst_Mcompar__n0089_inst_cy_147/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_82),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_146)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_821.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_821 (
    .ADR0(\DLX_IDinst_Imm[12] ),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[12]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_82)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_831.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_831 (
    .ADR0(\DLX_IDinst_Imm[13] ),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[13]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_83)
  );
  X_BUF \DLX_EXinst_Mcompar__n0089_inst_cy_147/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0089_inst_cy_147/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_147)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_147_863 (
    .IA(\DLX_IDinst_Imm[13] ),
    .IB(DLX_EXinst_Mcompar__n0089_inst_cy_146),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_83),
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_147/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0089_inst_cy_147/CYINIT_864  (
    .I(DLX_EXinst_Mcompar__n0089_inst_cy_145),
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_147/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_148_865 (
    .IA(\DLX_IDinst_Imm[14] ),
    .IB(\DLX_EXinst_Mcompar__n0089_inst_cy_149/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_84),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_148)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_841.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_841 (
    .ADR0(\DLX_IDinst_Imm[14] ),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[14]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_84)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_851.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_851 (
    .ADR0(\DLX_IDinst_Imm[15] ),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[15]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_85)
  );
  X_BUF \DLX_EXinst_Mcompar__n0089_inst_cy_149/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0089_inst_cy_149/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_149)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_149_866 (
    .IA(\DLX_IDinst_Imm[15] ),
    .IB(DLX_EXinst_Mcompar__n0089_inst_cy_148),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_85),
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_149/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0089_inst_cy_149/CYINIT_867  (
    .I(DLX_EXinst_Mcompar__n0089_inst_cy_147),
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_149/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_150_868 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(\DLX_EXinst_Mcompar__n0089_inst_cy_151/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_86),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_150)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_861.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_861 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(DLX_IDinst_reg_out_A[16]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_86)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_871.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_871 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[17]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_87)
  );
  X_BUF \DLX_EXinst_Mcompar__n0089_inst_cy_151/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0089_inst_cy_151/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_151)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_151_869 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(DLX_EXinst_Mcompar__n0089_inst_cy_150),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_87),
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_151/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0089_inst_cy_151/CYINIT_870  (
    .I(DLX_EXinst_Mcompar__n0089_inst_cy_149),
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_151/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_152_871 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(\DLX_EXinst_Mcompar__n0089_inst_cy_153/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_88),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_152)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_881.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_881 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[18]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_88)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_891.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_891 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(DLX_IDinst_reg_out_A[19]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_89)
  );
  X_BUF \DLX_EXinst_Mcompar__n0089_inst_cy_153/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0089_inst_cy_153/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_153)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_153_872 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(DLX_EXinst_Mcompar__n0089_inst_cy_152),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_89),
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_153/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0089_inst_cy_153/CYINIT_873  (
    .I(DLX_EXinst_Mcompar__n0089_inst_cy_151),
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_153/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_154_874 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(\DLX_EXinst_Mcompar__n0089_inst_cy_155/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_90),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_154)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_901.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_901 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[20]),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_90)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_911.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_911 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(DLX_IDinst_reg_out_A[21]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_91)
  );
  X_BUF \DLX_EXinst_Mcompar__n0089_inst_cy_155/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0089_inst_cy_155/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_155)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_155_875 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(DLX_EXinst_Mcompar__n0089_inst_cy_154),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_91),
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_155/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0089_inst_cy_155/CYINIT_876  (
    .I(DLX_EXinst_Mcompar__n0089_inst_cy_153),
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_155/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_156_877 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(\DLX_EXinst_Mcompar__n0089_inst_cy_157/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_92),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_156)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_921.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_921 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[22]),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_92)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_931.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_931 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[23]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_93)
  );
  X_BUF \DLX_EXinst_Mcompar__n0089_inst_cy_157/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0089_inst_cy_157/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_157)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_157_878 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(DLX_EXinst_Mcompar__n0089_inst_cy_156),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_93),
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_157/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0089_inst_cy_157/CYINIT_879  (
    .I(DLX_EXinst_Mcompar__n0089_inst_cy_155),
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_157/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_158_880 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(\DLX_EXinst_Mcompar__n0089_inst_cy_159/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_94),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_158)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_941.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_941 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(DLX_IDinst_reg_out_A[24]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_94)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_951.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_951 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(DLX_IDinst_reg_out_A[25]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_95)
  );
  X_BUF \DLX_EXinst_Mcompar__n0089_inst_cy_159/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0089_inst_cy_159/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_159)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_159_881 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(DLX_EXinst_Mcompar__n0089_inst_cy_158),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_95),
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_159/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0089_inst_cy_159/CYINIT_882  (
    .I(DLX_EXinst_Mcompar__n0089_inst_cy_157),
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_159/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_160_883 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(\DLX_EXinst_Mcompar__n0089_inst_cy_161/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_96),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_160)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_961.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_961 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[26]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_96)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_971.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_971 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[27]),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_97)
  );
  X_BUF \DLX_EXinst_Mcompar__n0089_inst_cy_161/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0089_inst_cy_161/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_161)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_161_884 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(DLX_EXinst_Mcompar__n0089_inst_cy_160),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_97),
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_161/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0089_inst_cy_161/CYINIT_885  (
    .I(DLX_EXinst_Mcompar__n0089_inst_cy_159),
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_161/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_162_886 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(\DLX_EXinst_Mcompar__n0089_inst_cy_163/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_98),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_162)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_981.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_981 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[28]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_98)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_991.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_991 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(DLX_IDinst_reg_out_A[29]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_99)
  );
  X_BUF \DLX_EXinst_Mcompar__n0089_inst_cy_163/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0089_inst_cy_163/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_163)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_163_887 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(DLX_EXinst_Mcompar__n0089_inst_cy_162),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_99),
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_163/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0089_inst_cy_163/CYINIT_888  (
    .I(DLX_EXinst_Mcompar__n0089_inst_cy_161),
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_163/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_164_889 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(\CHOICE5806/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_100),
    .O(\CHOICE5806/CYMUXF )
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_1001.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_1001 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(DLX_IDinst_reg_out_A[30]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_100)
  );
  defparam \DLX_EXinst__n0006<31>319 .INIT = 16'h88A0;
  X_LUT4 \DLX_EXinst__n0006<31>319  (
    .ADR0(DLX_IDinst_IR_function_field[0]),
    .ADR1(DLX_IDinst_reg_out_A[28]),
    .ADR2(DLX_IDinst_reg_out_A[30]),
    .ADR3(DLX_IDinst_IR_function_field[1]),
    .O(\CHOICE5806/GROM )
  );
  X_BUF \CHOICE5806/XBUSED  (
    .I(\CHOICE5806/CYMUXF ),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_164)
  );
  X_BUF \CHOICE5806/YUSED  (
    .I(\CHOICE5806/GROM ),
    .O(CHOICE5806)
  );
  X_BUF \CHOICE5806/CYINIT_890  (
    .I(DLX_EXinst_Mcompar__n0089_inst_cy_163),
    .O(\CHOICE5806/CYINIT )
  );
  X_ZERO \vga_top_vga1_gridvcounter<0>/LOGIC_ZERO_891  (
    .O(\vga_top_vga1_gridvcounter<0>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_0_892 (
    .IA(GLOBAL_LOGIC1_0),
    .IB(\vga_top_vga1_gridvcounter<0>/LOGIC_ZERO ),
    .SEL(vga_top_vga1_gridvcounter_Madd__n0000_inst_lut2_0),
    .O(vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_0)
  );
  defparam vga_top_vga1_gridvcounter_Madd__n0000_inst_lut2_01.INIT = 16'h00FF;
  X_LUT4 vga_top_vga1_gridvcounter_Madd__n0000_inst_lut2_01 (
    .ADR0(GLOBAL_LOGIC1_0),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_gridvcounter[0]),
    .O(vga_top_vga1_gridvcounter_Madd__n0000_inst_lut2_0)
  );
  defparam \vga_top_vga1_gridvcounter<0>/G .INIT = 16'hCCCC;
  X_LUT4 \vga_top_vga1_gridvcounter<0>/G  (
    .ADR0(GLOBAL_LOGIC0_8),
    .ADR1(vga_top_vga1_gridvcounter[1]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\vga_top_vga1_gridvcounter<0>/GROM )
  );
  X_BUF \vga_top_vga1_gridvcounter<0>/COUTUSED  (
    .I(\vga_top_vga1_gridvcounter<0>/CYMUXG ),
    .O(vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_1)
  );
  X_MUX2 vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_1_893 (
    .IA(GLOBAL_LOGIC0_8),
    .IB(vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_0),
    .SEL(\vga_top_vga1_gridvcounter<0>/GROM ),
    .O(\vga_top_vga1_gridvcounter<0>/CYMUXG )
  );
  X_XOR2 vga_top_vga1_gridvcounter_Madd__n0000_inst_sum_1 (
    .I0(vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_0),
    .I1(\vga_top_vga1_gridvcounter<0>/GROM ),
    .O(vga_top_vga1_gridvcounter__n0000[1])
  );
  X_ZERO \vga_top_vga1_gridvcounter<2>/LOGIC_ZERO_894  (
    .O(\vga_top_vga1_gridvcounter<2>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_2_895 (
    .IA(\vga_top_vga1_gridvcounter<2>/LOGIC_ZERO ),
    .IB(\vga_top_vga1_gridvcounter<2>/CYINIT ),
    .SEL(\vga_top_vga1_gridvcounter<2>/FROM ),
    .O(vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_2)
  );
  X_XOR2 vga_top_vga1_gridvcounter_Madd__n0000_inst_sum_2 (
    .I0(\vga_top_vga1_gridvcounter<2>/CYINIT ),
    .I1(\vga_top_vga1_gridvcounter<2>/FROM ),
    .O(vga_top_vga1_gridvcounter__n0000[2])
  );
  defparam \vga_top_vga1_gridvcounter<2>/F .INIT = 16'hFF00;
  X_LUT4 \vga_top_vga1_gridvcounter<2>/F  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_gridvcounter[2]),
    .O(\vga_top_vga1_gridvcounter<2>/FROM )
  );
  defparam \vga_top_vga1_gridvcounter<2>/G .INIT = 16'hFF00;
  X_LUT4 \vga_top_vga1_gridvcounter<2>/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_gridvcounter[3]),
    .O(\vga_top_vga1_gridvcounter<2>/GROM )
  );
  X_BUF \vga_top_vga1_gridvcounter<2>/COUTUSED  (
    .I(\vga_top_vga1_gridvcounter<2>/CYMUXG ),
    .O(vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_3)
  );
  X_MUX2 vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_3_896 (
    .IA(\vga_top_vga1_gridvcounter<2>/LOGIC_ZERO ),
    .IB(vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_2),
    .SEL(\vga_top_vga1_gridvcounter<2>/GROM ),
    .O(\vga_top_vga1_gridvcounter<2>/CYMUXG )
  );
  X_XOR2 vga_top_vga1_gridvcounter_Madd__n0000_inst_sum_3 (
    .I0(vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_2),
    .I1(\vga_top_vga1_gridvcounter<2>/GROM ),
    .O(vga_top_vga1_gridvcounter__n0000[3])
  );
  X_BUF \vga_top_vga1_gridvcounter<2>/CYINIT_897  (
    .I(vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_1),
    .O(\vga_top_vga1_gridvcounter<2>/CYINIT )
  );
  X_ZERO \vga_top_vga1_gridvcounter<4>/LOGIC_ZERO_898  (
    .O(\vga_top_vga1_gridvcounter<4>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_4_899 (
    .IA(\vga_top_vga1_gridvcounter<4>/LOGIC_ZERO ),
    .IB(\vga_top_vga1_gridvcounter<4>/CYINIT ),
    .SEL(\vga_top_vga1_gridvcounter<4>/FROM ),
    .O(vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_4)
  );
  X_XOR2 vga_top_vga1_gridvcounter_Madd__n0000_inst_sum_4 (
    .I0(\vga_top_vga1_gridvcounter<4>/CYINIT ),
    .I1(\vga_top_vga1_gridvcounter<4>/FROM ),
    .O(vga_top_vga1_gridvcounter__n0000[4])
  );
  defparam \vga_top_vga1_gridvcounter<4>/F .INIT = 16'hFF00;
  X_LUT4 \vga_top_vga1_gridvcounter<4>/F  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_gridvcounter[4]),
    .O(\vga_top_vga1_gridvcounter<4>/FROM )
  );
  defparam \vga_top_vga1_gridvcounter<4>/G .INIT = 16'hAAAA;
  X_LUT4 \vga_top_vga1_gridvcounter<4>/G  (
    .ADR0(vga_top_vga1_gridvcounter[5]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\vga_top_vga1_gridvcounter<4>/GROM )
  );
  X_BUF \vga_top_vga1_gridvcounter<4>/COUTUSED  (
    .I(\vga_top_vga1_gridvcounter<4>/CYMUXG ),
    .O(vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_5)
  );
  X_MUX2 vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_5_900 (
    .IA(\vga_top_vga1_gridvcounter<4>/LOGIC_ZERO ),
    .IB(vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_4),
    .SEL(\vga_top_vga1_gridvcounter<4>/GROM ),
    .O(\vga_top_vga1_gridvcounter<4>/CYMUXG )
  );
  X_XOR2 vga_top_vga1_gridvcounter_Madd__n0000_inst_sum_5 (
    .I0(vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_4),
    .I1(\vga_top_vga1_gridvcounter<4>/GROM ),
    .O(vga_top_vga1_gridvcounter__n0000[5])
  );
  X_BUF \vga_top_vga1_gridvcounter<4>/CYINIT_901  (
    .I(vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_3),
    .O(\vga_top_vga1_gridvcounter<4>/CYINIT )
  );
  defparam DLX_EXinst_ALU_result_0_1_902.INIT = 1'b0;
  X_FF DLX_EXinst_ALU_result_0_1_902 (
    .I(\DM_addr_eff<0>/OD ),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DM_addr_eff<0>/OFF/RST ),
    .O(DLX_EXinst_ALU_result_0_1)
  );
  X_OR2 \DM_addr_eff<0>/OFF/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DM_addr_eff<0>/OFF/RST )
  );
  X_ZERO \vga_top_vga1_gridvcounter<6>/LOGIC_ZERO_903  (
    .O(\vga_top_vga1_gridvcounter<6>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_6_904 (
    .IA(\vga_top_vga1_gridvcounter<6>/LOGIC_ZERO ),
    .IB(\vga_top_vga1_gridvcounter<6>/CYINIT ),
    .SEL(\vga_top_vga1_gridvcounter<6>/FROM ),
    .O(vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_6)
  );
  X_XOR2 vga_top_vga1_gridvcounter_Madd__n0000_inst_sum_6 (
    .I0(\vga_top_vga1_gridvcounter<6>/CYINIT ),
    .I1(\vga_top_vga1_gridvcounter<6>/FROM ),
    .O(vga_top_vga1_gridvcounter__n0000[6])
  );
  defparam \vga_top_vga1_gridvcounter<6>/F .INIT = 16'hFF00;
  X_LUT4 \vga_top_vga1_gridvcounter<6>/F  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_gridvcounter[6]),
    .O(\vga_top_vga1_gridvcounter<6>/FROM )
  );
  defparam \vga_top_vga1_gridvcounter<6>/G .INIT = 16'hF0F0;
  X_LUT4 \vga_top_vga1_gridvcounter<6>/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_gridvcounter[7]),
    .ADR3(VCC),
    .O(\vga_top_vga1_gridvcounter<6>/GROM )
  );
  X_BUF \vga_top_vga1_gridvcounter<6>/COUTUSED  (
    .I(\vga_top_vga1_gridvcounter<6>/CYMUXG ),
    .O(vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_7)
  );
  X_MUX2 vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_7_905 (
    .IA(\vga_top_vga1_gridvcounter<6>/LOGIC_ZERO ),
    .IB(vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_6),
    .SEL(\vga_top_vga1_gridvcounter<6>/GROM ),
    .O(\vga_top_vga1_gridvcounter<6>/CYMUXG )
  );
  X_XOR2 vga_top_vga1_gridvcounter_Madd__n0000_inst_sum_7 (
    .I0(vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_6),
    .I1(\vga_top_vga1_gridvcounter<6>/GROM ),
    .O(vga_top_vga1_gridvcounter__n0000[7])
  );
  X_BUF \vga_top_vga1_gridvcounter<6>/CYINIT_906  (
    .I(vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_5),
    .O(\vga_top_vga1_gridvcounter<6>/CYINIT )
  );
  X_XOR2 vga_top_vga1_gridvcounter_Madd__n0000_inst_sum_8 (
    .I0(\vga_top_vga1_gridvcounter<8>/CYINIT ),
    .I1(\vga_top_vga1_gridvcounter<8>_rt ),
    .O(vga_top_vga1_gridvcounter__n0000[8])
  );
  defparam \vga_top_vga1_gridvcounter<8>_rt_907 .INIT = 16'hFF00;
  X_LUT4 \vga_top_vga1_gridvcounter<8>_rt_907  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_gridvcounter[8]),
    .O(\vga_top_vga1_gridvcounter<8>_rt )
  );
  X_BUF \vga_top_vga1_gridvcounter<8>/CYINIT_908  (
    .I(vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_7),
    .O(\vga_top_vga1_gridvcounter<8>/CYINIT )
  );
  X_ONE \vga_top_vga1_Mcompar__n0033_inst_cy_344/LOGIC_ONE_909  (
    .O(\vga_top_vga1_Mcompar__n0033_inst_cy_344/LOGIC_ONE )
  );
  X_ZERO \vga_top_vga1_Mcompar__n0033_inst_cy_344/LOGIC_ZERO_910  (
    .O(\vga_top_vga1_Mcompar__n0033_inst_cy_344/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0033_inst_cy_343_911 (
    .IA(\vga_top_vga1_Mcompar__n0033_inst_cy_344/LOGIC_ZERO ),
    .IB(\vga_top_vga1_Mcompar__n0033_inst_cy_344/LOGIC_ONE ),
    .SEL(vga_top_vga1_Mcompar__n0033_inst_lut1_4),
    .O(vga_top_vga1_Mcompar__n0033_inst_cy_343)
  );
  defparam vga_top_vga1_Mcompar__n0033_inst_lut1_41.INIT = 16'h00FF;
  X_LUT4 vga_top_vga1_Mcompar__n0033_inst_lut1_41 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[0]),
    .O(vga_top_vga1_Mcompar__n0033_inst_lut1_4)
  );
  defparam vga_top_vga1_Mcompar__n0033_inst_lut1_51.INIT = 16'h5555;
  X_LUT4 vga_top_vga1_Mcompar__n0033_inst_lut1_51 (
    .ADR0(vga_top_vga1_hcounter[0]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(vga_top_vga1_Mcompar__n0033_inst_lut1_5)
  );
  X_BUF \vga_top_vga1_Mcompar__n0033_inst_cy_344/COUTUSED  (
    .I(\vga_top_vga1_Mcompar__n0033_inst_cy_344/CYMUXG ),
    .O(vga_top_vga1_Mcompar__n0033_inst_cy_344)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0033_inst_cy_344_912 (
    .IA(\vga_top_vga1_Mcompar__n0033_inst_cy_344/LOGIC_ZERO ),
    .IB(vga_top_vga1_Mcompar__n0033_inst_cy_343),
    .SEL(vga_top_vga1_Mcompar__n0033_inst_lut1_5),
    .O(\vga_top_vga1_Mcompar__n0033_inst_cy_344/CYMUXG )
  );
  X_ONE \vga_top_vga1_Mcompar__n0033_inst_cy_346/LOGIC_ONE_913  (
    .O(\vga_top_vga1_Mcompar__n0033_inst_cy_346/LOGIC_ONE )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0033_inst_cy_345_914 (
    .IA(\vga_top_vga1_Mcompar__n0033_inst_cy_346/LOGIC_ONE ),
    .IB(\vga_top_vga1_Mcompar__n0033_inst_cy_346/CYINIT ),
    .SEL(vga_top_vga1_Mcompar__n0033_inst_lut2_269),
    .O(vga_top_vga1_Mcompar__n0033_inst_cy_345)
  );
  defparam vga_top_vga1_Mcompar__n0033_inst_lut2_2691.INIT = 16'hF000;
  X_LUT4 vga_top_vga1_Mcompar__n0033_inst_lut2_2691 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_hcounter[2]),
    .ADR3(vga_top_vga1_hcounter[1]),
    .O(vga_top_vga1_Mcompar__n0033_inst_lut2_269)
  );
  defparam vga_top_vga1_Mcompar__n0033_inst_lut2_2701.INIT = 16'hF000;
  X_LUT4 vga_top_vga1_Mcompar__n0033_inst_lut2_2701 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_hcounter[1]),
    .ADR3(vga_top_vga1_hcounter[2]),
    .O(vga_top_vga1_Mcompar__n0033_inst_lut2_270)
  );
  X_BUF \vga_top_vga1_Mcompar__n0033_inst_cy_346/COUTUSED  (
    .I(\vga_top_vga1_Mcompar__n0033_inst_cy_346/CYMUXG ),
    .O(vga_top_vga1_Mcompar__n0033_inst_cy_346)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0033_inst_cy_346_915 (
    .IA(\vga_top_vga1_Mcompar__n0033_inst_cy_346/LOGIC_ONE ),
    .IB(vga_top_vga1_Mcompar__n0033_inst_cy_345),
    .SEL(vga_top_vga1_Mcompar__n0033_inst_lut2_270),
    .O(\vga_top_vga1_Mcompar__n0033_inst_cy_346/CYMUXG )
  );
  X_BUF \vga_top_vga1_Mcompar__n0033_inst_cy_346/CYINIT_916  (
    .I(vga_top_vga1_Mcompar__n0033_inst_cy_344),
    .O(\vga_top_vga1_Mcompar__n0033_inst_cy_346/CYINIT )
  );
  X_ZERO \vga_top_vga1_Mcompar__n0033_inst_cy_348/LOGIC_ZERO_917  (
    .O(\vga_top_vga1_Mcompar__n0033_inst_cy_348/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0033_inst_cy_347_918 (
    .IA(\vga_top_vga1_Mcompar__n0033_inst_cy_348/LOGIC_ZERO ),
    .IB(\vga_top_vga1_Mcompar__n0033_inst_cy_348/CYINIT ),
    .SEL(vga_top_vga1_Mcompar__n0033_inst_lut3_110),
    .O(vga_top_vga1_Mcompar__n0033_inst_cy_347)
  );
  defparam vga_top_vga1_Mcompar__n0033_inst_lut3_1101.INIT = 16'h0005;
  X_LUT4 vga_top_vga1_Mcompar__n0033_inst_lut3_1101 (
    .ADR0(vga_top_vga1_hcounter[3]),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_hcounter[4]),
    .ADR3(vga_top_vga1_hcounter[5]),
    .O(vga_top_vga1_Mcompar__n0033_inst_lut3_110)
  );
  defparam vga_top_vga1_Mcompar__n0033_inst_lut3_1111.INIT = 16'h0011;
  X_LUT4 vga_top_vga1_Mcompar__n0033_inst_lut3_1111 (
    .ADR0(vga_top_vga1_hcounter[3]),
    .ADR1(vga_top_vga1_hcounter[5]),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[4]),
    .O(vga_top_vga1_Mcompar__n0033_inst_lut3_111)
  );
  X_BUF \vga_top_vga1_Mcompar__n0033_inst_cy_348/COUTUSED  (
    .I(\vga_top_vga1_Mcompar__n0033_inst_cy_348/CYMUXG ),
    .O(vga_top_vga1_Mcompar__n0033_inst_cy_348)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0033_inst_cy_348_919 (
    .IA(\vga_top_vga1_Mcompar__n0033_inst_cy_348/LOGIC_ZERO ),
    .IB(vga_top_vga1_Mcompar__n0033_inst_cy_347),
    .SEL(vga_top_vga1_Mcompar__n0033_inst_lut3_111),
    .O(\vga_top_vga1_Mcompar__n0033_inst_cy_348/CYMUXG )
  );
  X_BUF \vga_top_vga1_Mcompar__n0033_inst_cy_348/CYINIT_920  (
    .I(vga_top_vga1_Mcompar__n0033_inst_cy_346),
    .O(\vga_top_vga1_Mcompar__n0033_inst_cy_348/CYINIT )
  );
  X_ONE \vga_top_vga1_Mcompar__n0033_inst_cy_350/LOGIC_ONE_921  (
    .O(\vga_top_vga1_Mcompar__n0033_inst_cy_350/LOGIC_ONE )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0033_inst_cy_349_922 (
    .IA(\vga_top_vga1_Mcompar__n0033_inst_cy_350/LOGIC_ONE ),
    .IB(\vga_top_vga1_Mcompar__n0033_inst_cy_350/CYINIT ),
    .SEL(vga_top_vga1_Mcompar__n0033_inst_lut2_271),
    .O(vga_top_vga1_Mcompar__n0033_inst_cy_349)
  );
  defparam vga_top_vga1_Mcompar__n0033_inst_lut2_2711.INIT = 16'h8888;
  X_LUT4 vga_top_vga1_Mcompar__n0033_inst_lut2_2711 (
    .ADR0(vga_top_vga1_hcounter[6]),
    .ADR1(vga_top_vga1_hcounter[7]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(vga_top_vga1_Mcompar__n0033_inst_lut2_271)
  );
  defparam vga_top_vga1_Mcompar__n0033_inst_lut2_2721.INIT = 16'hCC00;
  X_LUT4 vga_top_vga1_Mcompar__n0033_inst_lut2_2721 (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_hcounter[7]),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[6]),
    .O(vga_top_vga1_Mcompar__n0033_inst_lut2_272)
  );
  X_BUF \vga_top_vga1_Mcompar__n0033_inst_cy_350/COUTUSED  (
    .I(\vga_top_vga1_Mcompar__n0033_inst_cy_350/CYMUXG ),
    .O(vga_top_vga1_Mcompar__n0033_inst_cy_350)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0033_inst_cy_350_923 (
    .IA(\vga_top_vga1_Mcompar__n0033_inst_cy_350/LOGIC_ONE ),
    .IB(vga_top_vga1_Mcompar__n0033_inst_cy_349),
    .SEL(vga_top_vga1_Mcompar__n0033_inst_lut2_272),
    .O(\vga_top_vga1_Mcompar__n0033_inst_cy_350/CYMUXG )
  );
  X_BUF \vga_top_vga1_Mcompar__n0033_inst_cy_350/CYINIT_924  (
    .I(vga_top_vga1_Mcompar__n0033_inst_cy_348),
    .O(\vga_top_vga1_Mcompar__n0033_inst_cy_350/CYINIT )
  );
  X_ZERO \vga_top_vga1_Mcompar__n0033_inst_cy_352/LOGIC_ZERO_925  (
    .O(\vga_top_vga1_Mcompar__n0033_inst_cy_352/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0033_inst_cy_351_926 (
    .IA(\vga_top_vga1_Mcompar__n0033_inst_cy_352/LOGIC_ZERO ),
    .IB(\vga_top_vga1_Mcompar__n0033_inst_cy_352/CYINIT ),
    .SEL(vga_top_vga1_Mcompar__n0033_inst_lut1_6),
    .O(vga_top_vga1_Mcompar__n0033_inst_cy_351)
  );
  defparam vga_top_vga1_Mcompar__n0033_inst_lut1_61.INIT = 16'h3333;
  X_LUT4 vga_top_vga1_Mcompar__n0033_inst_lut1_61 (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_hcounter[8]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(vga_top_vga1_Mcompar__n0033_inst_lut1_6)
  );
  defparam vga_top_vga1_Mcompar__n0033_inst_lut1_71.INIT = 16'h00FF;
  X_LUT4 vga_top_vga1_Mcompar__n0033_inst_lut1_71 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[8]),
    .O(vga_top_vga1_Mcompar__n0033_inst_lut1_7)
  );
  X_BUF \vga_top_vga1_Mcompar__n0033_inst_cy_352/COUTUSED  (
    .I(\vga_top_vga1_Mcompar__n0033_inst_cy_352/CYMUXG ),
    .O(vga_top_vga1_Mcompar__n0033_inst_cy_352)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0033_inst_cy_352_927 (
    .IA(\vga_top_vga1_Mcompar__n0033_inst_cy_352/LOGIC_ZERO ),
    .IB(vga_top_vga1_Mcompar__n0033_inst_cy_351),
    .SEL(vga_top_vga1_Mcompar__n0033_inst_lut1_7),
    .O(\vga_top_vga1_Mcompar__n0033_inst_cy_352/CYMUXG )
  );
  X_BUF \vga_top_vga1_Mcompar__n0033_inst_cy_352/CYINIT_928  (
    .I(vga_top_vga1_Mcompar__n0033_inst_cy_350),
    .O(\vga_top_vga1_Mcompar__n0033_inst_cy_352/CYINIT )
  );
  X_ONE \vga_top_vga1_Mcompar__n0033_inst_cy_354/LOGIC_ONE_929  (
    .O(\vga_top_vga1_Mcompar__n0033_inst_cy_354/LOGIC_ONE )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0033_inst_cy_353_930 (
    .IA(\vga_top_vga1_Mcompar__n0033_inst_cy_354/LOGIC_ONE ),
    .IB(\vga_top_vga1_Mcompar__n0033_inst_cy_354/CYINIT ),
    .SEL(\$SIG_7 ),
    .O(vga_top_vga1_Mcompar__n0033_inst_cy_353)
  );
  defparam \$BEL_7 .INIT = 16'hF0F0;
  X_LUT4 \$BEL_7  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_hcounter[9]),
    .ADR3(VCC),
    .O(\$SIG_7 )
  );
  defparam \$BEL_8 .INIT = 16'hAAAA;
  X_LUT4 \$BEL_8  (
    .ADR0(vga_top_vga1_hcounter[9]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\$SIG_8 )
  );
  X_BUF \vga_top_vga1_Mcompar__n0033_inst_cy_354/COUTUSED  (
    .I(\vga_top_vga1_Mcompar__n0033_inst_cy_354/CYMUXG ),
    .O(vga_top_vga1_Mcompar__n0033_inst_cy_354)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0033_inst_cy_354_931 (
    .IA(\vga_top_vga1_Mcompar__n0033_inst_cy_354/LOGIC_ONE ),
    .IB(vga_top_vga1_Mcompar__n0033_inst_cy_353),
    .SEL(\$SIG_8 ),
    .O(\vga_top_vga1_Mcompar__n0033_inst_cy_354/CYMUXG )
  );
  X_BUF \vga_top_vga1_Mcompar__n0033_inst_cy_354/CYINIT_932  (
    .I(vga_top_vga1_Mcompar__n0033_inst_cy_352),
    .O(\vga_top_vga1_Mcompar__n0033_inst_cy_354/CYINIT )
  );
  X_ZERO \vga_top_vga1__n0033/LOGIC_ZERO_933  (
    .O(\vga_top_vga1__n0033/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0033_inst_cy_355_934 (
    .IA(\vga_top_vga1__n0033/LOGIC_ZERO ),
    .IB(\vga_top_vga1__n0033/CYINIT ),
    .SEL(vga_top_vga1_Mcompar__n0033_inst_lut4_47),
    .O(vga_top_vga1_Mcompar__n0033_inst_cy_355)
  );
  defparam vga_top_vga1_Mcompar__n0033_inst_lut4_471.INIT = 16'h0001;
  X_LUT4 vga_top_vga1_Mcompar__n0033_inst_lut4_471 (
    .ADR0(vga_top_vga1_hcounter[10]),
    .ADR1(vga_top_vga1_hcounter[13]),
    .ADR2(vga_top_vga1_hcounter[12]),
    .ADR3(vga_top_vga1_hcounter[11]),
    .O(vga_top_vga1_Mcompar__n0033_inst_lut4_47)
  );
  defparam vga_top_vga1_Mcompar__n0033_inst_lut2_2731.INIT = 16'h0505;
  X_LUT4 vga_top_vga1_Mcompar__n0033_inst_lut2_2731 (
    .ADR0(vga_top_vga1_hcounter[15]),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_hcounter[14]),
    .ADR3(VCC),
    .O(vga_top_vga1_Mcompar__n0033_inst_lut2_273)
  );
  X_BUF \vga_top_vga1__n0033/COUTUSED  (
    .I(\vga_top_vga1__n0033/CYMUXG ),
    .O(vga_top_vga1__n0033)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0033_inst_cy_356 (
    .IA(\vga_top_vga1__n0033/LOGIC_ZERO ),
    .IB(vga_top_vga1_Mcompar__n0033_inst_cy_355),
    .SEL(vga_top_vga1_Mcompar__n0033_inst_lut2_273),
    .O(\vga_top_vga1__n0033/CYMUXG )
  );
  X_BUF \vga_top_vga1__n0033/CYINIT_935  (
    .I(vga_top_vga1_Mcompar__n0033_inst_cy_354),
    .O(\vga_top_vga1__n0033/CYINIT )
  );
  X_ONE \vga_top_vga1_Mcompar__n0034_inst_cy_332/LOGIC_ONE_936  (
    .O(\vga_top_vga1_Mcompar__n0034_inst_cy_332/LOGIC_ONE )
  );
  X_ZERO \vga_top_vga1_Mcompar__n0034_inst_cy_332/LOGIC_ZERO_937  (
    .O(\vga_top_vga1_Mcompar__n0034_inst_cy_332/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0034_inst_cy_331_938 (
    .IA(\vga_top_vga1_Mcompar__n0034_inst_cy_332/LOGIC_ZERO ),
    .IB(\vga_top_vga1_Mcompar__n0034_inst_cy_332/LOGIC_ONE ),
    .SEL(\$SIG_9 ),
    .O(vga_top_vga1_Mcompar__n0034_inst_cy_331)
  );
  defparam \$BEL_9 .INIT = 16'hCCCC;
  X_LUT4 \$BEL_9  (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_hcounter[2]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\$SIG_9 )
  );
  defparam \$BEL_10 .INIT = 16'hCCCC;
  X_LUT4 \$BEL_10  (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_hcounter[2]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\$SIG_10 )
  );
  X_BUF \vga_top_vga1_Mcompar__n0034_inst_cy_332/COUTUSED  (
    .I(\vga_top_vga1_Mcompar__n0034_inst_cy_332/CYMUXG ),
    .O(vga_top_vga1_Mcompar__n0034_inst_cy_332)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0034_inst_cy_332_939 (
    .IA(\vga_top_vga1_Mcompar__n0034_inst_cy_332/LOGIC_ZERO ),
    .IB(vga_top_vga1_Mcompar__n0034_inst_cy_331),
    .SEL(\$SIG_10 ),
    .O(\vga_top_vga1_Mcompar__n0034_inst_cy_332/CYMUXG )
  );
  defparam DLX_EXinst_ALU_result_1_1_940.INIT = 1'b0;
  X_FF DLX_EXinst_ALU_result_1_1_940 (
    .I(\DM_addr_eff<1>/OD ),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DM_addr_eff<1>/OFF/RST ),
    .O(DLX_EXinst_ALU_result_1_1)
  );
  X_OR2 \DM_addr_eff<1>/OFF/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DM_addr_eff<1>/OFF/RST )
  );
  X_ONE \vga_top_vga1_Mcompar__n0034_inst_cy_334/LOGIC_ONE_941  (
    .O(\vga_top_vga1_Mcompar__n0034_inst_cy_334/LOGIC_ONE )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0034_inst_cy_333_942 (
    .IA(\vga_top_vga1_Mcompar__n0034_inst_cy_334/LOGIC_ONE ),
    .IB(\vga_top_vga1_Mcompar__n0034_inst_cy_334/CYINIT ),
    .SEL(vga_top_vga1_Mcompar__n0034_inst_lut2_262),
    .O(vga_top_vga1_Mcompar__n0034_inst_cy_333)
  );
  defparam vga_top_vga1_Mcompar__n0034_inst_lut2_2621.INIT = 16'h0303;
  X_LUT4 vga_top_vga1_Mcompar__n0034_inst_lut2_2621 (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_hcounter[4]),
    .ADR2(vga_top_vga1_hcounter[3]),
    .ADR3(VCC),
    .O(vga_top_vga1_Mcompar__n0034_inst_lut2_262)
  );
  defparam vga_top_vga1_Mcompar__n0034_inst_lut2_2631.INIT = 16'h1111;
  X_LUT4 vga_top_vga1_Mcompar__n0034_inst_lut2_2631 (
    .ADR0(vga_top_vga1_hcounter[3]),
    .ADR1(vga_top_vga1_hcounter[4]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(vga_top_vga1_Mcompar__n0034_inst_lut2_263)
  );
  X_BUF \vga_top_vga1_Mcompar__n0034_inst_cy_334/COUTUSED  (
    .I(\vga_top_vga1_Mcompar__n0034_inst_cy_334/CYMUXG ),
    .O(vga_top_vga1_Mcompar__n0034_inst_cy_334)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0034_inst_cy_334_943 (
    .IA(\vga_top_vga1_Mcompar__n0034_inst_cy_334/LOGIC_ONE ),
    .IB(vga_top_vga1_Mcompar__n0034_inst_cy_333),
    .SEL(vga_top_vga1_Mcompar__n0034_inst_lut2_263),
    .O(\vga_top_vga1_Mcompar__n0034_inst_cy_334/CYMUXG )
  );
  X_BUF \vga_top_vga1_Mcompar__n0034_inst_cy_334/CYINIT_944  (
    .I(vga_top_vga1_Mcompar__n0034_inst_cy_332),
    .O(\vga_top_vga1_Mcompar__n0034_inst_cy_334/CYINIT )
  );
  X_ZERO \vga_top_vga1_Mcompar__n0034_inst_cy_336/LOGIC_ZERO_945  (
    .O(\vga_top_vga1_Mcompar__n0034_inst_cy_336/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0034_inst_cy_335_946 (
    .IA(\vga_top_vga1_Mcompar__n0034_inst_cy_336/LOGIC_ZERO ),
    .IB(\vga_top_vga1_Mcompar__n0034_inst_cy_336/CYINIT ),
    .SEL(\$SIG_11 ),
    .O(vga_top_vga1_Mcompar__n0034_inst_cy_335)
  );
  defparam \$BEL_11 .INIT = 16'hAAAA;
  X_LUT4 \$BEL_11  (
    .ADR0(vga_top_vga1_hcounter[5]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\$SIG_11 )
  );
  defparam \$BEL_12 .INIT = 16'hCCCC;
  X_LUT4 \$BEL_12  (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_hcounter[5]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\$SIG_12 )
  );
  X_BUF \vga_top_vga1_Mcompar__n0034_inst_cy_336/COUTUSED  (
    .I(\vga_top_vga1_Mcompar__n0034_inst_cy_336/CYMUXG ),
    .O(vga_top_vga1_Mcompar__n0034_inst_cy_336)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0034_inst_cy_336_947 (
    .IA(\vga_top_vga1_Mcompar__n0034_inst_cy_336/LOGIC_ZERO ),
    .IB(vga_top_vga1_Mcompar__n0034_inst_cy_335),
    .SEL(\$SIG_12 ),
    .O(\vga_top_vga1_Mcompar__n0034_inst_cy_336/CYMUXG )
  );
  X_BUF \vga_top_vga1_Mcompar__n0034_inst_cy_336/CYINIT_948  (
    .I(vga_top_vga1_Mcompar__n0034_inst_cy_334),
    .O(\vga_top_vga1_Mcompar__n0034_inst_cy_336/CYINIT )
  );
  X_ONE \vga_top_vga1_Mcompar__n0034_inst_cy_338/LOGIC_ONE_949  (
    .O(\vga_top_vga1_Mcompar__n0034_inst_cy_338/LOGIC_ONE )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0034_inst_cy_337_950 (
    .IA(\vga_top_vga1_Mcompar__n0034_inst_cy_338/LOGIC_ONE ),
    .IB(\vga_top_vga1_Mcompar__n0034_inst_cy_338/CYINIT ),
    .SEL(vga_top_vga1_Mcompar__n0034_inst_lut2_264),
    .O(vga_top_vga1_Mcompar__n0034_inst_cy_337)
  );
  defparam vga_top_vga1_Mcompar__n0034_inst_lut2_2641.INIT = 16'h0505;
  X_LUT4 vga_top_vga1_Mcompar__n0034_inst_lut2_2641 (
    .ADR0(vga_top_vga1_hcounter[7]),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_hcounter[6]),
    .ADR3(VCC),
    .O(vga_top_vga1_Mcompar__n0034_inst_lut2_264)
  );
  defparam vga_top_vga1_Mcompar__n0034_inst_lut2_2651.INIT = 16'h0303;
  X_LUT4 vga_top_vga1_Mcompar__n0034_inst_lut2_2651 (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_hcounter[7]),
    .ADR2(vga_top_vga1_hcounter[6]),
    .ADR3(VCC),
    .O(vga_top_vga1_Mcompar__n0034_inst_lut2_265)
  );
  X_BUF \vga_top_vga1_Mcompar__n0034_inst_cy_338/COUTUSED  (
    .I(\vga_top_vga1_Mcompar__n0034_inst_cy_338/CYMUXG ),
    .O(vga_top_vga1_Mcompar__n0034_inst_cy_338)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0034_inst_cy_338_951 (
    .IA(\vga_top_vga1_Mcompar__n0034_inst_cy_338/LOGIC_ONE ),
    .IB(vga_top_vga1_Mcompar__n0034_inst_cy_337),
    .SEL(vga_top_vga1_Mcompar__n0034_inst_lut2_265),
    .O(\vga_top_vga1_Mcompar__n0034_inst_cy_338/CYMUXG )
  );
  X_BUF \vga_top_vga1_Mcompar__n0034_inst_cy_338/CYINIT_952  (
    .I(vga_top_vga1_Mcompar__n0034_inst_cy_336),
    .O(\vga_top_vga1_Mcompar__n0034_inst_cy_338/CYINIT )
  );
  X_ZERO \vga_top_vga1_Mcompar__n0034_inst_cy_340/LOGIC_ZERO_953  (
    .O(\vga_top_vga1_Mcompar__n0034_inst_cy_340/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0034_inst_cy_339_954 (
    .IA(\vga_top_vga1_Mcompar__n0034_inst_cy_340/LOGIC_ZERO ),
    .IB(\vga_top_vga1_Mcompar__n0034_inst_cy_340/CYINIT ),
    .SEL(vga_top_vga1_Mcompar__n0034_inst_lut2_266),
    .O(vga_top_vga1_Mcompar__n0034_inst_cy_339)
  );
  defparam vga_top_vga1_Mcompar__n0034_inst_lut2_2661.INIT = 16'hC0C0;
  X_LUT4 vga_top_vga1_Mcompar__n0034_inst_lut2_2661 (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_hcounter[8]),
    .ADR2(vga_top_vga1_hcounter[9]),
    .ADR3(VCC),
    .O(vga_top_vga1_Mcompar__n0034_inst_lut2_266)
  );
  defparam vga_top_vga1_Mcompar__n0034_inst_lut2_2671.INIT = 16'hCC00;
  X_LUT4 vga_top_vga1_Mcompar__n0034_inst_lut2_2671 (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_hcounter[8]),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[9]),
    .O(vga_top_vga1_Mcompar__n0034_inst_lut2_267)
  );
  X_BUF \vga_top_vga1_Mcompar__n0034_inst_cy_340/COUTUSED  (
    .I(\vga_top_vga1_Mcompar__n0034_inst_cy_340/CYMUXG ),
    .O(vga_top_vga1_Mcompar__n0034_inst_cy_340)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0034_inst_cy_340_955 (
    .IA(\vga_top_vga1_Mcompar__n0034_inst_cy_340/LOGIC_ZERO ),
    .IB(vga_top_vga1_Mcompar__n0034_inst_cy_339),
    .SEL(vga_top_vga1_Mcompar__n0034_inst_lut2_267),
    .O(\vga_top_vga1_Mcompar__n0034_inst_cy_340/CYMUXG )
  );
  X_BUF \vga_top_vga1_Mcompar__n0034_inst_cy_340/CYINIT_956  (
    .I(vga_top_vga1_Mcompar__n0034_inst_cy_338),
    .O(\vga_top_vga1_Mcompar__n0034_inst_cy_340/CYINIT )
  );
  X_ONE \vga_top_vga1__n0034/LOGIC_ONE_957  (
    .O(\vga_top_vga1__n0034/LOGIC_ONE )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0034_inst_cy_341_958 (
    .IA(\vga_top_vga1__n0034/LOGIC_ONE ),
    .IB(\vga_top_vga1__n0034/CYINIT ),
    .SEL(vga_top_vga1_Mcompar__n0034_inst_lut4_46),
    .O(vga_top_vga1_Mcompar__n0034_inst_cy_341)
  );
  defparam vga_top_vga1_Mcompar__n0034_inst_lut4_461.INIT = 16'h0001;
  X_LUT4 vga_top_vga1_Mcompar__n0034_inst_lut4_461 (
    .ADR0(vga_top_vga1_hcounter[13]),
    .ADR1(vga_top_vga1_hcounter[12]),
    .ADR2(vga_top_vga1_hcounter[11]),
    .ADR3(vga_top_vga1_hcounter[10]),
    .O(vga_top_vga1_Mcompar__n0034_inst_lut4_46)
  );
  defparam vga_top_vga1_Mcompar__n0034_inst_lut2_2681.INIT = 16'h0303;
  X_LUT4 vga_top_vga1_Mcompar__n0034_inst_lut2_2681 (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_hcounter[15]),
    .ADR2(vga_top_vga1_hcounter[14]),
    .ADR3(VCC),
    .O(vga_top_vga1_Mcompar__n0034_inst_lut2_268)
  );
  X_BUF \vga_top_vga1__n0034/COUTUSED  (
    .I(\vga_top_vga1__n0034/CYMUXG ),
    .O(vga_top_vga1__n0034)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0034_inst_cy_342 (
    .IA(\vga_top_vga1__n0034/LOGIC_ONE ),
    .IB(vga_top_vga1_Mcompar__n0034_inst_cy_341),
    .SEL(vga_top_vga1_Mcompar__n0034_inst_lut2_268),
    .O(\vga_top_vga1__n0034/CYMUXG )
  );
  X_BUF \vga_top_vga1__n0034/CYINIT_959  (
    .I(vga_top_vga1_Mcompar__n0034_inst_cy_340),
    .O(\vga_top_vga1__n0034/CYINIT )
  );
  X_ONE \DLX_IDinst__n0128<0>/LOGIC_ONE_960  (
    .O(\DLX_IDinst__n0128<0>/LOGIC_ONE )
  );
  X_MUX2 DLX_IDinst_Msub__n0128_inst_cy_299_961 (
    .IA(DLX_IDinst_Madd__n0129_inst_lut2_198),
    .IB(\DLX_IDinst__n0128<0>/CYINIT ),
    .SEL(DLX_IDinst_Msub__n0128_inst_lut2_230),
    .O(DLX_IDinst_Msub__n0128_inst_cy_299)
  );
  X_XOR2 DLX_IDinst_Msub__n0128_inst_sum_134 (
    .I0(\DLX_IDinst__n0128<0>/CYINIT ),
    .I1(DLX_IDinst_Msub__n0128_inst_lut2_230),
    .O(\DLX_IDinst__n0128<0>/XORF )
  );
  defparam DLX_IDinst_Msub__n0128_inst_lut2_2301.INIT = 16'hC3C3;
  X_LUT4 DLX_IDinst_Msub__n0128_inst_lut2_2301 (
    .ADR0(DLX_IDinst_Madd__n0129_inst_lut2_198),
    .ADR1(DLX_IFinst_NPC[0]),
    .ADR2(DLX_IDinst_jtarget[0]),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0128_inst_lut2_230)
  );
  defparam DLX_IDinst_Msub__n0128_inst_lut2_2311.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0128_inst_lut2_2311 (
    .ADR0(DLX_IDinst__n0129[1]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0128_inst_lut2_231)
  );
  X_BUF \DLX_IDinst__n0128<0>/COUTUSED  (
    .I(\DLX_IDinst__n0128<0>/CYMUXG ),
    .O(DLX_IDinst_Msub__n0128_inst_cy_300)
  );
  X_BUF \DLX_IDinst__n0128<0>/XUSED  (
    .I(\DLX_IDinst__n0128<0>/XORF ),
    .O(DLX_IDinst__n0128[0])
  );
  X_BUF \DLX_IDinst__n0128<0>/YUSED  (
    .I(\DLX_IDinst__n0128<0>/XORG ),
    .O(DLX_IDinst__n0128[1])
  );
  X_MUX2 DLX_IDinst_Msub__n0128_inst_cy_300_962 (
    .IA(DLX_IDinst__n0129[1]),
    .IB(DLX_IDinst_Msub__n0128_inst_cy_299),
    .SEL(DLX_IDinst_Msub__n0128_inst_lut2_231),
    .O(\DLX_IDinst__n0128<0>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Msub__n0128_inst_sum_135 (
    .I0(DLX_IDinst_Msub__n0128_inst_cy_299),
    .I1(DLX_IDinst_Msub__n0128_inst_lut2_231),
    .O(\DLX_IDinst__n0128<0>/XORG )
  );
  X_BUF \DLX_IDinst__n0128<0>/CYINIT_963  (
    .I(\DLX_IDinst__n0128<0>/LOGIC_ONE ),
    .O(\DLX_IDinst__n0128<0>/CYINIT )
  );
  X_MUX2 DLX_IDinst_Msub__n0128_inst_cy_301_964 (
    .IA(GLOBAL_LOGIC0_9),
    .IB(\DLX_IDinst__n0128<2>/CYINIT ),
    .SEL(\DLX_IDinst__n0128<2>/FROM ),
    .O(DLX_IDinst_Msub__n0128_inst_cy_301)
  );
  X_XOR2 DLX_IDinst_Msub__n0128_inst_sum_136 (
    .I0(\DLX_IDinst__n0128<2>/CYINIT ),
    .I1(\DLX_IDinst__n0128<2>/FROM ),
    .O(\DLX_IDinst__n0128<2>/XORF )
  );
  defparam \DLX_IDinst__n0128<2>/F .INIT = 16'hFF00;
  X_LUT4 \DLX_IDinst__n0128<2>/F  (
    .ADR0(GLOBAL_LOGIC0_9),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst__n0129[2]),
    .O(\DLX_IDinst__n0128<2>/FROM )
  );
  defparam DLX_IDinst_Msub__n0128_inst_lut2_2331.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0128_inst_lut2_2331 (
    .ADR0(DLX_IDinst__n0129[3]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0128_inst_lut2_233)
  );
  X_BUF \DLX_IDinst__n0128<2>/COUTUSED  (
    .I(\DLX_IDinst__n0128<2>/CYMUXG ),
    .O(DLX_IDinst_Msub__n0128_inst_cy_302)
  );
  X_BUF \DLX_IDinst__n0128<2>/XUSED  (
    .I(\DLX_IDinst__n0128<2>/XORF ),
    .O(DLX_IDinst__n0128[2])
  );
  X_BUF \DLX_IDinst__n0128<2>/YUSED  (
    .I(\DLX_IDinst__n0128<2>/XORG ),
    .O(DLX_IDinst__n0128[3])
  );
  X_MUX2 DLX_IDinst_Msub__n0128_inst_cy_302_965 (
    .IA(DLX_IDinst__n0129[3]),
    .IB(DLX_IDinst_Msub__n0128_inst_cy_301),
    .SEL(DLX_IDinst_Msub__n0128_inst_lut2_233),
    .O(\DLX_IDinst__n0128<2>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Msub__n0128_inst_sum_137 (
    .I0(DLX_IDinst_Msub__n0128_inst_cy_301),
    .I1(DLX_IDinst_Msub__n0128_inst_lut2_233),
    .O(\DLX_IDinst__n0128<2>/XORG )
  );
  X_BUF \DLX_IDinst__n0128<2>/CYINIT_966  (
    .I(DLX_IDinst_Msub__n0128_inst_cy_300),
    .O(\DLX_IDinst__n0128<2>/CYINIT )
  );
  X_MUX2 DLX_IDinst_Msub__n0128_inst_cy_303_967 (
    .IA(DLX_IDinst__n0129[4]),
    .IB(\DLX_IDinst__n0128<4>/CYINIT ),
    .SEL(DLX_IDinst_Msub__n0128_inst_lut2_234),
    .O(DLX_IDinst_Msub__n0128_inst_cy_303)
  );
  X_XOR2 DLX_IDinst_Msub__n0128_inst_sum_138 (
    .I0(\DLX_IDinst__n0128<4>/CYINIT ),
    .I1(DLX_IDinst_Msub__n0128_inst_lut2_234),
    .O(\DLX_IDinst__n0128<4>/XORF )
  );
  defparam DLX_IDinst_Msub__n0128_inst_lut2_2341.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0128_inst_lut2_2341 (
    .ADR0(DLX_IDinst__n0129[4]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0128_inst_lut2_234)
  );
  defparam DLX_IDinst_Msub__n0128_inst_lut2_2351.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0128_inst_lut2_2351 (
    .ADR0(DLX_IDinst__n0129[5]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0128_inst_lut2_235)
  );
  X_BUF \DLX_IDinst__n0128<4>/COUTUSED  (
    .I(\DLX_IDinst__n0128<4>/CYMUXG ),
    .O(DLX_IDinst_Msub__n0128_inst_cy_304)
  );
  X_BUF \DLX_IDinst__n0128<4>/XUSED  (
    .I(\DLX_IDinst__n0128<4>/XORF ),
    .O(DLX_IDinst__n0128[4])
  );
  X_BUF \DLX_IDinst__n0128<4>/YUSED  (
    .I(\DLX_IDinst__n0128<4>/XORG ),
    .O(DLX_IDinst__n0128[5])
  );
  X_MUX2 DLX_IDinst_Msub__n0128_inst_cy_304_968 (
    .IA(DLX_IDinst__n0129[5]),
    .IB(DLX_IDinst_Msub__n0128_inst_cy_303),
    .SEL(DLX_IDinst_Msub__n0128_inst_lut2_235),
    .O(\DLX_IDinst__n0128<4>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Msub__n0128_inst_sum_139 (
    .I0(DLX_IDinst_Msub__n0128_inst_cy_303),
    .I1(DLX_IDinst_Msub__n0128_inst_lut2_235),
    .O(\DLX_IDinst__n0128<4>/XORG )
  );
  X_BUF \DLX_IDinst__n0128<4>/CYINIT_969  (
    .I(DLX_IDinst_Msub__n0128_inst_cy_302),
    .O(\DLX_IDinst__n0128<4>/CYINIT )
  );
  X_MUX2 DLX_IDinst_Msub__n0128_inst_cy_305_970 (
    .IA(DLX_IDinst__n0129[6]),
    .IB(\DLX_IDinst__n0128<6>/CYINIT ),
    .SEL(DLX_IDinst_Msub__n0128_inst_lut2_236),
    .O(DLX_IDinst_Msub__n0128_inst_cy_305)
  );
  X_XOR2 DLX_IDinst_Msub__n0128_inst_sum_140 (
    .I0(\DLX_IDinst__n0128<6>/CYINIT ),
    .I1(DLX_IDinst_Msub__n0128_inst_lut2_236),
    .O(\DLX_IDinst__n0128<6>/XORF )
  );
  defparam DLX_IDinst_Msub__n0128_inst_lut2_2361.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0128_inst_lut2_2361 (
    .ADR0(DLX_IDinst__n0129[6]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0128_inst_lut2_236)
  );
  defparam DLX_IDinst_Msub__n0128_inst_lut2_2371.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0128_inst_lut2_2371 (
    .ADR0(DLX_IDinst__n0129[7]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0128_inst_lut2_237)
  );
  X_BUF \DLX_IDinst__n0128<6>/COUTUSED  (
    .I(\DLX_IDinst__n0128<6>/CYMUXG ),
    .O(DLX_IDinst_Msub__n0128_inst_cy_306)
  );
  X_BUF \DLX_IDinst__n0128<6>/XUSED  (
    .I(\DLX_IDinst__n0128<6>/XORF ),
    .O(DLX_IDinst__n0128[6])
  );
  X_BUF \DLX_IDinst__n0128<6>/YUSED  (
    .I(\DLX_IDinst__n0128<6>/XORG ),
    .O(DLX_IDinst__n0128[7])
  );
  X_MUX2 DLX_IDinst_Msub__n0128_inst_cy_306_971 (
    .IA(DLX_IDinst__n0129[7]),
    .IB(DLX_IDinst_Msub__n0128_inst_cy_305),
    .SEL(DLX_IDinst_Msub__n0128_inst_lut2_237),
    .O(\DLX_IDinst__n0128<6>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Msub__n0128_inst_sum_141 (
    .I0(DLX_IDinst_Msub__n0128_inst_cy_305),
    .I1(DLX_IDinst_Msub__n0128_inst_lut2_237),
    .O(\DLX_IDinst__n0128<6>/XORG )
  );
  X_BUF \DLX_IDinst__n0128<6>/CYINIT_972  (
    .I(DLX_IDinst_Msub__n0128_inst_cy_304),
    .O(\DLX_IDinst__n0128<6>/CYINIT )
  );
  X_MUX2 DLX_IDinst_Msub__n0128_inst_cy_307_973 (
    .IA(DLX_IDinst__n0129[8]),
    .IB(\DLX_IDinst__n0128<8>/CYINIT ),
    .SEL(DLX_IDinst_Msub__n0128_inst_lut2_238),
    .O(DLX_IDinst_Msub__n0128_inst_cy_307)
  );
  X_XOR2 DLX_IDinst_Msub__n0128_inst_sum_142 (
    .I0(\DLX_IDinst__n0128<8>/CYINIT ),
    .I1(DLX_IDinst_Msub__n0128_inst_lut2_238),
    .O(\DLX_IDinst__n0128<8>/XORF )
  );
  defparam DLX_IDinst_Msub__n0128_inst_lut2_2381.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0128_inst_lut2_2381 (
    .ADR0(DLX_IDinst__n0129[8]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0128_inst_lut2_238)
  );
  defparam DLX_IDinst_Msub__n0128_inst_lut2_2391.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0128_inst_lut2_2391 (
    .ADR0(DLX_IDinst__n0129[9]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0128_inst_lut2_239)
  );
  X_BUF \DLX_IDinst__n0128<8>/COUTUSED  (
    .I(\DLX_IDinst__n0128<8>/CYMUXG ),
    .O(DLX_IDinst_Msub__n0128_inst_cy_308)
  );
  X_BUF \DLX_IDinst__n0128<8>/XUSED  (
    .I(\DLX_IDinst__n0128<8>/XORF ),
    .O(DLX_IDinst__n0128[8])
  );
  X_BUF \DLX_IDinst__n0128<8>/YUSED  (
    .I(\DLX_IDinst__n0128<8>/XORG ),
    .O(DLX_IDinst__n0128[9])
  );
  X_MUX2 DLX_IDinst_Msub__n0128_inst_cy_308_974 (
    .IA(DLX_IDinst__n0129[9]),
    .IB(DLX_IDinst_Msub__n0128_inst_cy_307),
    .SEL(DLX_IDinst_Msub__n0128_inst_lut2_239),
    .O(\DLX_IDinst__n0128<8>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Msub__n0128_inst_sum_143 (
    .I0(DLX_IDinst_Msub__n0128_inst_cy_307),
    .I1(DLX_IDinst_Msub__n0128_inst_lut2_239),
    .O(\DLX_IDinst__n0128<8>/XORG )
  );
  X_BUF \DLX_IDinst__n0128<8>/CYINIT_975  (
    .I(DLX_IDinst_Msub__n0128_inst_cy_306),
    .O(\DLX_IDinst__n0128<8>/CYINIT )
  );
  X_MUX2 DLX_IDinst_Msub__n0128_inst_cy_309_976 (
    .IA(DLX_IDinst__n0129[10]),
    .IB(\DLX_IDinst__n0128<10>/CYINIT ),
    .SEL(DLX_IDinst_Msub__n0128_inst_lut2_240),
    .O(DLX_IDinst_Msub__n0128_inst_cy_309)
  );
  X_XOR2 DLX_IDinst_Msub__n0128_inst_sum_144 (
    .I0(\DLX_IDinst__n0128<10>/CYINIT ),
    .I1(DLX_IDinst_Msub__n0128_inst_lut2_240),
    .O(\DLX_IDinst__n0128<10>/XORF )
  );
  defparam DLX_IDinst_Msub__n0128_inst_lut2_2401.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0128_inst_lut2_2401 (
    .ADR0(DLX_IDinst__n0129[10]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0128_inst_lut2_240)
  );
  defparam DLX_IDinst_Msub__n0128_inst_lut2_2411.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0128_inst_lut2_2411 (
    .ADR0(DLX_IDinst__n0129[11]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0128_inst_lut2_241)
  );
  X_BUF \DLX_IDinst__n0128<10>/COUTUSED  (
    .I(\DLX_IDinst__n0128<10>/CYMUXG ),
    .O(DLX_IDinst_Msub__n0128_inst_cy_310)
  );
  X_BUF \DLX_IDinst__n0128<10>/XUSED  (
    .I(\DLX_IDinst__n0128<10>/XORF ),
    .O(DLX_IDinst__n0128[10])
  );
  X_BUF \DLX_IDinst__n0128<10>/YUSED  (
    .I(\DLX_IDinst__n0128<10>/XORG ),
    .O(DLX_IDinst__n0128[11])
  );
  X_MUX2 DLX_IDinst_Msub__n0128_inst_cy_310_977 (
    .IA(DLX_IDinst__n0129[11]),
    .IB(DLX_IDinst_Msub__n0128_inst_cy_309),
    .SEL(DLX_IDinst_Msub__n0128_inst_lut2_241),
    .O(\DLX_IDinst__n0128<10>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Msub__n0128_inst_sum_145 (
    .I0(DLX_IDinst_Msub__n0128_inst_cy_309),
    .I1(DLX_IDinst_Msub__n0128_inst_lut2_241),
    .O(\DLX_IDinst__n0128<10>/XORG )
  );
  X_BUF \DLX_IDinst__n0128<10>/CYINIT_978  (
    .I(DLX_IDinst_Msub__n0128_inst_cy_308),
    .O(\DLX_IDinst__n0128<10>/CYINIT )
  );
  X_MUX2 DLX_IDinst_Msub__n0128_inst_cy_311_979 (
    .IA(DLX_IDinst__n0129[12]),
    .IB(\DLX_IDinst__n0128<12>/CYINIT ),
    .SEL(DLX_IDinst_Msub__n0128_inst_lut2_242),
    .O(DLX_IDinst_Msub__n0128_inst_cy_311)
  );
  X_XOR2 DLX_IDinst_Msub__n0128_inst_sum_146 (
    .I0(\DLX_IDinst__n0128<12>/CYINIT ),
    .I1(DLX_IDinst_Msub__n0128_inst_lut2_242),
    .O(\DLX_IDinst__n0128<12>/XORF )
  );
  defparam DLX_IDinst_Msub__n0128_inst_lut2_2421.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0128_inst_lut2_2421 (
    .ADR0(DLX_IDinst__n0129[12]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0128_inst_lut2_242)
  );
  defparam DLX_IDinst_Msub__n0128_inst_lut2_2431.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0128_inst_lut2_2431 (
    .ADR0(DLX_IDinst__n0129[13]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0128_inst_lut2_243)
  );
  X_BUF \DLX_IDinst__n0128<12>/COUTUSED  (
    .I(\DLX_IDinst__n0128<12>/CYMUXG ),
    .O(DLX_IDinst_Msub__n0128_inst_cy_312)
  );
  X_BUF \DLX_IDinst__n0128<12>/XUSED  (
    .I(\DLX_IDinst__n0128<12>/XORF ),
    .O(DLX_IDinst__n0128[12])
  );
  X_BUF \DLX_IDinst__n0128<12>/YUSED  (
    .I(\DLX_IDinst__n0128<12>/XORG ),
    .O(DLX_IDinst__n0128[13])
  );
  X_MUX2 DLX_IDinst_Msub__n0128_inst_cy_312_980 (
    .IA(DLX_IDinst__n0129[13]),
    .IB(DLX_IDinst_Msub__n0128_inst_cy_311),
    .SEL(DLX_IDinst_Msub__n0128_inst_lut2_243),
    .O(\DLX_IDinst__n0128<12>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Msub__n0128_inst_sum_147 (
    .I0(DLX_IDinst_Msub__n0128_inst_cy_311),
    .I1(DLX_IDinst_Msub__n0128_inst_lut2_243),
    .O(\DLX_IDinst__n0128<12>/XORG )
  );
  X_BUF \DLX_IDinst__n0128<12>/CYINIT_981  (
    .I(DLX_IDinst_Msub__n0128_inst_cy_310),
    .O(\DLX_IDinst__n0128<12>/CYINIT )
  );
  X_MUX2 DLX_IDinst_Msub__n0128_inst_cy_313_982 (
    .IA(DLX_IDinst__n0129[14]),
    .IB(\DLX_IDinst__n0128<14>/CYINIT ),
    .SEL(DLX_IDinst_Msub__n0128_inst_lut2_244),
    .O(DLX_IDinst_Msub__n0128_inst_cy_313)
  );
  X_XOR2 DLX_IDinst_Msub__n0128_inst_sum_148 (
    .I0(\DLX_IDinst__n0128<14>/CYINIT ),
    .I1(DLX_IDinst_Msub__n0128_inst_lut2_244),
    .O(\DLX_IDinst__n0128<14>/XORF )
  );
  defparam DLX_IDinst_Msub__n0128_inst_lut2_2441.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0128_inst_lut2_2441 (
    .ADR0(DLX_IDinst__n0129[14]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0128_inst_lut2_244)
  );
  defparam DLX_IDinst_Msub__n0128_inst_lut2_2451.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0128_inst_lut2_2451 (
    .ADR0(DLX_IDinst__n0129[15]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0128_inst_lut2_245)
  );
  X_BUF \DLX_IDinst__n0128<14>/COUTUSED  (
    .I(\DLX_IDinst__n0128<14>/CYMUXG ),
    .O(DLX_IDinst_Msub__n0128_inst_cy_314)
  );
  X_BUF \DLX_IDinst__n0128<14>/XUSED  (
    .I(\DLX_IDinst__n0128<14>/XORF ),
    .O(DLX_IDinst__n0128[14])
  );
  X_BUF \DLX_IDinst__n0128<14>/YUSED  (
    .I(\DLX_IDinst__n0128<14>/XORG ),
    .O(DLX_IDinst__n0128[15])
  );
  X_MUX2 DLX_IDinst_Msub__n0128_inst_cy_314_983 (
    .IA(DLX_IDinst__n0129[15]),
    .IB(DLX_IDinst_Msub__n0128_inst_cy_313),
    .SEL(DLX_IDinst_Msub__n0128_inst_lut2_245),
    .O(\DLX_IDinst__n0128<14>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Msub__n0128_inst_sum_149 (
    .I0(DLX_IDinst_Msub__n0128_inst_cy_313),
    .I1(DLX_IDinst_Msub__n0128_inst_lut2_245),
    .O(\DLX_IDinst__n0128<14>/XORG )
  );
  X_BUF \DLX_IDinst__n0128<14>/CYINIT_984  (
    .I(DLX_IDinst_Msub__n0128_inst_cy_312),
    .O(\DLX_IDinst__n0128<14>/CYINIT )
  );
  X_MUX2 DLX_IDinst_Msub__n0128_inst_cy_315_985 (
    .IA(DLX_IDinst__n0129[16]),
    .IB(\DLX_IDinst__n0128<16>/CYINIT ),
    .SEL(DLX_IDinst_Msub__n0128_inst_lut2_246),
    .O(DLX_IDinst_Msub__n0128_inst_cy_315)
  );
  X_XOR2 DLX_IDinst_Msub__n0128_inst_sum_150 (
    .I0(\DLX_IDinst__n0128<16>/CYINIT ),
    .I1(DLX_IDinst_Msub__n0128_inst_lut2_246),
    .O(\DLX_IDinst__n0128<16>/XORF )
  );
  defparam DLX_IDinst_Msub__n0128_inst_lut2_2461.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0128_inst_lut2_2461 (
    .ADR0(DLX_IDinst__n0129[16]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0128_inst_lut2_246)
  );
  defparam DLX_IDinst_Msub__n0128_inst_lut2_2471.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0128_inst_lut2_2471 (
    .ADR0(DLX_IDinst__n0129[17]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0128_inst_lut2_247)
  );
  X_BUF \DLX_IDinst__n0128<16>/COUTUSED  (
    .I(\DLX_IDinst__n0128<16>/CYMUXG ),
    .O(DLX_IDinst_Msub__n0128_inst_cy_316)
  );
  X_BUF \DLX_IDinst__n0128<16>/XUSED  (
    .I(\DLX_IDinst__n0128<16>/XORF ),
    .O(DLX_IDinst__n0128[16])
  );
  X_BUF \DLX_IDinst__n0128<16>/YUSED  (
    .I(\DLX_IDinst__n0128<16>/XORG ),
    .O(DLX_IDinst__n0128[17])
  );
  X_MUX2 DLX_IDinst_Msub__n0128_inst_cy_316_986 (
    .IA(DLX_IDinst__n0129[17]),
    .IB(DLX_IDinst_Msub__n0128_inst_cy_315),
    .SEL(DLX_IDinst_Msub__n0128_inst_lut2_247),
    .O(\DLX_IDinst__n0128<16>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Msub__n0128_inst_sum_151 (
    .I0(DLX_IDinst_Msub__n0128_inst_cy_315),
    .I1(DLX_IDinst_Msub__n0128_inst_lut2_247),
    .O(\DLX_IDinst__n0128<16>/XORG )
  );
  X_BUF \DLX_IDinst__n0128<16>/CYINIT_987  (
    .I(DLX_IDinst_Msub__n0128_inst_cy_314),
    .O(\DLX_IDinst__n0128<16>/CYINIT )
  );
  defparam DLX_EXinst_ALU_result_2_1_988.INIT = 1'b0;
  X_FF DLX_EXinst_ALU_result_2_1_988 (
    .I(\DM_addr_eff<2>/OD ),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DM_addr_eff<2>/OFF/RST ),
    .O(DLX_EXinst_ALU_result_2_1)
  );
  X_OR2 \DM_addr_eff<2>/OFF/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DM_addr_eff<2>/OFF/RST )
  );
  X_MUX2 DLX_IDinst_Msub__n0128_inst_cy_317_989 (
    .IA(DLX_IDinst__n0129[18]),
    .IB(\DLX_IDinst__n0128<18>/CYINIT ),
    .SEL(DLX_IDinst_Msub__n0128_inst_lut2_248),
    .O(DLX_IDinst_Msub__n0128_inst_cy_317)
  );
  X_XOR2 DLX_IDinst_Msub__n0128_inst_sum_152 (
    .I0(\DLX_IDinst__n0128<18>/CYINIT ),
    .I1(DLX_IDinst_Msub__n0128_inst_lut2_248),
    .O(\DLX_IDinst__n0128<18>/XORF )
  );
  defparam DLX_IDinst_Msub__n0128_inst_lut2_2481.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0128_inst_lut2_2481 (
    .ADR0(DLX_IDinst__n0129[18]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0128_inst_lut2_248)
  );
  defparam DLX_IDinst_Msub__n0128_inst_lut2_2491.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0128_inst_lut2_2491 (
    .ADR0(DLX_IDinst__n0129[19]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0128_inst_lut2_249)
  );
  X_BUF \DLX_IDinst__n0128<18>/COUTUSED  (
    .I(\DLX_IDinst__n0128<18>/CYMUXG ),
    .O(DLX_IDinst_Msub__n0128_inst_cy_318)
  );
  X_BUF \DLX_IDinst__n0128<18>/XUSED  (
    .I(\DLX_IDinst__n0128<18>/XORF ),
    .O(DLX_IDinst__n0128[18])
  );
  X_BUF \DLX_IDinst__n0128<18>/YUSED  (
    .I(\DLX_IDinst__n0128<18>/XORG ),
    .O(DLX_IDinst__n0128[19])
  );
  X_MUX2 DLX_IDinst_Msub__n0128_inst_cy_318_990 (
    .IA(DLX_IDinst__n0129[19]),
    .IB(DLX_IDinst_Msub__n0128_inst_cy_317),
    .SEL(DLX_IDinst_Msub__n0128_inst_lut2_249),
    .O(\DLX_IDinst__n0128<18>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Msub__n0128_inst_sum_153 (
    .I0(DLX_IDinst_Msub__n0128_inst_cy_317),
    .I1(DLX_IDinst_Msub__n0128_inst_lut2_249),
    .O(\DLX_IDinst__n0128<18>/XORG )
  );
  X_BUF \DLX_IDinst__n0128<18>/CYINIT_991  (
    .I(DLX_IDinst_Msub__n0128_inst_cy_316),
    .O(\DLX_IDinst__n0128<18>/CYINIT )
  );
  X_MUX2 DLX_IDinst_Msub__n0128_inst_cy_319_992 (
    .IA(DLX_IDinst__n0129[20]),
    .IB(\DLX_IDinst__n0128<20>/CYINIT ),
    .SEL(DLX_IDinst_Msub__n0128_inst_lut2_250),
    .O(DLX_IDinst_Msub__n0128_inst_cy_319)
  );
  X_XOR2 DLX_IDinst_Msub__n0128_inst_sum_154 (
    .I0(\DLX_IDinst__n0128<20>/CYINIT ),
    .I1(DLX_IDinst_Msub__n0128_inst_lut2_250),
    .O(\DLX_IDinst__n0128<20>/XORF )
  );
  defparam DLX_IDinst_Msub__n0128_inst_lut2_2501.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0128_inst_lut2_2501 (
    .ADR0(DLX_IDinst__n0129[20]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0128_inst_lut2_250)
  );
  defparam DLX_IDinst_Msub__n0128_inst_lut2_2511.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0128_inst_lut2_2511 (
    .ADR0(DLX_IDinst__n0129[21]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0128_inst_lut2_251)
  );
  X_BUF \DLX_IDinst__n0128<20>/COUTUSED  (
    .I(\DLX_IDinst__n0128<20>/CYMUXG ),
    .O(DLX_IDinst_Msub__n0128_inst_cy_320)
  );
  X_BUF \DLX_IDinst__n0128<20>/XUSED  (
    .I(\DLX_IDinst__n0128<20>/XORF ),
    .O(DLX_IDinst__n0128[20])
  );
  X_BUF \DLX_IDinst__n0128<20>/YUSED  (
    .I(\DLX_IDinst__n0128<20>/XORG ),
    .O(DLX_IDinst__n0128[21])
  );
  X_MUX2 DLX_IDinst_Msub__n0128_inst_cy_320_993 (
    .IA(DLX_IDinst__n0129[21]),
    .IB(DLX_IDinst_Msub__n0128_inst_cy_319),
    .SEL(DLX_IDinst_Msub__n0128_inst_lut2_251),
    .O(\DLX_IDinst__n0128<20>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Msub__n0128_inst_sum_155 (
    .I0(DLX_IDinst_Msub__n0128_inst_cy_319),
    .I1(DLX_IDinst_Msub__n0128_inst_lut2_251),
    .O(\DLX_IDinst__n0128<20>/XORG )
  );
  X_BUF \DLX_IDinst__n0128<20>/CYINIT_994  (
    .I(DLX_IDinst_Msub__n0128_inst_cy_318),
    .O(\DLX_IDinst__n0128<20>/CYINIT )
  );
  X_MUX2 DLX_IDinst_Msub__n0128_inst_cy_321_995 (
    .IA(DLX_IDinst__n0129[22]),
    .IB(\DLX_IDinst__n0128<22>/CYINIT ),
    .SEL(DLX_IDinst_Msub__n0128_inst_lut2_252),
    .O(DLX_IDinst_Msub__n0128_inst_cy_321)
  );
  X_XOR2 DLX_IDinst_Msub__n0128_inst_sum_156 (
    .I0(\DLX_IDinst__n0128<22>/CYINIT ),
    .I1(DLX_IDinst_Msub__n0128_inst_lut2_252),
    .O(\DLX_IDinst__n0128<22>/XORF )
  );
  defparam DLX_IDinst_Msub__n0128_inst_lut2_2521.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0128_inst_lut2_2521 (
    .ADR0(DLX_IDinst__n0129[22]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0128_inst_lut2_252)
  );
  defparam DLX_IDinst_Msub__n0128_inst_lut2_2531.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0128_inst_lut2_2531 (
    .ADR0(DLX_IDinst__n0129[23]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0128_inst_lut2_253)
  );
  X_BUF \DLX_IDinst__n0128<22>/COUTUSED  (
    .I(\DLX_IDinst__n0128<22>/CYMUXG ),
    .O(DLX_IDinst_Msub__n0128_inst_cy_322)
  );
  X_BUF \DLX_IDinst__n0128<22>/XUSED  (
    .I(\DLX_IDinst__n0128<22>/XORF ),
    .O(DLX_IDinst__n0128[22])
  );
  X_BUF \DLX_IDinst__n0128<22>/YUSED  (
    .I(\DLX_IDinst__n0128<22>/XORG ),
    .O(DLX_IDinst__n0128[23])
  );
  X_MUX2 DLX_IDinst_Msub__n0128_inst_cy_322_996 (
    .IA(DLX_IDinst__n0129[23]),
    .IB(DLX_IDinst_Msub__n0128_inst_cy_321),
    .SEL(DLX_IDinst_Msub__n0128_inst_lut2_253),
    .O(\DLX_IDinst__n0128<22>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Msub__n0128_inst_sum_157 (
    .I0(DLX_IDinst_Msub__n0128_inst_cy_321),
    .I1(DLX_IDinst_Msub__n0128_inst_lut2_253),
    .O(\DLX_IDinst__n0128<22>/XORG )
  );
  X_BUF \DLX_IDinst__n0128<22>/CYINIT_997  (
    .I(DLX_IDinst_Msub__n0128_inst_cy_320),
    .O(\DLX_IDinst__n0128<22>/CYINIT )
  );
  X_MUX2 DLX_IDinst_Msub__n0128_inst_cy_323_998 (
    .IA(DLX_IDinst__n0129[24]),
    .IB(\DLX_IDinst__n0128<24>/CYINIT ),
    .SEL(DLX_IDinst_Msub__n0128_inst_lut2_254),
    .O(DLX_IDinst_Msub__n0128_inst_cy_323)
  );
  X_XOR2 DLX_IDinst_Msub__n0128_inst_sum_158 (
    .I0(\DLX_IDinst__n0128<24>/CYINIT ),
    .I1(DLX_IDinst_Msub__n0128_inst_lut2_254),
    .O(\DLX_IDinst__n0128<24>/XORF )
  );
  defparam DLX_IDinst_Msub__n0128_inst_lut2_2541.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0128_inst_lut2_2541 (
    .ADR0(DLX_IDinst__n0129[24]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0128_inst_lut2_254)
  );
  defparam DLX_IDinst_Msub__n0128_inst_lut2_2551.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0128_inst_lut2_2551 (
    .ADR0(DLX_IDinst__n0129[25]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0128_inst_lut2_255)
  );
  X_BUF \DLX_IDinst__n0128<24>/COUTUSED  (
    .I(\DLX_IDinst__n0128<24>/CYMUXG ),
    .O(DLX_IDinst_Msub__n0128_inst_cy_324)
  );
  X_BUF \DLX_IDinst__n0128<24>/XUSED  (
    .I(\DLX_IDinst__n0128<24>/XORF ),
    .O(DLX_IDinst__n0128[24])
  );
  X_BUF \DLX_IDinst__n0128<24>/YUSED  (
    .I(\DLX_IDinst__n0128<24>/XORG ),
    .O(DLX_IDinst__n0128[25])
  );
  X_MUX2 DLX_IDinst_Msub__n0128_inst_cy_324_999 (
    .IA(DLX_IDinst__n0129[25]),
    .IB(DLX_IDinst_Msub__n0128_inst_cy_323),
    .SEL(DLX_IDinst_Msub__n0128_inst_lut2_255),
    .O(\DLX_IDinst__n0128<24>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Msub__n0128_inst_sum_159 (
    .I0(DLX_IDinst_Msub__n0128_inst_cy_323),
    .I1(DLX_IDinst_Msub__n0128_inst_lut2_255),
    .O(\DLX_IDinst__n0128<24>/XORG )
  );
  X_BUF \DLX_IDinst__n0128<24>/CYINIT_1000  (
    .I(DLX_IDinst_Msub__n0128_inst_cy_322),
    .O(\DLX_IDinst__n0128<24>/CYINIT )
  );
  X_MUX2 DLX_IDinst_Msub__n0128_inst_cy_325_1001 (
    .IA(DLX_IDinst__n0129[26]),
    .IB(\DLX_IDinst__n0128<26>/CYINIT ),
    .SEL(DLX_IDinst_Msub__n0128_inst_lut2_256),
    .O(DLX_IDinst_Msub__n0128_inst_cy_325)
  );
  X_XOR2 DLX_IDinst_Msub__n0128_inst_sum_160 (
    .I0(\DLX_IDinst__n0128<26>/CYINIT ),
    .I1(DLX_IDinst_Msub__n0128_inst_lut2_256),
    .O(\DLX_IDinst__n0128<26>/XORF )
  );
  defparam DLX_IDinst_Msub__n0128_inst_lut2_2561.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0128_inst_lut2_2561 (
    .ADR0(DLX_IDinst__n0129[26]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0128_inst_lut2_256)
  );
  defparam DLX_IDinst_Msub__n0128_inst_lut2_2571.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0128_inst_lut2_2571 (
    .ADR0(DLX_IDinst__n0129[27]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0128_inst_lut2_257)
  );
  X_BUF \DLX_IDinst__n0128<26>/COUTUSED  (
    .I(\DLX_IDinst__n0128<26>/CYMUXG ),
    .O(DLX_IDinst_Msub__n0128_inst_cy_326)
  );
  X_BUF \DLX_IDinst__n0128<26>/XUSED  (
    .I(\DLX_IDinst__n0128<26>/XORF ),
    .O(DLX_IDinst__n0128[26])
  );
  X_BUF \DLX_IDinst__n0128<26>/YUSED  (
    .I(\DLX_IDinst__n0128<26>/XORG ),
    .O(DLX_IDinst__n0128[27])
  );
  X_MUX2 DLX_IDinst_Msub__n0128_inst_cy_326_1002 (
    .IA(DLX_IDinst__n0129[27]),
    .IB(DLX_IDinst_Msub__n0128_inst_cy_325),
    .SEL(DLX_IDinst_Msub__n0128_inst_lut2_257),
    .O(\DLX_IDinst__n0128<26>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Msub__n0128_inst_sum_161 (
    .I0(DLX_IDinst_Msub__n0128_inst_cy_325),
    .I1(DLX_IDinst_Msub__n0128_inst_lut2_257),
    .O(\DLX_IDinst__n0128<26>/XORG )
  );
  X_BUF \DLX_IDinst__n0128<26>/CYINIT_1003  (
    .I(DLX_IDinst_Msub__n0128_inst_cy_324),
    .O(\DLX_IDinst__n0128<26>/CYINIT )
  );
  X_MUX2 DLX_IDinst_Msub__n0128_inst_cy_327_1004 (
    .IA(DLX_IDinst__n0129[28]),
    .IB(\DLX_IDinst__n0128<28>/CYINIT ),
    .SEL(DLX_IDinst_Msub__n0128_inst_lut2_258),
    .O(DLX_IDinst_Msub__n0128_inst_cy_327)
  );
  X_XOR2 DLX_IDinst_Msub__n0128_inst_sum_162 (
    .I0(\DLX_IDinst__n0128<28>/CYINIT ),
    .I1(DLX_IDinst_Msub__n0128_inst_lut2_258),
    .O(\DLX_IDinst__n0128<28>/XORF )
  );
  defparam DLX_IDinst_Msub__n0128_inst_lut2_2581.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0128_inst_lut2_2581 (
    .ADR0(DLX_IDinst__n0129[28]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0128_inst_lut2_258)
  );
  defparam DLX_IDinst_Msub__n0128_inst_lut2_2591.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0128_inst_lut2_2591 (
    .ADR0(DLX_IDinst__n0129[29]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0128_inst_lut2_259)
  );
  X_BUF \DLX_IDinst__n0128<28>/COUTUSED  (
    .I(\DLX_IDinst__n0128<28>/CYMUXG ),
    .O(DLX_IDinst_Msub__n0128_inst_cy_328)
  );
  X_BUF \DLX_IDinst__n0128<28>/XUSED  (
    .I(\DLX_IDinst__n0128<28>/XORF ),
    .O(DLX_IDinst__n0128[28])
  );
  X_BUF \DLX_IDinst__n0128<28>/YUSED  (
    .I(\DLX_IDinst__n0128<28>/XORG ),
    .O(DLX_IDinst__n0128[29])
  );
  X_MUX2 DLX_IDinst_Msub__n0128_inst_cy_328_1005 (
    .IA(DLX_IDinst__n0129[29]),
    .IB(DLX_IDinst_Msub__n0128_inst_cy_327),
    .SEL(DLX_IDinst_Msub__n0128_inst_lut2_259),
    .O(\DLX_IDinst__n0128<28>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Msub__n0128_inst_sum_163 (
    .I0(DLX_IDinst_Msub__n0128_inst_cy_327),
    .I1(DLX_IDinst_Msub__n0128_inst_lut2_259),
    .O(\DLX_IDinst__n0128<28>/XORG )
  );
  X_BUF \DLX_IDinst__n0128<28>/CYINIT_1006  (
    .I(DLX_IDinst_Msub__n0128_inst_cy_326),
    .O(\DLX_IDinst__n0128<28>/CYINIT )
  );
  X_MUX2 DLX_IDinst_Msub__n0128_inst_cy_329_1007 (
    .IA(DLX_IDinst__n0129[30]),
    .IB(\DLX_IDinst__n0128<30>/CYINIT ),
    .SEL(DLX_IDinst_Msub__n0128_inst_lut2_260),
    .O(DLX_IDinst_Msub__n0128_inst_cy_329)
  );
  X_XOR2 DLX_IDinst_Msub__n0128_inst_sum_164 (
    .I0(\DLX_IDinst__n0128<30>/CYINIT ),
    .I1(DLX_IDinst_Msub__n0128_inst_lut2_260),
    .O(\DLX_IDinst__n0128<30>/XORF )
  );
  defparam DLX_IDinst_Msub__n0128_inst_lut2_2601.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0128_inst_lut2_2601 (
    .ADR0(DLX_IDinst__n0129[30]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0128_inst_lut2_260)
  );
  defparam DLX_IDinst_Msub__n0128_inst_lut2_2611.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0128_inst_lut2_2611 (
    .ADR0(DLX_IDinst__n0129[31]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0128_inst_lut2_261)
  );
  X_BUF \DLX_IDinst__n0128<30>/XUSED  (
    .I(\DLX_IDinst__n0128<30>/XORF ),
    .O(DLX_IDinst__n0128[30])
  );
  X_BUF \DLX_IDinst__n0128<30>/YUSED  (
    .I(\DLX_IDinst__n0128<30>/XORG ),
    .O(DLX_IDinst__n0128[31])
  );
  X_XOR2 DLX_IDinst_Msub__n0128_inst_sum_165 (
    .I0(DLX_IDinst_Msub__n0128_inst_cy_329),
    .I1(DLX_IDinst_Msub__n0128_inst_lut2_261),
    .O(\DLX_IDinst__n0128<30>/XORG )
  );
  X_BUF \DLX_IDinst__n0128<30>/CYINIT_1008  (
    .I(DLX_IDinst_Msub__n0128_inst_cy_328),
    .O(\DLX_IDinst__n0128<30>/CYINIT )
  );
  X_ONE \DLX_EXinst_Mcompar__n0053_inst_cy_103/LOGIC_ONE_1009  (
    .O(\DLX_EXinst_Mcompar__n0053_inst_cy_103/LOGIC_ONE )
  );
  X_ZERO \DLX_EXinst_Mcompar__n0053_inst_cy_103/LOGIC_ZERO_1010  (
    .O(\DLX_EXinst_Mcompar__n0053_inst_cy_103/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0053_inst_cy_102_1011 (
    .IA(\DLX_EXinst_Mcompar__n0053_inst_cy_103/LOGIC_ZERO ),
    .IB(\DLX_EXinst_Mcompar__n0053_inst_cy_103/LOGIC_ONE ),
    .SEL(DLX_EXinst_Mcompar__n0053_inst_lut4_0),
    .O(DLX_EXinst_Mcompar__n0053_inst_cy_102)
  );
  defparam DLX_EXinst_Mcompar__n0053_inst_lut4_01.INIT = 16'h8241;
  X_LUT4 DLX_EXinst_Mcompar__n0053_inst_lut4_01 (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(DLX_IDinst_reg_out_A[0]),
    .ADR2(DLX_IDinst_reg_out_B[0]),
    .ADR3(DLX_IDinst_reg_out_A[1]),
    .O(DLX_EXinst_Mcompar__n0053_inst_lut4_0)
  );
  defparam DLX_EXinst_Mcompar__n0053_inst_lut4_16.INIT = 16'h8421;
  X_LUT4 DLX_EXinst_Mcompar__n0053_inst_lut4_16 (
    .ADR0(DLX_IDinst_reg_out_A[3]),
    .ADR1(DLX_IDinst_reg_out_A[2]),
    .ADR2(DLX_IDinst_reg_out_B_3_1),
    .ADR3(DLX_IDinst_reg_out_B_2_1),
    .O(DLX_EXinst_Mcompar__n0053_inst_lut4_1)
  );
  X_BUF \DLX_EXinst_Mcompar__n0053_inst_cy_103/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0053_inst_cy_103/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0053_inst_cy_103)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0053_inst_cy_103_1012 (
    .IA(\DLX_EXinst_Mcompar__n0053_inst_cy_103/LOGIC_ZERO ),
    .IB(DLX_EXinst_Mcompar__n0053_inst_cy_102),
    .SEL(DLX_EXinst_Mcompar__n0053_inst_lut4_1),
    .O(\DLX_EXinst_Mcompar__n0053_inst_cy_103/CYMUXG )
  );
  X_ZERO \DLX_EXinst_Mcompar__n0053_inst_cy_105/LOGIC_ZERO_1013  (
    .O(\DLX_EXinst_Mcompar__n0053_inst_cy_105/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0053_inst_cy_104_1014 (
    .IA(\DLX_EXinst_Mcompar__n0053_inst_cy_105/LOGIC_ZERO ),
    .IB(\DLX_EXinst_Mcompar__n0053_inst_cy_105/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0053_inst_lut4_2),
    .O(DLX_EXinst_Mcompar__n0053_inst_cy_104)
  );
  defparam DLX_EXinst_Mcompar__n0053_inst_lut4_21.INIT = 16'h8421;
  X_LUT4 DLX_EXinst_Mcompar__n0053_inst_lut4_21 (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(DLX_IDinst_reg_out_B[5]),
    .ADR2(DLX_IDinst_reg_out_A[4]),
    .ADR3(DLX_IDinst_reg_out_A[5]),
    .O(DLX_EXinst_Mcompar__n0053_inst_lut4_2)
  );
  defparam DLX_EXinst_Mcompar__n0053_inst_lut4_31.INIT = 16'h8241;
  X_LUT4 DLX_EXinst_Mcompar__n0053_inst_lut4_31 (
    .ADR0(DLX_IDinst_reg_out_A[6]),
    .ADR1(DLX_IDinst_reg_out_B[7]),
    .ADR2(DLX_IDinst_reg_out_A[7]),
    .ADR3(DLX_IDinst_reg_out_B[6]),
    .O(DLX_EXinst_Mcompar__n0053_inst_lut4_3)
  );
  X_BUF \DLX_EXinst_Mcompar__n0053_inst_cy_105/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0053_inst_cy_105/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0053_inst_cy_105)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0053_inst_cy_105_1015 (
    .IA(\DLX_EXinst_Mcompar__n0053_inst_cy_105/LOGIC_ZERO ),
    .IB(DLX_EXinst_Mcompar__n0053_inst_cy_104),
    .SEL(DLX_EXinst_Mcompar__n0053_inst_lut4_3),
    .O(\DLX_EXinst_Mcompar__n0053_inst_cy_105/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0053_inst_cy_105/CYINIT_1016  (
    .I(DLX_EXinst_Mcompar__n0053_inst_cy_103),
    .O(\DLX_EXinst_Mcompar__n0053_inst_cy_105/CYINIT )
  );
  X_ZERO \DLX_EXinst_Mcompar__n0053_inst_cy_107/LOGIC_ZERO_1017  (
    .O(\DLX_EXinst_Mcompar__n0053_inst_cy_107/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0053_inst_cy_106_1018 (
    .IA(\DLX_EXinst_Mcompar__n0053_inst_cy_107/LOGIC_ZERO ),
    .IB(\DLX_EXinst_Mcompar__n0053_inst_cy_107/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0053_inst_lut4_4),
    .O(DLX_EXinst_Mcompar__n0053_inst_cy_106)
  );
  defparam DLX_EXinst_Mcompar__n0053_inst_lut4_41.INIT = 16'h8241;
  X_LUT4 DLX_EXinst_Mcompar__n0053_inst_lut4_41 (
    .ADR0(DLX_IDinst_reg_out_A[9]),
    .ADR1(DLX_IDinst_reg_out_B[8]),
    .ADR2(DLX_IDinst_reg_out_A[8]),
    .ADR3(DLX_IDinst_reg_out_B[9]),
    .O(DLX_EXinst_Mcompar__n0053_inst_lut4_4)
  );
  defparam DLX_EXinst_Mcompar__n0053_inst_lut4_51.INIT = 16'h8241;
  X_LUT4 DLX_EXinst_Mcompar__n0053_inst_lut4_51 (
    .ADR0(DLX_IDinst_reg_out_A[10]),
    .ADR1(DLX_IDinst_reg_out_B[11]),
    .ADR2(DLX_IDinst_reg_out_A[11]),
    .ADR3(DLX_IDinst_reg_out_B[10]),
    .O(DLX_EXinst_Mcompar__n0053_inst_lut4_5)
  );
  X_BUF \DLX_EXinst_Mcompar__n0053_inst_cy_107/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0053_inst_cy_107/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0053_inst_cy_107)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0053_inst_cy_107_1019 (
    .IA(\DLX_EXinst_Mcompar__n0053_inst_cy_107/LOGIC_ZERO ),
    .IB(DLX_EXinst_Mcompar__n0053_inst_cy_106),
    .SEL(DLX_EXinst_Mcompar__n0053_inst_lut4_5),
    .O(\DLX_EXinst_Mcompar__n0053_inst_cy_107/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0053_inst_cy_107/CYINIT_1020  (
    .I(DLX_EXinst_Mcompar__n0053_inst_cy_105),
    .O(\DLX_EXinst_Mcompar__n0053_inst_cy_107/CYINIT )
  );
  X_ZERO \DLX_EXinst_Mcompar__n0053_inst_cy_109/LOGIC_ZERO_1021  (
    .O(\DLX_EXinst_Mcompar__n0053_inst_cy_109/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0053_inst_cy_108_1022 (
    .IA(\DLX_EXinst_Mcompar__n0053_inst_cy_109/LOGIC_ZERO ),
    .IB(\DLX_EXinst_Mcompar__n0053_inst_cy_109/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0053_inst_lut4_6),
    .O(DLX_EXinst_Mcompar__n0053_inst_cy_108)
  );
  defparam DLX_EXinst_Mcompar__n0053_inst_lut4_61.INIT = 16'h8421;
  X_LUT4 DLX_EXinst_Mcompar__n0053_inst_lut4_61 (
    .ADR0(DLX_IDinst_reg_out_B[13]),
    .ADR1(DLX_IDinst_reg_out_B[12]),
    .ADR2(DLX_IDinst_reg_out_A[13]),
    .ADR3(DLX_IDinst_reg_out_A[12]),
    .O(DLX_EXinst_Mcompar__n0053_inst_lut4_6)
  );
  defparam DLX_EXinst_Mcompar__n0053_inst_lut4_71.INIT = 16'h8421;
  X_LUT4 DLX_EXinst_Mcompar__n0053_inst_lut4_71 (
    .ADR0(DLX_IDinst_reg_out_B[15]),
    .ADR1(DLX_IDinst_reg_out_B[14]),
    .ADR2(DLX_IDinst_reg_out_A[15]),
    .ADR3(DLX_IDinst_reg_out_A[14]),
    .O(DLX_EXinst_Mcompar__n0053_inst_lut4_7)
  );
  X_BUF \DLX_EXinst_Mcompar__n0053_inst_cy_109/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0053_inst_cy_109/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0053_inst_cy_109)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0053_inst_cy_109_1023 (
    .IA(\DLX_EXinst_Mcompar__n0053_inst_cy_109/LOGIC_ZERO ),
    .IB(DLX_EXinst_Mcompar__n0053_inst_cy_108),
    .SEL(DLX_EXinst_Mcompar__n0053_inst_lut4_7),
    .O(\DLX_EXinst_Mcompar__n0053_inst_cy_109/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0053_inst_cy_109/CYINIT_1024  (
    .I(DLX_EXinst_Mcompar__n0053_inst_cy_107),
    .O(\DLX_EXinst_Mcompar__n0053_inst_cy_109/CYINIT )
  );
  X_ZERO \DLX_EXinst_Mcompar__n0053_inst_cy_111/LOGIC_ZERO_1025  (
    .O(\DLX_EXinst_Mcompar__n0053_inst_cy_111/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0053_inst_cy_110_1026 (
    .IA(\DLX_EXinst_Mcompar__n0053_inst_cy_111/LOGIC_ZERO ),
    .IB(\DLX_EXinst_Mcompar__n0053_inst_cy_111/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0053_inst_lut4_8),
    .O(DLX_EXinst_Mcompar__n0053_inst_cy_110)
  );
  defparam DLX_EXinst_Mcompar__n0053_inst_lut4_81.INIT = 16'h9009;
  X_LUT4 DLX_EXinst_Mcompar__n0053_inst_lut4_81 (
    .ADR0(DLX_IDinst_reg_out_B[16]),
    .ADR1(DLX_IDinst_reg_out_A[16]),
    .ADR2(DLX_IDinst_reg_out_B[17]),
    .ADR3(DLX_IDinst_reg_out_A[17]),
    .O(DLX_EXinst_Mcompar__n0053_inst_lut4_8)
  );
  defparam DLX_EXinst_Mcompar__n0053_inst_lut4_91.INIT = 16'h8241;
  X_LUT4 DLX_EXinst_Mcompar__n0053_inst_lut4_91 (
    .ADR0(DLX_IDinst_reg_out_A[18]),
    .ADR1(DLX_IDinst_reg_out_A[19]),
    .ADR2(DLX_IDinst_reg_out_B[19]),
    .ADR3(DLX_IDinst_reg_out_B[18]),
    .O(DLX_EXinst_Mcompar__n0053_inst_lut4_9)
  );
  X_BUF \DLX_EXinst_Mcompar__n0053_inst_cy_111/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0053_inst_cy_111/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0053_inst_cy_111)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0053_inst_cy_111_1027 (
    .IA(\DLX_EXinst_Mcompar__n0053_inst_cy_111/LOGIC_ZERO ),
    .IB(DLX_EXinst_Mcompar__n0053_inst_cy_110),
    .SEL(DLX_EXinst_Mcompar__n0053_inst_lut4_9),
    .O(\DLX_EXinst_Mcompar__n0053_inst_cy_111/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0053_inst_cy_111/CYINIT_1028  (
    .I(DLX_EXinst_Mcompar__n0053_inst_cy_109),
    .O(\DLX_EXinst_Mcompar__n0053_inst_cy_111/CYINIT )
  );
  X_ZERO \DLX_EXinst_Mcompar__n0053_inst_cy_113/LOGIC_ZERO_1029  (
    .O(\DLX_EXinst_Mcompar__n0053_inst_cy_113/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0053_inst_cy_112_1030 (
    .IA(\DLX_EXinst_Mcompar__n0053_inst_cy_113/LOGIC_ZERO ),
    .IB(\DLX_EXinst_Mcompar__n0053_inst_cy_113/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0053_inst_lut4_10),
    .O(DLX_EXinst_Mcompar__n0053_inst_cy_112)
  );
  defparam DLX_EXinst_Mcompar__n0053_inst_lut4_101.INIT = 16'h9009;
  X_LUT4 DLX_EXinst_Mcompar__n0053_inst_lut4_101 (
    .ADR0(DLX_IDinst_reg_out_B[20]),
    .ADR1(DLX_IDinst_reg_out_A[20]),
    .ADR2(DLX_IDinst_reg_out_A[21]),
    .ADR3(DLX_IDinst_reg_out_B[21]),
    .O(DLX_EXinst_Mcompar__n0053_inst_lut4_10)
  );
  defparam DLX_EXinst_Mcompar__n0053_inst_lut4_111.INIT = 16'h9009;
  X_LUT4 DLX_EXinst_Mcompar__n0053_inst_lut4_111 (
    .ADR0(DLX_IDinst_reg_out_A[23]),
    .ADR1(DLX_IDinst_reg_out_B[23]),
    .ADR2(DLX_IDinst_reg_out_B[22]),
    .ADR3(DLX_IDinst_reg_out_A[22]),
    .O(DLX_EXinst_Mcompar__n0053_inst_lut4_11)
  );
  X_BUF \DLX_EXinst_Mcompar__n0053_inst_cy_113/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0053_inst_cy_113/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0053_inst_cy_113)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0053_inst_cy_113_1031 (
    .IA(\DLX_EXinst_Mcompar__n0053_inst_cy_113/LOGIC_ZERO ),
    .IB(DLX_EXinst_Mcompar__n0053_inst_cy_112),
    .SEL(DLX_EXinst_Mcompar__n0053_inst_lut4_11),
    .O(\DLX_EXinst_Mcompar__n0053_inst_cy_113/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0053_inst_cy_113/CYINIT_1032  (
    .I(DLX_EXinst_Mcompar__n0053_inst_cy_111),
    .O(\DLX_EXinst_Mcompar__n0053_inst_cy_113/CYINIT )
  );
  X_ZERO \DLX_EXinst_Mcompar__n0053_inst_cy_115/LOGIC_ZERO_1033  (
    .O(\DLX_EXinst_Mcompar__n0053_inst_cy_115/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0053_inst_cy_114_1034 (
    .IA(\DLX_EXinst_Mcompar__n0053_inst_cy_115/LOGIC_ZERO ),
    .IB(\DLX_EXinst_Mcompar__n0053_inst_cy_115/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0053_inst_lut4_12),
    .O(DLX_EXinst_Mcompar__n0053_inst_cy_114)
  );
  defparam DLX_EXinst_Mcompar__n0053_inst_lut4_121.INIT = 16'h8241;
  X_LUT4 DLX_EXinst_Mcompar__n0053_inst_lut4_121 (
    .ADR0(DLX_IDinst_reg_out_B[24]),
    .ADR1(DLX_IDinst_reg_out_A[25]),
    .ADR2(DLX_IDinst_reg_out_B[25]),
    .ADR3(DLX_IDinst_reg_out_A[24]),
    .O(DLX_EXinst_Mcompar__n0053_inst_lut4_12)
  );
  defparam DLX_EXinst_Mcompar__n0053_inst_lut4_131.INIT = 16'h8421;
  X_LUT4 DLX_EXinst_Mcompar__n0053_inst_lut4_131 (
    .ADR0(DLX_IDinst_reg_out_A[27]),
    .ADR1(DLX_IDinst_reg_out_B[26]),
    .ADR2(DLX_IDinst_reg_out_B[27]),
    .ADR3(DLX_IDinst_reg_out_A[26]),
    .O(DLX_EXinst_Mcompar__n0053_inst_lut4_13)
  );
  X_BUF \DLX_EXinst_Mcompar__n0053_inst_cy_115/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0053_inst_cy_115/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0053_inst_cy_115)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0053_inst_cy_115_1035 (
    .IA(\DLX_EXinst_Mcompar__n0053_inst_cy_115/LOGIC_ZERO ),
    .IB(DLX_EXinst_Mcompar__n0053_inst_cy_114),
    .SEL(DLX_EXinst_Mcompar__n0053_inst_lut4_13),
    .O(\DLX_EXinst_Mcompar__n0053_inst_cy_115/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0053_inst_cy_115/CYINIT_1036  (
    .I(DLX_EXinst_Mcompar__n0053_inst_cy_113),
    .O(\DLX_EXinst_Mcompar__n0053_inst_cy_115/CYINIT )
  );
  X_ZERO \DLX_EXinst__n0053/LOGIC_ZERO_1037  (
    .O(\DLX_EXinst__n0053/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0053_inst_cy_116_1038 (
    .IA(\DLX_EXinst__n0053/LOGIC_ZERO ),
    .IB(\DLX_EXinst__n0053/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0053_inst_lut4_14),
    .O(DLX_EXinst_Mcompar__n0053_inst_cy_116)
  );
  defparam DLX_EXinst_Mcompar__n0053_inst_lut4_141.INIT = 16'h8241;
  X_LUT4 DLX_EXinst_Mcompar__n0053_inst_lut4_141 (
    .ADR0(DLX_IDinst_reg_out_B[28]),
    .ADR1(DLX_IDinst_reg_out_A[29]),
    .ADR2(DLX_IDinst_reg_out_B[29]),
    .ADR3(DLX_IDinst_reg_out_A[28]),
    .O(DLX_EXinst_Mcompar__n0053_inst_lut4_14)
  );
  defparam DLX_EXinst_Mcompar__n0053_inst_lut4_151.INIT = 16'h8421;
  X_LUT4 DLX_EXinst_Mcompar__n0053_inst_lut4_151 (
    .ADR0(DLX_IDinst_reg_out_B[31]),
    .ADR1(DLX_IDinst_reg_out_A[30]),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(DLX_IDinst_reg_out_B[30]),
    .O(DLX_EXinst_Mcompar__n0053_inst_lut4_15)
  );
  X_BUF \DLX_EXinst__n0053/COUTUSED  (
    .I(\DLX_EXinst__n0053/CYMUXG ),
    .O(DLX_EXinst__n0053)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0053_inst_cy_117 (
    .IA(\DLX_EXinst__n0053/LOGIC_ZERO ),
    .IB(DLX_EXinst_Mcompar__n0053_inst_cy_116),
    .SEL(DLX_EXinst_Mcompar__n0053_inst_lut4_15),
    .O(\DLX_EXinst__n0053/CYMUXG )
  );
  X_BUF \DLX_EXinst__n0053/CYINIT_1039  (
    .I(DLX_EXinst_Mcompar__n0053_inst_cy_115),
    .O(\DLX_EXinst__n0053/CYINIT )
  );
  X_ZERO \DLX_EXinst_Mcompar__n0061_inst_cy_199/LOGIC_ZERO_1040  (
    .O(\DLX_EXinst_Mcompar__n0061_inst_cy_199/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0061_inst_cy_198_1041 (
    .IA(DLX_IDinst_reg_out_A[0]),
    .IB(\DLX_EXinst_Mcompar__n0061_inst_cy_199/LOGIC_ZERO ),
    .SEL(DLX_EXinst_Mcompar__n0061_inst_lut2_134),
    .O(DLX_EXinst_Mcompar__n0061_inst_cy_198)
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_lut2_1341.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_lut2_1341 (
    .ADR0(DLX_IDinst_reg_out_A[0]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[0]),
    .O(DLX_EXinst_Mcompar__n0061_inst_lut2_134)
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_lut2_1351.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_lut2_1351 (
    .ADR0(DLX_IDinst_reg_out_A[1]),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0061_inst_lut2_135)
  );
  X_BUF \DLX_EXinst_Mcompar__n0061_inst_cy_199/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0061_inst_cy_199/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0061_inst_cy_199)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0061_inst_cy_199_1042 (
    .IA(DLX_IDinst_reg_out_A[1]),
    .IB(DLX_EXinst_Mcompar__n0061_inst_cy_198),
    .SEL(DLX_EXinst_Mcompar__n0061_inst_lut2_135),
    .O(\DLX_EXinst_Mcompar__n0061_inst_cy_199/CYMUXG )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0061_inst_cy_200_1043 (
    .IA(DLX_IDinst_reg_out_A[2]),
    .IB(\DLX_EXinst_Mcompar__n0061_inst_cy_201/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0061_inst_lut2_136),
    .O(DLX_EXinst_Mcompar__n0061_inst_cy_200)
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_lut2_1361.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_lut2_1361 (
    .ADR0(DLX_IDinst_reg_out_A[2]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B_2_1),
    .O(DLX_EXinst_Mcompar__n0061_inst_lut2_136)
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_lut2_1371.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_lut2_1371 (
    .ADR0(DLX_IDinst_reg_out_A[3]),
    .ADR1(DLX_IDinst_reg_out_B_3_1),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0061_inst_lut2_137)
  );
  X_BUF \DLX_EXinst_Mcompar__n0061_inst_cy_201/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0061_inst_cy_201/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0061_inst_cy_201)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0061_inst_cy_201_1044 (
    .IA(DLX_IDinst_reg_out_A[3]),
    .IB(DLX_EXinst_Mcompar__n0061_inst_cy_200),
    .SEL(DLX_EXinst_Mcompar__n0061_inst_lut2_137),
    .O(\DLX_EXinst_Mcompar__n0061_inst_cy_201/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0061_inst_cy_201/CYINIT_1045  (
    .I(DLX_EXinst_Mcompar__n0061_inst_cy_199),
    .O(\DLX_EXinst_Mcompar__n0061_inst_cy_201/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0061_inst_cy_202_1046 (
    .IA(DLX_IDinst_reg_out_A[4]),
    .IB(\DLX_EXinst_Mcompar__n0061_inst_cy_203/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0061_inst_lut2_138),
    .O(DLX_EXinst_Mcompar__n0061_inst_cy_202)
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_lut2_1381.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_lut2_1381 (
    .ADR0(DLX_IDinst_reg_out_A[4]),
    .ADR1(DLX_IDinst_reg_out_B[4]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0061_inst_lut2_138)
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_lut2_1391.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_lut2_1391 (
    .ADR0(DLX_IDinst_reg_out_A[5]),
    .ADR1(DLX_IDinst_reg_out_B[5]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0061_inst_lut2_139)
  );
  X_BUF \DLX_EXinst_Mcompar__n0061_inst_cy_203/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0061_inst_cy_203/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0061_inst_cy_203)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0061_inst_cy_203_1047 (
    .IA(DLX_IDinst_reg_out_A[5]),
    .IB(DLX_EXinst_Mcompar__n0061_inst_cy_202),
    .SEL(DLX_EXinst_Mcompar__n0061_inst_lut2_139),
    .O(\DLX_EXinst_Mcompar__n0061_inst_cy_203/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0061_inst_cy_203/CYINIT_1048  (
    .I(DLX_EXinst_Mcompar__n0061_inst_cy_201),
    .O(\DLX_EXinst_Mcompar__n0061_inst_cy_203/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0061_inst_cy_204_1049 (
    .IA(DLX_IDinst_reg_out_A[6]),
    .IB(\DLX_EXinst_Mcompar__n0061_inst_cy_205/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0061_inst_lut2_140),
    .O(DLX_EXinst_Mcompar__n0061_inst_cy_204)
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_lut2_1401.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_lut2_1401 (
    .ADR0(DLX_IDinst_reg_out_A[6]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[6]),
    .O(DLX_EXinst_Mcompar__n0061_inst_lut2_140)
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_lut2_1411.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_lut2_1411 (
    .ADR0(DLX_IDinst_reg_out_A[7]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[7]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0061_inst_lut2_141)
  );
  X_BUF \DLX_EXinst_Mcompar__n0061_inst_cy_205/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0061_inst_cy_205/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0061_inst_cy_205)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0061_inst_cy_205_1050 (
    .IA(DLX_IDinst_reg_out_A[7]),
    .IB(DLX_EXinst_Mcompar__n0061_inst_cy_204),
    .SEL(DLX_EXinst_Mcompar__n0061_inst_lut2_141),
    .O(\DLX_EXinst_Mcompar__n0061_inst_cy_205/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0061_inst_cy_205/CYINIT_1051  (
    .I(DLX_EXinst_Mcompar__n0061_inst_cy_203),
    .O(\DLX_EXinst_Mcompar__n0061_inst_cy_205/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0061_inst_cy_206_1052 (
    .IA(DLX_IDinst_reg_out_A[8]),
    .IB(\DLX_EXinst_Mcompar__n0061_inst_cy_207/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0061_inst_lut2_142),
    .O(DLX_EXinst_Mcompar__n0061_inst_cy_206)
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_lut2_1421.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_lut2_1421 (
    .ADR0(DLX_IDinst_reg_out_A[8]),
    .ADR1(DLX_IDinst_reg_out_B[8]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0061_inst_lut2_142)
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_lut2_1431.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_lut2_1431 (
    .ADR0(DLX_IDinst_reg_out_A[9]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[9]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0061_inst_lut2_143)
  );
  X_BUF \DLX_EXinst_Mcompar__n0061_inst_cy_207/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0061_inst_cy_207/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0061_inst_cy_207)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0061_inst_cy_207_1053 (
    .IA(DLX_IDinst_reg_out_A[9]),
    .IB(DLX_EXinst_Mcompar__n0061_inst_cy_206),
    .SEL(DLX_EXinst_Mcompar__n0061_inst_lut2_143),
    .O(\DLX_EXinst_Mcompar__n0061_inst_cy_207/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0061_inst_cy_207/CYINIT_1054  (
    .I(DLX_EXinst_Mcompar__n0061_inst_cy_205),
    .O(\DLX_EXinst_Mcompar__n0061_inst_cy_207/CYINIT )
  );
  defparam DLX_EXinst_ALU_result_3_1_1055.INIT = 1'b0;
  X_FF DLX_EXinst_ALU_result_3_1_1055 (
    .I(\DM_addr_eff<3>/OD ),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DM_addr_eff<3>/OFF/RST ),
    .O(DLX_EXinst_ALU_result_3_1)
  );
  X_OR2 \DM_addr_eff<3>/OFF/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DM_addr_eff<3>/OFF/RST )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0061_inst_cy_208_1056 (
    .IA(DLX_IDinst_reg_out_A[10]),
    .IB(\DLX_EXinst_Mcompar__n0061_inst_cy_209/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0061_inst_lut2_144),
    .O(DLX_EXinst_Mcompar__n0061_inst_cy_208)
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_lut2_1441.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_lut2_1441 (
    .ADR0(DLX_IDinst_reg_out_A[10]),
    .ADR1(DLX_IDinst_reg_out_B[10]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0061_inst_lut2_144)
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_lut2_1451.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_lut2_1451 (
    .ADR0(DLX_IDinst_reg_out_A[11]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[11]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0061_inst_lut2_145)
  );
  X_BUF \DLX_EXinst_Mcompar__n0061_inst_cy_209/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0061_inst_cy_209/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0061_inst_cy_209)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0061_inst_cy_209_1057 (
    .IA(DLX_IDinst_reg_out_A[11]),
    .IB(DLX_EXinst_Mcompar__n0061_inst_cy_208),
    .SEL(DLX_EXinst_Mcompar__n0061_inst_lut2_145),
    .O(\DLX_EXinst_Mcompar__n0061_inst_cy_209/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0061_inst_cy_209/CYINIT_1058  (
    .I(DLX_EXinst_Mcompar__n0061_inst_cy_207),
    .O(\DLX_EXinst_Mcompar__n0061_inst_cy_209/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0061_inst_cy_210_1059 (
    .IA(DLX_IDinst_reg_out_A[12]),
    .IB(\DLX_EXinst_Mcompar__n0061_inst_cy_211/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0061_inst_lut2_146),
    .O(DLX_EXinst_Mcompar__n0061_inst_cy_210)
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_lut2_1461.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_lut2_1461 (
    .ADR0(DLX_IDinst_reg_out_A[12]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[12]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0061_inst_lut2_146)
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_lut2_1471.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_lut2_1471 (
    .ADR0(DLX_IDinst_reg_out_A[13]),
    .ADR1(DLX_IDinst_reg_out_B[13]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0061_inst_lut2_147)
  );
  X_BUF \DLX_EXinst_Mcompar__n0061_inst_cy_211/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0061_inst_cy_211/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0061_inst_cy_211)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0061_inst_cy_211_1060 (
    .IA(DLX_IDinst_reg_out_A[13]),
    .IB(DLX_EXinst_Mcompar__n0061_inst_cy_210),
    .SEL(DLX_EXinst_Mcompar__n0061_inst_lut2_147),
    .O(\DLX_EXinst_Mcompar__n0061_inst_cy_211/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0061_inst_cy_211/CYINIT_1061  (
    .I(DLX_EXinst_Mcompar__n0061_inst_cy_209),
    .O(\DLX_EXinst_Mcompar__n0061_inst_cy_211/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_232_1062 (
    .IA(DLX_IDinst_reg_out_B_2_1),
    .IB(\DLX_EXinst_Mcompar__n0063_inst_cy_233/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_168),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_232)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_1681.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_1681 (
    .ADR0(DLX_IDinst_reg_out_B_2_1),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[2]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_168)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_1691.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_1691 (
    .ADR0(DLX_IDinst_reg_out_B_3_1),
    .ADR1(DLX_IDinst_reg_out_A[3]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_169)
  );
  X_BUF \DLX_EXinst_Mcompar__n0063_inst_cy_233/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0063_inst_cy_233/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_233)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_233_1063 (
    .IA(DLX_IDinst_reg_out_B_3_1),
    .IB(DLX_EXinst_Mcompar__n0063_inst_cy_232),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_169),
    .O(\DLX_EXinst_Mcompar__n0063_inst_cy_233/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0063_inst_cy_233/CYINIT_1064  (
    .I(DLX_EXinst_Mcompar__n0063_inst_cy_231),
    .O(\DLX_EXinst_Mcompar__n0063_inst_cy_233/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_234_1065 (
    .IA(DLX_IDinst_reg_out_B[4]),
    .IB(\DLX_EXinst_Mcompar__n0063_inst_cy_235/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_170),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_234)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_1701.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_1701 (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(DLX_IDinst_reg_out_A[4]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_170)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_1711.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_1711 (
    .ADR0(DLX_IDinst_reg_out_B[5]),
    .ADR1(DLX_IDinst_reg_out_A[5]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_171)
  );
  X_BUF \DLX_EXinst_Mcompar__n0063_inst_cy_235/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0063_inst_cy_235/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_235)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_235_1066 (
    .IA(DLX_IDinst_reg_out_B[5]),
    .IB(DLX_EXinst_Mcompar__n0063_inst_cy_234),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_171),
    .O(\DLX_EXinst_Mcompar__n0063_inst_cy_235/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0063_inst_cy_235/CYINIT_1067  (
    .I(DLX_EXinst_Mcompar__n0063_inst_cy_233),
    .O(\DLX_EXinst_Mcompar__n0063_inst_cy_235/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_236_1068 (
    .IA(DLX_IDinst_reg_out_B[6]),
    .IB(\DLX_EXinst_Mcompar__n0063_inst_cy_237/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_172),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_236)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_1721.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_1721 (
    .ADR0(DLX_IDinst_reg_out_B[6]),
    .ADR1(DLX_IDinst_reg_out_A[6]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_172)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_1731.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_1731 (
    .ADR0(DLX_IDinst_reg_out_B[7]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[7]),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_173)
  );
  X_BUF \DLX_EXinst_Mcompar__n0063_inst_cy_237/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0063_inst_cy_237/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_237)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_237_1069 (
    .IA(DLX_IDinst_reg_out_B[7]),
    .IB(DLX_EXinst_Mcompar__n0063_inst_cy_236),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_173),
    .O(\DLX_EXinst_Mcompar__n0063_inst_cy_237/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0063_inst_cy_237/CYINIT_1070  (
    .I(DLX_EXinst_Mcompar__n0063_inst_cy_235),
    .O(\DLX_EXinst_Mcompar__n0063_inst_cy_237/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_238_1071 (
    .IA(DLX_IDinst_reg_out_B[8]),
    .IB(\DLX_EXinst_Mcompar__n0063_inst_cy_239/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_174),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_238)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_1741.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_1741 (
    .ADR0(DLX_IDinst_reg_out_B[8]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[8]),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_174)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_1751.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_1751 (
    .ADR0(DLX_IDinst_reg_out_B[9]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[9]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_175)
  );
  X_BUF \DLX_EXinst_Mcompar__n0063_inst_cy_239/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0063_inst_cy_239/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_239)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_239_1072 (
    .IA(DLX_IDinst_reg_out_B[9]),
    .IB(DLX_EXinst_Mcompar__n0063_inst_cy_238),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_175),
    .O(\DLX_EXinst_Mcompar__n0063_inst_cy_239/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0063_inst_cy_239/CYINIT_1073  (
    .I(DLX_EXinst_Mcompar__n0063_inst_cy_237),
    .O(\DLX_EXinst_Mcompar__n0063_inst_cy_239/CYINIT )
  );
  defparam DLX_EXinst_ALU_result_5_1_1074.INIT = 1'b0;
  X_FF DLX_EXinst_ALU_result_5_1_1074 (
    .I(\DM_addr_eff<5>/OD ),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DM_addr_eff<5>/OFF/RST ),
    .O(DLX_EXinst_ALU_result_5_1)
  );
  X_OR2 \DM_addr_eff<5>/OFF/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DM_addr_eff<5>/OFF/RST )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_240_1075 (
    .IA(DLX_IDinst_reg_out_B[10]),
    .IB(\DLX_EXinst_Mcompar__n0063_inst_cy_241/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_176),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_240)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_1761.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_1761 (
    .ADR0(DLX_IDinst_reg_out_B[10]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[10]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_176)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_1771.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_1771 (
    .ADR0(DLX_IDinst_reg_out_B[11]),
    .ADR1(DLX_IDinst_reg_out_A[11]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_177)
  );
  X_BUF \DLX_EXinst_Mcompar__n0063_inst_cy_241/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0063_inst_cy_241/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_241)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_241_1076 (
    .IA(DLX_IDinst_reg_out_B[11]),
    .IB(DLX_EXinst_Mcompar__n0063_inst_cy_240),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_177),
    .O(\DLX_EXinst_Mcompar__n0063_inst_cy_241/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0063_inst_cy_241/CYINIT_1077  (
    .I(DLX_EXinst_Mcompar__n0063_inst_cy_239),
    .O(\DLX_EXinst_Mcompar__n0063_inst_cy_241/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_242_1078 (
    .IA(DLX_IDinst_reg_out_B[12]),
    .IB(\DLX_EXinst_Mcompar__n0063_inst_cy_243/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_178),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_242)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_1781.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_1781 (
    .ADR0(DLX_IDinst_reg_out_B[12]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[12]),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_178)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_1791.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_1791 (
    .ADR0(DLX_IDinst_reg_out_B[13]),
    .ADR1(DLX_IDinst_reg_out_A[13]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_179)
  );
  X_BUF \DLX_EXinst_Mcompar__n0063_inst_cy_243/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0063_inst_cy_243/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_243)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_243_1079 (
    .IA(DLX_IDinst_reg_out_B[13]),
    .IB(DLX_EXinst_Mcompar__n0063_inst_cy_242),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_179),
    .O(\DLX_EXinst_Mcompar__n0063_inst_cy_243/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0063_inst_cy_243/CYINIT_1080  (
    .I(DLX_EXinst_Mcompar__n0063_inst_cy_241),
    .O(\DLX_EXinst_Mcompar__n0063_inst_cy_243/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_244_1081 (
    .IA(DLX_IDinst_reg_out_B[14]),
    .IB(\DLX_EXinst_Mcompar__n0063_inst_cy_245/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_180),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_244)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_1801.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_1801 (
    .ADR0(DLX_IDinst_reg_out_B[14]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[14]),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_180)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_1811.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_1811 (
    .ADR0(DLX_IDinst_reg_out_B[15]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[15]),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_181)
  );
  X_BUF \DLX_EXinst_Mcompar__n0063_inst_cy_245/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0063_inst_cy_245/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_245)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_245_1082 (
    .IA(DLX_IDinst_reg_out_B[15]),
    .IB(DLX_EXinst_Mcompar__n0063_inst_cy_244),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_181),
    .O(\DLX_EXinst_Mcompar__n0063_inst_cy_245/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0063_inst_cy_245/CYINIT_1083  (
    .I(DLX_EXinst_Mcompar__n0063_inst_cy_243),
    .O(\DLX_EXinst_Mcompar__n0063_inst_cy_245/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_246_1084 (
    .IA(DLX_IDinst_reg_out_B[16]),
    .IB(\DLX_EXinst_Mcompar__n0063_inst_cy_247/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_182),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_246)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_1821.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_1821 (
    .ADR0(DLX_IDinst_reg_out_B[16]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[16]),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_182)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_1831.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_1831 (
    .ADR0(DLX_IDinst_reg_out_B[17]),
    .ADR1(DLX_IDinst_reg_out_A[17]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_183)
  );
  X_BUF \DLX_EXinst_Mcompar__n0063_inst_cy_247/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0063_inst_cy_247/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_247)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_247_1085 (
    .IA(DLX_IDinst_reg_out_B[17]),
    .IB(DLX_EXinst_Mcompar__n0063_inst_cy_246),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_183),
    .O(\DLX_EXinst_Mcompar__n0063_inst_cy_247/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0063_inst_cy_247/CYINIT_1086  (
    .I(DLX_EXinst_Mcompar__n0063_inst_cy_245),
    .O(\DLX_EXinst_Mcompar__n0063_inst_cy_247/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_248_1087 (
    .IA(DLX_IDinst_reg_out_B[18]),
    .IB(\DLX_EXinst_Mcompar__n0063_inst_cy_249/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_184),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_248)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_1841.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_1841 (
    .ADR0(DLX_IDinst_reg_out_B[18]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[18]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_184)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_1851.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_1851 (
    .ADR0(DLX_IDinst_reg_out_B[19]),
    .ADR1(DLX_IDinst_reg_out_A[19]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_185)
  );
  X_BUF \DLX_EXinst_Mcompar__n0063_inst_cy_249/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0063_inst_cy_249/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_249)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_249_1088 (
    .IA(DLX_IDinst_reg_out_B[19]),
    .IB(DLX_EXinst_Mcompar__n0063_inst_cy_248),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_185),
    .O(\DLX_EXinst_Mcompar__n0063_inst_cy_249/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0063_inst_cy_249/CYINIT_1089  (
    .I(DLX_EXinst_Mcompar__n0063_inst_cy_247),
    .O(\DLX_EXinst_Mcompar__n0063_inst_cy_249/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_250_1090 (
    .IA(DLX_IDinst_reg_out_B[20]),
    .IB(\DLX_EXinst_Mcompar__n0063_inst_cy_251/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_186),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_250)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_1861.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_1861 (
    .ADR0(DLX_IDinst_reg_out_B[20]),
    .ADR1(DLX_IDinst_reg_out_A[20]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_186)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_1871.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_1871 (
    .ADR0(DLX_IDinst_reg_out_B[21]),
    .ADR1(DLX_IDinst_reg_out_A[21]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_187)
  );
  X_BUF \DLX_EXinst_Mcompar__n0063_inst_cy_251/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0063_inst_cy_251/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_251)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_251_1091 (
    .IA(DLX_IDinst_reg_out_B[21]),
    .IB(DLX_EXinst_Mcompar__n0063_inst_cy_250),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_187),
    .O(\DLX_EXinst_Mcompar__n0063_inst_cy_251/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0063_inst_cy_251/CYINIT_1092  (
    .I(DLX_EXinst_Mcompar__n0063_inst_cy_249),
    .O(\DLX_EXinst_Mcompar__n0063_inst_cy_251/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_252_1093 (
    .IA(DLX_IDinst_reg_out_B[22]),
    .IB(\DLX_EXinst_Mcompar__n0063_inst_cy_253/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_188),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_252)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_1881.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_1881 (
    .ADR0(DLX_IDinst_reg_out_B[22]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[22]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_188)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_1891.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_1891 (
    .ADR0(DLX_IDinst_reg_out_B[23]),
    .ADR1(DLX_IDinst_reg_out_A[23]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_189)
  );
  X_BUF \DLX_EXinst_Mcompar__n0063_inst_cy_253/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0063_inst_cy_253/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_253)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_253_1094 (
    .IA(DLX_IDinst_reg_out_B[23]),
    .IB(DLX_EXinst_Mcompar__n0063_inst_cy_252),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_189),
    .O(\DLX_EXinst_Mcompar__n0063_inst_cy_253/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0063_inst_cy_253/CYINIT_1095  (
    .I(DLX_EXinst_Mcompar__n0063_inst_cy_251),
    .O(\DLX_EXinst_Mcompar__n0063_inst_cy_253/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_254_1096 (
    .IA(DLX_IDinst_reg_out_B[24]),
    .IB(\DLX_EXinst_Mcompar__n0063_inst_cy_255/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_190),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_254)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_1901.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_1901 (
    .ADR0(DLX_IDinst_reg_out_B[24]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[24]),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_190)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_1911.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_1911 (
    .ADR0(DLX_IDinst_reg_out_B[25]),
    .ADR1(DLX_IDinst_reg_out_A[25]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_191)
  );
  X_BUF \DLX_EXinst_Mcompar__n0063_inst_cy_255/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0063_inst_cy_255/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_255)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_255_1097 (
    .IA(DLX_IDinst_reg_out_B[25]),
    .IB(DLX_EXinst_Mcompar__n0063_inst_cy_254),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_191),
    .O(\DLX_EXinst_Mcompar__n0063_inst_cy_255/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0063_inst_cy_255/CYINIT_1098  (
    .I(DLX_EXinst_Mcompar__n0063_inst_cy_253),
    .O(\DLX_EXinst_Mcompar__n0063_inst_cy_255/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_256_1099 (
    .IA(DLX_IDinst_reg_out_B[26]),
    .IB(\DLX_EXinst_Mcompar__n0063_inst_cy_257/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_192),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_256)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_1921.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_1921 (
    .ADR0(DLX_IDinst_reg_out_B[26]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[26]),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_192)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_1931.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_1931 (
    .ADR0(DLX_IDinst_reg_out_B[27]),
    .ADR1(DLX_IDinst_reg_out_A[27]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_193)
  );
  X_BUF \DLX_EXinst_Mcompar__n0063_inst_cy_257/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0063_inst_cy_257/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_257)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_257_1100 (
    .IA(DLX_IDinst_reg_out_B[27]),
    .IB(DLX_EXinst_Mcompar__n0063_inst_cy_256),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_193),
    .O(\DLX_EXinst_Mcompar__n0063_inst_cy_257/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0063_inst_cy_257/CYINIT_1101  (
    .I(DLX_EXinst_Mcompar__n0063_inst_cy_255),
    .O(\DLX_EXinst_Mcompar__n0063_inst_cy_257/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_258_1102 (
    .IA(DLX_IDinst_reg_out_B[28]),
    .IB(\DLX_EXinst_Mcompar__n0063_inst_cy_259/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_194),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_258)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_1941.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_1941 (
    .ADR0(DLX_IDinst_reg_out_B[28]),
    .ADR1(DLX_IDinst_reg_out_A[28]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_194)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_1951.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_1951 (
    .ADR0(DLX_IDinst_reg_out_B[29]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[29]),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_195)
  );
  X_BUF \DLX_EXinst_Mcompar__n0063_inst_cy_259/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0063_inst_cy_259/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_259)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_259_1103 (
    .IA(DLX_IDinst_reg_out_B[29]),
    .IB(DLX_EXinst_Mcompar__n0063_inst_cy_258),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_195),
    .O(\DLX_EXinst_Mcompar__n0063_inst_cy_259/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0063_inst_cy_259/CYINIT_1104  (
    .I(DLX_EXinst_Mcompar__n0063_inst_cy_257),
    .O(\DLX_EXinst_Mcompar__n0063_inst_cy_259/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_260_1105 (
    .IA(DLX_IDinst_reg_out_B[30]),
    .IB(\CHOICE5291/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_196),
    .O(\CHOICE5291/CYMUXF )
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_1961.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_1961 (
    .ADR0(DLX_IDinst_reg_out_B[30]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[30]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_196)
  );
  defparam \DLX_EXinst__n0006<30>166 .INIT = 16'hCC50;
  X_LUT4 \DLX_EXinst__n0006<30>166  (
    .ADR0(DLX_EXinst_N63157),
    .ADR1(\DLX_EXinst_Mshift__n0025_Sh[22] ),
    .ADR2(DLX_IDinst_reg_out_A[30]),
    .ADR3(DLX_IDinst_reg_out_B[3]),
    .O(\CHOICE5291/GROM )
  );
  X_BUF \CHOICE5291/XBUSED  (
    .I(\CHOICE5291/CYMUXF ),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_260)
  );
  X_BUF \CHOICE5291/YUSED  (
    .I(\CHOICE5291/GROM ),
    .O(CHOICE5291)
  );
  X_BUF \CHOICE5291/CYINIT_1106  (
    .I(DLX_EXinst_Mcompar__n0063_inst_cy_259),
    .O(\CHOICE5291/CYINIT )
  );
  X_ZERO \vga_top_vga1_gridhcounter<0>/LOGIC_ZERO_1107  (
    .O(\vga_top_vga1_gridhcounter<0>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_0_1108 (
    .IA(GLOBAL_LOGIC1_1),
    .IB(\vga_top_vga1_gridhcounter<0>/LOGIC_ZERO ),
    .SEL(vga_top_vga1_gridhcounter_Madd__n0000_inst_lut2_0),
    .O(vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_0)
  );
  defparam vga_top_vga1_gridhcounter_Madd__n0000_inst_lut2_01.INIT = 16'h3333;
  X_LUT4 vga_top_vga1_gridhcounter_Madd__n0000_inst_lut2_01 (
    .ADR0(GLOBAL_LOGIC1_1),
    .ADR1(vga_top_vga1_gridhcounter[0]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(vga_top_vga1_gridhcounter_Madd__n0000_inst_lut2_0)
  );
  defparam \vga_top_vga1_gridhcounter<0>/G .INIT = 16'hF0F0;
  X_LUT4 \vga_top_vga1_gridhcounter<0>/G  (
    .ADR0(GLOBAL_LOGIC0_7),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_gridhcounter[1]),
    .ADR3(VCC),
    .O(\vga_top_vga1_gridhcounter<0>/GROM )
  );
  X_BUF \vga_top_vga1_gridhcounter<0>/COUTUSED  (
    .I(\vga_top_vga1_gridhcounter<0>/CYMUXG ),
    .O(vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_1)
  );
  X_MUX2 vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_1_1109 (
    .IA(GLOBAL_LOGIC0_7),
    .IB(vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_0),
    .SEL(\vga_top_vga1_gridhcounter<0>/GROM ),
    .O(\vga_top_vga1_gridhcounter<0>/CYMUXG )
  );
  X_XOR2 vga_top_vga1_gridhcounter_Madd__n0000_inst_sum_1 (
    .I0(vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_0),
    .I1(\vga_top_vga1_gridhcounter<0>/GROM ),
    .O(vga_top_vga1_gridhcounter__n0000[1])
  );
  X_ZERO \vga_top_vga1_gridhcounter<2>/LOGIC_ZERO_1110  (
    .O(\vga_top_vga1_gridhcounter<2>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_2_1111 (
    .IA(\vga_top_vga1_gridhcounter<2>/LOGIC_ZERO ),
    .IB(\vga_top_vga1_gridhcounter<2>/CYINIT ),
    .SEL(\vga_top_vga1_gridhcounter<2>/FROM ),
    .O(vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_2)
  );
  X_XOR2 vga_top_vga1_gridhcounter_Madd__n0000_inst_sum_2 (
    .I0(\vga_top_vga1_gridhcounter<2>/CYINIT ),
    .I1(\vga_top_vga1_gridhcounter<2>/FROM ),
    .O(vga_top_vga1_gridhcounter__n0000[2])
  );
  defparam \vga_top_vga1_gridhcounter<2>/F .INIT = 16'hAAAA;
  X_LUT4 \vga_top_vga1_gridhcounter<2>/F  (
    .ADR0(vga_top_vga1_gridhcounter[2]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\vga_top_vga1_gridhcounter<2>/FROM )
  );
  defparam \vga_top_vga1_gridhcounter<2>/G .INIT = 16'hCCCC;
  X_LUT4 \vga_top_vga1_gridhcounter<2>/G  (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_gridhcounter[3]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\vga_top_vga1_gridhcounter<2>/GROM )
  );
  X_BUF \vga_top_vga1_gridhcounter<2>/COUTUSED  (
    .I(\vga_top_vga1_gridhcounter<2>/CYMUXG ),
    .O(vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_3)
  );
  X_MUX2 vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_3_1112 (
    .IA(\vga_top_vga1_gridhcounter<2>/LOGIC_ZERO ),
    .IB(vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_2),
    .SEL(\vga_top_vga1_gridhcounter<2>/GROM ),
    .O(\vga_top_vga1_gridhcounter<2>/CYMUXG )
  );
  X_XOR2 vga_top_vga1_gridhcounter_Madd__n0000_inst_sum_3 (
    .I0(vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_2),
    .I1(\vga_top_vga1_gridhcounter<2>/GROM ),
    .O(vga_top_vga1_gridhcounter__n0000[3])
  );
  X_BUF \vga_top_vga1_gridhcounter<2>/CYINIT_1113  (
    .I(vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_1),
    .O(\vga_top_vga1_gridhcounter<2>/CYINIT )
  );
  X_ZERO \vga_top_vga1_gridhcounter<4>/LOGIC_ZERO_1114  (
    .O(\vga_top_vga1_gridhcounter<4>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_4_1115 (
    .IA(\vga_top_vga1_gridhcounter<4>/LOGIC_ZERO ),
    .IB(\vga_top_vga1_gridhcounter<4>/CYINIT ),
    .SEL(\vga_top_vga1_gridhcounter<4>/FROM ),
    .O(vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_4)
  );
  X_XOR2 vga_top_vga1_gridhcounter_Madd__n0000_inst_sum_4 (
    .I0(\vga_top_vga1_gridhcounter<4>/CYINIT ),
    .I1(\vga_top_vga1_gridhcounter<4>/FROM ),
    .O(vga_top_vga1_gridhcounter__n0000[4])
  );
  defparam \vga_top_vga1_gridhcounter<4>/F .INIT = 16'hAAAA;
  X_LUT4 \vga_top_vga1_gridhcounter<4>/F  (
    .ADR0(vga_top_vga1_gridhcounter[4]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\vga_top_vga1_gridhcounter<4>/FROM )
  );
  defparam \vga_top_vga1_gridhcounter<4>/G .INIT = 16'hAAAA;
  X_LUT4 \vga_top_vga1_gridhcounter<4>/G  (
    .ADR0(vga_top_vga1_gridhcounter[5]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\vga_top_vga1_gridhcounter<4>/GROM )
  );
  X_BUF \vga_top_vga1_gridhcounter<4>/COUTUSED  (
    .I(\vga_top_vga1_gridhcounter<4>/CYMUXG ),
    .O(vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_5)
  );
  X_MUX2 vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_5_1116 (
    .IA(\vga_top_vga1_gridhcounter<4>/LOGIC_ZERO ),
    .IB(vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_4),
    .SEL(\vga_top_vga1_gridhcounter<4>/GROM ),
    .O(\vga_top_vga1_gridhcounter<4>/CYMUXG )
  );
  X_XOR2 vga_top_vga1_gridhcounter_Madd__n0000_inst_sum_5 (
    .I0(vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_4),
    .I1(\vga_top_vga1_gridhcounter<4>/GROM ),
    .O(vga_top_vga1_gridhcounter__n0000[5])
  );
  X_BUF \vga_top_vga1_gridhcounter<4>/CYINIT_1117  (
    .I(vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_3),
    .O(\vga_top_vga1_gridhcounter<4>/CYINIT )
  );
  X_ZERO \vga_top_vga1_gridhcounter<6>/LOGIC_ZERO_1118  (
    .O(\vga_top_vga1_gridhcounter<6>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_6_1119 (
    .IA(\vga_top_vga1_gridhcounter<6>/LOGIC_ZERO ),
    .IB(\vga_top_vga1_gridhcounter<6>/CYINIT ),
    .SEL(\vga_top_vga1_gridhcounter<6>/FROM ),
    .O(vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_6)
  );
  X_XOR2 vga_top_vga1_gridhcounter_Madd__n0000_inst_sum_6 (
    .I0(\vga_top_vga1_gridhcounter<6>/CYINIT ),
    .I1(\vga_top_vga1_gridhcounter<6>/FROM ),
    .O(vga_top_vga1_gridhcounter__n0000[6])
  );
  defparam \vga_top_vga1_gridhcounter<6>/F .INIT = 16'hCCCC;
  X_LUT4 \vga_top_vga1_gridhcounter<6>/F  (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_gridhcounter[6]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\vga_top_vga1_gridhcounter<6>/FROM )
  );
  defparam \vga_top_vga1_gridhcounter<6>/G .INIT = 16'hFF00;
  X_LUT4 \vga_top_vga1_gridhcounter<6>/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_gridhcounter[7]),
    .O(\vga_top_vga1_gridhcounter<6>/GROM )
  );
  X_BUF \vga_top_vga1_gridhcounter<6>/COUTUSED  (
    .I(\vga_top_vga1_gridhcounter<6>/CYMUXG ),
    .O(vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_7)
  );
  X_MUX2 vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_7_1120 (
    .IA(\vga_top_vga1_gridhcounter<6>/LOGIC_ZERO ),
    .IB(vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_6),
    .SEL(\vga_top_vga1_gridhcounter<6>/GROM ),
    .O(\vga_top_vga1_gridhcounter<6>/CYMUXG )
  );
  X_XOR2 vga_top_vga1_gridhcounter_Madd__n0000_inst_sum_7 (
    .I0(vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_6),
    .I1(\vga_top_vga1_gridhcounter<6>/GROM ),
    .O(vga_top_vga1_gridhcounter__n0000[7])
  );
  X_BUF \vga_top_vga1_gridhcounter<6>/CYINIT_1121  (
    .I(vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_5),
    .O(\vga_top_vga1_gridhcounter<6>/CYINIT )
  );
  X_XOR2 vga_top_vga1_gridhcounter_Madd__n0000_inst_sum_8 (
    .I0(\vga_top_vga1_gridhcounter<8>/CYINIT ),
    .I1(\vga_top_vga1_gridhcounter<8>_rt ),
    .O(vga_top_vga1_gridhcounter__n0000[8])
  );
  defparam \vga_top_vga1_gridhcounter<8>_rt_1122 .INIT = 16'hCCCC;
  X_LUT4 \vga_top_vga1_gridhcounter<8>_rt_1122  (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_gridhcounter[8]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\vga_top_vga1_gridhcounter<8>_rt )
  );
  X_BUF \vga_top_vga1_gridhcounter<8>/CYINIT_1123  (
    .I(vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_7),
    .O(\vga_top_vga1_gridhcounter<8>/CYINIT )
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<1>1 .INIT = 16'hAAAC;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<1>1  (
    .ADR0(DLX_IDinst_current_IR[1]),
    .ADR1(DLX_IFinst_IR_latched[1]),
    .ADR2(DLX_IDinst_counter[1]),
    .ADR3(DLX_IDinst_counter[0]),
    .O(\DLX_IDinst_current_IR<1>/FROM )
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<0>1 .INIT = 16'hFE04;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<0>1  (
    .ADR0(DLX_IDinst_counter[1]),
    .ADR1(DLX_IFinst_IR_latched[0]),
    .ADR2(DLX_IDinst_counter[0]),
    .ADR3(DLX_IDinst_current_IR[0]),
    .O(\DLX_IDinst_current_IR<1>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<1>/XUSED  (
    .I(\DLX_IDinst_current_IR<1>/FROM ),
    .O(DLX_IDinst_jtarget[1])
  );
  X_BUF \DLX_IDinst_current_IR<1>/YUSED  (
    .I(\DLX_IDinst_current_IR<1>/GROM ),
    .O(DLX_IDinst_jtarget[0])
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<3>1 .INIT = 16'hFE04;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<3>1  (
    .ADR0(DLX_IDinst_counter[0]),
    .ADR1(DLX_IFinst_IR_latched[3]),
    .ADR2(DLX_IDinst_counter[1]),
    .ADR3(DLX_IDinst_current_IR[3]),
    .O(\DLX_IDinst_current_IR<3>/FROM )
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<2>1 .INIT = 16'hFE04;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<2>1  (
    .ADR0(DLX_IDinst_counter[1]),
    .ADR1(DLX_IFinst_IR_latched[2]),
    .ADR2(DLX_IDinst_counter[0]),
    .ADR3(DLX_IDinst_current_IR[2]),
    .O(\DLX_IDinst_current_IR<3>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<3>/XUSED  (
    .I(\DLX_IDinst_current_IR<3>/FROM ),
    .O(DLX_IDinst_jtarget[3])
  );
  X_BUF \DLX_IDinst_current_IR<3>/YUSED  (
    .I(\DLX_IDinst_current_IR<3>/GROM ),
    .O(DLX_IDinst_jtarget[2])
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<5>1 .INIT = 16'hFE04;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<5>1  (
    .ADR0(DLX_IDinst_counter[1]),
    .ADR1(DLX_IFinst_IR_latched[5]),
    .ADR2(DLX_IDinst_counter[0]),
    .ADR3(DLX_IDinst_current_IR[5]),
    .O(\DLX_IDinst_current_IR<5>/FROM )
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<4>1 .INIT = 16'hCCCA;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<4>1  (
    .ADR0(DLX_IFinst_IR_latched[4]),
    .ADR1(DLX_IDinst_current_IR[4]),
    .ADR2(DLX_IDinst_counter[1]),
    .ADR3(DLX_IDinst_counter[0]),
    .O(\DLX_IDinst_current_IR<5>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<5>/XUSED  (
    .I(\DLX_IDinst_current_IR<5>/FROM ),
    .O(DLX_IDinst_jtarget[5])
  );
  X_BUF \DLX_IDinst_current_IR<5>/YUSED  (
    .I(\DLX_IDinst_current_IR<5>/GROM ),
    .O(DLX_IDinst_jtarget[4])
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<7>1 .INIT = 16'hCCCA;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<7>1  (
    .ADR0(DLX_IFinst_IR_latched[7]),
    .ADR1(DLX_IDinst_current_IR[7]),
    .ADR2(DLX_IDinst_counter[1]),
    .ADR3(DLX_IDinst_counter[0]),
    .O(\DLX_IDinst_current_IR<7>/FROM )
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<6>1 .INIT = 16'hAAAC;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<6>1  (
    .ADR0(DLX_IDinst_current_IR[6]),
    .ADR1(DLX_IFinst_IR_latched[6]),
    .ADR2(DLX_IDinst_counter[0]),
    .ADR3(DLX_IDinst_counter[1]),
    .O(\DLX_IDinst_current_IR<7>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<7>/XUSED  (
    .I(\DLX_IDinst_current_IR<7>/FROM ),
    .O(DLX_IDinst_jtarget[7])
  );
  X_BUF \DLX_IDinst_current_IR<7>/YUSED  (
    .I(\DLX_IDinst_current_IR<7>/GROM ),
    .O(DLX_IDinst_jtarget[6])
  );
  defparam DLX_EXinst_ALU_result_6_1_1124.INIT = 1'b0;
  X_FF DLX_EXinst_ALU_result_6_1_1124 (
    .I(\DM_addr_eff<6>/OD ),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DM_addr_eff<6>/OFF/RST ),
    .O(DLX_EXinst_ALU_result_6_1)
  );
  X_OR2 \DM_addr_eff<6>/OFF/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DM_addr_eff<6>/OFF/RST )
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<9>1 .INIT = 16'hCCCA;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<9>1  (
    .ADR0(DLX_IFinst_IR_latched[9]),
    .ADR1(DLX_IDinst_current_IR[9]),
    .ADR2(DLX_IDinst_counter[0]),
    .ADR3(DLX_IDinst_counter[1]),
    .O(\DLX_IDinst_current_IR<9>/FROM )
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<8>1 .INIT = 16'hABA8;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<8>1  (
    .ADR0(DLX_IDinst_current_IR[8]),
    .ADR1(DLX_IDinst_counter[0]),
    .ADR2(DLX_IDinst_counter[1]),
    .ADR3(DLX_IFinst_IR_latched[8]),
    .O(\DLX_IDinst_current_IR<9>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<9>/XUSED  (
    .I(\DLX_IDinst_current_IR<9>/FROM ),
    .O(DLX_IDinst_jtarget[9])
  );
  X_BUF \DLX_IDinst_current_IR<9>/YUSED  (
    .I(\DLX_IDinst_current_IR<9>/GROM ),
    .O(DLX_IDinst_jtarget[8])
  );
  defparam \DLX_IDinst_slot_num_FFd2-In10 .INIT = 16'hBBBA;
  X_LUT4 \DLX_IDinst_slot_num_FFd2-In10  (
    .ADR0(DLX_IDinst_slot_num_FFd2),
    .ADR1(DLX_IDinst_delay_slot),
    .ADR2(DLX_IDinst_slot_num_FFd3),
    .ADR3(DLX_IDinst_slot_num_FFd1),
    .O(\DLX_IDinst_slot_num_FFd1/FROM )
  );
  defparam \DLX_IDinst_slot_num_FFd1-In1 .INIT = 16'h0800;
  X_LUT4 \DLX_IDinst_slot_num_FFd1-In1  (
    .ADR0(N109741),
    .ADR1(DLX_IDinst_delay_slot),
    .ADR2(DLX_IDinst_N70570),
    .ADR3(DLX_IDinst_slot_num_FFd2),
    .O(\DLX_IDinst_slot_num_FFd1-In )
  );
  X_BUF \DLX_IDinst_slot_num_FFd1/XUSED  (
    .I(\DLX_IDinst_slot_num_FFd1/FROM ),
    .O(CHOICE2516)
  );
  defparam \DLX_IDinst_Mmux__n0123_Result<1>1 .INIT = 16'hAAE2;
  X_LUT4 \DLX_IDinst_Mmux__n0123_Result<1>1  (
    .ADR0(DLX_IDinst_EPC[1]),
    .ADR1(DLX_IDinst__n03641_1),
    .ADR2(DLX_IFinst_NPC[1]),
    .ADR3(DLX_IDinst_Ker709161_1),
    .O(DLX_IDinst__n0123[1])
  );
  defparam \DLX_IDinst_Mmux__n0123_Result<0>1 .INIT = 16'hF0D8;
  X_LUT4 \DLX_IDinst_Mmux__n0123_Result<0>1  (
    .ADR0(DLX_IDinst__n03641_1),
    .ADR1(DLX_IFinst_NPC[0]),
    .ADR2(DLX_IDinst_EPC[0]),
    .ADR3(DLX_IDinst_N70918),
    .O(DLX_IDinst__n0123[0])
  );
  defparam \DLX_IDinst_Mmux__n0123_Result<3>1 .INIT = 16'hAEA2;
  X_LUT4 \DLX_IDinst_Mmux__n0123_Result<3>1  (
    .ADR0(DLX_IDinst_EPC[3]),
    .ADR1(DLX_IDinst__n03641_1),
    .ADR2(DLX_IDinst_Ker709161_1),
    .ADR3(DLX_IFinst_NPC[3]),
    .O(DLX_IDinst__n0123[3])
  );
  defparam \DLX_IDinst_Mmux__n0123_Result<2>1 .INIT = 16'hCCAC;
  X_LUT4 \DLX_IDinst_Mmux__n0123_Result<2>1  (
    .ADR0(DLX_IFinst_NPC[2]),
    .ADR1(DLX_IDinst_EPC[2]),
    .ADR2(DLX_IDinst__n03641_1),
    .ADR3(DLX_IDinst_Ker709161_1),
    .O(DLX_IDinst__n0123[2])
  );
  defparam \DLX_IDinst_Mmux__n0123_Result<5>1 .INIT = 16'hF0B8;
  X_LUT4 \DLX_IDinst_Mmux__n0123_Result<5>1  (
    .ADR0(DLX_IFinst_NPC[5]),
    .ADR1(DLX_IDinst__n03641_1),
    .ADR2(DLX_IDinst_EPC[5]),
    .ADR3(DLX_IDinst_Ker709161_1),
    .O(DLX_IDinst__n0123[5])
  );
  defparam \DLX_IDinst_Mmux__n0123_Result<4>1 .INIT = 16'hCCE4;
  X_LUT4 \DLX_IDinst_Mmux__n0123_Result<4>1  (
    .ADR0(DLX_IDinst__n03641_1),
    .ADR1(DLX_IDinst_EPC[4]),
    .ADR2(DLX_IFinst_NPC[4]),
    .ADR3(DLX_IDinst_Ker709161_1),
    .O(DLX_IDinst__n0123[4])
  );
  defparam \DLX_IDinst_Mmux__n0123_Result<7>1 .INIT = 16'hFB08;
  X_LUT4 \DLX_IDinst_Mmux__n0123_Result<7>1  (
    .ADR0(DLX_IFinst_NPC[7]),
    .ADR1(DLX_IDinst__n03641_1),
    .ADR2(DLX_IDinst_Ker709161_1),
    .ADR3(DLX_IDinst_EPC[7]),
    .O(DLX_IDinst__n0123[7])
  );
  defparam \DLX_IDinst_Mmux__n0123_Result<6>1 .INIT = 16'hAEA2;
  X_LUT4 \DLX_IDinst_Mmux__n0123_Result<6>1  (
    .ADR0(DLX_IDinst_EPC[6]),
    .ADR1(DLX_IDinst__n03641_1),
    .ADR2(DLX_IDinst_Ker709161_1),
    .ADR3(DLX_IFinst_NPC[6]),
    .O(DLX_IDinst__n0123[6])
  );
  defparam \DLX_IDinst_Mmux__n0123_Result<9>1 .INIT = 16'hAAE2;
  X_LUT4 \DLX_IDinst_Mmux__n0123_Result<9>1  (
    .ADR0(DLX_IDinst_EPC[9]),
    .ADR1(DLX_IDinst__n03641_1),
    .ADR2(DLX_IFinst_NPC[9]),
    .ADR3(DLX_IDinst_Ker709161_1),
    .O(DLX_IDinst__n0123[9])
  );
  defparam \DLX_IDinst_Mmux__n0123_Result<8>1 .INIT = 16'hFB08;
  X_LUT4 \DLX_IDinst_Mmux__n0123_Result<8>1  (
    .ADR0(DLX_IFinst_NPC[8]),
    .ADR1(DLX_IDinst__n03641_1),
    .ADR2(DLX_IDinst_Ker709161_1),
    .ADR3(DLX_IDinst_EPC[8]),
    .O(DLX_IDinst__n0123[8])
  );
  X_OR2 \DLX_EXinst_mem_to_reg_EX/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_mem_to_reg_EX/FFY/RST )
  );
  defparam DLX_EXinst_mem_read_EX_1125.INIT = 1'b0;
  X_FF DLX_EXinst_mem_read_EX_1125 (
    .I(\DLX_EXinst_mem_to_reg_EX/GROM ),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_mem_to_reg_EX/FFY/RST ),
    .O(DLX_EXinst_mem_read_EX)
  );
  defparam DLX_EXinst__n00101.INIT = 16'h0022;
  X_LUT4 DLX_EXinst__n00101 (
    .ADR0(DLX_IDinst_mem_to_reg),
    .ADR1(DLX_IDinst_counter[1]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_counter[0]),
    .O(DLX_EXinst__n0010)
  );
  defparam DLX_EXinst__n00111.INIT = 16'h0022;
  X_LUT4 DLX_EXinst__n00111 (
    .ADR0(DLX_IDinst_mem_read),
    .ADR1(DLX_IDinst_counter[1]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_counter[0]),
    .O(\DLX_EXinst_mem_to_reg_EX/GROM )
  );
  X_BUF \DLX_EXinst_mem_to_reg_EX/YUSED  (
    .I(\DLX_EXinst_mem_to_reg_EX/GROM ),
    .O(DLX_EXinst__n0011)
  );
  defparam vga_top_vga1_helpcounter_2.INIT = 1'b0;
  X_SFF vga_top_vga1_helpcounter_2 (
    .I(vga_top_vga1_helpcounter__n0000[2]),
    .CE(VCC),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(vga_top_vga1__n0052),
    .SRST(reset_IBUF_1),
    .O(vga_top_vga1_helpcounter[2])
  );
  defparam vga_top_vga1__n00521.INIT = 16'hC0FF;
  X_LUT4 vga_top_vga1__n00521 (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_helpcounter[1]),
    .ADR2(vga_top_vga1_helpcounter[2]),
    .ADR3(vga_top_vga1_clockcounter_FFd1),
    .O(\vga_top_vga1_helpcounter<2>/FROM )
  );
  defparam \vga_top_vga1_helpcounter_Madd__n0000_Mxor_Result<2>_Result1 .INIT = 16'h5FA0;
  X_LUT4 \vga_top_vga1_helpcounter_Madd__n0000_Mxor_Result<2>_Result1  (
    .ADR0(vga_top_vga1_helpcounter[0]),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_helpcounter[1]),
    .ADR3(vga_top_vga1_helpcounter[2]),
    .O(vga_top_vga1_helpcounter__n0000[2])
  );
  X_BUF \vga_top_vga1_helpcounter<2>/XUSED  (
    .I(\vga_top_vga1_helpcounter<2>/FROM ),
    .O(vga_top_vga1__n0052)
  );
  defparam \DLX_IDinst__n0118<2>1 .INIT = 16'h8888;
  X_LUT4 \DLX_IDinst__n0118<2>1  (
    .ADR0(DLX_IDinst_regB_eff[2]),
    .ADR1(DLX_IDinst_N69711),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IDinst_reg_out_B_2_1/GROM )
  );
  X_BUF \DLX_IDinst_reg_out_B_2_1/YUSED  (
    .I(\DLX_IDinst_reg_out_B_2_1/GROM ),
    .O(DLX_IDinst__n0118[2])
  );
  defparam \DLX_IDinst__n0118<3>1 .INIT = 16'hF000;
  X_LUT4 \DLX_IDinst__n0118<3>1  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_regB_eff[3]),
    .ADR3(DLX_IDinst_N69711),
    .O(\DLX_IDinst_reg_out_B<3>/GROM )
  );
  X_BUF \DLX_IDinst_reg_out_B<3>/YUSED  (
    .I(\DLX_IDinst_reg_out_B<3>/GROM ),
    .O(DLX_IDinst__n0118[3])
  );
  defparam \DLX_EXinst__n0006<13>277 .INIT = 16'hFCEC;
  X_LUT4 \DLX_EXinst__n0006<13>277  (
    .ADR0(CHOICE4311),
    .ADR1(DLX_EXinst_N63689),
    .ADR2(DLX_EXinst__n0149),
    .ADR3(CHOICE4343),
    .O(\DLX_EXinst_ALU_result<13>/FROM )
  );
  defparam \DLX_EXinst__n0006<12>267 .INIT = 16'hFCEC;
  X_LUT4 \DLX_EXinst__n0006<12>267  (
    .ADR0(CHOICE3879),
    .ADR1(DLX_EXinst_N63689),
    .ADR2(DLX_EXinst__n0149),
    .ADR3(CHOICE3909),
    .O(\DLX_EXinst_ALU_result<13>/GROM )
  );
  X_BUF \DLX_EXinst_ALU_result<13>/XUSED  (
    .I(\DLX_EXinst_ALU_result<13>/FROM ),
    .O(N115578)
  );
  X_BUF \DLX_EXinst_ALU_result<13>/YUSED  (
    .I(\DLX_EXinst_ALU_result<13>/GROM ),
    .O(N112968)
  );
  X_OR2 \DLX_MEMinst_RF_data_in<11>/FFY/RSTOR  (
    .I0(reset_IBUF_1),
    .I1(GSR),
    .O(\DLX_MEMinst_RF_data_in<11>/FFY/RST )
  );
  defparam DLX_MEMinst_RF_data_in_10.INIT = 1'b0;
  X_FF DLX_MEMinst_RF_data_in_10 (
    .I(DLX_MEMinst__n0000[10]),
    .CE(VCC),
    .CLK(\DLX_MEMinst_RF_data_in<11>/CKMUXNOT ),
    .SET(GND),
    .RST(\DLX_MEMinst_RF_data_in<11>/FFY/RST ),
    .O(DLX_MEMinst_RF_data_in[10])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<11>1 .INIT = 16'hACAC;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<11>1  (
    .ADR0(DM_read_data[11]),
    .ADR1(DLX_EXinst_ALU_result[11]),
    .ADR2(DLX_EXinst_mem_to_reg_EX),
    .ADR3(VCC),
    .O(DLX_MEMinst__n0000[11])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<10>1 .INIT = 16'hD8D8;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<10>1  (
    .ADR0(DLX_EXinst_mem_to_reg_EX),
    .ADR1(DM_read_data[10]),
    .ADR2(DLX_EXinst_ALU_result[10]),
    .ADR3(VCC),
    .O(DLX_MEMinst__n0000[10])
  );
  X_INV \DLX_MEMinst_RF_data_in<11>/CKINV  (
    .I(DLX_MEMlc_master_ctrlMEM_l),
    .O(\DLX_MEMinst_RF_data_in<11>/CKMUXNOT )
  );
  X_OR2 \DLX_MEMinst_RF_data_in<21>/FFY/RSTOR  (
    .I0(reset_IBUF_1),
    .I1(GSR),
    .O(\DLX_MEMinst_RF_data_in<21>/FFY/RST )
  );
  defparam DLX_MEMinst_RF_data_in_20.INIT = 1'b0;
  X_FF DLX_MEMinst_RF_data_in_20 (
    .I(DLX_MEMinst__n0000[20]),
    .CE(VCC),
    .CLK(\DLX_MEMinst_RF_data_in<21>/CKMUXNOT ),
    .SET(GND),
    .RST(\DLX_MEMinst_RF_data_in<21>/FFY/RST ),
    .O(DLX_MEMinst_RF_data_in[20])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<21>1 .INIT = 16'hEE22;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<21>1  (
    .ADR0(DLX_EXinst_ALU_result[21]),
    .ADR1(DLX_EXinst_mem_to_reg_EX),
    .ADR2(VCC),
    .ADR3(DM_read_data[21]),
    .O(DLX_MEMinst__n0000[21])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<20>1 .INIT = 16'hCCF0;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<20>1  (
    .ADR0(VCC),
    .ADR1(DM_read_data[20]),
    .ADR2(DLX_EXinst_ALU_result[20]),
    .ADR3(DLX_EXinst_mem_to_reg_EX),
    .O(DLX_MEMinst__n0000[20])
  );
  X_INV \DLX_MEMinst_RF_data_in<21>/CKINV  (
    .I(DLX_MEMlc_master_ctrlMEM_l),
    .O(\DLX_MEMinst_RF_data_in<21>/CKMUXNOT )
  );
  defparam DLX_EXinst_ALU_result_7_1_1126.INIT = 1'b0;
  X_FF DLX_EXinst_ALU_result_7_1_1126 (
    .I(\DM_addr_eff<7>/OD ),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DM_addr_eff<7>/OFF/RST ),
    .O(DLX_EXinst_ALU_result_7_1)
  );
  X_OR2 \DM_addr_eff<7>/OFF/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DM_addr_eff<7>/OFF/RST )
  );
  X_OR2 \DLX_MEMinst_RF_data_in<13>/FFY/RSTOR  (
    .I0(reset_IBUF_1),
    .I1(GSR),
    .O(\DLX_MEMinst_RF_data_in<13>/FFY/RST )
  );
  defparam DLX_MEMinst_RF_data_in_12.INIT = 1'b0;
  X_FF DLX_MEMinst_RF_data_in_12 (
    .I(DLX_MEMinst__n0000[12]),
    .CE(VCC),
    .CLK(\DLX_MEMinst_RF_data_in<13>/CKMUXNOT ),
    .SET(GND),
    .RST(\DLX_MEMinst_RF_data_in<13>/FFY/RST ),
    .O(DLX_MEMinst_RF_data_in[12])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<13>1 .INIT = 16'hFA0A;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<13>1  (
    .ADR0(DLX_EXinst_ALU_result[13]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_mem_to_reg_EX),
    .ADR3(DM_read_data[13]),
    .O(DLX_MEMinst__n0000[13])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<12>1 .INIT = 16'hF0AA;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<12>1  (
    .ADR0(DLX_EXinst_ALU_result[12]),
    .ADR1(VCC),
    .ADR2(DM_read_data[12]),
    .ADR3(DLX_EXinst_mem_to_reg_EX),
    .O(DLX_MEMinst__n0000[12])
  );
  X_INV \DLX_MEMinst_RF_data_in<13>/CKINV  (
    .I(DLX_MEMlc_master_ctrlMEM_l),
    .O(\DLX_MEMinst_RF_data_in<13>/CKMUXNOT )
  );
  X_OR2 \DLX_MEMinst_RF_data_in<31>/FFY/RSTOR  (
    .I0(reset_IBUF_1),
    .I1(GSR),
    .O(\DLX_MEMinst_RF_data_in<31>/FFY/RST )
  );
  defparam DLX_MEMinst_RF_data_in_30.INIT = 1'b0;
  X_FF DLX_MEMinst_RF_data_in_30 (
    .I(DLX_MEMinst__n0000[30]),
    .CE(VCC),
    .CLK(\DLX_MEMinst_RF_data_in<31>/CKMUXNOT ),
    .SET(GND),
    .RST(\DLX_MEMinst_RF_data_in<31>/FFY/RST ),
    .O(DLX_MEMinst_RF_data_in[30])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<31>1 .INIT = 16'hE2E2;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<31>1  (
    .ADR0(DLX_EXinst_ALU_result[31]),
    .ADR1(DLX_EXinst_mem_to_reg_EX),
    .ADR2(DM_read_data[31]),
    .ADR3(VCC),
    .O(DLX_MEMinst__n0000[31])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<30>1 .INIT = 16'hE4E4;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<30>1  (
    .ADR0(DLX_EXinst_mem_to_reg_EX),
    .ADR1(DLX_EXinst_ALU_result[30]),
    .ADR2(DM_read_data[30]),
    .ADR3(VCC),
    .O(DLX_MEMinst__n0000[30])
  );
  X_INV \DLX_MEMinst_RF_data_in<31>/CKINV  (
    .I(DLX_MEMlc_master_ctrlMEM_l),
    .O(\DLX_MEMinst_RF_data_in<31>/CKMUXNOT )
  );
  X_OR2 \DLX_MEMinst_RF_data_in<23>/FFY/RSTOR  (
    .I0(reset_IBUF_1),
    .I1(GSR),
    .O(\DLX_MEMinst_RF_data_in<23>/FFY/RST )
  );
  defparam DLX_MEMinst_RF_data_in_22.INIT = 1'b0;
  X_FF DLX_MEMinst_RF_data_in_22 (
    .I(DLX_MEMinst__n0000[22]),
    .CE(VCC),
    .CLK(\DLX_MEMinst_RF_data_in<23>/CKMUXNOT ),
    .SET(GND),
    .RST(\DLX_MEMinst_RF_data_in<23>/FFY/RST ),
    .O(DLX_MEMinst_RF_data_in[22])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<23>1 .INIT = 16'hAACC;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<23>1  (
    .ADR0(DM_read_data[23]),
    .ADR1(DLX_EXinst_ALU_result[23]),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_mem_to_reg_EX),
    .O(DLX_MEMinst__n0000[23])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<22>1 .INIT = 16'hF0CC;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<22>1  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_ALU_result[22]),
    .ADR2(DM_read_data[22]),
    .ADR3(DLX_EXinst_mem_to_reg_EX),
    .O(DLX_MEMinst__n0000[22])
  );
  X_INV \DLX_MEMinst_RF_data_in<23>/CKINV  (
    .I(DLX_MEMlc_master_ctrlMEM_l),
    .O(\DLX_MEMinst_RF_data_in<23>/CKMUXNOT )
  );
  X_OR2 \DLX_MEMinst_RF_data_in<15>/FFY/RSTOR  (
    .I0(reset_IBUF_1),
    .I1(GSR),
    .O(\DLX_MEMinst_RF_data_in<15>/FFY/RST )
  );
  defparam DLX_MEMinst_RF_data_in_14.INIT = 1'b0;
  X_FF DLX_MEMinst_RF_data_in_14 (
    .I(DLX_MEMinst__n0000[14]),
    .CE(VCC),
    .CLK(\DLX_MEMinst_RF_data_in<15>/CKMUXNOT ),
    .SET(GND),
    .RST(\DLX_MEMinst_RF_data_in<15>/FFY/RST ),
    .O(DLX_MEMinst_RF_data_in[14])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<15>1 .INIT = 16'hD8D8;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<15>1  (
    .ADR0(DLX_EXinst_mem_to_reg_EX),
    .ADR1(DM_read_data[15]),
    .ADR2(DLX_EXinst_ALU_result[15]),
    .ADR3(VCC),
    .O(DLX_MEMinst__n0000[15])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<14>1 .INIT = 16'hEE44;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<14>1  (
    .ADR0(DLX_EXinst_mem_to_reg_EX),
    .ADR1(DLX_EXinst_ALU_result[14]),
    .ADR2(VCC),
    .ADR3(DM_read_data[14]),
    .O(DLX_MEMinst__n0000[14])
  );
  X_INV \DLX_MEMinst_RF_data_in<15>/CKINV  (
    .I(DLX_MEMlc_master_ctrlMEM_l),
    .O(\DLX_MEMinst_RF_data_in<15>/CKMUXNOT )
  );
  X_OR2 \DLX_MEMinst_RF_data_in<25>/FFY/RSTOR  (
    .I0(reset_IBUF_1),
    .I1(GSR),
    .O(\DLX_MEMinst_RF_data_in<25>/FFY/RST )
  );
  defparam DLX_MEMinst_RF_data_in_24.INIT = 1'b0;
  X_FF DLX_MEMinst_RF_data_in_24 (
    .I(DLX_MEMinst__n0000[24]),
    .CE(VCC),
    .CLK(\DLX_MEMinst_RF_data_in<25>/CKMUXNOT ),
    .SET(GND),
    .RST(\DLX_MEMinst_RF_data_in<25>/FFY/RST ),
    .O(DLX_MEMinst_RF_data_in[24])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<25>1 .INIT = 16'hD8D8;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<25>1  (
    .ADR0(DLX_EXinst_mem_to_reg_EX),
    .ADR1(DM_read_data[25]),
    .ADR2(DLX_EXinst_ALU_result[25]),
    .ADR3(VCC),
    .O(DLX_MEMinst__n0000[25])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<24>1 .INIT = 16'hEE22;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<24>1  (
    .ADR0(DLX_EXinst_ALU_result[24]),
    .ADR1(DLX_EXinst_mem_to_reg_EX),
    .ADR2(VCC),
    .ADR3(DM_read_data[24]),
    .O(DLX_MEMinst__n0000[24])
  );
  X_INV \DLX_MEMinst_RF_data_in<25>/CKINV  (
    .I(DLX_MEMlc_master_ctrlMEM_l),
    .O(\DLX_MEMinst_RF_data_in<25>/CKMUXNOT )
  );
  X_OR2 \DLX_MEMinst_RF_data_in<17>/FFY/RSTOR  (
    .I0(reset_IBUF_1),
    .I1(GSR),
    .O(\DLX_MEMinst_RF_data_in<17>/FFY/RST )
  );
  defparam DLX_MEMinst_RF_data_in_16.INIT = 1'b0;
  X_FF DLX_MEMinst_RF_data_in_16 (
    .I(DLX_MEMinst__n0000[16]),
    .CE(VCC),
    .CLK(\DLX_MEMinst_RF_data_in<17>/CKMUXNOT ),
    .SET(GND),
    .RST(\DLX_MEMinst_RF_data_in<17>/FFY/RST ),
    .O(DLX_MEMinst_RF_data_in[16])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<17>1 .INIT = 16'hEE44;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<17>1  (
    .ADR0(DLX_EXinst_mem_to_reg_EX),
    .ADR1(DLX_EXinst_ALU_result[17]),
    .ADR2(VCC),
    .ADR3(DM_read_data[17]),
    .O(DLX_MEMinst__n0000[17])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<16>1 .INIT = 16'hFC0C;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<16>1  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_ALU_result[16]),
    .ADR2(DLX_EXinst_mem_to_reg_EX),
    .ADR3(DM_read_data[16]),
    .O(DLX_MEMinst__n0000[16])
  );
  X_INV \DLX_MEMinst_RF_data_in<17>/CKINV  (
    .I(DLX_MEMlc_master_ctrlMEM_l),
    .O(\DLX_MEMinst_RF_data_in<17>/CKMUXNOT )
  );
  X_OR2 \DLX_MEMinst_RF_data_in<27>/FFY/RSTOR  (
    .I0(reset_IBUF_1),
    .I1(GSR),
    .O(\DLX_MEMinst_RF_data_in<27>/FFY/RST )
  );
  defparam DLX_MEMinst_RF_data_in_26.INIT = 1'b0;
  X_FF DLX_MEMinst_RF_data_in_26 (
    .I(DLX_MEMinst__n0000[26]),
    .CE(VCC),
    .CLK(\DLX_MEMinst_RF_data_in<27>/CKMUXNOT ),
    .SET(GND),
    .RST(\DLX_MEMinst_RF_data_in<27>/FFY/RST ),
    .O(DLX_MEMinst_RF_data_in[26])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<27>1 .INIT = 16'hFC0C;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<27>1  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_ALU_result[27]),
    .ADR2(DLX_EXinst_mem_to_reg_EX),
    .ADR3(DM_read_data[27]),
    .O(DLX_MEMinst__n0000[27])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<26>1 .INIT = 16'hCCAA;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<26>1  (
    .ADR0(DLX_EXinst_ALU_result[26]),
    .ADR1(DM_read_data[26]),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_mem_to_reg_EX),
    .O(DLX_MEMinst__n0000[26])
  );
  X_INV \DLX_MEMinst_RF_data_in<27>/CKINV  (
    .I(DLX_MEMlc_master_ctrlMEM_l),
    .O(\DLX_MEMinst_RF_data_in<27>/CKMUXNOT )
  );
  X_OR2 \DLX_MEMinst_RF_data_in<19>/FFY/RSTOR  (
    .I0(reset_IBUF_1),
    .I1(GSR),
    .O(\DLX_MEMinst_RF_data_in<19>/FFY/RST )
  );
  defparam DLX_MEMinst_RF_data_in_18.INIT = 1'b0;
  X_FF DLX_MEMinst_RF_data_in_18 (
    .I(DLX_MEMinst__n0000[18]),
    .CE(VCC),
    .CLK(\DLX_MEMinst_RF_data_in<19>/CKMUXNOT ),
    .SET(GND),
    .RST(\DLX_MEMinst_RF_data_in<19>/FFY/RST ),
    .O(DLX_MEMinst_RF_data_in[18])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<19>1 .INIT = 16'hEE22;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<19>1  (
    .ADR0(DLX_EXinst_ALU_result[19]),
    .ADR1(DLX_EXinst_mem_to_reg_EX),
    .ADR2(VCC),
    .ADR3(DM_read_data[19]),
    .O(DLX_MEMinst__n0000[19])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<18>1 .INIT = 16'hE2E2;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<18>1  (
    .ADR0(DLX_EXinst_ALU_result[18]),
    .ADR1(DLX_EXinst_mem_to_reg_EX),
    .ADR2(DM_read_data[18]),
    .ADR3(VCC),
    .O(DLX_MEMinst__n0000[18])
  );
  X_INV \DLX_MEMinst_RF_data_in<19>/CKINV  (
    .I(DLX_MEMlc_master_ctrlMEM_l),
    .O(\DLX_MEMinst_RF_data_in<19>/CKMUXNOT )
  );
  X_OR2 \DLX_MEMinst_RF_data_in<29>/FFY/RSTOR  (
    .I0(reset_IBUF_1),
    .I1(GSR),
    .O(\DLX_MEMinst_RF_data_in<29>/FFY/RST )
  );
  defparam DLX_MEMinst_RF_data_in_28.INIT = 1'b0;
  X_FF DLX_MEMinst_RF_data_in_28 (
    .I(DLX_MEMinst__n0000[28]),
    .CE(VCC),
    .CLK(\DLX_MEMinst_RF_data_in<29>/CKMUXNOT ),
    .SET(GND),
    .RST(\DLX_MEMinst_RF_data_in<29>/FFY/RST ),
    .O(DLX_MEMinst_RF_data_in[28])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<29>1 .INIT = 16'hAFA0;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<29>1  (
    .ADR0(DM_read_data[29]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_mem_to_reg_EX),
    .ADR3(DLX_EXinst_ALU_result[29]),
    .O(DLX_MEMinst__n0000[29])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<28>1 .INIT = 16'hBB88;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<28>1  (
    .ADR0(DM_read_data[28]),
    .ADR1(DLX_EXinst_mem_to_reg_EX),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_ALU_result[28]),
    .O(DLX_MEMinst__n0000[28])
  );
  X_INV \DLX_MEMinst_RF_data_in<29>/CKINV  (
    .I(DLX_MEMlc_master_ctrlMEM_l),
    .O(\DLX_MEMinst_RF_data_in<29>/CKMUXNOT )
  );
  X_OR2 \DLX_IDinst_current_IR<11>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_current_IR<11>/FFY/RST )
  );
  defparam DLX_IDinst_current_IR_10.INIT = 1'b0;
  X_FF DLX_IDinst_current_IR_10 (
    .I(\DLX_IDinst_current_IR<11>/GROM ),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_current_IR<11>/FFY/RST ),
    .O(DLX_IDinst_current_IR[10])
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<11>1 .INIT = 16'hF0E2;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<11>1  (
    .ADR0(DLX_IFinst_IR_latched[11]),
    .ADR1(DLX_IDinst_counter[1]),
    .ADR2(DLX_IDinst_current_IR[11]),
    .ADR3(DLX_IDinst_counter[0]),
    .O(\DLX_IDinst_current_IR<11>/FROM )
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<10>1 .INIT = 16'hF0E2;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<10>1  (
    .ADR0(DLX_IFinst_IR_latched[10]),
    .ADR1(DLX_IDinst_counter[1]),
    .ADR2(DLX_IDinst_current_IR[10]),
    .ADR3(DLX_IDinst_counter[0]),
    .O(\DLX_IDinst_current_IR<11>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<11>/XUSED  (
    .I(\DLX_IDinst_current_IR<11>/FROM ),
    .O(DLX_IDinst_jtarget[11])
  );
  X_BUF \DLX_IDinst_current_IR<11>/YUSED  (
    .I(\DLX_IDinst_current_IR<11>/GROM ),
    .O(DLX_IDinst_jtarget[10])
  );
  X_ZERO \DLX_IDinst_current_IR<20>/LOGIC_ZERO_1127  (
    .O(\DLX_IDinst_current_IR<20>/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mcompar__n0315_inst_cy_264 (
    .IA(\DLX_IDinst_current_IR<20>/LOGIC_ZERO ),
    .IB(\DLX_IDinst_current_IR<20>/CYINIT ),
    .SEL(DLX_IDinst_Mcompar__n0315_inst_lut4_42),
    .O(\DLX_IDinst_current_IR<20>/CYMUXF )
  );
  defparam DLX_IDinst_Mcompar__n0315_inst_lut4_421.INIT = 16'hA5A5;
  X_LUT4 DLX_IDinst_Mcompar__n0315_inst_lut4_421 (
    .ADR0(DLX_IDinst_regB_index[4]),
    .ADR1(VCC),
    .ADR2(DLX_MEMinst_reg_dst_out[4]),
    .ADR3(VCC),
    .O(DLX_IDinst_Mcompar__n0315_inst_lut4_42)
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<20>1 .INIT = 16'hF0E4;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<20>1  (
    .ADR0(DLX_IDinst_counter[0]),
    .ADR1(DLX_IFinst_IR_latched[20]),
    .ADR2(DLX_IDinst_current_IR[20]),
    .ADR3(DLX_IDinst_counter[1]),
    .O(\DLX_IDinst_current_IR<20>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<20>/XBUSED  (
    .I(\DLX_IDinst_current_IR<20>/CYMUXF ),
    .O(DLX_IDinst__n0315)
  );
  X_BUF \DLX_IDinst_current_IR<20>/YUSED  (
    .I(\DLX_IDinst_current_IR<20>/GROM ),
    .O(DLX_IDinst_regB_index[4])
  );
  X_BUF \DLX_IDinst_current_IR<20>/CYINIT_1128  (
    .I(DLX_IDinst_Mcompar__n0315_inst_cy_263),
    .O(\DLX_IDinst_current_IR<20>/CYINIT )
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<13>1 .INIT = 16'hFE02;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<13>1  (
    .ADR0(DLX_IFinst_IR_latched[13]),
    .ADR1(DLX_IDinst_counter[0]),
    .ADR2(DLX_IDinst_counter[1]),
    .ADR3(DLX_IDinst_current_IR[13]),
    .O(\DLX_IDinst_current_IR<13>/FROM )
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<12>1 .INIT = 16'hAAB8;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<12>1  (
    .ADR0(DLX_IDinst_current_IR[12]),
    .ADR1(DLX_IDinst_counter[1]),
    .ADR2(DLX_IFinst_IR_latched[12]),
    .ADR3(DLX_IDinst_counter[0]),
    .O(\DLX_IDinst_current_IR<13>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<13>/XUSED  (
    .I(\DLX_IDinst_current_IR<13>/FROM ),
    .O(DLX_IDinst_jtarget[13])
  );
  X_BUF \DLX_IDinst_current_IR<13>/YUSED  (
    .I(\DLX_IDinst_current_IR<13>/GROM ),
    .O(DLX_IDinst_jtarget[12])
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<21>1 .INIT = 16'hAAAC;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<21>1  (
    .ADR0(DLX_IDinst_current_IR[21]),
    .ADR1(DLX_IFinst_IR_latched[21]),
    .ADR2(DLX_IDinst_counter[1]),
    .ADR3(DLX_IDinst_counter[0]),
    .O(\DLX_IDinst_current_IR<21>/FROM )
  );
  defparam \DLX_IDinst__n0117<21>15 .INIT = 16'h3088;
  X_LUT4 \DLX_IDinst__n0117<21>15  (
    .ADR0(DLX_IDinst_EPC[21]),
    .ADR1(DLX_IDinst_regA_index[1]),
    .ADR2(DLX_IDinst_Cause_Reg[21]),
    .ADR3(DLX_IDinst_regA_index[0]),
    .O(\DLX_IDinst_current_IR<21>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<21>/XUSED  (
    .I(\DLX_IDinst_current_IR<21>/FROM ),
    .O(DLX_IDinst_regA_index[0])
  );
  X_BUF \DLX_IDinst_current_IR<21>/YUSED  (
    .I(\DLX_IDinst_current_IR<21>/GROM ),
    .O(CHOICE2398)
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<15>1 .INIT = 16'hFE02;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<15>1  (
    .ADR0(DLX_IFinst_IR_latched[15]),
    .ADR1(DLX_IDinst_counter[1]),
    .ADR2(DLX_IDinst_counter[0]),
    .ADR3(DLX_IDinst_current_IR[15]),
    .O(\DLX_IDinst_current_IR<15>/FROM )
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<14>1 .INIT = 16'hF0E2;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<14>1  (
    .ADR0(DLX_IFinst_IR_latched[14]),
    .ADR1(DLX_IDinst_counter[0]),
    .ADR2(DLX_IDinst_current_IR[14]),
    .ADR3(DLX_IDinst_counter[1]),
    .O(\DLX_IDinst_current_IR<15>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<15>/XUSED  (
    .I(\DLX_IDinst_current_IR<15>/FROM ),
    .O(DLX_IDinst_jtarget[15])
  );
  X_BUF \DLX_IDinst_current_IR<15>/YUSED  (
    .I(\DLX_IDinst_current_IR<15>/GROM ),
    .O(DLX_IDinst_jtarget[14])
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<23>1 .INIT = 16'hAAAC;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<23>1  (
    .ADR0(DLX_IDinst_current_IR[23]),
    .ADR1(DLX_IFinst_IR_latched[23]),
    .ADR2(DLX_IDinst_counter[0]),
    .ADR3(DLX_IDinst_counter[1]),
    .O(\DLX_IDinst_current_IR<23>/FROM )
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<22>1 .INIT = 16'hFE10;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<22>1  (
    .ADR0(DLX_IDinst_counter[0]),
    .ADR1(DLX_IDinst_counter[1]),
    .ADR2(DLX_IFinst_IR_latched[22]),
    .ADR3(DLX_IDinst_current_IR[22]),
    .O(\DLX_IDinst_current_IR<23>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<23>/XUSED  (
    .I(\DLX_IDinst_current_IR<23>/FROM ),
    .O(DLX_IDinst_regA_index[2])
  );
  X_BUF \DLX_IDinst_current_IR<23>/YUSED  (
    .I(\DLX_IDinst_current_IR<23>/GROM ),
    .O(DLX_IDinst_regA_index[1])
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<30>1 .INIT = 16'hF0E4;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<30>1  (
    .ADR0(DLX_IDinst_counter[0]),
    .ADR1(DLX_IFinst_IR_latched[30]),
    .ADR2(DLX_IDinst_current_IR[30]),
    .ADR3(DLX_IDinst_counter[1]),
    .O(\DLX_IDinst_current_IR<30>/FROM )
  );
  defparam DLX_IDinst_N700061.INIT = 16'h0040;
  X_LUT4 DLX_IDinst_N700061 (
    .ADR0(DLX_IDinst_IR_latched[27]),
    .ADR1(DLX_IDinst_IR_latched[30]),
    .ADR2(DLX_IDinst_N70991),
    .ADR3(DLX_IDinst__n03641_1),
    .O(\DLX_IDinst_current_IR<30>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<30>/XUSED  (
    .I(\DLX_IDinst_current_IR<30>/FROM ),
    .O(DLX_IDinst_IR_latched[30])
  );
  X_BUF \DLX_IDinst_current_IR<30>/YUSED  (
    .I(\DLX_IDinst_current_IR<30>/GROM ),
    .O(DLX_IDinst_N70006)
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<31>1 .INIT = 16'hF0E2;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<31>1  (
    .ADR0(DLX_IFinst_IR_latched[31]),
    .ADR1(DLX_IDinst_counter[0]),
    .ADR2(DLX_IDinst_current_IR[31]),
    .ADR3(DLX_IDinst_counter[1]),
    .O(\DLX_IDinst_current_IR<31>/FROM )
  );
  defparam DLX_IDinst__n00621.INIT = 16'hD0F0;
  X_LUT4 DLX_IDinst__n00621 (
    .ADR0(DLX_IDinst__n0338),
    .ADR1(DLX_IDinst_IR_latched[30]),
    .ADR2(DLX_IDinst__n0132),
    .ADR3(DLX_IDinst_IR_latched[31]),
    .O(\DLX_IDinst_current_IR<31>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<31>/XUSED  (
    .I(\DLX_IDinst_current_IR<31>/FROM ),
    .O(DLX_IDinst_IR_latched[31])
  );
  X_BUF \DLX_IDinst_current_IR<31>/YUSED  (
    .I(\DLX_IDinst_current_IR<31>/GROM ),
    .O(DLX_IDinst__n0062)
  );
  defparam DLX_EXinst_ALU_result_8_1_1129.INIT = 1'b0;
  X_FF DLX_EXinst_ALU_result_8_1_1129 (
    .I(\DM_addr_eff<8>/OD ),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DM_addr_eff<8>/OFF/RST ),
    .O(DLX_EXinst_ALU_result_8_1)
  );
  X_OR2 \DM_addr_eff<8>/OFF/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DM_addr_eff<8>/OFF/RST )
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<24>1 .INIT = 16'hCCD8;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<24>1  (
    .ADR0(DLX_IDinst_counter[0]),
    .ADR1(DLX_IDinst_current_IR[24]),
    .ADR2(DLX_IFinst_IR_latched[24]),
    .ADR3(DLX_IDinst_counter[1]),
    .O(\DLX_IDinst_current_IR<24>/FROM )
  );
  defparam DLX_IDinst_Ker706561.INIT = 16'h0005;
  X_LUT4 DLX_IDinst_Ker706561 (
    .ADR0(DLX_IDinst_regA_index[2]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_regA_index[4]),
    .ADR3(DLX_IDinst_regA_index[3]),
    .O(\DLX_IDinst_current_IR<24>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<24>/XUSED  (
    .I(\DLX_IDinst_current_IR<24>/FROM ),
    .O(DLX_IDinst_regA_index[3])
  );
  X_BUF \DLX_IDinst_current_IR<24>/YUSED  (
    .I(\DLX_IDinst_current_IR<24>/GROM ),
    .O(DLX_IDinst_N70658)
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<17>1 .INIT = 16'hF0E2;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<17>1  (
    .ADR0(DLX_IFinst_IR_latched[17]),
    .ADR1(DLX_IDinst_counter[0]),
    .ADR2(DLX_IDinst_current_IR[17]),
    .ADR3(DLX_IDinst_counter[1]),
    .O(\DLX_IDinst_current_IR<17>/FROM )
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<16>1 .INIT = 16'hF0E2;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<16>1  (
    .ADR0(DLX_IFinst_IR_latched[16]),
    .ADR1(DLX_IDinst_counter[1]),
    .ADR2(DLX_IDinst_current_IR[16]),
    .ADR3(DLX_IDinst_counter[0]),
    .O(\DLX_IDinst_current_IR<17>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<17>/XUSED  (
    .I(\DLX_IDinst_current_IR<17>/FROM ),
    .O(DLX_IDinst_regB_index[1])
  );
  X_BUF \DLX_IDinst_current_IR<17>/YUSED  (
    .I(\DLX_IDinst_current_IR<17>/GROM ),
    .O(DLX_IDinst_regB_index[0])
  );
  X_ZERO \DLX_IDinst_current_IR<25>/LOGIC_ZERO_1130  (
    .O(\DLX_IDinst_current_IR<25>/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mcompar__n0314_inst_cy_264 (
    .IA(\DLX_IDinst_current_IR<25>/LOGIC_ZERO ),
    .IB(\DLX_IDinst_current_IR<25>/CYINIT ),
    .SEL(DLX_IDinst_Mcompar__n0314_inst_lut4_42),
    .O(\DLX_IDinst_current_IR<25>/CYMUXF )
  );
  defparam DLX_IDinst_Mcompar__n0314_inst_lut4_421.INIT = 16'hC3C3;
  X_LUT4 DLX_IDinst_Mcompar__n0314_inst_lut4_421 (
    .ADR0(VCC),
    .ADR1(DLX_MEMinst_reg_dst_out[4]),
    .ADR2(DLX_IDinst_regA_index[4]),
    .ADR3(VCC),
    .O(DLX_IDinst_Mcompar__n0314_inst_lut4_42)
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<25>1 .INIT = 16'hCCCA;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<25>1  (
    .ADR0(DLX_IFinst_IR_latched[25]),
    .ADR1(DLX_IDinst_current_IR[25]),
    .ADR2(DLX_IDinst_counter[1]),
    .ADR3(DLX_IDinst_counter[0]),
    .O(\DLX_IDinst_current_IR<25>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<25>/XBUSED  (
    .I(\DLX_IDinst_current_IR<25>/CYMUXF ),
    .O(DLX_IDinst__n0314)
  );
  X_BUF \DLX_IDinst_current_IR<25>/YUSED  (
    .I(\DLX_IDinst_current_IR<25>/GROM ),
    .O(DLX_IDinst_regA_index[4])
  );
  X_BUF \DLX_IDinst_current_IR<25>/CYINIT_1131  (
    .I(DLX_IDinst_Mcompar__n0314_inst_cy_263),
    .O(\DLX_IDinst_current_IR<25>/CYINIT )
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<26>1 .INIT = 16'hFE04;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<26>1  (
    .ADR0(DLX_IDinst_counter[1]),
    .ADR1(DLX_IFinst_IR_latched[26]),
    .ADR2(DLX_IDinst_counter[0]),
    .ADR3(DLX_IDinst_current_IR[26]),
    .O(\DLX_IDinst_current_IR<26>/FROM )
  );
  defparam DLX_IDinst__n008912.INIT = 16'hAFFF;
  X_LUT4 DLX_IDinst__n008912 (
    .ADR0(DLX_IDinst_IR_latched[28]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_IR_latched[29]),
    .ADR3(DLX_IDinst_IR_latched[26]),
    .O(\DLX_IDinst_current_IR<26>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<26>/XUSED  (
    .I(\DLX_IDinst_current_IR<26>/FROM ),
    .O(DLX_IDinst_IR_latched[26])
  );
  X_BUF \DLX_IDinst_current_IR<26>/YUSED  (
    .I(\DLX_IDinst_current_IR<26>/GROM ),
    .O(CHOICE2847)
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<19>1 .INIT = 16'hCCD8;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<19>1  (
    .ADR0(DLX_IDinst_counter[0]),
    .ADR1(DLX_IDinst_current_IR[19]),
    .ADR2(DLX_IFinst_IR_latched[19]),
    .ADR3(DLX_IDinst_counter[1]),
    .O(\DLX_IDinst_current_IR<19>/FROM )
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<18>1 .INIT = 16'hF0E4;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<18>1  (
    .ADR0(DLX_IDinst_counter[0]),
    .ADR1(DLX_IFinst_IR_latched[18]),
    .ADR2(DLX_IDinst_current_IR[18]),
    .ADR3(DLX_IDinst_counter[1]),
    .O(\DLX_IDinst_current_IR<19>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<19>/XUSED  (
    .I(\DLX_IDinst_current_IR<19>/FROM ),
    .O(DLX_IDinst_regB_index[3])
  );
  X_BUF \DLX_IDinst_current_IR<19>/YUSED  (
    .I(\DLX_IDinst_current_IR<19>/GROM ),
    .O(DLX_IDinst_regB_index[2])
  );
  defparam DLX_IDinst__n02501_SW0.INIT = 16'hCCCA;
  X_LUT4 DLX_IDinst__n02501_SW0 (
    .ADR0(DLX_IFinst_IR_latched[27]),
    .ADR1(DLX_IDinst_current_IR[27]),
    .ADR2(DLX_IDinst_counter[0]),
    .ADR3(DLX_IDinst_counter[1]),
    .O(\DLX_IDinst_current_IR<27>/FROM )
  );
  defparam DLX_IDinst__n033915.INIT = 16'h0023;
  X_LUT4 DLX_IDinst__n033915 (
    .ADR0(DLX_IDinst_IR_latched[28]),
    .ADR1(DLX_IDinst_IR_latched[30]),
    .ADR2(DLX_IDinst_IR_latched[26]),
    .ADR3(DLX_IDinst_IR_latched[27]),
    .O(\DLX_IDinst_current_IR<27>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<27>/XUSED  (
    .I(\DLX_IDinst_current_IR<27>/FROM ),
    .O(DLX_IDinst_IR_latched[27])
  );
  X_BUF \DLX_IDinst_current_IR<27>/YUSED  (
    .I(\DLX_IDinst_current_IR<27>/GROM ),
    .O(CHOICE1387)
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<28>1 .INIT = 16'hFE04;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<28>1  (
    .ADR0(DLX_IDinst_counter[1]),
    .ADR1(DLX_IFinst_IR_latched[28]),
    .ADR2(DLX_IDinst_counter[0]),
    .ADR3(DLX_IDinst_current_IR[28]),
    .O(\DLX_IDinst_current_IR<28>/FROM )
  );
  defparam DLX_IDinst__n034241.INIT = 16'h0054;
  X_LUT4 DLX_IDinst__n034241 (
    .ADR0(DLX_IDinst_IR_latched[30]),
    .ADR1(CHOICE1796),
    .ADR2(CHOICE1800),
    .ADR3(DLX_IDinst_IR_latched[28]),
    .O(\DLX_IDinst_current_IR<28>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<28>/XUSED  (
    .I(\DLX_IDinst_current_IR<28>/FROM ),
    .O(DLX_IDinst_IR_latched[28])
  );
  X_BUF \DLX_IDinst_current_IR<28>/YUSED  (
    .I(\DLX_IDinst_current_IR<28>/GROM ),
    .O(N100686)
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<29>1 .INIT = 16'hFE10;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<29>1  (
    .ADR0(DLX_IDinst_counter[1]),
    .ADR1(DLX_IDinst_counter[0]),
    .ADR2(DLX_IFinst_IR_latched[29]),
    .ADR3(DLX_IDinst_current_IR[29]),
    .O(\DLX_IDinst_current_IR<29>/FROM )
  );
  defparam DLX_IDinst_Ker709071.INIT = 16'h0027;
  X_LUT4 DLX_IDinst_Ker709071 (
    .ADR0(DLX_EXinst__n0149),
    .ADR1(DLX_IFinst_IR_latched[31]),
    .ADR2(DLX_IDinst_current_IR[31]),
    .ADR3(DLX_IDinst_IR_latched[29]),
    .O(\DLX_IDinst_current_IR<29>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<29>/XUSED  (
    .I(\DLX_IDinst_current_IR<29>/FROM ),
    .O(DLX_IDinst_IR_latched[29])
  );
  X_BUF \DLX_IDinst_current_IR<29>/YUSED  (
    .I(\DLX_IDinst_current_IR<29>/GROM ),
    .O(DLX_IDinst_N70909)
  );
  defparam \DLX_IDinst_Mmux__n0123_Result<11>1 .INIT = 16'hF2D0;
  X_LUT4 \DLX_IDinst_Mmux__n0123_Result<11>1  (
    .ADR0(DLX_IDinst__n03641_1),
    .ADR1(DLX_IDinst_N70918),
    .ADR2(DLX_IDinst_EPC[11]),
    .ADR3(DLX_IFinst_NPC[11]),
    .O(DLX_IDinst__n0123[11])
  );
  defparam \DLX_IDinst_Mmux__n0123_Result<10>1 .INIT = 16'hCEC4;
  X_LUT4 \DLX_IDinst_Mmux__n0123_Result<10>1  (
    .ADR0(DLX_IDinst__n03641_1),
    .ADR1(DLX_IDinst_EPC[10]),
    .ADR2(DLX_IDinst_N70918),
    .ADR3(DLX_IFinst_NPC[10]),
    .O(DLX_IDinst__n0123[10])
  );
  defparam \DLX_IDinst_Mmux__n0123_Result<13>1 .INIT = 16'hFD20;
  X_LUT4 \DLX_IDinst_Mmux__n0123_Result<13>1  (
    .ADR0(DLX_IDinst__n03641_1),
    .ADR1(DLX_IDinst_Ker709161_1),
    .ADR2(DLX_IFinst_NPC[13]),
    .ADR3(DLX_IDinst_EPC[13]),
    .O(DLX_IDinst__n0123[13])
  );
  defparam \DLX_IDinst_Mmux__n0123_Result<12>1 .INIT = 16'hFB40;
  X_LUT4 \DLX_IDinst_Mmux__n0123_Result<12>1  (
    .ADR0(DLX_IDinst_Ker709161_1),
    .ADR1(DLX_IDinst__n03641_1),
    .ADR2(DLX_IFinst_NPC[12]),
    .ADR3(DLX_IDinst_EPC[12]),
    .O(DLX_IDinst__n0123[12])
  );
  defparam \DLX_IDinst_Mmux__n0123_Result<21>1 .INIT = 16'hBA8A;
  X_LUT4 \DLX_IDinst_Mmux__n0123_Result<21>1  (
    .ADR0(DLX_IDinst_EPC[21]),
    .ADR1(DLX_IDinst_Ker709161_1),
    .ADR2(DLX_IDinst__n03641_1),
    .ADR3(DLX_IFinst_NPC[21]),
    .O(DLX_IDinst__n0123[21])
  );
  defparam \DLX_IDinst_Mmux__n0123_Result<20>1 .INIT = 16'hEF40;
  X_LUT4 \DLX_IDinst_Mmux__n0123_Result<20>1  (
    .ADR0(DLX_IDinst_Ker709161_1),
    .ADR1(DLX_IFinst_NPC[20]),
    .ADR2(DLX_IDinst__n03641_1),
    .ADR3(DLX_IDinst_EPC[20]),
    .O(DLX_IDinst__n0123[20])
  );
  defparam \DLX_IDinst_Mmux__n0123_Result<15>1 .INIT = 16'hACAA;
  X_LUT4 \DLX_IDinst_Mmux__n0123_Result<15>1  (
    .ADR0(DLX_IDinst_EPC[15]),
    .ADR1(DLX_IFinst_NPC[15]),
    .ADR2(DLX_IDinst_Ker709161_1),
    .ADR3(DLX_IDinst__n03641_1),
    .O(DLX_IDinst__n0123[15])
  );
  defparam \DLX_IDinst_Mmux__n0123_Result<14>1 .INIT = 16'hF0D8;
  X_LUT4 \DLX_IDinst_Mmux__n0123_Result<14>1  (
    .ADR0(DLX_IDinst__n03641_1),
    .ADR1(DLX_IFinst_NPC[14]),
    .ADR2(DLX_IDinst_EPC[14]),
    .ADR3(DLX_IDinst_Ker709161_1),
    .O(DLX_IDinst__n0123[14])
  );
  defparam \DLX_IDinst_Mmux__n0123_Result<23>1 .INIT = 16'hB8AA;
  X_LUT4 \DLX_IDinst_Mmux__n0123_Result<23>1  (
    .ADR0(DLX_IDinst_EPC[23]),
    .ADR1(DLX_IDinst_Ker709161_1),
    .ADR2(DLX_IFinst_NPC[23]),
    .ADR3(DLX_IDinst__n03641_1),
    .O(DLX_IDinst__n0123[23])
  );
  defparam \DLX_IDinst_Mmux__n0123_Result<22>1 .INIT = 16'hAEA2;
  X_LUT4 \DLX_IDinst_Mmux__n0123_Result<22>1  (
    .ADR0(DLX_IDinst_EPC[22]),
    .ADR1(DLX_IDinst__n03641_1),
    .ADR2(DLX_IDinst_Ker709161_1),
    .ADR3(DLX_IFinst_NPC[22]),
    .O(DLX_IDinst__n0123[22])
  );
  defparam \DLX_IDinst_Mmux__n0123_Result<31>1 .INIT = 16'hF4B0;
  X_LUT4 \DLX_IDinst_Mmux__n0123_Result<31>1  (
    .ADR0(DLX_IDinst_Ker709161_1),
    .ADR1(DLX_IDinst__n03641_1),
    .ADR2(DLX_IDinst_EPC[31]),
    .ADR3(DLX_IFinst_NPC[31]),
    .O(DLX_IDinst__n0123[31])
  );
  defparam \DLX_IDinst_Mmux__n0123_Result<30>1 .INIT = 16'hF4B0;
  X_LUT4 \DLX_IDinst_Mmux__n0123_Result<30>1  (
    .ADR0(DLX_IDinst_Ker709161_1),
    .ADR1(DLX_IDinst__n03641_1),
    .ADR2(DLX_IDinst_EPC[30]),
    .ADR3(DLX_IFinst_NPC[30]),
    .O(DLX_IDinst__n0123[30])
  );
  defparam \DLX_IDinst_Mmux__n0123_Result<17>1 .INIT = 16'hE2F0;
  X_LUT4 \DLX_IDinst_Mmux__n0123_Result<17>1  (
    .ADR0(DLX_IFinst_NPC[17]),
    .ADR1(DLX_IDinst_Ker709161_1),
    .ADR2(DLX_IDinst_EPC[17]),
    .ADR3(DLX_IDinst__n03641_1),
    .O(DLX_IDinst__n0123[17])
  );
  defparam \DLX_IDinst_Mmux__n0123_Result<16>1 .INIT = 16'hFB08;
  X_LUT4 \DLX_IDinst_Mmux__n0123_Result<16>1  (
    .ADR0(DLX_IFinst_NPC[16]),
    .ADR1(DLX_IDinst__n03641_1),
    .ADR2(DLX_IDinst_Ker709161_1),
    .ADR3(DLX_IDinst_EPC[16]),
    .O(DLX_IDinst__n0123[16])
  );
  defparam \DLX_IDinst_Mmux__n0123_Result<25>1 .INIT = 16'hF4B0;
  X_LUT4 \DLX_IDinst_Mmux__n0123_Result<25>1  (
    .ADR0(DLX_IDinst_Ker709161_1),
    .ADR1(DLX_IDinst__n03641_1),
    .ADR2(DLX_IDinst_EPC[25]),
    .ADR3(DLX_IFinst_NPC[25]),
    .O(DLX_IDinst__n0123[25])
  );
  defparam \DLX_IDinst_Mmux__n0123_Result<24>1 .INIT = 16'hAACA;
  X_LUT4 \DLX_IDinst_Mmux__n0123_Result<24>1  (
    .ADR0(DLX_IDinst_EPC[24]),
    .ADR1(DLX_IFinst_NPC[24]),
    .ADR2(DLX_IDinst__n03641_1),
    .ADR3(DLX_IDinst_Ker709161_1),
    .O(DLX_IDinst__n0123[24])
  );
  defparam \DLX_IDinst_Mmux__n0123_Result<19>1 .INIT = 16'hEF20;
  X_LUT4 \DLX_IDinst_Mmux__n0123_Result<19>1  (
    .ADR0(DLX_IFinst_NPC[19]),
    .ADR1(DLX_IDinst_Ker709161_1),
    .ADR2(DLX_IDinst__n03641_1),
    .ADR3(DLX_IDinst_EPC[19]),
    .O(DLX_IDinst__n0123[19])
  );
  defparam \DLX_IDinst_Mmux__n0123_Result<18>1 .INIT = 16'hFD20;
  X_LUT4 \DLX_IDinst_Mmux__n0123_Result<18>1  (
    .ADR0(DLX_IDinst__n03641_1),
    .ADR1(DLX_IDinst_Ker709161_1),
    .ADR2(DLX_IFinst_NPC[18]),
    .ADR3(DLX_IDinst_EPC[18]),
    .O(DLX_IDinst__n0123[18])
  );
  defparam \DLX_IDinst_Mmux__n0123_Result<27>1 .INIT = 16'hFB40;
  X_LUT4 \DLX_IDinst_Mmux__n0123_Result<27>1  (
    .ADR0(DLX_IDinst_Ker709161_1),
    .ADR1(DLX_IDinst__n03641_1),
    .ADR2(DLX_IFinst_NPC[27]),
    .ADR3(DLX_IDinst_EPC[27]),
    .O(DLX_IDinst__n0123[27])
  );
  defparam \DLX_IDinst_Mmux__n0123_Result<26>1 .INIT = 16'hF0D8;
  X_LUT4 \DLX_IDinst_Mmux__n0123_Result<26>1  (
    .ADR0(DLX_IDinst__n03641_1),
    .ADR1(DLX_IFinst_NPC[26]),
    .ADR2(DLX_IDinst_EPC[26]),
    .ADR3(DLX_IDinst_Ker709161_1),
    .O(DLX_IDinst__n0123[26])
  );
  defparam \DLX_IDinst_Mmux__n0123_Result<29>1 .INIT = 16'hEF40;
  X_LUT4 \DLX_IDinst_Mmux__n0123_Result<29>1  (
    .ADR0(DLX_IDinst_Ker709161_1),
    .ADR1(DLX_IFinst_NPC[29]),
    .ADR2(DLX_IDinst__n03641_1),
    .ADR3(DLX_IDinst_EPC[29]),
    .O(DLX_IDinst__n0123[29])
  );
  defparam \DLX_IDinst_Mmux__n0123_Result<28>1 .INIT = 16'hE4F0;
  X_LUT4 \DLX_IDinst_Mmux__n0123_Result<28>1  (
    .ADR0(DLX_IDinst_Ker709161_1),
    .ADR1(DLX_IFinst_NPC[28]),
    .ADR2(DLX_IDinst_EPC[28]),
    .ADR3(DLX_IDinst__n03641_1),
    .O(DLX_IDinst__n0123[28])
  );
  defparam \DLX_Mmux_reg_dst_of_EX_Result<1>1 .INIT = 16'hE4E4;
  X_LUT4 \DLX_Mmux_reg_dst_of_EX_Result<1>1  (
    .ADR0(DLX_IDinst_reg_dst),
    .ADR1(DLX_IDinst_rt_addr[1]),
    .ADR2(DLX_IDinst_rd_addr[1]),
    .ADR3(VCC),
    .O(\DLX_reg_dst_of_MEM<1>/FROM )
  );
  defparam \DLX_Mmux_reg_dst_of_EX_Result<0>1 .INIT = 16'hFA50;
  X_LUT4 \DLX_Mmux_reg_dst_of_EX_Result<0>1  (
    .ADR0(DLX_IDinst_reg_dst),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_rt_addr[0]),
    .ADR3(DLX_IDinst_rd_addr[0]),
    .O(\DLX_reg_dst_of_MEM<1>/GROM )
  );
  X_BUF \DLX_reg_dst_of_MEM<1>/XUSED  (
    .I(\DLX_reg_dst_of_MEM<1>/FROM ),
    .O(DLX_reg_dst_of_EX[1])
  );
  X_BUF \DLX_reg_dst_of_MEM<1>/YUSED  (
    .I(\DLX_reg_dst_of_MEM<1>/GROM ),
    .O(DLX_reg_dst_of_EX[0])
  );
  defparam \DLX_Mmux_reg_dst_of_EX_Result<3>1 .INIT = 16'hAACC;
  X_LUT4 \DLX_Mmux_reg_dst_of_EX_Result<3>1  (
    .ADR0(DLX_IDinst_rd_addr[3]),
    .ADR1(DLX_IDinst_rt_addr[3]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_dst),
    .O(\DLX_reg_dst_of_MEM<3>/FROM )
  );
  defparam \DLX_Mmux_reg_dst_of_EX_Result<2>1 .INIT = 16'hDD88;
  X_LUT4 \DLX_Mmux_reg_dst_of_EX_Result<2>1  (
    .ADR0(DLX_IDinst_reg_dst),
    .ADR1(DLX_IDinst_rd_addr[2]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_rt_addr[2]),
    .O(\DLX_reg_dst_of_MEM<3>/GROM )
  );
  X_BUF \DLX_reg_dst_of_MEM<3>/XUSED  (
    .I(\DLX_reg_dst_of_MEM<3>/FROM ),
    .O(DLX_reg_dst_of_EX[3])
  );
  X_BUF \DLX_reg_dst_of_MEM<3>/YUSED  (
    .I(\DLX_reg_dst_of_MEM<3>/GROM ),
    .O(DLX_reg_dst_of_EX[2])
  );
  defparam DLX_IFinst_IR_curr_N36381.INIT = 16'h0005;
  X_LUT4 DLX_IFinst_IR_curr_N36381 (
    .ADR0(DLX_IDinst_stall),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_counter[0]),
    .ADR3(DLX_IDinst_counter[1]),
    .O(\DLX_IDinst_counter<1>/FROM )
  );
  defparam \DLX_IDinst__n0116<1>1 .INIT = 16'hC2C3;
  X_LUT4 \DLX_IDinst__n0116<1>1  (
    .ADR0(DLX_IDinst_intr_slot),
    .ADR1(DLX_IDinst_counter[1]),
    .ADR2(DLX_IDinst_counter[0]),
    .ADR3(N95693),
    .O(DLX_IDinst__n0116[1])
  );
  X_BUF \DLX_IDinst_counter<1>/XUSED  (
    .I(\DLX_IDinst_counter<1>/FROM ),
    .O(DLX_IFinst_IR_curr_N3638)
  );
  defparam DLX_EXinst_ALU_result_9_1_1132.INIT = 1'b0;
  X_FF DLX_EXinst_ALU_result_9_1_1132 (
    .I(\DM_addr_eff<9>/OD ),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DM_addr_eff<9>/OFF/RST ),
    .O(DLX_EXinst_ALU_result_9_1)
  );
  X_OR2 \DM_addr_eff<9>/OFF/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DM_addr_eff<9>/OFF/RST )
  );
  defparam DLX_EXinst__n00091.INIT = 16'h0404;
  X_LUT4 DLX_EXinst__n00091 (
    .ADR0(DLX_IDinst_counter[1]),
    .ADR1(DLX_IDinst_reg_write),
    .ADR2(DLX_IDinst_counter[0]),
    .ADR3(VCC),
    .O(DLX_EXinst__n0009)
  );
  defparam DLX_EXinst__n00121.INIT = 16'h0404;
  X_LUT4 DLX_EXinst__n00121 (
    .ADR0(DLX_IDinst_counter[1]),
    .ADR1(DLX_IDinst_mem_write),
    .ADR2(DLX_IDinst_counter[0]),
    .ADR3(VCC),
    .O(\DLX_EXinst_reg_write_EX/GROM )
  );
  X_BUF \DLX_EXinst_reg_write_EX/YUSED  (
    .I(\DLX_EXinst_reg_write_EX/GROM ),
    .O(DLX_EXinst__n0012)
  );
  defparam \DLX_IDinst_Mmux__n0127_Result<1>1 .INIT = 16'hAACA;
  X_LUT4 \DLX_IDinst_Mmux__n0127_Result<1>1  (
    .ADR0(DLX_IDinst_Cause_Reg[1]),
    .ADR1(DLX_IDinst_IR_function_field_1_1),
    .ADR2(DLX_IDinst__n03641_1),
    .ADR3(DLX_IDinst_Ker709161_1),
    .O(DLX_IDinst__n0127[1])
  );
  defparam \DLX_IDinst_Mmux__n0127_Result<0>1 .INIT = 16'hE2F0;
  X_LUT4 \DLX_IDinst_Mmux__n0127_Result<0>1  (
    .ADR0(DLX_IDinst_IR_function_field_0_1),
    .ADR1(DLX_IDinst_Ker709161_1),
    .ADR2(DLX_IDinst_Cause_Reg[0]),
    .ADR3(DLX_IDinst__n03641_1),
    .O(DLX_IDinst__n0127[0])
  );
  defparam \DLX_IDinst_Mmux__n0127_Result<3>1 .INIT = 16'hB8AA;
  X_LUT4 \DLX_IDinst_Mmux__n0127_Result<3>1  (
    .ADR0(DLX_IDinst_Cause_Reg[3]),
    .ADR1(DLX_IDinst_Ker709161_1),
    .ADR2(DLX_IDinst_IR_function_field_3_1),
    .ADR3(DLX_IDinst__n03641_1),
    .O(DLX_IDinst__n0127[3])
  );
  defparam \DLX_IDinst_Mmux__n0127_Result<2>1 .INIT = 16'hE4F0;
  X_LUT4 \DLX_IDinst_Mmux__n0127_Result<2>1  (
    .ADR0(DLX_IDinst_Ker709161_1),
    .ADR1(DLX_IDinst_IR_function_field_2_1),
    .ADR2(DLX_IDinst_Cause_Reg[2]),
    .ADR3(DLX_IDinst__n03641_1),
    .O(DLX_IDinst__n0127[2])
  );
  defparam \DLX_IDinst_Mmux__n0127_Result<5>1 .INIT = 16'hF0B8;
  X_LUT4 \DLX_IDinst_Mmux__n0127_Result<5>1  (
    .ADR0(\DLX_IDinst_Imm[5] ),
    .ADR1(DLX_IDinst__n03641_1),
    .ADR2(DLX_IDinst_Cause_Reg[5]),
    .ADR3(DLX_IDinst_Ker709161_1),
    .O(DLX_IDinst__n0127[5])
  );
  defparam \DLX_IDinst_Mmux__n0127_Result<4>1 .INIT = 16'hACAA;
  X_LUT4 \DLX_IDinst_Mmux__n0127_Result<4>1  (
    .ADR0(DLX_IDinst_Cause_Reg[4]),
    .ADR1(DLX_IDinst_IR_function_field[4]),
    .ADR2(DLX_IDinst_Ker709161_1),
    .ADR3(DLX_IDinst__n03641_1),
    .O(DLX_IDinst__n0127[4])
  );
  defparam \DLX_IDinst_Mmux__n0127_Result<7>1 .INIT = 16'hCCE4;
  X_LUT4 \DLX_IDinst_Mmux__n0127_Result<7>1  (
    .ADR0(DLX_IDinst__n03641_1),
    .ADR1(DLX_IDinst_Cause_Reg[7]),
    .ADR2(\DLX_IDinst_Imm[7] ),
    .ADR3(DLX_IDinst_Ker709161_1),
    .O(DLX_IDinst__n0127[7])
  );
  defparam \DLX_IDinst_Mmux__n0127_Result<6>1 .INIT = 16'hFB08;
  X_LUT4 \DLX_IDinst_Mmux__n0127_Result<6>1  (
    .ADR0(\DLX_IDinst_Imm[6] ),
    .ADR1(DLX_IDinst__n03641_1),
    .ADR2(DLX_IDinst_Ker709161_1),
    .ADR3(DLX_IDinst_Cause_Reg[6]),
    .O(DLX_IDinst__n0127[6])
  );
  defparam \DLX_IDinst_Mmux__n0127_Result<9>1 .INIT = 16'hCCAC;
  X_LUT4 \DLX_IDinst_Mmux__n0127_Result<9>1  (
    .ADR0(\DLX_IDinst_Imm[9] ),
    .ADR1(DLX_IDinst_Cause_Reg[9]),
    .ADR2(DLX_IDinst__n03641_1),
    .ADR3(DLX_IDinst_Ker709161_1),
    .O(DLX_IDinst__n0127[9])
  );
  defparam \DLX_IDinst_Mmux__n0127_Result<8>1 .INIT = 16'hAAE2;
  X_LUT4 \DLX_IDinst_Mmux__n0127_Result<8>1  (
    .ADR0(DLX_IDinst_Cause_Reg[8]),
    .ADR1(DLX_IDinst__n03641_1),
    .ADR2(\DLX_IDinst_Imm[8] ),
    .ADR3(DLX_IDinst_Ker709161_1),
    .O(DLX_IDinst__n0127[8])
  );
  defparam \DLX_EXinst__n0007<11>1 .INIT = 16'hCC00;
  X_LUT4 \DLX_EXinst__n0007<11>1  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_B[11]),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N66350),
    .O(DLX_EXinst__n0007[11])
  );
  defparam \DLX_EXinst__n0007<10>1 .INIT = 16'hA0A0;
  X_LUT4 \DLX_EXinst__n0007<10>1  (
    .ADR0(DLX_EXinst_N66350),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[10]),
    .ADR3(VCC),
    .O(DLX_EXinst__n0007[10])
  );
  defparam DLX_IDinst__n0105_1133.INIT = 16'hC800;
  X_LUT4 DLX_IDinst__n0105_1133 (
    .ADR0(N90703),
    .ADR1(DLX_IDinst_jtarget[0]),
    .ADR2(DLX_IDinst__n0364),
    .ADR3(DLX_IDinst_N70679),
    .O(\DLX_IDinst_IR_function_field<0>/GROM )
  );
  X_BUF \DLX_IDinst_IR_function_field<0>/YUSED  (
    .I(\DLX_IDinst_IR_function_field<0>/GROM ),
    .O(DLX_IDinst__n0105)
  );
  defparam \DLX_EXinst__n0007<13>1 .INIT = 16'hC0C0;
  X_LUT4 \DLX_EXinst__n0007<13>1  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N66350),
    .ADR2(DLX_IDinst_reg_out_B[13]),
    .ADR3(VCC),
    .O(DLX_EXinst__n0007[13])
  );
  defparam \DLX_EXinst__n0007<12>1 .INIT = 16'h8888;
  X_LUT4 \DLX_EXinst__n0007<12>1  (
    .ADR0(DLX_EXinst_N66350),
    .ADR1(DLX_IDinst_reg_out_B[12]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst__n0007[12])
  );
  defparam vga_top_vga1_vsyncout_1134.INIT = 1'b1;
  X_SFF vga_top_vga1_vsyncout_1134 (
    .I(\vsync/LOGIC_ZERO ),
    .CE(VCC),
    .CLK(clkdiv_vga),
    .SET(GSR),
    .RST(GND),
    .SSET(vga_top_vga1__n0011),
    .SRST(GND),
    .O(vga_top_vga1_vsyncout)
  );
  defparam \DLX_EXinst__n0007<21>1 .INIT = 16'hAA00;
  X_LUT4 \DLX_EXinst__n0007<21>1  (
    .ADR0(DLX_IDinst_reg_out_B[21]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N66271),
    .O(DLX_EXinst__n0007[21])
  );
  defparam \DLX_EXinst__n0007<20>1 .INIT = 16'h8888;
  X_LUT4 \DLX_EXinst__n0007<20>1  (
    .ADR0(DLX_EXinst_N66271),
    .ADR1(DLX_IDinst_reg_out_B[20]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst__n0007[20])
  );
  defparam \DLX_EXinst__n0007<23>1 .INIT = 16'hCC00;
  X_LUT4 \DLX_EXinst__n0007<23>1  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N66271),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[23]),
    .O(DLX_EXinst__n0007[23])
  );
  defparam \DLX_EXinst__n0007<22>1 .INIT = 16'hC0C0;
  X_LUT4 \DLX_EXinst__n0007<22>1  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N66271),
    .ADR2(DLX_IDinst_reg_out_B[22]),
    .ADR3(VCC),
    .O(DLX_EXinst__n0007[22])
  );
  defparam \DLX_EXinst__n0017<14>1 .INIT = 16'hDD88;
  X_LUT4 \DLX_EXinst__n0017<14>1  (
    .ADR0(DLX_EXinst__n0030_1),
    .ADR1(DLX_IDinst_reg_out_B[14]),
    .ADR2(VCC),
    .ADR3(\DLX_IDinst_Imm[14] ),
    .O(\DLX_EXinst_reg_out_B_EX<14>/FROM )
  );
  defparam \DLX_EXinst__n0007<14>1 .INIT = 16'h8888;
  X_LUT4 \DLX_EXinst__n0007<14>1  (
    .ADR0(DLX_IDinst_reg_out_B[14]),
    .ADR1(DLX_EXinst_N66350),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst__n0007[14])
  );
  X_BUF \DLX_EXinst_reg_out_B_EX<14>/XUSED  (
    .I(\DLX_EXinst_reg_out_B_EX<14>/FROM ),
    .O(DLX_EXinst__n0017[14])
  );
  defparam DLX_IDinst__n0104_1135.INIT = 16'hA800;
  X_LUT4 DLX_IDinst__n0104_1135 (
    .ADR0(DLX_IDinst_jtarget[1]),
    .ADR1(N90703),
    .ADR2(DLX_IDinst__n0364),
    .ADR3(DLX_IDinst_N70679),
    .O(\DLX_IDinst_IR_function_field<1>/GROM )
  );
  X_BUF \DLX_IDinst_IR_function_field<1>/YUSED  (
    .I(\DLX_IDinst_IR_function_field<1>/GROM ),
    .O(DLX_IDinst__n0104)
  );
  defparam \DLX_EXinst__n0007<25>1 .INIT = 16'hF000;
  X_LUT4 \DLX_EXinst__n0007<25>1  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[25]),
    .ADR3(DLX_EXinst_N66271),
    .O(DLX_EXinst__n0007[25])
  );
  defparam \DLX_EXinst__n0007<24>1 .INIT = 16'hCC00;
  X_LUT4 \DLX_EXinst__n0007<24>1  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_B[24]),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N66271),
    .O(DLX_EXinst__n0007[24])
  );
  defparam \DLX_EXinst__n0007<17>1 .INIT = 16'hCC00;
  X_LUT4 \DLX_EXinst__n0007<17>1  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N66271),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[17]),
    .O(DLX_EXinst__n0007[17])
  );
  defparam \DLX_EXinst__n0007<16>1 .INIT = 16'h8888;
  X_LUT4 \DLX_EXinst__n0007<16>1  (
    .ADR0(DLX_EXinst_N66271),
    .ADR1(DLX_IDinst_reg_out_B[16]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst__n0007[16])
  );
  defparam \DLX_EXinst__n0007<19>1 .INIT = 16'hF000;
  X_LUT4 \DLX_EXinst__n0007<19>1  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N66271),
    .ADR3(DLX_IDinst_reg_out_B[19]),
    .O(DLX_EXinst__n0007[19])
  );
  defparam \DLX_EXinst__n0007<18>1 .INIT = 16'hF000;
  X_LUT4 \DLX_EXinst__n0007<18>1  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[18]),
    .ADR3(DLX_EXinst_N66271),
    .O(DLX_EXinst__n0007[18])
  );
  defparam \DLX_EXinst__n0007<27>1 .INIT = 16'hA0A0;
  X_LUT4 \DLX_EXinst__n0007<27>1  (
    .ADR0(DLX_IDinst_reg_out_B[27]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N66271),
    .ADR3(VCC),
    .O(DLX_EXinst__n0007[27])
  );
  defparam \DLX_EXinst__n0007<26>1 .INIT = 16'h8888;
  X_LUT4 \DLX_EXinst__n0007<26>1  (
    .ADR0(DLX_EXinst_N66271),
    .ADR1(DLX_IDinst_reg_out_B[26]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst__n0007[26])
  );
  defparam DLX_IDinst__n0103_1136.INIT = 16'h8880;
  X_LUT4 DLX_IDinst__n0103_1136 (
    .ADR0(DLX_IDinst_jtarget[2]),
    .ADR1(DLX_IDinst_N70679),
    .ADR2(N90703),
    .ADR3(DLX_IDinst__n0364),
    .O(\DLX_IDinst_IR_function_field<2>/GROM )
  );
  X_BUF \DLX_IDinst_IR_function_field<2>/YUSED  (
    .I(\DLX_IDinst_IR_function_field<2>/GROM ),
    .O(DLX_IDinst__n0103)
  );
  defparam \DLX_EXinst__n0007<29>1 .INIT = 16'hA0A0;
  X_LUT4 \DLX_EXinst__n0007<29>1  (
    .ADR0(DLX_EXinst_N66271),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[29]),
    .ADR3(VCC),
    .O(DLX_EXinst__n0007[29])
  );
  defparam \DLX_EXinst__n0007<28>1 .INIT = 16'h8888;
  X_LUT4 \DLX_EXinst__n0007<28>1  (
    .ADR0(DLX_EXinst_N66271),
    .ADR1(DLX_IDinst_reg_out_B[28]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst__n0007[28])
  );
  defparam DLX_IDinst__n0102_1137.INIT = 16'hE000;
  X_LUT4 DLX_IDinst__n0102_1137 (
    .ADR0(N90703),
    .ADR1(DLX_IDinst__n0364),
    .ADR2(DLX_IDinst_jtarget[3]),
    .ADR3(DLX_IDinst_N70679),
    .O(\DLX_IDinst_IR_function_field<3>/GROM )
  );
  X_BUF \DLX_IDinst_IR_function_field<3>/YUSED  (
    .I(\DLX_IDinst_IR_function_field<3>/GROM ),
    .O(DLX_IDinst__n0102)
  );
  defparam \DLX_IDinst__n0118<11>1 .INIT = 16'hCC00;
  X_LUT4 \DLX_IDinst__n0118<11>1  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_regB_eff[11]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_N69711),
    .O(DLX_IDinst__n0118[11])
  );
  defparam \DLX_IDinst__n0118<10>1 .INIT = 16'hF000;
  X_LUT4 \DLX_IDinst__n0118<10>1  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_N69711),
    .ADR3(DLX_IDinst_regB_eff[10]),
    .O(DLX_IDinst__n0118[10])
  );
  defparam \DLX_IDinst__n0118<21>1 .INIT = 16'hA0A0;
  X_LUT4 \DLX_IDinst__n0118<21>1  (
    .ADR0(DLX_IDinst_regB_eff[21]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_N69711),
    .ADR3(VCC),
    .O(DLX_IDinst__n0118[21])
  );
  defparam \DLX_IDinst__n0118<20>1 .INIT = 16'hC0C0;
  X_LUT4 \DLX_IDinst__n0118<20>1  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_regB_eff[20]),
    .ADR2(DLX_IDinst_N69711),
    .ADR3(VCC),
    .O(DLX_IDinst__n0118[20])
  );
  defparam \DLX_IDinst__n0118<13>1 .INIT = 16'h8888;
  X_LUT4 \DLX_IDinst__n0118<13>1  (
    .ADR0(DLX_IDinst_regB_eff[13]),
    .ADR1(DLX_IDinst_N69711),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst__n0118[13])
  );
  defparam \DLX_IDinst__n0118<12>1 .INIT = 16'h8888;
  X_LUT4 \DLX_IDinst__n0118<12>1  (
    .ADR0(DLX_IDinst_regB_eff[12]),
    .ADR1(DLX_IDinst_N69711),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst__n0118[12])
  );
  defparam \DLX_IDinst__n0118<31>1 .INIT = 16'h8888;
  X_LUT4 \DLX_IDinst__n0118<31>1  (
    .ADR0(DLX_IDinst_N69711),
    .ADR1(DLX_IDinst_regB_eff[31]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst__n0118[31])
  );
  defparam \DLX_IDinst__n0118<30>1 .INIT = 16'h8888;
  X_LUT4 \DLX_IDinst__n0118<30>1  (
    .ADR0(DLX_IDinst_N69711),
    .ADR1(DLX_IDinst_regB_eff[30]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst__n0118[30])
  );
  defparam \DLX_IDinst__n0118<23>1 .INIT = 16'hF000;
  X_LUT4 \DLX_IDinst__n0118<23>1  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_N69711),
    .ADR3(DLX_IDinst_regB_eff[23]),
    .O(DLX_IDinst__n0118[23])
  );
  defparam \DLX_IDinst__n0118<22>1 .INIT = 16'hF000;
  X_LUT4 \DLX_IDinst__n0118<22>1  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_N69711),
    .ADR3(DLX_IDinst_regB_eff[22]),
    .O(DLX_IDinst__n0118[22])
  );
  defparam \DLX_IDinst__n0118<15>1 .INIT = 16'hA0A0;
  X_LUT4 \DLX_IDinst__n0118<15>1  (
    .ADR0(DLX_IDinst_N69711),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_regB_eff[15]),
    .ADR3(VCC),
    .O(DLX_IDinst__n0118[15])
  );
  defparam \DLX_IDinst__n0118<14>1 .INIT = 16'hAA00;
  X_LUT4 \DLX_IDinst__n0118<14>1  (
    .ADR0(DLX_IDinst_N69711),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_regB_eff[14]),
    .O(DLX_IDinst__n0118[14])
  );
  defparam \DLX_IDinst__n0118<25>1 .INIT = 16'hC0C0;
  X_LUT4 \DLX_IDinst__n0118<25>1  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_regB_eff[25]),
    .ADR2(DLX_IDinst_N69711),
    .ADR3(VCC),
    .O(DLX_IDinst__n0118[25])
  );
  defparam \DLX_IDinst__n0118<24>1 .INIT = 16'hA0A0;
  X_LUT4 \DLX_IDinst__n0118<24>1  (
    .ADR0(DLX_IDinst_regB_eff[24]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_N69711),
    .ADR3(VCC),
    .O(DLX_IDinst__n0118[24])
  );
  defparam \DLX_IDinst__n0118<17>1 .INIT = 16'hCC00;
  X_LUT4 \DLX_IDinst__n0118<17>1  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_N69711),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_regB_eff[17]),
    .O(DLX_IDinst__n0118[17])
  );
  defparam \DLX_IDinst__n0118<16>1 .INIT = 16'hAA00;
  X_LUT4 \DLX_IDinst__n0118<16>1  (
    .ADR0(DLX_IDinst_regB_eff[16]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_N69711),
    .O(DLX_IDinst__n0118[16])
  );
  defparam \DLX_IDinst__n0118<27>1 .INIT = 16'hA0A0;
  X_LUT4 \DLX_IDinst__n0118<27>1  (
    .ADR0(DLX_IDinst_regB_eff[27]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_N69711),
    .ADR3(VCC),
    .O(DLX_IDinst__n0118[27])
  );
  defparam \DLX_IDinst__n0118<26>1 .INIT = 16'hC0C0;
  X_LUT4 \DLX_IDinst__n0118<26>1  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_regB_eff[26]),
    .ADR2(DLX_IDinst_N69711),
    .ADR3(VCC),
    .O(DLX_IDinst__n0118[26])
  );
  defparam \DLX_IDinst__n0118<19>1 .INIT = 16'h8888;
  X_LUT4 \DLX_IDinst__n0118<19>1  (
    .ADR0(DLX_IDinst_N69711),
    .ADR1(DLX_IDinst_regB_eff[19]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst__n0118[19])
  );
  defparam \DLX_IDinst__n0118<18>1 .INIT = 16'hAA00;
  X_LUT4 \DLX_IDinst__n0118<18>1  (
    .ADR0(DLX_IDinst_N69711),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_regB_eff[18]),
    .O(DLX_IDinst__n0118[18])
  );
  defparam \DLX_IDinst__n0118<29>1 .INIT = 16'h8888;
  X_LUT4 \DLX_IDinst__n0118<29>1  (
    .ADR0(DLX_IDinst_N69711),
    .ADR1(DLX_IDinst_regB_eff[29]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst__n0118[29])
  );
  defparam \DLX_IDinst__n0118<28>1 .INIT = 16'hA0A0;
  X_LUT4 \DLX_IDinst__n0118<28>1  (
    .ADR0(DLX_IDinst_N69711),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_regB_eff[28]),
    .ADR3(VCC),
    .O(DLX_IDinst__n0118[28])
  );
  defparam DLX_EXinst_Ker63687_SW1.INIT = 16'h8000;
  X_LUT4 DLX_EXinst_Ker63687_SW1 (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(DLX_EXinst_N66078),
    .ADR2(DLX_IDinst_reg_out_B[5]),
    .ADR3(DLX_EXinst__n0149),
    .O(\DLX_EXinst_ALU_result<2>/FROM )
  );
  defparam \DLX_EXinst__n0006<2>412 .INIT = 16'hFAEA;
  X_LUT4 \DLX_EXinst__n0006<2>412  (
    .ADR0(DLX_EXinst_N63689),
    .ADR1(CHOICE5522),
    .ADR2(DLX_EXinst__n0149),
    .ADR3(CHOICE5567),
    .O(\DLX_EXinst_ALU_result<2>/GROM )
  );
  X_BUF \DLX_EXinst_ALU_result<2>/XUSED  (
    .I(\DLX_EXinst_ALU_result<2>/FROM ),
    .O(N101921)
  );
  X_BUF \DLX_EXinst_ALU_result<2>/YUSED  (
    .I(\DLX_EXinst_ALU_result<2>/GROM ),
    .O(N123038)
  );
  defparam \DLX_IDinst__n0113<2> .INIT = 16'hA080;
  X_LUT4 \DLX_IDinst__n0113<2>  (
    .ADR0(DLX_IDinst_N70679),
    .ADR1(DLX_IDinst__n0364),
    .ADR2(DLX_IDinst_IR_latched[28]),
    .ADR3(N90703),
    .O(DLX_IDinst__n0113[2])
  );
  defparam DLX_IDinst__n0099_1138.INIT = 16'hA080;
  X_LUT4 DLX_IDinst__n0099_1138 (
    .ADR0(DLX_IDinst_N70679),
    .ADR1(N90703),
    .ADR2(DLX_IDinst_jtarget[6]),
    .ADR3(DLX_IDinst__n0364),
    .O(DLX_IDinst__n0099)
  );
  defparam DLX_IDinst__n0097_1139.INIT = 16'hC800;
  X_LUT4 DLX_IDinst__n0097_1139 (
    .ADR0(DLX_IDinst__n0364),
    .ADR1(DLX_IDinst_jtarget[8]),
    .ADR2(N90703),
    .ADR3(DLX_IDinst_N70679),
    .O(DLX_IDinst__n0097)
  );
  defparam DLX_IDinst__n0098_1140.INIT = 16'h8880;
  X_LUT4 DLX_IDinst__n0098_1140 (
    .ADR0(DLX_IDinst_jtarget[7]),
    .ADR1(DLX_IDinst_N70679),
    .ADR2(N90703),
    .ADR3(DLX_IDinst__n0364),
    .O(DLX_IDinst__n0098)
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<1>1 .INIT = 16'hCCF0;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<1>1  (
    .ADR0(VCC),
    .ADR1(DM_read_data[1]),
    .ADR2(DLX_EXinst_ALU_result[1]),
    .ADR3(DLX_EXinst_mem_to_reg_EX),
    .O(DLX_MEMinst__n0000[1])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<0>1 .INIT = 16'hACAC;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<0>1  (
    .ADR0(DM_read_data[0]),
    .ADR1(DLX_EXinst_ALU_result[0]),
    .ADR2(DLX_EXinst_mem_to_reg_EX),
    .ADR3(VCC),
    .O(DLX_MEMinst__n0000[0])
  );
  X_INV \DLX_RF_data_in<1>/CKINV  (
    .I(DLX_MEMlc_master_ctrlMEM_l),
    .O(\DLX_RF_data_in<1>/CKMUXNOT )
  );
  defparam DLX_IDinst__n0095_1141.INIT = 16'hC080;
  X_LUT4 DLX_IDinst__n0095_1141 (
    .ADR0(DLX_IDinst__n0364),
    .ADR1(DLX_IDinst_jtarget[10]),
    .ADR2(DLX_IDinst_N70679),
    .ADR3(N90703),
    .O(DLX_IDinst__n0095)
  );
  defparam DLX_IDinst__n0096_1142.INIT = 16'hA800;
  X_LUT4 DLX_IDinst__n0096_1142 (
    .ADR0(DLX_IDinst_N70679),
    .ADR1(DLX_IDinst__n0364),
    .ADR2(N90703),
    .ADR3(DLX_IDinst_jtarget[9]),
    .O(DLX_IDinst__n0096)
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<3>1 .INIT = 16'hCACA;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<3>1  (
    .ADR0(DLX_EXinst_ALU_result[3]),
    .ADR1(DM_read_data[3]),
    .ADR2(DLX_EXinst_mem_to_reg_EX),
    .ADR3(VCC),
    .O(DLX_MEMinst__n0000[3])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<2>1 .INIT = 16'hAACC;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<2>1  (
    .ADR0(DM_read_data[2]),
    .ADR1(DLX_EXinst_ALU_result[2]),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_mem_to_reg_EX),
    .O(DLX_MEMinst__n0000[2])
  );
  X_INV \DLX_RF_data_in<3>/CKINV  (
    .I(DLX_MEMlc_master_ctrlMEM_l),
    .O(\DLX_RF_data_in<3>/CKMUXNOT )
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<5>1 .INIT = 16'hAAF0;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<5>1  (
    .ADR0(DM_read_data[5]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_ALU_result[5]),
    .ADR3(DLX_EXinst_mem_to_reg_EX),
    .O(DLX_MEMinst__n0000[5])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<4>1 .INIT = 16'hCFC0;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<4>1  (
    .ADR0(VCC),
    .ADR1(DM_read_data[4]),
    .ADR2(DLX_EXinst_mem_to_reg_EX),
    .ADR3(DLX_EXinst_ALU_result[4]),
    .O(DLX_MEMinst__n0000[4])
  );
  X_INV \DLX_RF_data_in<5>/CKINV  (
    .I(DLX_MEMlc_master_ctrlMEM_l),
    .O(\DLX_RF_data_in<5>/CKMUXNOT )
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<7>1 .INIT = 16'hCFC0;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<7>1  (
    .ADR0(VCC),
    .ADR1(DM_read_data[7]),
    .ADR2(DLX_EXinst_mem_to_reg_EX),
    .ADR3(DLX_EXinst_ALU_result[7]),
    .O(DLX_MEMinst__n0000[7])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<6>1 .INIT = 16'hFA50;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<6>1  (
    .ADR0(DLX_EXinst_mem_to_reg_EX),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_ALU_result[6]),
    .ADR3(DM_read_data[6]),
    .O(DLX_MEMinst__n0000[6])
  );
  X_INV \DLX_RF_data_in<7>/CKINV  (
    .I(DLX_MEMlc_master_ctrlMEM_l),
    .O(\DLX_RF_data_in<7>/CKMUXNOT )
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<9>1 .INIT = 16'hAACC;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<9>1  (
    .ADR0(DM_read_data[9]),
    .ADR1(DLX_EXinst_ALU_result[9]),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_mem_to_reg_EX),
    .O(DLX_MEMinst__n0000[9])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<8>1 .INIT = 16'hAFA0;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<8>1  (
    .ADR0(DM_read_data[8]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_mem_to_reg_EX),
    .ADR3(DLX_EXinst_ALU_result[8]),
    .O(DLX_MEMinst__n0000[8])
  );
  X_INV \DLX_MEMinst_RF_data_in<9>/CKINV  (
    .I(DLX_MEMlc_master_ctrlMEM_l),
    .O(\DLX_MEMinst_RF_data_in<9>/CKMUXNOT )
  );
  X_OR2 \DLX_IDinst_IR_opcode_field<5>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_IR_opcode_field<5>/FFY/RST )
  );
  defparam DLX_IDinst_IR_opcode_field_0.INIT = 1'b0;
  X_FF DLX_IDinst_IR_opcode_field_0 (
    .I(DLX_IDinst__n0113[0]),
    .CE(DLX_IDinst__n0422),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_IR_opcode_field<5>/FFY/RST ),
    .O(DLX_IDinst_IR_opcode_field[0])
  );
  defparam \DLX_IDinst__n0113<5> .INIT = 16'hC080;
  X_LUT4 \DLX_IDinst__n0113<5>  (
    .ADR0(N91278),
    .ADR1(DLX_IDinst_N70679),
    .ADR2(DLX_IDinst_IR_latched[31]),
    .ADR3(DLX_IDinst__n0364),
    .O(DLX_IDinst__n0113[5])
  );
  defparam \DLX_IDinst__n0113<0> .INIT = 16'hA080;
  X_LUT4 \DLX_IDinst__n0113<0>  (
    .ADR0(DLX_IDinst_N70679),
    .ADR1(N90703),
    .ADR2(DLX_IDinst_IR_latched[26]),
    .ADR3(DLX_IDinst__n0364),
    .O(DLX_IDinst__n0113[0])
  );
  defparam DLX_EXinst__n00151.INIT = 16'h20A0;
  X_LUT4 DLX_EXinst__n00151 (
    .ADR0(DLX_EXinst_N66130),
    .ADR1(DLX_IDinst_IR_opcode_field[2]),
    .ADR2(DLX_IDinst_IR_opcode_field[0]),
    .ADR3(DLX_IDinst_IR_opcode_field[3]),
    .O(DLX_EXinst__n0015)
  );
  defparam DLX_EXinst__n00141.INIT = 16'h0070;
  X_LUT4 DLX_EXinst__n00141 (
    .ADR0(DLX_IDinst_IR_opcode_field[2]),
    .ADR1(DLX_IDinst_IR_opcode_field[3]),
    .ADR2(DLX_EXinst_N66130),
    .ADR3(DLX_IDinst_IR_opcode_field[0]),
    .O(DLX_EXinst__n0014)
  );
  X_OR2 \DLX_IDinst_intr_slot/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_intr_slot/FFY/RST )
  );
  defparam DLX_IDinst_intr_slot_1143.INIT = 1'b0;
  X_FF DLX_IDinst_intr_slot_1143 (
    .I(DLX_IDinst__n0126),
    .CE(DLX_IDinst__n0443),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_intr_slot/FFY/RST ),
    .O(DLX_IDinst_intr_slot)
  );
  defparam DLX_IDinst__n03101.INIT = 16'h5000;
  X_LUT4 DLX_IDinst__n03101 (
    .ADR0(DLX_IDinst__n0331),
    .ADR1(VCC),
    .ADR2(DLX_IDinst__n0387),
    .ADR3(DLX_IDinst_N70918),
    .O(\DLX_IDinst_intr_slot/FROM )
  );
  defparam DLX_IDinst__n01261.INIT = 16'h0032;
  X_LUT4 DLX_IDinst__n01261 (
    .ADR0(DLX_IDinst__n03641_1),
    .ADR1(DLX_IDinst__n0331),
    .ADR2(DLX_IDinst__n0071),
    .ADR3(DLX_IDinst_N70918),
    .O(DLX_IDinst__n0126)
  );
  X_BUF \DLX_IDinst_intr_slot/XUSED  (
    .I(\DLX_IDinst_intr_slot/FROM ),
    .O(DLX_IDinst__n0310)
  );
  defparam DLX_IFinst_PC_ClkEn_INV1.INIT = 16'h0001;
  X_LUT4 DLX_IFinst_PC_ClkEn_INV1 (
    .ADR0(DLX_IDinst_stall),
    .ADR1(DLX_IDinst_counter[1]),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(DLX_IDinst_counter[0]),
    .O(\DLX_IFinst_stalled/FROM )
  );
  defparam DLX_IFinst__n00001.INIT = 16'hFFFC;
  X_LUT4 DLX_IFinst__n00001 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_stall),
    .ADR2(DLX_IDinst_counter[0]),
    .ADR3(DLX_IDinst_counter[1]),
    .O(\DLX_IFinst_stalled/GROM )
  );
  X_INV \DLX_IFinst_stalled/CEMUX  (
    .I(DLX_IDinst_branch_sig),
    .O(\DLX_IFinst_stalled/CEMUXNOT )
  );
  X_BUF \DLX_IFinst_stalled/XUSED  (
    .I(\DLX_IFinst_stalled/FROM ),
    .O(DLX_IFinst_PC_N3535)
  );
  X_BUF \DLX_IFinst_stalled/YUSED  (
    .I(\DLX_IFinst_stalled/GROM ),
    .O(DLX_IFinst__n0000)
  );
  defparam \DLX_IDinst__n0107<4>1 .INIT = 16'h00FC;
  X_LUT4 \DLX_IDinst__n0107<4>1  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst__n0023[4]),
    .ADR2(DLX_IDinst_N70918),
    .ADR3(DLX_IDinst__n0331),
    .O(DLX_IDinst__n0107[4])
  );
  defparam \DLX_IDinst__n0107<1>1 .INIT = 16'h3322;
  X_LUT4 \DLX_IDinst__n0107<1>1  (
    .ADR0(DLX_IDinst__n0023[1]),
    .ADR1(DLX_IDinst__n0331),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_N70918),
    .O(DLX_IDinst__n0107[1])
  );
  defparam \DLX_IDinst__n0107<3>1 .INIT = 16'h00FA;
  X_LUT4 \DLX_IDinst__n0107<3>1  (
    .ADR0(DLX_IDinst__n0023[3]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_N70918),
    .ADR3(DLX_IDinst__n0331),
    .O(DLX_IDinst__n0107[3])
  );
  defparam \DLX_IDinst__n0107<2>1 .INIT = 16'h00FA;
  X_LUT4 \DLX_IDinst__n0107<2>1  (
    .ADR0(DLX_IDinst__n0023[2]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_N70918),
    .ADR3(DLX_IDinst__n0331),
    .O(DLX_IDinst__n0107[2])
  );
  defparam \DLX_IDinst__n0118<1>1 .INIT = 16'hC0C0;
  X_LUT4 \DLX_IDinst__n0118<1>1  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_regB_eff[1]),
    .ADR2(DLX_IDinst_N69711),
    .ADR3(VCC),
    .O(DLX_IDinst__n0118[1])
  );
  defparam \DLX_IDinst__n0118<5>1 .INIT = 16'hA0A0;
  X_LUT4 \DLX_IDinst__n0118<5>1  (
    .ADR0(DLX_IDinst_N69711),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_regB_eff[5]),
    .ADR3(VCC),
    .O(DLX_IDinst__n0118[5])
  );
  defparam \DLX_IDinst__n0118<4>1 .INIT = 16'h8888;
  X_LUT4 \DLX_IDinst__n0118<4>1  (
    .ADR0(DLX_IDinst_regB_eff[4]),
    .ADR1(DLX_IDinst_N69711),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst__n0118[4])
  );
  defparam \DLX_IDinst__n0118<7>1 .INIT = 16'h8888;
  X_LUT4 \DLX_IDinst__n0118<7>1  (
    .ADR0(DLX_IDinst_regB_eff[7]),
    .ADR1(DLX_IDinst_N69711),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst__n0118[7])
  );
  defparam \DLX_IDinst__n0118<6>1 .INIT = 16'hCC00;
  X_LUT4 \DLX_IDinst__n0118<6>1  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_N69711),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_regB_eff[6]),
    .O(DLX_IDinst__n0118[6])
  );
  defparam \DLX_IDinst__n0118<9>1 .INIT = 16'hAA00;
  X_LUT4 \DLX_IDinst__n0118<9>1  (
    .ADR0(DLX_IDinst_N69711),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_regB_eff[9]),
    .O(DLX_IDinst__n0118[9])
  );
  defparam \DLX_IDinst__n0118<8>1 .INIT = 16'hA0A0;
  X_LUT4 \DLX_IDinst__n0118<8>1  (
    .ADR0(DLX_IDinst_N69711),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_regB_eff[8]),
    .ADR3(VCC),
    .O(DLX_IDinst__n0118[8])
  );
  defparam DLX_IDinst__n0108144.INIT = 16'hDDCC;
  X_LUT4 DLX_IDinst__n0108144 (
    .ADR0(DLX_IDinst__n0364),
    .ADR1(DLX_IDinst_N70918),
    .ADR2(VCC),
    .ADR3(DLX_IDinst__n0071),
    .O(\DLX_IDinst_rt_addr<1>/FROM )
  );
  defparam \DLX_IDinst__n0106<1> .INIT = 16'hA800;
  X_LUT4 \DLX_IDinst__n0106<1>  (
    .ADR0(DLX_IDinst_regB_index[1]),
    .ADR1(DLX_IDinst__n0364),
    .ADR2(N90703),
    .ADR3(DLX_IDinst_N70679),
    .O(DLX_IDinst__n0106[1])
  );
  X_BUF \DLX_IDinst_rt_addr<1>/XUSED  (
    .I(\DLX_IDinst_rt_addr<1>/FROM ),
    .O(CHOICE3460)
  );
  defparam \DLX_IDinst__n0106<3> .INIT = 16'hE000;
  X_LUT4 \DLX_IDinst__n0106<3>  (
    .ADR0(N90703),
    .ADR1(DLX_IDinst__n0364),
    .ADR2(DLX_IDinst_regB_index[3]),
    .ADR3(DLX_IDinst_N70679),
    .O(DLX_IDinst__n0106[3])
  );
  defparam \DLX_IDinst__n0106<2> .INIT = 16'hE000;
  X_LUT4 \DLX_IDinst__n0106<2>  (
    .ADR0(N90703),
    .ADR1(DLX_IDinst__n0364),
    .ADR2(DLX_IDinst_regB_index[2]),
    .ADR3(DLX_IDinst_N70679),
    .O(DLX_IDinst__n0106[2])
  );
  defparam DLX_IDinst__n0110_SW0.INIT = 16'hF077;
  X_LUT4 DLX_IDinst__n0110_SW0 (
    .ADR0(N102532),
    .ADR1(DLX_IDinst_N69568),
    .ADR2(DLX_IDinst__n0448[1]),
    .ADR3(DLX_IDinst__n0364),
    .O(\DLX_IDinst_mem_read/FROM )
  );
  defparam DLX_IDinst__n0111_1144.INIT = 16'h8000;
  X_LUT4 DLX_IDinst__n0111_1144 (
    .ADR0(N102532),
    .ADR1(DLX_IDinst__n0133),
    .ADR2(N90322),
    .ADR3(DLX_IDinst__n0132),
    .O(DLX_IDinst__n0111)
  );
  X_BUF \DLX_IDinst_mem_read/XUSED  (
    .I(\DLX_IDinst_mem_read/FROM ),
    .O(N100496)
  );
  defparam \DLX_IDinst_Mmux__n0127_Result<11>1 .INIT = 16'hAACA;
  X_LUT4 \DLX_IDinst_Mmux__n0127_Result<11>1  (
    .ADR0(DLX_IDinst_Cause_Reg[11]),
    .ADR1(\DLX_IDinst_Imm[11] ),
    .ADR2(DLX_IDinst__n03641_1),
    .ADR3(DLX_IDinst_Ker709161_1),
    .O(DLX_IDinst__n0127[11])
  );
  defparam \DLX_IDinst_Mmux__n0127_Result<10>1 .INIT = 16'hFD20;
  X_LUT4 \DLX_IDinst_Mmux__n0127_Result<10>1  (
    .ADR0(DLX_IDinst__n03641_1),
    .ADR1(DLX_IDinst_Ker709161_1),
    .ADR2(\DLX_IDinst_Imm[10] ),
    .ADR3(DLX_IDinst_Cause_Reg[10]),
    .O(DLX_IDinst__n0127[10])
  );
  defparam \DLX_IDinst_Mmux__n0127_Result<13>1 .INIT = 16'hFD08;
  X_LUT4 \DLX_IDinst_Mmux__n0127_Result<13>1  (
    .ADR0(DLX_IDinst__n03641_1),
    .ADR1(\DLX_IDinst_Imm[13] ),
    .ADR2(DLX_IDinst_Ker709161_1),
    .ADR3(DLX_IDinst_Cause_Reg[13]),
    .O(DLX_IDinst__n0127[13])
  );
  defparam \DLX_IDinst_Mmux__n0127_Result<12>1 .INIT = 16'hF4B0;
  X_LUT4 \DLX_IDinst_Mmux__n0127_Result<12>1  (
    .ADR0(DLX_IDinst_Ker709161_1),
    .ADR1(DLX_IDinst__n03641_1),
    .ADR2(DLX_IDinst_Cause_Reg[12]),
    .ADR3(\DLX_IDinst_Imm[12] ),
    .O(DLX_IDinst__n0127[12])
  );
  defparam \DLX_IDinst_Mmux__n0127_Result<21>1 .INIT = 16'hFD08;
  X_LUT4 \DLX_IDinst_Mmux__n0127_Result<21>1  (
    .ADR0(DLX_IDinst__n03641_1),
    .ADR1(DLX_IDinst_Imm_31_1),
    .ADR2(DLX_IDinst_Ker709161_1),
    .ADR3(DLX_IDinst_Cause_Reg[21]),
    .O(DLX_IDinst__n0127[21])
  );
  defparam \DLX_IDinst_Mmux__n0127_Result<20>1 .INIT = 16'hCCAC;
  X_LUT4 \DLX_IDinst_Mmux__n0127_Result<20>1  (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(DLX_IDinst_Cause_Reg[20]),
    .ADR2(DLX_IDinst__n03641_1),
    .ADR3(DLX_IDinst_Ker709161_1),
    .O(DLX_IDinst__n0127[20])
  );
  defparam DLX_IDinst_Ker6963328_SW0.INIT = 16'h77FF;
  X_LUT4 DLX_IDinst_Ker6963328_SW0 (
    .ADR0(DLX_IDinst_IR_latched[26]),
    .ADR1(DLX_IDinst_N70673),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_IR_latched[31]),
    .O(\DLX_IDinst_mem_write/FROM )
  );
  defparam DLX_IDinst__n0112_1145.INIT = 16'h2000;
  X_LUT4 DLX_IDinst__n0112_1145 (
    .ADR0(DLX_IDinst_N70821),
    .ADR1(N100243),
    .ADR2(DLX_IDinst_IR_latched[31]),
    .ADR3(DLX_IDinst_N70679),
    .O(DLX_IDinst__n0112)
  );
  X_BUF \DLX_IDinst_mem_write/XUSED  (
    .I(\DLX_IDinst_mem_write/FROM ),
    .O(N127551)
  );
  defparam \DLX_IDinst_Mmux__n0127_Result<15>1 .INIT = 16'hCCAC;
  X_LUT4 \DLX_IDinst_Mmux__n0127_Result<15>1  (
    .ADR0(\DLX_IDinst_Imm[15] ),
    .ADR1(DLX_IDinst_Cause_Reg[15]),
    .ADR2(DLX_IDinst__n03641_1),
    .ADR3(DLX_IDinst_Ker709161_1),
    .O(DLX_IDinst__n0127[15])
  );
  defparam \DLX_IDinst_Mmux__n0127_Result<14>1 .INIT = 16'hFD08;
  X_LUT4 \DLX_IDinst_Mmux__n0127_Result<14>1  (
    .ADR0(DLX_IDinst__n03641_1),
    .ADR1(\DLX_IDinst_Imm[14] ),
    .ADR2(DLX_IDinst_Ker709161_1),
    .ADR3(DLX_IDinst_Cause_Reg[14]),
    .O(DLX_IDinst__n0127[14])
  );
  defparam \DLX_IDinst_Mmux__n0127_Result<23>1 .INIT = 16'hAEA2;
  X_LUT4 \DLX_IDinst_Mmux__n0127_Result<23>1  (
    .ADR0(DLX_IDinst_Cause_Reg[23]),
    .ADR1(DLX_IDinst__n03641_1),
    .ADR2(DLX_IDinst_Ker709161_1),
    .ADR3(DLX_IDinst_Imm_31_1),
    .O(DLX_IDinst__n0127[23])
  );
  defparam \DLX_IDinst_Mmux__n0127_Result<22>1 .INIT = 16'hCACC;
  X_LUT4 \DLX_IDinst_Mmux__n0127_Result<22>1  (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(DLX_IDinst_Cause_Reg[22]),
    .ADR2(DLX_IDinst_Ker709161_1),
    .ADR3(DLX_IDinst__n03641_1),
    .O(DLX_IDinst__n0127[22])
  );
  defparam \DLX_IDinst_Mmux__n0127_Result<31>1 .INIT = 16'hF0B8;
  X_LUT4 \DLX_IDinst_Mmux__n0127_Result<31>1  (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(DLX_IDinst__n03641_1),
    .ADR2(DLX_IDinst_Cause_Reg[31]),
    .ADR3(DLX_IDinst_Ker709161_1),
    .O(DLX_IDinst__n0127[31])
  );
  defparam \DLX_IDinst_Mmux__n0127_Result<30>1 .INIT = 16'hF2D0;
  X_LUT4 \DLX_IDinst_Mmux__n0127_Result<30>1  (
    .ADR0(DLX_IDinst__n03641_1),
    .ADR1(DLX_IDinst_Ker709161_1),
    .ADR2(DLX_IDinst_Cause_Reg[30]),
    .ADR3(DLX_IDinst_Imm_31_1),
    .O(DLX_IDinst__n0127[30])
  );
  defparam \DLX_IDinst_Mmux__n0127_Result<17>1 .INIT = 16'hF0D8;
  X_LUT4 \DLX_IDinst_Mmux__n0127_Result<17>1  (
    .ADR0(DLX_IDinst__n03641_1),
    .ADR1(DLX_IDinst_Imm_31_1),
    .ADR2(DLX_IDinst_Cause_Reg[17]),
    .ADR3(DLX_IDinst_Ker709161_1),
    .O(DLX_IDinst__n0127[17])
  );
  defparam \DLX_IDinst_Mmux__n0127_Result<16>1 .INIT = 16'hEF40;
  X_LUT4 \DLX_IDinst_Mmux__n0127_Result<16>1  (
    .ADR0(DLX_IDinst_Ker709161_1),
    .ADR1(DLX_IDinst_Imm_31_1),
    .ADR2(DLX_IDinst__n03641_1),
    .ADR3(DLX_IDinst_Cause_Reg[16]),
    .O(DLX_IDinst__n0127[16])
  );
  defparam \DLX_IDinst_Mmux__n0127_Result<25>1 .INIT = 16'hBA8A;
  X_LUT4 \DLX_IDinst_Mmux__n0127_Result<25>1  (
    .ADR0(DLX_IDinst_Cause_Reg[25]),
    .ADR1(DLX_IDinst_Ker709161_1),
    .ADR2(DLX_IDinst__n03641_1),
    .ADR3(DLX_IDinst_Imm_31_1),
    .O(DLX_IDinst__n0127[25])
  );
  defparam \DLX_IDinst_Mmux__n0127_Result<24>1 .INIT = 16'hB8AA;
  X_LUT4 \DLX_IDinst_Mmux__n0127_Result<24>1  (
    .ADR0(DLX_IDinst_Cause_Reg[24]),
    .ADR1(DLX_IDinst_Ker709161_1),
    .ADR2(DLX_IDinst_Imm_31_1),
    .ADR3(DLX_IDinst__n03641_1),
    .O(DLX_IDinst__n0127[24])
  );
  defparam \DLX_IDinst_Mmux__n0127_Result<19>1 .INIT = 16'hCCE4;
  X_LUT4 \DLX_IDinst_Mmux__n0127_Result<19>1  (
    .ADR0(DLX_IDinst__n03641_1),
    .ADR1(DLX_IDinst_Cause_Reg[19]),
    .ADR2(DLX_IDinst_Imm_31_1),
    .ADR3(DLX_IDinst_Ker709161_1),
    .O(DLX_IDinst__n0127[19])
  );
  defparam \DLX_IDinst_Mmux__n0127_Result<18>1 .INIT = 16'hF2D0;
  X_LUT4 \DLX_IDinst_Mmux__n0127_Result<18>1  (
    .ADR0(DLX_IDinst__n03641_1),
    .ADR1(DLX_IDinst_Ker709161_1),
    .ADR2(DLX_IDinst_Cause_Reg[18]),
    .ADR3(DLX_IDinst_Imm_31_1),
    .O(DLX_IDinst__n0127[18])
  );
  defparam \DLX_IDinst_Mmux__n0127_Result<27>1 .INIT = 16'hCCAC;
  X_LUT4 \DLX_IDinst_Mmux__n0127_Result<27>1  (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(DLX_IDinst_Cause_Reg[27]),
    .ADR2(DLX_IDinst__n03641_1),
    .ADR3(DLX_IDinst_Ker709161_1),
    .O(DLX_IDinst__n0127[27])
  );
  defparam \DLX_IDinst_Mmux__n0127_Result<26>1 .INIT = 16'hDC8C;
  X_LUT4 \DLX_IDinst_Mmux__n0127_Result<26>1  (
    .ADR0(DLX_IDinst_Ker709161_1),
    .ADR1(DLX_IDinst_Cause_Reg[26]),
    .ADR2(DLX_IDinst__n03641_1),
    .ADR3(DLX_IDinst_Imm_31_1),
    .O(DLX_IDinst__n0127[26])
  );
  defparam \DLX_IDinst_Mmux__n0127_Result<29>1 .INIT = 16'hACAA;
  X_LUT4 \DLX_IDinst_Mmux__n0127_Result<29>1  (
    .ADR0(DLX_IDinst_Cause_Reg[29]),
    .ADR1(DLX_IDinst_Imm_31_1),
    .ADR2(DLX_IDinst_Ker709161_1),
    .ADR3(DLX_IDinst__n03641_1),
    .O(DLX_IDinst__n0127[29])
  );
  defparam \DLX_IDinst_Mmux__n0127_Result<28>1 .INIT = 16'hB8AA;
  X_LUT4 \DLX_IDinst_Mmux__n0127_Result<28>1  (
    .ADR0(DLX_IDinst_Cause_Reg[28]),
    .ADR1(DLX_IDinst_Ker709161_1),
    .ADR2(DLX_IDinst_Imm_31_1),
    .ADR3(DLX_IDinst__n03641_1),
    .O(DLX_IDinst__n0127[28])
  );
  defparam \DLX_EXinst__n0007<1>1 .INIT = 16'h000A;
  X_LUT4 \DLX_EXinst__n0007<1>1  (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_counter[1]),
    .ADR3(DLX_IDinst_counter[0]),
    .O(DLX_EXinst__n0007[1])
  );
  defparam \DLX_EXinst__n0007<0>1 .INIT = 16'h000A;
  X_LUT4 \DLX_EXinst__n0007<0>1  (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_counter[0]),
    .ADR3(DLX_IDinst_counter[1]),
    .O(\DLX_EXinst_reg_out_B_EX<1>/GROM )
  );
  X_BUF \DLX_EXinst_reg_out_B_EX<1>/YUSED  (
    .I(\DLX_EXinst_reg_out_B_EX<1>/GROM ),
    .O(DLX_EXinst__n0007[0])
  );
  defparam \DLX_EXinst__n0007<3>1 .INIT = 16'h0030;
  X_LUT4 \DLX_EXinst__n0007<3>1  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_counter[1]),
    .ADR2(DLX_IDinst_reg_out_B[3]),
    .ADR3(DLX_IDinst_counter[0]),
    .O(DLX_EXinst__n0007[3])
  );
  defparam \DLX_EXinst__n0007<2>1 .INIT = 16'h1100;
  X_LUT4 \DLX_EXinst__n0007<2>1  (
    .ADR0(DLX_IDinst_counter[0]),
    .ADR1(DLX_IDinst_counter[1]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[2]),
    .O(DLX_EXinst__n0007[2])
  );
  defparam \DLX_EXinst__n0007<5>1 .INIT = 16'h1010;
  X_LUT4 \DLX_EXinst__n0007<5>1  (
    .ADR0(DLX_IDinst_counter[0]),
    .ADR1(DLX_IDinst_counter[1]),
    .ADR2(DLX_IDinst_reg_out_B[5]),
    .ADR3(VCC),
    .O(DLX_EXinst__n0007[5])
  );
  defparam \DLX_EXinst__n0007<4>1 .INIT = 16'h0404;
  X_LUT4 \DLX_EXinst__n0007<4>1  (
    .ADR0(DLX_IDinst_counter[0]),
    .ADR1(DLX_IDinst_reg_out_B[4]),
    .ADR2(DLX_IDinst_counter[1]),
    .ADR3(VCC),
    .O(DLX_EXinst__n0007[4])
  );
  defparam \DLX_EXinst__n0007<7>1 .INIT = 16'h0030;
  X_LUT4 \DLX_EXinst__n0007<7>1  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_counter[0]),
    .ADR2(DLX_IDinst_reg_out_B[7]),
    .ADR3(DLX_IDinst_counter[1]),
    .O(DLX_EXinst__n0007[7])
  );
  defparam \DLX_EXinst__n0007<6>1 .INIT = 16'h1010;
  X_LUT4 \DLX_EXinst__n0007<6>1  (
    .ADR0(DLX_IDinst_counter[0]),
    .ADR1(DLX_IDinst_counter[1]),
    .ADR2(DLX_IDinst_reg_out_B[6]),
    .ADR3(VCC),
    .O(DLX_EXinst__n0007[6])
  );
  defparam \DLX_EXinst__n0007<9>1 .INIT = 16'h8888;
  X_LUT4 \DLX_EXinst__n0007<9>1  (
    .ADR0(DLX_EXinst_N66350),
    .ADR1(DLX_IDinst_reg_out_B[9]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst__n0007[9])
  );
  defparam \DLX_EXinst__n0007<8>1 .INIT = 16'h8888;
  X_LUT4 \DLX_EXinst__n0007<8>1  (
    .ADR0(DLX_IDinst_reg_out_B[8]),
    .ADR1(DLX_EXinst_N66350),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst__n0007[8])
  );
  defparam \DLX_EXinst__n0008<1>1 .INIT = 16'hA088;
  X_LUT4 \DLX_EXinst__n0008<1>1  (
    .ADR0(DLX_EXinst__n0149),
    .ADR1(DLX_IDinst_rt_addr[1]),
    .ADR2(DLX_IDinst_rd_addr[1]),
    .ADR3(DLX_IDinst_reg_dst),
    .O(DLX_EXinst__n0008[1])
  );
  defparam \DLX_EXinst__n0008<0>1 .INIT = 16'hA088;
  X_LUT4 \DLX_EXinst__n0008<0>1  (
    .ADR0(DLX_EXinst__n0149),
    .ADR1(DLX_IDinst_rt_addr[0]),
    .ADR2(DLX_IDinst_rd_addr[0]),
    .ADR3(DLX_IDinst_reg_dst),
    .O(DLX_EXinst__n0008[0])
  );
  X_OR2 \DLX_EXinst_reg_dst_out<3>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_reg_dst_out<3>/FFY/RST )
  );
  defparam DLX_EXinst_reg_dst_out_2.INIT = 1'b0;
  X_FF DLX_EXinst_reg_dst_out_2 (
    .I(DLX_EXinst__n0008[2]),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_reg_dst_out<3>/FFY/RST ),
    .O(DLX_EXinst_reg_dst_out[2])
  );
  defparam \DLX_EXinst__n0008<3>1 .INIT = 16'hE040;
  X_LUT4 \DLX_EXinst__n0008<3>1  (
    .ADR0(DLX_IDinst_reg_dst),
    .ADR1(DLX_IDinst_rt_addr[3]),
    .ADR2(DLX_EXinst__n0149),
    .ADR3(DLX_IDinst_rd_addr[3]),
    .O(DLX_EXinst__n0008[3])
  );
  defparam \DLX_EXinst__n0008<2>1 .INIT = 16'hA088;
  X_LUT4 \DLX_EXinst__n0008<2>1  (
    .ADR0(DLX_EXinst__n0149),
    .ADR1(DLX_IDinst_rt_addr[2]),
    .ADR2(DLX_IDinst_rd_addr[2]),
    .ADR3(DLX_IDinst_reg_dst),
    .O(DLX_EXinst__n0008[2])
  );
  X_OR2 \DLX_IDinst_IR_function_field<5>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_IR_function_field<5>/FFY/RST )
  );
  defparam DLX_IDinst_IR_function_field_4.INIT = 1'b0;
  X_FF DLX_IDinst_IR_function_field_4 (
    .I(DLX_IDinst__n0101),
    .CE(DLX_IDinst__n0422),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_IR_function_field<5>/FFY/RST ),
    .O(DLX_IDinst_IR_function_field[4])
  );
  defparam \DLX_IDinst__n0114<5>1 .INIT = 16'h3232;
  X_LUT4 \DLX_IDinst__n0114<5>1  (
    .ADR0(DLX_IDinst_N70918),
    .ADR1(DLX_IDinst__n0331),
    .ADR2(DLX_IDinst__n0030[5]),
    .ADR3(VCC),
    .O(DLX_IDinst__n0114[5])
  );
  defparam DLX_IDinst__n0101_1146.INIT = 16'h8880;
  X_LUT4 DLX_IDinst__n0101_1146 (
    .ADR0(DLX_IDinst_N70679),
    .ADR1(DLX_IDinst_jtarget[4]),
    .ADR2(DLX_IDinst__n0364),
    .ADR3(N90703),
    .O(DLX_IDinst__n0101)
  );
  defparam DLX_EXinst_Ker64872125.INIT = 16'h3020;
  X_LUT4 DLX_EXinst_Ker64872125 (
    .ADR0(CHOICE3205),
    .ADR1(N110935),
    .ADR2(DLX_EXinst__n0049),
    .ADR3(CHOICE3208),
    .O(\CHOICE3210/FROM )
  );
  defparam DLX_EXinst_Ker64872136.INIT = 16'hFFA0;
  X_LUT4 DLX_EXinst_Ker64872136 (
    .ADR0(N111221),
    .ADR1(VCC),
    .ADR2(CHOICE3198),
    .ADR3(CHOICE3210),
    .O(\CHOICE3210/GROM )
  );
  X_BUF \CHOICE3210/XUSED  (
    .I(\CHOICE3210/FROM ),
    .O(CHOICE3210)
  );
  X_BUF \CHOICE3210/YUSED  (
    .I(\CHOICE3210/GROM ),
    .O(N108909)
  );
  defparam \DLX_IDinst__n0117<28>29 .INIT = 16'hEAC0;
  X_LUT4 \DLX_IDinst__n0117<28>29  (
    .ADR0(N101161),
    .ADR1(DLX_IDinst_N69914),
    .ADR2(DLX_IDinst_regA_eff[28]),
    .ADR3(CHOICE2458),
    .O(\DLX_IDinst_reg_out_A<28>/FROM )
  );
  defparam \DLX_IDinst__n0117<28>39 .INIT = 16'hFFA0;
  X_LUT4 \DLX_IDinst__n0117<28>39  (
    .ADR0(DLX_IFinst_NPC[28]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst__n0310),
    .ADR3(CHOICE2461),
    .O(N104508)
  );
  X_BUF \DLX_IDinst_reg_out_A<28>/XUSED  (
    .I(\DLX_IDinst_reg_out_A<28>/FROM ),
    .O(CHOICE2461)
  );
  defparam \DLX_IDinst__n0117<5>29 .INIT = 16'hEAC0;
  X_LUT4 \DLX_IDinst__n0117<5>29  (
    .ADR0(DLX_IDinst_N69914),
    .ADR1(CHOICE2194),
    .ADR2(N101161),
    .ADR3(DLX_IDinst_regA_eff[5]),
    .O(\DLX_IDinst_reg_out_A<5>/FROM )
  );
  defparam \DLX_IDinst__n0117<5>39 .INIT = 16'hFF88;
  X_LUT4 \DLX_IDinst__n0117<5>39  (
    .ADR0(DLX_IFinst_NPC[5]),
    .ADR1(DLX_IDinst__n0310),
    .ADR2(VCC),
    .ADR3(CHOICE2197),
    .O(N103012)
  );
  X_BUF \DLX_IDinst_reg_out_A<5>/XUSED  (
    .I(\DLX_IDinst_reg_out_A<5>/FROM ),
    .O(CHOICE2197)
  );
  defparam \DLX_IDinst__n0117<22>15 .INIT = 16'h3808;
  X_LUT4 \DLX_IDinst__n0117<22>15  (
    .ADR0(DLX_IDinst_Cause_Reg[22]),
    .ADR1(DLX_IDinst_regA_index[0]),
    .ADR2(DLX_IDinst_regA_index[1]),
    .ADR3(DLX_IDinst_EPC[22]),
    .O(\CHOICE2386/FROM )
  );
  defparam \DLX_IDinst__n0117<29>15 .INIT = 16'h6420;
  X_LUT4 \DLX_IDinst__n0117<29>15  (
    .ADR0(DLX_IDinst_regA_index[1]),
    .ADR1(DLX_IDinst_regA_index[0]),
    .ADR2(DLX_IDinst_EPC[29]),
    .ADR3(DLX_IDinst_Cause_Reg[29]),
    .O(\CHOICE2386/GROM )
  );
  X_BUF \CHOICE2386/XUSED  (
    .I(\CHOICE2386/FROM ),
    .O(CHOICE2386)
  );
  X_BUF \CHOICE2386/YUSED  (
    .I(\CHOICE2386/GROM ),
    .O(CHOICE2482)
  );
  defparam \DLX_IDinst__n0117<16>15 .INIT = 16'h2C20;
  X_LUT4 \DLX_IDinst__n0117<16>15  (
    .ADR0(DLX_IDinst_Cause_Reg[16]),
    .ADR1(DLX_IDinst_regA_index[1]),
    .ADR2(DLX_IDinst_regA_index[0]),
    .ADR3(DLX_IDinst_EPC[16]),
    .O(\CHOICE2338/FROM )
  );
  defparam \DLX_IDinst__n0117<6>15 .INIT = 16'h5088;
  X_LUT4 \DLX_IDinst__n0117<6>15  (
    .ADR0(DLX_IDinst_regA_index[1]),
    .ADR1(DLX_IDinst_EPC[6]),
    .ADR2(DLX_IDinst_Cause_Reg[6]),
    .ADR3(DLX_IDinst_regA_index[0]),
    .O(\CHOICE2338/GROM )
  );
  X_BUF \CHOICE2338/XUSED  (
    .I(\CHOICE2338/FROM ),
    .O(CHOICE2338)
  );
  X_BUF \CHOICE2338/YUSED  (
    .I(\CHOICE2338/GROM ),
    .O(CHOICE2218)
  );
  defparam DLX_MEMlc_ridp31.INIT = 16'h00FF;
  X_LUT4 DLX_MEMlc_ridp31 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_MEMlc_pd_wint1),
    .O(\DLX_MEMlc_ridp3/FROM )
  );
  defparam DLX_MEMlc_md_mda2_a1.INIT = 16'h00AA;
  X_LUT4 DLX_MEMlc_md_mda2_a1 (
    .ADR0(DLX_MEMlc_md_wint1),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_MEMlc_pd_wint1),
    .O(\DLX_MEMlc_ridp3/GROM )
  );
  X_BUF \DLX_MEMlc_ridp3/XUSED  (
    .I(\DLX_MEMlc_ridp3/FROM ),
    .O(DLX_MEMlc_ridp3)
  );
  X_BUF \DLX_MEMlc_ridp3/YUSED  (
    .I(\DLX_MEMlc_ridp3/GROM ),
    .O(DLX_MEMlc_md_wint2)
  );
  defparam \DLX_EXinst_Mshift__n0025_Sh<46>_SW0 .INIT = 16'h03CF;
  X_LUT4 \DLX_EXinst_Mshift__n0025_Sh<46>_SW0  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_B_2_1),
    .ADR2(\DLX_EXinst_Mshift__n0025_Sh[14] ),
    .ADR3(\DLX_EXinst_Mshift__n0025_Sh[10] ),
    .O(\N93747/FROM )
  );
  defparam \DLX_EXinst__n0006<14>176 .INIT = 16'h880A;
  X_LUT4 \DLX_EXinst__n0006<14>176  (
    .ADR0(DLX_EXinst_N66535),
    .ADR1(DLX_EXinst_N62911),
    .ADR2(N93747),
    .ADR3(DLX_IDinst_reg_out_B[3]),
    .O(\N93747/GROM )
  );
  X_BUF \N93747/XUSED  (
    .I(\N93747/FROM ),
    .O(N93747)
  );
  X_BUF \N93747/YUSED  (
    .I(\N93747/GROM ),
    .O(CHOICE4276)
  );
  defparam \DLX_EXinst__n0006<22>41_SW0 .INIT = 16'hFF3F;
  X_LUT4 \DLX_EXinst__n0006<22>41_SW0  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N62826),
    .ADR2(DLX_IDinst_IR_function_field[4]),
    .ADR3(DLX_IDinst_IR_function_field[3]),
    .O(\N127155/FROM )
  );
  defparam \DLX_EXinst__n0006<31>395_SW0 .INIT = 16'hF3E2;
  X_LUT4 \DLX_EXinst__n0006<31>395_SW0  (
    .ADR0(CHOICE5806),
    .ADR1(DLX_IDinst_IR_function_field[3]),
    .ADR2(\DLX_EXinst_Mshift__n0027_Sh[23] ),
    .ADR3(CHOICE5801),
    .O(\N127155/GROM )
  );
  X_BUF \N127155/XUSED  (
    .I(\N127155/FROM ),
    .O(N127155)
  );
  X_BUF \N127155/YUSED  (
    .I(\N127155/GROM ),
    .O(N126154)
  );
  defparam \DLX_EXinst__n0006<23>100_SW0 .INIT = 16'hB3A0;
  X_LUT4 \DLX_EXinst__n0006<23>100_SW0  (
    .ADR0(\DLX_IDinst_Imm[7] ),
    .ADR1(DLX_IDinst_IR_function_field[4]),
    .ADR2(DLX_EXinst__n0077),
    .ADR3(N107780),
    .O(\N126593/FROM )
  );
  defparam \DLX_EXinst__n0006<21>100_SW0 .INIT = 16'hA0EC;
  X_LUT4 \DLX_EXinst__n0006<21>100_SW0  (
    .ADR0(\DLX_IDinst_Imm[5] ),
    .ADR1(N108266),
    .ADR2(DLX_EXinst__n0077),
    .ADR3(DLX_IDinst_IR_function_field[4]),
    .O(\N126593/GROM )
  );
  X_BUF \N126593/XUSED  (
    .I(\N126593/FROM ),
    .O(N126593)
  );
  X_BUF \N126593/YUSED  (
    .I(\N126593/GROM ),
    .O(N126451)
  );
  defparam \DLX_IDinst__n0117<29>29 .INIT = 16'hEAC0;
  X_LUT4 \DLX_IDinst__n0117<29>29  (
    .ADR0(DLX_IDinst_N69914),
    .ADR1(CHOICE2482),
    .ADR2(N101161),
    .ADR3(DLX_IDinst_regA_eff[29]),
    .O(\DLX_IDinst_reg_out_A<29>/FROM )
  );
  defparam \DLX_IDinst__n0117<29>39 .INIT = 16'hFFA0;
  X_LUT4 \DLX_IDinst__n0117<29>39  (
    .ADR0(DLX_IFinst_NPC[29]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst__n0310),
    .ADR3(CHOICE2485),
    .O(N104644)
  );
  X_BUF \DLX_IDinst_reg_out_A<29>/XUSED  (
    .I(\DLX_IDinst_reg_out_A<29>/FROM ),
    .O(CHOICE2485)
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<5>1 .INIT = 16'hBB88;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<5>1  (
    .ADR0(DLX_EXinst_N62946),
    .ADR1(DLX_IDinst_reg_out_B[0]),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N63284),
    .O(\DLX_EXinst_Mshift__n0023_Sh<5>/FROM )
  );
  defparam \DLX_EXinst__n0006<5>162 .INIT = 16'h3120;
  X_LUT4 \DLX_EXinst__n0006<5>162  (
    .ADR0(DLX_IDinst_reg_out_B[2]),
    .ADR1(DLX_IDinst_reg_out_B[3]),
    .ADR2(\DLX_EXinst_Mshift__n0023_Sh[9] ),
    .ADR3(\DLX_EXinst_Mshift__n0023_Sh[5] ),
    .O(\DLX_EXinst_Mshift__n0023_Sh<5>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0023_Sh<5>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0023_Sh<5>/FROM ),
    .O(\DLX_EXinst_Mshift__n0023_Sh[5] )
  );
  X_BUF \DLX_EXinst_Mshift__n0023_Sh<5>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0023_Sh<5>/GROM ),
    .O(CHOICE4459)
  );
  X_OR2 \DLX_IDinst_reg_out_A<6>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_A<6>/FFY/RST )
  );
  defparam DLX_IDinst_reg_out_A_6.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_A_6 (
    .I(N103148),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_A<6>/FFY/RST ),
    .O(DLX_IDinst_reg_out_A[6])
  );
  defparam \DLX_IDinst__n0117<6>29 .INIT = 16'hEAC0;
  X_LUT4 \DLX_IDinst__n0117<6>29  (
    .ADR0(DLX_IDinst_N69914),
    .ADR1(N101161),
    .ADR2(CHOICE2218),
    .ADR3(DLX_IDinst_regA_eff[6]),
    .O(\DLX_IDinst_reg_out_A<6>/FROM )
  );
  defparam \DLX_IDinst__n0117<6>39 .INIT = 16'hFFC0;
  X_LUT4 \DLX_IDinst__n0117<6>39  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst__n0310),
    .ADR2(DLX_IFinst_NPC[6]),
    .ADR3(CHOICE2221),
    .O(N103148)
  );
  X_BUF \DLX_IDinst_reg_out_A<6>/XUSED  (
    .I(\DLX_IDinst_reg_out_A<6>/FROM ),
    .O(CHOICE2221)
  );
  defparam \DLX_EXinst__n0006<7>16_SW0 .INIT = 16'h0505;
  X_LUT4 \DLX_EXinst__n0006<7>16_SW0  (
    .ADR0(DLX_IDinst_IR_opcode_field[0]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[7]),
    .ADR3(VCC),
    .O(\N127392/FROM )
  );
  defparam \DLX_EXinst__n0006<28>88_SW0 .INIT = 16'h1111;
  X_LUT4 \DLX_EXinst__n0006<28>88_SW0  (
    .ADR0(DLX_IDinst_IR_opcode_field[0]),
    .ADR1(DLX_IDinst_reg_out_A[28]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\N127392/GROM )
  );
  X_BUF \N127392/XUSED  (
    .I(\N127392/FROM ),
    .O(N127392)
  );
  X_BUF \N127392/YUSED  (
    .I(\N127392/GROM ),
    .O(N127298)
  );
  defparam \DLX_IDinst__n0117<5>15 .INIT = 16'h6420;
  X_LUT4 \DLX_IDinst__n0117<5>15  (
    .ADR0(DLX_IDinst_regA_index[0]),
    .ADR1(DLX_IDinst_regA_index[1]),
    .ADR2(DLX_IDinst_Cause_Reg[5]),
    .ADR3(DLX_IDinst_EPC[5]),
    .O(\CHOICE2194/FROM )
  );
  defparam \DLX_IDinst__n0117<7>15 .INIT = 16'h2C20;
  X_LUT4 \DLX_IDinst__n0117<7>15  (
    .ADR0(DLX_IDinst_EPC[7]),
    .ADR1(DLX_IDinst_regA_index[0]),
    .ADR2(DLX_IDinst_regA_index[1]),
    .ADR3(DLX_IDinst_Cause_Reg[7]),
    .O(\CHOICE2194/GROM )
  );
  X_BUF \CHOICE2194/XUSED  (
    .I(\CHOICE2194/FROM ),
    .O(CHOICE2194)
  );
  X_BUF \CHOICE2194/YUSED  (
    .I(\CHOICE2194/GROM ),
    .O(CHOICE2206)
  );
  defparam DLX_MEMlc_md_mda13_a1.INIT = 16'h0A0A;
  X_LUT4 DLX_MEMlc_md_mda13_a1 (
    .ADR0(DLX_MEMlc_md_wint12),
    .ADR1(VCC),
    .ADR2(DLX_MEMlc_pd_wint1),
    .ADR3(VCC),
    .O(\DLX_MEMlc_md_wint13/FROM )
  );
  defparam DLX_MEMlc_md_mda3_a1.INIT = 16'h00F0;
  X_LUT4 DLX_MEMlc_md_mda3_a1 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_MEMlc_md_wint2),
    .ADR3(DLX_MEMlc_pd_wint1),
    .O(\DLX_MEMlc_md_wint13/GROM )
  );
  X_BUF \DLX_MEMlc_md_wint13/XUSED  (
    .I(\DLX_MEMlc_md_wint13/FROM ),
    .O(DLX_MEMlc_md_wint13)
  );
  X_BUF \DLX_MEMlc_md_wint13/YUSED  (
    .I(\DLX_MEMlc_md_wint13/GROM ),
    .O(DLX_MEMlc_md_wint3)
  );
  defparam \DLX_IDinst__n0117<7>29 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst__n0117<7>29  (
    .ADR0(DLX_IDinst_N69914),
    .ADR1(DLX_IDinst_regA_eff[7]),
    .ADR2(N101161),
    .ADR3(CHOICE2206),
    .O(\DLX_IDinst_reg_out_A<7>/FROM )
  );
  defparam \DLX_IDinst__n0117<7>39 .INIT = 16'hFFC0;
  X_LUT4 \DLX_IDinst__n0117<7>39  (
    .ADR0(VCC),
    .ADR1(DLX_IFinst_NPC[7]),
    .ADR2(DLX_IDinst__n0310),
    .ADR3(CHOICE2209),
    .O(N103080)
  );
  X_BUF \DLX_IDinst_reg_out_A<7>/XUSED  (
    .I(\DLX_IDinst_reg_out_A<7>/FROM ),
    .O(CHOICE2209)
  );
  defparam DLX_MEMlc_slave_ctrlMEM__n0001_SW111.INIT = 16'hBA30;
  X_LUT4 DLX_MEMlc_slave_ctrlMEM__n0001_SW111 (
    .ADR0(DLX_reqout_MEM),
    .ADR1(reset_IBUF_1),
    .ADR2(DLX_MEMlc_slave_ctrlMEM_l),
    .ADR3(DLX_ackin_ID),
    .O(\CHOICE39/FROM )
  );
  defparam DLX_MEMlc_slave_ctrlMEM__n0001_SW112.INIT = 16'hCC00;
  X_LUT4 DLX_MEMlc_slave_ctrlMEM__n0001_SW112 (
    .ADR0(VCC),
    .ADR1(DLX_MEMlc_master_ctrlMEM_nro),
    .ADR2(VCC),
    .ADR3(CHOICE39),
    .O(\CHOICE39/GROM )
  );
  X_BUF \CHOICE39/XUSED  (
    .I(\CHOICE39/FROM ),
    .O(CHOICE39)
  );
  X_BUF \CHOICE39/YUSED  (
    .I(\CHOICE39/GROM ),
    .O(DLX_MEMlc_slave_ctrlMEM_l)
  );
  defparam \DLX_IDinst__n0117<25>15 .INIT = 16'h44A0;
  X_LUT4 \DLX_IDinst__n0117<25>15  (
    .ADR0(DLX_IDinst_regA_index[1]),
    .ADR1(DLX_IDinst_Cause_Reg[25]),
    .ADR2(DLX_IDinst_EPC[25]),
    .ADR3(DLX_IDinst_regA_index[0]),
    .O(\CHOICE2422/FROM )
  );
  defparam \DLX_IDinst__n0117<8>15 .INIT = 16'h6240;
  X_LUT4 \DLX_IDinst__n0117<8>15  (
    .ADR0(DLX_IDinst_regA_index[1]),
    .ADR1(DLX_IDinst_regA_index[0]),
    .ADR2(DLX_IDinst_Cause_Reg[8]),
    .ADR3(DLX_IDinst_EPC[8]),
    .O(\CHOICE2422/GROM )
  );
  X_BUF \CHOICE2422/XUSED  (
    .I(\CHOICE2422/FROM ),
    .O(CHOICE2422)
  );
  X_BUF \CHOICE2422/YUSED  (
    .I(\CHOICE2422/GROM ),
    .O(CHOICE2230)
  );
  defparam DLX_MEMlc_md_mda12_a1.INIT = 16'h0C0C;
  X_LUT4 DLX_MEMlc_md_mda12_a1 (
    .ADR0(VCC),
    .ADR1(DLX_MEMlc_md_wint11),
    .ADR2(DLX_MEMlc_pd_wint1),
    .ADR3(VCC),
    .O(\DLX_MEMlc_md_wint12/FROM )
  );
  defparam DLX_MEMlc_md_mda4_a1.INIT = 16'h00CC;
  X_LUT4 DLX_MEMlc_md_mda4_a1 (
    .ADR0(VCC),
    .ADR1(DLX_MEMlc_md_wint3),
    .ADR2(VCC),
    .ADR3(DLX_MEMlc_pd_wint1),
    .O(\DLX_MEMlc_md_wint12/GROM )
  );
  X_BUF \DLX_MEMlc_md_wint12/XUSED  (
    .I(\DLX_MEMlc_md_wint12/FROM ),
    .O(DLX_MEMlc_md_wint12)
  );
  X_BUF \DLX_MEMlc_md_wint12/YUSED  (
    .I(\DLX_MEMlc_md_wint12/GROM ),
    .O(DLX_MEMlc_md_wint4)
  );
  defparam DLX_EXinst_Ker661751.INIT = 16'hF000;
  X_LUT4 DLX_EXinst_Ker661751 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[4]),
    .ADR3(N111221),
    .O(\DLX_EXinst_N66177/FROM )
  );
  defparam DLX_EXinst_Ker64867108.INIT = 16'hEEAA;
  X_LUT4 DLX_EXinst_Ker64867108 (
    .ADR0(CHOICE3132),
    .ADR1(CHOICE3124),
    .ADR2(VCC),
    .ADR3(N111221),
    .O(\DLX_EXinst_N66177/GROM )
  );
  X_BUF \DLX_EXinst_N66177/XUSED  (
    .I(\DLX_EXinst_N66177/FROM ),
    .O(DLX_EXinst_N66177)
  );
  X_BUF \DLX_EXinst_N66177/YUSED  (
    .I(\DLX_EXinst_N66177/GROM ),
    .O(N108433)
  );
  defparam \DLX_EXinst__n0006<30>335_SW0 .INIT = 16'hFFEA;
  X_LUT4 \DLX_EXinst__n0006<30>335_SW0  (
    .ADR0(CHOICE5316),
    .ADR1(N95120),
    .ADR2(DLX_EXinst_N66078),
    .ADR3(CHOICE5307),
    .O(\N126519/FROM )
  );
  defparam \DLX_EXinst__n0006<28>331_SW0 .INIT = 16'hFFEA;
  X_LUT4 \DLX_EXinst__n0006<28>331_SW0  (
    .ADR0(CHOICE5239),
    .ADR1(DLX_EXinst_N66078),
    .ADR2(N95810),
    .ADR3(CHOICE5230),
    .O(\N126519/GROM )
  );
  X_BUF \N126519/XUSED  (
    .I(\N126519/FROM ),
    .O(N126519)
  );
  X_BUF \N126519/YUSED  (
    .I(\N126519/GROM ),
    .O(N126584)
  );
  defparam \DLX_EXinst__n0006<19>387_SW0 .INIT = 16'h3332;
  X_LUT4 \DLX_EXinst__n0006<19>387_SW0  (
    .ADR0(CHOICE4973),
    .ADR1(DLX_EXinst__n0030),
    .ADR2(CHOICE4944),
    .ADR3(CHOICE4941),
    .O(\DLX_EXinst_ALU_result<19>/FROM )
  );
  defparam \DLX_EXinst__n0006<19>387 .INIT = 16'hAAA8;
  X_LUT4 \DLX_EXinst__n0006<19>387  (
    .ADR0(DLX_EXinst__n0149),
    .ADR1(N100490),
    .ADR2(CHOICE5011),
    .ADR3(N126461),
    .O(N119626)
  );
  X_BUF \DLX_EXinst_ALU_result<19>/XUSED  (
    .I(\DLX_EXinst_ALU_result<19>/FROM ),
    .O(N126461)
  );
  defparam DLX_reqin_IF1.INIT = 16'h0C0C;
  X_LUT4 DLX_reqin_IF1 (
    .ADR0(VCC),
    .ADR1(DLX_reqout_ID),
    .ADR2(STOP_fetch_IBUF),
    .ADR3(VCC),
    .O(\DLX_reqin_IF/GROM )
  );
  X_BUF \DLX_reqin_IF/YUSED  (
    .I(\DLX_reqin_IF/GROM ),
    .O(DLX_reqin_IF)
  );
  defparam \DLX_IDinst__n0117<8>29 .INIT = 16'hECA0;
  X_LUT4 \DLX_IDinst__n0117<8>29  (
    .ADR0(CHOICE2230),
    .ADR1(DLX_IDinst_regA_eff[8]),
    .ADR2(N101161),
    .ADR3(DLX_IDinst_N69914),
    .O(\DLX_IDinst_reg_out_A<8>/FROM )
  );
  defparam \DLX_IDinst__n0117<8>39 .INIT = 16'hFFA0;
  X_LUT4 \DLX_IDinst__n0117<8>39  (
    .ADR0(DLX_IFinst_NPC[8]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst__n0310),
    .ADR3(CHOICE2233),
    .O(N103216)
  );
  X_BUF \DLX_IDinst_reg_out_A<8>/XUSED  (
    .I(\DLX_IDinst_reg_out_A<8>/FROM ),
    .O(CHOICE2233)
  );
  defparam \DLX_EXinst__n0006<2>129_SW0 .INIT = 16'hFAAA;
  X_LUT4 \DLX_EXinst__n0006<2>129_SW0  (
    .ADR0(CHOICE5509),
    .ADR1(VCC),
    .ADR2(N97521),
    .ADR3(DLX_IDinst_IR_function_field[2]),
    .O(\N126297/FROM )
  );
  defparam \DLX_EXinst__n0006<3>129_SW0 .INIT = 16'hFCAC;
  X_LUT4 \DLX_EXinst__n0006<3>129_SW0  (
    .ADR0(CHOICE1090),
    .ADR1(N127440),
    .ADR2(DLX_IDinst_IR_function_field[2]),
    .ADR3(CHOICE1096),
    .O(\N126297/GROM )
  );
  X_BUF \N126297/XUSED  (
    .I(\N126297/FROM ),
    .O(N126297)
  );
  X_BUF \N126297/YUSED  (
    .I(\N126297/GROM ),
    .O(N126393)
  );
  defparam DLX_IDinst_Ker706511.INIT = 16'h0070;
  X_LUT4 DLX_IDinst_Ker706511 (
    .ADR0(DLX_IDinst_slot_num_FFd1),
    .ADR1(DLX_IDinst_delay_slot),
    .ADR2(FREEZE_IBUF),
    .ADR3(DLX_IDinst_intr_slot),
    .O(\DLX_IDinst_N70653/FROM )
  );
  defparam DLX_IDinst__n0420_SW0.INIT = 16'hFFF0;
  X_LUT4 DLX_IDinst__n0420_SW0 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_delay_slot),
    .ADR3(DLX_IDinst_intr_slot),
    .O(\DLX_IDinst_N70653/GROM )
  );
  X_BUF \DLX_IDinst_N70653/XUSED  (
    .I(\DLX_IDinst_N70653/FROM ),
    .O(DLX_IDinst_N70653)
  );
  X_BUF \DLX_IDinst_N70653/YUSED  (
    .I(\DLX_IDinst_N70653/GROM ),
    .O(N90148)
  );
  defparam \DLX_IDinst__n0117<12>15 .INIT = 16'h6420;
  X_LUT4 \DLX_IDinst__n0117<12>15  (
    .ADR0(DLX_IDinst_regA_index[0]),
    .ADR1(DLX_IDinst_regA_index[1]),
    .ADR2(DLX_IDinst_Cause_Reg[12]),
    .ADR3(DLX_IDinst_EPC[12]),
    .O(\CHOICE2266/FROM )
  );
  defparam \DLX_IDinst__n0117<9>15 .INIT = 16'h6240;
  X_LUT4 \DLX_IDinst__n0117<9>15  (
    .ADR0(DLX_IDinst_regA_index[0]),
    .ADR1(DLX_IDinst_regA_index[1]),
    .ADR2(DLX_IDinst_EPC[9]),
    .ADR3(DLX_IDinst_Cause_Reg[9]),
    .O(\CHOICE2266/GROM )
  );
  X_BUF \CHOICE2266/XUSED  (
    .I(\CHOICE2266/FROM ),
    .O(CHOICE2266)
  );
  X_BUF \CHOICE2266/YUSED  (
    .I(\CHOICE2266/GROM ),
    .O(CHOICE2242)
  );
  defparam \DLX_EXinst__n0006<22>85_SW0 .INIT = 16'h1111;
  X_LUT4 \DLX_EXinst__n0006<22>85_SW0  (
    .ADR0(DLX_IDinst_IR_opcode_field[0]),
    .ADR1(DLX_IDinst_reg_out_A[22]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\N127388/FROM )
  );
  defparam \DLX_EXinst__n0006<5>16_SW0 .INIT = 16'h0505;
  X_LUT4 \DLX_EXinst__n0006<5>16_SW0  (
    .ADR0(DLX_IDinst_IR_opcode_field[0]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[5]),
    .ADR3(VCC),
    .O(\N127388/GROM )
  );
  X_BUF \N127388/XUSED  (
    .I(\N127388/FROM ),
    .O(N127388)
  );
  X_BUF \N127388/YUSED  (
    .I(\N127388/GROM ),
    .O(N127318)
  );
  defparam DLX_MEMlc_md_mda7_a1.INIT = 16'h0F00;
  X_LUT4 DLX_MEMlc_md_mda7_a1 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_MEMlc_pd_wint1),
    .ADR3(DLX_MEMlc_md_wint6),
    .O(\DLX_MEMlc_md_wint7/FROM )
  );
  defparam DLX_MEMlc_md_mda5_a1.INIT = 16'h0F00;
  X_LUT4 DLX_MEMlc_md_mda5_a1 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_MEMlc_pd_wint1),
    .ADR3(DLX_MEMlc_md_wint4),
    .O(\DLX_MEMlc_md_wint7/GROM )
  );
  X_BUF \DLX_MEMlc_md_wint7/XUSED  (
    .I(\DLX_MEMlc_md_wint7/FROM ),
    .O(DLX_MEMlc_md_wint7)
  );
  X_BUF \DLX_MEMlc_md_wint7/YUSED  (
    .I(\DLX_MEMlc_md_wint7/GROM ),
    .O(DLX_MEMlc_md_wint5)
  );
  defparam \DLX_IDinst__n0117<9>29 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst__n0117<9>29  (
    .ADR0(N101161),
    .ADR1(CHOICE2242),
    .ADR2(DLX_IDinst_regA_eff[9]),
    .ADR3(DLX_IDinst_N69914),
    .O(\DLX_IDinst_reg_out_A<9>/FROM )
  );
  defparam \DLX_IDinst__n0117<9>39 .INIT = 16'hFFA0;
  X_LUT4 \DLX_IDinst__n0117<9>39  (
    .ADR0(DLX_IDinst__n0310),
    .ADR1(VCC),
    .ADR2(DLX_IFinst_NPC[9]),
    .ADR3(CHOICE2245),
    .O(N103284)
  );
  X_BUF \DLX_IDinst_reg_out_A<9>/XUSED  (
    .I(\DLX_IDinst_reg_out_A<9>/FROM ),
    .O(CHOICE2245)
  );
  defparam DLX_EXinst_Ker64060.INIT = 16'hF3C0;
  X_LUT4 DLX_EXinst_Ker64060 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_IR_function_field[3]),
    .ADR2(\DLX_EXinst_Mshift__n0027_Sh[9] ),
    .ADR3(N93127),
    .O(\DLX_EXinst_N64062/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0027_Sh<45>_SW0 .INIT = 16'hF3C0;
  X_LUT4 \DLX_EXinst_Mshift__n0027_Sh<45>_SW0  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_IR_function_field_2_1),
    .ADR2(\DLX_EXinst_Mshift__n0027_Sh[9] ),
    .ADR3(\DLX_EXinst_Mshift__n0027_Sh[13] ),
    .O(\DLX_EXinst_N64062/GROM )
  );
  X_BUF \DLX_EXinst_N64062/XUSED  (
    .I(\DLX_EXinst_N64062/FROM ),
    .O(DLX_EXinst_N64062)
  );
  X_BUF \DLX_EXinst_N64062/YUSED  (
    .I(\DLX_EXinst_N64062/GROM ),
    .O(N93279)
  );
  defparam DLX_EXinst_Ker64877107.INIT = 16'hECA0;
  X_LUT4 DLX_EXinst_Ker64877107 (
    .ADR0(N126268),
    .ADR1(CHOICE2997),
    .ADR2(N111221),
    .ADR3(DLX_EXinst_N66494),
    .O(\N107613/FROM )
  );
  defparam \DLX_EXinst__n0006<23>236 .INIT = 16'hF5F0;
  X_LUT4 \DLX_EXinst__n0006<23>236  (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(VCC),
    .ADR2(CHOICE4087),
    .ADR3(N107613),
    .O(\N107613/GROM )
  );
  X_BUF \N107613/XUSED  (
    .I(\N107613/FROM ),
    .O(N107613)
  );
  X_BUF \N107613/YUSED  (
    .I(\N107613/GROM ),
    .O(CHOICE4088)
  );
  defparam DLX_IDinst__n012052.INIT = 16'hF0FE;
  X_LUT4 DLX_IDinst__n012052 (
    .ADR0(CHOICE3494),
    .ADR1(CHOICE3493),
    .ADR2(CHOICE3499),
    .ADR3(DLX_IDinst__n0135),
    .O(\CHOICE3500/FROM )
  );
  defparam DLX_IDinst__n0120111_SW0.INIT = 16'h4000;
  X_LUT4 DLX_IDinst__n0120111_SW0 (
    .ADR0(DLX_IDinst__n0364),
    .ADR1(DLX_IDinst_N69568),
    .ADR2(DLX_IDinst_N70679),
    .ADR3(CHOICE3500),
    .O(\CHOICE3500/GROM )
  );
  X_BUF \CHOICE3500/XUSED  (
    .I(\CHOICE3500/FROM ),
    .O(CHOICE3500)
  );
  X_BUF \CHOICE3500/YUSED  (
    .I(\CHOICE3500/GROM ),
    .O(N126293)
  );
  defparam DLX_MEMlc_md_mda1_a1.INIT = 16'h0A0A;
  X_LUT4 DLX_MEMlc_md_mda1_a1 (
    .ADR0(DLX_MEMlc_ridp3),
    .ADR1(VCC),
    .ADR2(DLX_MEMlc_pd_wint1),
    .ADR3(VCC),
    .O(\DLX_MEMlc_md_wint1/FROM )
  );
  defparam DLX_MEMlc_md_mda6_a1.INIT = 16'h0F00;
  X_LUT4 DLX_MEMlc_md_mda6_a1 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_MEMlc_pd_wint1),
    .ADR3(DLX_MEMlc_md_wint5),
    .O(\DLX_MEMlc_md_wint1/GROM )
  );
  X_BUF \DLX_MEMlc_md_wint1/XUSED  (
    .I(\DLX_MEMlc_md_wint1/FROM ),
    .O(DLX_MEMlc_md_wint1)
  );
  X_BUF \DLX_MEMlc_md_wint1/YUSED  (
    .I(\DLX_MEMlc_md_wint1/GROM ),
    .O(DLX_MEMlc_md_wint6)
  );
  defparam DLX_EXinst_Ker64065_SW0.INIT = 16'hACAC;
  X_LUT4 DLX_EXinst_Ker64065_SW0 (
    .ADR0(DLX_EXinst_N62791),
    .ADR1(DLX_EXinst_N63459),
    .ADR2(DLX_IDinst_IR_function_field[0]),
    .ADR3(VCC),
    .O(\N93229/FROM )
  );
  defparam DLX_EXinst_Ker64060_SW0.INIT = 16'hE2E2;
  X_LUT4 DLX_EXinst_Ker64060_SW0 (
    .ADR0(DLX_EXinst_N62791),
    .ADR1(DLX_IDinst_IR_function_field[0]),
    .ADR2(DLX_EXinst_N63454),
    .ADR3(VCC),
    .O(\N93229/GROM )
  );
  X_BUF \N93229/XUSED  (
    .I(\N93229/FROM ),
    .O(N93229)
  );
  X_BUF \N93229/YUSED  (
    .I(\N93229/GROM ),
    .O(N93127)
  );
  defparam DLX_EXlc_slave_ctrlEX__n0001_SW110.INIT = 16'h4F44;
  X_LUT4 DLX_EXlc_slave_ctrlEX__n0001_SW110 (
    .ADR0(DLX_MEMlc_master_ctrlMEM_l),
    .ADR1(DLX_reqout_EX),
    .ADR2(reset_IBUF),
    .ADR3(DLX_EXlc_slave_ctrlEX_l),
    .O(\CHOICE45/FROM )
  );
  defparam DLX_MEMlc_master_ctrlMEM__n00021.INIT = 16'hF0FA;
  X_LUT4 DLX_MEMlc_master_ctrlMEM__n00021 (
    .ADR0(DLX_MEMlc_master_ctrlMEM_nro),
    .ADR1(VCC),
    .ADR2(DLX_MEMlc_master_ctrlMEM_l),
    .ADR3(DLX_MEMlc_slave_ctrlMEM_l),
    .O(\CHOICE45/GROM )
  );
  X_BUF \CHOICE45/XUSED  (
    .I(\CHOICE45/FROM ),
    .O(CHOICE45)
  );
  X_BUF \CHOICE45/YUSED  (
    .I(\CHOICE45/GROM ),
    .O(DLX_MEMlc_master_ctrlMEM_nro)
  );
  defparam \DLX_EXinst_Mshift__n0025_Sh<47>_SW0 .INIT = 16'h11DD;
  X_LUT4 \DLX_EXinst_Mshift__n0025_Sh<47>_SW0  (
    .ADR0(\DLX_EXinst_Mshift__n0025_Sh[15] ),
    .ADR1(DLX_IDinst_reg_out_B_2_1),
    .ADR2(VCC),
    .ADR3(\DLX_EXinst_Mshift__n0025_Sh[11] ),
    .O(\N93695/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0025_Sh<47> .INIT = 16'hC0F3;
  X_LUT4 \DLX_EXinst_Mshift__n0025_Sh<47>  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_B_3_1),
    .ADR2(DLX_EXinst_N62916),
    .ADR3(N93695),
    .O(\N93695/GROM )
  );
  X_BUF \N93695/XUSED  (
    .I(\N93695/FROM ),
    .O(N93695)
  );
  X_BUF \N93695/YUSED  (
    .I(\N93695/GROM ),
    .O(\DLX_EXinst_Mshift__n0025_Sh[47] )
  );
  defparam DLX_RF_delay_inst_wint101.INIT = 16'h5555;
  X_LUT4 DLX_RF_delay_inst_wint101 (
    .ADR0(DLX_RF_delay_inst_wint9),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_RF_delay_inst_wint10/GROM )
  );
  X_BUF \DLX_RF_delay_inst_wint10/YUSED  (
    .I(\DLX_RF_delay_inst_wint10/GROM ),
    .O(DLX_RF_delay_inst_wint10)
  );
  defparam DLX_IDinst__n010813.INIT = 16'h002A;
  X_LUT4 DLX_IDinst__n010813 (
    .ADR0(DLX_IDinst__n0135),
    .ADR1(DLX_IDinst_N70647),
    .ADR2(N98420),
    .ADR3(N98613),
    .O(\CHOICE3436/FROM )
  );
  defparam DLX_IDinst__n012048.INIT = 16'hA888;
  X_LUT4 DLX_IDinst__n012048 (
    .ADR0(DLX_IDinst__n0135),
    .ADR1(N98613),
    .ADR2(N98420),
    .ADR3(DLX_IDinst_N70647),
    .O(\CHOICE3436/GROM )
  );
  X_BUF \CHOICE3436/XUSED  (
    .I(\CHOICE3436/FROM ),
    .O(CHOICE3436)
  );
  X_BUF \CHOICE3436/YUSED  (
    .I(\CHOICE3436/GROM ),
    .O(CHOICE3499)
  );
  defparam vga_top_vga1_Ker733611.INIT = 16'h0300;
  X_LUT4 vga_top_vga1_Ker733611 (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_vcounter[5]),
    .ADR2(vga_top_vga1_vcounter[4]),
    .ADR3(vga_top_vga1_N73394),
    .O(\vga_top_vga1_N73363/FROM )
  );
  defparam vga_top_vga1__n000819.INIT = 16'h7F00;
  X_LUT4 vga_top_vga1__n000819 (
    .ADR0(vga_top_vga1_vcounter[1]),
    .ADR1(vga_top_vga1_vcounter[3]),
    .ADR2(vga_top_vga1_vcounter[2]),
    .ADR3(vga_top_vga1_N73363),
    .O(\vga_top_vga1_N73363/GROM )
  );
  X_BUF \vga_top_vga1_N73363/XUSED  (
    .I(\vga_top_vga1_N73363/FROM ),
    .O(vga_top_vga1_N73363)
  );
  X_BUF \vga_top_vga1_N73363/YUSED  (
    .I(\vga_top_vga1_N73363/GROM ),
    .O(CHOICE3221)
  );
  defparam DLX_RF_delay_inst_wint111.INIT = 16'h3333;
  X_LUT4 DLX_RF_delay_inst_wint111 (
    .ADR0(VCC),
    .ADR1(DLX_RF_delay_inst_wint10),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_RF_delay_inst_wint11/GROM )
  );
  X_BUF \DLX_RF_delay_inst_wint11/YUSED  (
    .I(\DLX_RF_delay_inst_wint11/GROM ),
    .O(DLX_RF_delay_inst_wint11)
  );
  defparam DLX_IDinst__n04211.INIT = 16'h4505;
  X_LUT4 DLX_IDinst__n04211 (
    .ADR0(DLX_IDinst__n0331),
    .ADR1(DLX_IDinst_slot_num_FFd2),
    .ADR2(DLX_IDinst_stall),
    .ADR3(DLX_IDinst_delay_slot),
    .O(\DLX_IDinst__n0421/FROM )
  );
  defparam DLX_IDinst__n0085_SW1.INIT = 16'hFF2A;
  X_LUT4 DLX_IDinst__n0085_SW1 (
    .ADR0(DLX_IDinst_stall),
    .ADR1(DLX_IDinst_delay_slot),
    .ADR2(DLX_IDinst_slot_num_FFd2),
    .ADR3(reset_IBUF),
    .O(\DLX_IDinst__n0421/GROM )
  );
  X_BUF \DLX_IDinst__n0421/XUSED  (
    .I(\DLX_IDinst__n0421/FROM ),
    .O(DLX_IDinst__n0421)
  );
  X_BUF \DLX_IDinst__n0421/YUSED  (
    .I(\DLX_IDinst__n0421/GROM ),
    .O(N127098)
  );
  defparam DLX_RF_delay_inst_wint121.INIT = 16'h3333;
  X_LUT4 DLX_RF_delay_inst_wint121 (
    .ADR0(VCC),
    .ADR1(DLX_RF_delay_inst_wint11),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_RF_delay_inst_wint12/GROM )
  );
  X_BUF \DLX_RF_delay_inst_wint12/YUSED  (
    .I(\DLX_RF_delay_inst_wint12/GROM ),
    .O(DLX_RF_delay_inst_wint12)
  );
  defparam DLX_RF_delay_inst_wint201.INIT = 16'h00FF;
  X_LUT4 DLX_RF_delay_inst_wint201 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_RF_delay_inst_wint19),
    .O(\DLX_RF_delay_inst_wint20/FROM )
  );
  defparam DLX_RF_delay_inst_wint211.INIT = 16'h00FF;
  X_LUT4 DLX_RF_delay_inst_wint211 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_RF_delay_inst_wint20),
    .O(\DLX_RF_delay_inst_wint20/GROM )
  );
  X_BUF \DLX_RF_delay_inst_wint20/XUSED  (
    .I(\DLX_RF_delay_inst_wint20/FROM ),
    .O(DLX_RF_delay_inst_wint20)
  );
  X_BUF \DLX_RF_delay_inst_wint20/YUSED  (
    .I(\DLX_RF_delay_inst_wint20/GROM ),
    .O(DLX_RF_delay_inst_wint21)
  );
  defparam vga_top_vga1_Ker733551.INIT = 16'h0010;
  X_LUT4 vga_top_vga1_Ker733551 (
    .ADR0(vga_top_vga1_hcounter[4]),
    .ADR1(vga_top_vga1_hcounter[1]),
    .ADR2(vga_top_vga1_N73379),
    .ADR3(vga_top_vga1_hcounter[7]),
    .O(\vga_top_vga1_N73357/FROM )
  );
  defparam vga_top_vga1_Ker733871.INIT = 16'hA000;
  X_LUT4 vga_top_vga1_Ker733871 (
    .ADR0(vga_top_vga1_hcounter[5]),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_hcounter[2]),
    .ADR3(vga_top_vga1_N73357),
    .O(\vga_top_vga1_N73357/GROM )
  );
  X_BUF \vga_top_vga1_N73357/XUSED  (
    .I(\vga_top_vga1_N73357/FROM ),
    .O(vga_top_vga1_N73357)
  );
  X_BUF \vga_top_vga1_N73357/YUSED  (
    .I(\vga_top_vga1_N73357/GROM ),
    .O(vga_top_vga1_N73389)
  );
  defparam DLX_RF_delay_inst_wint131.INIT = 16'h0F0F;
  X_LUT4 DLX_RF_delay_inst_wint131 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_RF_delay_inst_wint12),
    .ADR3(VCC),
    .O(\DLX_RF_delay_inst_wint13/GROM )
  );
  X_BUF \DLX_RF_delay_inst_wint13/YUSED  (
    .I(\DLX_RF_delay_inst_wint13/GROM ),
    .O(DLX_RF_delay_inst_wint13)
  );
  defparam DM_delay_inst_wint11_1147.INIT = 16'h00FF;
  X_LUT4 DM_delay_inst_wint11_1147 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_clk_EX),
    .O(\DM_delay_inst_wint1/GROM )
  );
  X_BUF \DM_delay_inst_wint1/YUSED  (
    .I(\DM_delay_inst_wint1/GROM ),
    .O(DM_delay_inst_wint1)
  );
  defparam vga_top_vga1_Ker733721.INIT = 16'h0101;
  X_LUT4 vga_top_vga1_Ker733721 (
    .ADR0(vga_top_vga1_vcounter[2]),
    .ADR1(vga_top_vga1_vcounter[4]),
    .ADR2(vga_top_vga1_vcounter[3]),
    .ADR3(VCC),
    .O(\vga_top_vga1_N73374/FROM )
  );
  defparam vga_top_vga1__n000954.INIT = 16'h1303;
  X_LUT4 vga_top_vga1__n000954 (
    .ADR0(vga_top_vga1_vcounter[1]),
    .ADR1(vga_top_vga1_vcounter[9]),
    .ADR2(vga_top_vga1_vcounter[5]),
    .ADR3(vga_top_vga1_N73374),
    .O(\vga_top_vga1_N73374/GROM )
  );
  X_BUF \vga_top_vga1_N73374/XUSED  (
    .I(\vga_top_vga1_N73374/FROM ),
    .O(vga_top_vga1_N73374)
  );
  X_BUF \vga_top_vga1_N73374/YUSED  (
    .I(\vga_top_vga1_N73374/GROM ),
    .O(CHOICE3425)
  );
  defparam DLX_IDinst__n010830.INIT = 16'h1B0A;
  X_LUT4 DLX_IDinst__n010830 (
    .ADR0(DLX_IDinst__n0136),
    .ADR1(DLX_IDinst__n0347),
    .ADR2(DLX_IDinst__n0344),
    .ADR3(DLX_IDinst__n0345),
    .O(\CHOICE3444/FROM )
  );
  defparam DLX_IDinst__n010834.INIT = 16'hF300;
  X_LUT4 DLX_IDinst__n010834 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst__n0073),
    .ADR2(DLX_IDinst__n0002),
    .ADR3(CHOICE3444),
    .O(\CHOICE3444/GROM )
  );
  X_BUF \CHOICE3444/XUSED  (
    .I(\CHOICE3444/FROM ),
    .O(CHOICE3444)
  );
  X_BUF \CHOICE3444/YUSED  (
    .I(\CHOICE3444/GROM ),
    .O(CHOICE3445)
  );
  defparam DLX_RF_delay_inst_wint141.INIT = 16'h3333;
  X_LUT4 DLX_RF_delay_inst_wint141 (
    .ADR0(VCC),
    .ADR1(DLX_RF_delay_inst_wint13),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_RF_delay_inst_wint14/FROM )
  );
  defparam DLX_RF_delay_inst_wint151.INIT = 16'h00FF;
  X_LUT4 DLX_RF_delay_inst_wint151 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_RF_delay_inst_wint14),
    .O(\DLX_RF_delay_inst_wint14/GROM )
  );
  X_BUF \DLX_RF_delay_inst_wint14/XUSED  (
    .I(\DLX_RF_delay_inst_wint14/FROM ),
    .O(DLX_RF_delay_inst_wint14)
  );
  X_BUF \DLX_RF_delay_inst_wint14/YUSED  (
    .I(\DLX_RF_delay_inst_wint14/GROM ),
    .O(DLX_RF_delay_inst_wint15)
  );
  defparam DLX_RF_delay_inst_wint221.INIT = 16'h3333;
  X_LUT4 DLX_RF_delay_inst_wint221 (
    .ADR0(VCC),
    .ADR1(DLX_RF_delay_inst_wint21),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_RF_delay_inst_wint22/GROM )
  );
  X_BUF \DLX_RF_delay_inst_wint22/YUSED  (
    .I(\DLX_RF_delay_inst_wint22/GROM ),
    .O(DLX_RF_delay_inst_wint22)
  );
  defparam DLX_RF_delay_inst_wint301.INIT = 16'h3333;
  X_LUT4 DLX_RF_delay_inst_wint301 (
    .ADR0(VCC),
    .ADR1(DLX_RF_delay_inst_wint29),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_RF_delay_inst_wint30/GROM )
  );
  X_BUF \DLX_RF_delay_inst_wint30/YUSED  (
    .I(\DLX_RF_delay_inst_wint30/GROM ),
    .O(DLX_RF_delay_inst_wint30)
  );
  defparam DM_delay_inst_wint21_1148.INIT = 16'h0F0F;
  X_LUT4 DM_delay_inst_wint21_1148 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DM_delay_inst_wint1),
    .ADR3(VCC),
    .O(\DM_delay_inst_wint2/GROM )
  );
  X_BUF \DM_delay_inst_wint2/YUSED  (
    .I(\DM_delay_inst_wint2/GROM ),
    .O(DM_delay_inst_wint2)
  );
  defparam DLX_RF_delay_inst_wint231.INIT = 16'h00FF;
  X_LUT4 DLX_RF_delay_inst_wint231 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_RF_delay_inst_wint22),
    .O(\DLX_RF_delay_inst_wint23/GROM )
  );
  X_BUF \DLX_RF_delay_inst_wint23/YUSED  (
    .I(\DLX_RF_delay_inst_wint23/GROM ),
    .O(DLX_RF_delay_inst_wint23)
  );
  defparam DM_delay_inst_wint31_1149.INIT = 16'h0F0F;
  X_LUT4 DM_delay_inst_wint31_1149 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DM_delay_inst_wint2),
    .ADR3(VCC),
    .O(\DM_delay_inst_wint3/GROM )
  );
  X_BUF \DM_delay_inst_wint3/YUSED  (
    .I(\DM_delay_inst_wint3/GROM ),
    .O(DM_delay_inst_wint3)
  );
  defparam DLX_IDinst__n010922.INIT = 16'hEE66;
  X_LUT4 DLX_IDinst__n010922 (
    .ADR0(DLX_IDinst_IR_latched[30]),
    .ADR1(DLX_IDinst_IR_latched[27]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_IR_latched[28]),
    .O(\CHOICE3518/FROM )
  );
  defparam DLX_IDinst__n010927.INIT = 16'hFF5D;
  X_LUT4 DLX_IDinst__n010927 (
    .ADR0(DLX_IDinst_N70909),
    .ADR1(DLX_IDinst_IR_latched[26]),
    .ADR2(DLX_IDinst_IR_latched[28]),
    .ADR3(CHOICE3518),
    .O(\CHOICE3518/GROM )
  );
  X_BUF \CHOICE3518/XUSED  (
    .I(\CHOICE3518/FROM ),
    .O(CHOICE3518)
  );
  X_BUF \CHOICE3518/YUSED  (
    .I(\CHOICE3518/GROM ),
    .O(CHOICE3519)
  );
  defparam \DLX_EXinst__n0006<7>204 .INIT = 16'hEAC0;
  X_LUT4 \DLX_EXinst__n0006<7>204  (
    .ADR0(N107613),
    .ADR1(N101725),
    .ADR2(DLX_EXinst_ALU_result[7]),
    .ADR3(DLX_IDinst_reg_out_B[4]),
    .O(\CHOICE3847/FROM )
  );
  defparam \DLX_EXinst__n0006<7>228_SW0 .INIT = 16'hFF0E;
  X_LUT4 \DLX_EXinst__n0006<7>228_SW0  (
    .ADR0(CHOICE3836),
    .ADR1(CHOICE3833),
    .ADR2(DLX_IDinst_reg_out_B[4]),
    .ADR3(CHOICE3847),
    .O(\CHOICE3847/GROM )
  );
  X_BUF \CHOICE3847/XUSED  (
    .I(\CHOICE3847/FROM ),
    .O(CHOICE3847)
  );
  X_BUF \CHOICE3847/YUSED  (
    .I(\CHOICE3847/GROM ),
    .O(N126465)
  );
  defparam DLX_EXinst__n001810.INIT = 16'hFFFB;
  X_LUT4 DLX_EXinst__n001810 (
    .ADR0(DLX_IDinst_IR_opcode_field[0]),
    .ADR1(DLX_IDinst_IR_function_field[5]),
    .ADR2(DLX_IDinst_IR_function_field[4]),
    .ADR3(DLX_IDinst_IR_function_field[1]),
    .O(\CHOICE3166/FROM )
  );
  defparam DLX_EXinst__n001820.INIT = 16'h0F0E;
  X_LUT4 DLX_EXinst__n001820 (
    .ADR0(DLX_IDinst_IR_function_field[2]),
    .ADR1(DLX_IDinst_IR_function_field[3]),
    .ADR2(DLX_IDinst_IR_opcode_field[3]),
    .ADR3(CHOICE3166),
    .O(\CHOICE3166/GROM )
  );
  X_BUF \CHOICE3166/XUSED  (
    .I(\CHOICE3166/FROM ),
    .O(CHOICE3166)
  );
  X_BUF \CHOICE3166/YUSED  (
    .I(\CHOICE3166/GROM ),
    .O(CHOICE3168)
  );
  defparam DLX_EXinst_Ker6582050.INIT = 16'hFFA8;
  X_LUT4 DLX_EXinst_Ker6582050 (
    .ADR0(N110065),
    .ADR1(CHOICE2043),
    .ADR2(CHOICE2046),
    .ADR3(CHOICE2051),
    .O(\N102162/FROM )
  );
  defparam \DLX_EXinst__n0006<29>115 .INIT = 16'hFDFC;
  X_LUT4 \DLX_EXinst__n0006<29>115  (
    .ADR0(DLX_IDinst_IR_function_field[4]),
    .ADR1(CHOICE5355),
    .ADR2(CHOICE5333),
    .ADR3(N102162),
    .O(\N102162/GROM )
  );
  X_BUF \N102162/XUSED  (
    .I(\N102162/FROM ),
    .O(N102162)
  );
  X_BUF \N102162/YUSED  (
    .I(\N102162/GROM ),
    .O(CHOICE5356)
  );
  defparam DLX_IDinst_Ker699798.INIT = 16'h00CC;
  X_LUT4 DLX_IDinst_Ker699798 (
    .ADR0(VCC),
    .ADR1(DLX_opcode_of_MEM[4]),
    .ADR2(VCC),
    .ADR3(DLX_opcode_of_MEM[5]),
    .O(\CHOICE1452/FROM )
  );
  defparam DLX_IDinst_Ker6997912.INIT = 16'hC400;
  X_LUT4 DLX_IDinst_Ker6997912 (
    .ADR0(DLX_opcode_of_MEM[0]),
    .ADR1(DLX_opcode_of_MEM[2]),
    .ADR2(DLX_opcode_of_MEM[1]),
    .ADR3(CHOICE1452),
    .O(\CHOICE1452/GROM )
  );
  X_BUF \CHOICE1452/XUSED  (
    .I(\CHOICE1452/FROM ),
    .O(CHOICE1452)
  );
  X_BUF \CHOICE1452/YUSED  (
    .I(\CHOICE1452/GROM ),
    .O(CHOICE1453)
  );
  defparam DLX_cg3_c1.INIT = 16'hFBB0;
  X_LUT4 DLX_cg3_c1 (
    .ADR0(DLX_EXlc_md_outp2),
    .ADR1(CHOICE12),
    .ADR2(DLX_clk_IF),
    .ADR3(DLX_ackout_ID),
    .O(\DLX_ackout_ID/FROM )
  );
  defparam DLX_EXlc_master_ctrlEX__n0001_SW111.INIT = 16'hFF33;
  X_LUT4 DLX_EXlc_master_ctrlEX__n0001_SW111 (
    .ADR0(VCC),
    .ADR1(CHOICE12),
    .ADR2(VCC),
    .ADR3(DLX_EXlc_md_outp2),
    .O(\DLX_ackout_ID/GROM )
  );
  X_BUF \DLX_ackout_ID/XUSED  (
    .I(\DLX_ackout_ID/FROM ),
    .O(DLX_ackout_ID)
  );
  X_BUF \DLX_ackout_ID/YUSED  (
    .I(\DLX_ackout_ID/GROM ),
    .O(DLX_ackin_EX)
  );
  defparam DLX_EXlc_md_mda20_a1.INIT = 16'h0A0A;
  X_LUT4 DLX_EXlc_md_mda20_a1 (
    .ADR0(DLX_EXlc_md_wint19),
    .ADR1(VCC),
    .ADR2(DLX_EXlc_pd_wint5),
    .ADR3(VCC),
    .O(\DLX_EXlc_md_wint20/FROM )
  );
  defparam DLX_EXlc_md_mda11_a1.INIT = 16'h3300;
  X_LUT4 DLX_EXlc_md_mda11_a1 (
    .ADR0(VCC),
    .ADR1(DLX_EXlc_pd_wint5),
    .ADR2(VCC),
    .ADR3(DLX_EXlc_md_wint10),
    .O(\DLX_EXlc_md_wint20/GROM )
  );
  X_BUF \DLX_EXlc_md_wint20/XUSED  (
    .I(\DLX_EXlc_md_wint20/FROM ),
    .O(DLX_EXlc_md_wint20)
  );
  X_BUF \DLX_EXlc_md_wint20/YUSED  (
    .I(\DLX_EXlc_md_wint20/GROM ),
    .O(DLX_EXlc_md_wint11)
  );
  defparam \DLX_EXinst__n0006<31>524 .INIT = 16'h5D0C;
  X_LUT4 \DLX_EXinst__n0006<31>524  (
    .ADR0(\DLX_IDinst_Imm[31] ),
    .ADR1(N110065),
    .ADR2(\DLX_IDinst_Imm[5] ),
    .ADR3(DLX_EXinst__n0080),
    .O(\CHOICE5839/FROM )
  );
  defparam DLX_EXinst_Ker63687_SW0.INIT = 16'h7FFF;
  X_LUT4 DLX_EXinst_Ker63687_SW0 (
    .ADR0(\DLX_IDinst_Imm[5] ),
    .ADR1(N110065),
    .ADR2(DLX_EXinst__n0149),
    .ADR3(DLX_IDinst_reg_out_A[31]),
    .O(\CHOICE5839/GROM )
  );
  X_BUF \CHOICE5839/XUSED  (
    .I(\CHOICE5839/FROM ),
    .O(CHOICE5839)
  );
  X_BUF \CHOICE5839/YUSED  (
    .I(\CHOICE5839/GROM ),
    .O(N101919)
  );
  defparam DLX_EXinst_Ker6538950.INIT = 16'hFFA8;
  X_LUT4 DLX_EXinst_Ker6538950 (
    .ADR0(N110065),
    .ADR1(CHOICE1359),
    .ADR2(CHOICE1356),
    .ADR3(CHOICE1364),
    .O(\N98127/FROM )
  );
  defparam \DLX_EXinst__n0006<8>84 .INIT = 16'hFEEE;
  X_LUT4 \DLX_EXinst__n0006<8>84  (
    .ADR0(CHOICE3684),
    .ADR1(CHOICE3699),
    .ADR2(DLX_IDinst_IR_function_field[4]),
    .ADR3(N98127),
    .O(\N98127/GROM )
  );
  X_BUF \N98127/XUSED  (
    .I(\N98127/FROM ),
    .O(N98127)
  );
  X_BUF \N98127/YUSED  (
    .I(\N98127/GROM ),
    .O(CHOICE3700)
  );
  defparam \DLX_EXinst_Mshift__n0028_Sh<51>1 .INIT = 16'hE2E2;
  X_LUT4 \DLX_EXinst_Mshift__n0028_Sh<51>1  (
    .ADR0(DLX_EXinst_N64849),
    .ADR1(DLX_IDinst_IR_function_field_2_1),
    .ADR2(DLX_EXinst_N63031),
    .ADR3(VCC),
    .O(\DLX_EXinst_Mshift__n0028_Sh<51>/FROM )
  );
  defparam DLX_EXinst_Ker6582047.INIT = 16'h0008;
  X_LUT4 DLX_EXinst_Ker6582047 (
    .ADR0(\DLX_EXinst_Mshift__n0028_Sh[29] ),
    .ADR1(DLX_EXinst_N66507),
    .ADR2(DLX_IDinst_IR_function_field_2_1),
    .ADR3(DLX_IDinst_IR_function_field_3_1),
    .O(\DLX_EXinst_Mshift__n0028_Sh<51>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0028_Sh<51>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0028_Sh<51>/FROM ),
    .O(\DLX_EXinst_Mshift__n0028_Sh[51] )
  );
  X_BUF \DLX_EXinst_Mshift__n0028_Sh<51>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0028_Sh<51>/GROM ),
    .O(CHOICE2051)
  );
  defparam DLX_EXinst__n003512.INIT = 16'hFFFE;
  X_LUT4 DLX_EXinst__n003512 (
    .ADR0(DLX_IDinst_reg_out_B[27]),
    .ADR1(DLX_IDinst_reg_out_B[24]),
    .ADR2(DLX_IDinst_reg_out_B[25]),
    .ADR3(DLX_IDinst_reg_out_B[26]),
    .O(\CHOICE3539/FROM )
  );
  defparam DLX_EXinst__n003515.INIT = 16'hFFFE;
  X_LUT4 DLX_EXinst__n003515 (
    .ADR0(DLX_IDinst_reg_out_B[29]),
    .ADR1(DLX_IDinst_reg_out_B[28]),
    .ADR2(DLX_IDinst_reg_out_B[30]),
    .ADR3(CHOICE3539),
    .O(\CHOICE3539/GROM )
  );
  X_BUF \CHOICE3539/XUSED  (
    .I(\CHOICE3539/FROM ),
    .O(CHOICE3539)
  );
  X_BUF \CHOICE3539/YUSED  (
    .I(\CHOICE3539/GROM ),
    .O(CHOICE3540)
  );
  defparam \DLX_EXinst__n0006<24>223_SW0 .INIT = 16'hD5C0;
  X_LUT4 \DLX_EXinst__n0006<24>223_SW0  (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(DLX_EXinst_ALU_result[24]),
    .ADR2(N101725),
    .ADR3(N98218),
    .O(\N126546/FROM )
  );
  defparam \DLX_EXinst__n0006<26>240_SW0 .INIT = 16'h88F8;
  X_LUT4 \DLX_EXinst__n0006<26>240_SW0  (
    .ADR0(DLX_EXinst_ALU_result[26]),
    .ADR1(N101725),
    .ADR2(N107934),
    .ADR3(DLX_IDinst_reg_out_B[4]),
    .O(\N126546/GROM )
  );
  X_BUF \N126546/XUSED  (
    .I(\N126546/FROM ),
    .O(N126546)
  );
  X_BUF \N126546/YUSED  (
    .I(\N126546/GROM ),
    .O(N126354)
  );
  defparam \DLX_EXinst__n0006<11>161 .INIT = 16'hAC00;
  X_LUT4 \DLX_EXinst__n0006<11>161  (
    .ADR0(N97449),
    .ADR1(DLX_EXinst_N65160),
    .ADR2(DLX_IDinst_reg_out_B[2]),
    .ADR3(DLX_EXinst_N62631),
    .O(\CHOICE3957/FROM )
  );
  defparam \DLX_EXinst__n0006<7>147 .INIT = 16'h8A80;
  X_LUT4 \DLX_EXinst__n0006<7>147  (
    .ADR0(DLX_EXinst_N62631),
    .ADR1(DLX_EXinst_N65160),
    .ADR2(DLX_IDinst_reg_out_B[2]),
    .ADR3(N96945),
    .O(\CHOICE3957/GROM )
  );
  X_BUF \CHOICE3957/XUSED  (
    .I(\CHOICE3957/FROM ),
    .O(CHOICE3957)
  );
  X_BUF \CHOICE3957/YUSED  (
    .I(\CHOICE3957/GROM ),
    .O(CHOICE3833)
  );
  defparam DLX_EXinst_Ker6581513.INIT = 16'h8000;
  X_LUT4 DLX_EXinst_Ker6581513 (
    .ADR0(CHOICE3377),
    .ADR1(\DLX_IDinst_Imm[5] ),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(CHOICE3408),
    .O(\CHOICE2077/FROM )
  );
  defparam DLX_EXinst_Ker6581535.INIT = 16'h0302;
  X_LUT4 DLX_EXinst_Ker6581535 (
    .ADR0(CHOICE2075),
    .ADR1(DLX_IDinst_IR_function_field_3_1),
    .ADR2(DLX_IDinst_IR_function_field_2_1),
    .ADR3(CHOICE2077),
    .O(\CHOICE2077/GROM )
  );
  X_BUF \CHOICE2077/XUSED  (
    .I(\CHOICE2077/FROM ),
    .O(CHOICE2077)
  );
  X_BUF \CHOICE2077/YUSED  (
    .I(\CHOICE2077/GROM ),
    .O(CHOICE2081)
  );
  defparam \DLX_EXinst__n0006<7>228 .INIT = 16'hFE00;
  X_LUT4 \DLX_EXinst__n0006<7>228  (
    .ADR0(N126465),
    .ADR1(CHOICE3828),
    .ADR2(CHOICE3844),
    .ADR3(DLX_EXinst__n0030_1),
    .O(\CHOICE3850/FROM )
  );
  defparam \DLX_EXinst__n0006<7>240 .INIT = 16'hFF88;
  X_LUT4 \DLX_EXinst__n0006<7>240  (
    .ADR0(DLX_EXinst_N63836),
    .ADR1(DLX_EXinst__n0016[7]),
    .ADR2(VCC),
    .ADR3(CHOICE3850),
    .O(\CHOICE3850/GROM )
  );
  X_BUF \CHOICE3850/XUSED  (
    .I(\CHOICE3850/FROM ),
    .O(CHOICE3850)
  );
  X_BUF \CHOICE3850/YUSED  (
    .I(\CHOICE3850/GROM ),
    .O(CHOICE3851)
  );
  defparam DLX_IDinst_Mmux__n0148_inst_mux_f5_301.INIT = 16'hF022;
  X_LUT4 DLX_IDinst_Mmux__n0148_inst_mux_f5_301 (
    .ADR0(DLX_RF_data_in[7]),
    .ADR1(DLX_opcode_of_WB[2]),
    .ADR2(DLX_MEMinst_RF_data_in[15]),
    .ADR3(DLX_opcode_of_WB[0]),
    .O(\DLX_IDinst__n0445<47>/FROM )
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<15>1 .INIT = 16'hEE44;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<15>1  (
    .ADR0(DLX_IDinst__n0147),
    .ADR1(DLX_MEMinst_RF_data_in[15]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst__n0445[47]),
    .O(\DLX_IDinst__n0445<47>/GROM )
  );
  X_BUF \DLX_IDinst__n0445<47>/XUSED  (
    .I(\DLX_IDinst__n0445<47>/FROM ),
    .O(DLX_IDinst__n0445[47])
  );
  X_BUF \DLX_IDinst__n0445<47>/YUSED  (
    .I(\DLX_IDinst__n0445<47>/GROM ),
    .O(DLX_IDinst_WB_data_eff[15])
  );
  defparam DLX_EXlc_md_mda19_a1.INIT = 16'h0A0A;
  X_LUT4 DLX_EXlc_md_mda19_a1 (
    .ADR0(DLX_EXlc_md_wint18),
    .ADR1(VCC),
    .ADR2(DLX_EXlc_pd_wint5),
    .ADR3(VCC),
    .O(\DLX_EXlc_md_wint19/FROM )
  );
  defparam DLX_EXlc_md_mda12_a1.INIT = 16'h0C0C;
  X_LUT4 DLX_EXlc_md_mda12_a1 (
    .ADR0(VCC),
    .ADR1(DLX_EXlc_md_wint11),
    .ADR2(DLX_EXlc_pd_wint5),
    .ADR3(VCC),
    .O(\DLX_EXlc_md_wint19/GROM )
  );
  X_BUF \DLX_EXlc_md_wint19/XUSED  (
    .I(\DLX_EXlc_md_wint19/FROM ),
    .O(DLX_EXlc_md_wint19)
  );
  X_BUF \DLX_EXlc_md_wint19/YUSED  (
    .I(\DLX_EXlc_md_wint19/GROM ),
    .O(DLX_EXlc_md_wint12)
  );
  defparam DLX_EXinst_Ker6581550.INIT = 16'hFFCC;
  X_LUT4 DLX_EXinst_Ker6581550 (
    .ADR0(VCC),
    .ADR1(CHOICE2081),
    .ADR2(VCC),
    .ADR3(CHOICE2085),
    .O(\N102358/FROM )
  );
  defparam \DLX_EXinst__n0006<28>115 .INIT = 16'hEEFE;
  X_LUT4 \DLX_EXinst__n0006<28>115  (
    .ADR0(CHOICE5181),
    .ADR1(CHOICE5203),
    .ADR2(N102358),
    .ADR3(DLX_IDinst_IR_function_field[4]),
    .O(\N102358/GROM )
  );
  X_BUF \N102358/XUSED  (
    .I(\N102358/FROM ),
    .O(N102358)
  );
  X_BUF \N102358/YUSED  (
    .I(\N102358/GROM ),
    .O(CHOICE5204)
  );
  defparam DLX_IDinst_Mmux__n0148_inst_mux_f5_231.INIT = 16'hA0AC;
  X_LUT4 DLX_IDinst_Mmux__n0148_inst_mux_f5_231 (
    .ADR0(DLX_MEMinst_RF_data_in[8]),
    .ADR1(DLX_RF_data_in[7]),
    .ADR2(DLX_opcode_of_WB[0]),
    .ADR3(DLX_opcode_of_WB[2]),
    .O(\DLX_IDinst__n0445<40>/FROM )
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<8>1 .INIT = 16'hFA0A;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<8>1  (
    .ADR0(DLX_MEMinst_RF_data_in[8]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst__n0147),
    .ADR3(DLX_IDinst__n0445[40]),
    .O(\DLX_IDinst__n0445<40>/GROM )
  );
  X_BUF \DLX_IDinst__n0445<40>/XUSED  (
    .I(\DLX_IDinst__n0445<40>/FROM ),
    .O(DLX_IDinst__n0445[40])
  );
  X_BUF \DLX_IDinst__n0445<40>/YUSED  (
    .I(\DLX_IDinst__n0445<40>/GROM ),
    .O(DLX_IDinst_WB_data_eff[8])
  );
  defparam DLX_IDinst_Mmux__n0148_inst_mux_f5_241.INIT = 16'hAA30;
  X_LUT4 DLX_IDinst_Mmux__n0148_inst_mux_f5_241 (
    .ADR0(DLX_MEMinst_RF_data_in[9]),
    .ADR1(DLX_opcode_of_WB[2]),
    .ADR2(DLX_RF_data_in[7]),
    .ADR3(DLX_opcode_of_WB[0]),
    .O(\DLX_IDinst__n0445<41>/FROM )
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<9>1 .INIT = 16'hEE44;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<9>1  (
    .ADR0(DLX_IDinst__n0147),
    .ADR1(DLX_MEMinst_RF_data_in[9]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst__n0445[41]),
    .O(\DLX_IDinst__n0445<41>/GROM )
  );
  X_BUF \DLX_IDinst__n0445<41>/XUSED  (
    .I(\DLX_IDinst__n0445<41>/FROM ),
    .O(DLX_IDinst__n0445[41])
  );
  X_BUF \DLX_IDinst__n0445<41>/YUSED  (
    .I(\DLX_IDinst__n0445<41>/GROM ),
    .O(DLX_IDinst_WB_data_eff[9])
  );
  defparam DLX_IDinst__n00021.INIT = 16'h0404;
  X_LUT4 DLX_IDinst__n00021 (
    .ADR0(DLX_IDinst_regA_index[0]),
    .ADR1(DLX_IDinst_N70658),
    .ADR2(DLX_IDinst_regA_index[1]),
    .ADR3(VCC),
    .O(\DLX_IDinst__n0002/FROM )
  );
  defparam DLX_IDinst_Ker7066682.INIT = 16'hF010;
  X_LUT4 DLX_IDinst_Ker7066682 (
    .ADR0(DLX_IDinst__n0077),
    .ADR1(DLX_IDinst__n0073),
    .ADR2(CHOICE3274),
    .ADR3(DLX_IDinst__n0002),
    .O(\DLX_IDinst__n0002/GROM )
  );
  X_BUF \DLX_IDinst__n0002/XUSED  (
    .I(\DLX_IDinst__n0002/FROM ),
    .O(DLX_IDinst__n0002)
  );
  X_BUF \DLX_IDinst__n0002/YUSED  (
    .I(\DLX_IDinst__n0002/GROM ),
    .O(CHOICE3275)
  );
  defparam \DLX_EXinst__n0006<8>115 .INIT = 16'hEECC;
  X_LUT4 \DLX_EXinst__n0006<8>115  (
    .ADR0(DLX_IDinst_reg_out_B[8]),
    .ADR1(DLX_EXinst_N64448),
    .ADR2(VCC),
    .ADR3(DLX_EXinst__n0045),
    .O(\CHOICE3706/FROM )
  );
  defparam \DLX_EXinst__n0006<8>124 .INIT = 16'hF020;
  X_LUT4 \DLX_EXinst__n0006<8>124  (
    .ADR0(DLX_EXinst__n0047),
    .ADR1(DLX_IDinst_reg_out_B[8]),
    .ADR2(DLX_IDinst_reg_out_A[8]),
    .ADR3(CHOICE3706),
    .O(\CHOICE3706/GROM )
  );
  X_BUF \CHOICE3706/XUSED  (
    .I(\CHOICE3706/FROM ),
    .O(CHOICE3706)
  );
  X_BUF \CHOICE3706/YUSED  (
    .I(\CHOICE3706/GROM ),
    .O(CHOICE3708)
  );
  defparam \DLX_EXinst__n0006<7>268 .INIT = 16'hCE00;
  X_LUT4 \DLX_EXinst__n0006<7>268  (
    .ADR0(CHOICE3820),
    .ADR1(CHOICE3851),
    .ADR2(DLX_EXinst__n0030_1),
    .ADR3(DLX_EXinst__n0149),
    .O(\DLX_EXinst_ALU_result<7>/FROM )
  );
  defparam \DLX_EXinst__n0006<7>278 .INIT = 16'hFFF0;
  X_LUT4 \DLX_EXinst__n0006<7>278  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N63689),
    .ADR3(CHOICE3853),
    .O(\DLX_EXinst_ALU_result<7>/GROM )
  );
  X_BUF \DLX_EXinst_ALU_result<7>/XUSED  (
    .I(\DLX_EXinst_ALU_result<7>/FROM ),
    .O(CHOICE3853)
  );
  X_BUF \DLX_EXinst_ALU_result<7>/YUSED  (
    .I(\DLX_EXinst_ALU_result<7>/GROM ),
    .O(N112616)
  );
  defparam DLX_EXinst_Ker66248116.INIT = 16'h0001;
  X_LUT4 DLX_EXinst_Ker66248116 (
    .ADR0(\DLX_IDinst_Imm[13] ),
    .ADR1(\DLX_IDinst_Imm[11] ),
    .ADR2(\DLX_IDinst_Imm[12] ),
    .ADR3(\DLX_IDinst_Imm[14] ),
    .O(\CHOICE3399/FROM )
  );
  defparam DLX_EXinst__n003650.INIT = 16'hFFFE;
  X_LUT4 DLX_EXinst__n003650 (
    .ADR0(\DLX_IDinst_Imm[12] ),
    .ADR1(\DLX_IDinst_Imm[13] ),
    .ADR2(\DLX_IDinst_Imm[14] ),
    .ADR3(\DLX_IDinst_Imm[15] ),
    .O(\CHOICE3399/GROM )
  );
  X_BUF \CHOICE3399/XUSED  (
    .I(\CHOICE3399/FROM ),
    .O(CHOICE3399)
  );
  X_BUF \CHOICE3399/YUSED  (
    .I(\CHOICE3399/GROM ),
    .O(CHOICE3246)
  );
  defparam DLX_IDinst_Mmux__n0148_inst_mux_f5_251.INIT = 16'hC0E2;
  X_LUT4 DLX_IDinst_Mmux__n0148_inst_mux_f5_251 (
    .ADR0(DLX_RF_data_in[7]),
    .ADR1(DLX_opcode_of_WB[0]),
    .ADR2(DLX_MEMinst_RF_data_in[10]),
    .ADR3(DLX_opcode_of_WB[2]),
    .O(\DLX_IDinst__n0445<42>/FROM )
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<10>1 .INIT = 16'hFA50;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<10>1  (
    .ADR0(DLX_IDinst__n0147),
    .ADR1(VCC),
    .ADR2(DLX_MEMinst_RF_data_in[10]),
    .ADR3(DLX_IDinst__n0445[42]),
    .O(\DLX_IDinst__n0445<42>/GROM )
  );
  X_BUF \DLX_IDinst__n0445<42>/XUSED  (
    .I(\DLX_IDinst__n0445<42>/FROM ),
    .O(DLX_IDinst__n0445[42])
  );
  X_BUF \DLX_IDinst__n0445<42>/YUSED  (
    .I(\DLX_IDinst__n0445<42>/GROM ),
    .O(DLX_IDinst_WB_data_eff[10])
  );
  defparam DLX_EXinst__n003555.INIT = 16'hFFFE;
  X_LUT4 DLX_EXinst__n003555 (
    .ADR0(DLX_IDinst_reg_out_B[11]),
    .ADR1(DLX_IDinst_reg_out_B[9]),
    .ADR2(DLX_IDinst_reg_out_B[8]),
    .ADR3(DLX_IDinst_reg_out_B[10]),
    .O(\CHOICE3554/FROM )
  );
  defparam DLX_EXinst__n003564_SW0.INIT = 16'hFFFE;
  X_LUT4 DLX_EXinst__n003564_SW0 (
    .ADR0(DLX_IDinst_reg_out_B[20]),
    .ADR1(CHOICE3551),
    .ADR2(CHOICE3547),
    .ADR3(CHOICE3554),
    .O(\CHOICE3554/GROM )
  );
  X_BUF \CHOICE3554/XUSED  (
    .I(\CHOICE3554/FROM ),
    .O(CHOICE3554)
  );
  X_BUF \CHOICE3554/YUSED  (
    .I(\CHOICE3554/GROM ),
    .O(N126510)
  );
  defparam DLX_EXinst_Ker6628835.INIT = 16'h0504;
  X_LUT4 DLX_EXinst_Ker6628835 (
    .ADR0(DLX_EXinst__n0030_1),
    .ADR1(CHOICE1757),
    .ADR2(DLX_IDinst_IR_opcode_field[4]),
    .ADR3(CHOICE1758),
    .O(\N100440/FROM )
  );
  defparam \DLX_EXinst__n0017<16>1 .INIT = 16'hF888;
  X_LUT4 \DLX_EXinst__n0017<16>1  (
    .ADR0(DLX_IDinst_reg_out_B[16]),
    .ADR1(DLX_EXinst__n0030_1),
    .ADR2(\DLX_IDinst_Imm[31] ),
    .ADR3(N100440),
    .O(\N100440/GROM )
  );
  X_BUF \N100440/XUSED  (
    .I(\N100440/FROM ),
    .O(N100440)
  );
  X_BUF \N100440/YUSED  (
    .I(\N100440/GROM ),
    .O(DLX_EXinst__n0017[16])
  );
  defparam DLX_EXinst__n003564.INIT = 16'hFFFE;
  X_LUT4 DLX_EXinst__n003564 (
    .ADR0(DLX_IDinst_reg_out_B[21]),
    .ADR1(DLX_IDinst_reg_out_B[22]),
    .ADR2(DLX_IDinst_reg_out_B[23]),
    .ADR3(N126510),
    .O(\CHOICE3556/FROM )
  );
  defparam DLX_EXinst__n003575.INIT = 16'hFFEE;
  X_LUT4 DLX_EXinst__n003575 (
    .ADR0(CHOICE3534),
    .ADR1(CHOICE3540),
    .ADR2(VCC),
    .ADR3(CHOICE3556),
    .O(\CHOICE3556/GROM )
  );
  X_BUF \CHOICE3556/XUSED  (
    .I(\CHOICE3556/FROM ),
    .O(CHOICE3556)
  );
  X_BUF \CHOICE3556/YUSED  (
    .I(\CHOICE3556/GROM ),
    .O(N110935)
  );
  defparam DLX_IDinst_Mmux__n0148_inst_mux_f5_261.INIT = 16'hC5C0;
  X_LUT4 DLX_IDinst_Mmux__n0148_inst_mux_f5_261 (
    .ADR0(DLX_opcode_of_WB[2]),
    .ADR1(DLX_MEMinst_RF_data_in[11]),
    .ADR2(DLX_opcode_of_WB[0]),
    .ADR3(DLX_RF_data_in[7]),
    .O(\DLX_IDinst__n0445<43>/FROM )
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<11>1 .INIT = 16'hEE22;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<11>1  (
    .ADR0(DLX_MEMinst_RF_data_in[11]),
    .ADR1(DLX_IDinst__n0147),
    .ADR2(VCC),
    .ADR3(DLX_IDinst__n0445[43]),
    .O(\DLX_IDinst__n0445<43>/GROM )
  );
  X_BUF \DLX_IDinst__n0445<43>/XUSED  (
    .I(\DLX_IDinst__n0445<43>/FROM ),
    .O(DLX_IDinst__n0445[43])
  );
  X_BUF \DLX_IDinst__n0445<43>/YUSED  (
    .I(\DLX_IDinst__n0445<43>/GROM ),
    .O(DLX_IDinst_WB_data_eff[11])
  );
  defparam DLX_EXinst_Ker6486711.INIT = 16'hE400;
  X_LUT4 DLX_EXinst_Ker6486711 (
    .ADR0(DLX_IDinst_reg_out_B_3_1),
    .ADR1(\DLX_EXinst_Mshift__n0023_Sh[25] ),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(DLX_IDinst_reg_out_B_2_1),
    .O(\CHOICE3112/FROM )
  );
  defparam DLX_EXinst_Ker6488212.INIT = 16'h8C80;
  X_LUT4 DLX_EXinst_Ker6488212 (
    .ADR0(\DLX_EXinst_Mshift__n0023_Sh[61] ),
    .ADR1(DLX_IDinst_reg_out_B[5]),
    .ADR2(DLX_IDinst_reg_out_B_2_1),
    .ADR3(DLX_IDinst_reg_out_A[31]),
    .O(\CHOICE3112/GROM )
  );
  X_BUF \CHOICE3112/XUSED  (
    .I(\CHOICE3112/FROM ),
    .O(CHOICE3112)
  );
  X_BUF \CHOICE3112/YUSED  (
    .I(\CHOICE3112/GROM ),
    .O(CHOICE3139)
  );
  defparam DLX_EXlc_md_mda18_a1.INIT = 16'h3300;
  X_LUT4 DLX_EXlc_md_mda18_a1 (
    .ADR0(VCC),
    .ADR1(DLX_EXlc_pd_wint5),
    .ADR2(VCC),
    .ADR3(DLX_EXlc_md_wint17),
    .O(\DLX_EXlc_md_wint18/FROM )
  );
  defparam DLX_EXlc_md_mda13_a1.INIT = 16'h5500;
  X_LUT4 DLX_EXlc_md_mda13_a1 (
    .ADR0(DLX_EXlc_pd_wint5),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_EXlc_md_wint12),
    .O(\DLX_EXlc_md_wint18/GROM )
  );
  X_BUF \DLX_EXlc_md_wint18/XUSED  (
    .I(\DLX_EXlc_md_wint18/FROM ),
    .O(DLX_EXlc_md_wint18)
  );
  X_BUF \DLX_EXlc_md_wint18/YUSED  (
    .I(\DLX_EXlc_md_wint18/GROM ),
    .O(DLX_EXlc_md_wint13)
  );
  defparam DLX_IDinst_Mmux__n0148_inst_mux_f5_271.INIT = 16'hF202;
  X_LUT4 DLX_IDinst_Mmux__n0148_inst_mux_f5_271 (
    .ADR0(DLX_RF_data_in[7]),
    .ADR1(DLX_opcode_of_WB[2]),
    .ADR2(DLX_opcode_of_WB[0]),
    .ADR3(DLX_MEMinst_RF_data_in[12]),
    .O(\DLX_IDinst__n0445<44>/FROM )
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<12>1 .INIT = 16'hFA50;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<12>1  (
    .ADR0(DLX_IDinst__n0147),
    .ADR1(VCC),
    .ADR2(DLX_MEMinst_RF_data_in[12]),
    .ADR3(DLX_IDinst__n0445[44]),
    .O(\DLX_IDinst__n0445<44>/GROM )
  );
  X_BUF \DLX_IDinst__n0445<44>/XUSED  (
    .I(\DLX_IDinst__n0445<44>/FROM ),
    .O(DLX_IDinst__n0445[44])
  );
  X_BUF \DLX_IDinst__n0445<44>/YUSED  (
    .I(\DLX_IDinst__n0445<44>/GROM ),
    .O(DLX_IDinst_WB_data_eff[12])
  );
  defparam \DLX_EXinst__n0006<8>209 .INIT = 16'hCCC8;
  X_LUT4 \DLX_EXinst__n0006<8>209  (
    .ADR0(CHOICE3717),
    .ADR1(DLX_EXinst__n0030_1),
    .ADR2(CHOICE3726),
    .ADR3(CHOICE3708),
    .O(\CHOICE3728/FROM )
  );
  defparam \DLX_EXinst__n0006<8>221 .INIT = 16'hFFC0;
  X_LUT4 \DLX_EXinst__n0006<8>221  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst__n0016[8]),
    .ADR2(DLX_EXinst_N63836),
    .ADR3(CHOICE3728),
    .O(\CHOICE3728/GROM )
  );
  X_BUF \CHOICE3728/XUSED  (
    .I(\CHOICE3728/FROM ),
    .O(CHOICE3728)
  );
  X_BUF \CHOICE3728/YUSED  (
    .I(\CHOICE3728/GROM ),
    .O(CHOICE3729)
  );
  defparam DLX_EXinst__n003655.INIT = 16'hFFFE;
  X_LUT4 DLX_EXinst__n003655 (
    .ADR0(\DLX_IDinst_Imm[11] ),
    .ADR1(\DLX_IDinst_Imm[9] ),
    .ADR2(\DLX_IDinst_Imm[8] ),
    .ADR3(\DLX_IDinst_Imm[10] ),
    .O(\CHOICE3249/GROM )
  );
  X_BUF \CHOICE3249/YUSED  (
    .I(\CHOICE3249/GROM ),
    .O(CHOICE3249)
  );
  defparam \DLX_EXinst__n0006<8>137 .INIT = 16'hC0A0;
  X_LUT4 \DLX_EXinst__n0006<8>137  (
    .ADR0(DLX_EXinst_N64804),
    .ADR1(N97375),
    .ADR2(DLX_EXinst_N62631),
    .ADR3(DLX_IDinst_reg_out_B[2]),
    .O(\CHOICE3713/FROM )
  );
  defparam \DLX_EXinst__n0006<8>151 .INIT = 16'h5540;
  X_LUT4 \DLX_EXinst__n0006<8>151  (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(DLX_EXinst_N66226),
    .ADR2(\DLX_EXinst_Mshift__n0025_Sh[40] ),
    .ADR3(CHOICE3713),
    .O(\CHOICE3713/GROM )
  );
  X_BUF \CHOICE3713/XUSED  (
    .I(\CHOICE3713/FROM ),
    .O(CHOICE3713)
  );
  X_BUF \CHOICE3713/YUSED  (
    .I(\CHOICE3713/GROM ),
    .O(CHOICE3717)
  );
  defparam DLX_IDinst_Mmux__n0148_inst_mux_f5_281.INIT = 16'hDC10;
  X_LUT4 DLX_IDinst_Mmux__n0148_inst_mux_f5_281 (
    .ADR0(DLX_opcode_of_WB[2]),
    .ADR1(DLX_opcode_of_WB[0]),
    .ADR2(DLX_RF_data_in[7]),
    .ADR3(DLX_MEMinst_RF_data_in[13]),
    .O(\DLX_IDinst__n0445<45>/FROM )
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<13>1 .INIT = 16'hEE44;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<13>1  (
    .ADR0(DLX_IDinst__n0147),
    .ADR1(DLX_MEMinst_RF_data_in[13]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst__n0445[45]),
    .O(\DLX_IDinst__n0445<45>/GROM )
  );
  X_BUF \DLX_IDinst__n0445<45>/XUSED  (
    .I(\DLX_IDinst__n0445<45>/FROM ),
    .O(DLX_IDinst__n0445[45])
  );
  X_BUF \DLX_IDinst__n0445<45>/YUSED  (
    .I(\DLX_IDinst__n0445<45>/GROM ),
    .O(DLX_IDinst_WB_data_eff[13])
  );
  defparam \DLX_EXinst__n0006<21>152 .INIT = 16'hF040;
  X_LUT4 \DLX_EXinst__n0006<21>152  (
    .ADR0(DLX_IDinst_reg_out_A[21]),
    .ADR1(DLX_EXinst__n0047),
    .ADR2(DLX_IDinst_reg_out_B[21]),
    .ADR3(DLX_EXinst__n0046),
    .O(\CHOICE4196/FROM )
  );
  defparam \DLX_EXinst__n0006<8>180 .INIT = 16'hA2A0;
  X_LUT4 \DLX_EXinst__n0006<8>180  (
    .ADR0(DLX_IDinst_reg_out_B[8]),
    .ADR1(DLX_IDinst_reg_out_A[8]),
    .ADR2(DLX_EXinst__n0046),
    .ADR3(DLX_EXinst__n0047),
    .O(\CHOICE4196/GROM )
  );
  X_BUF \CHOICE4196/XUSED  (
    .I(\CHOICE4196/FROM ),
    .O(CHOICE4196)
  );
  X_BUF \CHOICE4196/YUSED  (
    .I(\CHOICE4196/GROM ),
    .O(CHOICE3722)
  );
  defparam DLX_IDinst_Mmux__n0148_inst_mux_f5_291.INIT = 16'h8B88;
  X_LUT4 DLX_IDinst_Mmux__n0148_inst_mux_f5_291 (
    .ADR0(DLX_MEMinst_RF_data_in[14]),
    .ADR1(DLX_opcode_of_WB[0]),
    .ADR2(DLX_opcode_of_WB[2]),
    .ADR3(DLX_RF_data_in[7]),
    .O(\DLX_IDinst__n0445<46>/FROM )
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<14>1 .INIT = 16'hEE22;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<14>1  (
    .ADR0(DLX_MEMinst_RF_data_in[14]),
    .ADR1(DLX_IDinst__n0147),
    .ADR2(VCC),
    .ADR3(DLX_IDinst__n0445[46]),
    .O(\DLX_IDinst__n0445<46>/GROM )
  );
  X_BUF \DLX_IDinst__n0445<46>/XUSED  (
    .I(\DLX_IDinst__n0445<46>/FROM ),
    .O(DLX_IDinst__n0445[46])
  );
  X_BUF \DLX_IDinst__n0445<46>/YUSED  (
    .I(\DLX_IDinst__n0445<46>/GROM ),
    .O(DLX_IDinst_WB_data_eff[14])
  );
  defparam DLX_EXlc_md_mda30_a1.INIT = 16'h0F00;
  X_LUT4 DLX_EXlc_md_mda30_a1 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_EXlc_pd_wint5),
    .ADR3(DLX_EXlc_md_wint29),
    .O(\DLX_EXlc_md_wint30/FROM )
  );
  defparam DLX_EXlc_md_mda31_a1.INIT = 16'h0F00;
  X_LUT4 DLX_EXlc_md_mda31_a1 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_EXlc_pd_wint5),
    .ADR3(DLX_EXlc_md_wint30),
    .O(\DLX_EXlc_md_wint30/GROM )
  );
  X_BUF \DLX_EXlc_md_wint30/XUSED  (
    .I(\DLX_EXlc_md_wint30/FROM ),
    .O(DLX_EXlc_md_wint30)
  );
  X_BUF \DLX_EXlc_md_wint30/YUSED  (
    .I(\DLX_EXlc_md_wint30/GROM ),
    .O(DLX_EXlc_md_wint31)
  );
  defparam DLX_EXlc_md_mda17_a1.INIT = 16'h4444;
  X_LUT4 DLX_EXlc_md_mda17_a1 (
    .ADR0(DLX_EXlc_pd_wint5),
    .ADR1(DLX_EXlc_md_wint16),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_EXlc_md_wint17/FROM )
  );
  defparam DLX_EXlc_md_mda14_a1.INIT = 16'h5500;
  X_LUT4 DLX_EXlc_md_mda14_a1 (
    .ADR0(DLX_EXlc_pd_wint5),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_EXlc_md_wint13),
    .O(\DLX_EXlc_md_wint17/GROM )
  );
  X_BUF \DLX_EXlc_md_wint17/XUSED  (
    .I(\DLX_EXlc_md_wint17/FROM ),
    .O(DLX_EXlc_md_wint17)
  );
  X_BUF \DLX_EXlc_md_wint17/YUSED  (
    .I(\DLX_EXlc_md_wint17/GROM ),
    .O(DLX_EXlc_md_wint14)
  );
  defparam \DLX_IDinst__n0086<10>25 .INIT = 16'hCDCC;
  X_LUT4 \DLX_IDinst__n0086<10>25  (
    .ADR0(DLX_IDinst__n0364),
    .ADR1(CHOICE2672),
    .ADR2(DLX_IDinst_N70918),
    .ADR3(CHOICE2668),
    .O(\DLX_IDinst_branch_address<10>/FROM )
  );
  defparam \DLX_IDinst__n0086<10>31 .INIT = 16'hFFC0;
  X_LUT4 \DLX_IDinst__n0086<10>31  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst__n0128[10]),
    .ADR2(N100609),
    .ADR3(CHOICE2673),
    .O(N105724)
  );
  X_BUF \DLX_IDinst_branch_address<10>/XUSED  (
    .I(\DLX_IDinst_branch_address<10>/FROM ),
    .O(CHOICE2673)
  );
  defparam DLX_EXinst_Ker6582566.INIT = 16'hFFA8;
  X_LUT4 DLX_EXinst_Ker6582566 (
    .ADR0(N110065),
    .ADR1(CHOICE2064),
    .ADR2(CHOICE2060),
    .ADR3(CHOICE2069),
    .O(\N102270/FROM )
  );
  defparam \DLX_EXinst__n0006<30>115 .INIT = 16'hEFEE;
  X_LUT4 \DLX_EXinst__n0006<30>115  (
    .ADR0(CHOICE5256),
    .ADR1(CHOICE5278),
    .ADR2(DLX_IDinst_IR_function_field[4]),
    .ADR3(N102270),
    .O(\N102270/GROM )
  );
  X_BUF \N102270/XUSED  (
    .I(\N102270/FROM ),
    .O(N102270)
  );
  X_BUF \N102270/YUSED  (
    .I(\N102270/GROM ),
    .O(CHOICE5279)
  );
  defparam DLX_EXinst__n012743.INIT = 16'hFFF8;
  X_LUT4 DLX_EXinst__n012743 (
    .ADR0(CHOICE1972),
    .ADR1(DLX_IDinst_IR_function_field[4]),
    .ADR2(N126528),
    .ADR3(CHOICE1977),
    .O(\N101725/FROM )
  );
  defparam \DLX_EXinst__n0006<15>224 .INIT = 16'hFEEE;
  X_LUT4 \DLX_EXinst__n0006<15>224  (
    .ADR0(CHOICE4849),
    .ADR1(CHOICE4862),
    .ADR2(DLX_EXinst_ALU_result[15]),
    .ADR3(N101725),
    .O(\N101725/GROM )
  );
  X_BUF \N101725/XUSED  (
    .I(\N101725/FROM ),
    .O(N101725)
  );
  X_BUF \N101725/YUSED  (
    .I(\N101725/GROM ),
    .O(CHOICE4863)
  );
  defparam \DLX_EXinst__n0006<8>249 .INIT = 16'hCE00;
  X_LUT4 \DLX_EXinst__n0006<8>249  (
    .ADR0(CHOICE3700),
    .ADR1(CHOICE3729),
    .ADR2(DLX_EXinst__n0030_1),
    .ADR3(DLX_EXinst__n0149),
    .O(\DLX_EXinst_ALU_result<8>/FROM )
  );
  defparam \DLX_EXinst__n0006<8>259 .INIT = 16'hFFF0;
  X_LUT4 \DLX_EXinst__n0006<8>259  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N63689),
    .ADR3(CHOICE3731),
    .O(\DLX_EXinst_ALU_result<8>/GROM )
  );
  X_BUF \DLX_EXinst_ALU_result<8>/XUSED  (
    .I(\DLX_EXinst_ALU_result<8>/FROM ),
    .O(CHOICE3731)
  );
  X_BUF \DLX_EXinst_ALU_result<8>/YUSED  (
    .I(\DLX_EXinst_ALU_result<8>/GROM ),
    .O(N111878)
  );
  defparam \DLX_EXinst__n0006<8>185 .INIT = 16'hEAC0;
  X_LUT4 \DLX_EXinst__n0006<8>185  (
    .ADR0(DLX_EXinst_ALU_result[8]),
    .ADR1(DLX_IDinst_reg_out_B[4]),
    .ADR2(N98218),
    .ADR3(N101725),
    .O(\CHOICE3725/FROM )
  );
  defparam \DLX_EXinst__n0006<8>186 .INIT = 16'hFFAA;
  X_LUT4 \DLX_EXinst__n0006<8>186  (
    .ADR0(CHOICE3722),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(CHOICE3725),
    .O(\CHOICE3725/GROM )
  );
  X_BUF \CHOICE3725/XUSED  (
    .I(\CHOICE3725/FROM ),
    .O(CHOICE3725)
  );
  X_BUF \CHOICE3725/YUSED  (
    .I(\CHOICE3725/GROM ),
    .O(CHOICE3726)
  );
  defparam DLX_EXinst__n012728.INIT = 16'hF000;
  X_LUT4 DLX_EXinst__n012728 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_IR_function_field[2]),
    .ADR3(DLX_IDinst_IR_function_field[1]),
    .O(\CHOICE1976/FROM )
  );
  defparam DLX_EXinst__n012731.INIT = 16'hEA00;
  X_LUT4 DLX_EXinst__n012731 (
    .ADR0(DLX_IDinst_IR_function_field[3]),
    .ADR1(DLX_IDinst_IR_function_field[5]),
    .ADR2(DLX_IDinst_IR_function_field[0]),
    .ADR3(CHOICE1976),
    .O(\CHOICE1976/GROM )
  );
  X_BUF \CHOICE1976/XUSED  (
    .I(\CHOICE1976/FROM ),
    .O(CHOICE1976)
  );
  X_BUF \CHOICE1976/YUSED  (
    .I(\CHOICE1976/GROM ),
    .O(CHOICE1977)
  );
  defparam \DLX_EXinst__n0006<31>24 .INIT = 16'hEAC0;
  X_LUT4 \DLX_EXinst__n0006<31>24  (
    .ADR0(DLX_EXinst__n0016[31]),
    .ADR1(DLX_EXinst_ALU_result[31]),
    .ADR2(N101725),
    .ADR3(DLX_EXinst__n0114),
    .O(\CHOICE5746/FROM )
  );
  defparam \DLX_EXinst__n0006<0>4 .INIT = 16'hF888;
  X_LUT4 \DLX_EXinst__n0006<0>4  (
    .ADR0(N101725),
    .ADR1(DLX_EXinst_ALU_result[0]),
    .ADR2(DLX_EXinst__n0016[0]),
    .ADR3(DLX_EXinst__n0114),
    .O(\CHOICE5746/GROM )
  );
  X_BUF \CHOICE5746/XUSED  (
    .I(\CHOICE5746/FROM ),
    .O(CHOICE5746)
  );
  X_BUF \CHOICE5746/YUSED  (
    .I(\CHOICE5746/GROM ),
    .O(CHOICE5850)
  );
  defparam DLX_RF_delay_inst_wint161.INIT = 16'h3333;
  X_LUT4 DLX_RF_delay_inst_wint161 (
    .ADR0(VCC),
    .ADR1(DLX_RF_delay_inst_wint15),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_RF_delay_inst_wint16/GROM )
  );
  X_BUF \DLX_RF_delay_inst_wint16/YUSED  (
    .I(\DLX_RF_delay_inst_wint16/GROM ),
    .O(DLX_RF_delay_inst_wint16)
  );
  defparam DLX_RF_delay_inst_wint241.INIT = 16'h3333;
  X_LUT4 DLX_RF_delay_inst_wint241 (
    .ADR0(VCC),
    .ADR1(DLX_RF_delay_inst_wint23),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_RF_delay_inst_wint24/FROM )
  );
  defparam DLX_RF_delay_inst_wint251.INIT = 16'h00FF;
  X_LUT4 DLX_RF_delay_inst_wint251 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_RF_delay_inst_wint24),
    .O(\DLX_RF_delay_inst_wint24/GROM )
  );
  X_BUF \DLX_RF_delay_inst_wint24/XUSED  (
    .I(\DLX_RF_delay_inst_wint24/FROM ),
    .O(DLX_RF_delay_inst_wint24)
  );
  X_BUF \DLX_RF_delay_inst_wint24/YUSED  (
    .I(\DLX_RF_delay_inst_wint24/GROM ),
    .O(DLX_RF_delay_inst_wint25)
  );
  defparam DM_delay_inst_wint41.INIT = 16'h0F0F;
  X_LUT4 DM_delay_inst_wint41 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DM_delay_inst_wint3),
    .ADR3(VCC),
    .O(\DM_delay_inst_wint4/GROM )
  );
  X_BUF \DM_delay_inst_wint4/YUSED  (
    .I(\DM_delay_inst_wint4/GROM ),
    .O(DM_delay_inst_wint4)
  );
  defparam DLX_MEMlc_md_mda8_a1.INIT = 16'h00AA;
  X_LUT4 DLX_MEMlc_md_mda8_a1 (
    .ADR0(DLX_MEMlc_md_wint7),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_MEMlc_pd_wint1),
    .O(\DLX_MEMlc_md_wint8/FROM )
  );
  defparam DLX_MEMlc_md_mda9_a1.INIT = 16'h0F00;
  X_LUT4 DLX_MEMlc_md_mda9_a1 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_MEMlc_pd_wint1),
    .ADR3(DLX_MEMlc_md_wint8),
    .O(\DLX_MEMlc_md_wint8/GROM )
  );
  X_BUF \DLX_MEMlc_md_wint8/XUSED  (
    .I(\DLX_MEMlc_md_wint8/FROM ),
    .O(DLX_MEMlc_md_wint8)
  );
  X_BUF \DLX_MEMlc_md_wint8/YUSED  (
    .I(\DLX_MEMlc_md_wint8/GROM ),
    .O(DLX_MEMlc_md_wint9)
  );
  defparam DLX_RF_delay_inst_wint171.INIT = 16'h00FF;
  X_LUT4 DLX_RF_delay_inst_wint171 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_RF_delay_inst_wint16),
    .O(\DLX_RF_delay_inst_wint17/GROM )
  );
  X_BUF \DLX_RF_delay_inst_wint17/YUSED  (
    .I(\DLX_RF_delay_inst_wint17/GROM ),
    .O(DLX_RF_delay_inst_wint17)
  );
  defparam DM_delay_inst_wint51.INIT = 16'h00FF;
  X_LUT4 DM_delay_inst_wint51 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DM_delay_inst_wint4),
    .O(\DM_delay_inst_wint5/GROM )
  );
  X_BUF \DM_delay_inst_wint5/YUSED  (
    .I(\DM_delay_inst_wint5/GROM ),
    .O(DM_delay_inst_wint5)
  );
  defparam vga_top_vga1_Ker733921.INIT = 16'h0101;
  X_LUT4 vga_top_vga1_Ker733921 (
    .ADR0(vga_top_vga1_vcounter[7]),
    .ADR1(vga_top_vga1_vcounter[6]),
    .ADR2(vga_top_vga1_vcounter[8]),
    .ADR3(VCC),
    .O(\vga_top_vga1_N73394/GROM )
  );
  X_BUF \vga_top_vga1_N73394/YUSED  (
    .I(\vga_top_vga1_N73394/GROM ),
    .O(vga_top_vga1_N73394)
  );
  defparam DLX_RF_delay_inst_wint181.INIT = 16'h3333;
  X_LUT4 DLX_RF_delay_inst_wint181 (
    .ADR0(VCC),
    .ADR1(DLX_RF_delay_inst_wint17),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_RF_delay_inst_wint18/GROM )
  );
  X_BUF \DLX_RF_delay_inst_wint18/YUSED  (
    .I(\DLX_RF_delay_inst_wint18/GROM ),
    .O(DLX_RF_delay_inst_wint18)
  );
  defparam DLX_RF_delay_inst_wint261.INIT = 16'h0F0F;
  X_LUT4 DLX_RF_delay_inst_wint261 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_RF_delay_inst_wint25),
    .ADR3(VCC),
    .O(\DLX_RF_delay_inst_wint26/GROM )
  );
  X_BUF \DLX_RF_delay_inst_wint26/YUSED  (
    .I(\DLX_RF_delay_inst_wint26/GROM ),
    .O(DLX_RF_delay_inst_wint26)
  );
  defparam DM_delay_inst_wint61.INIT = 16'h0F0F;
  X_LUT4 DM_delay_inst_wint61 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DM_delay_inst_wint5),
    .ADR3(VCC),
    .O(\DM_delay_inst_wint6/GROM )
  );
  X_BUF \DM_delay_inst_wint6/YUSED  (
    .I(\DM_delay_inst_wint6/GROM ),
    .O(DM_delay_inst_wint6)
  );
  defparam DLX_IDinst_Ker700751.INIT = 16'hFFFA;
  X_LUT4 DLX_IDinst_Ker700751 (
    .ADR0(DLX_IDinst_slot_num_FFd3),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_slot_num_FFd1),
    .ADR3(DLX_IDinst_slot_num_FFd2),
    .O(\DLX_IDinst_N70077/FROM )
  );
  defparam \DLX_IDinst_slot_num_FFd3-In15_SW0 .INIT = 16'hFDFC;
  X_LUT4 \DLX_IDinst_slot_num_FFd3-In15_SW0  (
    .ADR0(DLX_IDinst_delay_slot),
    .ADR1(DLX_IDinst_slot_num_FFd3),
    .ADR2(DLX_IDinst_slot_num_FFd1),
    .ADR3(DLX_IDinst_slot_num_FFd2),
    .O(\DLX_IDinst_N70077/GROM )
  );
  X_BUF \DLX_IDinst_N70077/XUSED  (
    .I(\DLX_IDinst_N70077/FROM ),
    .O(DLX_IDinst_N70077)
  );
  X_BUF \DLX_IDinst_N70077/YUSED  (
    .I(\DLX_IDinst_N70077/GROM ),
    .O(N126589)
  );
  defparam DLX_RF_delay_inst_wint191.INIT = 16'h00FF;
  X_LUT4 DLX_RF_delay_inst_wint191 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_RF_delay_inst_wint18),
    .O(\DLX_RF_delay_inst_wint19/GROM )
  );
  X_BUF \DLX_RF_delay_inst_wint19/YUSED  (
    .I(\DLX_RF_delay_inst_wint19/GROM ),
    .O(DLX_RF_delay_inst_wint19)
  );
  defparam DLX_RF_delay_inst_wint271.INIT = 16'h0F0F;
  X_LUT4 DLX_RF_delay_inst_wint271 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_RF_delay_inst_wint26),
    .ADR3(VCC),
    .O(\DLX_RF_delay_inst_wint27/GROM )
  );
  X_BUF \DLX_RF_delay_inst_wint27/YUSED  (
    .I(\DLX_RF_delay_inst_wint27/GROM ),
    .O(DLX_RF_delay_inst_wint27)
  );
  defparam DM_delay_inst_wint71.INIT = 16'h0F0F;
  X_LUT4 DM_delay_inst_wint71 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DM_delay_inst_wint6),
    .ADR3(VCC),
    .O(\DM_delay_inst_wint7/GROM )
  );
  X_BUF \DM_delay_inst_wint7/YUSED  (
    .I(\DM_delay_inst_wint7/GROM ),
    .O(DM_delay_inst_wint7)
  );
  defparam \DLX_EXinst__n0006<1>7 .INIT = 16'h0040;
  X_LUT4 \DLX_EXinst__n0006<1>7  (
    .ADR0(DLX_IDinst_IR_function_field[2]),
    .ADR1(DLX_EXinst_N66525),
    .ADR2(\DLX_EXinst_Mshift__n0027_Sh[1] ),
    .ADR3(DLX_IDinst_IR_function_field[3]),
    .O(\CHOICE5657/FROM )
  );
  defparam \DLX_EXinst__n0006<1>16 .INIT = 16'h3320;
  X_LUT4 \DLX_EXinst__n0006<1>16  (
    .ADR0(DLX_EXinst_N66373),
    .ADR1(N109130),
    .ADR2(\DLX_EXinst_Mshift__n0028_Sh[49] ),
    .ADR3(CHOICE5657),
    .O(\CHOICE5657/GROM )
  );
  X_BUF \CHOICE5657/XUSED  (
    .I(\CHOICE5657/FROM ),
    .O(CHOICE5657)
  );
  X_BUF \CHOICE5657/YUSED  (
    .I(\CHOICE5657/GROM ),
    .O(CHOICE5659)
  );
  defparam \DLX_IDinst__n0113<1>_SW0 .INIT = 16'hE0EE;
  X_LUT4 \DLX_IDinst__n0113<1>_SW0  (
    .ADR0(CHOICE2100),
    .ADR1(DLX_IDinst_N69963),
    .ADR2(DLX_IDinst_IR_latched[30]),
    .ADR3(DLX_IDinst_N70991),
    .O(\DLX_IDinst_IR_opcode_field<1>/FROM )
  );
  defparam \DLX_IDinst__n0113<1> .INIT = 16'hA080;
  X_LUT4 \DLX_IDinst__n0113<1>  (
    .ADR0(DLX_IDinst_IR_latched[27]),
    .ADR1(DLX_IDinst__n0364),
    .ADR2(DLX_IDinst_N70679),
    .ADR3(N95527),
    .O(DLX_IDinst__n0113[1])
  );
  X_BUF \DLX_IDinst_IR_opcode_field<1>/XUSED  (
    .I(\DLX_IDinst_IR_opcode_field<1>/FROM ),
    .O(N95527)
  );
  defparam DLX_RF_delay_inst_wint281.INIT = 16'h3333;
  X_LUT4 DLX_RF_delay_inst_wint281 (
    .ADR0(VCC),
    .ADR1(DLX_RF_delay_inst_wint27),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_RF_delay_inst_wint28/GROM )
  );
  X_BUF \DLX_RF_delay_inst_wint28/YUSED  (
    .I(\DLX_RF_delay_inst_wint28/GROM ),
    .O(DLX_RF_delay_inst_wint28)
  );
  defparam DM_delay_inst_wint81.INIT = 16'h3333;
  X_LUT4 DM_delay_inst_wint81 (
    .ADR0(VCC),
    .ADR1(DM_delay_inst_wint7),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DM_delay_inst_wint8/GROM )
  );
  X_BUF \DM_delay_inst_wint8/YUSED  (
    .I(\DM_delay_inst_wint8/GROM ),
    .O(DM_delay_inst_wint8)
  );
  defparam DLX_IDlc_slave_ctrlID__n0001_SW110.INIT = 16'h88F8;
  X_LUT4 DLX_IDlc_slave_ctrlID__n0001_SW110 (
    .ADR0(DLX_reqout_ID),
    .ADR1(DLX_ackout_ID),
    .ADR2(DLX_IDlc_slave_ctrlID_l),
    .ADR3(reset_IBUF_3),
    .O(\CHOICE51/FROM )
  );
  defparam DLX_IDlc_slave_ctrlID__n0001_SW111.INIT = 16'hCC00;
  X_LUT4 DLX_IDlc_slave_ctrlID__n0001_SW111 (
    .ADR0(VCC),
    .ADR1(DLX_IDlc_master_ctrlID_nro),
    .ADR2(VCC),
    .ADR3(CHOICE51),
    .O(\CHOICE51/GROM )
  );
  X_BUF \CHOICE51/XUSED  (
    .I(\CHOICE51/FROM ),
    .O(CHOICE51)
  );
  X_BUF \CHOICE51/YUSED  (
    .I(\CHOICE51/GROM ),
    .O(DLX_IDlc_slave_ctrlID_l)
  );
  defparam DLX_RF_delay_inst_wint291.INIT = 16'h0F0F;
  X_LUT4 DLX_RF_delay_inst_wint291 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_RF_delay_inst_wint28),
    .ADR3(VCC),
    .O(\DLX_RF_delay_inst_wint29/GROM )
  );
  X_BUF \DLX_RF_delay_inst_wint29/YUSED  (
    .I(\DLX_RF_delay_inst_wint29/GROM ),
    .O(DLX_RF_delay_inst_wint29)
  );
  defparam DM_delay_inst_wint91.INIT = 16'h0F0F;
  X_LUT4 DM_delay_inst_wint91 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DM_delay_inst_wint8),
    .ADR3(VCC),
    .O(\DM_delay_inst_wint9/GROM )
  );
  X_BUF \DM_delay_inst_wint9/YUSED  (
    .I(\DM_delay_inst_wint9/GROM ),
    .O(DM_delay_inst_wint9)
  );
  defparam \DLX_EXinst__n0006<18>14 .INIT = 16'h0008;
  X_LUT4 \DLX_EXinst__n0006<18>14  (
    .ADR0(DLX_EXinst_N66087),
    .ADR1(\DLX_EXinst_Mshift__n0027_Sh[2] ),
    .ADR2(DLX_IDinst_IR_function_field[3]),
    .ADR3(DLX_IDinst_IR_function_field[2]),
    .O(\CHOICE5411/FROM )
  );
  defparam \DLX_EXinst__n0006<2>7 .INIT = 16'h0040;
  X_LUT4 \DLX_EXinst__n0006<2>7  (
    .ADR0(DLX_IDinst_IR_function_field[2]),
    .ADR1(DLX_EXinst_N66525),
    .ADR2(\DLX_EXinst_Mshift__n0027_Sh[2] ),
    .ADR3(DLX_IDinst_IR_function_field[3]),
    .O(\CHOICE5411/GROM )
  );
  X_BUF \CHOICE5411/XUSED  (
    .I(\CHOICE5411/FROM ),
    .O(CHOICE5411)
  );
  X_BUF \CHOICE5411/YUSED  (
    .I(\CHOICE5411/GROM ),
    .O(CHOICE5491)
  );
  defparam \DLX_IDinst__n0113<3>_SW0_SW0 .INIT = 16'h2F0F;
  X_LUT4 \DLX_IDinst__n0113<3>_SW0_SW0  (
    .ADR0(DLX_IDinst__n0350),
    .ADR1(DLX_IDinst__n0004),
    .ADR2(DLX_IDinst_N70610),
    .ADR3(DLX_IDinst__n0078),
    .O(\N127139/FROM )
  );
  defparam DLX_IDinst__n010959.INIT = 16'h50C0;
  X_LUT4 DLX_IDinst__n010959 (
    .ADR0(DLX_IDinst__n0350),
    .ADR1(CHOICE3519),
    .ADR2(DLX_IDinst__n0062),
    .ADR3(DLX_IDinst__n0348),
    .O(\N127139/GROM )
  );
  X_BUF \N127139/XUSED  (
    .I(\N127139/FROM ),
    .O(N127139)
  );
  X_BUF \N127139/YUSED  (
    .I(\N127139/GROM ),
    .O(CHOICE3523)
  );
  defparam DLX_IDinst__n010984.INIT = 16'hCC88;
  X_LUT4 DLX_IDinst__n010984 (
    .ADR0(CHOICE3523),
    .ADR1(DLX_IDinst_N70610),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_N70035),
    .O(\CHOICE3525/FROM )
  );
  defparam DLX_IDinst__n0109100.INIT = 16'hFFC8;
  X_LUT4 DLX_IDinst__n0109100 (
    .ADR0(DLX_IDinst__n0448[1]),
    .ADR1(DLX_IDinst_N69963),
    .ADR2(DLX_IDinst__n0062),
    .ADR3(CHOICE3525),
    .O(\CHOICE3525/GROM )
  );
  X_BUF \CHOICE3525/XUSED  (
    .I(\CHOICE3525/FROM ),
    .O(CHOICE3525)
  );
  X_BUF \CHOICE3525/YUSED  (
    .I(\CHOICE3525/GROM ),
    .O(CHOICE3526)
  );
  defparam vga_top_vga1_Ker733971.INIT = 16'h0001;
  X_LUT4 vga_top_vga1_Ker733971 (
    .ADR0(vga_top_vga1_hcounter[2]),
    .ADR1(vga_top_vga1_hcounter[3]),
    .ADR2(vga_top_vga1_hcounter[0]),
    .ADR3(vga_top_vga1_hcounter[8]),
    .O(\vga_top_vga1_N73399/FROM )
  );
  defparam vga_top_vga1__n000835.INIT = 16'hF000;
  X_LUT4 vga_top_vga1__n000835 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_N73379),
    .ADR3(vga_top_vga1_N73399),
    .O(\vga_top_vga1_N73399/GROM )
  );
  X_BUF \vga_top_vga1_N73399/XUSED  (
    .I(\vga_top_vga1_N73399/FROM ),
    .O(vga_top_vga1_N73399)
  );
  X_BUF \vga_top_vga1_N73399/YUSED  (
    .I(\vga_top_vga1_N73399/GROM ),
    .O(CHOICE3224)
  );
  defparam \DLX_EXinst__n0006<3>7 .INIT = 16'h0200;
  X_LUT4 \DLX_EXinst__n0006<3>7  (
    .ADR0(DLX_EXinst_N66525),
    .ADR1(DLX_IDinst_IR_function_field[3]),
    .ADR2(DLX_IDinst_IR_function_field[2]),
    .ADR3(\DLX_EXinst_Mshift__n0027_Sh[3] ),
    .O(\CHOICE5020/FROM )
  );
  defparam \DLX_EXinst__n0006<3>16 .INIT = 16'h3320;
  X_LUT4 \DLX_EXinst__n0006<3>16  (
    .ADR0(DLX_EXinst_N66373),
    .ADR1(N109130),
    .ADR2(\DLX_EXinst_Mshift__n0028_Sh[51] ),
    .ADR3(CHOICE5020),
    .O(\CHOICE5020/GROM )
  );
  X_BUF \CHOICE5020/XUSED  (
    .I(\CHOICE5020/FROM ),
    .O(CHOICE5020)
  );
  X_BUF \CHOICE5020/YUSED  (
    .I(\CHOICE5020/GROM ),
    .O(CHOICE5022)
  );
  defparam \DLX_EXinst__n0006<9>59_SW0 .INIT = 16'h1111;
  X_LUT4 \DLX_EXinst__n0006<9>59_SW0  (
    .ADR0(DLX_IDinst_IR_opcode_field[0]),
    .ADR1(DLX_IDinst_reg_out_A[9]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\N127378/FROM )
  );
  defparam \DLX_EXinst__n0006<21>85_SW0 .INIT = 16'h000F;
  X_LUT4 \DLX_EXinst__n0006<21>85_SW0  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_IR_opcode_field[0]),
    .ADR3(DLX_IDinst_reg_out_A[21]),
    .O(\N127378/GROM )
  );
  X_BUF \N127378/XUSED  (
    .I(\N127378/FROM ),
    .O(N127378)
  );
  X_BUF \N127378/YUSED  (
    .I(\N127378/GROM ),
    .O(N127370)
  );
  defparam DLX_IFlc_md_mda33_a1.INIT = 16'h2222;
  X_LUT4 DLX_IFlc_md_mda33_a1 (
    .ADR0(DLX_IFlc_md_wint32),
    .ADR1(DLX_IFlc_pd_wint1),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IFlc_md_wint33/FROM )
  );
  defparam DLX_IFlc_md_mda10_a1.INIT = 16'h00CC;
  X_LUT4 DLX_IFlc_md_mda10_a1 (
    .ADR0(VCC),
    .ADR1(DLX_IFlc_md_wint9),
    .ADR2(VCC),
    .ADR3(DLX_IFlc_pd_wint1),
    .O(\DLX_IFlc_md_wint33/GROM )
  );
  X_BUF \DLX_IFlc_md_wint33/XUSED  (
    .I(\DLX_IFlc_md_wint33/FROM ),
    .O(DLX_IFlc_md_wint33)
  );
  X_BUF \DLX_IFlc_md_wint33/YUSED  (
    .I(\DLX_IFlc_md_wint33/GROM ),
    .O(DLX_IFlc_md_wint10)
  );
  defparam DLX_IDinst__n03381.INIT = 16'h4500;
  X_LUT4 DLX_IDinst__n03381 (
    .ADR0(DLX_IDinst_IR_latched[28]),
    .ADR1(DLX_IDinst_IR_latched[26]),
    .ADR2(DLX_IDinst_IR_latched[27]),
    .ADR3(DLX_IDinst_IR_latched[29]),
    .O(\DLX_IDinst__n0338/FROM )
  );
  defparam DLX_IDinst__n034210.INIT = 16'h8A00;
  X_LUT4 DLX_IDinst__n034210 (
    .ADR0(DLX_IDinst_IR_latched[29]),
    .ADR1(DLX_IDinst_IR_latched[26]),
    .ADR2(DLX_IDinst_IR_latched[27]),
    .ADR3(DLX_IDinst_IR_latched[31]),
    .O(\DLX_IDinst__n0338/GROM )
  );
  X_BUF \DLX_IDinst__n0338/XUSED  (
    .I(\DLX_IDinst__n0338/FROM ),
    .O(DLX_IDinst__n0338)
  );
  X_BUF \DLX_IDinst__n0338/YUSED  (
    .I(\DLX_IDinst__n0338/GROM ),
    .O(CHOICE1796)
  );
  defparam DLX_IFlc_md_mda32_a1.INIT = 16'h5050;
  X_LUT4 DLX_IFlc_md_mda32_a1 (
    .ADR0(DLX_IFlc_pd_wint1),
    .ADR1(VCC),
    .ADR2(DLX_IFlc_md_wint31),
    .ADR3(VCC),
    .O(\DLX_IFlc_md_wint32/FROM )
  );
  defparam DLX_IFlc_md_mda11_a1.INIT = 16'h00CC;
  X_LUT4 DLX_IFlc_md_mda11_a1 (
    .ADR0(VCC),
    .ADR1(DLX_IFlc_md_wint10),
    .ADR2(VCC),
    .ADR3(DLX_IFlc_pd_wint1),
    .O(\DLX_IFlc_md_wint32/GROM )
  );
  X_BUF \DLX_IFlc_md_wint32/XUSED  (
    .I(\DLX_IFlc_md_wint32/FROM ),
    .O(DLX_IFlc_md_wint32)
  );
  X_BUF \DLX_IFlc_md_wint32/YUSED  (
    .I(\DLX_IFlc_md_wint32/GROM ),
    .O(DLX_IFlc_md_wint11)
  );
  defparam \DLX_EXinst__n0006<16>360_SW0 .INIT = 16'hFEFA;
  X_LUT4 \DLX_EXinst__n0006<16>360_SW0  (
    .ADR0(CHOICE5140),
    .ADR1(DLX_EXinst__n0016[16]),
    .ADR2(CHOICE5169),
    .ADR3(DLX_EXinst__n0114),
    .O(\N126847/FROM )
  );
  defparam \DLX_EXinst__n0006<16>360 .INIT = 16'hF808;
  X_LUT4 \DLX_EXinst__n0006<16>360  (
    .ADR0(DLX_EXinst__n0016[16]),
    .ADR1(DLX_EXinst__n0128),
    .ADR2(DLX_EXinst__n0030),
    .ADR3(N126847),
    .O(\N126847/GROM )
  );
  X_BUF \N126847/XUSED  (
    .I(\N126847/FROM ),
    .O(N126847)
  );
  X_BUF \N126847/YUSED  (
    .I(\N126847/GROM ),
    .O(CHOICE5172)
  );
  defparam DLX_IDinst__n0122115.INIT = 16'h0800;
  X_LUT4 DLX_IDinst__n0122115 (
    .ADR0(DLX_IDinst_IR_latched[26]),
    .ADR1(DLX_IDinst_N70909),
    .ADR2(DLX_IDinst_IR_latched[28]),
    .ADR3(DLX_IDinst_IR_latched[27]),
    .O(\CHOICE3317/FROM )
  );
  defparam DLX_IDinst__n034217.INIT = 16'h0030;
  X_LUT4 DLX_IDinst__n034217 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_IR_latched[27]),
    .ADR2(DLX_IDinst_N70909),
    .ADR3(DLX_IDinst_IR_latched[26]),
    .O(\CHOICE3317/GROM )
  );
  X_BUF \CHOICE3317/XUSED  (
    .I(\CHOICE3317/FROM ),
    .O(CHOICE3317)
  );
  X_BUF \CHOICE3317/YUSED  (
    .I(\CHOICE3317/GROM ),
    .O(CHOICE1800)
  );
  X_OR2 \DLX_IFinst_PC<9>/FFY/RSTOR  (
    .I0(reset_IBUF_1),
    .I1(GSR),
    .O(\DLX_IFinst_PC<9>/FFY/RST )
  );
  defparam DLX_IFinst_PC_8.INIT = 1'b0;
  X_FF DLX_IFinst_PC_8 (
    .I(DLX_IFinst_NPC[8]),
    .CE(DLX_IFinst_PC_N3535),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_PC<9>/FFY/RST ),
    .O(DLX_IFinst_PC[8])
  );
  defparam DLX_IFlc_md_mda29_a1.INIT = 16'h5500;
  X_LUT4 DLX_IFlc_md_mda29_a1 (
    .ADR0(DLX_IFlc_pd_wint1),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IFlc_md_wint28),
    .O(\DLX_IFlc_md_wint29/FROM )
  );
  defparam DLX_IFlc_md_mda20_a1.INIT = 16'h00AA;
  X_LUT4 DLX_IFlc_md_mda20_a1 (
    .ADR0(DLX_IFlc_md_wint19),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IFlc_pd_wint1),
    .O(\DLX_IFlc_md_wint29/GROM )
  );
  X_BUF \DLX_IFlc_md_wint29/XUSED  (
    .I(\DLX_IFlc_md_wint29/FROM ),
    .O(DLX_IFlc_md_wint29)
  );
  X_BUF \DLX_IFlc_md_wint29/YUSED  (
    .I(\DLX_IFlc_md_wint29/GROM ),
    .O(DLX_IFlc_md_wint20)
  );
  defparam DLX_IFlc_md_mda28_a1.INIT = 16'h4444;
  X_LUT4 DLX_IFlc_md_mda28_a1 (
    .ADR0(DLX_IFlc_pd_wint1),
    .ADR1(DLX_IFlc_md_wint27),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IFlc_md_wint28/FROM )
  );
  defparam DLX_IFlc_md_mda12_a1.INIT = 16'h0F00;
  X_LUT4 DLX_IFlc_md_mda12_a1 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IFlc_pd_wint1),
    .ADR3(DLX_IFlc_md_wint11),
    .O(\DLX_IFlc_md_wint28/GROM )
  );
  X_BUF \DLX_IFlc_md_wint28/XUSED  (
    .I(\DLX_IFlc_md_wint28/FROM ),
    .O(DLX_IFlc_md_wint28)
  );
  X_BUF \DLX_IFlc_md_wint28/YUSED  (
    .I(\DLX_IFlc_md_wint28/GROM ),
    .O(DLX_IFlc_md_wint12)
  );
  defparam DLX_IDinst_Ker6974431_SW0.INIT = 16'hF8F8;
  X_LUT4 DLX_IDinst_Ker6974431_SW0 (
    .ADR0(DLX_IDinst_N70924),
    .ADR1(DLX_IDinst_N70610),
    .ADR2(DLX_IDinst_N69963),
    .ADR3(VCC),
    .O(\N126580/FROM )
  );
  defparam DLX_IDinst__n008816.INIT = 16'hF800;
  X_LUT4 DLX_IDinst__n008816 (
    .ADR0(DLX_IDinst_N70924),
    .ADR1(DLX_IDinst_N70610),
    .ADR2(DLX_IDinst_N69963),
    .ADR3(DLX_IDinst_branch_sig),
    .O(\N126580/GROM )
  );
  X_BUF \N126580/XUSED  (
    .I(\N126580/FROM ),
    .O(N126580)
  );
  X_BUF \N126580/YUSED  (
    .I(\N126580/GROM ),
    .O(CHOICE3470)
  );
  defparam DLX_EXinst_Ker631271.INIT = 16'hFAFA;
  X_LUT4 DLX_EXinst_Ker631271 (
    .ADR0(DLX_IDinst_IR_function_field[0]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_IR_function_field[1]),
    .ADR3(VCC),
    .O(\DLX_EXinst_N63129/FROM )
  );
  defparam \DLX_EXinst__n0017<0>1 .INIT = 16'hB8B8;
  X_LUT4 \DLX_EXinst__n0017<0>1  (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(DLX_EXinst__n0030_1),
    .ADR2(DLX_IDinst_IR_function_field[0]),
    .ADR3(VCC),
    .O(\DLX_EXinst_N63129/GROM )
  );
  X_BUF \DLX_EXinst_N63129/XUSED  (
    .I(\DLX_EXinst_N63129/FROM ),
    .O(DLX_EXinst_N63129)
  );
  X_BUF \DLX_EXinst_N63129/YUSED  (
    .I(\DLX_EXinst_N63129/GROM ),
    .O(DLX_EXinst__n0017[0])
  );
  defparam DLX_IDinst__n008921.INIT = 16'hCCC8;
  X_LUT4 DLX_IDinst__n008921 (
    .ADR0(DLX_IDinst_IR_latched[30]),
    .ADR1(N126776),
    .ADR2(DLX_IDinst_IR_latched[31]),
    .ADR3(CHOICE2847),
    .O(\DLX_IDinst_Imm_31_1/FROM )
  );
  defparam DLX_IDinst__n008929.INIT = 16'h1000;
  X_LUT4 DLX_IDinst__n008929 (
    .ADR0(DLX_IDinst__n0331),
    .ADR1(DLX_IDinst_N70918),
    .ADR2(DLX_IDinst_jtarget[15]),
    .ADR3(CHOICE2849),
    .O(\DLX_IDinst_Imm_31_1/GROM )
  );
  X_BUF \DLX_IDinst_Imm_31_1/XUSED  (
    .I(\DLX_IDinst_Imm_31_1/FROM ),
    .O(CHOICE2849)
  );
  X_BUF \DLX_IDinst_Imm_31_1/YUSED  (
    .I(\DLX_IDinst_Imm_31_1/GROM ),
    .O(N106726)
  );
  defparam \DLX_EXinst_Mshift__n0027_Sh<47>_SW0 .INIT = 16'hF3C0;
  X_LUT4 \DLX_EXinst_Mshift__n0027_Sh<47>_SW0  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_IR_function_field_2_1),
    .ADR2(\DLX_EXinst_Mshift__n0027_Sh[11] ),
    .ADR3(\DLX_EXinst_Mshift__n0027_Sh[15] ),
    .O(\N93383/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0027_Sh<47> .INIT = 16'hAFA0;
  X_LUT4 \DLX_EXinst_Mshift__n0027_Sh<47>  (
    .ADR0(DLX_EXinst_N62831),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_IR_function_field_3_1),
    .ADR3(N93383),
    .O(\N93383/GROM )
  );
  X_BUF \N93383/XUSED  (
    .I(\N93383/FROM ),
    .O(N93383)
  );
  X_BUF \N93383/YUSED  (
    .I(\N93383/GROM ),
    .O(\DLX_EXinst_Mshift__n0027_Sh[47] )
  );
  defparam DLX_IDinst__n02501.INIT = 16'h0020;
  X_LUT4 DLX_IDinst__n02501 (
    .ADR0(DLX_IDinst_IR_latched[27]),
    .ADR1(DLX_IDinst_IR_latched[26]),
    .ADR2(DLX_IDinst_IR_latched[30]),
    .ADR3(DLX_IDinst_IR_latched[28]),
    .O(\DLX_IDinst__n0250/FROM )
  );
  defparam DLX_IDinst__n008850.INIT = 16'h9A9A;
  X_LUT4 DLX_IDinst__n008850 (
    .ADR0(DLX_IDinst_IR_latched[27]),
    .ADR1(DLX_IDinst_IR_latched[26]),
    .ADR2(DLX_IDinst_IR_latched[30]),
    .ADR3(VCC),
    .O(\DLX_IDinst__n0250/GROM )
  );
  X_BUF \DLX_IDinst__n0250/XUSED  (
    .I(\DLX_IDinst__n0250/FROM ),
    .O(DLX_IDinst__n0250)
  );
  X_BUF \DLX_IDinst__n0250/YUSED  (
    .I(\DLX_IDinst__n0250/GROM ),
    .O(CHOICE3480)
  );
  defparam DLX_EXinst_Ker634821.INIT = 16'hCFC0;
  X_LUT4 DLX_EXinst_Ker634821 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[6]),
    .ADR2(DLX_IDinst_IR_function_field[1]),
    .ADR3(DLX_IDinst_reg_out_A[8]),
    .O(\DLX_EXinst_N63484/FROM )
  );
  defparam \DLX_EXinst__n0017<1>1 .INIT = 16'hE2E2;
  X_LUT4 \DLX_EXinst__n0017<1>1  (
    .ADR0(DLX_IDinst_IR_function_field[1]),
    .ADR1(DLX_EXinst__n0030_1),
    .ADR2(DLX_IDinst_reg_out_B[1]),
    .ADR3(VCC),
    .O(\DLX_EXinst_N63484/GROM )
  );
  X_BUF \DLX_EXinst_N63484/XUSED  (
    .I(\DLX_EXinst_N63484/FROM ),
    .O(DLX_EXinst_N63484)
  );
  X_BUF \DLX_EXinst_N63484/YUSED  (
    .I(\DLX_EXinst_N63484/GROM ),
    .O(DLX_EXinst__n0017[1])
  );
  defparam DLX_IDinst__n008854.INIT = 16'h00A0;
  X_LUT4 DLX_IDinst__n008854 (
    .ADR0(DLX_IDinst_N70909),
    .ADR1(VCC),
    .ADR2(CHOICE3480),
    .ADR3(DLX_IDinst_IR_latched[28]),
    .O(\DLX_IDinst_branch_sig/FROM )
  );
  defparam DLX_IDinst__n008887.INIT = 16'h0F0E;
  X_LUT4 DLX_IDinst__n008887 (
    .ADR0(CHOICE3472),
    .ADR1(DLX_IDinst__n0364),
    .ADR2(DLX_IDinst__n0331),
    .ADR3(CHOICE3481),
    .O(\DLX_IDinst_branch_sig/GROM )
  );
  X_BUF \DLX_IDinst_branch_sig/XUSED  (
    .I(\DLX_IDinst_branch_sig/FROM ),
    .O(CHOICE3481)
  );
  X_BUF \DLX_IDinst_branch_sig/YUSED  (
    .I(\DLX_IDinst_branch_sig/GROM ),
    .O(N110516)
  );
  defparam DLX_IFlc_md_mda25_a1.INIT = 16'h2222;
  X_LUT4 DLX_IFlc_md_mda25_a1 (
    .ADR0(DLX_IFlc_md_wint24),
    .ADR1(DLX_IFlc_pd_wint1),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IFlc_md_wint25/FROM )
  );
  defparam DLX_IFlc_md_mda21_a1.INIT = 16'h3030;
  X_LUT4 DLX_IFlc_md_mda21_a1 (
    .ADR0(VCC),
    .ADR1(DLX_IFlc_pd_wint1),
    .ADR2(DLX_IFlc_md_wint20),
    .ADR3(VCC),
    .O(\DLX_IFlc_md_wint25/GROM )
  );
  X_BUF \DLX_IFlc_md_wint25/XUSED  (
    .I(\DLX_IFlc_md_wint25/FROM ),
    .O(DLX_IFlc_md_wint25)
  );
  X_BUF \DLX_IFlc_md_wint25/YUSED  (
    .I(\DLX_IFlc_md_wint25/GROM ),
    .O(DLX_IFlc_md_wint21)
  );
  defparam DLX_IFlc_md_mda24_a1.INIT = 16'h0C0C;
  X_LUT4 DLX_IFlc_md_mda24_a1 (
    .ADR0(VCC),
    .ADR1(DLX_IFlc_md_wint23),
    .ADR2(DLX_IFlc_pd_wint1),
    .ADR3(VCC),
    .O(\DLX_IFlc_md_wint24/FROM )
  );
  defparam DLX_IFlc_md_mda13_a1.INIT = 16'h0A0A;
  X_LUT4 DLX_IFlc_md_mda13_a1 (
    .ADR0(DLX_IFlc_md_wint12),
    .ADR1(VCC),
    .ADR2(DLX_IFlc_pd_wint1),
    .ADR3(VCC),
    .O(\DLX_IFlc_md_wint24/GROM )
  );
  X_BUF \DLX_IFlc_md_wint24/XUSED  (
    .I(\DLX_IFlc_md_wint24/FROM ),
    .O(DLX_IFlc_md_wint24)
  );
  X_BUF \DLX_IFlc_md_wint24/YUSED  (
    .I(\DLX_IFlc_md_wint24/GROM ),
    .O(DLX_IFlc_md_wint13)
  );
  defparam \DLX_EXinst__n0017<9>1 .INIT = 16'hF0AA;
  X_LUT4 \DLX_EXinst__n0017<9>1  (
    .ADR0(\DLX_IDinst_Imm[9] ),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[9]),
    .ADR3(DLX_EXinst__n0030_1),
    .O(\DLX_EXinst__n0017<9>/FROM )
  );
  defparam \DLX_EXinst__n0017<2>1 .INIT = 16'hAACC;
  X_LUT4 \DLX_EXinst__n0017<2>1  (
    .ADR0(DLX_IDinst_reg_out_B[2]),
    .ADR1(DLX_IDinst_IR_function_field[2]),
    .ADR2(VCC),
    .ADR3(DLX_EXinst__n0030_1),
    .O(\DLX_EXinst__n0017<9>/GROM )
  );
  X_BUF \DLX_EXinst__n0017<9>/XUSED  (
    .I(\DLX_EXinst__n0017<9>/FROM ),
    .O(DLX_EXinst__n0017[9])
  );
  X_BUF \DLX_EXinst__n0017<9>/YUSED  (
    .I(\DLX_EXinst__n0017<9>/GROM ),
    .O(DLX_EXinst__n0017[2])
  );
  defparam \mask<1>_SW117 .INIT = 16'h585D;
  X_LUT4 \mask<1>_SW117  (
    .ADR0(DLX_EXinst_byte),
    .ADR1(DLX_EXinst_ALU_result[1]),
    .ADR2(DLX_EXinst_ALU_result[0]),
    .ADR3(DLX_EXinst_word),
    .O(\CHOICE292/FROM )
  );
  defparam \mask<1>_SW122 .INIT = 16'hAA00;
  X_LUT4 \mask<1>_SW122  (
    .ADR0(vga_select_6[0]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(CHOICE292),
    .O(\CHOICE292/GROM )
  );
  X_BUF \CHOICE292/XUSED  (
    .I(\CHOICE292/FROM ),
    .O(CHOICE292)
  );
  X_BUF \CHOICE292/YUSED  (
    .I(\CHOICE292/GROM ),
    .O(mask_1_OBUF)
  );
  defparam DLX_EXinst_Ker628041.INIT = 16'hAFA0;
  X_LUT4 DLX_EXinst_Ker628041 (
    .ADR0(DLX_IDinst_reg_out_A[21]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_IR_function_field[1]),
    .ADR3(DLX_IDinst_reg_out_A[23]),
    .O(\DLX_EXinst_N62806/FROM )
  );
  defparam DLX_EXinst_Ker630041.INIT = 16'hAFA0;
  X_LUT4 DLX_EXinst_Ker630041 (
    .ADR0(DLX_IDinst_reg_out_A[21]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_IR_function_field[1]),
    .ADR3(DLX_IDinst_reg_out_A[19]),
    .O(\DLX_EXinst_N62806/GROM )
  );
  X_BUF \DLX_EXinst_N62806/XUSED  (
    .I(\DLX_EXinst_N62806/FROM ),
    .O(DLX_EXinst_N62806)
  );
  X_BUF \DLX_EXinst_N62806/YUSED  (
    .I(\DLX_EXinst_N62806/GROM ),
    .O(DLX_EXinst_N63006)
  );
  defparam \DLX_EXinst__n0006<6>194 .INIT = 16'h5000;
  X_LUT4 \DLX_EXinst__n0006<6>194  (
    .ADR0(DLX_IDinst_reg_out_B[3]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N66226),
    .ADR3(DLX_EXinst_N62911),
    .O(\CHOICE4396/FROM )
  );
  defparam \DLX_EXinst__n0017<3>1 .INIT = 16'hFA0A;
  X_LUT4 \DLX_EXinst__n0017<3>1  (
    .ADR0(DLX_IDinst_IR_function_field[3]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst__n0030_1),
    .ADR3(DLX_IDinst_reg_out_B[3]),
    .O(\CHOICE4396/GROM )
  );
  X_BUF \CHOICE4396/XUSED  (
    .I(\CHOICE4396/FROM ),
    .O(CHOICE4396)
  );
  X_BUF \CHOICE4396/YUSED  (
    .I(\CHOICE4396/GROM ),
    .O(DLX_EXinst__n0017[3])
  );
  defparam DLX_IFlc_md_mda30_a1.INIT = 16'h5050;
  X_LUT4 DLX_IFlc_md_mda30_a1 (
    .ADR0(DLX_IFlc_pd_wint1),
    .ADR1(VCC),
    .ADR2(DLX_IFlc_md_wint29),
    .ADR3(VCC),
    .O(\DLX_IFlc_md_wint30/FROM )
  );
  defparam DLX_IFlc_md_mda31_a1.INIT = 16'h3300;
  X_LUT4 DLX_IFlc_md_mda31_a1 (
    .ADR0(VCC),
    .ADR1(DLX_IFlc_pd_wint1),
    .ADR2(VCC),
    .ADR3(DLX_IFlc_md_wint30),
    .O(\DLX_IFlc_md_wint30/GROM )
  );
  X_BUF \DLX_IFlc_md_wint30/XUSED  (
    .I(\DLX_IFlc_md_wint30/FROM ),
    .O(DLX_IFlc_md_wint30)
  );
  X_BUF \DLX_IFlc_md_wint30/YUSED  (
    .I(\DLX_IFlc_md_wint30/GROM ),
    .O(DLX_IFlc_md_wint31)
  );
  defparam DLX_IFlc_md_mda19_a1.INIT = 16'h4444;
  X_LUT4 DLX_IFlc_md_mda19_a1 (
    .ADR0(DLX_IFlc_pd_wint1),
    .ADR1(DLX_IFlc_md_wint18),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IFlc_md_wint19/FROM )
  );
  defparam DLX_IFlc_md_mda22_a1.INIT = 16'h5500;
  X_LUT4 DLX_IFlc_md_mda22_a1 (
    .ADR0(DLX_IFlc_pd_wint1),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IFlc_md_wint21),
    .O(\DLX_IFlc_md_wint19/GROM )
  );
  X_BUF \DLX_IFlc_md_wint19/XUSED  (
    .I(\DLX_IFlc_md_wint19/FROM ),
    .O(DLX_IFlc_md_wint19)
  );
  X_BUF \DLX_IFlc_md_wint19/YUSED  (
    .I(\DLX_IFlc_md_wint19/GROM ),
    .O(DLX_IFlc_md_wint22)
  );
  defparam DLX_IFlc_md_mda23_a1.INIT = 16'h00F0;
  X_LUT4 DLX_IFlc_md_mda23_a1 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IFlc_md_wint22),
    .ADR3(DLX_IFlc_pd_wint1),
    .O(\DLX_IFlc_md_wint23/FROM )
  );
  defparam DLX_IFlc_md_mda14_a1.INIT = 16'h3300;
  X_LUT4 DLX_IFlc_md_mda14_a1 (
    .ADR0(VCC),
    .ADR1(DLX_IFlc_pd_wint1),
    .ADR2(VCC),
    .ADR3(DLX_IFlc_md_wint13),
    .O(\DLX_IFlc_md_wint23/GROM )
  );
  X_BUF \DLX_IFlc_md_wint23/XUSED  (
    .I(\DLX_IFlc_md_wint23/FROM ),
    .O(DLX_IFlc_md_wint23)
  );
  X_BUF \DLX_IFlc_md_wint23/YUSED  (
    .I(\DLX_IFlc_md_wint23/GROM ),
    .O(DLX_IFlc_md_wint14)
  );
  defparam DLX_EXinst_Ker628091.INIT = 16'hBB88;
  X_LUT4 DLX_EXinst_Ker628091 (
    .ADR0(DLX_IDinst_reg_out_A[23]),
    .ADR1(DLX_IDinst_IR_function_field[1]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[25]),
    .O(\DLX_EXinst_N62811/FROM )
  );
  defparam DLX_EXinst_Ker630141.INIT = 16'hFC0C;
  X_LUT4 DLX_EXinst_Ker630141 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[23]),
    .ADR2(DLX_IDinst_IR_function_field[1]),
    .ADR3(DLX_IDinst_reg_out_A[25]),
    .O(\DLX_EXinst_N62811/GROM )
  );
  X_BUF \DLX_EXinst_N62811/XUSED  (
    .I(\DLX_EXinst_N62811/FROM ),
    .O(DLX_EXinst_N62811)
  );
  X_BUF \DLX_EXinst_N62811/YUSED  (
    .I(\DLX_EXinst_N62811/GROM ),
    .O(DLX_EXinst_N63016)
  );
  defparam DLX_EXinst_Ker664831.INIT = 16'h5500;
  X_LUT4 DLX_EXinst_Ker664831 (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N62631),
    .O(\DLX_EXinst_N66485/FROM )
  );
  defparam \DLX_EXinst__n0017<4>1 .INIT = 16'hB8B8;
  X_LUT4 \DLX_EXinst__n0017<4>1  (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(DLX_EXinst__n0030_1),
    .ADR2(DLX_IDinst_IR_function_field[4]),
    .ADR3(VCC),
    .O(\DLX_EXinst_N66485/GROM )
  );
  X_BUF \DLX_EXinst_N66485/XUSED  (
    .I(\DLX_EXinst_N66485/FROM ),
    .O(DLX_EXinst_N66485)
  );
  X_BUF \DLX_EXinst_N66485/YUSED  (
    .I(\DLX_EXinst_N66485/GROM ),
    .O(DLX_EXinst__n0017[4])
  );
  defparam DLX_EXinst_Ker630241.INIT = 16'hE2E2;
  X_LUT4 DLX_EXinst_Ker630241 (
    .ADR0(\DLX_EXinst_Mshift__n0028_Sh[22] ),
    .ADR1(DLX_IDinst_IR_function_field[3]),
    .ADR2(\DLX_EXinst_Mshift__n0028_Sh[30] ),
    .ADR3(VCC),
    .O(\DLX_EXinst_N63026/FROM )
  );
  defparam DLX_EXinst_Ker6515396.INIT = 16'h3B08;
  X_LUT4 DLX_EXinst_Ker6515396 (
    .ADR0(\DLX_EXinst_Mshift__n0024_Sh[26] ),
    .ADR1(DLX_IDinst_IR_function_field_2_1),
    .ADR2(DLX_IDinst_IR_function_field_3_1),
    .ADR3(DLX_EXinst_N63026),
    .O(\DLX_EXinst_N63026/GROM )
  );
  X_BUF \DLX_EXinst_N63026/XUSED  (
    .I(\DLX_EXinst_N63026/FROM ),
    .O(DLX_EXinst_N63026)
  );
  X_BUF \DLX_EXinst_N63026/YUSED  (
    .I(\DLX_EXinst_N63026/GROM ),
    .O(CHOICE3077)
  );
  defparam DLX_EXinst_Ker6615530.INIT = 16'h0F00;
  X_LUT4 DLX_EXinst_Ker6615530 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(\DLX_IDinst_Imm[5] ),
    .ADR3(\DLX_EXinst_Mshift__n0028_Sh[52] ),
    .O(\CHOICE1324/FROM )
  );
  defparam \DLX_EXinst__n0017<5>1 .INIT = 16'hF3C0;
  X_LUT4 \DLX_EXinst__n0017<5>1  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst__n0030_1),
    .ADR2(DLX_IDinst_reg_out_B[5]),
    .ADR3(\DLX_IDinst_Imm[5] ),
    .O(\CHOICE1324/GROM )
  );
  X_BUF \CHOICE1324/XUSED  (
    .I(\CHOICE1324/FROM ),
    .O(CHOICE1324)
  );
  X_BUF \CHOICE1324/YUSED  (
    .I(\CHOICE1324/GROM ),
    .O(DLX_EXinst__n0017[5])
  );
  defparam DLX_EXinst_Ker630091.INIT = 16'hACAC;
  X_LUT4 DLX_EXinst_Ker630091 (
    .ADR0(DLX_IDinst_reg_out_A[23]),
    .ADR1(DLX_IDinst_reg_out_A[21]),
    .ADR2(DLX_IDinst_IR_function_field[1]),
    .ADR3(VCC),
    .O(\DLX_EXinst_N63011/FROM )
  );
  defparam DLX_EXinst_Ker62713_SW0.INIT = 16'hEE22;
  X_LUT4 DLX_EXinst_Ker62713_SW0 (
    .ADR0(DLX_EXinst_N63514),
    .ADR1(DLX_IDinst_IR_function_field[0]),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N63011),
    .O(\DLX_EXinst_N63011/GROM )
  );
  X_BUF \DLX_EXinst_N63011/XUSED  (
    .I(\DLX_EXinst_N63011/FROM ),
    .O(DLX_EXinst_N63011)
  );
  X_BUF \DLX_EXinst_N63011/YUSED  (
    .I(\DLX_EXinst_N63011/GROM ),
    .O(N94007)
  );
  defparam DLX_EXinst__n003675_SW0.INIT = 16'hFFEE;
  X_LUT4 DLX_EXinst__n003675_SW0 (
    .ADR0(\DLX_IDinst_Imm[31] ),
    .ADR1(CHOICE3249),
    .ADR2(VCC),
    .ADR3(CHOICE3246),
    .O(\N125959/FROM )
  );
  defparam DLX_EXinst__n003675.INIT = 16'hFFFE;
  X_LUT4 DLX_EXinst__n003675 (
    .ADR0(\DLX_IDinst_Imm[6] ),
    .ADR1(\DLX_IDinst_Imm[5] ),
    .ADR2(\DLX_IDinst_Imm[7] ),
    .ADR3(N125959),
    .O(\N125959/GROM )
  );
  X_BUF \N125959/XUSED  (
    .I(\N125959/FROM ),
    .O(N125959)
  );
  X_BUF \N125959/YUSED  (
    .I(\N125959/GROM ),
    .O(N109130)
  );
  defparam DLX_IDinst_PIPEEMPTY1.INIT = 16'hC000;
  X_LUT4 DLX_IDinst_PIPEEMPTY1 (
    .ADR0(VCC),
    .ADR1(DLX_MEMinst_noop),
    .ADR2(FREEZE_IBUF),
    .ADR3(DLX_EXinst_noop),
    .O(\PIPEEMPTY_OBUF/GROM )
  );
  X_BUF \PIPEEMPTY_OBUF/YUSED  (
    .I(\PIPEEMPTY_OBUF/GROM ),
    .O(PIPEEMPTY_OBUF)
  );
  defparam DLX_IFlc_md_mda18_a1.INIT = 16'h4444;
  X_LUT4 DLX_IFlc_md_mda18_a1 (
    .ADR0(DLX_IFlc_pd_wint1),
    .ADR1(DLX_IFlc_md_wint17),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IFlc_md_wint18/FROM )
  );
  defparam DLX_IFlc_md_mda15_a1.INIT = 16'h4444;
  X_LUT4 DLX_IFlc_md_mda15_a1 (
    .ADR0(DLX_IFlc_pd_wint1),
    .ADR1(DLX_IFlc_md_wint14),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IFlc_md_wint18/GROM )
  );
  X_BUF \DLX_IFlc_md_wint18/XUSED  (
    .I(\DLX_IFlc_md_wint18/FROM ),
    .O(DLX_IFlc_md_wint18)
  );
  X_BUF \DLX_IFlc_md_wint18/YUSED  (
    .I(\DLX_IFlc_md_wint18/GROM ),
    .O(DLX_IFlc_md_wint15)
  );
  defparam \DLX_EXinst_Mshift__n0024_Sh<25> .INIT = 16'hAFA0;
  X_LUT4 \DLX_EXinst_Mshift__n0024_Sh<25>  (
    .ADR0(N94205),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_IR_function_field_0_1),
    .ADR3(DLX_EXinst_N63790),
    .O(\DLX_EXinst_Mshift__n0024_Sh<25>/FROM )
  );
  defparam DLX_EXinst_Ker648521.INIT = 16'hFC0C;
  X_LUT4 DLX_EXinst_Ker648521 (
    .ADR0(VCC),
    .ADR1(\DLX_EXinst_Mshift__n0028_Sh[17] ),
    .ADR2(DLX_IDinst_IR_function_field_3_1),
    .ADR3(\DLX_EXinst_Mshift__n0024_Sh[25] ),
    .O(\DLX_EXinst_Mshift__n0024_Sh<25>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0024_Sh<25>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0024_Sh<25>/FROM ),
    .O(\DLX_EXinst_Mshift__n0024_Sh[25] )
  );
  X_BUF \DLX_EXinst_Mshift__n0024_Sh<25>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0024_Sh<25>/GROM ),
    .O(DLX_EXinst_N64854)
  );
  defparam \DLX_EXinst__n0006<24>290_SW0 .INIT = 16'h5554;
  X_LUT4 \DLX_EXinst__n0006<24>290_SW0  (
    .ADR0(DLX_EXinst__n0030),
    .ADR1(CHOICE3759),
    .ADR2(CHOICE3736),
    .ADR3(CHOICE3745),
    .O(\DLX_EXinst_ALU_result<24>/FROM )
  );
  defparam \DLX_EXinst__n0006<24>290 .INIT = 16'hCCC8;
  X_LUT4 \DLX_EXinst__n0006<24>290  (
    .ADR0(CHOICE3791),
    .ADR1(DLX_EXinst__n0149),
    .ADR2(N100490),
    .ADR3(N126534),
    .O(N112254)
  );
  X_BUF \DLX_EXinst_ALU_result<24>/XUSED  (
    .I(\DLX_EXinst_ALU_result<24>/FROM ),
    .O(N126534)
  );
  defparam DLX_EXinst_Ker630341.INIT = 16'hFC30;
  X_LUT4 DLX_EXinst_Ker630341 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(DLX_IDinst_reg_out_A[11]),
    .ADR3(DLX_IDinst_reg_out_A[13]),
    .O(\DLX_EXinst_N63036/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0026_Sh<10>1 .INIT = 16'hFC0C;
  X_LUT4 \DLX_EXinst_Mshift__n0026_Sh<10>1  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N63329),
    .ADR2(DLX_IDinst_reg_out_B[0]),
    .ADR3(DLX_EXinst_N63036),
    .O(\DLX_EXinst_N63036/GROM )
  );
  X_BUF \DLX_EXinst_N63036/XUSED  (
    .I(\DLX_EXinst_N63036/FROM ),
    .O(DLX_EXinst_N63036)
  );
  X_BUF \DLX_EXinst_N63036/YUSED  (
    .I(\DLX_EXinst_N63036/GROM ),
    .O(\DLX_EXinst_Mshift__n0026_Sh[10] )
  );
  defparam \DLX_EXinst__n0017<10>1 .INIT = 16'hE4E4;
  X_LUT4 \DLX_EXinst__n0017<10>1  (
    .ADR0(DLX_EXinst__n0030_1),
    .ADR1(\DLX_IDinst_Imm[10] ),
    .ADR2(DLX_IDinst_reg_out_B[10]),
    .ADR3(VCC),
    .O(\DLX_EXinst__n0017<10>/FROM )
  );
  defparam \DLX_EXinst__n0017<6>1 .INIT = 16'hBB88;
  X_LUT4 \DLX_EXinst__n0017<6>1  (
    .ADR0(DLX_IDinst_reg_out_B[6]),
    .ADR1(DLX_EXinst__n0030_1),
    .ADR2(VCC),
    .ADR3(\DLX_IDinst_Imm[6] ),
    .O(\DLX_EXinst__n0017<10>/GROM )
  );
  X_BUF \DLX_EXinst__n0017<10>/XUSED  (
    .I(\DLX_EXinst__n0017<10>/FROM ),
    .O(DLX_EXinst__n0017[10])
  );
  X_BUF \DLX_EXinst__n0017<10>/YUSED  (
    .I(\DLX_EXinst__n0017<10>/GROM ),
    .O(DLX_EXinst__n0017[6])
  );
  defparam \DLX_IDinst__n0113<3>_SW0 .INIT = 16'h2300;
  X_LUT4 \DLX_IDinst__n0113<3>_SW0  (
    .ADR0(DLX_IDinst_N69963),
    .ADR1(DLX_IDinst__n0364),
    .ADR2(N127139),
    .ADR3(DLX_IDinst_N69568),
    .O(\DLX_IDinst_IR_opcode_field<3>/FROM )
  );
  defparam \DLX_IDinst__n0113<3> .INIT = 16'hA080;
  X_LUT4 \DLX_IDinst__n0113<3>  (
    .ADR0(DLX_IDinst_N70679),
    .ADR1(DLX_IDinst__n0364),
    .ADR2(DLX_IDinst_IR_latched[29]),
    .ADR3(N91278),
    .O(DLX_IDinst__n0113[3])
  );
  X_BUF \DLX_IDinst_IR_opcode_field<3>/XUSED  (
    .I(\DLX_IDinst_IR_opcode_field<3>/FROM ),
    .O(N91278)
  );
  defparam \DLX_EXinst_Mshift__n0024_Sh<27> .INIT = 16'hF3C0;
  X_LUT4 \DLX_EXinst_Mshift__n0024_Sh<27>  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_IR_function_field_1_1),
    .ADR2(DLX_EXinst_N62709),
    .ADR3(N93799),
    .O(\DLX_EXinst_Mshift__n0024_Sh<27>/FROM )
  );
  defparam DLX_EXinst_Ker648471.INIT = 16'hFC0C;
  X_LUT4 DLX_EXinst_Ker648471 (
    .ADR0(VCC),
    .ADR1(\DLX_EXinst_Mshift__n0028_Sh[19] ),
    .ADR2(DLX_IDinst_IR_function_field_3_1),
    .ADR3(\DLX_EXinst_Mshift__n0024_Sh[27] ),
    .O(\DLX_EXinst_Mshift__n0024_Sh<27>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0024_Sh<27>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0024_Sh<27>/FROM ),
    .O(\DLX_EXinst_Mshift__n0024_Sh[27] )
  );
  X_BUF \DLX_EXinst_Mshift__n0024_Sh<27>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0024_Sh<27>/GROM ),
    .O(DLX_EXinst_N64849)
  );
  defparam DLX_EXinst_Ker630441.INIT = 16'hCFC0;
  X_LUT4 DLX_EXinst_Ker630441 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[17]),
    .ADR2(DLX_IDinst_reg_out_B[1]),
    .ADR3(DLX_IDinst_reg_out_A[15]),
    .O(\DLX_EXinst_N63046/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0026_Sh<14>1 .INIT = 16'hEE22;
  X_LUT4 \DLX_EXinst_Mshift__n0026_Sh<14>1  (
    .ADR0(DLX_EXinst_N63414),
    .ADR1(DLX_IDinst_reg_out_B[0]),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N63046),
    .O(\DLX_EXinst_N63046/GROM )
  );
  X_BUF \DLX_EXinst_N63046/XUSED  (
    .I(\DLX_EXinst_N63046/FROM ),
    .O(DLX_EXinst_N63046)
  );
  X_BUF \DLX_EXinst_N63046/YUSED  (
    .I(\DLX_EXinst_N63046/GROM ),
    .O(\DLX_EXinst_Mshift__n0026_Sh[14] )
  );
  defparam \DLX_EXinst__n0017<13>1 .INIT = 16'hF5A0;
  X_LUT4 \DLX_EXinst__n0017<13>1  (
    .ADR0(DLX_EXinst__n0030_1),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[13]),
    .ADR3(\DLX_IDinst_Imm[13] ),
    .O(\DLX_EXinst__n0017<13>/FROM )
  );
  defparam \DLX_EXinst__n0017<7>1 .INIT = 16'hAACC;
  X_LUT4 \DLX_EXinst__n0017<7>1  (
    .ADR0(DLX_IDinst_reg_out_B[7]),
    .ADR1(\DLX_IDinst_Imm[7] ),
    .ADR2(VCC),
    .ADR3(DLX_EXinst__n0030_1),
    .O(\DLX_EXinst__n0017<13>/GROM )
  );
  X_BUF \DLX_EXinst__n0017<13>/XUSED  (
    .I(\DLX_EXinst__n0017<13>/FROM ),
    .O(DLX_EXinst__n0017[13])
  );
  X_BUF \DLX_EXinst__n0017<13>/YUSED  (
    .I(\DLX_EXinst__n0017<13>/GROM ),
    .O(DLX_EXinst__n0017[7])
  );
  defparam DLX_IFlc_md_mda9_a1.INIT = 16'h0A0A;
  X_LUT4 DLX_IFlc_md_mda9_a1 (
    .ADR0(DLX_IFlc_md_wint8),
    .ADR1(VCC),
    .ADR2(DLX_IFlc_pd_wint1),
    .ADR3(VCC),
    .O(\DLX_IFlc_md_wint9/FROM )
  );
  defparam DLX_IFlc_md_mda16_a1.INIT = 16'h0F00;
  X_LUT4 DLX_IFlc_md_mda16_a1 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IFlc_pd_wint1),
    .ADR3(DLX_IFlc_md_wint15),
    .O(\DLX_IFlc_md_wint9/GROM )
  );
  X_BUF \DLX_IFlc_md_wint9/XUSED  (
    .I(\DLX_IFlc_md_wint9/FROM ),
    .O(DLX_IFlc_md_wint9)
  );
  X_BUF \DLX_IFlc_md_wint9/YUSED  (
    .I(\DLX_IFlc_md_wint9/GROM ),
    .O(DLX_IFlc_md_wint16)
  );
  defparam DLX_IFlc_md_mda17_a1.INIT = 16'h00CC;
  X_LUT4 DLX_IFlc_md_mda17_a1 (
    .ADR0(VCC),
    .ADR1(DLX_IFlc_md_wint16),
    .ADR2(VCC),
    .ADR3(DLX_IFlc_pd_wint1),
    .O(\DLX_IFlc_md_wint17/FROM )
  );
  defparam DLX_IFlc_md_mda40_a1.INIT = 16'h2222;
  X_LUT4 DLX_IFlc_md_mda40_a1 (
    .ADR0(DLX_IFlc_md_wint39),
    .ADR1(DLX_IFlc_pd_wint1),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IFlc_md_wint17/GROM )
  );
  X_BUF \DLX_IFlc_md_wint17/XUSED  (
    .I(\DLX_IFlc_md_wint17/FROM ),
    .O(DLX_IFlc_md_wint17)
  );
  X_BUF \DLX_IFlc_md_wint17/YUSED  (
    .I(\DLX_IFlc_md_wint17/GROM ),
    .O(DLX_IFlc_md_wint40)
  );
  defparam DLX_EXinst_Ker630541.INIT = 16'hF5A0;
  X_LUT4 DLX_EXinst_Ker630541 (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[21]),
    .ADR3(DLX_IDinst_reg_out_A[19]),
    .O(\DLX_EXinst_N63056/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0026_Sh<18>1 .INIT = 16'hEE44;
  X_LUT4 \DLX_EXinst_Mshift__n0026_Sh<18>1  (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(DLX_EXinst_N63424),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N63056),
    .O(\DLX_EXinst_N63056/GROM )
  );
  X_BUF \DLX_EXinst_N63056/XUSED  (
    .I(\DLX_EXinst_N63056/FROM ),
    .O(DLX_EXinst_N63056)
  );
  X_BUF \DLX_EXinst_N63056/YUSED  (
    .I(\DLX_EXinst_N63056/GROM ),
    .O(\DLX_EXinst_Mshift__n0026_Sh[18] )
  );
  defparam \DLX_EXinst__n0006<19>219 .INIT = 16'hC808;
  X_LUT4 \DLX_EXinst__n0006<19>219  (
    .ADR0(\DLX_EXinst_Mshift__n0025_Sh[15] ),
    .ADR1(DLX_IDinst_reg_out_B[2]),
    .ADR2(DLX_IDinst_reg_out_B[3]),
    .ADR3(\DLX_EXinst_Mshift__n0025_Sh[7] ),
    .O(\CHOICE4990/FROM )
  );
  defparam DLX_EXinst_Ker641021.INIT = 16'hE4E4;
  X_LUT4 DLX_EXinst_Ker641021 (
    .ADR0(DLX_IDinst_reg_out_B[3]),
    .ADR1(\DLX_EXinst_Mshift__n0025_Sh[23] ),
    .ADR2(\DLX_EXinst_Mshift__n0025_Sh[15] ),
    .ADR3(VCC),
    .O(\CHOICE4990/GROM )
  );
  X_BUF \CHOICE4990/XUSED  (
    .I(\CHOICE4990/FROM ),
    .O(CHOICE4990)
  );
  X_BUF \CHOICE4990/YUSED  (
    .I(\CHOICE4990/GROM ),
    .O(DLX_EXinst_N64104)
  );
  defparam DLX_EXinst_Ker633371.INIT = 16'hACAC;
  X_LUT4 DLX_EXinst_Ker633371 (
    .ADR0(DLX_IDinst_reg_out_A[10]),
    .ADR1(DLX_IDinst_reg_out_A[8]),
    .ADR2(DLX_IDinst_IR_function_field[1]),
    .ADR3(VCC),
    .O(\DLX_EXinst_N63339/FROM )
  );
  defparam DLX_EXinst_Ker633021.INIT = 16'hB8B8;
  X_LUT4 DLX_EXinst_Ker633021 (
    .ADR0(DLX_IDinst_reg_out_A[10]),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(DLX_IDinst_reg_out_A[8]),
    .ADR3(VCC),
    .O(\DLX_EXinst_N63339/GROM )
  );
  X_BUF \DLX_EXinst_N63339/XUSED  (
    .I(\DLX_EXinst_N63339/FROM ),
    .O(DLX_EXinst_N63339)
  );
  X_BUF \DLX_EXinst_N63339/YUSED  (
    .I(\DLX_EXinst_N63339/GROM ),
    .O(DLX_EXinst_N63304)
  );
  defparam \DLX_EXinst__n0017<15>1 .INIT = 16'hD8D8;
  X_LUT4 \DLX_EXinst__n0017<15>1  (
    .ADR0(DLX_EXinst__n0030_1),
    .ADR1(DLX_IDinst_reg_out_B[15]),
    .ADR2(\DLX_IDinst_Imm[15] ),
    .ADR3(VCC),
    .O(\DLX_EXinst__n0017<15>/FROM )
  );
  defparam \DLX_EXinst__n0017<8>1 .INIT = 16'hFA50;
  X_LUT4 \DLX_EXinst__n0017<8>1  (
    .ADR0(DLX_EXinst__n0030_1),
    .ADR1(VCC),
    .ADR2(\DLX_IDinst_Imm[8] ),
    .ADR3(DLX_IDinst_reg_out_B[8]),
    .O(\DLX_EXinst__n0017<15>/GROM )
  );
  X_BUF \DLX_EXinst__n0017<15>/XUSED  (
    .I(\DLX_EXinst__n0017<15>/FROM ),
    .O(DLX_EXinst__n0017[15])
  );
  X_BUF \DLX_EXinst__n0017<15>/YUSED  (
    .I(\DLX_EXinst__n0017<15>/GROM ),
    .O(DLX_EXinst__n0017[8])
  );
  defparam DLX_EXinst_Ker630391.INIT = 16'hF3C0;
  X_LUT4 DLX_EXinst_Ker630391 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(DLX_IDinst_reg_out_A[15]),
    .ADR3(DLX_IDinst_reg_out_A[13]),
    .O(\DLX_EXinst_N63041/FROM )
  );
  defparam DLX_EXinst_Ker6426211.INIT = 16'hA820;
  X_LUT4 DLX_EXinst_Ker6426211 (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(DLX_IDinst_reg_out_B[3]),
    .ADR2(DLX_EXinst_N63284),
    .ADR3(DLX_EXinst_N63041),
    .O(\DLX_EXinst_N63041/GROM )
  );
  X_BUF \DLX_EXinst_N63041/XUSED  (
    .I(\DLX_EXinst_N63041/FROM ),
    .O(DLX_EXinst_N63041)
  );
  X_BUF \DLX_EXinst_N63041/YUSED  (
    .I(\DLX_EXinst_N63041/GROM ),
    .O(CHOICE1030)
  );
  defparam \DLX_EXinst__n0006<11>6 .INIT = 16'hECA0;
  X_LUT4 \DLX_EXinst__n0006<11>6  (
    .ADR0(DLX_EXinst_N66525),
    .ADR1(\DLX_EXinst_Mshift__n0028_Sh[59] ),
    .ADR2(\DLX_EXinst_Mshift__n0027_Sh[43] ),
    .ADR3(DLX_EXinst_N66373),
    .O(\CHOICE3917/FROM )
  );
  defparam \DLX_EXinst__n0006<10>6 .INIT = 16'hF888;
  X_LUT4 \DLX_EXinst__n0006<10>6  (
    .ADR0(DLX_EXinst_N66373),
    .ADR1(\DLX_EXinst_Mshift__n0028_Sh[58] ),
    .ADR2(DLX_EXinst_N66525),
    .ADR3(\DLX_EXinst_Mshift__n0027_Sh[42] ),
    .O(\CHOICE3917/GROM )
  );
  X_BUF \CHOICE3917/XUSED  (
    .I(\CHOICE3917/FROM ),
    .O(CHOICE3917)
  );
  X_BUF \CHOICE3917/YUSED  (
    .I(\CHOICE3917/GROM ),
    .O(CHOICE4487)
  );
  defparam \vga_top_vga1_helpcounter_Madd__n0000_Mxor_Result<1>_Result1 .INIT = 16'h0FF0;
  X_LUT4 \vga_top_vga1_helpcounter_Madd__n0000_Mxor_Result<1>_Result1  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_helpcounter[1]),
    .ADR3(vga_top_vga1_helpcounter[0]),
    .O(vga_top_vga1_helpcounter__n0000[1])
  );
  X_INV \vga_top_vga1_helpcounter<0>/BXMUX  (
    .I(vga_top_vga1_helpcounter[0]),
    .O(\vga_top_vga1_helpcounter<0>/BXMUXNOT )
  );
  defparam DLX_EXinst_Ker630641.INIT = 16'hF3C0;
  X_LUT4 DLX_EXinst_Ker630641 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(DLX_IDinst_reg_out_A[25]),
    .ADR3(DLX_IDinst_reg_out_A[23]),
    .O(\DLX_EXinst_N63066/FROM )
  );
  defparam DLX_EXinst_Ker664291.INIT = 16'h3120;
  X_LUT4 DLX_EXinst_Ker664291 (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(DLX_IDinst_reg_out_B_3_1),
    .ADR2(DLX_EXinst_N63780),
    .ADR3(DLX_EXinst_N63066),
    .O(\DLX_EXinst_N63066/GROM )
  );
  X_BUF \DLX_EXinst_N63066/XUSED  (
    .I(\DLX_EXinst_N63066/FROM ),
    .O(DLX_EXinst_N63066)
  );
  X_BUF \DLX_EXinst_N63066/YUSED  (
    .I(\DLX_EXinst_N63066/GROM ),
    .O(DLX_EXinst_N66431)
  );
  defparam \DLX_EXinst__n0006<19>42_SW0 .INIT = 16'h1111;
  X_LUT4 \DLX_EXinst__n0006<19>42_SW0  (
    .ADR0(DLX_IDinst_IR_opcode_field[0]),
    .ADR1(DLX_IDinst_reg_out_A[19]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\N127404/FROM )
  );
  defparam DLX_EXinst_Ker630491.INIT = 16'hB8B8;
  X_LUT4 DLX_EXinst_Ker630491 (
    .ADR0(DLX_IDinst_reg_out_A[19]),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(DLX_IDinst_reg_out_A[17]),
    .ADR3(VCC),
    .O(\N127404/GROM )
  );
  X_BUF \N127404/XUSED  (
    .I(\N127404/FROM ),
    .O(N127404)
  );
  X_BUF \N127404/YUSED  (
    .I(\N127404/GROM ),
    .O(DLX_EXinst_N63051)
  );
  defparam DLX_EXinst_Ker634021.INIT = 16'hE4E4;
  X_LUT4 DLX_EXinst_Ker634021 (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(DLX_IDinst_reg_out_A[8]),
    .ADR2(DLX_IDinst_reg_out_A[6]),
    .ADR3(VCC),
    .O(\DLX_EXinst_N63404/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0025_Sh<9>1 .INIT = 16'hEE44;
  X_LUT4 \DLX_EXinst_Mshift__n0025_Sh<9>1  (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(DLX_EXinst_N62856),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N63404),
    .O(\DLX_EXinst_N63404/GROM )
  );
  X_BUF \DLX_EXinst_N63404/XUSED  (
    .I(\DLX_EXinst_N63404/FROM ),
    .O(DLX_EXinst_N63404)
  );
  X_BUF \DLX_EXinst_N63404/YUSED  (
    .I(\DLX_EXinst_N63404/GROM ),
    .O(\DLX_EXinst_Mshift__n0025_Sh[9] )
  );
  defparam DLX_EXinst_Ker631551.INIT = 16'hFCFC;
  X_LUT4 DLX_EXinst_Ker631551 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_B[0]),
    .ADR2(DLX_IDinst_reg_out_B[1]),
    .ADR3(VCC),
    .O(\DLX_EXinst_N63157/GROM )
  );
  X_BUF \DLX_EXinst_N63157/YUSED  (
    .I(\DLX_EXinst_N63157/GROM ),
    .O(DLX_EXinst_N63157)
  );
  defparam DLX_EXinst_Ker630591.INIT = 16'hCACA;
  X_LUT4 DLX_EXinst_Ker630591 (
    .ADR0(DLX_IDinst_reg_out_A[21]),
    .ADR1(DLX_IDinst_reg_out_A[23]),
    .ADR2(DLX_IDinst_reg_out_B[1]),
    .ADR3(VCC),
    .O(\DLX_EXinst_N63061/FROM )
  );
  defparam DLX_EXinst_Ker62725_SW0.INIT = 16'hFA50;
  X_LUT4 DLX_EXinst_Ker62725_SW0 (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N63429),
    .ADR3(DLX_EXinst_N63061),
    .O(\DLX_EXinst_N63061/GROM )
  );
  X_BUF \DLX_EXinst_N63061/XUSED  (
    .I(\DLX_EXinst_N63061/FROM ),
    .O(DLX_EXinst_N63061)
  );
  X_BUF \DLX_EXinst_N63061/YUSED  (
    .I(\DLX_EXinst_N63061/GROM ),
    .O(N94057)
  );
  defparam DLX_EXinst_Ker632771.INIT = 16'hFA0A;
  X_LUT4 DLX_EXinst_Ker632771 (
    .ADR0(DLX_IDinst_reg_out_A[24]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_IR_function_field[1]),
    .ADR3(DLX_IDinst_reg_out_A[26]),
    .O(\DLX_EXinst_N63279/FROM )
  );
  defparam DLX_EXinst_Ker633071.INIT = 16'hF0AA;
  X_LUT4 DLX_EXinst_Ker633071 (
    .ADR0(DLX_IDinst_reg_out_A[26]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[24]),
    .ADR3(DLX_IDinst_IR_function_field[1]),
    .O(\DLX_EXinst_N63279/GROM )
  );
  X_BUF \DLX_EXinst_N63279/XUSED  (
    .I(\DLX_EXinst_N63279/FROM ),
    .O(DLX_EXinst_N63279)
  );
  X_BUF \DLX_EXinst_N63279/YUSED  (
    .I(\DLX_EXinst_N63279/GROM ),
    .O(DLX_EXinst_N63309)
  );
  defparam \DLX_EXinst__n0006<17>42_SW0 .INIT = 16'h0303;
  X_LUT4 \DLX_EXinst__n0006<17>42_SW0  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[17]),
    .ADR2(DLX_IDinst_IR_opcode_field[0]),
    .ADR3(VCC),
    .O(\N127322/FROM )
  );
  defparam \DLX_EXinst__n0006<29>88_SW0 .INIT = 16'h0303;
  X_LUT4 \DLX_EXinst__n0006<29>88_SW0  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[29]),
    .ADR2(DLX_IDinst_IR_opcode_field[0]),
    .ADR3(VCC),
    .O(\N127322/GROM )
  );
  X_BUF \N127322/XUSED  (
    .I(\N127322/FROM ),
    .O(N127322)
  );
  X_BUF \N127322/YUSED  (
    .I(\N127322/GROM ),
    .O(N127374)
  );
  defparam DLX_IDinst__n04421.INIT = 16'h2033;
  X_LUT4 DLX_IDinst__n04421 (
    .ADR0(DLX_IDinst_slot_num_FFd1),
    .ADR1(DLX_IDinst__n0335),
    .ADR2(DLX_IDinst_delay_slot),
    .ADR3(DLX_IDinst__n0331),
    .O(\DLX_IDinst__n0442/FROM )
  );
  defparam DLX_IDinst__n0443_SW0.INIT = 16'hCFCF;
  X_LUT4 DLX_IDinst__n0443_SW0 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_delay_slot),
    .ADR2(DLX_IDinst_slot_num_FFd1),
    .ADR3(VCC),
    .O(\DLX_IDinst__n0442/GROM )
  );
  X_BUF \DLX_IDinst__n0442/XUSED  (
    .I(\DLX_IDinst__n0442/FROM ),
    .O(DLX_IDinst__n0442)
  );
  X_BUF \DLX_IDinst__n0442/YUSED  (
    .I(\DLX_IDinst__n0442/GROM ),
    .O(N90101)
  );
  defparam DLX_EXinst_Ker634121.INIT = 16'hF3C0;
  X_LUT4 DLX_EXinst_Ker634121 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(DLX_IDinst_reg_out_A[16]),
    .ADR3(DLX_IDinst_reg_out_A[14]),
    .O(\DLX_EXinst_N63414/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0026_Sh<13>1 .INIT = 16'hFC0C;
  X_LUT4 \DLX_EXinst_Mshift__n0026_Sh<13>1  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N63041),
    .ADR2(DLX_IDinst_reg_out_B[0]),
    .ADR3(DLX_EXinst_N63414),
    .O(\DLX_EXinst_N63414/GROM )
  );
  X_BUF \DLX_EXinst_N63414/XUSED  (
    .I(\DLX_EXinst_N63414/FROM ),
    .O(DLX_EXinst_N63414)
  );
  X_BUF \DLX_EXinst_N63414/YUSED  (
    .I(\DLX_EXinst_N63414/GROM ),
    .O(\DLX_EXinst_Mshift__n0026_Sh[13] )
  );
  defparam DLX_EXinst_Ker629441.INIT = 16'hFA50;
  X_LUT4 DLX_EXinst_Ker629441 (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[6]),
    .ADR3(DLX_IDinst_reg_out_A[8]),
    .O(\DLX_EXinst_N62946/FROM )
  );
  defparam DLX_EXinst_Ker633321.INIT = 16'hEE22;
  X_LUT4 DLX_EXinst_Ker633321 (
    .ADR0(DLX_IDinst_reg_out_A[6]),
    .ADR1(DLX_IDinst_IR_function_field[1]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[8]),
    .O(\DLX_EXinst_N62946/GROM )
  );
  X_BUF \DLX_EXinst_N62946/XUSED  (
    .I(\DLX_EXinst_N62946/FROM ),
    .O(DLX_EXinst_N62946)
  );
  X_BUF \DLX_EXinst_N62946/YUSED  (
    .I(\DLX_EXinst_N62946/GROM ),
    .O(DLX_EXinst_N63334)
  );
  defparam \DLX_EXinst__n0006<21>41_SW0 .INIT = 16'hDFDF;
  X_LUT4 \DLX_EXinst__n0006<21>41_SW0  (
    .ADR0(DLX_EXinst_N62821),
    .ADR1(DLX_IDinst_IR_function_field[3]),
    .ADR2(DLX_IDinst_IR_function_field[4]),
    .ADR3(VCC),
    .O(\N127126/FROM )
  );
  defparam \DLX_EXinst__n0006<23>41_SW0 .INIT = 16'hAFFF;
  X_LUT4 \DLX_EXinst__n0006<23>41_SW0  (
    .ADR0(DLX_IDinst_IR_function_field[3]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N62831),
    .ADR3(DLX_IDinst_IR_function_field[4]),
    .O(\N127126/GROM )
  );
  X_BUF \N127126/XUSED  (
    .I(\N127126/FROM ),
    .O(N127126)
  );
  X_BUF \N127126/YUSED  (
    .I(\N127126/GROM ),
    .O(N127189)
  );
  defparam DLX_IDinst_Ker70883.INIT = 16'h0040;
  X_LUT4 DLX_IDinst_Ker70883 (
    .ADR0(N90255),
    .ADR1(DLX_IDinst_N70610),
    .ADR2(DLX_IDinst_N70909),
    .ADR3(DLX_IDinst__n0348),
    .O(\DLX_IDinst_N70885/FROM )
  );
  defparam DLX_IDinst_Ker70070.INIT = 16'hAE0C;
  X_LUT4 DLX_IDinst_Ker70070 (
    .ADR0(DLX_IDinst_N70635),
    .ADR1(N100191),
    .ADR2(DLX_IDinst_IR_latched[30]),
    .ADR3(DLX_IDinst_N70885),
    .O(\DLX_IDinst_N70885/GROM )
  );
  X_BUF \DLX_IDinst_N70885/XUSED  (
    .I(\DLX_IDinst_N70885/FROM ),
    .O(DLX_IDinst_N70885)
  );
  X_BUF \DLX_IDinst_N70885/YUSED  (
    .I(\DLX_IDinst_N70885/GROM ),
    .O(DLX_IDinst_N70072)
  );
  defparam DM_delay_inst_wint101.INIT = 16'h00FF;
  X_LUT4 DM_delay_inst_wint101 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DM_delay_inst_wint9),
    .O(\DM_delay_inst_wint10/GROM )
  );
  X_BUF \DM_delay_inst_wint10/YUSED  (
    .I(\DM_delay_inst_wint10/GROM ),
    .O(DM_delay_inst_wint10)
  );
  defparam \DLX_IDinst_regB_eff<1>1 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst_regB_eff<1>1  (
    .ADR0(DLX_IDinst_reg_out_B_RF[1]),
    .ADR1(DLX_IDinst_N70716),
    .ADR2(DLX_RF_data_in[1]),
    .ADR3(DLX_IDinst__n0145),
    .O(\DLX_IDinst_regB_eff<1>/FROM )
  );
  defparam \DLX_IDinst_regB_eff<10>1 .INIT = 16'hEAC0;
  X_LUT4 \DLX_IDinst_regB_eff<10>1  (
    .ADR0(DLX_MEMinst_RF_data_in[10]),
    .ADR1(DLX_IDinst_N70716),
    .ADR2(DLX_IDinst_reg_out_B_RF[10]),
    .ADR3(DLX_IDinst__n0145),
    .O(\DLX_IDinst_regB_eff<1>/GROM )
  );
  X_BUF \DLX_IDinst_regB_eff<1>/XUSED  (
    .I(\DLX_IDinst_regB_eff<1>/FROM ),
    .O(DLX_IDinst_regB_eff[1])
  );
  X_BUF \DLX_IDinst_regB_eff<1>/YUSED  (
    .I(\DLX_IDinst_regB_eff<1>/GROM ),
    .O(DLX_IDinst_regB_eff[10])
  );
  defparam DLX_IFlc_md_mda34_a1.INIT = 16'h2222;
  X_LUT4 DLX_IFlc_md_mda34_a1 (
    .ADR0(DLX_IFlc_md_wint33),
    .ADR1(DLX_IFlc_pd_wint1),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IFlc_md_wint34/FROM )
  );
  defparam DLX_IFlc_md_mda35_a1.INIT = 16'h5500;
  X_LUT4 DLX_IFlc_md_mda35_a1 (
    .ADR0(DLX_IFlc_pd_wint1),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IFlc_md_wint34),
    .O(\DLX_IFlc_md_wint34/GROM )
  );
  X_BUF \DLX_IFlc_md_wint34/XUSED  (
    .I(\DLX_IFlc_md_wint34/FROM ),
    .O(DLX_IFlc_md_wint34)
  );
  X_BUF \DLX_IFlc_md_wint34/YUSED  (
    .I(\DLX_IFlc_md_wint34/GROM ),
    .O(DLX_IFlc_md_wint35)
  );
  defparam DLX_IFlc_md_mda26_a1.INIT = 16'h3300;
  X_LUT4 DLX_IFlc_md_mda26_a1 (
    .ADR0(VCC),
    .ADR1(DLX_IFlc_pd_wint1),
    .ADR2(VCC),
    .ADR3(DLX_IFlc_md_wint25),
    .O(\DLX_IFlc_md_wint26/FROM )
  );
  defparam DLX_IFlc_md_mda27_a1.INIT = 16'h5500;
  X_LUT4 DLX_IFlc_md_mda27_a1 (
    .ADR0(DLX_IFlc_pd_wint1),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IFlc_md_wint26),
    .O(\DLX_IFlc_md_wint26/GROM )
  );
  X_BUF \DLX_IFlc_md_wint26/XUSED  (
    .I(\DLX_IFlc_md_wint26/FROM ),
    .O(DLX_IFlc_md_wint26)
  );
  X_BUF \DLX_IFlc_md_wint26/YUSED  (
    .I(\DLX_IFlc_md_wint26/GROM ),
    .O(DLX_IFlc_md_wint27)
  );
  defparam DLX_IDinst_Ker6960436.INIT = 16'hB0BB;
  X_LUT4 DLX_IDinst_Ker6960436 (
    .ADR0(DLX_IDinst__n0002),
    .ADR1(DLX_IDinst__n0077),
    .ADR2(DLX_IDinst__n0004),
    .ADR3(DLX_IDinst__n0075),
    .O(\CHOICE2099/FROM )
  );
  defparam DLX_IDinst__n0108123.INIT = 16'h80C0;
  X_LUT4 DLX_IDinst__n0108123 (
    .ADR0(DLX_IDinst__n0002),
    .ADR1(DLX_IDinst_N70035),
    .ADR2(CHOICE3457),
    .ADR3(DLX_IDinst__n0077),
    .O(\CHOICE2099/GROM )
  );
  X_BUF \CHOICE2099/XUSED  (
    .I(\CHOICE2099/FROM ),
    .O(CHOICE2099)
  );
  X_BUF \CHOICE2099/YUSED  (
    .I(\CHOICE2099/GROM ),
    .O(CHOICE3458)
  );
  defparam DM_delay_inst_wint111.INIT = 16'h00FF;
  X_LUT4 DM_delay_inst_wint111 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DM_delay_inst_wint10),
    .O(\DM_delay_inst_wint11/GROM )
  );
  X_BUF \DM_delay_inst_wint11/YUSED  (
    .I(\DM_delay_inst_wint11/GROM ),
    .O(DM_delay_inst_wint11)
  );
  defparam DLX_EXinst_Ker634221.INIT = 16'hCCAA;
  X_LUT4 DLX_EXinst_Ker634221 (
    .ADR0(DLX_IDinst_reg_out_A[18]),
    .ADR1(DLX_IDinst_reg_out_A[20]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[1]),
    .O(\DLX_EXinst_N63424/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0026_Sh<17>1 .INIT = 16'hFA50;
  X_LUT4 \DLX_EXinst_Mshift__n0026_Sh<17>1  (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N63051),
    .ADR3(DLX_EXinst_N63424),
    .O(\DLX_EXinst_N63424/GROM )
  );
  X_BUF \DLX_EXinst_N63424/XUSED  (
    .I(\DLX_EXinst_N63424/FROM ),
    .O(DLX_EXinst_N63424)
  );
  X_BUF \DLX_EXinst_N63424/YUSED  (
    .I(\DLX_EXinst_N63424/GROM ),
    .O(\DLX_EXinst_Mshift__n0026_Sh[17] )
  );
  defparam DLX_EXinst_Ker64558.INIT = 16'hF3C0;
  X_LUT4 DLX_EXinst_Ker64558 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_IR_function_field[3]),
    .ADR2(\DLX_EXinst_Mshift__n0028_Sh[21] ),
    .ADR3(N93955),
    .O(\DLX_EXinst_N64560/FROM )
  );
  defparam DLX_EXinst_Ker640701.INIT = 16'hEE44;
  X_LUT4 DLX_EXinst_Ker640701 (
    .ADR0(DLX_IDinst_IR_function_field[3]),
    .ADR1(\DLX_EXinst_Mshift__n0027_Sh[19] ),
    .ADR2(VCC),
    .ADR3(\DLX_EXinst_Mshift__n0027_Sh[11] ),
    .O(\DLX_EXinst_N64560/GROM )
  );
  X_BUF \DLX_EXinst_N64560/XUSED  (
    .I(\DLX_EXinst_N64560/FROM ),
    .O(DLX_EXinst_N64560)
  );
  X_BUF \DLX_EXinst_N64560/YUSED  (
    .I(\DLX_EXinst_N64560/GROM ),
    .O(DLX_EXinst_N64072)
  );
  defparam DLX_EXinst_Ker635021.INIT = 16'hD8D8;
  X_LUT4 DLX_EXinst_Ker635021 (
    .ADR0(DLX_IDinst_IR_function_field_1_1),
    .ADR1(DLX_IDinst_reg_out_A[18]),
    .ADR2(DLX_IDinst_reg_out_A[16]),
    .ADR3(VCC),
    .O(\DLX_EXinst_N63504/FROM )
  );
  defparam DLX_EXinst_Ker6480710.INIT = 16'hA820;
  X_LUT4 DLX_EXinst_Ker6480710 (
    .ADR0(DLX_IDinst_IR_function_field[3]),
    .ADR1(DLX_IDinst_IR_function_field[0]),
    .ADR2(DLX_EXinst_N62996),
    .ADR3(DLX_EXinst_N63504),
    .O(\DLX_EXinst_N63504/GROM )
  );
  X_BUF \DLX_EXinst_N63504/XUSED  (
    .I(\DLX_EXinst_N63504/FROM ),
    .O(DLX_EXinst_N63504)
  );
  X_BUF \DLX_EXinst_N63504/YUSED  (
    .I(\DLX_EXinst_N63504/GROM ),
    .O(CHOICE1090)
  );
  defparam DM_delay_inst_wint121.INIT = 16'h3333;
  X_LUT4 DM_delay_inst_wint121 (
    .ADR0(VCC),
    .ADR1(DM_delay_inst_wint11),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DM_delay_inst_wint12/GROM )
  );
  X_BUF \DM_delay_inst_wint12/YUSED  (
    .I(\DM_delay_inst_wint12/GROM ),
    .O(DM_delay_inst_wint12)
  );
  defparam DM_delay_inst_wint201.INIT = 16'h3333;
  X_LUT4 DM_delay_inst_wint201 (
    .ADR0(VCC),
    .ADR1(DM_delay_inst_wint19),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DM_delay_inst_wint20/FROM )
  );
  defparam DM_delay_inst_wint211.INIT = 16'h00FF;
  X_LUT4 DM_delay_inst_wint211 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DM_delay_inst_wint20),
    .O(\DM_delay_inst_wint20/GROM )
  );
  X_BUF \DM_delay_inst_wint20/XUSED  (
    .I(\DM_delay_inst_wint20/FROM ),
    .O(DM_delay_inst_wint20)
  );
  X_BUF \DM_delay_inst_wint20/YUSED  (
    .I(\DM_delay_inst_wint20/GROM ),
    .O(DM_delay_inst_wint21)
  );
  defparam DLX_EXlc_slave_ctrlEX__n0001_SW111.INIT = 16'hF000;
  X_LUT4 DLX_EXlc_slave_ctrlEX__n0001_SW111 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_EXlc_master_ctrlEX_nro),
    .ADR3(CHOICE45),
    .O(\DLX_EXlc_slave_ctrlEX_l/GROM )
  );
  X_BUF \DLX_EXlc_slave_ctrlEX_l/YUSED  (
    .I(\DLX_EXlc_slave_ctrlEX_l/GROM ),
    .O(DLX_EXlc_slave_ctrlEX_l)
  );
  defparam \DLX_IDinst_regB_eff<2>1 .INIT = 16'hECA0;
  X_LUT4 \DLX_IDinst_regB_eff<2>1  (
    .ADR0(DLX_IDinst_N70716),
    .ADR1(DLX_RF_data_in[2]),
    .ADR2(DLX_IDinst_reg_out_B_RF[2]),
    .ADR3(DLX_IDinst__n0145),
    .O(\DLX_IDinst_regB_eff<2>/FROM )
  );
  defparam \DLX_IDinst_regB_eff<11>1 .INIT = 16'hEAC0;
  X_LUT4 \DLX_IDinst_regB_eff<11>1  (
    .ADR0(DLX_MEMinst_RF_data_in[11]),
    .ADR1(DLX_IDinst_reg_out_B_RF[11]),
    .ADR2(DLX_IDinst_N70716),
    .ADR3(DLX_IDinst__n0145),
    .O(\DLX_IDinst_regB_eff<2>/GROM )
  );
  X_BUF \DLX_IDinst_regB_eff<2>/XUSED  (
    .I(\DLX_IDinst_regB_eff<2>/FROM ),
    .O(DLX_IDinst_regB_eff[2])
  );
  X_BUF \DLX_IDinst_regB_eff<2>/YUSED  (
    .I(\DLX_IDinst_regB_eff<2>/GROM ),
    .O(DLX_IDinst_regB_eff[11])
  );
  defparam \DLX_EXinst__n0006<0>697_SW0 .INIT = 16'h8000;
  X_LUT4 \DLX_EXinst__n0006<0>697_SW0  (
    .ADR0(\DLX_IDinst_Imm[5] ),
    .ADR1(DLX_IDinst_reg_out_A[31]),
    .ADR2(CHOICE3408),
    .ADR3(CHOICE3377),
    .O(\N126811/FROM )
  );
  defparam DLX_EXinst_Ker631831.INIT = 16'hFF40;
  X_LUT4 DLX_EXinst_Ker631831 (
    .ADR0(\DLX_IDinst_Imm[5] ),
    .ADR1(CHOICE3377),
    .ADR2(CHOICE3408),
    .ADR3(DLX_EXinst_N66507),
    .O(\N126811/GROM )
  );
  X_BUF \N126811/XUSED  (
    .I(\N126811/FROM ),
    .O(N126811)
  );
  X_BUF \N126811/YUSED  (
    .I(\N126811/GROM ),
    .O(DLX_EXinst_N63185)
  );
  defparam DLX_EXinst_Ker6615516.INIT = 16'h66AA;
  X_LUT4 DLX_EXinst_Ker6615516 (
    .ADR0(\DLX_IDinst_Imm[5] ),
    .ADR1(DLX_IDinst_IR_function_field_3_1),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_IR_function_field_2_1),
    .O(\CHOICE1321/FROM )
  );
  defparam DLX_EXinst_Ker651031.INIT = 16'hFC0C;
  X_LUT4 DLX_EXinst_Ker651031 (
    .ADR0(VCC),
    .ADR1(\DLX_EXinst_Mshift__n0028_Sh[8] ),
    .ADR2(DLX_IDinst_IR_function_field_3_1),
    .ADR3(\DLX_EXinst_Mshift__n0028_Sh[16] ),
    .O(\CHOICE1321/GROM )
  );
  X_BUF \CHOICE1321/XUSED  (
    .I(\CHOICE1321/FROM ),
    .O(CHOICE1321)
  );
  X_BUF \CHOICE1321/YUSED  (
    .I(\CHOICE1321/GROM ),
    .O(DLX_EXinst_N65105)
  );
  defparam DLX_EXinst_Ker630791.INIT = 16'hAEAA;
  X_LUT4 DLX_EXinst_Ker630791 (
    .ADR0(DLX_EXinst_N66431),
    .ADR1(DLX_IDinst_reg_out_A[31]),
    .ADR2(DLX_EXinst_N63157),
    .ADR3(DLX_IDinst_reg_out_B[3]),
    .O(\DLX_EXinst_N63081/FROM )
  );
  defparam DLX_EXinst_Ker6487795.INIT = 16'h7520;
  X_LUT4 DLX_EXinst_Ker6487795 (
    .ADR0(DLX_IDinst_reg_out_B_2_1),
    .ADR1(DLX_IDinst_reg_out_B_3_1),
    .ADR2(\DLX_EXinst_Mshift__n0023_Sh[27] ),
    .ADR3(DLX_EXinst_N63081),
    .O(\DLX_EXinst_N63081/GROM )
  );
  X_BUF \DLX_EXinst_N63081/XUSED  (
    .I(\DLX_EXinst_N63081/FROM ),
    .O(DLX_EXinst_N63081)
  );
  X_BUF \DLX_EXinst_N63081/YUSED  (
    .I(\DLX_EXinst_N63081/GROM ),
    .O(CHOICE2997)
  );
  defparam DLX_EXinst_Ker634071.INIT = 16'hBB88;
  X_LUT4 DLX_EXinst_Ker634071 (
    .ADR0(DLX_IDinst_reg_out_A[14]),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[12]),
    .O(\DLX_EXinst_N63409/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0026_Sh<11>1 .INIT = 16'hEE22;
  X_LUT4 \DLX_EXinst_Mshift__n0026_Sh<11>1  (
    .ADR0(DLX_EXinst_N63036),
    .ADR1(DLX_IDinst_reg_out_B[0]),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N63409),
    .O(\DLX_EXinst_N63409/GROM )
  );
  X_BUF \DLX_EXinst_N63409/XUSED  (
    .I(\DLX_EXinst_N63409/FROM ),
    .O(DLX_EXinst_N63409)
  );
  X_BUF \DLX_EXinst_N63409/YUSED  (
    .I(\DLX_EXinst_N63409/GROM ),
    .O(\DLX_EXinst_Mshift__n0026_Sh[11] )
  );
  defparam DLX_EXinst_Ker633271.INIT = 16'hD8D8;
  X_LUT4 DLX_EXinst_Ker633271 (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(DLX_IDinst_reg_out_A[12]),
    .ADR2(DLX_IDinst_reg_out_A[10]),
    .ADR3(VCC),
    .O(\DLX_EXinst_N63329/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<9>1 .INIT = 16'hFC0C;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<9>1  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N62951),
    .ADR2(DLX_IDinst_reg_out_B[0]),
    .ADR3(DLX_EXinst_N63329),
    .O(\DLX_EXinst_N63329/GROM )
  );
  X_BUF \DLX_EXinst_N63329/XUSED  (
    .I(\DLX_EXinst_N63329/FROM ),
    .O(DLX_EXinst_N63329)
  );
  X_BUF \DLX_EXinst_N63329/YUSED  (
    .I(\DLX_EXinst_N63329/GROM ),
    .O(\DLX_EXinst_Mshift__n0023_Sh[9] )
  );
  defparam \DLX_EXinst__n0006<24>9 .INIT = 16'hF020;
  X_LUT4 \DLX_EXinst__n0006<24>9  (
    .ADR0(DLX_EXinst__n0080),
    .ADR1(\DLX_IDinst_Imm[31] ),
    .ADR2(DLX_IDinst_reg_out_A[24]),
    .ADR3(DLX_EXinst__n0079),
    .O(\CHOICE3736/FROM )
  );
  defparam \DLX_EXinst__n0006<21>9 .INIT = 16'hA2A0;
  X_LUT4 \DLX_EXinst__n0006<21>9  (
    .ADR0(DLX_IDinst_reg_out_A[21]),
    .ADR1(\DLX_IDinst_Imm[31] ),
    .ADR2(DLX_EXinst__n0079),
    .ADR3(DLX_EXinst__n0080),
    .O(\CHOICE3736/GROM )
  );
  X_BUF \CHOICE3736/XUSED  (
    .I(\CHOICE3736/FROM ),
    .O(CHOICE3736)
  );
  X_BUF \CHOICE3736/YUSED  (
    .I(\CHOICE3736/GROM ),
    .O(CHOICE4164)
  );
  defparam DM_delay_inst_wint131.INIT = 16'h00FF;
  X_LUT4 DM_delay_inst_wint131 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DM_delay_inst_wint12),
    .O(\DM_delay_inst_wint13/GROM )
  );
  X_BUF \DM_delay_inst_wint13/YUSED  (
    .I(\DM_delay_inst_wint13/GROM ),
    .O(DM_delay_inst_wint13)
  );
  defparam DLX_EXinst_Ker651733.INIT = 16'h5404;
  X_LUT4 DLX_EXinst_Ker651733 (
    .ADR0(DLX_IDinst_reg_out_B_3_1),
    .ADR1(DLX_IDinst_reg_out_A[24]),
    .ADR2(DLX_IDinst_reg_out_B[1]),
    .ADR3(DLX_IDinst_reg_out_A[22]),
    .O(\CHOICE1184/FROM )
  );
  defparam DLX_EXinst_Ker634321.INIT = 16'hD8D8;
  X_LUT4 DLX_EXinst_Ker634321 (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(DLX_IDinst_reg_out_A[24]),
    .ADR2(DLX_IDinst_reg_out_A[22]),
    .ADR3(VCC),
    .O(\CHOICE1184/GROM )
  );
  X_BUF \CHOICE1184/XUSED  (
    .I(\CHOICE1184/FROM ),
    .O(CHOICE1184)
  );
  X_BUF \CHOICE1184/YUSED  (
    .I(\CHOICE1184/GROM ),
    .O(DLX_EXinst_N63434)
  );
  defparam DLX_EXinst_Ker637781.INIT = 16'hF5A0;
  X_LUT4 DLX_EXinst_Ker637781 (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[26]),
    .ADR3(DLX_IDinst_reg_out_A[24]),
    .O(\DLX_EXinst_N63780/FROM )
  );
  defparam DLX_EXinst_Ker632721.INIT = 16'hCACA;
  X_LUT4 DLX_EXinst_Ker632721 (
    .ADR0(DLX_IDinst_reg_out_A[26]),
    .ADR1(DLX_IDinst_reg_out_A[24]),
    .ADR2(DLX_IDinst_reg_out_B[1]),
    .ADR3(VCC),
    .O(\DLX_EXinst_N63780/GROM )
  );
  X_BUF \DLX_EXinst_N63780/XUSED  (
    .I(\DLX_EXinst_N63780/FROM ),
    .O(DLX_EXinst_N63780)
  );
  X_BUF \DLX_EXinst_N63780/YUSED  (
    .I(\DLX_EXinst_N63780/GROM ),
    .O(DLX_EXinst_N63274)
  );
  defparam DLX_EXinst_Ker643121.INIT = 16'hF3C0;
  X_LUT4 DLX_EXinst_Ker643121 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_IR_function_field[3]),
    .ADR2(\DLX_EXinst_Mshift__n0027_Sh[15] ),
    .ADR3(\DLX_EXinst_Mshift__n0027_Sh[23] ),
    .O(\DLX_EXinst_N64314/FROM )
  );
  defparam \DLX_EXinst__n0006<27>51 .INIT = 16'hC808;
  X_LUT4 \DLX_EXinst__n0006<27>51  (
    .ADR0(N100919),
    .ADR1(DLX_EXinst__n0081),
    .ADR2(DLX_IDinst_IR_function_field[2]),
    .ADR3(DLX_EXinst_N64314),
    .O(\DLX_EXinst_N64314/GROM )
  );
  X_BUF \DLX_EXinst_N64314/XUSED  (
    .I(\DLX_EXinst_N64314/FROM ),
    .O(DLX_EXinst_N64314)
  );
  X_BUF \DLX_EXinst_N64314/YUSED  (
    .I(\DLX_EXinst_N64314/GROM ),
    .O(CHOICE4628)
  );
  defparam DLX_EXinst_Ker635121.INIT = 16'hDD88;
  X_LUT4 DLX_EXinst_Ker635121 (
    .ADR0(DLX_IDinst_IR_function_field_1_1),
    .ADR1(DLX_IDinst_reg_out_A[22]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[20]),
    .O(\DLX_EXinst_N63514/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0028_Sh<19>1 .INIT = 16'hFA50;
  X_LUT4 \DLX_EXinst_Mshift__n0028_Sh<19>1  (
    .ADR0(DLX_IDinst_IR_function_field_0_1),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N63006),
    .ADR3(DLX_EXinst_N63514),
    .O(\DLX_EXinst_N63514/GROM )
  );
  X_BUF \DLX_EXinst_N63514/XUSED  (
    .I(\DLX_EXinst_N63514/FROM ),
    .O(DLX_EXinst_N63514)
  );
  X_BUF \DLX_EXinst_N63514/YUSED  (
    .I(\DLX_EXinst_N63514/GROM ),
    .O(\DLX_EXinst_Mshift__n0028_Sh[19] )
  );
  defparam DM_delay_inst_wint141.INIT = 16'h0F0F;
  X_LUT4 DM_delay_inst_wint141 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DM_delay_inst_wint13),
    .ADR3(VCC),
    .O(\DM_delay_inst_wint14/GROM )
  );
  X_BUF \DM_delay_inst_wint14/YUSED  (
    .I(\DM_delay_inst_wint14/GROM ),
    .O(DM_delay_inst_wint14)
  );
  defparam DLX_EXinst_mem_read_EX_1_1150.INIT = 1'b0;
  X_FF DLX_EXinst_mem_read_EX_1_1150 (
    .I(\DM_read/OD ),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DM_read/OFF/RST ),
    .O(DLX_EXinst_mem_read_EX_1)
  );
  X_OR2 \DM_read/OFF/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DM_read/OFF/RST )
  );
  defparam DM_delay_inst_wint221.INIT = 16'h3333;
  X_LUT4 DM_delay_inst_wint221 (
    .ADR0(VCC),
    .ADR1(DM_delay_inst_wint21),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DM_delay_inst_wint22/GROM )
  );
  X_BUF \DM_delay_inst_wint22/YUSED  (
    .I(\DM_delay_inst_wint22/GROM ),
    .O(DM_delay_inst_wint22)
  );
  defparam DM_delay_inst_wint301.INIT = 16'h3333;
  X_LUT4 DM_delay_inst_wint301 (
    .ADR0(VCC),
    .ADR1(DM_delay_inst_wint29),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DM_delay_inst_wint30/GROM )
  );
  X_BUF \DM_delay_inst_wint30/YUSED  (
    .I(\DM_delay_inst_wint30/GROM ),
    .O(DM_delay_inst_wint30)
  );
  defparam \DLX_IDinst_regB_eff<3>1 .INIT = 16'hEAC0;
  X_LUT4 \DLX_IDinst_regB_eff<3>1  (
    .ADR0(DLX_IDinst_N70716),
    .ADR1(DLX_IDinst__n0145),
    .ADR2(DLX_RF_data_in[3]),
    .ADR3(DLX_IDinst_reg_out_B_RF[3]),
    .O(\DLX_IDinst_regB_eff<3>/FROM )
  );
  defparam \DLX_IDinst_regB_eff<12>1 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst_regB_eff<12>1  (
    .ADR0(DLX_IDinst_N70716),
    .ADR1(DLX_IDinst_reg_out_B_RF[12]),
    .ADR2(DLX_MEMinst_RF_data_in[12]),
    .ADR3(DLX_IDinst__n0145),
    .O(\DLX_IDinst_regB_eff<3>/GROM )
  );
  X_BUF \DLX_IDinst_regB_eff<3>/XUSED  (
    .I(\DLX_IDinst_regB_eff<3>/FROM ),
    .O(DLX_IDinst_regB_eff[3])
  );
  X_BUF \DLX_IDinst_regB_eff<3>/YUSED  (
    .I(\DLX_IDinst_regB_eff<3>/GROM ),
    .O(DLX_IDinst_regB_eff[12])
  );
  defparam \DLX_IDinst_regB_eff<4>1 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst_regB_eff<4>1  (
    .ADR0(DLX_IDinst__n0145),
    .ADR1(DLX_RF_data_in[4]),
    .ADR2(DLX_IDinst_N70716),
    .ADR3(DLX_IDinst_reg_out_B_RF[4]),
    .O(\DLX_IDinst_regB_eff<4>/FROM )
  );
  defparam \DLX_IDinst_regB_eff<20>1 .INIT = 16'hECA0;
  X_LUT4 \DLX_IDinst_regB_eff<20>1  (
    .ADR0(DLX_IDinst__n0145),
    .ADR1(DLX_IDinst_reg_out_B_RF[20]),
    .ADR2(DLX_MEMinst_RF_data_in[20]),
    .ADR3(DLX_IDinst_N70716),
    .O(\DLX_IDinst_regB_eff<4>/GROM )
  );
  X_BUF \DLX_IDinst_regB_eff<4>/XUSED  (
    .I(\DLX_IDinst_regB_eff<4>/FROM ),
    .O(DLX_IDinst_regB_eff[4])
  );
  X_BUF \DLX_IDinst_regB_eff<4>/YUSED  (
    .I(\DLX_IDinst_regB_eff<4>/GROM ),
    .O(DLX_IDinst_regB_eff[20])
  );
  defparam DLX_EXinst_Ker634171.INIT = 16'hFA0A;
  X_LUT4 DLX_EXinst_Ker634171 (
    .ADR0(DLX_IDinst_reg_out_A[16]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[1]),
    .ADR3(DLX_IDinst_reg_out_A[18]),
    .O(\DLX_EXinst_N63419/FROM )
  );
  defparam DLX_EXinst_Ker6489710.INIT = 16'hE020;
  X_LUT4 DLX_EXinst_Ker6489710 (
    .ADR0(DLX_EXinst_N63304),
    .ADR1(DLX_IDinst_reg_out_B_3_1),
    .ADR2(DLX_IDinst_reg_out_B[0]),
    .ADR3(DLX_EXinst_N63419),
    .O(\DLX_EXinst_N63419/GROM )
  );
  X_BUF \DLX_EXinst_N63419/XUSED  (
    .I(\DLX_EXinst_N63419/FROM ),
    .O(DLX_EXinst_N63419)
  );
  X_BUF \DLX_EXinst_N63419/YUSED  (
    .I(\DLX_EXinst_N63419/GROM ),
    .O(CHOICE1162)
  );
  defparam \DLX_EXinst__n0006<28>331 .INIT = 16'hECA0;
  X_LUT4 \DLX_EXinst__n0006<28>331  (
    .ADR0(N126584),
    .ADR1(DLX_IDinst_reg_out_A[25]),
    .ADR2(DLX_EXinst__n0030),
    .ADR3(DLX_EXinst_N63712),
    .O(\CHOICE5244/FROM )
  );
  defparam \DLX_EXinst__n0006<28>363_SW0 .INIT = 16'hFFCE;
  X_LUT4 \DLX_EXinst__n0006<28>363_SW0  (
    .ADR0(CHOICE5204),
    .ADR1(CHOICE5247),
    .ADR2(DLX_EXinst__n0030),
    .ADR3(CHOICE5244),
    .O(\CHOICE5244/GROM )
  );
  X_BUF \CHOICE5244/XUSED  (
    .I(\CHOICE5244/FROM ),
    .O(CHOICE5244)
  );
  X_BUF \CHOICE5244/YUSED  (
    .I(\CHOICE5244/GROM ),
    .O(N126576)
  );
  defparam \DLX_EXinst__n0006<29>12 .INIT = 16'hF020;
  X_LUT4 \DLX_EXinst__n0006<29>12  (
    .ADR0(DLX_EXinst__n0080),
    .ADR1(\DLX_IDinst_Imm[31] ),
    .ADR2(DLX_IDinst_reg_out_A[29]),
    .ADR3(DLX_EXinst__n0079),
    .O(\CHOICE5333/FROM )
  );
  defparam \DLX_EXinst__n0006<22>9 .INIT = 16'h8A88;
  X_LUT4 \DLX_EXinst__n0006<22>9  (
    .ADR0(DLX_IDinst_reg_out_A[22]),
    .ADR1(DLX_EXinst__n0079),
    .ADR2(\DLX_IDinst_Imm[31] ),
    .ADR3(DLX_EXinst__n0080),
    .O(\CHOICE5333/GROM )
  );
  X_BUF \CHOICE5333/XUSED  (
    .I(\CHOICE5333/FROM ),
    .O(CHOICE5333)
  );
  X_BUF \CHOICE5333/YUSED  (
    .I(\CHOICE5333/GROM ),
    .O(CHOICE4098)
  );
  defparam DM_delay_inst_wint151.INIT = 16'h3333;
  X_LUT4 DM_delay_inst_wint151 (
    .ADR0(VCC),
    .ADR1(DM_delay_inst_wint14),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DM_delay_inst_wint15/GROM )
  );
  X_BUF \DM_delay_inst_wint15/YUSED  (
    .I(\DM_delay_inst_wint15/GROM ),
    .O(DM_delay_inst_wint15)
  );
  defparam DM_delay_inst_wint231.INIT = 16'h00FF;
  X_LUT4 DM_delay_inst_wint231 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DM_delay_inst_wint22),
    .O(\DM_delay_inst_wint23/GROM )
  );
  X_BUF \DM_delay_inst_wint23/YUSED  (
    .I(\DM_delay_inst_wint23/GROM ),
    .O(DM_delay_inst_wint23)
  );
  defparam DM_delay_inst_wint311.INIT = 16'h00FF;
  X_LUT4 DM_delay_inst_wint311 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DM_delay_inst_wint30),
    .O(\DM_delay_inst_wint31/GROM )
  );
  X_BUF \DM_delay_inst_wint31/YUSED  (
    .I(\DM_delay_inst_wint31/GROM ),
    .O(DM_delay_inst_wint31)
  );
  defparam DLX_EXinst_Ker629741.INIT = 16'hEE44;
  X_LUT4 DLX_EXinst_Ker629741 (
    .ADR0(DLX_IDinst_IR_function_field[1]),
    .ADR1(DLX_IDinst_reg_out_A[5]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[7]),
    .O(\DLX_EXinst_N62976/FROM )
  );
  defparam DLX_EXinst_Ker632821.INIT = 16'hDD88;
  X_LUT4 DLX_EXinst_Ker632821 (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(DLX_IDinst_reg_out_A[7]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[5]),
    .O(\DLX_EXinst_N62976/GROM )
  );
  X_BUF \DLX_EXinst_N62976/XUSED  (
    .I(\DLX_EXinst_N62976/FROM ),
    .O(DLX_EXinst_N62976)
  );
  X_BUF \DLX_EXinst_N62976/YUSED  (
    .I(\DLX_EXinst_N62976/GROM ),
    .O(DLX_EXinst_N63284)
  );
  defparam DLX_EXinst_Ker633621.INIT = 16'hCCF0;
  X_LUT4 DLX_EXinst_Ker633621 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[10]),
    .ADR2(DLX_IDinst_reg_out_A[12]),
    .ADR3(DLX_IDinst_reg_out_B[1]),
    .O(\DLX_EXinst_N63364/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0025_Sh<13>1 .INIT = 16'hFA50;
  X_LUT4 \DLX_EXinst_Mshift__n0025_Sh<13>1  (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N62866),
    .ADR3(DLX_EXinst_N63364),
    .O(\DLX_EXinst_N63364/GROM )
  );
  X_BUF \DLX_EXinst_N63364/XUSED  (
    .I(\DLX_EXinst_N63364/FROM ),
    .O(DLX_EXinst_N63364)
  );
  X_BUF \DLX_EXinst_N63364/YUSED  (
    .I(\DLX_EXinst_N63364/GROM ),
    .O(\DLX_EXinst_Mshift__n0025_Sh[13] )
  );
  defparam DLX_EXinst_Ker643221.INIT = 16'hE4E4;
  X_LUT4 DLX_EXinst_Ker643221 (
    .ADR0(DLX_IDinst_reg_out_B_3_1),
    .ADR1(\DLX_EXinst_Mshift__n0026_Sh[19] ),
    .ADR2(\DLX_EXinst_Mshift__n0023_Sh[27] ),
    .ADR3(VCC),
    .O(\DLX_EXinst_N64324/FROM )
  );
  defparam \DLX_EXinst__n0006<15>148 .INIT = 16'hC840;
  X_LUT4 \DLX_EXinst__n0006<15>148  (
    .ADR0(DLX_IDinst_reg_out_B[2]),
    .ADR1(DLX_EXinst_N66485),
    .ADR2(N97449),
    .ADR3(DLX_EXinst_N64324),
    .O(\DLX_EXinst_N64324/GROM )
  );
  X_BUF \DLX_EXinst_N64324/XUSED  (
    .I(\DLX_EXinst_N64324/FROM ),
    .O(DLX_EXinst_N64324)
  );
  X_BUF \DLX_EXinst_N64324/YUSED  (
    .I(\DLX_EXinst_N64324/GROM ),
    .O(CHOICE4842)
  );
  defparam \DLX_EXinst__n0006<10>59_SW0 .INIT = 16'h0055;
  X_LUT4 \DLX_EXinst__n0006<10>59_SW0  (
    .ADR0(DLX_IDinst_IR_opcode_field[0]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[10]),
    .O(\N127396/FROM )
  );
  defparam DLX_EXinst_Ker634421.INIT = 16'hFC0C;
  X_LUT4 DLX_EXinst_Ker634421 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[12]),
    .ADR2(DLX_IDinst_IR_function_field[1]),
    .ADR3(DLX_IDinst_reg_out_A[10]),
    .O(\N127396/GROM )
  );
  X_BUF \N127396/XUSED  (
    .I(\N127396/FROM ),
    .O(N127396)
  );
  X_BUF \N127396/YUSED  (
    .I(\N127396/GROM ),
    .O(DLX_EXinst_N63444)
  );
  defparam DLX_IFlc_master_ctrlIF_nl1.INIT = 16'h0F0F;
  X_LUT4 DLX_IFlc_master_ctrlIF_nl1 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IFlc_master_ctrlIF_l),
    .ADR3(VCC),
    .O(\DLX_clk_IF/FROM )
  );
  defparam DLX_RF_delay_inst_wint31.INIT = 16'h00FF;
  X_LUT4 DLX_RF_delay_inst_wint31 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_clk_IF),
    .O(\DLX_clk_IF/GROM )
  );
  X_BUF \DLX_clk_IF/XUSED  (
    .I(\DLX_clk_IF/FROM ),
    .O(DLX_clk_IF)
  );
  X_BUF \DLX_clk_IF/YUSED  (
    .I(\DLX_clk_IF/GROM ),
    .O(DLX_RF_delay_inst_wint3)
  );
  defparam DM_delay_inst_wint161.INIT = 16'h5555;
  X_LUT4 DM_delay_inst_wint161 (
    .ADR0(DM_delay_inst_wint15),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DM_delay_inst_wint16/GROM )
  );
  X_BUF \DM_delay_inst_wint16/YUSED  (
    .I(\DM_delay_inst_wint16/GROM ),
    .O(DM_delay_inst_wint16)
  );
  defparam DM_delay_inst_wint241.INIT = 16'h0F0F;
  X_LUT4 DM_delay_inst_wint241 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DM_delay_inst_wint23),
    .ADR3(VCC),
    .O(\DM_delay_inst_wint24/GROM )
  );
  X_BUF \DM_delay_inst_wint24/YUSED  (
    .I(\DM_delay_inst_wint24/GROM ),
    .O(DM_delay_inst_wint24)
  );
  defparam DM_delay_inst_wint321.INIT = 16'h3333;
  X_LUT4 DM_delay_inst_wint321 (
    .ADR0(VCC),
    .ADR1(DM_delay_inst_wint31),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DM_delay_inst_wint32/GROM )
  );
  X_BUF \DM_delay_inst_wint32/YUSED  (
    .I(\DM_delay_inst_wint32/GROM ),
    .O(DM_delay_inst_wint32)
  );
  defparam DM_delay_inst_wint401.INIT = 16'h3333;
  X_LUT4 DM_delay_inst_wint401 (
    .ADR0(VCC),
    .ADR1(DM_delay_inst_wint39),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DM_delay_inst_wint40/GROM )
  );
  X_BUF \DM_delay_inst_wint40/YUSED  (
    .I(\DM_delay_inst_wint40/GROM ),
    .O(DM_delay_inst_wint40)
  );
  defparam \DLX_IDinst_regB_eff<5>1 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst_regB_eff<5>1  (
    .ADR0(DLX_IDinst_N70716),
    .ADR1(DLX_IDinst_reg_out_B_RF[5]),
    .ADR2(DLX_RF_data_in[5]),
    .ADR3(DLX_IDinst__n0145),
    .O(\DLX_IDinst_regB_eff<5>/FROM )
  );
  defparam \DLX_IDinst_regB_eff<13>1 .INIT = 16'hEAC0;
  X_LUT4 \DLX_IDinst_regB_eff<13>1  (
    .ADR0(DLX_IDinst_reg_out_B_RF[13]),
    .ADR1(DLX_IDinst__n0145),
    .ADR2(DLX_MEMinst_RF_data_in[13]),
    .ADR3(DLX_IDinst_N70716),
    .O(\DLX_IDinst_regB_eff<5>/GROM )
  );
  X_BUF \DLX_IDinst_regB_eff<5>/XUSED  (
    .I(\DLX_IDinst_regB_eff<5>/FROM ),
    .O(DLX_IDinst_regB_eff[5])
  );
  X_BUF \DLX_IDinst_regB_eff<5>/YUSED  (
    .I(\DLX_IDinst_regB_eff<5>/GROM ),
    .O(DLX_IDinst_regB_eff[13])
  );
  defparam \DLX_IDinst_regB_eff<6>1 .INIT = 16'hEAC0;
  X_LUT4 \DLX_IDinst_regB_eff<6>1  (
    .ADR0(DLX_IDinst_N70716),
    .ADR1(DLX_IDinst__n0145),
    .ADR2(DLX_RF_data_in[6]),
    .ADR3(DLX_IDinst_reg_out_B_RF[6]),
    .O(\DLX_IDinst_regB_eff<6>/FROM )
  );
  defparam \DLX_IDinst_regB_eff<21>1 .INIT = 16'hECA0;
  X_LUT4 \DLX_IDinst_regB_eff<21>1  (
    .ADR0(DLX_IDinst_N70716),
    .ADR1(DLX_IDinst__n0145),
    .ADR2(DLX_IDinst_reg_out_B_RF[21]),
    .ADR3(DLX_MEMinst_RF_data_in[21]),
    .O(\DLX_IDinst_regB_eff<6>/GROM )
  );
  X_BUF \DLX_IDinst_regB_eff<6>/XUSED  (
    .I(\DLX_IDinst_regB_eff<6>/FROM ),
    .O(DLX_IDinst_regB_eff[6])
  );
  X_BUF \DLX_IDinst_regB_eff<6>/YUSED  (
    .I(\DLX_IDinst_regB_eff<6>/GROM ),
    .O(DLX_IDinst_regB_eff[21])
  );
  defparam DLX_EXinst_Ker627311.INIT = 16'hEEEE;
  X_LUT4 DLX_EXinst_Ker627311 (
    .ADR0(DLX_IDinst_IR_function_field[2]),
    .ADR1(DLX_IDinst_IR_function_field[3]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_EXinst_N62733/FROM )
  );
  defparam DLX_EXinst_Ker6581549.INIT = 16'h2000;
  X_LUT4 DLX_EXinst_Ker6581549 (
    .ADR0(N110065),
    .ADR1(\DLX_IDinst_Imm[5] ),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(DLX_EXinst_N62733),
    .O(\DLX_EXinst_N62733/GROM )
  );
  X_BUF \DLX_EXinst_N62733/XUSED  (
    .I(\DLX_EXinst_N62733/FROM ),
    .O(DLX_EXinst_N62733)
  );
  X_BUF \DLX_EXinst_N62733/YUSED  (
    .I(\DLX_EXinst_N62733/GROM ),
    .O(CHOICE2085)
  );
  defparam DLX_EXinst_Ker627071.INIT = 16'hCCF0;
  X_LUT4 DLX_EXinst_Ker627071 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[30]),
    .ADR2(DLX_IDinst_reg_out_A[29]),
    .ADR3(DLX_IDinst_IR_function_field[0]),
    .O(\DLX_EXinst_N62709/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0028_Sh<29>1 .INIT = 16'h2F20;
  X_LUT4 \DLX_EXinst_Mshift__n0028_Sh<29>1  (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(DLX_IDinst_IR_function_field_0_1),
    .ADR2(DLX_IDinst_IR_function_field_1_1),
    .ADR3(DLX_EXinst_N62709),
    .O(\DLX_EXinst_N62709/GROM )
  );
  X_BUF \DLX_EXinst_N62709/XUSED  (
    .I(\DLX_EXinst_N62709/FROM ),
    .O(DLX_EXinst_N62709)
  );
  X_BUF \DLX_EXinst_N62709/YUSED  (
    .I(\DLX_EXinst_N62709/GROM ),
    .O(\DLX_EXinst_Mshift__n0028_Sh[29] )
  );
  defparam DLX_EXinst_Ker632671.INIT = 16'h0B3B;
  X_LUT4 DLX_EXinst_Ker632671 (
    .ADR0(DLX_IDinst_IR_opcode_field[0]),
    .ADR1(DLX_IDinst_IR_opcode_field[1]),
    .ADR2(DLX_IDinst_IR_opcode_field[2]),
    .ADR3(DLX_IDinst_IR_opcode_field[3]),
    .O(\DLX_EXinst_N63269/FROM )
  );
  defparam DLX_EXinst_Ker6628813.INIT = 16'hAA00;
  X_LUT4 DLX_EXinst_Ker6628813 (
    .ADR0(DLX_IDinst_IR_opcode_field[5]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N63269),
    .O(\DLX_EXinst_N63269/GROM )
  );
  X_BUF \DLX_EXinst_N63269/XUSED  (
    .I(\DLX_EXinst_N63269/FROM ),
    .O(DLX_EXinst_N63269)
  );
  X_BUF \DLX_EXinst_N63269/YUSED  (
    .I(\DLX_EXinst_N63269/GROM ),
    .O(CHOICE1758)
  );
  defparam DLX_EXinst_Ker634271.INIT = 16'hD8D8;
  X_LUT4 DLX_EXinst_Ker634271 (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(DLX_IDinst_reg_out_A[22]),
    .ADR2(DLX_IDinst_reg_out_A[20]),
    .ADR3(VCC),
    .O(\DLX_EXinst_N63429/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0026_Sh<19>1 .INIT = 16'hFC30;
  X_LUT4 \DLX_EXinst_Mshift__n0026_Sh<19>1  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_B[0]),
    .ADR2(DLX_EXinst_N63056),
    .ADR3(DLX_EXinst_N63429),
    .O(\DLX_EXinst_N63429/GROM )
  );
  X_BUF \DLX_EXinst_N63429/XUSED  (
    .I(\DLX_EXinst_N63429/FROM ),
    .O(DLX_EXinst_N63429)
  );
  X_BUF \DLX_EXinst_N63429/YUSED  (
    .I(\DLX_EXinst_N63429/GROM ),
    .O(\DLX_EXinst_Mshift__n0026_Sh[19] )
  );
  defparam DLX_EXinst_Ker635071.INIT = 16'hF0AA;
  X_LUT4 DLX_EXinst_Ker635071 (
    .ADR0(DLX_IDinst_reg_out_A[18]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[20]),
    .ADR3(DLX_IDinst_IR_function_field_1_1),
    .O(\DLX_EXinst_N63509/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0028_Sh<17>1 .INIT = 16'hFA50;
  X_LUT4 \DLX_EXinst_Mshift__n0028_Sh<17>1  (
    .ADR0(DLX_IDinst_IR_function_field_0_1),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N63001),
    .ADR3(DLX_EXinst_N63509),
    .O(\DLX_EXinst_N63509/GROM )
  );
  X_BUF \DLX_EXinst_N63509/XUSED  (
    .I(\DLX_EXinst_N63509/FROM ),
    .O(DLX_EXinst_N63509)
  );
  X_BUF \DLX_EXinst_N63509/YUSED  (
    .I(\DLX_EXinst_N63509/GROM ),
    .O(\DLX_EXinst_Mshift__n0028_Sh[17] )
  );
  defparam \DLX_EXinst__n0006<16>306_SW0 .INIT = 16'hDCDC;
  X_LUT4 \DLX_EXinst__n0006<16>306_SW0  (
    .ADR0(DLX_IDinst_reg_out_A[16]),
    .ADR1(DLX_EXinst__n0046),
    .ADR2(DLX_EXinst__n0047),
    .ADR3(VCC),
    .O(\N126263/FROM )
  );
  defparam \DLX_EXinst__n0006<31>9 .INIT = 16'hD0C0;
  X_LUT4 \DLX_EXinst__n0006<31>9  (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(DLX_EXinst__n0046),
    .ADR2(DLX_IDinst_reg_out_B[31]),
    .ADR3(DLX_EXinst__n0047),
    .O(\N126263/GROM )
  );
  X_BUF \N126263/XUSED  (
    .I(\N126263/FROM ),
    .O(N126263)
  );
  X_BUF \N126263/YUSED  (
    .I(\N126263/GROM ),
    .O(CHOICE5740)
  );
  defparam \DLX_EXinst__n0006<27>9 .INIT = 16'h88C8;
  X_LUT4 \DLX_EXinst__n0006<27>9  (
    .ADR0(DLX_EXinst__n0079),
    .ADR1(DLX_IDinst_reg_out_A[27]),
    .ADR2(DLX_EXinst__n0080),
    .ADR3(\DLX_IDinst_Imm[31] ),
    .O(\CHOICE4610/FROM )
  );
  defparam \DLX_EXinst__n0006<23>9 .INIT = 16'hBA00;
  X_LUT4 \DLX_EXinst__n0006<23>9  (
    .ADR0(DLX_EXinst__n0079),
    .ADR1(\DLX_IDinst_Imm[31] ),
    .ADR2(DLX_EXinst__n0080),
    .ADR3(DLX_IDinst_reg_out_A[23]),
    .O(\CHOICE4610/GROM )
  );
  X_BUF \CHOICE4610/XUSED  (
    .I(\CHOICE4610/FROM ),
    .O(CHOICE4610)
  );
  X_BUF \CHOICE4610/YUSED  (
    .I(\CHOICE4610/GROM ),
    .O(CHOICE4032)
  );
  defparam DLX_IFinst_NPC_10_1_1151.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_10_1_1151 (
    .I(\NPC_eff<10>/OD ),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\NPC_eff<10>/OFF/RST ),
    .O(DLX_IFinst_NPC_10_1)
  );
  X_OR2 \NPC_eff<10>/OFF/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\NPC_eff<10>/OFF/RST )
  );
  defparam DM_delay_inst_wint171.INIT = 16'h00FF;
  X_LUT4 DM_delay_inst_wint171 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DM_delay_inst_wint16),
    .O(\DM_delay_inst_wint17/GROM )
  );
  X_BUF \DM_delay_inst_wint17/YUSED  (
    .I(\DM_delay_inst_wint17/GROM ),
    .O(DM_delay_inst_wint17)
  );
  defparam DM_delay_inst_wint251.INIT = 16'h00FF;
  X_LUT4 DM_delay_inst_wint251 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DM_delay_inst_wint24),
    .O(\DM_delay_inst_wint25/GROM )
  );
  X_BUF \DM_delay_inst_wint25/YUSED  (
    .I(\DM_delay_inst_wint25/GROM ),
    .O(DM_delay_inst_wint25)
  );
  defparam DM_delay_inst_wint331.INIT = 16'h0F0F;
  X_LUT4 DM_delay_inst_wint331 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DM_delay_inst_wint32),
    .ADR3(VCC),
    .O(\DM_delay_inst_wint33/GROM )
  );
  X_BUF \DM_delay_inst_wint33/YUSED  (
    .I(\DM_delay_inst_wint33/GROM ),
    .O(DM_delay_inst_wint33)
  );
  defparam \DLX_IDinst__n0106<0>_SW0 .INIT = 16'h3200;
  X_LUT4 \DLX_IDinst__n0106<0>_SW0  (
    .ADR0(DLX_IDinst_N69963),
    .ADR1(DLX_IDinst__n0364),
    .ADR2(CHOICE2100),
    .ADR3(DLX_IDinst_N69568),
    .O(\DLX_IDinst_rt_addr<0>/FROM )
  );
  defparam \DLX_IDinst__n0106<0> .INIT = 16'h8880;
  X_LUT4 \DLX_IDinst__n0106<0>  (
    .ADR0(DLX_IDinst_regB_index[0]),
    .ADR1(DLX_IDinst_N70679),
    .ADR2(DLX_IDinst__n0364),
    .ADR3(N90703),
    .O(DLX_IDinst__n0106[0])
  );
  X_BUF \DLX_IDinst_rt_addr<0>/XUSED  (
    .I(\DLX_IDinst_rt_addr<0>/FROM ),
    .O(N90703)
  );
  defparam DLX_EXinst_Ker633721.INIT = 16'hFC30;
  X_LUT4 DLX_EXinst_Ker633721 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(DLX_IDinst_reg_out_A[16]),
    .ADR3(DLX_IDinst_reg_out_A[14]),
    .O(\DLX_EXinst_N63374/FROM )
  );
  defparam DLX_EXinst_Ker63908_SW0.INIT = 16'hEE22;
  X_LUT4 DLX_EXinst_Ker63908_SW0 (
    .ADR0(DLX_EXinst_N62876),
    .ADR1(DLX_IDinst_reg_out_B[0]),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N63374),
    .O(\DLX_EXinst_N63374/GROM )
  );
  X_BUF \DLX_EXinst_N63374/XUSED  (
    .I(\DLX_EXinst_N63374/FROM ),
    .O(DLX_EXinst_N63374)
  );
  X_BUF \DLX_EXinst_N63374/YUSED  (
    .I(\DLX_EXinst_N63374/GROM ),
    .O(N93487)
  );
  defparam \DLX_IDinst__n0113<4>_SW0 .INIT = 16'hA8FC;
  X_LUT4 \DLX_IDinst__n0113<4>_SW0  (
    .ADR0(DLX_IDinst_IR_latched[27]),
    .ADR1(DLX_IDinst_N69963),
    .ADR2(CHOICE2100),
    .ADR3(DLX_IDinst_N70991),
    .O(\DLX_IDinst_IR_opcode_field<4>/FROM )
  );
  defparam \DLX_IDinst__n0113<4> .INIT = 16'hC080;
  X_LUT4 \DLX_IDinst__n0113<4>  (
    .ADR0(DLX_IDinst__n0364),
    .ADR1(DLX_IDinst_N70679),
    .ADR2(DLX_IDinst_IR_latched[30]),
    .ADR3(N95569),
    .O(DLX_IDinst__n0113[4])
  );
  X_BUF \DLX_IDinst_IR_opcode_field<4>/XUSED  (
    .I(\DLX_IDinst_IR_opcode_field<4>/FROM ),
    .O(N95569)
  );
  defparam DLX_EXinst_Ker632921.INIT = 16'hFACC;
  X_LUT4 DLX_EXinst_Ker632921 (
    .ADR0(CHOICE1132),
    .ADR1(\DLX_EXinst_Mshift__n0028_Sh[24] ),
    .ADR2(CHOICE1126),
    .ADR3(DLX_IDinst_IR_function_field_2_1),
    .O(\DLX_EXinst_N63294/FROM )
  );
  defparam DLX_EXinst_Ker6538912.INIT = 16'h00AC;
  X_LUT4 DLX_EXinst_Ker6538912 (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(DLX_EXinst_N63294),
    .ADR2(DLX_IDinst_IR_function_field_3_1),
    .ADR3(\DLX_IDinst_Imm[5] ),
    .O(\DLX_EXinst_N63294/GROM )
  );
  X_BUF \DLX_EXinst_N63294/XUSED  (
    .I(\DLX_EXinst_N63294/FROM ),
    .O(DLX_EXinst_N63294)
  );
  X_BUF \DLX_EXinst_N63294/YUSED  (
    .I(\DLX_EXinst_N63294/GROM ),
    .O(CHOICE1356)
  );
  defparam DLX_IFinst_NPC_11_1_1152.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_11_1_1152 (
    .I(\NPC_eff<11>/OD ),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\NPC_eff<11>/OFF/RST ),
    .O(DLX_IFinst_NPC_11_1)
  );
  X_OR2 \NPC_eff<11>/OFF/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\NPC_eff<11>/OFF/RST )
  );
  defparam DLX_EXinst_Ker643321.INIT = 16'hFDA8;
  X_LUT4 DLX_EXinst_Ker643321 (
    .ADR0(DLX_IDinst_reg_out_B_3_1),
    .ADR1(CHOICE1138),
    .ADR2(CHOICE1144),
    .ADR3(\DLX_EXinst_Mshift__n0026_Sh[18] ),
    .O(\DLX_EXinst_N64334/FROM )
  );
  defparam \DLX_EXinst__n0006<14>130 .INIT = 16'hA820;
  X_LUT4 \DLX_EXinst__n0006<14>130  (
    .ADR0(DLX_EXinst_N66485),
    .ADR1(DLX_IDinst_reg_out_B[2]),
    .ADR2(DLX_EXinst_N64530),
    .ADR3(DLX_EXinst_N64334),
    .O(\DLX_EXinst_N64334/GROM )
  );
  X_BUF \DLX_EXinst_N64334/XUSED  (
    .I(\DLX_EXinst_N64334/FROM ),
    .O(DLX_EXinst_N64334)
  );
  X_BUF \DLX_EXinst_N64334/YUSED  (
    .I(\DLX_EXinst_N64334/GROM ),
    .O(CHOICE4261)
  );
  defparam DLX_EXinst_Ker634521.INIT = 16'hFC30;
  X_LUT4 DLX_EXinst_Ker634521 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_IR_function_field[1]),
    .ADR2(DLX_IDinst_reg_out_A[16]),
    .ADR3(DLX_IDinst_reg_out_A[14]),
    .O(\DLX_EXinst_N63454/FROM )
  );
  defparam DLX_EXinst_Ker6540910.INIT = 16'hA808;
  X_LUT4 DLX_EXinst_Ker6540910 (
    .ADR0(DLX_IDinst_IR_function_field_3_1),
    .ADR1(DLX_EXinst_N62791),
    .ADR2(DLX_IDinst_IR_function_field[0]),
    .ADR3(DLX_EXinst_N63454),
    .O(\DLX_EXinst_N63454/GROM )
  );
  X_BUF \DLX_EXinst_N63454/XUSED  (
    .I(\DLX_EXinst_N63454/FROM ),
    .O(DLX_EXinst_N63454)
  );
  X_BUF \DLX_EXinst_N63454/YUSED  (
    .I(\DLX_EXinst_N63454/GROM ),
    .O(CHOICE1282)
  );
  defparam DLX_EXinst_Ker640921.INIT = 16'hEE22;
  X_LUT4 DLX_EXinst_Ker640921 (
    .ADR0(\DLX_EXinst_Mshift__n0025_Sh[21] ),
    .ADR1(DLX_IDinst_reg_out_B[3]),
    .ADR2(VCC),
    .ADR3(\DLX_EXinst_Mshift__n0025_Sh[13] ),
    .O(\DLX_EXinst_N64094/FROM )
  );
  defparam \DLX_EXinst__n0006<25>172 .INIT = 16'h5404;
  X_LUT4 \DLX_EXinst__n0006<25>172  (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(N97089),
    .ADR2(DLX_IDinst_reg_out_B[2]),
    .ADR3(DLX_EXinst_N64094),
    .O(\DLX_EXinst_N64094/GROM )
  );
  X_BUF \DLX_EXinst_N64094/XUSED  (
    .I(\DLX_EXinst_N64094/FROM ),
    .O(DLX_EXinst_N64094)
  );
  X_BUF \DLX_EXinst_N64094/YUSED  (
    .I(\DLX_EXinst_N64094/GROM ),
    .O(CHOICE4780)
  );
  defparam \DLX_EXinst__n0006<1>117_SW0 .INIT = 16'h0505;
  X_LUT4 \DLX_EXinst__n0006<1>117_SW0  (
    .ADR0(DLX_IDinst_reg_out_A[1]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_IR_opcode_field[0]),
    .ADR3(VCC),
    .O(\N127314/FROM )
  );
  defparam \DLX_EXinst__n0006<6>16_SW0 .INIT = 16'h0505;
  X_LUT4 \DLX_EXinst__n0006<6>16_SW0  (
    .ADR0(DLX_IDinst_IR_opcode_field[0]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[6]),
    .ADR3(VCC),
    .O(\N127314/GROM )
  );
  X_BUF \N127314/XUSED  (
    .I(\N127314/FROM ),
    .O(N127314)
  );
  X_BUF \N127314/YUSED  (
    .I(\N127314/GROM ),
    .O(N127286)
  );
  defparam DM_delay_inst_wint181.INIT = 16'h3333;
  X_LUT4 DM_delay_inst_wint181 (
    .ADR0(VCC),
    .ADR1(DM_delay_inst_wint17),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DM_delay_inst_wint18/GROM )
  );
  X_BUF \DM_delay_inst_wint18/YUSED  (
    .I(\DM_delay_inst_wint18/GROM ),
    .O(DM_delay_inst_wint18)
  );
  defparam DM_delay_inst_wint261.INIT = 16'h5555;
  X_LUT4 DM_delay_inst_wint261 (
    .ADR0(DM_delay_inst_wint25),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DM_delay_inst_wint26/FROM )
  );
  defparam DM_delay_inst_wint271.INIT = 16'h00FF;
  X_LUT4 DM_delay_inst_wint271 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DM_delay_inst_wint26),
    .O(\DM_delay_inst_wint26/GROM )
  );
  X_BUF \DM_delay_inst_wint26/XUSED  (
    .I(\DM_delay_inst_wint26/FROM ),
    .O(DM_delay_inst_wint26)
  );
  X_BUF \DM_delay_inst_wint26/YUSED  (
    .I(\DM_delay_inst_wint26/GROM ),
    .O(DM_delay_inst_wint27)
  );
  defparam DM_delay_inst_wint341.INIT = 16'h00FF;
  X_LUT4 DM_delay_inst_wint341 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DM_delay_inst_wint33),
    .O(\DM_delay_inst_wint34/FROM )
  );
  defparam DM_delay_inst_wint351.INIT = 16'h00FF;
  X_LUT4 DM_delay_inst_wint351 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DM_delay_inst_wint34),
    .O(\DM_delay_inst_wint34/GROM )
  );
  X_BUF \DM_delay_inst_wint34/XUSED  (
    .I(\DM_delay_inst_wint34/FROM ),
    .O(DM_delay_inst_wint34)
  );
  X_BUF \DM_delay_inst_wint34/YUSED  (
    .I(\DM_delay_inst_wint34/GROM ),
    .O(DM_delay_inst_wint35)
  );
  defparam \DLX_EXinst__n0006<0>36 .INIT = 16'h2320;
  X_LUT4 \DLX_EXinst__n0006<0>36  (
    .ADR0(DLX_EXinst_N64864),
    .ADR1(DLX_IDinst_reg_out_B[3]),
    .ADR2(DLX_IDinst_reg_out_B[0]),
    .ADR3(N126134),
    .O(\CHOICE5864/FROM )
  );
  defparam \DLX_EXinst__n0006<0>59 .INIT = 16'h3320;
  X_LUT4 \DLX_EXinst__n0006<0>59  (
    .ADR0(DLX_IDinst_reg_out_B[3]),
    .ADR1(DLX_IDinst_reg_out_B[2]),
    .ADR2(\DLX_EXinst_Mshift__n0023_Sh[8] ),
    .ADR3(CHOICE5864),
    .O(\CHOICE5864/GROM )
  );
  X_BUF \CHOICE5864/XUSED  (
    .I(\CHOICE5864/FROM ),
    .O(CHOICE5864)
  );
  X_BUF \CHOICE5864/YUSED  (
    .I(\CHOICE5864/GROM ),
    .O(CHOICE5866)
  );
  defparam \DLX_IDinst_regB_eff<7>1 .INIT = 16'hEAC0;
  X_LUT4 \DLX_IDinst_regB_eff<7>1  (
    .ADR0(DLX_RF_data_in[7]),
    .ADR1(DLX_IDinst_N70716),
    .ADR2(DLX_IDinst_reg_out_B_RF[7]),
    .ADR3(DLX_IDinst__n0145),
    .O(\DLX_IDinst_regB_eff<7>/FROM )
  );
  defparam \DLX_IDinst_regB_eff<14>1 .INIT = 16'hECA0;
  X_LUT4 \DLX_IDinst_regB_eff<14>1  (
    .ADR0(DLX_IDinst_N70716),
    .ADR1(DLX_IDinst__n0145),
    .ADR2(DLX_IDinst_reg_out_B_RF[14]),
    .ADR3(DLX_MEMinst_RF_data_in[14]),
    .O(\DLX_IDinst_regB_eff<7>/GROM )
  );
  X_BUF \DLX_IDinst_regB_eff<7>/XUSED  (
    .I(\DLX_IDinst_regB_eff<7>/FROM ),
    .O(DLX_IDinst_regB_eff[7])
  );
  X_BUF \DLX_IDinst_regB_eff<7>/YUSED  (
    .I(\DLX_IDinst_regB_eff<7>/GROM ),
    .O(DLX_IDinst_regB_eff[14])
  );
  defparam \DLX_IDinst_regB_eff<8>1 .INIT = 16'hEAC0;
  X_LUT4 \DLX_IDinst_regB_eff<8>1  (
    .ADR0(DLX_IDinst_N70716),
    .ADR1(DLX_IDinst__n0145),
    .ADR2(DLX_MEMinst_RF_data_in[8]),
    .ADR3(DLX_IDinst_reg_out_B_RF[8]),
    .O(\DLX_IDinst_regB_eff<8>/FROM )
  );
  defparam \DLX_IDinst_regB_eff<22>1 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst_regB_eff<22>1  (
    .ADR0(DLX_IDinst_reg_out_B_RF[22]),
    .ADR1(DLX_IDinst_N70716),
    .ADR2(DLX_MEMinst_RF_data_in[22]),
    .ADR3(DLX_IDinst__n0145),
    .O(\DLX_IDinst_regB_eff<8>/GROM )
  );
  X_BUF \DLX_IDinst_regB_eff<8>/XUSED  (
    .I(\DLX_IDinst_regB_eff<8>/FROM ),
    .O(DLX_IDinst_regB_eff[8])
  );
  X_BUF \DLX_IDinst_regB_eff<8>/YUSED  (
    .I(\DLX_IDinst_regB_eff<8>/GROM ),
    .O(DLX_IDinst_regB_eff[22])
  );
  defparam \DLX_IDinst_regB_eff<9>1 .INIT = 16'hECA0;
  X_LUT4 \DLX_IDinst_regB_eff<9>1  (
    .ADR0(DLX_IDinst_reg_out_B_RF[9]),
    .ADR1(DLX_IDinst__n0145),
    .ADR2(DLX_IDinst_N70716),
    .ADR3(DLX_MEMinst_RF_data_in[9]),
    .O(\DLX_IDinst_regB_eff<9>/FROM )
  );
  defparam \DLX_IDinst_regB_eff<30>1 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst_regB_eff<30>1  (
    .ADR0(DLX_MEMinst_RF_data_in[30]),
    .ADR1(DLX_IDinst__n0145),
    .ADR2(DLX_IDinst_N70716),
    .ADR3(DLX_IDinst_reg_out_B_RF[30]),
    .O(\DLX_IDinst_regB_eff<9>/GROM )
  );
  X_BUF \DLX_IDinst_regB_eff<9>/XUSED  (
    .I(\DLX_IDinst_regB_eff<9>/FROM ),
    .O(DLX_IDinst_regB_eff[9])
  );
  X_BUF \DLX_IDinst_regB_eff<9>/YUSED  (
    .I(\DLX_IDinst_regB_eff<9>/GROM ),
    .O(DLX_IDinst_regB_eff[30])
  );
  defparam DLX_IFlc_md_mda8_a1.INIT = 16'h2222;
  X_LUT4 DLX_IFlc_md_mda8_a1 (
    .ADR0(DLX_IFlc_md_wint7),
    .ADR1(DLX_IFlc_pd_wint1),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IFlc_md_wint8/FROM )
  );
  defparam DLX_IFlc_md_mda1_a1.INIT = 16'h0F00;
  X_LUT4 DLX_IFlc_md_mda1_a1 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IFlc_pd_wint1),
    .ADR3(DLX_IFlc_ridp3),
    .O(\DLX_IFlc_md_wint8/GROM )
  );
  X_BUF \DLX_IFlc_md_wint8/XUSED  (
    .I(\DLX_IFlc_md_wint8/FROM ),
    .O(DLX_IFlc_md_wint8)
  );
  X_BUF \DLX_IFlc_md_wint8/YUSED  (
    .I(\DLX_IFlc_md_wint8/GROM ),
    .O(DLX_IFlc_md_wint1)
  );
  defparam DLX_EXinst_Ker626291.INIT = 16'h5D0C;
  X_LUT4 DLX_EXinst_Ker626291 (
    .ADR0(DLX_IDinst_reg_out_B[5]),
    .ADR1(DLX_EXinst__n0049),
    .ADR2(N110935),
    .ADR3(N111221),
    .O(\DLX_EXinst_N62631/FROM )
  );
  defparam \DLX_EXinst__n0006<4>177 .INIT = 16'hE200;
  X_LUT4 \DLX_EXinst__n0006<4>177  (
    .ADR0(N96153),
    .ADR1(DLX_IDinst_reg_out_B[2]),
    .ADR2(DLX_EXinst_N64804),
    .ADR3(DLX_EXinst_N62631),
    .O(\DLX_EXinst_N62631/GROM )
  );
  X_BUF \DLX_EXinst_N62631/XUSED  (
    .I(\DLX_EXinst_N62631/FROM ),
    .O(DLX_EXinst_N62631)
  );
  X_BUF \DLX_EXinst_N62631/YUSED  (
    .I(\DLX_EXinst_N62631/GROM ),
    .O(CHOICE4016)
  );
  defparam \DLX_EXinst_Mshift__n0027_Sh<6>_SW0 .INIT = 16'hCACA;
  X_LUT4 \DLX_EXinst_Mshift__n0027_Sh<6>_SW0  (
    .ADR0(DLX_IDinst_reg_out_A[5]),
    .ADR1(DLX_IDinst_reg_out_A[3]),
    .ADR2(DLX_IDinst_IR_function_field_1_1),
    .ADR3(VCC),
    .O(\N94155/FROM )
  );
  defparam DLX_EXinst_Ker651331.INIT = 16'hCFC0;
  X_LUT4 DLX_EXinst_Ker651331 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[3]),
    .ADR2(DLX_IDinst_IR_function_field_1_1),
    .ADR3(DLX_IDinst_reg_out_A[1]),
    .O(\N94155/GROM )
  );
  X_BUF \N94155/XUSED  (
    .I(\N94155/FROM ),
    .O(N94155)
  );
  X_BUF \N94155/YUSED  (
    .I(\N94155/GROM ),
    .O(DLX_EXinst_N65135)
  );
  defparam DLX_EXinst_Ker633571.INIT = 16'hEE22;
  X_LUT4 DLX_EXinst_Ker633571 (
    .ADR0(DLX_IDinst_reg_out_A[10]),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[8]),
    .O(\DLX_EXinst_N63359/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0025_Sh<11>1 .INIT = 16'hFA0A;
  X_LUT4 \DLX_EXinst_Mshift__n0025_Sh<11>1  (
    .ADR0(DLX_EXinst_N62861),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[0]),
    .ADR3(DLX_EXinst_N63359),
    .O(\DLX_EXinst_N63359/GROM )
  );
  X_BUF \DLX_EXinst_N63359/XUSED  (
    .I(\DLX_EXinst_N63359/FROM ),
    .O(DLX_EXinst_N63359)
  );
  X_BUF \DLX_EXinst_N63359/YUSED  (
    .I(\DLX_EXinst_N63359/GROM ),
    .O(\DLX_EXinst_Mshift__n0025_Sh[11] )
  );
  defparam DLX_EXinst_Ker634721.INIT = 16'hFC0C;
  X_LUT4 DLX_EXinst_Ker634721 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[24]),
    .ADR2(DLX_IDinst_IR_function_field[1]),
    .ADR3(DLX_IDinst_reg_out_A[22]),
    .O(\DLX_EXinst_N63474/FROM )
  );
  defparam DLX_EXinst_Ker635171.INIT = 16'hF5A0;
  X_LUT4 DLX_EXinst_Ker635171 (
    .ADR0(DLX_IDinst_IR_function_field_1_1),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[24]),
    .ADR3(DLX_IDinst_reg_out_A[22]),
    .O(\DLX_EXinst_N63474/GROM )
  );
  X_BUF \DLX_EXinst_N63474/XUSED  (
    .I(\DLX_EXinst_N63474/FROM ),
    .O(DLX_EXinst_N63474)
  );
  X_BUF \DLX_EXinst_N63474/YUSED  (
    .I(\DLX_EXinst_N63474/GROM ),
    .O(DLX_EXinst_N63519)
  );
  defparam DLX_EXinst_Ker643171.INIT = 16'hEE22;
  X_LUT4 DLX_EXinst_Ker643171 (
    .ADR0(\DLX_EXinst_Mshift__n0026_Sh[16] ),
    .ADR1(DLX_IDinst_reg_out_B_3_1),
    .ADR2(VCC),
    .ADR3(\DLX_EXinst_Mshift__n0026_Sh[24] ),
    .O(\DLX_EXinst_N64319/FROM )
  );
  defparam \DLX_EXinst__n0006<12>130 .INIT = 16'hA820;
  X_LUT4 \DLX_EXinst__n0006<12>130  (
    .ADR0(DLX_EXinst_N66485),
    .ADR1(DLX_IDinst_reg_out_B[2]),
    .ADR2(N97375),
    .ADR3(DLX_EXinst_N64319),
    .O(\DLX_EXinst_N64319/GROM )
  );
  X_BUF \DLX_EXinst_N64319/XUSED  (
    .I(\DLX_EXinst_N64319/FROM ),
    .O(DLX_EXinst_N64319)
  );
  X_BUF \DLX_EXinst_N64319/YUSED  (
    .I(\DLX_EXinst_N64319/GROM ),
    .O(CHOICE3889)
  );
  defparam DLX_IFinst_NPC_12_1_1153.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_12_1_1153 (
    .I(\NPC_eff<12>/OD ),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\NPC_eff<12>/OFF/RST ),
    .O(DLX_IFinst_NPC_12_1)
  );
  X_OR2 \NPC_eff<12>/OFF/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\NPC_eff<12>/OFF/RST )
  );
  defparam \DLX_EXinst_Mshift__n0025_Sh<7>_SW0 .INIT = 16'hF5A0;
  X_LUT4 \DLX_EXinst_Mshift__n0025_Sh<7>_SW0  (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[4]),
    .ADR3(DLX_IDinst_reg_out_A[6]),
    .O(\N94305/FROM )
  );
  defparam DLX_EXinst_Ker642531.INIT = 16'hAFA0;
  X_LUT4 DLX_EXinst_Ker642531 (
    .ADR0(DLX_IDinst_reg_out_A[4]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[1]),
    .ADR3(DLX_IDinst_reg_out_A[2]),
    .O(\N94305/GROM )
  );
  X_BUF \N94305/XUSED  (
    .I(\N94305/FROM ),
    .O(N94305)
  );
  X_BUF \N94305/YUSED  (
    .I(\N94305/GROM ),
    .O(DLX_EXinst_N64255)
  );
  defparam DLX_EXinst_Ker634371.INIT = 16'hF0CC;
  X_LUT4 DLX_EXinst_Ker634371 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[10]),
    .ADR2(DLX_IDinst_reg_out_A[8]),
    .ADR3(DLX_IDinst_IR_function_field[1]),
    .O(\DLX_EXinst_N63439/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0027_Sh<11>1 .INIT = 16'hEE22;
  X_LUT4 \DLX_EXinst_Mshift__n0027_Sh<11>1  (
    .ADR0(DLX_EXinst_N62776),
    .ADR1(DLX_IDinst_IR_function_field_0_1),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N63439),
    .O(\DLX_EXinst_N63439/GROM )
  );
  X_BUF \DLX_EXinst_N63439/XUSED  (
    .I(\DLX_EXinst_N63439/FROM ),
    .O(DLX_EXinst_N63439)
  );
  X_BUF \DLX_EXinst_N63439/YUSED  (
    .I(\DLX_EXinst_N63439/GROM ),
    .O(\DLX_EXinst_Mshift__n0027_Sh[11] )
  );
  defparam Ker57310.INIT = 16'h0001;
  X_LUT4 Ker57310 (
    .ADR0(vga_select_6[0]),
    .ADR1(N95202),
    .ADR2(vga_select_6[2]),
    .ADR3(vga_select_6[1]),
    .O(\N57312/FROM )
  );
  defparam \DM_read_data<30>1 .INIT = 16'hFFC0;
  X_LUT4 \DM_read_data<30>1  (
    .ADR0(VCC),
    .ADR1(vga_select_6[0]),
    .ADR2(RAM_read_data[30]),
    .ADR3(N57312),
    .O(\N57312/GROM )
  );
  X_BUF \N57312/XUSED  (
    .I(\N57312/FROM ),
    .O(N57312)
  );
  X_BUF \N57312/YUSED  (
    .I(\N57312/GROM ),
    .O(DM_read_data[30])
  );
  defparam DLX_IFlc_md_mda7_a1.INIT = 16'h4444;
  X_LUT4 DLX_IFlc_md_mda7_a1 (
    .ADR0(DLX_IFlc_pd_wint1),
    .ADR1(DLX_IFlc_md_wint6),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IFlc_md_wint7/FROM )
  );
  defparam DLX_IFlc_md_mda36_a1.INIT = 16'h3300;
  X_LUT4 DLX_IFlc_md_mda36_a1 (
    .ADR0(VCC),
    .ADR1(DLX_IFlc_pd_wint1),
    .ADR2(VCC),
    .ADR3(DLX_IFlc_md_wint35),
    .O(\DLX_IFlc_md_wint7/GROM )
  );
  X_BUF \DLX_IFlc_md_wint7/XUSED  (
    .I(\DLX_IFlc_md_wint7/FROM ),
    .O(DLX_IFlc_md_wint7)
  );
  X_BUF \DLX_IFlc_md_wint7/YUSED  (
    .I(\DLX_IFlc_md_wint7/GROM ),
    .O(DLX_IFlc_md_wint36)
  );
  defparam DM_delay_inst_wint191.INIT = 16'h00FF;
  X_LUT4 DM_delay_inst_wint191 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DM_delay_inst_wint18),
    .O(\DM_delay_inst_wint19/GROM )
  );
  X_BUF \DM_delay_inst_wint19/YUSED  (
    .I(\DM_delay_inst_wint19/GROM ),
    .O(DM_delay_inst_wint19)
  );
  defparam DLX_EXinst_Ker661101.INIT = 16'h0008;
  X_LUT4 DLX_EXinst_Ker661101 (
    .ADR0(DLX_IDinst_IR_opcode_field[4]),
    .ADR1(DLX_IDinst_IR_opcode_field[2]),
    .ADR2(DLX_IDinst_IR_opcode_field[3]),
    .ADR3(DLX_IDinst_IR_opcode_field[5]),
    .O(\DLX_EXinst_N66112/FROM )
  );
  defparam DLX_EXinst_Ker665051.INIT = 16'h1000;
  X_LUT4 DLX_EXinst_Ker665051 (
    .ADR0(N109130),
    .ADR1(DLX_IDinst_IR_opcode_field[0]),
    .ADR2(DLX_IDinst_IR_opcode_field[1]),
    .ADR3(DLX_EXinst_N66112),
    .O(\DLX_EXinst_N66112/GROM )
  );
  X_BUF \DLX_EXinst_N66112/XUSED  (
    .I(\DLX_EXinst_N66112/FROM ),
    .O(DLX_EXinst_N66112)
  );
  X_BUF \DLX_EXinst_N66112/YUSED  (
    .I(\DLX_EXinst_N66112/GROM ),
    .O(DLX_EXinst_N66507)
  );
  defparam DLX_EXinst_Ker633821.INIT = 16'hFC30;
  X_LUT4 DLX_EXinst_Ker633821 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(DLX_IDinst_reg_out_A[20]),
    .ADR3(DLX_IDinst_reg_out_A[18]),
    .O(\DLX_EXinst_N63384/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0025_Sh<21>1 .INIT = 16'hFC0C;
  X_LUT4 \DLX_EXinst_Mshift__n0025_Sh<21>1  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N62886),
    .ADR2(DLX_IDinst_reg_out_B[0]),
    .ADR3(DLX_EXinst_N63384),
    .O(\DLX_EXinst_N63384/GROM )
  );
  X_BUF \DLX_EXinst_N63384/XUSED  (
    .I(\DLX_EXinst_N63384/FROM ),
    .O(DLX_EXinst_N63384)
  );
  X_BUF \DLX_EXinst_N63384/YUSED  (
    .I(\DLX_EXinst_N63384/GROM ),
    .O(\DLX_EXinst_Mshift__n0025_Sh[21] )
  );
  defparam DLX_EXinst_Ker634621.INIT = 16'hCFC0;
  X_LUT4 DLX_EXinst_Ker634621 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[18]),
    .ADR2(DLX_IDinst_IR_function_field[1]),
    .ADR3(DLX_IDinst_reg_out_A[20]),
    .O(\DLX_EXinst_N63464/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0027_Sh<21>1 .INIT = 16'hEE44;
  X_LUT4 \DLX_EXinst_Mshift__n0027_Sh<21>1  (
    .ADR0(DLX_IDinst_IR_function_field_0_1),
    .ADR1(DLX_EXinst_N62801),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N63464),
    .O(\DLX_EXinst_N63464/GROM )
  );
  X_BUF \DLX_EXinst_N63464/XUSED  (
    .I(\DLX_EXinst_N63464/FROM ),
    .O(DLX_EXinst_N63464)
  );
  X_BUF \DLX_EXinst_N63464/YUSED  (
    .I(\DLX_EXinst_N63464/GROM ),
    .O(\DLX_EXinst_Mshift__n0027_Sh[21] )
  );
  defparam DM_delay_inst_wint281.INIT = 16'h3333;
  X_LUT4 DM_delay_inst_wint281 (
    .ADR0(VCC),
    .ADR1(DM_delay_inst_wint27),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DM_delay_inst_wint28/GROM )
  );
  X_BUF \DM_delay_inst_wint28/YUSED  (
    .I(\DM_delay_inst_wint28/GROM ),
    .O(DM_delay_inst_wint28)
  );
  defparam DM_delay_inst_wint361.INIT = 16'h00FF;
  X_LUT4 DM_delay_inst_wint361 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DM_delay_inst_wint35),
    .O(\DM_delay_inst_wint36/GROM )
  );
  X_BUF \DM_delay_inst_wint36/YUSED  (
    .I(\DM_delay_inst_wint36/GROM ),
    .O(DM_delay_inst_wint36)
  );
  defparam reset_IBUF_1_1154.INIT = 16'hAAAA;
  X_LUT4 reset_IBUF_1_1154 (
    .ADR0(reset_IBUF),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\reset_IBUF_1/FROM )
  );
  defparam \vga_top_vga1_greenout<1>1 .INIT = 16'h000C;
  X_LUT4 \vga_top_vga1_greenout<1>1  (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_videoon),
    .ADR2(vram_out_vga_eff),
    .ADR3(reset_IBUF_1),
    .O(\reset_IBUF_1/GROM )
  );
  X_BUF \reset_IBUF_1/XUSED  (
    .I(\reset_IBUF_1/FROM ),
    .O(reset_IBUF_1)
  );
  X_BUF \reset_IBUF_1/YUSED  (
    .I(\reset_IBUF_1/GROM ),
    .O(green_1_OBUF)
  );
  defparam \DLX_IDinst_regB_eff<16>1 .INIT = 16'hECA0;
  X_LUT4 \DLX_IDinst_regB_eff<16>1  (
    .ADR0(DLX_IDinst__n0145),
    .ADR1(DLX_IDinst_N70716),
    .ADR2(DLX_MEMinst_RF_data_in[16]),
    .ADR3(DLX_IDinst_reg_out_B_RF[16]),
    .O(\DLX_IDinst_regB_eff<16>/FROM )
  );
  defparam \DLX_IDinst_regB_eff<15>1 .INIT = 16'hEAC0;
  X_LUT4 \DLX_IDinst_regB_eff<15>1  (
    .ADR0(DLX_IDinst_reg_out_B_RF[15]),
    .ADR1(DLX_IDinst__n0145),
    .ADR2(DLX_MEMinst_RF_data_in[15]),
    .ADR3(DLX_IDinst_N70716),
    .O(\DLX_IDinst_regB_eff<16>/GROM )
  );
  X_BUF \DLX_IDinst_regB_eff<16>/XUSED  (
    .I(\DLX_IDinst_regB_eff<16>/FROM ),
    .O(DLX_IDinst_regB_eff[16])
  );
  X_BUF \DLX_IDinst_regB_eff<16>/YUSED  (
    .I(\DLX_IDinst_regB_eff<16>/GROM ),
    .O(DLX_IDinst_regB_eff[15])
  );
  defparam \DLX_IDinst_regB_eff<17>1 .INIT = 16'hECA0;
  X_LUT4 \DLX_IDinst_regB_eff<17>1  (
    .ADR0(DLX_IDinst__n0145),
    .ADR1(DLX_IDinst_N70716),
    .ADR2(DLX_MEMinst_RF_data_in[17]),
    .ADR3(DLX_IDinst_reg_out_B_RF[17]),
    .O(\DLX_IDinst_regB_eff<17>/FROM )
  );
  defparam \DLX_IDinst_regB_eff<23>1 .INIT = 16'hEAC0;
  X_LUT4 \DLX_IDinst_regB_eff<23>1  (
    .ADR0(DLX_IDinst__n0145),
    .ADR1(DLX_IDinst_reg_out_B_RF[23]),
    .ADR2(DLX_IDinst_N70716),
    .ADR3(DLX_MEMinst_RF_data_in[23]),
    .O(\DLX_IDinst_regB_eff<17>/GROM )
  );
  X_BUF \DLX_IDinst_regB_eff<17>/XUSED  (
    .I(\DLX_IDinst_regB_eff<17>/FROM ),
    .O(DLX_IDinst_regB_eff[17])
  );
  X_BUF \DLX_IDinst_regB_eff<17>/YUSED  (
    .I(\DLX_IDinst_regB_eff<17>/GROM ),
    .O(DLX_IDinst_regB_eff[23])
  );
  defparam \DLX_IDinst_regB_eff<18>1 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst_regB_eff<18>1  (
    .ADR0(DLX_IDinst_N70716),
    .ADR1(DLX_IDinst_reg_out_B_RF[18]),
    .ADR2(DLX_IDinst__n0145),
    .ADR3(DLX_MEMinst_RF_data_in[18]),
    .O(\DLX_IDinst_regB_eff<18>/FROM )
  );
  defparam \DLX_IDinst_regB_eff<31>1 .INIT = 16'hEAC0;
  X_LUT4 \DLX_IDinst_regB_eff<31>1  (
    .ADR0(DLX_IDinst__n0145),
    .ADR1(DLX_IDinst_reg_out_B_RF[31]),
    .ADR2(DLX_IDinst_N70716),
    .ADR3(DLX_MEMinst_RF_data_in[31]),
    .O(\DLX_IDinst_regB_eff<18>/GROM )
  );
  X_BUF \DLX_IDinst_regB_eff<18>/XUSED  (
    .I(\DLX_IDinst_regB_eff<18>/FROM ),
    .O(DLX_IDinst_regB_eff[18])
  );
  X_BUF \DLX_IDinst_regB_eff<18>/YUSED  (
    .I(\DLX_IDinst_regB_eff<18>/GROM ),
    .O(DLX_IDinst_regB_eff[31])
  );
  defparam DLX_EXinst_Ker633671.INIT = 16'hFC0C;
  X_LUT4 DLX_EXinst_Ker633671 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[14]),
    .ADR2(DLX_IDinst_reg_out_B[1]),
    .ADR3(DLX_IDinst_reg_out_A[12]),
    .O(\DLX_EXinst_N63369/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0025_Sh<15>1 .INIT = 16'hEE44;
  X_LUT4 \DLX_EXinst_Mshift__n0025_Sh<15>1  (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(DLX_EXinst_N62871),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N63369),
    .O(\DLX_EXinst_N63369/GROM )
  );
  X_BUF \DLX_EXinst_N63369/XUSED  (
    .I(\DLX_EXinst_N63369/FROM ),
    .O(DLX_EXinst_N63369)
  );
  X_BUF \DLX_EXinst_N63369/YUSED  (
    .I(\DLX_EXinst_N63369/GROM ),
    .O(\DLX_EXinst_Mshift__n0025_Sh[15] )
  );
  defparam DLX_EXinst_Ker661031.INIT = 16'h0008;
  X_LUT4 DLX_EXinst_Ker661031 (
    .ADR0(DLX_IDinst_IR_opcode_field[3]),
    .ADR1(DLX_IDinst_IR_opcode_field[2]),
    .ADR2(DLX_IDinst_IR_opcode_field[5]),
    .ADR3(DLX_IDinst_IR_opcode_field[4]),
    .O(\DLX_EXinst_N66105/FROM )
  );
  defparam DLX_EXinst__n00801.INIT = 16'h2200;
  X_LUT4 DLX_EXinst__n00801 (
    .ADR0(DLX_IDinst_IR_opcode_field[1]),
    .ADR1(DLX_IDinst_IR_opcode_field[0]),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N66105),
    .O(\DLX_EXinst_N66105/GROM )
  );
  X_BUF \DLX_EXinst_N66105/XUSED  (
    .I(\DLX_EXinst_N66105/FROM ),
    .O(DLX_EXinst_N66105)
  );
  X_BUF \DLX_EXinst_N66105/YUSED  (
    .I(\DLX_EXinst_N66105/GROM ),
    .O(DLX_EXinst__n0080)
  );
  defparam DLX_EXinst_Ker627191.INIT = 16'hF3C0;
  X_LUT4 DLX_EXinst_Ker627191 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_B[0]),
    .ADR2(DLX_IDinst_reg_out_A[30]),
    .ADR3(DLX_IDinst_reg_out_A[29]),
    .O(\DLX_EXinst_N62721/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0026_Sh<29>1 .INIT = 16'h2F20;
  X_LUT4 \DLX_EXinst_Mshift__n0026_Sh<29>1  (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(DLX_IDinst_reg_out_B[0]),
    .ADR2(DLX_IDinst_reg_out_B[1]),
    .ADR3(DLX_EXinst_N62721),
    .O(\DLX_EXinst_N62721/GROM )
  );
  X_BUF \DLX_EXinst_N62721/XUSED  (
    .I(\DLX_EXinst_N62721/FROM ),
    .O(DLX_EXinst_N62721)
  );
  X_BUF \DLX_EXinst_N62721/YUSED  (
    .I(\DLX_EXinst_N62721/GROM ),
    .O(\DLX_EXinst_Mshift__n0026_Sh[29] )
  );
  defparam DLX_IFinst_NPC_13_1_1155.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_13_1_1155 (
    .I(\NPC_eff<13>/OD ),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\NPC_eff<13>/OFF/RST ),
    .O(DLX_IFinst_NPC_13_1)
  );
  X_OR2 \NPC_eff<13>/OFF/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\NPC_eff<13>/OFF/RST )
  );
  defparam DLX_EXinst_Ker634471.INIT = 16'hFA0A;
  X_LUT4 DLX_EXinst_Ker634471 (
    .ADR0(DLX_IDinst_reg_out_A[14]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_IR_function_field[1]),
    .ADR3(DLX_IDinst_reg_out_A[12]),
    .O(\DLX_EXinst_N63449/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0027_Sh<15>1 .INIT = 16'hFA0A;
  X_LUT4 \DLX_EXinst_Mshift__n0027_Sh<15>1  (
    .ADR0(DLX_EXinst_N62786),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_IR_function_field_0_1),
    .ADR3(DLX_EXinst_N63449),
    .O(\DLX_EXinst_N63449/GROM )
  );
  X_BUF \DLX_EXinst_N63449/XUSED  (
    .I(\DLX_EXinst_N63449/FROM ),
    .O(DLX_EXinst_N63449)
  );
  X_BUF \DLX_EXinst_N63449/YUSED  (
    .I(\DLX_EXinst_N63449/GROM ),
    .O(\DLX_EXinst_Mshift__n0027_Sh[15] )
  );
  defparam DLX_EXinst_Ker643271.INIT = 16'hEEE4;
  X_LUT4 DLX_EXinst_Ker643271 (
    .ADR0(DLX_IDinst_reg_out_B_3_1),
    .ADR1(\DLX_EXinst_Mshift__n0026_Sh[17] ),
    .ADR2(CHOICE1312),
    .ADR3(CHOICE1306),
    .O(\DLX_EXinst_N64329/FROM )
  );
  defparam \DLX_EXinst__n0006<13>130 .INIT = 16'hE040;
  X_LUT4 \DLX_EXinst__n0006<13>130  (
    .ADR0(DLX_IDinst_reg_out_B[2]),
    .ADR1(DLX_EXinst_N64545),
    .ADR2(DLX_EXinst_N66485),
    .ADR3(DLX_EXinst_N64329),
    .O(\DLX_EXinst_N64329/GROM )
  );
  X_BUF \DLX_EXinst_N64329/XUSED  (
    .I(\DLX_EXinst_N64329/FROM ),
    .O(DLX_EXinst_N64329)
  );
  X_BUF \DLX_EXinst_N64329/YUSED  (
    .I(\DLX_EXinst_N64329/GROM ),
    .O(CHOICE4321)
  );
  defparam reset_IBUF_2_1156.INIT = 16'hFF00;
  X_LUT4 reset_IBUF_2_1156 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(reset_IBUF),
    .O(\reset_IBUF_2/GROM )
  );
  X_BUF \reset_IBUF_2/YUSED  (
    .I(\reset_IBUF_2/GROM ),
    .O(reset_IBUF_2)
  );
  defparam \DLX_EXinst__n0006<18>9 .INIT = 16'h8C88;
  X_LUT4 \DLX_EXinst__n0006<18>9  (
    .ADR0(DLX_EXinst__n0079),
    .ADR1(DLX_IDinst_reg_out_A[18]),
    .ADR2(\DLX_IDinst_Imm[31] ),
    .ADR3(DLX_EXinst__n0080),
    .O(\CHOICE5408/FROM )
  );
  defparam \DLX_EXinst__n0006<25>9 .INIT = 16'h88C8;
  X_LUT4 \DLX_EXinst__n0006<25>9  (
    .ADR0(DLX_EXinst__n0079),
    .ADR1(DLX_IDinst_reg_out_A[25]),
    .ADR2(DLX_EXinst__n0080),
    .ADR3(\DLX_IDinst_Imm[31] ),
    .O(\CHOICE5408/GROM )
  );
  X_BUF \CHOICE5408/XUSED  (
    .I(\CHOICE5408/FROM ),
    .O(CHOICE5408)
  );
  X_BUF \CHOICE5408/YUSED  (
    .I(\CHOICE5408/GROM ),
    .O(CHOICE4740)
  );
  defparam \DLX_EXinst__n0006<26>9 .INIT = 16'hAA08;
  X_LUT4 \DLX_EXinst__n0006<26>9  (
    .ADR0(DLX_IDinst_reg_out_A[26]),
    .ADR1(DLX_EXinst__n0080),
    .ADR2(\DLX_IDinst_Imm[31] ),
    .ADR3(DLX_EXinst__n0079),
    .O(\CHOICE4675/FROM )
  );
  defparam \DLX_EXinst__n0006<17>9 .INIT = 16'hB0A0;
  X_LUT4 \DLX_EXinst__n0006<17>9  (
    .ADR0(DLX_EXinst__n0079),
    .ADR1(\DLX_IDinst_Imm[31] ),
    .ADR2(DLX_IDinst_reg_out_A[17]),
    .ADR3(DLX_EXinst__n0080),
    .O(\CHOICE4675/GROM )
  );
  X_BUF \CHOICE4675/XUSED  (
    .I(\CHOICE4675/FROM ),
    .O(CHOICE4675)
  );
  X_BUF \CHOICE4675/YUSED  (
    .I(\CHOICE4675/GROM ),
    .O(CHOICE5574)
  );
  defparam DM_delay_inst_wint291.INIT = 16'h3333;
  X_LUT4 DM_delay_inst_wint291 (
    .ADR0(VCC),
    .ADR1(DM_delay_inst_wint28),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DM_delay_inst_wint29/GROM )
  );
  X_BUF \DM_delay_inst_wint29/YUSED  (
    .I(\DM_delay_inst_wint29/GROM ),
    .O(DM_delay_inst_wint29)
  );
  defparam DM_delay_inst_wint371.INIT = 16'h3333;
  X_LUT4 DM_delay_inst_wint371 (
    .ADR0(VCC),
    .ADR1(DM_delay_inst_wint36),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DM_delay_inst_wint37/GROM )
  );
  X_BUF \DM_delay_inst_wint37/YUSED  (
    .I(\DM_delay_inst_wint37/GROM ),
    .O(DM_delay_inst_wint37)
  );
  defparam reset_IBUF_3_1157.INIT = 16'hCCCC;
  X_LUT4 reset_IBUF_3_1157 (
    .ADR0(VCC),
    .ADR1(reset_IBUF),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\reset_IBUF_3/GROM )
  );
  X_BUF \reset_IBUF_3/YUSED  (
    .I(\reset_IBUF_3/GROM ),
    .O(reset_IBUF_3)
  );
  defparam DLX_EXinst_Ker662001.INIT = 16'h0004;
  X_LUT4 DLX_EXinst_Ker662001 (
    .ADR0(DLX_IDinst_IR_opcode_field[0]),
    .ADR1(DLX_EXinst_N66112),
    .ADR2(N109130),
    .ADR3(DLX_IDinst_IR_opcode_field[1]),
    .O(\DLX_EXinst_N66202/FROM )
  );
  defparam \DLX_EXinst__n0006<0>635 .INIT = 16'h0400;
  X_LUT4 \DLX_EXinst__n0006<0>635  (
    .ADR0(DLX_IDinst_IR_function_field[2]),
    .ADR1(\DLX_EXinst_Mshift__n0027_Sh[0] ),
    .ADR2(DLX_IDinst_IR_function_field[3]),
    .ADR3(DLX_EXinst_N66202),
    .O(\DLX_EXinst_N66202/GROM )
  );
  X_BUF \DLX_EXinst_N66202/XUSED  (
    .I(\DLX_EXinst_N66202/FROM ),
    .O(DLX_EXinst_N66202)
  );
  X_BUF \DLX_EXinst_N66202/YUSED  (
    .I(\DLX_EXinst_N66202/GROM ),
    .O(CHOICE5976)
  );
  defparam reset_IBUF_4_1158.INIT = 16'hF0F0;
  X_LUT4 reset_IBUF_4_1158 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(reset_IBUF),
    .ADR3(VCC),
    .O(\reset_IBUF_4/GROM )
  );
  X_BUF \reset_IBUF_4/YUSED  (
    .I(\reset_IBUF_4/GROM ),
    .O(reset_IBUF_4)
  );
  defparam DM_delay_inst_wint381.INIT = 16'h00FF;
  X_LUT4 DM_delay_inst_wint381 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DM_delay_inst_wint37),
    .O(\DM_delay_inst_wint38/GROM )
  );
  X_BUF \DM_delay_inst_wint38/YUSED  (
    .I(\DM_delay_inst_wint38/GROM ),
    .O(DM_delay_inst_wint38)
  );
  defparam reset_IBUF_5_1159.INIT = 16'hCCCC;
  X_LUT4 reset_IBUF_5_1159 (
    .ADR0(VCC),
    .ADR1(reset_IBUF),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\reset_IBUF_5/GROM )
  );
  X_BUF \reset_IBUF_5/YUSED  (
    .I(\reset_IBUF_5/GROM ),
    .O(reset_IBUF_5)
  );
  defparam \DLX_IDinst_regB_eff<19>1 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst_regB_eff<19>1  (
    .ADR0(DLX_IDinst_N70716),
    .ADR1(DLX_IDinst_reg_out_B_RF[19]),
    .ADR2(DLX_IDinst__n0145),
    .ADR3(DLX_MEMinst_RF_data_in[19]),
    .O(\DLX_IDinst_regB_eff<19>/FROM )
  );
  defparam \DLX_IDinst_regB_eff<24>1 .INIT = 16'hECA0;
  X_LUT4 \DLX_IDinst_regB_eff<24>1  (
    .ADR0(DLX_IDinst_reg_out_B_RF[24]),
    .ADR1(DLX_IDinst__n0145),
    .ADR2(DLX_IDinst_N70716),
    .ADR3(DLX_MEMinst_RF_data_in[24]),
    .O(\DLX_IDinst_regB_eff<19>/GROM )
  );
  X_BUF \DLX_IDinst_regB_eff<19>/XUSED  (
    .I(\DLX_IDinst_regB_eff<19>/FROM ),
    .O(DLX_IDinst_regB_eff[19])
  );
  X_BUF \DLX_IDinst_regB_eff<19>/YUSED  (
    .I(\DLX_IDinst_regB_eff<19>/GROM ),
    .O(DLX_IDinst_regB_eff[24])
  );
  defparam DLX_IFlc_md_mda6_a1.INIT = 16'h3300;
  X_LUT4 DLX_IFlc_md_mda6_a1 (
    .ADR0(VCC),
    .ADR1(DLX_IFlc_pd_wint1),
    .ADR2(VCC),
    .ADR3(DLX_IFlc_md_wint5),
    .O(\DLX_IFlc_md_wint6/FROM )
  );
  defparam DLX_IFlc_md_mda2_a1.INIT = 16'h0F00;
  X_LUT4 DLX_IFlc_md_mda2_a1 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IFlc_pd_wint1),
    .ADR3(DLX_IFlc_md_wint1),
    .O(\DLX_IFlc_md_wint6/GROM )
  );
  X_BUF \DLX_IFlc_md_wint6/XUSED  (
    .I(\DLX_IFlc_md_wint6/FROM ),
    .O(DLX_IFlc_md_wint6)
  );
  X_BUF \DLX_IFlc_md_wint6/YUSED  (
    .I(\DLX_IFlc_md_wint6/GROM ),
    .O(DLX_IFlc_md_wint2)
  );
  defparam DLX_EXinst_Ker633771.INIT = 16'hCACA;
  X_LUT4 DLX_EXinst_Ker633771 (
    .ADR0(DLX_IDinst_reg_out_A[18]),
    .ADR1(DLX_IDinst_reg_out_A[16]),
    .ADR2(DLX_IDinst_reg_out_B[1]),
    .ADR3(VCC),
    .O(\DLX_EXinst_N63379/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0025_Sh<19>1 .INIT = 16'hFA50;
  X_LUT4 \DLX_EXinst_Mshift__n0025_Sh<19>1  (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N62881),
    .ADR3(DLX_EXinst_N63379),
    .O(\DLX_EXinst_N63379/GROM )
  );
  X_BUF \DLX_EXinst_N63379/XUSED  (
    .I(\DLX_EXinst_N63379/FROM ),
    .O(DLX_EXinst_N63379)
  );
  X_BUF \DLX_EXinst_N63379/YUSED  (
    .I(\DLX_EXinst_N63379/GROM ),
    .O(\DLX_EXinst_Mshift__n0025_Sh[19] )
  );
  defparam \DLX_EXinst__n0006<7>154 .INIT = 16'h5000;
  X_LUT4 \DLX_EXinst__n0006<7>154  (
    .ADR0(DLX_IDinst_reg_out_B[3]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N66226),
    .ADR3(DLX_EXinst_N62916),
    .O(\CHOICE3836/FROM )
  );
  defparam DLX_EXinst_Ker640971.INIT = 16'hF0CC;
  X_LUT4 DLX_EXinst_Ker640971 (
    .ADR0(VCC),
    .ADR1(\DLX_EXinst_Mshift__n0025_Sh[22] ),
    .ADR2(\DLX_EXinst_Mshift__n0025_Sh[14] ),
    .ADR3(DLX_IDinst_reg_out_B[3]),
    .O(\CHOICE3836/GROM )
  );
  X_BUF \CHOICE3836/XUSED  (
    .I(\CHOICE3836/FROM ),
    .O(CHOICE3836)
  );
  X_BUF \CHOICE3836/YUSED  (
    .I(\CHOICE3836/GROM ),
    .O(DLX_EXinst_N64099)
  );
  defparam DLX_EXinst_Ker634571.INIT = 16'hAACC;
  X_LUT4 DLX_EXinst_Ker634571 (
    .ADR0(DLX_IDinst_reg_out_A[16]),
    .ADR1(DLX_IDinst_reg_out_A[18]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_IR_function_field[1]),
    .O(\DLX_EXinst_N63459/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0027_Sh<19>1 .INIT = 16'hEE22;
  X_LUT4 \DLX_EXinst_Mshift__n0027_Sh<19>1  (
    .ADR0(DLX_EXinst_N62796),
    .ADR1(DLX_IDinst_IR_function_field_0_1),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N63459),
    .O(\DLX_EXinst_N63459/GROM )
  );
  X_BUF \DLX_EXinst_N63459/XUSED  (
    .I(\DLX_EXinst_N63459/FROM ),
    .O(DLX_EXinst_N63459)
  );
  X_BUF \DLX_EXinst_N63459/YUSED  (
    .I(\DLX_EXinst_N63459/GROM ),
    .O(\DLX_EXinst_Mshift__n0027_Sh[19] )
  );
  defparam DLX_IFinst_NPC_14_1_1160.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_14_1_1160 (
    .I(\NPC_eff<14>/OD ),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\NPC_eff<14>/OFF/RST ),
    .O(DLX_IFinst_NPC_14_1)
  );
  X_OR2 \NPC_eff<14>/OFF/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\NPC_eff<14>/OFF/RST )
  );
  defparam \DLX_EXinst__n0006<7>76 .INIT = 16'hC4C0;
  X_LUT4 \DLX_EXinst__n0006<7>76  (
    .ADR0(\DLX_IDinst_Imm[7] ),
    .ADR1(DLX_IDinst_reg_out_A[7]),
    .ADR2(DLX_EXinst__n0079),
    .ADR3(DLX_EXinst__n0080),
    .O(\CHOICE3818/FROM )
  );
  defparam \DLX_EXinst__n0006<1>29 .INIT = 16'hF200;
  X_LUT4 \DLX_EXinst__n0006<1>29  (
    .ADR0(DLX_EXinst__n0080),
    .ADR1(DLX_IDinst_IR_function_field[1]),
    .ADR2(DLX_EXinst__n0079),
    .ADR3(DLX_IDinst_reg_out_A[1]),
    .O(\CHOICE3818/GROM )
  );
  X_BUF \CHOICE3818/XUSED  (
    .I(\CHOICE3818/FROM ),
    .O(CHOICE3818)
  );
  X_BUF \CHOICE3818/YUSED  (
    .I(\CHOICE3818/GROM ),
    .O(CHOICE5663)
  );
  defparam DLX_IFlc_md_mda5_a1.INIT = 16'h3300;
  X_LUT4 DLX_IFlc_md_mda5_a1 (
    .ADR0(VCC),
    .ADR1(DLX_IFlc_pd_wint1),
    .ADR2(VCC),
    .ADR3(DLX_IFlc_md_wint4),
    .O(\DLX_IFlc_md_wint5/FROM )
  );
  defparam DLX_IFlc_md_mda37_a1.INIT = 16'h0F00;
  X_LUT4 DLX_IFlc_md_mda37_a1 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IFlc_pd_wint1),
    .ADR3(DLX_IFlc_md_wint36),
    .O(\DLX_IFlc_md_wint5/GROM )
  );
  X_BUF \DLX_IFlc_md_wint5/XUSED  (
    .I(\DLX_IFlc_md_wint5/FROM ),
    .O(DLX_IFlc_md_wint5)
  );
  X_BUF \DLX_IFlc_md_wint5/YUSED  (
    .I(\DLX_IFlc_md_wint5/GROM ),
    .O(DLX_IFlc_md_wint37)
  );
  defparam DM_delay_inst_wint391.INIT = 16'h0F0F;
  X_LUT4 DM_delay_inst_wint391 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DM_delay_inst_wint38),
    .ADR3(VCC),
    .O(\DM_delay_inst_wint39/GROM )
  );
  X_BUF \DM_delay_inst_wint39/YUSED  (
    .I(\DM_delay_inst_wint39/GROM ),
    .O(DM_delay_inst_wint39)
  );
  defparam DLX_EXinst_Ker627381.INIT = 16'hFFAA;
  X_LUT4 DLX_EXinst_Ker627381 (
    .ADR0(DLX_IDinst_reg_out_B[2]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[3]),
    .O(\DLX_EXinst_N62740/FROM )
  );
  defparam DLX_EXinst_Ker6509321.INIT = 16'h4408;
  X_LUT4 DLX_EXinst_Ker6509321 (
    .ADR0(DLX_IDinst_reg_out_B[5]),
    .ADR1(DLX_IDinst_reg_out_A[31]),
    .ADR2(DLX_IDinst_reg_out_B[1]),
    .ADR3(DLX_EXinst_N62740),
    .O(\DLX_EXinst_N62740/GROM )
  );
  X_BUF \DLX_EXinst_N62740/XUSED  (
    .I(\DLX_EXinst_N62740/FROM ),
    .O(DLX_EXinst_N62740)
  );
  X_BUF \DLX_EXinst_N62740/YUSED  (
    .I(\DLX_EXinst_N62740/GROM ),
    .O(CHOICE859)
  );
  defparam \DLX_EXinst__n0006<8>41 .INIT = 16'h0808;
  X_LUT4 \DLX_EXinst__n0006<8>41  (
    .ADR0(DLX_EXinst__n0081),
    .ADR1(\DLX_EXinst_Mshift__n0027_Sh[40] ),
    .ADR2(N109130),
    .ADR3(VCC),
    .O(\CHOICE3692/FROM )
  );
  defparam \DLX_EXinst__n0006<2>16 .INIT = 16'h5450;
  X_LUT4 \DLX_EXinst__n0006<2>16  (
    .ADR0(N109130),
    .ADR1(DLX_EXinst_N66373),
    .ADR2(CHOICE5491),
    .ADR3(\DLX_EXinst_Mshift__n0028_Sh[50] ),
    .O(\CHOICE3692/GROM )
  );
  X_BUF \CHOICE3692/XUSED  (
    .I(\CHOICE3692/FROM ),
    .O(CHOICE3692)
  );
  X_BUF \CHOICE3692/YUSED  (
    .I(\CHOICE3692/GROM ),
    .O(CHOICE5493)
  );
  defparam \DLX_IDinst_regB_eff<26>1 .INIT = 16'hECA0;
  X_LUT4 \DLX_IDinst_regB_eff<26>1  (
    .ADR0(DLX_IDinst_reg_out_B_RF[26]),
    .ADR1(DLX_MEMinst_RF_data_in[26]),
    .ADR2(DLX_IDinst_N70716),
    .ADR3(DLX_IDinst__n0145),
    .O(\DLX_IDinst_regB_eff<26>/FROM )
  );
  defparam \DLX_IDinst_regB_eff<25>1 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst_regB_eff<25>1  (
    .ADR0(DLX_IDinst_N70716),
    .ADR1(DLX_IDinst_reg_out_B_RF[25]),
    .ADR2(DLX_MEMinst_RF_data_in[25]),
    .ADR3(DLX_IDinst__n0145),
    .O(\DLX_IDinst_regB_eff<26>/GROM )
  );
  X_BUF \DLX_IDinst_regB_eff<26>/XUSED  (
    .I(\DLX_IDinst_regB_eff<26>/FROM ),
    .O(DLX_IDinst_regB_eff[26])
  );
  X_BUF \DLX_IDinst_regB_eff<26>/YUSED  (
    .I(\DLX_IDinst_regB_eff<26>/GROM ),
    .O(DLX_IDinst_regB_eff[25])
  );
  defparam DLX_EXinst_Ker628191.INIT = 16'hF0EE;
  X_LUT4 DLX_EXinst_Ker628191 (
    .ADR0(CHOICE1024),
    .ADR1(CHOICE1018),
    .ADR2(\DLX_EXinst_Mshift__n0027_Sh[1] ),
    .ADR3(DLX_IDinst_IR_function_field[2]),
    .O(\DLX_EXinst_N62821/FROM )
  );
  defparam \DLX_EXinst__n0006<5>46 .INIT = 16'h0200;
  X_LUT4 \DLX_EXinst__n0006<5>46  (
    .ADR0(DLX_EXinst__n0081),
    .ADR1(N109130),
    .ADR2(DLX_IDinst_IR_function_field[3]),
    .ADR3(DLX_EXinst_N62821),
    .O(\DLX_EXinst_N62821/GROM )
  );
  X_BUF \DLX_EXinst_N62821/XUSED  (
    .I(\DLX_EXinst_N62821/FROM ),
    .O(DLX_EXinst_N62821)
  );
  X_BUF \DLX_EXinst_N62821/YUSED  (
    .I(\DLX_EXinst_N62821/GROM ),
    .O(CHOICE4432)
  );
  defparam \DLX_EXinst_Mshift__n0025_Sh<6>10 .INIT = 16'hE040;
  X_LUT4 \DLX_EXinst_Mshift__n0025_Sh<6>10  (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(DLX_IDinst_reg_out_A[5]),
    .ADR2(DLX_IDinst_reg_out_B[0]),
    .ADR3(DLX_IDinst_reg_out_A[3]),
    .O(\CHOICE1294/FROM )
  );
  defparam DLX_EXinst_Ker651631.INIT = 16'hCCAA;
  X_LUT4 DLX_EXinst_Ker651631 (
    .ADR0(DLX_IDinst_reg_out_A[3]),
    .ADR1(DLX_IDinst_reg_out_A[5]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_IR_function_field_1_1),
    .O(\CHOICE1294/GROM )
  );
  X_BUF \CHOICE1294/XUSED  (
    .I(\CHOICE1294/FROM ),
    .O(CHOICE1294)
  );
  X_BUF \CHOICE1294/YUSED  (
    .I(\CHOICE1294/GROM ),
    .O(DLX_EXinst_N65165)
  );
  defparam DLX_EXinst_Ker634671.INIT = 16'hCACA;
  X_LUT4 DLX_EXinst_Ker634671 (
    .ADR0(DLX_IDinst_reg_out_A[22]),
    .ADR1(DLX_IDinst_reg_out_A[20]),
    .ADR2(DLX_IDinst_IR_function_field[1]),
    .ADR3(VCC),
    .O(\DLX_EXinst_N63469/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0027_Sh<23>1 .INIT = 16'hEE22;
  X_LUT4 \DLX_EXinst_Mshift__n0027_Sh<23>1  (
    .ADR0(DLX_EXinst_N62806),
    .ADR1(DLX_IDinst_IR_function_field_0_1),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N63469),
    .O(\DLX_EXinst_N63469/GROM )
  );
  X_BUF \DLX_EXinst_N63469/XUSED  (
    .I(\DLX_EXinst_N63469/FROM ),
    .O(DLX_EXinst_N63469)
  );
  X_BUF \DLX_EXinst_N63469/YUSED  (
    .I(\DLX_EXinst_N63469/GROM ),
    .O(\DLX_EXinst_Mshift__n0027_Sh[23] )
  );
  defparam DLX_EXinst_Ker633871.INIT = 16'hFC0C;
  X_LUT4 DLX_EXinst_Ker633871 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[22]),
    .ADR2(DLX_IDinst_reg_out_B[1]),
    .ADR3(DLX_IDinst_reg_out_A[20]),
    .O(\DLX_EXinst_N63389/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0025_Sh<23>1 .INIT = 16'hEE22;
  X_LUT4 \DLX_EXinst_Mshift__n0025_Sh<23>1  (
    .ADR0(DLX_EXinst_N62891),
    .ADR1(DLX_IDinst_reg_out_B[0]),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N63389),
    .O(\DLX_EXinst_N63389/GROM )
  );
  X_BUF \DLX_EXinst_N63389/XUSED  (
    .I(\DLX_EXinst_N63389/FROM ),
    .O(DLX_EXinst_N63389)
  );
  X_BUF \DLX_EXinst_N63389/YUSED  (
    .I(\DLX_EXinst_N63389/GROM ),
    .O(\DLX_EXinst_Mshift__n0025_Sh[23] )
  );
  defparam \DLX_EXinst__n0006<30>12 .INIT = 16'hC4C0;
  X_LUT4 \DLX_EXinst__n0006<30>12  (
    .ADR0(\DLX_IDinst_Imm[31] ),
    .ADR1(DLX_IDinst_reg_out_A[30]),
    .ADR2(DLX_EXinst__n0079),
    .ADR3(DLX_EXinst__n0080),
    .O(\CHOICE5256/FROM )
  );
  defparam \DLX_EXinst__n0006<19>9 .INIT = 16'hCC08;
  X_LUT4 \DLX_EXinst__n0006<19>9  (
    .ADR0(DLX_EXinst__n0080),
    .ADR1(DLX_IDinst_reg_out_A[19]),
    .ADR2(\DLX_IDinst_Imm[31] ),
    .ADR3(DLX_EXinst__n0079),
    .O(\CHOICE5256/GROM )
  );
  X_BUF \CHOICE5256/XUSED  (
    .I(\CHOICE5256/FROM ),
    .O(CHOICE5256)
  );
  X_BUF \CHOICE5256/YUSED  (
    .I(\CHOICE5256/GROM ),
    .O(CHOICE4941)
  );
  defparam DLX_EXinst_Ker627641.INIT = 16'hAAF0;
  X_LUT4 DLX_EXinst_Ker627641 (
    .ADR0(DLX_IDinst_reg_out_A[5]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[7]),
    .ADR3(DLX_IDinst_IR_function_field[1]),
    .O(\DLX_EXinst_N62766/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0027_Sh<8>1 .INIT = 16'hFA50;
  X_LUT4 \DLX_EXinst_Mshift__n0027_Sh<8>1  (
    .ADR0(DLX_IDinst_IR_function_field_0_1),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N63484),
    .ADR3(DLX_EXinst_N62766),
    .O(\DLX_EXinst_N62766/GROM )
  );
  X_BUF \DLX_EXinst_N62766/XUSED  (
    .I(\DLX_EXinst_N62766/FROM ),
    .O(DLX_EXinst_N62766)
  );
  X_BUF \DLX_EXinst_N62766/YUSED  (
    .I(\DLX_EXinst_N62766/GROM ),
    .O(\DLX_EXinst_Mshift__n0027_Sh[8] )
  );
  defparam DLX_EXinst_Ker634921.INIT = 16'hD8D8;
  X_LUT4 DLX_EXinst_Ker634921 (
    .ADR0(DLX_IDinst_IR_function_field[1]),
    .ADR1(DLX_IDinst_reg_out_A[14]),
    .ADR2(DLX_IDinst_reg_out_A[12]),
    .ADR3(VCC),
    .O(\DLX_EXinst_N63494/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0028_Sh<11>1 .INIT = 16'hEE22;
  X_LUT4 \DLX_EXinst_Mshift__n0028_Sh<11>1  (
    .ADR0(DLX_EXinst_N62986),
    .ADR1(DLX_IDinst_IR_function_field_0_1),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N63494),
    .O(\DLX_EXinst_N63494/GROM )
  );
  X_BUF \DLX_EXinst_N63494/XUSED  (
    .I(\DLX_EXinst_N63494/FROM ),
    .O(DLX_EXinst_N63494)
  );
  X_BUF \DLX_EXinst_N63494/YUSED  (
    .I(\DLX_EXinst_N63494/GROM ),
    .O(\DLX_EXinst_Mshift__n0028_Sh[11] )
  );
  defparam DLX_IFlc_md_mda38_a1.INIT = 16'h5050;
  X_LUT4 DLX_IFlc_md_mda38_a1 (
    .ADR0(DLX_IFlc_pd_wint1),
    .ADR1(VCC),
    .ADR2(DLX_IFlc_md_wint37),
    .ADR3(VCC),
    .O(\DLX_IFlc_md_wint38/FROM )
  );
  defparam DLX_IFlc_md_mda3_a1.INIT = 16'h00AA;
  X_LUT4 DLX_IFlc_md_mda3_a1 (
    .ADR0(DLX_IFlc_md_wint2),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IFlc_pd_wint1),
    .O(\DLX_IFlc_md_wint38/GROM )
  );
  X_BUF \DLX_IFlc_md_wint38/XUSED  (
    .I(\DLX_IFlc_md_wint38/FROM ),
    .O(DLX_IFlc_md_wint38)
  );
  X_BUF \DLX_IFlc_md_wint38/YUSED  (
    .I(\DLX_IFlc_md_wint38/GROM ),
    .O(DLX_IFlc_md_wint3)
  );
  defparam DLX_EXinst_Ker645851.INIT = 16'hAACC;
  X_LUT4 DLX_EXinst_Ker645851 (
    .ADR0(DLX_IDinst_reg_out_A[6]),
    .ADR1(DLX_IDinst_reg_out_A[4]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[1]),
    .O(\DLX_EXinst_N64587/FROM )
  );
  defparam DLX_EXinst_Ker634771.INIT = 16'hCFC0;
  X_LUT4 DLX_EXinst_Ker634771 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[4]),
    .ADR2(DLX_IDinst_IR_function_field[1]),
    .ADR3(DLX_IDinst_reg_out_A[6]),
    .O(\DLX_EXinst_N64587/GROM )
  );
  X_BUF \DLX_EXinst_N64587/XUSED  (
    .I(\DLX_EXinst_N64587/FROM ),
    .O(DLX_EXinst_N64587)
  );
  X_BUF \DLX_EXinst_N64587/YUSED  (
    .I(\DLX_EXinst_N64587/GROM ),
    .O(DLX_EXinst_N63479)
  );
  defparam \DLX_EXinst__n0006<5>76 .INIT = 16'hC0C8;
  X_LUT4 \DLX_EXinst__n0006<5>76  (
    .ADR0(DLX_EXinst__n0080),
    .ADR1(DLX_IDinst_reg_out_A[5]),
    .ADR2(DLX_EXinst__n0079),
    .ADR3(\DLX_IDinst_Imm[5] ),
    .O(\CHOICE4438/FROM )
  );
  defparam \DLX_EXinst__n0006<2>29 .INIT = 16'hCE00;
  X_LUT4 \DLX_EXinst__n0006<2>29  (
    .ADR0(DLX_EXinst__n0080),
    .ADR1(DLX_EXinst__n0079),
    .ADR2(DLX_IDinst_IR_function_field[2]),
    .ADR3(DLX_IDinst_reg_out_A[2]),
    .O(\CHOICE4438/GROM )
  );
  X_BUF \CHOICE4438/XUSED  (
    .I(\CHOICE4438/FROM ),
    .O(CHOICE4438)
  );
  X_BUF \CHOICE4438/YUSED  (
    .I(\CHOICE4438/GROM ),
    .O(CHOICE5497)
  );
  defparam DLX_EXinst_Ker64548.INIT = 16'hAFA0;
  X_LUT4 DLX_EXinst_Ker64548 (
    .ADR0(\DLX_EXinst_Mshift__n0028_Sh[22] ),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_IR_function_field[3]),
    .ADR3(N93905),
    .O(\DLX_EXinst_N64550/FROM )
  );
  defparam DLX_EXinst_Ker629341.INIT = 16'hFA50;
  X_LUT4 DLX_EXinst_Ker629341 (
    .ADR0(DLX_IDinst_IR_function_field[3]),
    .ADR1(VCC),
    .ADR2(\DLX_EXinst_Mshift__n0028_Sh[21] ),
    .ADR3(\DLX_EXinst_Mshift__n0024_Sh[29] ),
    .O(\DLX_EXinst_N64550/GROM )
  );
  X_BUF \DLX_EXinst_N64550/XUSED  (
    .I(\DLX_EXinst_N64550/FROM ),
    .O(DLX_EXinst_N64550)
  );
  X_BUF \DLX_EXinst_N64550/YUSED  (
    .I(\DLX_EXinst_N64550/GROM ),
    .O(DLX_EXinst_N62936)
  );
  defparam DLX_EXinst_Ker628541.INIT = 16'hACAC;
  X_LUT4 DLX_EXinst_Ker628541 (
    .ADR0(DLX_IDinst_reg_out_A[7]),
    .ADR1(DLX_IDinst_reg_out_A[9]),
    .ADR2(DLX_IDinst_reg_out_B[1]),
    .ADR3(VCC),
    .O(\DLX_EXinst_N62856/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0025_Sh<10>1 .INIT = 16'hFA50;
  X_LUT4 \DLX_EXinst_Mshift__n0025_Sh<10>1  (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N63359),
    .ADR3(DLX_EXinst_N62856),
    .O(\DLX_EXinst_N62856/GROM )
  );
  X_BUF \DLX_EXinst_N62856/XUSED  (
    .I(\DLX_EXinst_N62856/FROM ),
    .O(DLX_EXinst_N62856)
  );
  X_BUF \DLX_EXinst_N62856/YUSED  (
    .I(\DLX_EXinst_N62856/GROM ),
    .O(\DLX_EXinst_Mshift__n0025_Sh[10] )
  );
  defparam DLX_EXinst_Ker629191.INIT = 16'hFC0C;
  X_LUT4 DLX_EXinst_Ker629191 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[7]),
    .ADR2(DLX_IDinst_IR_function_field[1]),
    .ADR3(DLX_IDinst_reg_out_A[9]),
    .O(\DLX_EXinst_N62921/FROM )
  );
  defparam DLX_EXinst_Ker627741.INIT = 16'hFA0A;
  X_LUT4 DLX_EXinst_Ker627741 (
    .ADR0(DLX_IDinst_reg_out_A[11]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_IR_function_field[1]),
    .ADR3(DLX_IDinst_reg_out_A[9]),
    .O(\DLX_EXinst_N62921/GROM )
  );
  X_BUF \DLX_EXinst_N62921/XUSED  (
    .I(\DLX_EXinst_N62921/FROM ),
    .O(DLX_EXinst_N62921)
  );
  X_BUF \DLX_EXinst_N62921/YUSED  (
    .I(\DLX_EXinst_N62921/GROM ),
    .O(DLX_EXinst_N62776)
  );
  defparam \DLX_EXinst_Mshift__n0026_Sh<50>_SW0 .INIT = 16'hF5A0;
  X_LUT4 \DLX_EXinst_Mshift__n0026_Sh<50>_SW0  (
    .ADR0(DLX_IDinst_reg_out_B_3_1),
    .ADR1(VCC),
    .ADR2(\DLX_EXinst_Mshift__n0026_Sh[30] ),
    .ADR3(\DLX_EXinst_Mshift__n0026_Sh[22] ),
    .O(\N94255/FROM )
  );
  defparam DLX_EXinst_Ker651581.INIT = 16'hF0AA;
  X_LUT4 DLX_EXinst_Ker651581 (
    .ADR0(\DLX_EXinst_Mshift__n0026_Sh[11] ),
    .ADR1(VCC),
    .ADR2(\DLX_EXinst_Mshift__n0026_Sh[19] ),
    .ADR3(DLX_IDinst_reg_out_B_3_1),
    .O(\N94255/GROM )
  );
  X_BUF \N94255/XUSED  (
    .I(\N94255/FROM ),
    .O(N94255)
  );
  X_BUF \N94255/YUSED  (
    .I(\N94255/GROM ),
    .O(DLX_EXinst_N65160)
  );
  defparam \DLX_IDinst_regB_eff<28>1 .INIT = 16'hECA0;
  X_LUT4 \DLX_IDinst_regB_eff<28>1  (
    .ADR0(DLX_IDinst__n0145),
    .ADR1(DLX_IDinst_N70716),
    .ADR2(DLX_MEMinst_RF_data_in[28]),
    .ADR3(DLX_IDinst_reg_out_B_RF[28]),
    .O(\DLX_IDinst_regB_eff<28>/FROM )
  );
  defparam \DLX_IDinst_regB_eff<27>1 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst_regB_eff<27>1  (
    .ADR0(DLX_MEMinst_RF_data_in[27]),
    .ADR1(DLX_IDinst__n0145),
    .ADR2(DLX_IDinst_reg_out_B_RF[27]),
    .ADR3(DLX_IDinst_N70716),
    .O(\DLX_IDinst_regB_eff<28>/GROM )
  );
  X_BUF \DLX_IDinst_regB_eff<28>/XUSED  (
    .I(\DLX_IDinst_regB_eff<28>/FROM ),
    .O(DLX_IDinst_regB_eff[28])
  );
  X_BUF \DLX_IDinst_regB_eff<28>/YUSED  (
    .I(\DLX_IDinst_regB_eff<28>/GROM ),
    .O(DLX_IDinst_regB_eff[27])
  );
  defparam DLX_IDinst__n0133_SW0.INIT = 16'hFCFF;
  X_LUT4 DLX_IDinst__n0133_SW0 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_IR_latched[29]),
    .ADR2(DLX_IDinst_IR_latched[30]),
    .ADR3(DLX_IDinst_IR_latched[31]),
    .O(\N95468/FROM )
  );
  defparam DLX_IDinst__n0133_1161.INIT = 16'h0075;
  X_LUT4 DLX_IDinst__n0133_1161 (
    .ADR0(DLX_IDinst_IR_latched[27]),
    .ADR1(DLX_IDinst_IR_latched[28]),
    .ADR2(DLX_IDinst_IR_latched[26]),
    .ADR3(N95468),
    .O(\N95468/GROM )
  );
  X_BUF \N95468/XUSED  (
    .I(\N95468/FROM ),
    .O(N95468)
  );
  X_BUF \N95468/YUSED  (
    .I(\N95468/GROM ),
    .O(DLX_IDinst__n0133)
  );
  defparam DLX_IDinst_Ker69955112.INIT = 16'h0E0A;
  X_LUT4 DLX_IDinst_Ker69955112 (
    .ADR0(CHOICE1444),
    .ADR1(CHOICE1436),
    .ADR2(DLX_IDinst_IR_opcode_field[5]),
    .ADR3(DLX_IDinst_IR_opcode_field[3]),
    .O(\CHOICE1446/FROM )
  );
  defparam DLX_IDinst_Ker69955126.INIT = 16'hFF54;
  X_LUT4 DLX_IDinst_Ker69955126 (
    .ADR0(DLX_IDinst_IR_opcode_field[3]),
    .ADR1(CHOICE1425),
    .ADR2(CHOICE1418),
    .ADR3(CHOICE1446),
    .O(\CHOICE1446/GROM )
  );
  X_BUF \CHOICE1446/XUSED  (
    .I(\CHOICE1446/FROM ),
    .O(CHOICE1446)
  );
  X_BUF \CHOICE1446/YUSED  (
    .I(\CHOICE1446/GROM ),
    .O(N98613)
  );
  defparam DLX_IDlc_md_mda4_a1.INIT = 16'h00CC;
  X_LUT4 DLX_IDlc_md_mda4_a1 (
    .ADR0(VCC),
    .ADR1(DLX_IDlc_md_wint3),
    .ADR2(VCC),
    .ADR3(DLX_IDlc_pd_wint1),
    .O(\DLX_IDlc_md_wint4/FROM )
  );
  defparam DLX_IDlc_md_mda1_a1.INIT = 16'h00AA;
  X_LUT4 DLX_IDlc_md_mda1_a1 (
    .ADR0(DLX_IDlc_ridp3),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDlc_pd_wint1),
    .O(\DLX_IDlc_md_wint4/GROM )
  );
  X_BUF \DLX_IDlc_md_wint4/XUSED  (
    .I(\DLX_IDlc_md_wint4/FROM ),
    .O(DLX_IDlc_md_wint4)
  );
  X_BUF \DLX_IDlc_md_wint4/YUSED  (
    .I(\DLX_IDlc_md_wint4/GROM ),
    .O(DLX_IDlc_md_wint1)
  );
  defparam \DLX_IDinst__n0117<10>29 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst__n0117<10>29  (
    .ADR0(CHOICE2254),
    .ADR1(N101161),
    .ADR2(DLX_IDinst_N69914),
    .ADR3(DLX_IDinst_regA_eff[10]),
    .O(\DLX_IDinst_reg_out_A<10>/FROM )
  );
  defparam \DLX_IDinst__n0117<10>39 .INIT = 16'hFFA0;
  X_LUT4 \DLX_IDinst__n0117<10>39  (
    .ADR0(DLX_IDinst__n0310),
    .ADR1(VCC),
    .ADR2(DLX_IFinst_NPC[10]),
    .ADR3(CHOICE2257),
    .O(N103352)
  );
  X_BUF \DLX_IDinst_reg_out_A<10>/XUSED  (
    .I(\DLX_IDinst_reg_out_A<10>/FROM ),
    .O(CHOICE2257)
  );
  defparam \DLX_IDinst__n0117<26>15 .INIT = 16'h3808;
  X_LUT4 \DLX_IDinst__n0117<26>15  (
    .ADR0(DLX_IDinst_Cause_Reg[26]),
    .ADR1(DLX_IDinst_regA_index[0]),
    .ADR2(DLX_IDinst_regA_index[1]),
    .ADR3(DLX_IDinst_EPC[26]),
    .O(\CHOICE2446/FROM )
  );
  defparam \DLX_IDinst__n0117<11>15 .INIT = 16'h0AC0;
  X_LUT4 \DLX_IDinst__n0117<11>15  (
    .ADR0(DLX_IDinst_EPC[11]),
    .ADR1(DLX_IDinst_Cause_Reg[11]),
    .ADR2(DLX_IDinst_regA_index[0]),
    .ADR3(DLX_IDinst_regA_index[1]),
    .O(\CHOICE2446/GROM )
  );
  X_BUF \CHOICE2446/XUSED  (
    .I(\CHOICE2446/FROM ),
    .O(CHOICE2446)
  );
  X_BUF \CHOICE2446/YUSED  (
    .I(\CHOICE2446/GROM ),
    .O(CHOICE2278)
  );
  defparam \DLX_IDinst__n0116<0>14 .INIT = 16'hA808;
  X_LUT4 \DLX_IDinst__n0116<0>14  (
    .ADR0(DLX_IDinst_N70647),
    .ADR1(N100686),
    .ADR2(DLX_IDinst__n0135),
    .ADR3(N98420),
    .O(\CHOICE2924/FROM )
  );
  defparam \DLX_IDinst__n0116<0>25 .INIT = 16'hEEE0;
  X_LUT4 \DLX_IDinst__n0116<0>25  (
    .ADR0(DLX_IDinst__n0136),
    .ADR1(DLX_IDinst__n0135),
    .ADR2(N98613),
    .ADR3(CHOICE2924),
    .O(\CHOICE2924/GROM )
  );
  X_BUF \CHOICE2924/XUSED  (
    .I(\CHOICE2924/FROM ),
    .O(CHOICE2924)
  );
  X_BUF \CHOICE2924/YUSED  (
    .I(\CHOICE2924/GROM ),
    .O(CHOICE2927)
  );
  defparam \DLX_EXinst_Mshift__n0027_Sh<6> .INIT = 16'hFC0C;
  X_LUT4 \DLX_EXinst_Mshift__n0027_Sh<6>  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N63479),
    .ADR2(DLX_IDinst_IR_function_field_0_1),
    .ADR3(N94155),
    .O(\DLX_EXinst_Mshift__n0027_Sh<6>/FROM )
  );
  defparam DLX_EXinst_Ker628241.INIT = 16'hDD88;
  X_LUT4 DLX_EXinst_Ker628241 (
    .ADR0(DLX_IDinst_IR_function_field[2]),
    .ADR1(\DLX_EXinst_Mshift__n0027_Sh[2] ),
    .ADR2(VCC),
    .ADR3(\DLX_EXinst_Mshift__n0027_Sh[6] ),
    .O(\DLX_EXinst_Mshift__n0027_Sh<6>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0027_Sh<6>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0027_Sh<6>/FROM ),
    .O(\DLX_EXinst_Mshift__n0027_Sh[6] )
  );
  X_BUF \DLX_EXinst_Mshift__n0027_Sh<6>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0027_Sh<6>/GROM ),
    .O(DLX_EXinst_N62826)
  );
  defparam \DLX_EXinst_Mshift__n0024_Sh<61>1 .INIT = 16'h4C4C;
  X_LUT4 \DLX_EXinst_Mshift__n0024_Sh<61>1  (
    .ADR0(DLX_IDinst_IR_function_field_0_1),
    .ADR1(DLX_IDinst_reg_out_A[31]),
    .ADR2(DLX_IDinst_IR_function_field_1_1),
    .ADR3(VCC),
    .O(\DLX_EXinst_Mshift__n0024_Sh<61>/FROM )
  );
  defparam DLX_EXinst_Ker6511312.INIT = 16'hA808;
  X_LUT4 DLX_EXinst_Ker6511312 (
    .ADR0(\DLX_IDinst_Imm[5] ),
    .ADR1(DLX_IDinst_reg_out_A[31]),
    .ADR2(DLX_IDinst_IR_function_field_2_1),
    .ADR3(\DLX_EXinst_Mshift__n0024_Sh[61] ),
    .O(\DLX_EXinst_Mshift__n0024_Sh<61>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0024_Sh<61>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0024_Sh<61>/FROM ),
    .O(\DLX_EXinst_Mshift__n0024_Sh[61] )
  );
  X_BUF \DLX_EXinst_Mshift__n0024_Sh<61>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0024_Sh<61>/GROM ),
    .O(CHOICE1985)
  );
  defparam \DLX_EXinst_Mshift__n0024_Sh<29>1 .INIT = 16'hF3C0;
  X_LUT4 \DLX_EXinst_Mshift__n0024_Sh<29>1  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_IR_function_field_1_1),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(DLX_EXinst_N62709),
    .O(\DLX_EXinst_Mshift__n0024_Sh<29>/FROM )
  );
  defparam DLX_EXinst_Ker6582012.INIT = 16'h4540;
  X_LUT4 DLX_EXinst_Ker6582012 (
    .ADR0(\DLX_IDinst_Imm[5] ),
    .ADR1(DLX_IDinst_reg_out_A[31]),
    .ADR2(DLX_EXinst_N62733),
    .ADR3(\DLX_EXinst_Mshift__n0024_Sh[29] ),
    .O(\DLX_EXinst_Mshift__n0024_Sh<29>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0024_Sh<29>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0024_Sh<29>/FROM ),
    .O(\DLX_EXinst_Mshift__n0024_Sh[29] )
  );
  X_BUF \DLX_EXinst_Mshift__n0024_Sh<29>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0024_Sh<29>/GROM ),
    .O(CHOICE2043)
  );
  defparam DLX_IDlc_md_mda2_a1.INIT = 16'h00AA;
  X_LUT4 DLX_IDlc_md_mda2_a1 (
    .ADR0(DLX_IDlc_md_wint1),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDlc_pd_wint1),
    .O(\DLX_IDlc_md_wint2/GROM )
  );
  X_BUF \DLX_IDlc_md_wint2/YUSED  (
    .I(\DLX_IDlc_md_wint2/GROM ),
    .O(DLX_IDlc_md_wint2)
  );
  defparam \DLX_EXinst_Mshift__n0028_Sh<50>1 .INIT = 16'hF3C0;
  X_LUT4 \DLX_EXinst_Mshift__n0028_Sh<50>1  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_IR_function_field_2_1),
    .ADR2(DLX_EXinst_N63026),
    .ADR3(DLX_EXinst_N64859),
    .O(\DLX_EXinst_Mshift__n0028_Sh<50>/FROM )
  );
  defparam \DLX_EXinst__n0006<18>109_SW0 .INIT = 16'hEECC;
  X_LUT4 \DLX_EXinst__n0006<18>109_SW0  (
    .ADR0(DLX_EXinst__n0082),
    .ADR1(CHOICE5432),
    .ADR2(VCC),
    .ADR3(\DLX_EXinst_Mshift__n0028_Sh[50] ),
    .O(\DLX_EXinst_Mshift__n0028_Sh<50>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0028_Sh<50>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0028_Sh<50>/FROM ),
    .O(\DLX_EXinst_Mshift__n0028_Sh[50] )
  );
  X_BUF \DLX_EXinst_Mshift__n0028_Sh<50>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0028_Sh<50>/GROM ),
    .O(N126407)
  );
  defparam \DLX_EXinst_Mshift__n0028_Sh<18>1 .INIT = 16'hEE22;
  X_LUT4 \DLX_EXinst_Mshift__n0028_Sh<18>1  (
    .ADR0(DLX_EXinst_N63509),
    .ADR1(DLX_IDinst_IR_function_field_0_1),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N63006),
    .O(\DLX_EXinst_Mshift__n0028_Sh<18>/FROM )
  );
  defparam DLX_EXinst_Ker648571.INIT = 16'hFDA8;
  X_LUT4 DLX_EXinst_Ker648571 (
    .ADR0(DLX_IDinst_IR_function_field_3_1),
    .ADR1(CHOICE1114),
    .ADR2(CHOICE1120),
    .ADR3(\DLX_EXinst_Mshift__n0028_Sh[18] ),
    .O(\DLX_EXinst_Mshift__n0028_Sh<18>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0028_Sh<18>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0028_Sh<18>/FROM ),
    .O(\DLX_EXinst_Mshift__n0028_Sh[18] )
  );
  X_BUF \DLX_EXinst_Mshift__n0028_Sh<18>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0028_Sh<18>/GROM ),
    .O(DLX_EXinst_N64859)
  );
  defparam \DLX_IDinst__n0117<11>29 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst__n0117<11>29  (
    .ADR0(DLX_IDinst_regA_eff[11]),
    .ADR1(DLX_IDinst_N69914),
    .ADR2(N101161),
    .ADR3(CHOICE2278),
    .O(\DLX_IDinst_reg_out_A<11>/FROM )
  );
  defparam \DLX_IDinst__n0117<11>39 .INIT = 16'hFFC0;
  X_LUT4 \DLX_IDinst__n0117<11>39  (
    .ADR0(VCC),
    .ADR1(DLX_IFinst_NPC[11]),
    .ADR2(DLX_IDinst__n0310),
    .ADR3(CHOICE2281),
    .O(N103488)
  );
  X_BUF \DLX_IDinst_reg_out_A<11>/XUSED  (
    .I(\DLX_IDinst_reg_out_A<11>/FROM ),
    .O(CHOICE2281)
  );
  defparam \DLX_IDinst__n0117<17>15 .INIT = 16'h5808;
  X_LUT4 \DLX_IDinst__n0117<17>15  (
    .ADR0(DLX_IDinst_regA_index[0]),
    .ADR1(DLX_IDinst_Cause_Reg[17]),
    .ADR2(DLX_IDinst_regA_index[1]),
    .ADR3(DLX_IDinst_EPC[17]),
    .O(\CHOICE2326/FROM )
  );
  defparam \DLX_IDinst__n0117<20>15 .INIT = 16'h22C0;
  X_LUT4 \DLX_IDinst__n0117<20>15  (
    .ADR0(DLX_IDinst_Cause_Reg[20]),
    .ADR1(DLX_IDinst_regA_index[1]),
    .ADR2(DLX_IDinst_EPC[20]),
    .ADR3(DLX_IDinst_regA_index[0]),
    .O(\CHOICE2326/GROM )
  );
  X_BUF \CHOICE2326/XUSED  (
    .I(\CHOICE2326/FROM ),
    .O(CHOICE2326)
  );
  X_BUF \CHOICE2326/YUSED  (
    .I(\CHOICE2326/GROM ),
    .O(CHOICE2374)
  );
  defparam DLX_EXinst_Ker66307161_SW0_SW0.INIT = 16'hA000;
  X_LUT4 DLX_EXinst_Ker66307161_SW0_SW0 (
    .ADR0(CHOICE3595),
    .ADR1(VCC),
    .ADR2(CHOICE3610),
    .ADR3(CHOICE3603),
    .O(\N127257/FROM )
  );
  defparam DLX_EXinst_Ker66307161_SW0.INIT = 16'h7FFF;
  X_LUT4 DLX_EXinst_Ker66307161_SW0 (
    .ADR0(CHOICE3588),
    .ADR1(CHOICE3572),
    .ADR2(CHOICE3579),
    .ADR3(N127257),
    .O(\N127257/GROM )
  );
  X_BUF \N127257/XUSED  (
    .I(\N127257/FROM ),
    .O(N127257)
  );
  X_BUF \N127257/YUSED  (
    .I(\N127257/GROM ),
    .O(N126424)
  );
  defparam DLX_EXinst_Ker65384107.INIT = 16'hF888;
  X_LUT4 DLX_EXinst_Ker65384107 (
    .ADR0(N110065),
    .ADR1(N126272),
    .ADR2(DLX_EXinst_N66507),
    .ADR3(CHOICE3024),
    .O(\N107780/FROM )
  );
  defparam \DLX_EXinst__n0006<7>93 .INIT = 16'hFEFC;
  X_LUT4 \DLX_EXinst__n0006<7>93  (
    .ADR0(DLX_IDinst_IR_function_field[4]),
    .ADR1(CHOICE3802),
    .ADR2(CHOICE3819),
    .ADR3(N107780),
    .O(\N107780/GROM )
  );
  X_BUF \N107780/XUSED  (
    .I(\N107780/FROM ),
    .O(N107780)
  );
  X_BUF \N107780/YUSED  (
    .I(\N107780/GROM ),
    .O(CHOICE3820)
  );
  defparam DLX_IDlc_md_mda3_a1.INIT = 16'h00F0;
  X_LUT4 DLX_IDlc_md_mda3_a1 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IDlc_md_wint2),
    .ADR3(DLX_IDlc_pd_wint1),
    .O(\DLX_IDlc_md_wint3/GROM )
  );
  X_BUF \DLX_IDlc_md_wint3/YUSED  (
    .I(\DLX_IDlc_md_wint3/GROM ),
    .O(DLX_IDlc_md_wint3)
  );
  defparam \DLX_EXinst_Mshift__n0024_Sh<80>1 .INIT = 16'hFA50;
  X_LUT4 \DLX_EXinst_Mshift__n0024_Sh<80>1  (
    .ADR0(DLX_IDinst_IR_function_field_2_1),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N64565),
    .ADR3(DLX_EXinst_N62715),
    .O(\DLX_EXinst_Mshift__n0024_Sh<80>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0024_Sh<80>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0024_Sh<80>/GROM ),
    .O(\DLX_EXinst_Mshift__n0024_Sh[80] )
  );
  defparam \DLX_IDinst__n0117<12>29 .INIT = 16'hEAC0;
  X_LUT4 \DLX_IDinst__n0117<12>29  (
    .ADR0(CHOICE2266),
    .ADR1(DLX_IDinst_regA_eff[12]),
    .ADR2(DLX_IDinst_N69914),
    .ADR3(N101161),
    .O(\DLX_IDinst_reg_out_A<12>/FROM )
  );
  defparam \DLX_IDinst__n0117<12>39 .INIT = 16'hFFA0;
  X_LUT4 \DLX_IDinst__n0117<12>39  (
    .ADR0(DLX_IDinst__n0310),
    .ADR1(VCC),
    .ADR2(DLX_IFinst_NPC[12]),
    .ADR3(CHOICE2269),
    .O(N103420)
  );
  X_BUF \DLX_IDinst_reg_out_A<12>/XUSED  (
    .I(\DLX_IDinst_reg_out_A<12>/FROM ),
    .O(CHOICE2269)
  );
  defparam \DLX_IDinst__n0117<20>29 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst__n0117<20>29  (
    .ADR0(N101161),
    .ADR1(CHOICE2374),
    .ADR2(DLX_IDinst_regA_eff[20]),
    .ADR3(DLX_IDinst_N69914),
    .O(\DLX_IDinst_reg_out_A<20>/FROM )
  );
  defparam \DLX_IDinst__n0117<20>39 .INIT = 16'hFF88;
  X_LUT4 \DLX_IDinst__n0117<20>39  (
    .ADR0(DLX_IFinst_NPC[20]),
    .ADR1(DLX_IDinst__n0310),
    .ADR2(VCC),
    .ADR3(CHOICE2377),
    .O(N104032)
  );
  X_BUF \DLX_IDinst_reg_out_A<20>/XUSED  (
    .I(\DLX_IDinst_reg_out_A<20>/FROM ),
    .O(CHOICE2377)
  );
  defparam DLX_EXinst_Ker66248129.INIT = 16'h0001;
  X_LUT4 DLX_EXinst_Ker66248129 (
    .ADR0(\DLX_IDinst_Imm[8] ),
    .ADR1(\DLX_IDinst_Imm[10] ),
    .ADR2(\DLX_IDinst_Imm[9] ),
    .ADR3(\DLX_IDinst_Imm[7] ),
    .O(\CHOICE3406/FROM )
  );
  defparam DLX_EXinst_Ker66248153.INIT = 16'h1000;
  X_LUT4 DLX_EXinst_Ker66248153 (
    .ADR0(\DLX_IDinst_Imm[15] ),
    .ADR1(\DLX_IDinst_Imm[31] ),
    .ADR2(CHOICE3399),
    .ADR3(CHOICE3406),
    .O(\CHOICE3406/GROM )
  );
  X_BUF \CHOICE3406/XUSED  (
    .I(\CHOICE3406/FROM ),
    .O(CHOICE3406)
  );
  X_BUF \CHOICE3406/YUSED  (
    .I(\CHOICE3406/GROM ),
    .O(CHOICE3408)
  );
  defparam DLX_IDinst_Ker6995525.INIT = 16'h00CC;
  X_LUT4 DLX_IDinst_Ker6995525 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_IR_opcode_field[5]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_IR_opcode_field[4]),
    .O(\CHOICE1424/FROM )
  );
  defparam DLX_IDinst_Ker6995530.INIT = 16'h5D00;
  X_LUT4 DLX_IDinst_Ker6995530 (
    .ADR0(DLX_IDinst_IR_opcode_field[1]),
    .ADR1(DLX_IDinst_IR_opcode_field[0]),
    .ADR2(DLX_IDinst_IR_opcode_field[2]),
    .ADR3(CHOICE1424),
    .O(\CHOICE1424/GROM )
  );
  X_BUF \CHOICE1424/XUSED  (
    .I(\CHOICE1424/FROM ),
    .O(CHOICE1424)
  );
  X_BUF \CHOICE1424/YUSED  (
    .I(\CHOICE1424/GROM ),
    .O(CHOICE1425)
  );
  defparam \DLX_IDinst__n0117<30>15 .INIT = 16'h4A40;
  X_LUT4 \DLX_IDinst__n0117<30>15  (
    .ADR0(DLX_IDinst_regA_index[1]),
    .ADR1(DLX_IDinst_Cause_Reg[30]),
    .ADR2(DLX_IDinst_regA_index[0]),
    .ADR3(DLX_IDinst_EPC[30]),
    .O(\CHOICE2494/FROM )
  );
  defparam \DLX_IDinst__n0117<13>15 .INIT = 16'h0CA0;
  X_LUT4 \DLX_IDinst__n0117<13>15  (
    .ADR0(DLX_IDinst_EPC[13]),
    .ADR1(DLX_IDinst_Cause_Reg[13]),
    .ADR2(DLX_IDinst_regA_index[1]),
    .ADR3(DLX_IDinst_regA_index[0]),
    .O(\CHOICE2494/GROM )
  );
  X_BUF \CHOICE2494/XUSED  (
    .I(\CHOICE2494/FROM ),
    .O(CHOICE2494)
  );
  X_BUF \CHOICE2494/YUSED  (
    .I(\CHOICE2494/GROM ),
    .O(CHOICE2290)
  );
  defparam DLX_IFlc_pd_wint11.INIT = 16'h00FF;
  X_LUT4 DLX_IFlc_pd_wint11 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_reqin_IF),
    .O(\DLX_IFlc_pd_wint1/FROM )
  );
  defparam DLX_IFlc_ridp21.INIT = 16'hFF00;
  X_LUT4 DLX_IFlc_ridp21 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IFlc_pd_wint1),
    .O(\DLX_IFlc_pd_wint1/GROM )
  );
  X_BUF \DLX_IFlc_pd_wint1/XUSED  (
    .I(\DLX_IFlc_pd_wint1/FROM ),
    .O(DLX_IFlc_pd_wint1)
  );
  X_BUF \DLX_IFlc_pd_wint1/YUSED  (
    .I(\DLX_IFlc_pd_wint1/GROM ),
    .O(DLX_IFlc_ridp2)
  );
  defparam DLX_EXinst__n001880_SW0.INIT = 16'hFFFC;
  X_LUT4 DLX_EXinst__n001880_SW0 (
    .ADR0(VCC),
    .ADR1(CHOICE3168),
    .ADR2(DLX_IDinst_IR_opcode_field[1]),
    .ADR3(DLX_IDinst_IR_opcode_field[2]),
    .O(\N126205/FROM )
  );
  defparam DLX_EXinst__n001880.INIT = 16'hEFEC;
  X_LUT4 DLX_EXinst__n001880 (
    .ADR0(N126207),
    .ADR1(DLX_IDinst_IR_opcode_field[4]),
    .ADR2(DLX_IDinst_IR_opcode_field[5]),
    .ADR3(N126205),
    .O(\N126205/GROM )
  );
  X_BUF \N126205/XUSED  (
    .I(\N126205/FROM ),
    .O(N126205)
  );
  X_BUF \N126205/YUSED  (
    .I(\N126205/GROM ),
    .O(N108704)
  );
  defparam \DLX_EXinst_Mshift__n0025_Sh<44>_SW0 .INIT = 16'h03F3;
  X_LUT4 \DLX_EXinst_Mshift__n0025_Sh<44>_SW0  (
    .ADR0(VCC),
    .ADR1(\DLX_EXinst_Mshift__n0025_Sh[12] ),
    .ADR2(DLX_IDinst_reg_out_B_2_1),
    .ADR3(\DLX_EXinst_Mshift__n0025_Sh[8] ),
    .O(\N93587/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0025_Sh<44> .INIT = 16'h88BB;
  X_LUT4 \DLX_EXinst_Mshift__n0025_Sh<44>  (
    .ADR0(DLX_EXinst_N62901),
    .ADR1(DLX_IDinst_reg_out_B_3_1),
    .ADR2(VCC),
    .ADR3(N93587),
    .O(\N93587/GROM )
  );
  X_BUF \N93587/XUSED  (
    .I(\N93587/FROM ),
    .O(N93587)
  );
  X_BUF \N93587/YUSED  (
    .I(\N93587/GROM ),
    .O(\DLX_EXinst_Mshift__n0025_Sh[44] )
  );
  defparam \DLX_IDinst__n0117<21>29 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst__n0117<21>29  (
    .ADR0(DLX_IDinst_N69914),
    .ADR1(DLX_IDinst_regA_eff[21]),
    .ADR2(CHOICE2398),
    .ADR3(N101161),
    .O(\DLX_IDinst_reg_out_A<21>/FROM )
  );
  defparam \DLX_IDinst__n0117<21>39 .INIT = 16'hFFC0;
  X_LUT4 \DLX_IDinst__n0117<21>39  (
    .ADR0(VCC),
    .ADR1(DLX_IFinst_NPC[21]),
    .ADR2(DLX_IDinst__n0310),
    .ADR3(CHOICE2401),
    .O(N104168)
  );
  X_BUF \DLX_IDinst_reg_out_A<21>/XUSED  (
    .I(\DLX_IDinst_reg_out_A<21>/FROM ),
    .O(CHOICE2401)
  );
  defparam \DLX_IDinst__n0117<13>29 .INIT = 16'hECA0;
  X_LUT4 \DLX_IDinst__n0117<13>29  (
    .ADR0(DLX_IDinst_N69914),
    .ADR1(N101161),
    .ADR2(DLX_IDinst_regA_eff[13]),
    .ADR3(CHOICE2290),
    .O(\DLX_IDinst_reg_out_A<13>/FROM )
  );
  defparam \DLX_IDinst__n0117<13>39 .INIT = 16'hFFA0;
  X_LUT4 \DLX_IDinst__n0117<13>39  (
    .ADR0(DLX_IDinst__n0310),
    .ADR1(VCC),
    .ADR2(DLX_IFinst_NPC[13]),
    .ADR3(CHOICE2293),
    .O(N103556)
  );
  X_BUF \DLX_IDinst_reg_out_A<13>/XUSED  (
    .I(\DLX_IDinst_reg_out_A<13>/FROM ),
    .O(CHOICE2293)
  );
  defparam \DLX_IDinst__n0117<4>15 .INIT = 16'h6420;
  X_LUT4 \DLX_IDinst__n0117<4>15  (
    .ADR0(DLX_IDinst_regA_index[1]),
    .ADR1(DLX_IDinst_regA_index[0]),
    .ADR2(DLX_IDinst_EPC[4]),
    .ADR3(DLX_IDinst_Cause_Reg[4]),
    .O(\CHOICE2170/FROM )
  );
  defparam \DLX_IDinst__n0117<14>15 .INIT = 16'h0CA0;
  X_LUT4 \DLX_IDinst__n0117<14>15  (
    .ADR0(DLX_IDinst_Cause_Reg[14]),
    .ADR1(DLX_IDinst_EPC[14]),
    .ADR2(DLX_IDinst_regA_index[0]),
    .ADR3(DLX_IDinst_regA_index[1]),
    .O(\CHOICE2170/GROM )
  );
  X_BUF \CHOICE2170/XUSED  (
    .I(\CHOICE2170/FROM ),
    .O(CHOICE2170)
  );
  X_BUF \CHOICE2170/YUSED  (
    .I(\CHOICE2170/GROM ),
    .O(CHOICE2302)
  );
  defparam \DLX_EXinst__n0006<2>372_SW0 .INIT = 16'hFEFA;
  X_LUT4 \DLX_EXinst__n0006<2>372_SW0  (
    .ADR0(CHOICE5564),
    .ADR1(DLX_EXinst__n0114),
    .ADR2(CHOICE5543),
    .ADR3(DLX_EXinst__n0016[2]),
    .O(\N126816/FROM )
  );
  defparam \DLX_EXinst__n0006<2>372 .INIT = 16'hE4A0;
  X_LUT4 \DLX_EXinst__n0006<2>372  (
    .ADR0(DLX_EXinst__n0030),
    .ADR1(DLX_EXinst__n0016[2]),
    .ADR2(N126816),
    .ADR3(DLX_EXinst__n0128),
    .O(\N126816/GROM )
  );
  X_BUF \N126816/XUSED  (
    .I(\N126816/FROM ),
    .O(N126816)
  );
  X_BUF \N126816/YUSED  (
    .I(\N126816/GROM ),
    .O(CHOICE5567)
  );
  defparam \DLX_IDinst__n0117<22>29 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst__n0117<22>29  (
    .ADR0(CHOICE2386),
    .ADR1(N101161),
    .ADR2(DLX_IDinst_N69914),
    .ADR3(DLX_IDinst_regA_eff[22]),
    .O(\DLX_IDinst_reg_out_A<22>/FROM )
  );
  defparam \DLX_IDinst__n0117<22>39 .INIT = 16'hFFA0;
  X_LUT4 \DLX_IDinst__n0117<22>39  (
    .ADR0(DLX_IDinst__n0310),
    .ADR1(VCC),
    .ADR2(DLX_IFinst_NPC[22]),
    .ADR3(CHOICE2389),
    .O(N104100)
  );
  X_BUF \DLX_IDinst_reg_out_A<22>/XUSED  (
    .I(\DLX_IDinst_reg_out_A<22>/FROM ),
    .O(CHOICE2389)
  );
  defparam \DLX_IDinst__n0117<14>29 .INIT = 16'hECA0;
  X_LUT4 \DLX_IDinst__n0117<14>29  (
    .ADR0(N101161),
    .ADR1(DLX_IDinst_regA_eff[14]),
    .ADR2(CHOICE2302),
    .ADR3(DLX_IDinst_N69914),
    .O(\DLX_IDinst_reg_out_A<14>/FROM )
  );
  defparam \DLX_IDinst__n0117<14>39 .INIT = 16'hFF88;
  X_LUT4 \DLX_IDinst__n0117<14>39  (
    .ADR0(DLX_IFinst_NPC[14]),
    .ADR1(DLX_IDinst__n0310),
    .ADR2(VCC),
    .ADR3(CHOICE2305),
    .O(N103624)
  );
  X_BUF \DLX_IDinst_reg_out_A<14>/XUSED  (
    .I(\DLX_IDinst_reg_out_A<14>/FROM ),
    .O(CHOICE2305)
  );
  defparam \DLX_IDinst__n0117<30>29 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst__n0117<30>29  (
    .ADR0(DLX_IDinst_regA_eff[30]),
    .ADR1(DLX_IDinst_N69914),
    .ADR2(CHOICE2494),
    .ADR3(N101161),
    .O(\DLX_IDinst_reg_out_A<30>/FROM )
  );
  defparam \DLX_IDinst__n0117<30>39 .INIT = 16'hFF88;
  X_LUT4 \DLX_IDinst__n0117<30>39  (
    .ADR0(DLX_IDinst__n0310),
    .ADR1(DLX_IFinst_NPC[30]),
    .ADR2(VCC),
    .ADR3(CHOICE2497),
    .O(N104712)
  );
  X_BUF \DLX_IDinst_reg_out_A<30>/XUSED  (
    .I(\DLX_IDinst_reg_out_A<30>/FROM ),
    .O(CHOICE2497)
  );
  defparam DLX_EXinst_Ker629641.INIT = 16'hACAC;
  X_LUT4 DLX_EXinst_Ker629641 (
    .ADR0(\DLX_EXinst_Mshift__n0023_Sh[29] ),
    .ADR1(\DLX_EXinst_Mshift__n0026_Sh[21] ),
    .ADR2(DLX_IDinst_reg_out_B[3]),
    .ADR3(VCC),
    .O(\DLX_EXinst_N62966/FROM )
  );
  defparam DLX_EXinst_Ker645431.INIT = 16'hCCAA;
  X_LUT4 DLX_EXinst_Ker645431 (
    .ADR0(\DLX_EXinst_Mshift__n0026_Sh[13] ),
    .ADR1(\DLX_EXinst_Mshift__n0026_Sh[21] ),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B_3_1),
    .O(\DLX_EXinst_N62966/GROM )
  );
  X_BUF \DLX_EXinst_N62966/XUSED  (
    .I(\DLX_EXinst_N62966/FROM ),
    .O(DLX_EXinst_N62966)
  );
  X_BUF \DLX_EXinst_N62966/YUSED  (
    .I(\DLX_EXinst_N62966/GROM ),
    .O(DLX_EXinst_N64545)
  );
  defparam DLX_EXinst_Ker634871.INIT = 16'hEE22;
  X_LUT4 DLX_EXinst_Ker634871 (
    .ADR0(DLX_IDinst_reg_out_A[10]),
    .ADR1(DLX_IDinst_IR_function_field[1]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[12]),
    .O(\DLX_EXinst_N63489/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0028_Sh<9>1 .INIT = 16'hEE22;
  X_LUT4 \DLX_EXinst_Mshift__n0028_Sh<9>1  (
    .ADR0(DLX_EXinst_N62981),
    .ADR1(DLX_IDinst_IR_function_field_0_1),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N63489),
    .O(\DLX_EXinst_N63489/GROM )
  );
  X_BUF \DLX_EXinst_N63489/XUSED  (
    .I(\DLX_EXinst_N63489/FROM ),
    .O(DLX_EXinst_N63489)
  );
  X_BUF \DLX_EXinst_N63489/YUSED  (
    .I(\DLX_EXinst_N63489/GROM ),
    .O(\DLX_EXinst_Mshift__n0028_Sh[9] )
  );
  defparam DLX_EXinst_Ker628641.INIT = 16'hFC30;
  X_LUT4 DLX_EXinst_Ker628641 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(DLX_IDinst_reg_out_A[13]),
    .ADR3(DLX_IDinst_reg_out_A[11]),
    .O(\DLX_EXinst_N62866/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0025_Sh<14>1 .INIT = 16'hFC30;
  X_LUT4 \DLX_EXinst_Mshift__n0025_Sh<14>1  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_B[0]),
    .ADR2(DLX_EXinst_N63369),
    .ADR3(DLX_EXinst_N62866),
    .O(\DLX_EXinst_N62866/GROM )
  );
  X_BUF \DLX_EXinst_N62866/XUSED  (
    .I(\DLX_EXinst_N62866/FROM ),
    .O(DLX_EXinst_N62866)
  );
  X_BUF \DLX_EXinst_N62866/YUSED  (
    .I(\DLX_EXinst_N62866/GROM ),
    .O(\DLX_EXinst_Mshift__n0025_Sh[14] )
  );
  defparam DLX_EXinst_Ker627841.INIT = 16'hFA50;
  X_LUT4 DLX_EXinst_Ker627841 (
    .ADR0(DLX_IDinst_IR_function_field[1]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[15]),
    .ADR3(DLX_IDinst_reg_out_A[13]),
    .O(\DLX_EXinst_N62786/FROM )
  );
  defparam DLX_EXinst_Ker64917_SW0.INIT = 16'hFC30;
  X_LUT4 DLX_EXinst_Ker64917_SW0 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_IR_function_field[0]),
    .ADR2(DLX_EXinst_N63454),
    .ADR3(DLX_EXinst_N62786),
    .O(\DLX_EXinst_N62786/GROM )
  );
  X_BUF \DLX_EXinst_N62786/XUSED  (
    .I(\DLX_EXinst_N62786/FROM ),
    .O(DLX_EXinst_N62786)
  );
  X_BUF \DLX_EXinst_N62786/YUSED  (
    .I(\DLX_EXinst_N62786/GROM ),
    .O(N93179)
  );
  defparam \DLX_EXinst_Mshift__n0027_Sh<5>10 .INIT = 16'hE040;
  X_LUT4 \DLX_EXinst_Mshift__n0027_Sh<5>10  (
    .ADR0(DLX_IDinst_IR_function_field_1_1),
    .ADR1(DLX_IDinst_reg_out_A[4]),
    .ADR2(DLX_IDinst_IR_function_field_0_1),
    .ADR3(DLX_IDinst_reg_out_A[2]),
    .O(\CHOICE1018/FROM )
  );
  defparam DLX_EXinst_Ker644721.INIT = 16'hFA0A;
  X_LUT4 DLX_EXinst_Ker644721 (
    .ADR0(DLX_IDinst_reg_out_A[2]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_IR_function_field_1_1),
    .ADR3(DLX_IDinst_reg_out_A[4]),
    .O(\CHOICE1018/GROM )
  );
  X_BUF \CHOICE1018/XUSED  (
    .I(\CHOICE1018/FROM ),
    .O(CHOICE1018)
  );
  X_BUF \CHOICE1018/YUSED  (
    .I(\CHOICE1018/GROM ),
    .O(DLX_EXinst_N64474)
  );
  defparam DLX_EXinst_Ker64912.INIT = 16'hEE44;
  X_LUT4 DLX_EXinst_Ker64912 (
    .ADR0(DLX_IDinst_reg_out_B_3_1),
    .ADR1(N93435),
    .ADR2(VCC),
    .ADR3(\DLX_EXinst_Mshift__n0025_Sh[8] ),
    .O(\DLX_EXinst_N64914/FROM )
  );
  defparam DLX_EXinst_Ker645281.INIT = 16'hD8D8;
  X_LUT4 DLX_EXinst_Ker645281 (
    .ADR0(DLX_IDinst_reg_out_B_3_1),
    .ADR1(\DLX_EXinst_Mshift__n0026_Sh[22] ),
    .ADR2(\DLX_EXinst_Mshift__n0026_Sh[14] ),
    .ADR3(VCC),
    .O(\DLX_EXinst_N64914/GROM )
  );
  X_BUF \DLX_EXinst_N64914/XUSED  (
    .I(\DLX_EXinst_N64914/FROM ),
    .O(DLX_EXinst_N64914)
  );
  X_BUF \DLX_EXinst_N64914/YUSED  (
    .I(\DLX_EXinst_N64914/GROM ),
    .O(DLX_EXinst_N64530)
  );
  defparam DLX_IFinst_NPC_15_1_1162.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_15_1_1162 (
    .I(\NPC_eff<15>/OD ),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\NPC_eff<15>/OFF/RST ),
    .O(DLX_IFinst_NPC_15_1)
  );
  X_OR2 \NPC_eff<15>/OFF/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\NPC_eff<15>/OFF/RST )
  );
  defparam DLX_EXinst_Ker661281.INIT = 16'h0050;
  X_LUT4 DLX_EXinst_Ker661281 (
    .ADR0(DLX_IDinst_IR_opcode_field[4]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_IR_opcode_field[5]),
    .ADR3(DLX_IDinst_IR_opcode_field[1]),
    .O(\DLX_EXinst_N66130/FROM )
  );
  defparam DLX_EXinst__n01471.INIT = 16'h0A00;
  X_LUT4 DLX_EXinst__n01471 (
    .ADR0(DLX_IDinst_IR_opcode_field[3]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_IR_opcode_field[2]),
    .ADR3(DLX_EXinst_N66130),
    .O(\DLX_EXinst_N66130/GROM )
  );
  X_BUF \DLX_EXinst_N66130/XUSED  (
    .I(\DLX_EXinst_N66130/FROM ),
    .O(DLX_EXinst_N66130)
  );
  X_BUF \DLX_EXinst_N66130/YUSED  (
    .I(\DLX_EXinst_N66130/GROM ),
    .O(DLX_EXinst__n0147)
  );
  defparam DLX_IDinst_Mmux__n0148_inst_lut3_1081.INIT = 16'hCFC0;
  X_LUT4 DLX_IDinst_Mmux__n0148_inst_lut3_1081 (
    .ADR0(VCC),
    .ADR1(DLX_MEMinst_RF_data_in[15]),
    .ADR2(DLX_opcode_of_WB[0]),
    .ADR3(DLX_RF_data_in[7]),
    .O(\DLX_IDinst_Mmux__n0148__net123/GROM )
  );
  X_BUF \DLX_IDinst_Mmux__n0148__net123/YUSED  (
    .I(\DLX_IDinst_Mmux__n0148__net123/GROM ),
    .O(DLX_IDinst_Mmux__n0148__net123)
  );
  defparam \DLX_EXinst__n0006<0>36_SW0 .INIT = 16'hAFA0;
  X_LUT4 \DLX_EXinst__n0006<0>36_SW0  (
    .ADR0(DLX_IDinst_reg_out_A[2]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[1]),
    .ADR3(DLX_IDinst_reg_out_A[0]),
    .O(\N126134/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0025_Sh<3>11 .INIT = 16'hE020;
  X_LUT4 \DLX_EXinst_Mshift__n0025_Sh<3>11  (
    .ADR0(DLX_IDinst_reg_out_A[2]),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(DLX_IDinst_reg_out_B[0]),
    .ADR3(DLX_IDinst_reg_out_A[0]),
    .O(\N126134/GROM )
  );
  X_BUF \N126134/XUSED  (
    .I(\N126134/FROM ),
    .O(N126134)
  );
  X_BUF \N126134/YUSED  (
    .I(\N126134/GROM ),
    .O(CHOICE1054)
  );
  defparam DLX_IFlc_md_mda39_a1.INIT = 16'h2222;
  X_LUT4 DLX_IFlc_md_mda39_a1 (
    .ADR0(DLX_IFlc_md_wint38),
    .ADR1(DLX_IFlc_pd_wint1),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IFlc_md_wint39/FROM )
  );
  defparam DLX_IFlc_md_mda4_a1.INIT = 16'h00CC;
  X_LUT4 DLX_IFlc_md_mda4_a1 (
    .ADR0(VCC),
    .ADR1(DLX_IFlc_md_wint3),
    .ADR2(VCC),
    .ADR3(DLX_IFlc_pd_wint1),
    .O(\DLX_IFlc_md_wint39/GROM )
  );
  X_BUF \DLX_IFlc_md_wint39/XUSED  (
    .I(\DLX_IFlc_md_wint39/FROM ),
    .O(DLX_IFlc_md_wint39)
  );
  X_BUF \DLX_IFlc_md_wint39/YUSED  (
    .I(\DLX_IFlc_md_wint39/GROM ),
    .O(DLX_IFlc_md_wint4)
  );
  defparam DLX_EXinst_Ker628491.INIT = 16'hB8B8;
  X_LUT4 DLX_EXinst_Ker628491 (
    .ADR0(DLX_IDinst_reg_out_A[5]),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(DLX_IDinst_reg_out_A[7]),
    .ADR3(VCC),
    .O(\DLX_EXinst_N62851/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0025_Sh<8>1 .INIT = 16'hEE22;
  X_LUT4 \DLX_EXinst_Mshift__n0025_Sh<8>1  (
    .ADR0(DLX_EXinst_N63404),
    .ADR1(DLX_IDinst_reg_out_B[0]),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N62851),
    .O(\DLX_EXinst_N62851/GROM )
  );
  X_BUF \DLX_EXinst_N62851/XUSED  (
    .I(\DLX_EXinst_N62851/FROM ),
    .O(DLX_EXinst_N62851)
  );
  X_BUF \DLX_EXinst_N62851/YUSED  (
    .I(\DLX_EXinst_N62851/GROM ),
    .O(\DLX_EXinst_Mshift__n0025_Sh[8] )
  );
  defparam DLX_EXinst_Ker637831.INIT = 16'hAAF0;
  X_LUT4 DLX_EXinst_Ker637831 (
    .ADR0(DLX_IDinst_reg_out_A[9]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[7]),
    .ADR3(DLX_IDinst_reg_out_B[1]),
    .O(\DLX_EXinst_N63785/FROM )
  );
  defparam DLX_EXinst_Ker627691.INIT = 16'hF0AA;
  X_LUT4 DLX_EXinst_Ker627691 (
    .ADR0(DLX_IDinst_reg_out_A[9]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[7]),
    .ADR3(DLX_IDinst_IR_function_field[1]),
    .O(\DLX_EXinst_N63785/GROM )
  );
  X_BUF \DLX_EXinst_N63785/XUSED  (
    .I(\DLX_EXinst_N63785/FROM ),
    .O(DLX_EXinst_N63785)
  );
  X_BUF \DLX_EXinst_N63785/YUSED  (
    .I(\DLX_EXinst_N63785/GROM ),
    .O(DLX_EXinst_N62771)
  );
  defparam DLX_EXinst_Ker634971.INIT = 16'hFA0A;
  X_LUT4 DLX_EXinst_Ker634971 (
    .ADR0(DLX_IDinst_reg_out_A[14]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_IR_function_field_1_1),
    .ADR3(DLX_IDinst_reg_out_A[16]),
    .O(\DLX_EXinst_N63499/FROM )
  );
  defparam DLX_EXinst_Ker64558_SW0.INIT = 16'hEE44;
  X_LUT4 DLX_EXinst_Ker64558_SW0 (
    .ADR0(DLX_IDinst_IR_function_field[0]),
    .ADR1(DLX_EXinst_N62991),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N63499),
    .O(\DLX_EXinst_N63499/GROM )
  );
  X_BUF \DLX_EXinst_N63499/XUSED  (
    .I(\DLX_EXinst_N63499/FROM ),
    .O(DLX_EXinst_N63499)
  );
  X_BUF \DLX_EXinst_N63499/YUSED  (
    .I(\DLX_EXinst_N63499/GROM ),
    .O(N93955)
  );
  defparam \DLX_EXinst__n0006<9>21 .INIT = 16'h8C88;
  X_LUT4 \DLX_EXinst__n0006<9>21  (
    .ADR0(DLX_EXinst__n0079),
    .ADR1(DLX_IDinst_reg_out_A[9]),
    .ADR2(\DLX_IDinst_Imm[9] ),
    .ADR3(DLX_EXinst__n0080),
    .O(\CHOICE4554/FROM )
  );
  defparam \DLX_EXinst__n0006<3>29 .INIT = 16'hC0E0;
  X_LUT4 \DLX_EXinst__n0006<3>29  (
    .ADR0(DLX_EXinst__n0080),
    .ADR1(DLX_EXinst__n0079),
    .ADR2(DLX_IDinst_reg_out_A[3]),
    .ADR3(DLX_IDinst_IR_function_field[3]),
    .O(\CHOICE4554/GROM )
  );
  X_BUF \CHOICE4554/XUSED  (
    .I(\CHOICE4554/FROM ),
    .O(CHOICE4554)
  );
  X_BUF \CHOICE4554/YUSED  (
    .I(\CHOICE4554/GROM ),
    .O(CHOICE5026)
  );
  defparam \DLX_EXinst__n0006<4>13 .INIT = 16'h88C0;
  X_LUT4 \DLX_EXinst__n0006<4>13  (
    .ADR0(DLX_EXinst_N65105),
    .ADR1(DLX_EXinst_N63185),
    .ADR2(N97593),
    .ADR3(DLX_IDinst_IR_function_field[2]),
    .O(\CHOICE3978/FROM )
  );
  defparam \DLX_EXinst__n0006<4>25 .INIT = 16'hFFF8;
  X_LUT4 \DLX_EXinst__n0006<4>25  (
    .ADR0(DLX_IDinst_reg_out_A[4]),
    .ADR1(DLX_EXinst__n0080),
    .ADR2(DLX_EXinst_N66152),
    .ADR3(CHOICE3978),
    .O(\CHOICE3978/GROM )
  );
  X_BUF \CHOICE3978/XUSED  (
    .I(\CHOICE3978/FROM ),
    .O(CHOICE3978)
  );
  X_BUF \CHOICE3978/YUSED  (
    .I(\CHOICE3978/GROM ),
    .O(CHOICE3980)
  );
  defparam vga_top_vga1__n00101.INIT = 16'hFFFA;
  X_LUT4 vga_top_vga1__n00101 (
    .ADR0(vga_top_vga1__n0034),
    .ADR1(VCC),
    .ADR2(vga_top_vga1__n0033),
    .ADR3(vga_top_vga1_helpme),
    .O(\vga_top_vga1__n0010/FROM )
  );
  defparam vga_top_vga1__n0007_1163.INIT = 16'hF4F0;
  X_LUT4 vga_top_vga1__n0007_1163 (
    .ADR0(N100333),
    .ADR1(vga_top_vga1_vcounter[9]),
    .ADR2(vga_top_vga1_helpme),
    .ADR3(vga_top_vga1_N73363),
    .O(\vga_top_vga1__n0010/GROM )
  );
  X_BUF \vga_top_vga1__n0010/XUSED  (
    .I(\vga_top_vga1__n0010/FROM ),
    .O(vga_top_vga1__n0010)
  );
  X_BUF \vga_top_vga1__n0010/YUSED  (
    .I(\vga_top_vga1__n0010/GROM ),
    .O(vga_top_vga1__n0007)
  );
  defparam DLX_EXinst_Ker628741.INIT = 16'hBB88;
  X_LUT4 DLX_EXinst_Ker628741 (
    .ADR0(DLX_IDinst_reg_out_A[15]),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[17]),
    .O(\DLX_EXinst_N62876/FROM )
  );
  defparam DLX_EXinst_Ker63913_SW0.INIT = 16'hFA0A;
  X_LUT4 DLX_EXinst_Ker63913_SW0 (
    .ADR0(DLX_EXinst_N63379),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[0]),
    .ADR3(DLX_EXinst_N62876),
    .O(\DLX_EXinst_N62876/GROM )
  );
  X_BUF \DLX_EXinst_N62876/XUSED  (
    .I(\DLX_EXinst_N62876/FROM ),
    .O(DLX_EXinst_N62876)
  );
  X_BUF \DLX_EXinst_N62876/YUSED  (
    .I(\DLX_EXinst_N62876/GROM ),
    .O(N93537)
  );
  defparam DLX_EXinst_Ker627941.INIT = 16'hE2E2;
  X_LUT4 DLX_EXinst_Ker627941 (
    .ADR0(DLX_IDinst_reg_out_A[19]),
    .ADR1(DLX_IDinst_IR_function_field[1]),
    .ADR2(DLX_IDinst_reg_out_A[17]),
    .ADR3(VCC),
    .O(\DLX_EXinst_N62796/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0027_Sh<20>1 .INIT = 16'hFA0A;
  X_LUT4 \DLX_EXinst_Mshift__n0027_Sh<20>1  (
    .ADR0(DLX_EXinst_N63464),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_IR_function_field_0_1),
    .ADR3(DLX_EXinst_N62796),
    .O(\DLX_EXinst_N62796/GROM )
  );
  X_BUF \DLX_EXinst_N62796/XUSED  (
    .I(\DLX_EXinst_N62796/FROM ),
    .O(DLX_EXinst_N62796)
  );
  X_BUF \DLX_EXinst_N62796/YUSED  (
    .I(\DLX_EXinst_N62796/GROM ),
    .O(\DLX_EXinst_Mshift__n0027_Sh[20] )
  );
  defparam DLX_EXinst_Ker6538947.INIT = 16'h0088;
  X_LUT4 DLX_EXinst_Ker6538947 (
    .ADR0(DLX_EXinst_N63294),
    .ADR1(DLX_EXinst_N66507),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_IR_function_field_3_1),
    .O(\CHOICE1364/FROM )
  );
  defparam DLX_EXinst_Ker650981.INIT = 16'hB8B8;
  X_LUT4 DLX_EXinst_Ker650981 (
    .ADR0(\DLX_EXinst_Mshift__n0028_Sh[19] ),
    .ADR1(DLX_IDinst_IR_function_field_3_1),
    .ADR2(\DLX_EXinst_Mshift__n0028_Sh[11] ),
    .ADR3(VCC),
    .O(\CHOICE1364/GROM )
  );
  X_BUF \CHOICE1364/XUSED  (
    .I(\CHOICE1364/FROM ),
    .O(CHOICE1364)
  );
  X_BUF \CHOICE1364/YUSED  (
    .I(\CHOICE1364/GROM ),
    .O(DLX_EXinst_N65100)
  );
  defparam \DLX_EXinst__n0006<9>62 .INIT = 16'h8000;
  X_LUT4 \DLX_EXinst__n0006<9>62  (
    .ADR0(CHOICE3377),
    .ADR1(CHOICE3408),
    .ADR2(DLX_IDinst_IR_function_field[4]),
    .ADR3(N101839),
    .O(\CHOICE4567/FROM )
  );
  defparam DLX_EXinst_Ker660581.INIT = 16'hA000;
  X_LUT4 DLX_EXinst_Ker660581 (
    .ADR0(CHOICE3377),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_IR_function_field[4]),
    .ADR3(CHOICE3408),
    .O(\CHOICE4567/GROM )
  );
  X_BUF \CHOICE4567/XUSED  (
    .I(\CHOICE4567/FROM ),
    .O(CHOICE4567)
  );
  X_BUF \CHOICE4567/YUSED  (
    .I(\CHOICE4567/GROM ),
    .O(DLX_EXinst_N66060)
  );
  defparam \DLX_EXinst__n0017<12>1 .INIT = 16'hAAF0;
  X_LUT4 \DLX_EXinst__n0017<12>1  (
    .ADR0(DLX_IDinst_reg_out_B[12]),
    .ADR1(VCC),
    .ADR2(\DLX_IDinst_Imm[12] ),
    .ADR3(DLX_EXinst__n0030_1),
    .O(\DLX_EXinst__n0017<12>/FROM )
  );
  defparam DLX_EXinst_Ker638341.INIT = 16'hFC30;
  X_LUT4 DLX_EXinst_Ker638341 (
    .ADR0(VCC),
    .ADR1(DLX_EXinst__n0030_1),
    .ADR2(DLX_EXinst__n0128),
    .ADR3(DLX_EXinst__n0114),
    .O(\DLX_EXinst__n0017<12>/GROM )
  );
  X_BUF \DLX_EXinst__n0017<12>/XUSED  (
    .I(\DLX_EXinst__n0017<12>/FROM ),
    .O(DLX_EXinst__n0017[12])
  );
  X_BUF \DLX_EXinst__n0017<12>/YUSED  (
    .I(\DLX_EXinst__n0017<12>/GROM ),
    .O(DLX_EXinst_N63836)
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<29>1 .INIT = 16'h30AA;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<29>1  (
    .ADR0(DLX_MEMinst_RF_data_in[29]),
    .ADR1(DLX_opcode_of_WB[2]),
    .ADR2(DLX_IDinst_Mmux__n0148__net123),
    .ADR3(DLX_IDinst__n0147),
    .O(\DLX_IDinst_WB_data_eff<29>/FROM )
  );
  defparam \DLX_IDinst_regB_eff<29>1 .INIT = 16'hEAC0;
  X_LUT4 \DLX_IDinst_regB_eff<29>1  (
    .ADR0(DLX_IDinst_N70716),
    .ADR1(DLX_MEMinst_RF_data_in[29]),
    .ADR2(DLX_IDinst__n0145),
    .ADR3(DLX_IDinst_reg_out_B_RF[29]),
    .O(\DLX_IDinst_WB_data_eff<29>/GROM )
  );
  X_BUF \DLX_IDinst_WB_data_eff<29>/XUSED  (
    .I(\DLX_IDinst_WB_data_eff<29>/FROM ),
    .O(DLX_IDinst_WB_data_eff[29])
  );
  X_BUF \DLX_IDinst_WB_data_eff<29>/YUSED  (
    .I(\DLX_IDinst_WB_data_eff<29>/GROM ),
    .O(DLX_IDinst_regB_eff[29])
  );
  defparam DLX_EXinst_Ker628591.INIT = 16'hCCAA;
  X_LUT4 DLX_EXinst_Ker628591 (
    .ADR0(DLX_IDinst_reg_out_A[11]),
    .ADR1(DLX_IDinst_reg_out_A[9]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[1]),
    .O(\DLX_EXinst_N62861/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0025_Sh<12>1 .INIT = 16'hFC0C;
  X_LUT4 \DLX_EXinst_Mshift__n0025_Sh<12>1  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N63364),
    .ADR2(DLX_IDinst_reg_out_B[0]),
    .ADR3(DLX_EXinst_N62861),
    .O(\DLX_EXinst_N62861/GROM )
  );
  X_BUF \DLX_EXinst_N62861/XUSED  (
    .I(\DLX_EXinst_N62861/FROM ),
    .O(DLX_EXinst_N62861)
  );
  X_BUF \DLX_EXinst_N62861/YUSED  (
    .I(\DLX_EXinst_N62861/GROM ),
    .O(\DLX_EXinst_Mshift__n0025_Sh[12] )
  );
  defparam \DLX_EXinst__n0006<11>59_SW0 .INIT = 16'h0055;
  X_LUT4 \DLX_EXinst__n0006<11>59_SW0  (
    .ADR0(DLX_IDinst_reg_out_A[11]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_IR_opcode_field[0]),
    .O(\N127334/FROM )
  );
  defparam DLX_EXinst_Ker627791.INIT = 16'hACAC;
  X_LUT4 DLX_EXinst_Ker627791 (
    .ADR0(DLX_IDinst_reg_out_A[11]),
    .ADR1(DLX_IDinst_reg_out_A[13]),
    .ADR2(DLX_IDinst_IR_function_field[1]),
    .ADR3(VCC),
    .O(\N127334/GROM )
  );
  X_BUF \N127334/XUSED  (
    .I(\N127334/FROM ),
    .O(N127334)
  );
  X_BUF \N127334/YUSED  (
    .I(\N127334/GROM ),
    .O(DLX_EXinst_N62781)
  );
  defparam \DLX_EXinst__n0006<28>166 .INIT = 16'hCC0A;
  X_LUT4 \DLX_EXinst__n0006<28>166  (
    .ADR0(DLX_IDinst_reg_out_A[28]),
    .ADR1(\DLX_EXinst_Mshift__n0025_Sh[20] ),
    .ADR2(DLX_EXinst_N63157),
    .ADR3(DLX_IDinst_reg_out_B[3]),
    .O(\CHOICE5216/FROM )
  );
  defparam DLX_EXinst_Ker639231.INIT = 16'hE2E2;
  X_LUT4 DLX_EXinst_Ker639231 (
    .ADR0(\DLX_EXinst_Mshift__n0025_Sh[20] ),
    .ADR1(DLX_IDinst_reg_out_B[3]),
    .ADR2(\DLX_EXinst_Mshift__n0025_Sh[12] ),
    .ADR3(VCC),
    .O(\CHOICE5216/GROM )
  );
  X_BUF \CHOICE5216/XUSED  (
    .I(\CHOICE5216/FROM ),
    .O(CHOICE5216)
  );
  X_BUF \CHOICE5216/YUSED  (
    .I(\CHOICE5216/GROM ),
    .O(DLX_EXinst_N63925)
  );
  defparam DLX_EXinst_Ker645631.INIT = 16'hAAF0;
  X_LUT4 DLX_EXinst_Ker645631 (
    .ADR0(\DLX_EXinst_Mshift__n0028_Sh[24] ),
    .ADR1(VCC),
    .ADR2(\DLX_EXinst_Mshift__n0028_Sh[16] ),
    .ADR3(DLX_IDinst_IR_function_field[3]),
    .O(\DLX_EXinst_N64565/FROM )
  );
  defparam \DLX_EXinst__n0006<12>38 .INIT = 16'hE020;
  X_LUT4 \DLX_EXinst__n0006<12>38  (
    .ADR0(N97233),
    .ADR1(DLX_IDinst_IR_function_field[2]),
    .ADR2(DLX_EXinst_N63185),
    .ADR3(DLX_EXinst_N64565),
    .O(\DLX_EXinst_N64565/GROM )
  );
  X_BUF \DLX_EXinst_N64565/XUSED  (
    .I(\DLX_EXinst_N64565/FROM ),
    .O(DLX_EXinst_N64565)
  );
  X_BUF \DLX_EXinst_N64565/YUSED  (
    .I(\DLX_EXinst_N64565/GROM ),
    .O(CHOICE3869)
  );
  defparam DLX_EXinst_reg_out_B_EX_0_1_1164.INIT = 1'b0;
  X_FF DLX_EXinst_reg_out_B_EX_0_1_1164 (
    .I(\DM_write_data<0>/OD ),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DM_write_data<0>/OFF/RST ),
    .O(DLX_EXinst_reg_out_B_EX_0_1)
  );
  X_OR2 \DM_write_data<0>/OFF/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DM_write_data<0>/OFF/RST )
  );
  defparam \DLX_EXinst_Mshift__n0025_Sh<3>25 .INIT = 16'h2230;
  X_LUT4 \DLX_EXinst_Mshift__n0025_Sh<3>25  (
    .ADR0(DLX_IDinst_reg_out_A[1]),
    .ADR1(DLX_IDinst_reg_out_B[0]),
    .ADR2(DLX_IDinst_reg_out_A[3]),
    .ADR3(DLX_IDinst_reg_out_B[1]),
    .O(\CHOICE1060/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0025_Sh<3>28 .INIT = 16'hFFCC;
  X_LUT4 \DLX_EXinst_Mshift__n0025_Sh<3>28  (
    .ADR0(VCC),
    .ADR1(CHOICE1054),
    .ADR2(VCC),
    .ADR3(CHOICE1060),
    .O(\CHOICE1060/GROM )
  );
  X_BUF \CHOICE1060/XUSED  (
    .I(\CHOICE1060/FROM ),
    .O(CHOICE1060)
  );
  X_BUF \CHOICE1060/YUSED  (
    .I(\CHOICE1060/GROM ),
    .O(\DLX_EXinst_Mshift__n0025_Sh[3] )
  );
  defparam DLX_EXinst_Ker628841.INIT = 16'hDD88;
  X_LUT4 DLX_EXinst_Ker628841 (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(DLX_IDinst_reg_out_A[19]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[21]),
    .O(\DLX_EXinst_N62886/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0025_Sh<22>1 .INIT = 16'hFC30;
  X_LUT4 \DLX_EXinst_Mshift__n0025_Sh<22>1  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_B[0]),
    .ADR2(DLX_EXinst_N63389),
    .ADR3(DLX_EXinst_N62886),
    .O(\DLX_EXinst_N62886/GROM )
  );
  X_BUF \DLX_EXinst_N62886/XUSED  (
    .I(\DLX_EXinst_N62886/FROM ),
    .O(DLX_EXinst_N62886)
  );
  X_BUF \DLX_EXinst_N62886/YUSED  (
    .I(\DLX_EXinst_N62886/GROM ),
    .O(\DLX_EXinst_Mshift__n0025_Sh[22] )
  );
  defparam DLX_EXinst_Ker64065.INIT = 16'hDD88;
  X_LUT4 DLX_EXinst_Ker64065 (
    .ADR0(DLX_IDinst_IR_function_field[3]),
    .ADR1(\DLX_EXinst_Mshift__n0027_Sh[10] ),
    .ADR2(VCC),
    .ADR3(N93229),
    .O(\DLX_EXinst_N64067/FROM )
  );
  defparam DLX_EXinst_Ker648121.INIT = 16'hF5A0;
  X_LUT4 DLX_EXinst_Ker648121 (
    .ADR0(DLX_IDinst_IR_function_field[3]),
    .ADR1(VCC),
    .ADR2(\DLX_EXinst_Mshift__n0028_Sh[18] ),
    .ADR3(\DLX_EXinst_Mshift__n0028_Sh[10] ),
    .O(\DLX_EXinst_N64067/GROM )
  );
  X_BUF \DLX_EXinst_N64067/XUSED  (
    .I(\DLX_EXinst_N64067/FROM ),
    .O(DLX_EXinst_N64067)
  );
  X_BUF \DLX_EXinst_N64067/YUSED  (
    .I(\DLX_EXinst_N64067/GROM ),
    .O(DLX_EXinst_N64814)
  );
  defparam DLX_EXinst_Ker660761.INIT = 16'h0C0C;
  X_LUT4 DLX_EXinst_Ker660761 (
    .ADR0(VCC),
    .ADR1(N111221),
    .ADR2(DLX_IDinst_reg_out_B[4]),
    .ADR3(VCC),
    .O(\DLX_EXinst_N66078/FROM )
  );
  defparam \DLX_EXinst__n0006<29>335_SW0 .INIT = 16'hFEEE;
  X_LUT4 \DLX_EXinst__n0006<29>335_SW0  (
    .ADR0(CHOICE5393),
    .ADR1(CHOICE5384),
    .ADR2(DLX_EXinst_N65090),
    .ADR3(DLX_EXinst_N66078),
    .O(\DLX_EXinst_N66078/GROM )
  );
  X_BUF \DLX_EXinst_N66078/XUSED  (
    .I(\DLX_EXinst_N66078/FROM ),
    .O(DLX_EXinst_N66078)
  );
  X_BUF \DLX_EXinst_N66078/YUSED  (
    .I(\DLX_EXinst_N66078/GROM ),
    .O(N126442)
  );
  defparam vga_top_vga1__n0011_SW1.INIT = 16'hEFAF;
  X_LUT4 vga_top_vga1__n0011_SW1 (
    .ADR0(vga_top_vga1_vcounter[5]),
    .ADR1(vga_top_vga1_vcounter[3]),
    .ADR2(vga_top_vga1_N73394),
    .ADR3(vga_top_vga1_vcounter[2]),
    .O(\N127107/FROM )
  );
  defparam vga_top_vga1__n0011_1165.INIT = 16'hF3F7;
  X_LUT4 vga_top_vga1__n0011_1165 (
    .ADR0(vga_top_vga1_vcounter[4]),
    .ADR1(vga_top_vga1_vcounter[9]),
    .ADR2(vga_top_vga1_helpme),
    .ADR3(N127107),
    .O(\N127107/GROM )
  );
  X_BUF \N127107/XUSED  (
    .I(\N127107/FROM ),
    .O(N127107)
  );
  X_BUF \N127107/YUSED  (
    .I(\N127107/GROM ),
    .O(vga_top_vga1__n0011)
  );
  defparam DLX_EXinst_Ker648621.INIT = 16'hEE44;
  X_LUT4 DLX_EXinst_Ker648621 (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(DLX_IDinst_reg_out_A[1]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[3]),
    .O(\DLX_EXinst_N64864/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0025_Sh<4>11 .INIT = 16'hA0C0;
  X_LUT4 \DLX_EXinst_Mshift__n0025_Sh<4>11  (
    .ADR0(DLX_IDinst_reg_out_A[1]),
    .ADR1(DLX_IDinst_reg_out_A[3]),
    .ADR2(DLX_IDinst_reg_out_B[0]),
    .ADR3(DLX_IDinst_reg_out_B[1]),
    .O(\DLX_EXinst_N64864/GROM )
  );
  X_BUF \DLX_EXinst_N64864/XUSED  (
    .I(\DLX_EXinst_N64864/FROM ),
    .O(DLX_EXinst_N64864)
  );
  X_BUF \DLX_EXinst_N64864/YUSED  (
    .I(\DLX_EXinst_N64864/GROM ),
    .O(CHOICE1078)
  );
  defparam DLX_EXinst_Ker629491.INIT = 16'hE2E2;
  X_LUT4 DLX_EXinst_Ker629491 (
    .ADR0(DLX_IDinst_reg_out_A[9]),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(DLX_IDinst_reg_out_A[11]),
    .ADR3(VCC),
    .O(\DLX_EXinst_N62951/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<8>1 .INIT = 16'hFA50;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<8>1  (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N63304),
    .ADR3(DLX_EXinst_N62951),
    .O(\DLX_EXinst_N62951/GROM )
  );
  X_BUF \DLX_EXinst_N62951/XUSED  (
    .I(\DLX_EXinst_N62951/FROM ),
    .O(DLX_EXinst_N62951)
  );
  X_BUF \DLX_EXinst_N62951/YUSED  (
    .I(\DLX_EXinst_N62951/GROM ),
    .O(\DLX_EXinst_Mshift__n0023_Sh[8] )
  );
  defparam DLX_EXinst_Ker628691.INIT = 16'hCCF0;
  X_LUT4 DLX_EXinst_Ker628691 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[13]),
    .ADR2(DLX_IDinst_reg_out_A[15]),
    .ADR3(DLX_IDinst_reg_out_B[1]),
    .O(\DLX_EXinst_N62871/FROM )
  );
  defparam DLX_EXinst_Ker64912_SW0.INIT = 16'hFA0A;
  X_LUT4 DLX_EXinst_Ker64912_SW0 (
    .ADR0(DLX_EXinst_N63374),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[0]),
    .ADR3(DLX_EXinst_N62871),
    .O(\DLX_EXinst_N62871/GROM )
  );
  X_BUF \DLX_EXinst_N62871/XUSED  (
    .I(\DLX_EXinst_N62871/FROM ),
    .O(DLX_EXinst_N62871)
  );
  X_BUF \DLX_EXinst_N62871/YUSED  (
    .I(\DLX_EXinst_N62871/GROM ),
    .O(N93435)
  );
  defparam DLX_EXinst_Ker627891.INIT = 16'hFC0C;
  X_LUT4 DLX_EXinst_Ker627891 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[17]),
    .ADR2(DLX_IDinst_IR_function_field[1]),
    .ADR3(DLX_IDinst_reg_out_A[15]),
    .O(\DLX_EXinst_N62791/FROM )
  );
  defparam DLX_EXinst_Ker6540411.INIT = 16'hC808;
  X_LUT4 DLX_EXinst_Ker6540411 (
    .ADR0(DLX_EXinst_N63459),
    .ADR1(DLX_IDinst_IR_function_field_3_1),
    .ADR2(DLX_IDinst_IR_function_field[0]),
    .ADR3(DLX_EXinst_N62791),
    .O(\DLX_EXinst_N62791/GROM )
  );
  X_BUF \DLX_EXinst_N62791/XUSED  (
    .I(\DLX_EXinst_N62791/FROM ),
    .O(DLX_EXinst_N62791)
  );
  X_BUF \DLX_EXinst_N62791/YUSED  (
    .I(\DLX_EXinst_N62791/GROM ),
    .O(CHOICE1343)
  );
  defparam DLX_EXinst_Ker660851.INIT = 16'h0C00;
  X_LUT4 DLX_EXinst_Ker660851 (
    .ADR0(VCC),
    .ADR1(DLX_EXinst__n0081),
    .ADR2(N109130),
    .ADR3(DLX_IDinst_IR_function_field[4]),
    .O(\DLX_EXinst_N66087/FROM )
  );
  defparam \DLX_EXinst__n0006<17>14 .INIT = 16'h0200;
  X_LUT4 \DLX_EXinst__n0006<17>14  (
    .ADR0(\DLX_EXinst_Mshift__n0027_Sh[1] ),
    .ADR1(DLX_IDinst_IR_function_field[3]),
    .ADR2(DLX_IDinst_IR_function_field[2]),
    .ADR3(DLX_EXinst_N66087),
    .O(\DLX_EXinst_N66087/GROM )
  );
  X_BUF \DLX_EXinst_N66087/XUSED  (
    .I(\DLX_EXinst_N66087/FROM ),
    .O(DLX_EXinst_N66087)
  );
  X_BUF \DLX_EXinst_N66087/YUSED  (
    .I(\DLX_EXinst_N66087/GROM ),
    .O(CHOICE5577)
  );
  defparam DLX_EXinst_Ker649021.INIT = 16'hCCF0;
  X_LUT4 DLX_EXinst_Ker649021 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[5]),
    .ADR2(DLX_IDinst_reg_out_A[3]),
    .ADR3(DLX_IDinst_reg_out_B[1]),
    .O(\DLX_EXinst_N64904/FROM )
  );
  defparam \DLX_EXinst__n0006<3>227 .INIT = 16'h0B08;
  X_LUT4 \DLX_EXinst__n0006<3>227  (
    .ADR0(DLX_EXinst_N64587),
    .ADR1(DLX_IDinst_reg_out_B[0]),
    .ADR2(DLX_IDinst_reg_out_B[3]),
    .ADR3(DLX_EXinst_N64904),
    .O(\DLX_EXinst_N64904/GROM )
  );
  X_BUF \DLX_EXinst_N64904/XUSED  (
    .I(\DLX_EXinst_N64904/FROM ),
    .O(DLX_EXinst_N64904)
  );
  X_BUF \DLX_EXinst_N64904/YUSED  (
    .I(\DLX_EXinst_N64904/GROM ),
    .O(CHOICE5073)
  );
  defparam DLX_EXinst_Ker628891.INIT = 16'hCCF0;
  X_LUT4 DLX_EXinst_Ker628891 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[21]),
    .ADR2(DLX_IDinst_reg_out_A[23]),
    .ADR3(DLX_IDinst_reg_out_B[1]),
    .O(\DLX_EXinst_N62891/FROM )
  );
  defparam DLX_EXinst_Ker628941.INIT = 16'hCCF0;
  X_LUT4 DLX_EXinst_Ker628941 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[23]),
    .ADR2(DLX_IDinst_reg_out_A[25]),
    .ADR3(DLX_IDinst_reg_out_B[1]),
    .O(\DLX_EXinst_N62891/GROM )
  );
  X_BUF \DLX_EXinst_N62891/XUSED  (
    .I(\DLX_EXinst_N62891/FROM ),
    .O(DLX_EXinst_N62891)
  );
  X_BUF \DLX_EXinst_N62891/YUSED  (
    .I(\DLX_EXinst_N62891/GROM ),
    .O(DLX_EXinst_N62896)
  );
  defparam DLX_EXinst_Ker660941.INIT = 16'h000C;
  X_LUT4 DLX_EXinst_Ker660941 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_IR_function_field_2_1),
    .ADR2(DLX_IDinst_IR_function_field[4]),
    .ADR3(DLX_IDinst_IR_function_field_3_1),
    .O(\DLX_EXinst_N66096/FROM )
  );
  defparam DLX_EXinst__n00451.INIT = 16'h0200;
  X_LUT4 DLX_EXinst__n00451 (
    .ADR0(DLX_IDinst_IR_function_field[5]),
    .ADR1(DLX_IDinst_IR_function_field[1]),
    .ADR2(DLX_IDinst_IR_function_field[0]),
    .ADR3(DLX_EXinst_N66096),
    .O(\DLX_EXinst_N66096/GROM )
  );
  X_BUF \DLX_EXinst_N66096/XUSED  (
    .I(\DLX_EXinst_N66096/FROM ),
    .O(DLX_EXinst_N66096)
  );
  X_BUF \DLX_EXinst_N66096/YUSED  (
    .I(\DLX_EXinst_N66096/GROM ),
    .O(DLX_EXinst__n0045)
  );
  defparam DLX_EXinst_Ker6538920.INIT = 16'h0C00;
  X_LUT4 DLX_EXinst_Ker6538920 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[31]),
    .ADR2(DLX_IDinst_IR_function_field_3_1),
    .ADR3(\DLX_IDinst_Imm[5] ),
    .O(\CHOICE1359/FROM )
  );
  defparam DLX_EXinst_Ker648221.INIT = 16'hFA0A;
  X_LUT4 DLX_EXinst_Ker648221 (
    .ADR0(\DLX_EXinst_Mshift__n0028_Sh[9] ),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_IR_function_field_3_1),
    .ADR3(\DLX_EXinst_Mshift__n0028_Sh[17] ),
    .O(\CHOICE1359/GROM )
  );
  X_BUF \CHOICE1359/XUSED  (
    .I(\CHOICE1359/FROM ),
    .O(CHOICE1359)
  );
  X_BUF \CHOICE1359/YUSED  (
    .I(\CHOICE1359/GROM ),
    .O(DLX_EXinst_N64824)
  );
  defparam DLX_EXinst_Ker63913.INIT = 16'hEE22;
  X_LUT4 DLX_EXinst_Ker63913 (
    .ADR0(N93537),
    .ADR1(DLX_IDinst_reg_out_B[3]),
    .ADR2(VCC),
    .ADR3(\DLX_EXinst_Mshift__n0025_Sh[10] ),
    .O(\DLX_EXinst_N63915/FROM )
  );
  defparam DLX_EXinst_Ker639181.INIT = 16'hEE22;
  X_LUT4 DLX_EXinst_Ker639181 (
    .ADR0(\DLX_EXinst_Mshift__n0025_Sh[19] ),
    .ADR1(DLX_IDinst_reg_out_B[3]),
    .ADR2(VCC),
    .ADR3(\DLX_EXinst_Mshift__n0025_Sh[11] ),
    .O(\DLX_EXinst_N63915/GROM )
  );
  X_BUF \DLX_EXinst_N63915/XUSED  (
    .I(\DLX_EXinst_N63915/FROM ),
    .O(DLX_EXinst_N63915)
  );
  X_BUF \DLX_EXinst_N63915/YUSED  (
    .I(\DLX_EXinst_N63915/GROM ),
    .O(DLX_EXinst_N63920)
  );
  defparam \DLX_EXinst__n0006<10>59 .INIT = 16'h8200;
  X_LUT4 \DLX_EXinst__n0006<10>59  (
    .ADR0(DLX_EXinst_N66105),
    .ADR1(DLX_IDinst_IR_opcode_field[1]),
    .ADR2(N127396),
    .ADR3(\DLX_IDinst_Imm[10] ),
    .O(\CHOICE4504/FROM )
  );
  defparam \DLX_EXinst__n0006<5>16 .INIT = 16'h8020;
  X_LUT4 \DLX_EXinst__n0006<5>16  (
    .ADR0(DLX_EXinst_N66105),
    .ADR1(DLX_IDinst_IR_opcode_field[1]),
    .ADR2(\DLX_IDinst_Imm[5] ),
    .ADR3(N127318),
    .O(\CHOICE4504/GROM )
  );
  X_BUF \CHOICE4504/XUSED  (
    .I(\CHOICE4504/FROM ),
    .O(CHOICE4504)
  );
  X_BUF \CHOICE4504/YUSED  (
    .I(\CHOICE4504/GROM ),
    .O(CHOICE4422)
  );
  defparam DLX_EXinst_Ker628791.INIT = 16'hEE22;
  X_LUT4 DLX_EXinst_Ker628791 (
    .ADR0(DLX_IDinst_reg_out_A[19]),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[17]),
    .O(\DLX_EXinst_N62881/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0025_Sh<20>1 .INIT = 16'hFC30;
  X_LUT4 \DLX_EXinst_Mshift__n0025_Sh<20>1  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_B[0]),
    .ADR2(DLX_EXinst_N63384),
    .ADR3(DLX_EXinst_N62881),
    .O(\DLX_EXinst_N62881/GROM )
  );
  X_BUF \DLX_EXinst_N62881/XUSED  (
    .I(\DLX_EXinst_N62881/FROM ),
    .O(DLX_EXinst_N62881)
  );
  X_BUF \DLX_EXinst_N62881/YUSED  (
    .I(\DLX_EXinst_N62881/GROM ),
    .O(\DLX_EXinst_Mshift__n0025_Sh[20] )
  );
  defparam DLX_EXinst_Ker627991.INIT = 16'hFA0A;
  X_LUT4 DLX_EXinst_Ker627991 (
    .ADR0(DLX_IDinst_reg_out_A[21]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_IR_function_field[1]),
    .ADR3(DLX_IDinst_reg_out_A[19]),
    .O(\DLX_EXinst_N62801/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0027_Sh<22>1 .INIT = 16'hFC30;
  X_LUT4 \DLX_EXinst_Mshift__n0027_Sh<22>1  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_IR_function_field_0_1),
    .ADR2(DLX_EXinst_N63469),
    .ADR3(DLX_EXinst_N62801),
    .O(\DLX_EXinst_N62801/GROM )
  );
  X_BUF \DLX_EXinst_N62801/XUSED  (
    .I(\DLX_EXinst_N62801/FROM ),
    .O(DLX_EXinst_N62801)
  );
  X_BUF \DLX_EXinst_N62801/YUSED  (
    .I(\DLX_EXinst_N62801/GROM ),
    .O(\DLX_EXinst_Mshift__n0027_Sh[22] )
  );
  defparam \DLX_EXinst_Mshift__n0025_Sh<4>25 .INIT = 16'h5410;
  X_LUT4 \DLX_EXinst_Mshift__n0025_Sh<4>25  (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(DLX_IDinst_reg_out_A[4]),
    .ADR3(DLX_IDinst_reg_out_A[2]),
    .O(\CHOICE1084/FROM )
  );
  defparam DLX_EXinst_Ker628991.INIT = 16'hBBB8;
  X_LUT4 DLX_EXinst_Ker628991 (
    .ADR0(\DLX_EXinst_Mshift__n0025_Sh[0] ),
    .ADR1(DLX_IDinst_reg_out_B[2]),
    .ADR2(CHOICE1078),
    .ADR3(CHOICE1084),
    .O(\CHOICE1084/GROM )
  );
  X_BUF \CHOICE1084/XUSED  (
    .I(\CHOICE1084/FROM ),
    .O(CHOICE1084)
  );
  X_BUF \CHOICE1084/YUSED  (
    .I(\CHOICE1084/GROM ),
    .O(DLX_EXinst_N62901)
  );
  defparam DLX_EXinst_Ker629841.INIT = 16'hB8B8;
  X_LUT4 DLX_EXinst_Ker629841 (
    .ADR0(DLX_IDinst_reg_out_A[13]),
    .ADR1(DLX_IDinst_IR_function_field[1]),
    .ADR2(DLX_IDinst_reg_out_A[11]),
    .ADR3(VCC),
    .O(\DLX_EXinst_N62986/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0028_Sh<10>1 .INIT = 16'hFA0A;
  X_LUT4 \DLX_EXinst_Mshift__n0028_Sh<10>1  (
    .ADR0(DLX_EXinst_N63489),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_IR_function_field_0_1),
    .ADR3(DLX_EXinst_N62986),
    .O(\DLX_EXinst_N62986/GROM )
  );
  X_BUF \DLX_EXinst_N62986/XUSED  (
    .I(\DLX_EXinst_N62986/FROM ),
    .O(DLX_EXinst_N62986)
  );
  X_BUF \DLX_EXinst_N62986/YUSED  (
    .I(\DLX_EXinst_N62986/GROM ),
    .O(\DLX_EXinst_Mshift__n0028_Sh[10] )
  );
  defparam \DLX_EXinst__n0006<4>74 .INIT = 16'hEAC0;
  X_LUT4 \DLX_EXinst__n0006<4>74  (
    .ADR0(DLX_IDinst_reg_out_A[4]),
    .ADR1(CHOICE3990),
    .ADR2(DLX_IDinst_IR_function_field[4]),
    .ADR3(DLX_EXinst__n0079),
    .O(\CHOICE3992/FROM )
  );
  defparam \DLX_EXinst__n0006<4>100 .INIT = 16'h0F04;
  X_LUT4 \DLX_EXinst__n0006<4>100  (
    .ADR0(DLX_IDinst_IR_function_field[4]),
    .ADR1(CHOICE3980),
    .ADR2(DLX_EXinst__n0030_1),
    .ADR3(CHOICE3992),
    .O(\CHOICE3992/GROM )
  );
  X_BUF \CHOICE3992/XUSED  (
    .I(\CHOICE3992/FROM ),
    .O(CHOICE3992)
  );
  X_BUF \CHOICE3992/YUSED  (
    .I(\CHOICE3992/GROM ),
    .O(CHOICE3994)
  );
  defparam \DLX_EXinst__n0006<2>117_SW0 .INIT = 16'h0033;
  X_LUT4 \DLX_EXinst__n0006<2>117_SW0  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_IR_opcode_field[0]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[2]),
    .O(\N127306/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0025_Sh<5>10 .INIT = 16'h88A0;
  X_LUT4 \DLX_EXinst_Mshift__n0025_Sh<5>10  (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(DLX_IDinst_reg_out_A[2]),
    .ADR2(DLX_IDinst_reg_out_A[3]),
    .ADR3(DLX_IDinst_reg_out_B[0]),
    .O(\N127306/GROM )
  );
  X_BUF \N127306/XUSED  (
    .I(\N127306/FROM ),
    .O(N127306)
  );
  X_BUF \N127306/YUSED  (
    .I(\N127306/GROM ),
    .O(CHOICE1066)
  );
  defparam DLX_IDinst__n0146153.INIT = 16'hCC00;
  X_LUT4 DLX_IDinst__n0146153 (
    .ADR0(VCC),
    .ADR1(CHOICE3673),
    .ADR2(VCC),
    .ADR3(CHOICE3666),
    .O(\CHOICE3674/FROM )
  );
  defparam DLX_IDinst__n0146182_SW0.INIT = 16'h8000;
  X_LUT4 DLX_IDinst__n0146182_SW0 (
    .ADR0(CHOICE3658),
    .ADR1(CHOICE3642),
    .ADR2(CHOICE3651),
    .ADR3(CHOICE3674),
    .O(\CHOICE3674/GROM )
  );
  X_BUF \CHOICE3674/XUSED  (
    .I(\CHOICE3674/FROM ),
    .O(CHOICE3674)
  );
  X_BUF \CHOICE3674/YUSED  (
    .I(\CHOICE3674/GROM ),
    .O(N126289)
  );
  defparam DLX_EXinst_Ker63710_SW0.INIT = 16'hC000;
  X_LUT4 DLX_EXinst_Ker63710_SW0 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_IR_function_field[0]),
    .ADR2(DLX_IDinst_IR_function_field_1_1),
    .ADR3(DLX_EXinst_N66519),
    .O(\N95300/FROM )
  );
  defparam DLX_EXinst_Ker63710.INIT = 16'hFF80;
  X_LUT4 DLX_EXinst_Ker63710 (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(DLX_IDinst_reg_out_B[0]),
    .ADR2(DLX_EXinst_N66072),
    .ADR3(N95300),
    .O(\N95300/GROM )
  );
  X_BUF \N95300/XUSED  (
    .I(\N95300/FROM ),
    .O(N95300)
  );
  X_BUF \N95300/YUSED  (
    .I(\N95300/GROM ),
    .O(DLX_EXinst_N63712)
  );
  defparam DLX_EXinst_Ker629691.INIT = 16'hCCAA;
  X_LUT4 DLX_EXinst_Ker629691 (
    .ADR0(\DLX_EXinst_Mshift__n0026_Sh[22] ),
    .ADR1(\DLX_EXinst_Mshift__n0023_Sh[30] ),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[3]),
    .O(\DLX_EXinst_N62971/FROM )
  );
  defparam DLX_EXinst_Ker6487252.INIT = 16'h7520;
  X_LUT4 DLX_EXinst_Ker6487252 (
    .ADR0(DLX_IDinst_reg_out_B_2_1),
    .ADR1(DLX_IDinst_reg_out_B_3_1),
    .ADR2(\DLX_EXinst_Mshift__n0023_Sh[26] ),
    .ADR3(DLX_EXinst_N62971),
    .O(\DLX_EXinst_N62971/GROM )
  );
  X_BUF \DLX_EXinst_N62971/XUSED  (
    .I(\DLX_EXinst_N62971/FROM ),
    .O(DLX_EXinst_N62971)
  );
  X_BUF \DLX_EXinst_N62971/YUSED  (
    .I(\DLX_EXinst_N62971/GROM ),
    .O(CHOICE3196)
  );
  defparam DLX_EXinst__n0128_SW0.INIT = 16'h0050;
  X_LUT4 DLX_EXinst__n0128_SW0 (
    .ADR0(DLX_IDinst_IR_opcode_field[2]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_IR_opcode_field[3]),
    .ADR3(DLX_IDinst_IR_opcode_field[5]),
    .O(\N89980/FROM )
  );
  defparam DLX_EXinst_Ker664411.INIT = 16'h00F0;
  X_LUT4 DLX_EXinst_Ker664411 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_IR_opcode_field[3]),
    .ADR3(DLX_IDinst_IR_opcode_field[5]),
    .O(\N89980/GROM )
  );
  X_BUF \N89980/XUSED  (
    .I(\N89980/FROM ),
    .O(N89980)
  );
  X_BUF \N89980/YUSED  (
    .I(\N89980/GROM ),
    .O(DLX_EXinst_N66443)
  );
  defparam \DLX_EXinst_Mshift__n0025_Sh<4>28 .INIT = 16'hFCFC;
  X_LUT4 \DLX_EXinst_Mshift__n0025_Sh<4>28  (
    .ADR0(VCC),
    .ADR1(CHOICE1078),
    .ADR2(CHOICE1084),
    .ADR3(VCC),
    .O(\DLX_EXinst_Mshift__n0025_Sh<4>/FROM )
  );
  defparam \DLX_EXinst__n0006<16>256 .INIT = 16'hA808;
  X_LUT4 \DLX_EXinst__n0006<16>256  (
    .ADR0(DLX_IDinst_reg_out_B[2]),
    .ADR1(\DLX_EXinst_Mshift__n0025_Sh[12] ),
    .ADR2(DLX_IDinst_reg_out_B[3]),
    .ADR3(\DLX_EXinst_Mshift__n0025_Sh[4] ),
    .O(\DLX_EXinst_Mshift__n0025_Sh<4>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0025_Sh<4>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0025_Sh<4>/FROM ),
    .O(\DLX_EXinst_Mshift__n0025_Sh[4] )
  );
  X_BUF \DLX_EXinst_Mshift__n0025_Sh<4>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0025_Sh<4>/GROM ),
    .O(CHOICE5162)
  );
  defparam \DLX_EXinst__n0006<5>38 .INIT = 16'hE020;
  X_LUT4 \DLX_EXinst__n0006<5>38  (
    .ADR0(N96585),
    .ADR1(DLX_IDinst_IR_function_field[2]),
    .ADR2(DLX_EXinst_N63185),
    .ADR3(DLX_EXinst_N64824),
    .O(\CHOICE4429/FROM )
  );
  defparam \DLX_EXinst__n0006<5>80 .INIT = 16'hAFAE;
  X_LUT4 \DLX_EXinst__n0006<5>80  (
    .ADR0(CHOICE4438),
    .ADR1(CHOICE4432),
    .ADR2(DLX_IDinst_IR_function_field[4]),
    .ADR3(CHOICE4429),
    .O(\CHOICE4429/GROM )
  );
  X_BUF \CHOICE4429/XUSED  (
    .I(\CHOICE4429/FROM ),
    .O(CHOICE4429)
  );
  X_BUF \CHOICE4429/YUSED  (
    .I(\CHOICE4429/GROM ),
    .O(CHOICE4439)
  );
  defparam DLX_EXinst_Ker629941.INIT = 16'hAACC;
  X_LUT4 DLX_EXinst_Ker629941 (
    .ADR0(DLX_IDinst_reg_out_A[17]),
    .ADR1(DLX_IDinst_reg_out_A[15]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_IR_function_field[1]),
    .O(\DLX_EXinst_N62996/FROM )
  );
  defparam DLX_EXinst_Ker64548_SW0.INIT = 16'hEE22;
  X_LUT4 DLX_EXinst_Ker64548_SW0 (
    .ADR0(DLX_EXinst_N63499),
    .ADR1(DLX_IDinst_IR_function_field[0]),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N62996),
    .O(\DLX_EXinst_N62996/GROM )
  );
  X_BUF \DLX_EXinst_N62996/XUSED  (
    .I(\DLX_EXinst_N62996/FROM ),
    .O(DLX_EXinst_N62996)
  );
  X_BUF \DLX_EXinst_N62996/YUSED  (
    .I(\DLX_EXinst_N62996/GROM ),
    .O(N93905)
  );
  defparam \DLX_EXinst__n0006<21>312_SW0 .INIT = 16'h3332;
  X_LUT4 \DLX_EXinst__n0006<21>312_SW0  (
    .ADR0(CHOICE4189),
    .ADR1(DLX_EXinst__n0030),
    .ADR2(CHOICE4164),
    .ADR3(CHOICE4175),
    .O(\DLX_EXinst_ALU_result<21>/FROM )
  );
  defparam \DLX_EXinst__n0006<21>312 .INIT = 16'hCCC8;
  X_LUT4 \DLX_EXinst__n0006<21>312  (
    .ADR0(N100490),
    .ADR1(DLX_EXinst__n0149),
    .ADR2(CHOICE4223),
    .ADR3(N126415),
    .O(N114850)
  );
  X_BUF \DLX_EXinst_ALU_result<21>/XUSED  (
    .I(\DLX_EXinst_ALU_result<21>/FROM ),
    .O(N126415)
  );
  defparam DLX_IDinst__n0146182.INIT = 16'h8000;
  X_LUT4 DLX_IDinst__n0146182 (
    .ADR0(CHOICE3620),
    .ADR1(N126289),
    .ADR2(CHOICE3635),
    .ADR3(CHOICE3627),
    .O(\DLX_IDinst_zflag/FROM )
  );
  defparam DLX_IDinst_Ker7066629.INIT = 16'h1144;
  X_LUT4 DLX_IDinst_Ker7066629 (
    .ADR0(DLX_IFinst_IR_latched[30]),
    .ADR1(DLX_IFinst_IR_latched[26]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_zflag),
    .O(\DLX_IDinst_zflag/GROM )
  );
  X_BUF \DLX_IDinst_zflag/XUSED  (
    .I(\DLX_IDinst_zflag/FROM ),
    .O(DLX_IDinst_zflag)
  );
  X_BUF \DLX_IDinst_zflag/YUSED  (
    .I(\DLX_IDinst_zflag/GROM ),
    .O(CHOICE3267)
  );
  defparam DLX_EXinst__n00821.INIT = 16'h0088;
  X_LUT4 DLX_EXinst__n00821 (
    .ADR0(DLX_EXinst_N66112),
    .ADR1(DLX_IDinst_IR_opcode_field[1]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_IR_opcode_field[0]),
    .O(\DLX_EXinst__n0082/FROM )
  );
  defparam DLX_EXinst_Ker663711.INIT = 16'h0800;
  X_LUT4 DLX_EXinst_Ker663711 (
    .ADR0(DLX_EXinst_N66112),
    .ADR1(DLX_IDinst_IR_opcode_field[1]),
    .ADR2(DLX_IDinst_IR_opcode_field[0]),
    .ADR3(DLX_IDinst_IR_function_field[4]),
    .O(\DLX_EXinst__n0082/GROM )
  );
  X_BUF \DLX_EXinst__n0082/XUSED  (
    .I(\DLX_EXinst__n0082/FROM ),
    .O(DLX_EXinst__n0082)
  );
  X_BUF \DLX_EXinst__n0082/YUSED  (
    .I(\DLX_EXinst__n0082/GROM ),
    .O(DLX_EXinst_N66373)
  );
  defparam DLX_EXinst_Ker629791.INIT = 16'hD8D8;
  X_LUT4 DLX_EXinst_Ker629791 (
    .ADR0(DLX_IDinst_IR_function_field[1]),
    .ADR1(DLX_IDinst_reg_out_A[11]),
    .ADR2(DLX_IDinst_reg_out_A[9]),
    .ADR3(VCC),
    .O(\DLX_EXinst_N62981/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0028_Sh<8>1 .INIT = 16'hFA50;
  X_LUT4 \DLX_EXinst_Mshift__n0028_Sh<8>1  (
    .ADR0(DLX_IDinst_IR_function_field_0_1),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N63339),
    .ADR3(DLX_EXinst_N62981),
    .O(\DLX_EXinst_N62981/GROM )
  );
  X_BUF \DLX_EXinst_N62981/XUSED  (
    .I(\DLX_EXinst_N62981/FROM ),
    .O(DLX_EXinst_N62981)
  );
  X_BUF \DLX_EXinst_N62981/YUSED  (
    .I(\DLX_EXinst_N62981/GROM ),
    .O(\DLX_EXinst_Mshift__n0028_Sh[8] )
  );
  defparam DLX_EXinst_Ker664191.INIT = 16'h0D08;
  X_LUT4 DLX_EXinst_Ker664191 (
    .ADR0(DLX_IDinst_IR_function_field_0_1),
    .ADR1(DLX_EXinst_N63279),
    .ADR2(DLX_IDinst_IR_function_field_3_1),
    .ADR3(DLX_EXinst_N63016),
    .O(\DLX_EXinst_N66421/FROM )
  );
  defparam DLX_EXinst_Ker630291.INIT = 16'hFF08;
  X_LUT4 DLX_EXinst_Ker630291 (
    .ADR0(DLX_IDinst_IR_function_field[3]),
    .ADR1(DLX_IDinst_reg_out_A[31]),
    .ADR2(DLX_EXinst_N63129),
    .ADR3(DLX_EXinst_N66421),
    .O(\DLX_EXinst_N66421/GROM )
  );
  X_BUF \DLX_EXinst_N66421/XUSED  (
    .I(\DLX_EXinst_N66421/FROM ),
    .O(DLX_EXinst_N66421)
  );
  X_BUF \DLX_EXinst_N66421/YUSED  (
    .I(\DLX_EXinst_N66421/GROM ),
    .O(DLX_EXinst_N63031)
  );
  defparam DLX_EXinst_Ker665231.INIT = 16'h0002;
  X_LUT4 DLX_EXinst_Ker665231 (
    .ADR0(DLX_EXinst_N66112),
    .ADR1(DLX_IDinst_IR_opcode_field[1]),
    .ADR2(DLX_IDinst_IR_opcode_field[0]),
    .ADR3(DLX_IDinst_IR_function_field[4]),
    .O(\DLX_EXinst_N66525/FROM )
  );
  defparam \DLX_EXinst__n0006<15>6 .INIT = 16'hECA0;
  X_LUT4 \DLX_EXinst__n0006<15>6  (
    .ADR0(\DLX_EXinst_Mshift__n0024_Sh[127] ),
    .ADR1(\DLX_EXinst_Mshift__n0027_Sh[47] ),
    .ADR2(DLX_EXinst_N66373),
    .ADR3(DLX_EXinst_N66525),
    .O(\DLX_EXinst_N66525/GROM )
  );
  X_BUF \DLX_EXinst_N66525/XUSED  (
    .I(\DLX_EXinst_N66525/FROM ),
    .O(DLX_EXinst_N66525)
  );
  X_BUF \DLX_EXinst_N66525/YUSED  (
    .I(\DLX_EXinst_N66525/GROM ),
    .O(CHOICE4806)
  );
  defparam DLX_EXinst_Ker664351.INIT = 16'h00CC;
  X_LUT4 DLX_EXinst_Ker664351 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_IR_function_field_0_1),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_IR_function_field_1_1),
    .O(\DLX_EXinst_N66437/FROM )
  );
  defparam DLX_EXinst__n012743_SW0.INIT = 16'h5551;
  X_LUT4 DLX_EXinst__n012743_SW0 (
    .ADR0(DLX_IDinst_IR_function_field[5]),
    .ADR1(DLX_IDinst_IR_function_field[2]),
    .ADR2(DLX_IDinst_IR_function_field[3]),
    .ADR3(DLX_EXinst_N66437),
    .O(\DLX_EXinst_N66437/GROM )
  );
  X_BUF \DLX_EXinst_N66437/XUSED  (
    .I(\DLX_EXinst_N66437/FROM ),
    .O(DLX_EXinst_N66437)
  );
  X_BUF \DLX_EXinst_N66437/YUSED  (
    .I(\DLX_EXinst_N66437/GROM ),
    .O(N126528)
  );
  defparam \DLX_EXinst_Mshift__n0027_Sh<4>25 .INIT = 16'h4450;
  X_LUT4 \DLX_EXinst_Mshift__n0027_Sh<4>25  (
    .ADR0(DLX_IDinst_IR_function_field_1_1),
    .ADR1(DLX_IDinst_reg_out_A[3]),
    .ADR2(DLX_IDinst_reg_out_A[4]),
    .ADR3(DLX_IDinst_IR_function_field_0_1),
    .O(\CHOICE1012/FROM )
  );
  defparam DLX_EXinst_Ker649071.INIT = 16'hD8D8;
  X_LUT4 DLX_EXinst_Ker649071 (
    .ADR0(DLX_IDinst_IR_function_field_1_1),
    .ADR1(DLX_IDinst_reg_out_A[6]),
    .ADR2(DLX_IDinst_reg_out_A[4]),
    .ADR3(VCC),
    .O(\CHOICE1012/GROM )
  );
  X_BUF \CHOICE1012/XUSED  (
    .I(\CHOICE1012/FROM ),
    .O(CHOICE1012)
  );
  X_BUF \CHOICE1012/YUSED  (
    .I(\CHOICE1012/GROM ),
    .O(DLX_EXinst_N64909)
  );
  defparam \DLX_EXinst__n0006<7>16 .INIT = 16'h8008;
  X_LUT4 \DLX_EXinst__n0006<7>16  (
    .ADR0(DLX_EXinst_N66105),
    .ADR1(\DLX_IDinst_Imm[7] ),
    .ADR2(N127392),
    .ADR3(DLX_IDinst_IR_opcode_field[1]),
    .O(\CHOICE3802/FROM )
  );
  defparam \DLX_EXinst__n0006<6>16 .INIT = 16'h8040;
  X_LUT4 \DLX_EXinst__n0006<6>16  (
    .ADR0(DLX_IDinst_IR_opcode_field[1]),
    .ADR1(\DLX_IDinst_Imm[6] ),
    .ADR2(DLX_EXinst_N66105),
    .ADR3(N127286),
    .O(\CHOICE3802/GROM )
  );
  X_BUF \CHOICE3802/XUSED  (
    .I(\CHOICE3802/FROM ),
    .O(CHOICE3802)
  );
  X_BUF \CHOICE3802/YUSED  (
    .I(\CHOICE3802/GROM ),
    .O(CHOICE4354)
  );
  defparam vga_top_vga1__n0012_SW0.INIT = 16'h5F5F;
  X_LUT4 vga_top_vga1__n0012_SW0 (
    .ADR0(vga_top_vga1_N73399),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_N73357),
    .ADR3(VCC),
    .O(\N90461/FROM )
  );
  defparam vga_top_vga1__n0012_1166.INIT = 16'hAAAB;
  X_LUT4 vga_top_vga1__n0012_1166 (
    .ADR0(reset_IBUF_1),
    .ADR1(vga_top_vga1_hcounter[5]),
    .ADR2(vga_top_vga1_hcounter[9]),
    .ADR3(N90461),
    .O(\N90461/GROM )
  );
  X_BUF \N90461/XUSED  (
    .I(\N90461/FROM ),
    .O(N90461)
  );
  X_BUF \N90461/YUSED  (
    .I(\N90461/GROM ),
    .O(vga_top_vga1__n0012)
  );
  defparam DLX_EXinst_Ker637881.INIT = 16'hCFC0;
  X_LUT4 DLX_EXinst_Ker637881 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[27]),
    .ADR2(DLX_IDinst_IR_function_field_1_1),
    .ADR3(DLX_IDinst_reg_out_A[25]),
    .O(\DLX_EXinst_N63790/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0028_Sh<24>1 .INIT = 16'hEE22;
  X_LUT4 \DLX_EXinst_Mshift__n0028_Sh<24>1  (
    .ADR0(DLX_EXinst_N63279),
    .ADR1(DLX_IDinst_IR_function_field_0_1),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N63790),
    .O(\DLX_EXinst_N63790/GROM )
  );
  X_BUF \DLX_EXinst_N63790/XUSED  (
    .I(\DLX_EXinst_N63790/FROM ),
    .O(DLX_EXinst_N63790)
  );
  X_BUF \DLX_EXinst_N63790/YUSED  (
    .I(\DLX_EXinst_N63790/GROM ),
    .O(\DLX_EXinst_Mshift__n0028_Sh[24] )
  );
  defparam DLX_EXinst_Ker663481.INIT = 16'hAA8A;
  X_LUT4 DLX_EXinst_Ker663481 (
    .ADR0(DLX_EXinst__n0149),
    .ADR1(DLX_IDinst_reg_dst),
    .ADR2(DLX_EXinst__n0147),
    .ADR3(DLX_IDinst_IR_opcode_field[0]),
    .O(\DLX_EXinst_reg_out_B_EX<15>/FROM )
  );
  defparam \DLX_EXinst__n0007<15>1 .INIT = 16'hCC00;
  X_LUT4 \DLX_EXinst__n0007<15>1  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_B[15]),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N66350),
    .O(DLX_EXinst__n0007[15])
  );
  X_BUF \DLX_EXinst_reg_out_B_EX<15>/XUSED  (
    .I(\DLX_EXinst_reg_out_B_EX<15>/FROM ),
    .O(DLX_EXinst_N66350)
  );
  defparam \DLX_EXinst_Mshift__n0025_Sh<5>26 .INIT = 16'h5140;
  X_LUT4 \DLX_EXinst_Mshift__n0025_Sh<5>26  (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(DLX_IDinst_reg_out_B[0]),
    .ADR2(DLX_IDinst_reg_out_A[4]),
    .ADR3(DLX_IDinst_reg_out_A[5]),
    .O(\CHOICE1072/FROM )
  );
  defparam DLX_EXinst_Ker629041.INIT = 16'hF3E2;
  X_LUT4 DLX_EXinst_Ker629041 (
    .ADR0(CHOICE1066),
    .ADR1(DLX_IDinst_reg_out_B_2_1),
    .ADR2(\DLX_EXinst_Mshift__n0025_Sh[1] ),
    .ADR3(CHOICE1072),
    .O(\CHOICE1072/GROM )
  );
  X_BUF \CHOICE1072/XUSED  (
    .I(\CHOICE1072/FROM ),
    .O(CHOICE1072)
  );
  X_BUF \CHOICE1072/YUSED  (
    .I(\CHOICE1072/GROM ),
    .O(DLX_EXinst_N62906)
  );
  defparam \mask<0>_SW0 .INIT = 16'hAF03;
  X_LUT4 \mask<0>_SW0  (
    .ADR0(DLX_EXinst_ALU_result[1]),
    .ADR1(DLX_EXinst_word),
    .ADR2(DLX_EXinst_byte),
    .ADR3(DLX_EXinst_ALU_result[0]),
    .O(\N90557/FROM )
  );
  defparam \mask<0> .INIT = 16'hF000;
  X_LUT4 \mask<0>  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(vga_select_6[0]),
    .ADR3(N90557),
    .O(\N90557/GROM )
  );
  X_BUF \N90557/XUSED  (
    .I(\N90557/FROM ),
    .O(N90557)
  );
  X_BUF \N90557/YUSED  (
    .I(\N90557/GROM ),
    .O(mask_0_OBUF)
  );
  defparam DLX_EXinst_Ker629891.INIT = 16'hAACC;
  X_LUT4 DLX_EXinst_Ker629891 (
    .ADR0(DLX_IDinst_reg_out_A[15]),
    .ADR1(DLX_IDinst_reg_out_A[13]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_IR_function_field[1]),
    .O(\DLX_EXinst_N62991/FROM )
  );
  defparam DLX_EXinst_Ker6450311.INIT = 16'hA820;
  X_LUT4 DLX_EXinst_Ker6450311 (
    .ADR0(DLX_IDinst_IR_function_field[3]),
    .ADR1(DLX_IDinst_IR_function_field[0]),
    .ADR2(DLX_EXinst_N63494),
    .ADR3(DLX_EXinst_N62991),
    .O(\DLX_EXinst_N62991/GROM )
  );
  X_BUF \DLX_EXinst_N62991/XUSED  (
    .I(\DLX_EXinst_N62991/FROM ),
    .O(DLX_EXinst_N62991)
  );
  X_BUF \DLX_EXinst_N62991/YUSED  (
    .I(\DLX_EXinst_N62991/GROM ),
    .O(CHOICE1270)
  );
  defparam DLX_EXinst_Ker665331.INIT = 16'h0C0C;
  X_LUT4 DLX_EXinst_Ker665331 (
    .ADR0(VCC),
    .ADR1(DLX_EXinst__n0048),
    .ADR2(DLX_IDinst_reg_out_B[4]),
    .ADR3(VCC),
    .O(\DLX_EXinst_N66535/FROM )
  );
  defparam \DLX_EXinst__n0006<2>298 .INIT = 16'h0008;
  X_LUT4 \DLX_EXinst__n0006<2>298  (
    .ADR0(\DLX_EXinst_Mshift__n0025_Sh[2] ),
    .ADR1(DLX_EXinst_N66535),
    .ADR2(DLX_IDinst_reg_out_B[2]),
    .ADR3(DLX_IDinst_reg_out_B[3]),
    .O(\DLX_EXinst_N66535/GROM )
  );
  X_BUF \DLX_EXinst_N66535/XUSED  (
    .I(\DLX_EXinst_N66535/FROM ),
    .O(DLX_EXinst_N66535)
  );
  X_BUF \DLX_EXinst_N66535/YUSED  (
    .I(\DLX_EXinst_N66535/GROM ),
    .O(CHOICE5556)
  );
  defparam DLX_EXinst_Ker662691.INIT = 16'h0203;
  X_LUT4 DLX_EXinst_Ker662691 (
    .ADR0(DLX_IDinst_reg_dst),
    .ADR1(DLX_IDinst_counter[1]),
    .ADR2(DLX_IDinst_counter[0]),
    .ADR3(DLX_EXinst__n0147),
    .O(\DLX_EXinst_reg_out_B_EX<31>/FROM )
  );
  defparam \DLX_EXinst__n0007<31>1 .INIT = 16'hAA00;
  X_LUT4 \DLX_EXinst__n0007<31>1  (
    .ADR0(DLX_IDinst_reg_out_B[31]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N66271),
    .O(DLX_EXinst__n0007[31])
  );
  X_BUF \DLX_EXinst_reg_out_B_EX<31>/XUSED  (
    .I(\DLX_EXinst_reg_out_B_EX<31>/FROM ),
    .O(DLX_EXinst_N66271)
  );
  defparam \DLX_EXinst__n0006<28>212 .INIT = 16'h4400;
  X_LUT4 \DLX_EXinst__n0006<28>212  (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(DLX_EXinst__n0049),
    .ADR2(VCC),
    .ADR3(\DLX_EXinst_Mshift__n0026_Sh[60] ),
    .O(\CHOICE5223/FROM )
  );
  defparam DLX_EXinst_Ker663811.INIT = 16'hC0C0;
  X_LUT4 DLX_EXinst_Ker663811 (
    .ADR0(VCC),
    .ADR1(DLX_EXinst__n0049),
    .ADR2(DLX_IDinst_reg_out_B[4]),
    .ADR3(VCC),
    .O(\CHOICE5223/GROM )
  );
  X_BUF \CHOICE5223/XUSED  (
    .I(\CHOICE5223/FROM ),
    .O(CHOICE5223)
  );
  X_BUF \CHOICE5223/YUSED  (
    .I(\CHOICE5223/GROM ),
    .O(DLX_EXinst_N66383)
  );
  defparam \DLX_EXinst_Mshift__n0025_Sh<5>28 .INIT = 16'hFCFC;
  X_LUT4 \DLX_EXinst_Mshift__n0025_Sh<5>28  (
    .ADR0(VCC),
    .ADR1(CHOICE1066),
    .ADR2(CHOICE1072),
    .ADR3(VCC),
    .O(\DLX_EXinst_Mshift__n0025_Sh<5>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0025_Sh<5>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0025_Sh<5>/GROM ),
    .O(\DLX_EXinst_Mshift__n0025_Sh[5] )
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_inv_01.INIT = 16'h50F5;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_inv_01 (
    .ADR0(DLX_EXinst_Mcompar__n0061_inst_cy_228),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(DLX_IDinst_reg_out_B[31]),
    .O(\DLX_EXinst__n0061/FROM )
  );
  defparam \DLX_EXinst__n0006<0>235 .INIT = 16'h0E02;
  X_LUT4 \DLX_EXinst__n0006<0>235  (
    .ADR0(DLX_EXinst__n0053),
    .ADR1(DLX_IDinst_IR_function_field[2]),
    .ADR2(DLX_IDinst_IR_function_field[0]),
    .ADR3(DLX_EXinst__n0061),
    .O(\DLX_EXinst__n0061/GROM )
  );
  X_BUF \DLX_EXinst__n0061/XUSED  (
    .I(\DLX_EXinst__n0061/FROM ),
    .O(DLX_EXinst__n0061)
  );
  X_BUF \DLX_EXinst__n0061/YUSED  (
    .I(\DLX_EXinst__n0061/GROM ),
    .O(CHOICE5905)
  );
  defparam \DLX_EXinst__n0006<7>46 .INIT = 16'h0200;
  X_LUT4 \DLX_EXinst__n0006<7>46  (
    .ADR0(DLX_EXinst_N62831),
    .ADR1(DLX_IDinst_IR_function_field[3]),
    .ADR2(N109130),
    .ADR3(DLX_EXinst__n0081),
    .O(\CHOICE3812/FROM )
  );
  defparam \DLX_EXinst__n0006<6>46 .INIT = 16'h0020;
  X_LUT4 \DLX_EXinst__n0006<6>46  (
    .ADR0(DLX_EXinst__n0081),
    .ADR1(N109130),
    .ADR2(DLX_EXinst_N62826),
    .ADR3(DLX_IDinst_IR_function_field[3]),
    .O(\CHOICE3812/GROM )
  );
  X_BUF \CHOICE3812/XUSED  (
    .I(\CHOICE3812/FROM ),
    .O(CHOICE3812)
  );
  X_BUF \CHOICE3812/YUSED  (
    .I(\CHOICE3812/GROM ),
    .O(CHOICE4364)
  );
  defparam \DLX_EXinst__n0006<6>38 .INIT = 16'hD080;
  X_LUT4 \DLX_EXinst__n0006<6>38  (
    .ADR0(DLX_IDinst_IR_function_field[2]),
    .ADR1(DLX_EXinst_N64814),
    .ADR2(DLX_EXinst_N63185),
    .ADR3(N97521),
    .O(\CHOICE4361/FROM )
  );
  defparam \DLX_EXinst__n0006<6>80 .INIT = 16'hF5F4;
  X_LUT4 \DLX_EXinst__n0006<6>80  (
    .ADR0(DLX_IDinst_IR_function_field[4]),
    .ADR1(CHOICE4364),
    .ADR2(CHOICE4370),
    .ADR3(CHOICE4361),
    .O(\CHOICE4361/GROM )
  );
  X_BUF \CHOICE4361/XUSED  (
    .I(\CHOICE4361/FROM ),
    .O(CHOICE4361)
  );
  X_BUF \CHOICE4361/YUSED  (
    .I(\CHOICE4361/GROM ),
    .O(CHOICE4371)
  );
  defparam DLX_EXinst__n01141.INIT = 16'h0100;
  X_LUT4 DLX_EXinst__n01141 (
    .ADR0(DLX_IDinst_IR_function_field[2]),
    .ADR1(DLX_IDinst_IR_function_field[4]),
    .ADR2(DLX_IDinst_IR_function_field[3]),
    .ADR3(DLX_IDinst_IR_function_field[5]),
    .O(\DLX_EXinst__n0114/FROM )
  );
  defparam \DLX_EXinst__n0006<25>240 .INIT = 16'hFEFC;
  X_LUT4 \DLX_EXinst__n0006<25>240  (
    .ADR0(DLX_EXinst__n0016[25]),
    .ADR1(CHOICE4792),
    .ADR2(N126281),
    .ADR3(DLX_EXinst__n0114),
    .O(\DLX_EXinst__n0114/GROM )
  );
  X_BUF \DLX_EXinst__n0114/XUSED  (
    .I(\DLX_EXinst__n0114/FROM ),
    .O(DLX_EXinst__n0114)
  );
  X_BUF \DLX_EXinst__n0114/YUSED  (
    .I(\DLX_EXinst__n0114/GROM ),
    .O(CHOICE4796)
  );
  defparam DLX_EXinst_Ker663901.INIT = 16'h0C0C;
  X_LUT4 DLX_EXinst_Ker663901 (
    .ADR0(VCC),
    .ADR1(DLX_EXinst__n0049),
    .ADR2(DLX_IDinst_reg_out_B[4]),
    .ADR3(VCC),
    .O(\DLX_EXinst_N66392/FROM )
  );
  defparam \DLX_EXinst__n0006<29>216 .INIT = 16'h0400;
  X_LUT4 \DLX_EXinst__n0006<29>216  (
    .ADR0(DLX_IDinst_reg_out_B[3]),
    .ADR1(DLX_EXinst_N66392),
    .ADR2(DLX_IDinst_reg_out_B[2]),
    .ADR3(\DLX_EXinst_Mshift__n0026_Sh[29] ),
    .O(\DLX_EXinst_N66392/GROM )
  );
  X_BUF \DLX_EXinst_N66392/XUSED  (
    .I(\DLX_EXinst_N66392/FROM ),
    .O(DLX_EXinst_N66392)
  );
  X_BUF \DLX_EXinst_N66392/YUSED  (
    .I(\DLX_EXinst_N66392/GROM ),
    .O(CHOICE5377)
  );
  defparam DLX_EXinst_Ker629991.INIT = 16'hEE44;
  X_LUT4 DLX_EXinst_Ker629991 (
    .ADR0(DLX_IDinst_IR_function_field[1]),
    .ADR1(DLX_IDinst_reg_out_A[17]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[19]),
    .O(\DLX_EXinst_N63001/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0028_Sh<16>1 .INIT = 16'hFA0A;
  X_LUT4 \DLX_EXinst_Mshift__n0028_Sh<16>1  (
    .ADR0(DLX_EXinst_N63504),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_IR_function_field_0_1),
    .ADR3(DLX_EXinst_N63001),
    .O(\DLX_EXinst_N63001/GROM )
  );
  X_BUF \DLX_EXinst_N63001/XUSED  (
    .I(\DLX_EXinst_N63001/FROM ),
    .O(DLX_EXinst_N63001)
  );
  X_BUF \DLX_EXinst_N63001/YUSED  (
    .I(\DLX_EXinst_N63001/GROM ),
    .O(\DLX_EXinst_Mshift__n0028_Sh[16] )
  );
  defparam \DLX_EXinst_Mshift__n0025_Sh<6>25 .INIT = 16'h00E2;
  X_LUT4 \DLX_EXinst_Mshift__n0025_Sh<6>25  (
    .ADR0(DLX_IDinst_reg_out_A[6]),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(DLX_IDinst_reg_out_A[4]),
    .ADR3(DLX_IDinst_reg_out_B[0]),
    .O(\CHOICE1300/FROM )
  );
  defparam DLX_EXinst_Ker629091.INIT = 16'hF5E4;
  X_LUT4 DLX_EXinst_Ker629091 (
    .ADR0(DLX_IDinst_reg_out_B_2_1),
    .ADR1(CHOICE1294),
    .ADR2(\DLX_EXinst_Mshift__n0025_Sh[2] ),
    .ADR3(CHOICE1300),
    .O(\CHOICE1300/GROM )
  );
  X_BUF \CHOICE1300/XUSED  (
    .I(\CHOICE1300/FROM ),
    .O(CHOICE1300)
  );
  X_BUF \CHOICE1300/YUSED  (
    .I(\CHOICE1300/GROM ),
    .O(DLX_EXinst_N62911)
  );
  defparam DLX_EXinst_Ker66307133.INIT = 16'h0001;
  X_LUT4 DLX_EXinst_Ker66307133 (
    .ADR0(DLX_IDinst_reg_out_B[6]),
    .ADR1(DLX_IDinst_reg_out_B[7]),
    .ADR2(DLX_IDinst_reg_out_B[8]),
    .ADR3(DLX_IDinst_reg_out_B[9]),
    .O(\CHOICE3610/FROM )
  );
  defparam DLX_EXinst__n00354.INIT = 16'hFFFE;
  X_LUT4 DLX_EXinst__n00354 (
    .ADR0(DLX_IDinst_reg_out_B[7]),
    .ADR1(DLX_IDinst_reg_out_B[6]),
    .ADR2(DLX_IDinst_reg_out_B[5]),
    .ADR3(DLX_IDinst_reg_out_B[31]),
    .O(\CHOICE3610/GROM )
  );
  X_BUF \CHOICE3610/XUSED  (
    .I(\CHOICE3610/FROM ),
    .O(CHOICE3610)
  );
  X_BUF \CHOICE3610/YUSED  (
    .I(\CHOICE3610/GROM ),
    .O(CHOICE3534)
  );
  defparam \DLX_EXinst__n0006<10>21 .INIT = 16'hA2A0;
  X_LUT4 \DLX_EXinst__n0006<10>21  (
    .ADR0(DLX_IDinst_reg_out_A[10]),
    .ADR1(\DLX_IDinst_Imm[10] ),
    .ADR2(DLX_EXinst__n0079),
    .ADR3(DLX_EXinst__n0080),
    .O(\CHOICE4492/FROM )
  );
  defparam \DLX_EXinst__n0006<6>76 .INIT = 16'hD0C0;
  X_LUT4 \DLX_EXinst__n0006<6>76  (
    .ADR0(\DLX_IDinst_Imm[6] ),
    .ADR1(DLX_EXinst__n0079),
    .ADR2(DLX_IDinst_reg_out_A[6]),
    .ADR3(DLX_EXinst__n0080),
    .O(\CHOICE4492/GROM )
  );
  X_BUF \CHOICE4492/XUSED  (
    .I(\CHOICE4492/FROM ),
    .O(CHOICE4492)
  );
  X_BUF \CHOICE4492/YUSED  (
    .I(\CHOICE4492/GROM ),
    .O(CHOICE4370)
  );
  defparam DLX_EXinst_Ker6581510.INIT = 16'h8C88;
  X_LUT4 DLX_EXinst_Ker6581510 (
    .ADR0(DLX_EXinst_N66507),
    .ADR1(\DLX_EXinst_Mshift__n0024_Sh[28] ),
    .ADR2(\DLX_IDinst_Imm[5] ),
    .ADR3(N110065),
    .O(\CHOICE2075/FROM )
  );
  defparam DLX_EXinst_Ker664731.INIT = 16'h00AE;
  X_LUT4 DLX_EXinst_Ker664731 (
    .ADR0(DLX_EXinst_N66507),
    .ADR1(N110065),
    .ADR2(\DLX_IDinst_Imm[5] ),
    .ADR3(DLX_IDinst_IR_function_field[4]),
    .O(\CHOICE2075/GROM )
  );
  X_BUF \CHOICE2075/XUSED  (
    .I(\CHOICE2075/FROM ),
    .O(CHOICE2075)
  );
  X_BUF \CHOICE2075/YUSED  (
    .I(\CHOICE2075/GROM ),
    .O(DLX_EXinst_N66475)
  );
  defparam \DLX_EXinst_Mshift__n0025_Sh<6>28 .INIT = 16'hFAFA;
  X_LUT4 \DLX_EXinst_Mshift__n0025_Sh<6>28  (
    .ADR0(CHOICE1300),
    .ADR1(VCC),
    .ADR2(CHOICE1294),
    .ADR3(VCC),
    .O(\DLX_EXinst_Mshift__n0025_Sh<6>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0025_Sh<6>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0025_Sh<6>/GROM ),
    .O(\DLX_EXinst_Mshift__n0025_Sh[6] )
  );
  defparam \DLX_EXinst__n0006<7>38 .INIT = 16'hE020;
  X_LUT4 \DLX_EXinst__n0006<7>38  (
    .ADR0(N96513),
    .ADR1(DLX_IDinst_IR_function_field[2]),
    .ADR2(DLX_EXinst_N63185),
    .ADR3(DLX_EXinst_N65100),
    .O(\CHOICE3809/FROM )
  );
  defparam \DLX_EXinst__n0006<7>80 .INIT = 16'hBBBA;
  X_LUT4 \DLX_EXinst__n0006<7>80  (
    .ADR0(CHOICE3818),
    .ADR1(DLX_IDinst_IR_function_field[4]),
    .ADR2(CHOICE3812),
    .ADR3(CHOICE3809),
    .O(\CHOICE3809/GROM )
  );
  X_BUF \CHOICE3809/XUSED  (
    .I(\CHOICE3809/FROM ),
    .O(CHOICE3809)
  );
  X_BUF \CHOICE3809/YUSED  (
    .I(\CHOICE3809/GROM ),
    .O(CHOICE3819)
  );
  defparam \DLX_EXinst__n0006<9>215 .INIT = 16'hEAC0;
  X_LUT4 \DLX_EXinst__n0006<9>215  (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(DLX_EXinst_ALU_result[9]),
    .ADR2(N101725),
    .ADR3(N108593),
    .O(\CHOICE4599/FROM )
  );
  defparam \DLX_EXinst__n0006<25>240_SW0 .INIT = 16'hF444;
  X_LUT4 \DLX_EXinst__n0006<25>240_SW0  (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(N108593),
    .ADR2(N101725),
    .ADR3(DLX_EXinst_ALU_result[25]),
    .O(\CHOICE4599/GROM )
  );
  X_BUF \CHOICE4599/XUSED  (
    .I(\CHOICE4599/FROM ),
    .O(CHOICE4599)
  );
  X_BUF \CHOICE4599/YUSED  (
    .I(\CHOICE4599/GROM ),
    .O(N126281)
  );
  defparam DLX_EXinst__n00461.INIT = 16'h2000;
  X_LUT4 DLX_EXinst__n00461 (
    .ADR0(DLX_IDinst_IR_function_field[0]),
    .ADR1(DLX_IDinst_IR_function_field[1]),
    .ADR2(DLX_EXinst_N66096),
    .ADR3(DLX_IDinst_IR_function_field[5]),
    .O(\DLX_EXinst__n0046/FROM )
  );
  defparam \DLX_EXinst__n0006<28>249 .INIT = 16'hF020;
  X_LUT4 \DLX_EXinst__n0006<28>249  (
    .ADR0(DLX_EXinst__n0047),
    .ADR1(DLX_IDinst_reg_out_A[28]),
    .ADR2(DLX_IDinst_reg_out_B[28]),
    .ADR3(DLX_EXinst__n0046),
    .O(\DLX_EXinst__n0046/GROM )
  );
  X_BUF \DLX_EXinst__n0046/XUSED  (
    .I(\DLX_EXinst__n0046/FROM ),
    .O(DLX_EXinst__n0046)
  );
  X_BUF \DLX_EXinst__n0046/YUSED  (
    .I(\DLX_EXinst__n0046/GROM ),
    .O(CHOICE5229)
  );
  defparam \DLX_EXinst__n0006<22>85 .INIT = 16'h9000;
  X_LUT4 \DLX_EXinst__n0006<22>85  (
    .ADR0(N127388),
    .ADR1(DLX_IDinst_IR_opcode_field[1]),
    .ADR2(DLX_EXinst_N66105),
    .ADR3(\DLX_IDinst_Imm[31] ),
    .O(\CHOICE4119/FROM )
  );
  defparam \DLX_EXinst__n0006<8>16 .INIT = 16'h9000;
  X_LUT4 \DLX_EXinst__n0006<8>16  (
    .ADR0(DLX_IDinst_IR_opcode_field[1]),
    .ADR1(N127302),
    .ADR2(\DLX_IDinst_Imm[8] ),
    .ADR3(DLX_EXinst_N66105),
    .O(\CHOICE4119/GROM )
  );
  X_BUF \CHOICE4119/XUSED  (
    .I(\CHOICE4119/FROM ),
    .O(CHOICE4119)
  );
  X_BUF \CHOICE4119/YUSED  (
    .I(\CHOICE4119/GROM ),
    .O(CHOICE3684)
  );
  defparam DLX_EXinst_Ker64446_SW0.INIT = 16'hF7F7;
  X_LUT4 DLX_EXinst_Ker64446_SW0 (
    .ADR0(DLX_IDinst_IR_function_field[0]),
    .ADR1(DLX_IDinst_IR_function_field[5]),
    .ADR2(DLX_IDinst_IR_function_field_1_1),
    .ADR3(VCC),
    .O(\N127412/FROM )
  );
  defparam DLX_EXinst__n00471.INIT = 16'h0800;
  X_LUT4 DLX_EXinst__n00471 (
    .ADR0(DLX_IDinst_IR_function_field[5]),
    .ADR1(DLX_IDinst_IR_function_field[1]),
    .ADR2(DLX_IDinst_IR_function_field[0]),
    .ADR3(DLX_EXinst_N66096),
    .O(\N127412/GROM )
  );
  X_BUF \N127412/XUSED  (
    .I(\N127412/FROM ),
    .O(N127412)
  );
  X_BUF \N127412/YUSED  (
    .I(\N127412/GROM ),
    .O(DLX_EXinst__n0047)
  );
  defparam DLX_EXinst__n00481.INIT = 16'h0100;
  X_LUT4 DLX_EXinst__n00481 (
    .ADR0(DLX_IDinst_IR_function_field[0]),
    .ADR1(DLX_IDinst_IR_function_field[5]),
    .ADR2(DLX_IDinst_IR_function_field[1]),
    .ADR3(DLX_EXinst_N66096),
    .O(\DLX_EXinst__n0048/FROM )
  );
  defparam DLX_EXinst_Ker662241.INIT = 16'h0100;
  X_LUT4 DLX_EXinst_Ker662241 (
    .ADR0(CHOICE3540),
    .ADR1(CHOICE3534),
    .ADR2(CHOICE3556),
    .ADR3(DLX_EXinst__n0048),
    .O(\DLX_EXinst__n0048/GROM )
  );
  X_BUF \DLX_EXinst__n0048/XUSED  (
    .I(\DLX_EXinst__n0048/FROM ),
    .O(DLX_EXinst__n0048)
  );
  X_BUF \DLX_EXinst__n0048/YUSED  (
    .I(\DLX_EXinst__n0048/GROM ),
    .O(DLX_EXinst_N66226)
  );
  defparam DLX_IDinst_Ker70293_SW0.INIT = 16'hAAFF;
  X_LUT4 DLX_IDinst_Ker70293_SW0 (
    .ADR0(DLX_IDinst__n03641_1),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst__n0250),
    .O(\N90344/FROM )
  );
  defparam DLX_IDinst_Ker70293.INIT = 16'hA0EC;
  X_LUT4 DLX_IDinst_Ker70293 (
    .ADR0(DLX_IDinst_N70918),
    .ADR1(DLX_IDinst_N70885),
    .ADR2(DLX_IDinst_IR_latched[30]),
    .ADR3(N90344),
    .O(\N90344/GROM )
  );
  X_BUF \N90344/XUSED  (
    .I(\N90344/FROM ),
    .O(N90344)
  );
  X_BUF \N90344/YUSED  (
    .I(\N90344/GROM ),
    .O(DLX_IDinst_N70295)
  );
  defparam DLX_EXinst__n00491.INIT = 16'h1000;
  X_LUT4 DLX_EXinst__n00491 (
    .ADR0(DLX_IDinst_IR_function_field[0]),
    .ADR1(DLX_IDinst_IR_function_field[5]),
    .ADR2(DLX_IDinst_IR_function_field[1]),
    .ADR3(DLX_EXinst_N66096),
    .O(\DLX_EXinst__n0049/FROM )
  );
  defparam DLX_EXinst_Ker664921.INIT = 16'h0100;
  X_LUT4 DLX_EXinst_Ker664921 (
    .ADR0(CHOICE3540),
    .ADR1(CHOICE3534),
    .ADR2(CHOICE3556),
    .ADR3(DLX_EXinst__n0049),
    .O(\DLX_EXinst__n0049/GROM )
  );
  X_BUF \DLX_EXinst__n0049/XUSED  (
    .I(\DLX_EXinst__n0049/FROM ),
    .O(DLX_EXinst__n0049)
  );
  X_BUF \DLX_EXinst__n0049/YUSED  (
    .I(\DLX_EXinst__n0049/GROM ),
    .O(DLX_EXinst_N66494)
  );
  defparam DLX_EXinst__n00811.INIT = 16'h0022;
  X_LUT4 DLX_EXinst__n00811 (
    .ADR0(DLX_EXinst_N66112),
    .ADR1(DLX_IDinst_IR_opcode_field[1]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_IR_opcode_field[0]),
    .O(\DLX_EXinst__n0081/FROM )
  );
  defparam DLX_EXinst_Ker66517_SW1.INIT = 16'hFAFF;
  X_LUT4 DLX_EXinst_Ker66517_SW1 (
    .ADR0(DLX_IDinst_IR_function_field_2_1),
    .ADR1(VCC),
    .ADR2(N109130),
    .ADR3(DLX_EXinst__n0081),
    .O(\DLX_EXinst__n0081/GROM )
  );
  X_BUF \DLX_EXinst__n0081/XUSED  (
    .I(\DLX_EXinst__n0081/FROM ),
    .O(DLX_EXinst__n0081)
  );
  X_BUF \DLX_EXinst__n0081/YUSED  (
    .I(\DLX_EXinst__n0081/GROM ),
    .O(N127093)
  );
  defparam vga_top_vga1_helpme_1167.INIT = 1'b1;
  X_SFF vga_top_vga1_helpme_1167 (
    .I(\vga_top_vga1_helpme/LOGIC_ZERO ),
    .CE(vga_top_vga1__n0052),
    .CLK(clkdiv_vga),
    .SET(GSR),
    .RST(GND),
    .SSET(reset_IBUF_1),
    .SRST(GND),
    .O(vga_top_vga1_helpme)
  );
  X_ZERO \vga_top_vga1_helpme/LOGIC_ZERO_1168  (
    .O(\vga_top_vga1_helpme/LOGIC_ZERO )
  );
  defparam \DLX_EXinst__n0006<8>38 .INIT = 16'hC480;
  X_LUT4 \DLX_EXinst__n0006<8>38  (
    .ADR0(DLX_IDinst_IR_function_field[2]),
    .ADR1(DLX_EXinst_N63185),
    .ADR2(N97233),
    .ADR3(DLX_EXinst_N65105),
    .O(\CHOICE3691/FROM )
  );
  defparam \DLX_EXinst__n0006<8>71 .INIT = 16'hF5F4;
  X_LUT4 \DLX_EXinst__n0006<8>71  (
    .ADR0(DLX_IDinst_IR_function_field[4]),
    .ADR1(CHOICE3692),
    .ADR2(CHOICE3698),
    .ADR3(CHOICE3691),
    .O(\CHOICE3691/GROM )
  );
  X_BUF \CHOICE3691/XUSED  (
    .I(\CHOICE3691/FROM ),
    .O(CHOICE3691)
  );
  X_BUF \CHOICE3691/YUSED  (
    .I(\CHOICE3691/GROM ),
    .O(CHOICE3699)
  );
  X_OR2 \DLX_IFinst_PC<13>/FFY/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_PC<13>/FFY/RST )
  );
  defparam DLX_IFinst_PC_12.INIT = 1'b0;
  X_FF DLX_IFinst_PC_12 (
    .I(DLX_IFinst_NPC[12]),
    .CE(DLX_IFinst_PC_N3535),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_PC<13>/FFY/RST ),
    .O(DLX_IFinst_PC[12])
  );
  defparam DLX_IFinst_IR_previous_28.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_28 (
    .I(DLX_IFinst_IR_latched[28]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[28])
  );
  X_OR2 \DLX_IFinst_PC<23>/FFY/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_PC<23>/FFY/RST )
  );
  defparam DLX_IFinst_PC_22.INIT = 1'b0;
  X_FF DLX_IFinst_PC_22 (
    .I(DLX_IFinst_NPC[22]),
    .CE(DLX_IFinst_PC_N3535),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_PC<23>/FFY/RST ),
    .O(DLX_IFinst_PC[22])
  );
  X_OR2 \DLX_IFinst_PC<15>/FFY/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_PC<15>/FFY/RST )
  );
  defparam DLX_IFinst_PC_14.INIT = 1'b0;
  X_FF DLX_IFinst_PC_14 (
    .I(DLX_IFinst_NPC[14]),
    .CE(DLX_IFinst_PC_N3535),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_PC<15>/FFY/RST ),
    .O(DLX_IFinst_PC[14])
  );
  defparam \DLX_IDinst__n0086<0>6 .INIT = 16'hECA0;
  X_LUT4 \DLX_IDinst__n0086<0>6  (
    .ADR0(DLX_IDinst_EPC[0]),
    .ADR1(DLX_IDinst_N70786),
    .ADR2(DLX_IDinst__n0071),
    .ADR3(DLX_IDinst_branch_address[0]),
    .O(\CHOICE2558/FROM )
  );
  defparam \DLX_IDinst__n0086<11>6 .INIT = 16'hECA0;
  X_LUT4 \DLX_IDinst__n0086<11>6  (
    .ADR0(DLX_IDinst__n0071),
    .ADR1(DLX_IDinst_N70786),
    .ADR2(DLX_IDinst_EPC[11]),
    .ADR3(DLX_IDinst_branch_address[11]),
    .O(\CHOICE2558/GROM )
  );
  X_BUF \CHOICE2558/XUSED  (
    .I(\CHOICE2558/FROM ),
    .O(CHOICE2558)
  );
  X_BUF \CHOICE2558/YUSED  (
    .I(\CHOICE2558/GROM ),
    .O(CHOICE2679)
  );
  defparam DLX_EXinst_Ker66307120.INIT = 16'h0001;
  X_LUT4 DLX_EXinst_Ker66307120 (
    .ADR0(DLX_IDinst_reg_out_B[10]),
    .ADR1(DLX_IDinst_reg_out_B[11]),
    .ADR2(DLX_IDinst_reg_out_B[13]),
    .ADR3(DLX_IDinst_reg_out_B[12]),
    .O(\CHOICE3603/FROM )
  );
  defparam \DLX_EXinst__n0017<11>1 .INIT = 16'hAAF0;
  X_LUT4 \DLX_EXinst__n0017<11>1  (
    .ADR0(DLX_IDinst_reg_out_B[11]),
    .ADR1(VCC),
    .ADR2(\DLX_IDinst_Imm[11] ),
    .ADR3(DLX_EXinst__n0030_1),
    .O(\CHOICE3603/GROM )
  );
  X_BUF \CHOICE3603/XUSED  (
    .I(\CHOICE3603/FROM ),
    .O(CHOICE3603)
  );
  X_BUF \CHOICE3603/YUSED  (
    .I(\CHOICE3603/GROM ),
    .O(DLX_EXinst__n0017[11])
  );
  defparam \DLX_EXinst__n0006<9>42 .INIT = 16'hCA00;
  X_LUT4 \DLX_EXinst__n0006<9>42  (
    .ADR0(DLX_EXinst_N64824),
    .ADR1(DLX_EXinst_N64560),
    .ADR2(DLX_IDinst_IR_function_field[2]),
    .ADR3(DLX_EXinst_N66475),
    .O(\CHOICE4560/FROM )
  );
  defparam \DLX_EXinst__n0006<9>71 .INIT = 16'hFEFE;
  X_LUT4 \DLX_EXinst__n0006<9>71  (
    .ADR0(CHOICE4567),
    .ADR1(CHOICE4566),
    .ADR2(CHOICE4560),
    .ADR3(VCC),
    .O(\CHOICE4560/GROM )
  );
  X_BUF \CHOICE4560/XUSED  (
    .I(\CHOICE4560/FROM ),
    .O(CHOICE4560)
  );
  X_BUF \CHOICE4560/YUSED  (
    .I(\CHOICE4560/GROM ),
    .O(CHOICE4569)
  );
  X_OR2 \DLX_IFinst_PC<17>/FFY/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_PC<17>/FFY/RST )
  );
  defparam DLX_IFinst_PC_16.INIT = 1'b0;
  X_FF DLX_IFinst_PC_16 (
    .I(DLX_IFinst_NPC[16]),
    .CE(DLX_IFinst_PC_N3535),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_PC<17>/FFY/RST ),
    .O(DLX_IFinst_PC[16])
  );
  defparam \DLX_EXinst__n0006<12>67 .INIT = 16'hAE00;
  X_LUT4 \DLX_EXinst__n0006<12>67  (
    .ADR0(DLX_EXinst__n0079),
    .ADR1(DLX_EXinst__n0080),
    .ADR2(\DLX_IDinst_Imm[12] ),
    .ADR3(DLX_IDinst_reg_out_A[12]),
    .O(\CHOICE3876/FROM )
  );
  defparam \DLX_EXinst__n0006<8>67 .INIT = 16'h88A8;
  X_LUT4 \DLX_EXinst__n0006<8>67  (
    .ADR0(DLX_IDinst_reg_out_A[8]),
    .ADR1(DLX_EXinst__n0079),
    .ADR2(DLX_EXinst__n0080),
    .ADR3(\DLX_IDinst_Imm[8] ),
    .O(\CHOICE3876/GROM )
  );
  X_BUF \CHOICE3876/XUSED  (
    .I(\CHOICE3876/FROM ),
    .O(CHOICE3876)
  );
  X_BUF \CHOICE3876/YUSED  (
    .I(\CHOICE3876/GROM ),
    .O(CHOICE3698)
  );
  defparam DLX_EXinst__n01491.INIT = 16'h0505;
  X_LUT4 DLX_EXinst__n01491 (
    .ADR0(DLX_IDinst_counter[0]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_counter[1]),
    .ADR3(VCC),
    .O(\DLX_IDinst_slot_num_FFd2/FROM )
  );
  defparam \DLX_IDinst_slot_num_FFd2-In66 .INIT = 16'h0E00;
  X_LUT4 \DLX_IDinst_slot_num_FFd2-In66  (
    .ADR0(CHOICE2523),
    .ADR1(CHOICE2525),
    .ADR2(DLX_IDinst_intr_slot),
    .ADR3(DLX_EXinst__n0149),
    .O(\DLX_IDinst_slot_num_FFd2-In )
  );
  X_BUF \DLX_IDinst_slot_num_FFd2/XUSED  (
    .I(\DLX_IDinst_slot_num_FFd2/FROM ),
    .O(DLX_EXinst__n0149)
  );
  defparam DLX_EXinst__n00771.INIT = 16'h8080;
  X_LUT4 DLX_EXinst__n00771 (
    .ADR0(DLX_EXinst_N66105),
    .ADR1(DLX_IDinst_IR_opcode_field[1]),
    .ADR2(DLX_IDinst_IR_opcode_field[0]),
    .ADR3(VCC),
    .O(\DLX_EXinst__n0077/FROM )
  );
  defparam \DLX_EXinst__n0006<16>142 .INIT = 16'hFEFC;
  X_LUT4 \DLX_EXinst__n0006<16>142  (
    .ADR0(DLX_IDinst_IR_function_field[0]),
    .ADR1(CHOICE5107),
    .ADR2(CHOICE5128),
    .ADR3(DLX_EXinst__n0077),
    .O(\DLX_EXinst__n0077/GROM )
  );
  X_BUF \DLX_EXinst__n0077/XUSED  (
    .I(\DLX_EXinst__n0077/FROM ),
    .O(DLX_EXinst__n0077)
  );
  X_BUF \DLX_EXinst__n0077/YUSED  (
    .I(\DLX_EXinst__n0077/GROM ),
    .O(CHOICE5129)
  );
  X_OR2 \DLX_IFinst_PC<19>/FFY/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_PC<19>/FFY/RST )
  );
  defparam DLX_IFinst_PC_18.INIT = 1'b0;
  X_FF DLX_IFinst_PC_18 (
    .I(DLX_IFinst_NPC[18]),
    .CE(DLX_IFinst_PC_N3535),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_PC<19>/FFY/RST ),
    .O(DLX_IFinst_PC[18])
  );
  defparam \DLX_IDinst__n0086<6>6 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst__n0086<6>6  (
    .ADR0(DLX_IDinst_N70786),
    .ADR1(DLX_IDinst_branch_address[6]),
    .ADR2(DLX_IDinst_EPC[6]),
    .ADR3(DLX_IDinst__n0071),
    .O(\CHOICE2635/FROM )
  );
  defparam \DLX_IDinst__n0086<12>6 .INIT = 16'hECA0;
  X_LUT4 \DLX_IDinst__n0086<12>6  (
    .ADR0(DLX_IDinst_EPC[12]),
    .ADR1(DLX_IDinst_branch_address[12]),
    .ADR2(DLX_IDinst__n0071),
    .ADR3(DLX_IDinst_N70786),
    .O(\CHOICE2635/GROM )
  );
  X_BUF \CHOICE2635/XUSED  (
    .I(\CHOICE2635/FROM ),
    .O(CHOICE2635)
  );
  X_BUF \CHOICE2635/YUSED  (
    .I(\CHOICE2635/GROM ),
    .O(CHOICE2690)
  );
  defparam \DLX_IDinst__n0086<27>6 .INIT = 16'hEAC0;
  X_LUT4 \DLX_IDinst__n0086<27>6  (
    .ADR0(DLX_IDinst_N70786),
    .ADR1(DLX_IDinst__n0071),
    .ADR2(DLX_IDinst_EPC[27]),
    .ADR3(DLX_IDinst_branch_address[27]),
    .O(\CHOICE2877/FROM )
  );
  defparam \DLX_IDinst__n0086<20>6 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst__n0086<20>6  (
    .ADR0(DLX_IDinst_N70786),
    .ADR1(DLX_IDinst_branch_address[20]),
    .ADR2(DLX_IDinst__n0071),
    .ADR3(DLX_IDinst_EPC[20]),
    .O(\CHOICE2877/GROM )
  );
  X_BUF \CHOICE2877/XUSED  (
    .I(\CHOICE2877/FROM ),
    .O(CHOICE2877)
  );
  X_BUF \CHOICE2877/YUSED  (
    .I(\CHOICE2877/GROM ),
    .O(CHOICE2778)
  );
  defparam \DLX_EXinst__n0017<24>1 .INIT = 16'hECA0;
  X_LUT4 \DLX_EXinst__n0017<24>1  (
    .ADR0(DLX_EXinst__n0030_1),
    .ADR1(\DLX_IDinst_Imm[31] ),
    .ADR2(DLX_IDinst_reg_out_B[24]),
    .ADR3(N100440),
    .O(\DLX_EXinst__n0017<24>/FROM )
  );
  defparam \DLX_EXinst__n0017<20>1 .INIT = 16'hEAC0;
  X_LUT4 \DLX_EXinst__n0017<20>1  (
    .ADR0(\DLX_IDinst_Imm[31] ),
    .ADR1(DLX_EXinst__n0030_1),
    .ADR2(DLX_IDinst_reg_out_B[20]),
    .ADR3(N100440),
    .O(\DLX_EXinst__n0017<24>/GROM )
  );
  X_BUF \DLX_EXinst__n0017<24>/XUSED  (
    .I(\DLX_EXinst__n0017<24>/FROM ),
    .O(DLX_EXinst__n0017[24])
  );
  X_BUF \DLX_EXinst__n0017<24>/YUSED  (
    .I(\DLX_EXinst__n0017<24>/GROM ),
    .O(DLX_EXinst__n0017[20])
  );
  defparam DLX_IDinst__n0331_1169.INIT = 16'hFFFB;
  X_LUT4 DLX_IDinst__n0331_1169 (
    .ADR0(DLX_IDinst_counter[0]),
    .ADR1(N95693),
    .ADR2(DLX_IDinst_counter[1]),
    .ADR3(DLX_IDinst_intr_slot),
    .O(\DLX_IDinst__n0331/FROM )
  );
  defparam DLX_IDinst_Ker706771.INIT = 16'h007F;
  X_LUT4 DLX_IDinst_Ker706771 (
    .ADR0(DLX_IDinst_IR_latched[26]),
    .ADR1(DLX_IDinst_IR_latched[27]),
    .ADR2(DLX_IDinst_N70623),
    .ADR3(DLX_IDinst__n0331),
    .O(\DLX_IDinst__n0331/GROM )
  );
  X_BUF \DLX_IDinst__n0331/XUSED  (
    .I(\DLX_IDinst__n0331/FROM ),
    .O(DLX_IDinst__n0331)
  );
  X_BUF \DLX_IDinst__n0331/YUSED  (
    .I(\DLX_IDinst__n0331/GROM ),
    .O(DLX_IDinst_N70679)
  );
  defparam DLX_EXinst__n00781.INIT = 16'h0022;
  X_LUT4 DLX_EXinst__n00781 (
    .ADR0(DLX_EXinst_N66105),
    .ADR1(DLX_IDinst_IR_opcode_field[1]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_IR_opcode_field[0]),
    .O(\DLX_EXinst__n0078/FROM )
  );
  defparam \DLX_EXinst__n0006<4>57 .INIT = 16'hFEDC;
  X_LUT4 \DLX_EXinst__n0006<4>57  (
    .ADR0(DLX_IDinst_reg_out_A[4]),
    .ADR1(N126038),
    .ADR2(DLX_EXinst__n0080),
    .ADR3(DLX_EXinst__n0078),
    .O(\DLX_EXinst__n0078/GROM )
  );
  X_BUF \DLX_EXinst__n0078/XUSED  (
    .I(\DLX_EXinst__n0078/FROM ),
    .O(DLX_EXinst__n0078)
  );
  X_BUF \DLX_EXinst__n0078/YUSED  (
    .I(\DLX_EXinst__n0078/GROM ),
    .O(CHOICE3990)
  );
  defparam DLX_IDinst__n0443_1170.INIT = 16'h0075;
  X_LUT4 DLX_IDinst__n0443_1170 (
    .ADR0(DLX_IDinst__n0331),
    .ADR1(N90101),
    .ADR2(DLX_IDinst_intr_slot),
    .ADR3(DLX_IDinst__n0335),
    .O(\DLX_IDinst__n0443/FROM )
  );
  defparam DLX_IDinst__n0420_1171.INIT = 16'h00D5;
  X_LUT4 DLX_IDinst__n0420_1171 (
    .ADR0(DLX_IDinst__n0331),
    .ADR1(N90148),
    .ADR2(DLX_IDinst_slot_num_FFd1),
    .ADR3(DLX_IDinst__n0335),
    .O(\DLX_IDinst__n0443/GROM )
  );
  X_BUF \DLX_IDinst__n0443/XUSED  (
    .I(\DLX_IDinst__n0443/FROM ),
    .O(DLX_IDinst__n0443)
  );
  X_BUF \DLX_IDinst__n0443/YUSED  (
    .I(\DLX_IDinst__n0443/GROM ),
    .O(DLX_IDinst__n0420)
  );
  defparam \mask<2>_SW117 .INIT = 16'h07A7;
  X_LUT4 \mask<2>_SW117  (
    .ADR0(DLX_EXinst_ALU_result[0]),
    .ADR1(DLX_EXinst_word),
    .ADR2(DLX_EXinst_byte),
    .ADR3(DLX_EXinst_ALU_result[1]),
    .O(\CHOICE283/FROM )
  );
  defparam \mask<2>_SW122 .INIT = 16'hCC00;
  X_LUT4 \mask<2>_SW122  (
    .ADR0(VCC),
    .ADR1(vga_select_6[0]),
    .ADR2(VCC),
    .ADR3(CHOICE283),
    .O(\CHOICE283/GROM )
  );
  X_BUF \CHOICE283/XUSED  (
    .I(\CHOICE283/FROM ),
    .O(CHOICE283)
  );
  X_BUF \CHOICE283/YUSED  (
    .I(\CHOICE283/GROM ),
    .O(mask_2_OBUF)
  );
  defparam DLX_IDinst__n0440_1172.INIT = 16'h0075;
  X_LUT4 DLX_IDinst__n0440_1172 (
    .ADR0(DLX_EXinst__n0149),
    .ADR1(DLX_IDinst_intr_slot),
    .ADR2(N95693),
    .ADR3(DLX_IDinst__n0335),
    .O(\DLX_IDinst__n0440/FROM )
  );
  defparam DLX_IDinst__n0085_1173.INIT = 16'h0200;
  X_LUT4 DLX_IDinst__n0085_1173 (
    .ADR0(DLX_EXinst__n0149),
    .ADR1(DLX_IDinst_intr_slot),
    .ADR2(N127098),
    .ADR3(N95693),
    .O(\DLX_IDinst__n0440/GROM )
  );
  X_BUF \DLX_IDinst__n0440/XUSED  (
    .I(\DLX_IDinst__n0440/FROM ),
    .O(DLX_IDinst__n0440)
  );
  X_BUF \DLX_IDinst__n0440/YUSED  (
    .I(\DLX_IDinst__n0440/GROM ),
    .O(DLX_IDinst__n0085)
  );
  defparam DLX_EXinst__n00791.INIT = 16'h0A00;
  X_LUT4 DLX_EXinst__n00791 (
    .ADR0(DLX_EXinst_N66105),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_IR_opcode_field[1]),
    .ADR3(DLX_IDinst_IR_opcode_field[0]),
    .O(\DLX_EXinst__n0079/FROM )
  );
  defparam \DLX_EXinst__n0006<28>12 .INIT = 16'hAA08;
  X_LUT4 \DLX_EXinst__n0006<28>12  (
    .ADR0(DLX_IDinst_reg_out_A[28]),
    .ADR1(DLX_EXinst__n0080),
    .ADR2(\DLX_IDinst_Imm[31] ),
    .ADR3(DLX_EXinst__n0079),
    .O(\DLX_EXinst__n0079/GROM )
  );
  X_BUF \DLX_EXinst__n0079/XUSED  (
    .I(\DLX_EXinst__n0079/FROM ),
    .O(DLX_EXinst__n0079)
  );
  X_BUF \DLX_EXinst__n0079/YUSED  (
    .I(\DLX_EXinst__n0079/GROM ),
    .O(CHOICE5181)
  );
  defparam \DLX_IDinst__n0086<14>6 .INIT = 16'hECA0;
  X_LUT4 \DLX_IDinst__n0086<14>6  (
    .ADR0(DLX_IDinst_N70786),
    .ADR1(DLX_IDinst__n0071),
    .ADR2(DLX_IDinst_branch_address[14]),
    .ADR3(DLX_IDinst_EPC[14]),
    .O(\CHOICE2712/FROM )
  );
  defparam \DLX_IDinst__n0086<21>6 .INIT = 16'hEAC0;
  X_LUT4 \DLX_IDinst__n0086<21>6  (
    .ADR0(DLX_IDinst_branch_address[21]),
    .ADR1(DLX_IDinst_EPC[21]),
    .ADR2(DLX_IDinst__n0071),
    .ADR3(DLX_IDinst_N70786),
    .O(\CHOICE2712/GROM )
  );
  X_BUF \CHOICE2712/XUSED  (
    .I(\CHOICE2712/FROM ),
    .O(CHOICE2712)
  );
  X_BUF \CHOICE2712/YUSED  (
    .I(\CHOICE2712/GROM ),
    .O(CHOICE2800)
  );
  defparam \DLX_IDinst__n0086<19>6 .INIT = 16'hECA0;
  X_LUT4 \DLX_IDinst__n0086<19>6  (
    .ADR0(DLX_IDinst_branch_address[19]),
    .ADR1(DLX_IDinst__n0071),
    .ADR2(DLX_IDinst_N70786),
    .ADR3(DLX_IDinst_EPC[19]),
    .O(\CHOICE2756/FROM )
  );
  defparam \DLX_IDinst__n0086<13>6 .INIT = 16'hEAC0;
  X_LUT4 \DLX_IDinst__n0086<13>6  (
    .ADR0(DLX_IDinst_branch_address[13]),
    .ADR1(DLX_IDinst__n0071),
    .ADR2(DLX_IDinst_EPC[13]),
    .ADR3(DLX_IDinst_N70786),
    .O(\CHOICE2756/GROM )
  );
  X_BUF \CHOICE2756/XUSED  (
    .I(\CHOICE2756/FROM ),
    .O(CHOICE2756)
  );
  X_BUF \CHOICE2756/YUSED  (
    .I(\CHOICE2756/GROM ),
    .O(CHOICE2701)
  );
  defparam \DLX_EXinst__n0017<22>1 .INIT = 16'hF888;
  X_LUT4 \DLX_EXinst__n0017<22>1  (
    .ADR0(\DLX_IDinst_Imm[31] ),
    .ADR1(N100440),
    .ADR2(DLX_IDinst_reg_out_B[22]),
    .ADR3(DLX_EXinst__n0030_1),
    .O(\DLX_EXinst__n0017<22>/FROM )
  );
  defparam \DLX_EXinst__n0017<21>1 .INIT = 16'hEAC0;
  X_LUT4 \DLX_EXinst__n0017<21>1  (
    .ADR0(DLX_IDinst_reg_out_B[21]),
    .ADR1(\DLX_IDinst_Imm[31] ),
    .ADR2(N100440),
    .ADR3(DLX_EXinst__n0030_1),
    .O(\DLX_EXinst__n0017<22>/GROM )
  );
  X_BUF \DLX_EXinst__n0017<22>/XUSED  (
    .I(\DLX_EXinst__n0017<22>/FROM ),
    .O(DLX_EXinst__n0017[22])
  );
  X_BUF \DLX_EXinst__n0017<22>/YUSED  (
    .I(\DLX_EXinst__n0017<22>/GROM ),
    .O(DLX_EXinst__n0017[21])
  );
  defparam vga_top_vga1__n0006_SW0.INIT = 16'hFFF3;
  X_LUT4 vga_top_vga1__n0006_SW0 (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_N73389),
    .ADR2(vga_top_vga1_hcounter[0]),
    .ADR3(vga_top_vga1_hcounter[3]),
    .O(\N95654/FROM )
  );
  defparam vga_top_vga1__n0006_1174.INIT = 16'hAAEA;
  X_LUT4 vga_top_vga1__n0006_1174 (
    .ADR0(vga_top_vga1_helpme),
    .ADR1(vga_top_vga1_hcounter[9]),
    .ADR2(vga_top_vga1_hcounter[8]),
    .ADR3(N95654),
    .O(\N95654/GROM )
  );
  X_BUF \N95654/XUSED  (
    .I(\N95654/FROM ),
    .O(N95654)
  );
  X_BUF \N95654/YUSED  (
    .I(\N95654/GROM ),
    .O(vga_top_vga1__n0006)
  );
  defparam vga_top_vga1__n0014_SW0.INIT = 16'hFF5F;
  X_LUT4 vga_top_vga1__n0014_SW0 (
    .ADR0(vga_top_vga1_N73384),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_N73394),
    .ADR3(vga_top_vga1_vcounter[9]),
    .O(\N95611/FROM )
  );
  defparam vga_top_vga1__n0014_1175.INIT = 16'hF0FB;
  X_LUT4 vga_top_vga1__n0014_1175 (
    .ADR0(vga_top_vga1_N73374),
    .ADR1(vga_top_vga1_vcounter[5]),
    .ADR2(reset_IBUF_1),
    .ADR3(N95611),
    .O(\N95611/GROM )
  );
  X_BUF \N95611/XUSED  (
    .I(\N95611/FROM ),
    .O(N95611)
  );
  X_BUF \N95611/YUSED  (
    .I(\N95611/GROM ),
    .O(vga_top_vga1__n0014)
  );
  defparam \DLX_EXinst__n0006<19>42 .INIT = 16'h8200;
  X_LUT4 \DLX_EXinst__n0006<19>42  (
    .ADR0(\DLX_IDinst_Imm[31] ),
    .ADR1(N127404),
    .ADR2(DLX_IDinst_IR_opcode_field[1]),
    .ADR3(DLX_EXinst_N66105),
    .O(\CHOICE4954/FROM )
  );
  defparam \DLX_EXinst__n0006<9>59 .INIT = 16'h8200;
  X_LUT4 \DLX_EXinst__n0006<9>59  (
    .ADR0(\DLX_IDinst_Imm[9] ),
    .ADR1(DLX_IDinst_IR_opcode_field[1]),
    .ADR2(N127378),
    .ADR3(DLX_EXinst_N66105),
    .O(\CHOICE4954/GROM )
  );
  X_BUF \CHOICE4954/XUSED  (
    .I(\CHOICE4954/FROM ),
    .O(CHOICE4954)
  );
  X_BUF \CHOICE4954/YUSED  (
    .I(\CHOICE4954/GROM ),
    .O(CHOICE4566)
  );
  defparam \DLX_IDinst__n0086<23>6 .INIT = 16'hEAC0;
  X_LUT4 \DLX_IDinst__n0086<23>6  (
    .ADR0(DLX_IDinst_N70786),
    .ADR1(DLX_IDinst_EPC[23]),
    .ADR2(DLX_IDinst__n0071),
    .ADR3(DLX_IDinst_branch_address[23]),
    .O(\CHOICE2811/FROM )
  );
  defparam \DLX_IDinst__n0086<22>6 .INIT = 16'hEAC0;
  X_LUT4 \DLX_IDinst__n0086<22>6  (
    .ADR0(DLX_IDinst__n0071),
    .ADR1(DLX_IDinst_N70786),
    .ADR2(DLX_IDinst_branch_address[22]),
    .ADR3(DLX_IDinst_EPC[22]),
    .O(\CHOICE2811/GROM )
  );
  X_BUF \CHOICE2811/XUSED  (
    .I(\CHOICE2811/FROM ),
    .O(CHOICE2811)
  );
  X_BUF \CHOICE2811/YUSED  (
    .I(\CHOICE2811/GROM ),
    .O(CHOICE2822)
  );
  defparam \DLX_IDinst__n0086<9>6 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst__n0086<9>6  (
    .ADR0(DLX_IDinst_N70786),
    .ADR1(DLX_IDinst_branch_address[9]),
    .ADR2(DLX_IDinst__n0071),
    .ADR3(DLX_IDinst_EPC[9]),
    .O(\CHOICE2657/FROM )
  );
  defparam \DLX_IDinst__n0086<30>6 .INIT = 16'hEAC0;
  X_LUT4 \DLX_IDinst__n0086<30>6  (
    .ADR0(DLX_IDinst_branch_address[30]),
    .ADR1(DLX_IDinst_EPC[30]),
    .ADR2(DLX_IDinst__n0071),
    .ADR3(DLX_IDinst_N70786),
    .O(\CHOICE2657/GROM )
  );
  X_BUF \CHOICE2657/XUSED  (
    .I(\CHOICE2657/FROM ),
    .O(CHOICE2657)
  );
  X_BUF \CHOICE2657/YUSED  (
    .I(\CHOICE2657/GROM ),
    .O(CHOICE2789)
  );
  defparam \DLX_EXinst__n0017<17>1 .INIT = 16'hECA0;
  X_LUT4 \DLX_EXinst__n0017<17>1  (
    .ADR0(N100440),
    .ADR1(DLX_EXinst__n0030_1),
    .ADR2(\DLX_IDinst_Imm[31] ),
    .ADR3(DLX_IDinst_reg_out_B[17]),
    .O(\DLX_EXinst__n0017<17>/FROM )
  );
  defparam \DLX_EXinst__n0017<30>1 .INIT = 16'hEAC0;
  X_LUT4 \DLX_EXinst__n0017<30>1  (
    .ADR0(N100440),
    .ADR1(DLX_IDinst_reg_out_B[30]),
    .ADR2(DLX_EXinst__n0030_1),
    .ADR3(\DLX_IDinst_Imm[31] ),
    .O(\DLX_EXinst__n0017<17>/GROM )
  );
  X_BUF \DLX_EXinst__n0017<17>/XUSED  (
    .I(\DLX_EXinst__n0017<17>/FROM ),
    .O(DLX_EXinst__n0017[17])
  );
  X_BUF \DLX_EXinst__n0017<17>/YUSED  (
    .I(\DLX_EXinst__n0017<17>/GROM ),
    .O(DLX_EXinst__n0017[30])
  );
  defparam \DLX_EXinst__n0006<10>87 .INIT = 16'hFBFA;
  X_LUT4 \DLX_EXinst__n0006<10>87  (
    .ADR0(CHOICE4507),
    .ADR1(N109130),
    .ADR2(CHOICE4492),
    .ADR3(CHOICE4487),
    .O(\CHOICE4508/FROM )
  );
  defparam \DLX_EXinst__n0006<9>87 .INIT = 16'hFDFC;
  X_LUT4 \DLX_EXinst__n0006<9>87  (
    .ADR0(N109130),
    .ADR1(CHOICE4569),
    .ADR2(CHOICE4554),
    .ADR3(CHOICE4549),
    .O(\CHOICE4508/GROM )
  );
  X_BUF \CHOICE4508/XUSED  (
    .I(\CHOICE4508/FROM ),
    .O(CHOICE4508)
  );
  X_BUF \CHOICE4508/YUSED  (
    .I(\CHOICE4508/GROM ),
    .O(CHOICE4570)
  );
  defparam \vga_top_vga1_blueout<2>1 .INIT = 16'h000A;
  X_LUT4 \vga_top_vga1_blueout<2>1  (
    .ADR0(vga_top_vga1_videoon),
    .ADR1(VCC),
    .ADR2(vram_out_vga_eff),
    .ADR3(reset_IBUF_1),
    .O(\blue_2_OBUF/FROM )
  );
  defparam \vga_top_vga1_greenout<0>1 .INIT = 16'h0050;
  X_LUT4 \vga_top_vga1_greenout<0>1  (
    .ADR0(vram_out_vga_eff),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_videoon),
    .ADR3(reset_IBUF_1),
    .O(\blue_2_OBUF/GROM )
  );
  X_BUF \blue_2_OBUF/XUSED  (
    .I(\blue_2_OBUF/FROM ),
    .O(blue_2_OBUF)
  );
  X_BUF \blue_2_OBUF/YUSED  (
    .I(\blue_2_OBUF/GROM ),
    .O(green_0_OBUF)
  );
  defparam \DLX_IDinst__n0086<2>6 .INIT = 16'hEAC0;
  X_LUT4 \DLX_IDinst__n0086<2>6  (
    .ADR0(DLX_IDinst_EPC[2]),
    .ADR1(DLX_IDinst_N70786),
    .ADR2(DLX_IDinst_branch_address[2]),
    .ADR3(DLX_IDinst__n0071),
    .O(\CHOICE2569/FROM )
  );
  defparam \DLX_IDinst__n0086<15>6 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst__n0086<15>6  (
    .ADR0(DLX_IDinst_EPC[15]),
    .ADR1(DLX_IDinst__n0071),
    .ADR2(DLX_IDinst_branch_address[15]),
    .ADR3(DLX_IDinst_N70786),
    .O(\CHOICE2569/GROM )
  );
  X_BUF \CHOICE2569/XUSED  (
    .I(\CHOICE2569/FROM ),
    .O(CHOICE2569)
  );
  X_BUF \CHOICE2569/YUSED  (
    .I(\CHOICE2569/GROM ),
    .O(CHOICE2723)
  );
  defparam \DLX_EXinst__n0017<18>1 .INIT = 16'hECA0;
  X_LUT4 \DLX_EXinst__n0017<18>1  (
    .ADR0(N100440),
    .ADR1(DLX_IDinst_reg_out_B[18]),
    .ADR2(\DLX_IDinst_Imm[31] ),
    .ADR3(DLX_EXinst__n0030_1),
    .O(\DLX_EXinst__n0017<18>/FROM )
  );
  defparam \DLX_EXinst__n0017<23>1 .INIT = 16'hF888;
  X_LUT4 \DLX_EXinst__n0017<23>1  (
    .ADR0(N100440),
    .ADR1(\DLX_IDinst_Imm[31] ),
    .ADR2(DLX_IDinst_reg_out_B[23]),
    .ADR3(DLX_EXinst__n0030_1),
    .O(\DLX_EXinst__n0017<18>/GROM )
  );
  X_BUF \DLX_EXinst__n0017<18>/XUSED  (
    .I(\DLX_EXinst__n0017<18>/FROM ),
    .O(DLX_EXinst__n0017[18])
  );
  X_BUF \DLX_EXinst__n0017<18>/YUSED  (
    .I(\DLX_EXinst__n0017<18>/GROM ),
    .O(DLX_EXinst__n0017[23])
  );
  defparam \DLX_EXinst__n0017<28>1 .INIT = 16'hEAC0;
  X_LUT4 \DLX_EXinst__n0017<28>1  (
    .ADR0(\DLX_IDinst_Imm[31] ),
    .ADR1(DLX_IDinst_reg_out_B[28]),
    .ADR2(DLX_EXinst__n0030_1),
    .ADR3(N100440),
    .O(\DLX_EXinst__n0017<28>/FROM )
  );
  defparam \DLX_EXinst__n0017<31>1 .INIT = 16'hF888;
  X_LUT4 \DLX_EXinst__n0017<31>1  (
    .ADR0(\DLX_IDinst_Imm[31] ),
    .ADR1(N100440),
    .ADR2(DLX_EXinst__n0030_1),
    .ADR3(DLX_IDinst_reg_out_B[31]),
    .O(\DLX_EXinst__n0017<28>/GROM )
  );
  X_BUF \DLX_EXinst__n0017<28>/XUSED  (
    .I(\DLX_EXinst__n0017<28>/FROM ),
    .O(DLX_EXinst__n0017[28])
  );
  X_BUF \DLX_EXinst__n0017<28>/YUSED  (
    .I(\DLX_EXinst__n0017<28>/GROM ),
    .O(DLX_EXinst__n0017[31])
  );
  defparam \DLX_EXinst_Mshift__n0025_Sh<1>1 .INIT = 16'h0C0A;
  X_LUT4 \DLX_EXinst_Mshift__n0025_Sh<1>1  (
    .ADR0(DLX_IDinst_reg_out_A[1]),
    .ADR1(DLX_IDinst_reg_out_A[0]),
    .ADR2(DLX_IDinst_reg_out_B[1]),
    .ADR3(DLX_IDinst_reg_out_B[0]),
    .O(\DLX_EXinst_Mshift__n0025_Sh<1>/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0025_Sh<0>1 .INIT = 16'h0300;
  X_LUT4 \DLX_EXinst_Mshift__n0025_Sh<0>1  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(DLX_IDinst_reg_out_B[0]),
    .ADR3(DLX_IDinst_reg_out_A[0]),
    .O(\DLX_EXinst_Mshift__n0025_Sh<1>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0025_Sh<1>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0025_Sh<1>/FROM ),
    .O(\DLX_EXinst_Mshift__n0025_Sh[1] )
  );
  X_BUF \DLX_EXinst_Mshift__n0025_Sh<1>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0025_Sh<1>/GROM ),
    .O(\DLX_EXinst_Mshift__n0025_Sh[0] )
  );
  defparam \DLX_IDinst__n0086<0>25 .INIT = 16'hAABA;
  X_LUT4 \DLX_IDinst__n0086<0>25  (
    .ADR0(CHOICE2562),
    .ADR1(DLX_IDinst_N70918),
    .ADR2(CHOICE2558),
    .ADR3(DLX_IDinst__n0364),
    .O(\DLX_IDinst_branch_address<0>/FROM )
  );
  defparam \DLX_IDinst__n0086<0>31 .INIT = 16'hFFA0;
  X_LUT4 \DLX_IDinst__n0086<0>31  (
    .ADR0(DLX_IDinst__n0128[0]),
    .ADR1(VCC),
    .ADR2(N100609),
    .ADR3(CHOICE2563),
    .O(N105098)
  );
  X_BUF \DLX_IDinst_branch_address<0>/XUSED  (
    .I(\DLX_IDinst_branch_address<0>/FROM ),
    .O(CHOICE2563)
  );
  defparam \DLX_IDinst__n0086<3>6 .INIT = 16'hECA0;
  X_LUT4 \DLX_IDinst__n0086<3>6  (
    .ADR0(DLX_IDinst_branch_address[3]),
    .ADR1(DLX_IDinst__n0071),
    .ADR2(DLX_IDinst_N70786),
    .ADR3(DLX_IDinst_EPC[3]),
    .O(\CHOICE2591/FROM )
  );
  defparam \DLX_IDinst__n0086<24>6 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst__n0086<24>6  (
    .ADR0(DLX_IDinst_branch_address[24]),
    .ADR1(DLX_IDinst_N70786),
    .ADR2(DLX_IDinst__n0071),
    .ADR3(DLX_IDinst_EPC[24]),
    .O(\CHOICE2591/GROM )
  );
  X_BUF \CHOICE2591/XUSED  (
    .I(\CHOICE2591/FROM ),
    .O(CHOICE2591)
  );
  X_BUF \CHOICE2591/YUSED  (
    .I(\CHOICE2591/GROM ),
    .O(CHOICE2833)
  );
  defparam \DLX_IDinst__n0086<28>6 .INIT = 16'hEAC0;
  X_LUT4 \DLX_IDinst__n0086<28>6  (
    .ADR0(DLX_IDinst_branch_address[28]),
    .ADR1(DLX_IDinst__n0071),
    .ADR2(DLX_IDinst_EPC[28]),
    .ADR3(DLX_IDinst_N70786),
    .O(\CHOICE2888/FROM )
  );
  defparam \DLX_IDinst__n0086<16>6 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst__n0086<16>6  (
    .ADR0(DLX_IDinst__n0071),
    .ADR1(DLX_IDinst_EPC[16]),
    .ADR2(DLX_IDinst_N70786),
    .ADR3(DLX_IDinst_branch_address[16]),
    .O(\CHOICE2888/GROM )
  );
  X_BUF \CHOICE2888/XUSED  (
    .I(\CHOICE2888/FROM ),
    .O(CHOICE2888)
  );
  X_BUF \CHOICE2888/YUSED  (
    .I(\CHOICE2888/GROM ),
    .O(CHOICE2734)
  );
  defparam \DLX_EXinst__n0006<17>410_SW0 .INIT = 16'h3332;
  X_LUT4 \DLX_EXinst__n0006<17>410_SW0  (
    .ADR0(CHOICE5574),
    .ADR1(DLX_EXinst__n0030),
    .ADR2(CHOICE5577),
    .ADR3(CHOICE5606),
    .O(\DLX_EXinst_ALU_result<17>/FROM )
  );
  defparam \DLX_EXinst__n0006<17>410 .INIT = 16'hF0E0;
  X_LUT4 \DLX_EXinst__n0006<17>410  (
    .ADR0(CHOICE5648),
    .ADR1(N100490),
    .ADR2(DLX_EXinst__n0149),
    .ADR3(N126601),
    .O(N123529)
  );
  X_BUF \DLX_EXinst_ALU_result<17>/XUSED  (
    .I(\DLX_EXinst_ALU_result<17>/FROM ),
    .O(N126601)
  );
  defparam \DLX_EXinst__n0006<25>306_SW0 .INIT = 16'h00FE;
  X_LUT4 \DLX_EXinst__n0006<25>306_SW0  (
    .ADR0(CHOICE4740),
    .ADR1(CHOICE4741),
    .ADR2(CHOICE4766),
    .ADR3(DLX_EXinst__n0030),
    .O(\DLX_EXinst_ALU_result<25>/FROM )
  );
  defparam \DLX_EXinst__n0006<25>306 .INIT = 16'hAAA8;
  X_LUT4 \DLX_EXinst__n0006<25>306  (
    .ADR0(DLX_EXinst__n0149),
    .ADR1(CHOICE4798),
    .ADR2(N100490),
    .ADR3(N126276),
    .O(N118327)
  );
  X_BUF \DLX_EXinst_ALU_result<25>/XUSED  (
    .I(\DLX_EXinst_ALU_result<25>/FROM ),
    .O(N126276)
  );
  defparam \vga_top_vga1_blueout<1>1 .INIT = 16'h0022;
  X_LUT4 \vga_top_vga1_blueout<1>1  (
    .ADR0(vga_top_vga1_videoon),
    .ADR1(vram_out_vga_eff),
    .ADR2(VCC),
    .ADR3(reset_IBUF_1),
    .O(\blue_1_OBUF/FROM )
  );
  defparam \vga_top_vga1_greenout<2>1 .INIT = 16'h0404;
  X_LUT4 \vga_top_vga1_greenout<2>1  (
    .ADR0(reset_IBUF_1),
    .ADR1(vga_top_vga1_videoon),
    .ADR2(vram_out_vga_eff),
    .ADR3(VCC),
    .O(\blue_1_OBUF/GROM )
  );
  X_BUF \blue_1_OBUF/XUSED  (
    .I(\blue_1_OBUF/FROM ),
    .O(blue_1_OBUF)
  );
  X_BUF \blue_1_OBUF/YUSED  (
    .I(\blue_1_OBUF/GROM ),
    .O(green_2_OBUF)
  );
  defparam DLX_EXlc_slave_ctrlEX__n00021.INIT = 16'h0032;
  X_LUT4 DLX_EXlc_slave_ctrlEX__n00021 (
    .ADR0(DLX_MEMlc_master_ctrlMEM_l),
    .ADR1(DLX_EXlc_slave_ctrlEX_l),
    .ADR2(DLX_reqout_EX),
    .ADR3(reset_IBUF),
    .O(\DLX_reqout_EX/GROM )
  );
  X_BUF \DLX_reqout_EX/YUSED  (
    .I(\DLX_reqout_EX/GROM ),
    .O(DLX_reqout_EX)
  );
  defparam \DLX_IDinst__n0086<1>6 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst__n0086<1>6  (
    .ADR0(DLX_IDinst_N70786),
    .ADR1(DLX_IDinst_branch_address[1]),
    .ADR2(DLX_IDinst__n0071),
    .ADR3(DLX_IDinst_EPC[1]),
    .O(\CHOICE2580/FROM )
  );
  defparam \DLX_IDinst__n0086<17>6 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst__n0086<17>6  (
    .ADR0(DLX_IDinst__n0071),
    .ADR1(DLX_IDinst_EPC[17]),
    .ADR2(DLX_IDinst_N70786),
    .ADR3(DLX_IDinst_branch_address[17]),
    .O(\CHOICE2580/GROM )
  );
  X_BUF \CHOICE2580/XUSED  (
    .I(\CHOICE2580/FROM ),
    .O(CHOICE2580)
  );
  X_BUF \CHOICE2580/YUSED  (
    .I(\CHOICE2580/GROM ),
    .O(CHOICE2745)
  );
  defparam \DLX_IDinst__n0086<29>6 .INIT = 16'hECA0;
  X_LUT4 \DLX_IDinst__n0086<29>6  (
    .ADR0(DLX_IDinst_N70786),
    .ADR1(DLX_IDinst__n0071),
    .ADR2(DLX_IDinst_branch_address[29]),
    .ADR3(DLX_IDinst_EPC[29]),
    .O(\CHOICE2899/FROM )
  );
  defparam \DLX_IDinst__n0086<25>6 .INIT = 16'hECA0;
  X_LUT4 \DLX_IDinst__n0086<25>6  (
    .ADR0(DLX_IDinst_N70786),
    .ADR1(DLX_IDinst_EPC[25]),
    .ADR2(DLX_IDinst_branch_address[25]),
    .ADR3(DLX_IDinst__n0071),
    .O(\CHOICE2899/GROM )
  );
  X_BUF \CHOICE2899/XUSED  (
    .I(\CHOICE2899/FROM ),
    .O(CHOICE2899)
  );
  X_BUF \CHOICE2899/YUSED  (
    .I(\CHOICE2899/GROM ),
    .O(CHOICE2855)
  );
  defparam \DLX_EXinst__n0017<27>1 .INIT = 16'hF888;
  X_LUT4 \DLX_EXinst__n0017<27>1  (
    .ADR0(DLX_EXinst__n0030_1),
    .ADR1(DLX_IDinst_reg_out_B[27]),
    .ADR2(\DLX_IDinst_Imm[31] ),
    .ADR3(N100440),
    .O(\DLX_EXinst__n0017<27>/FROM )
  );
  defparam \DLX_EXinst__n0017<25>1 .INIT = 16'hECA0;
  X_LUT4 \DLX_EXinst__n0017<25>1  (
    .ADR0(DLX_IDinst_reg_out_B[25]),
    .ADR1(\DLX_IDinst_Imm[31] ),
    .ADR2(DLX_EXinst__n0030_1),
    .ADR3(N100440),
    .O(\DLX_EXinst__n0017<27>/GROM )
  );
  X_BUF \DLX_EXinst__n0017<27>/XUSED  (
    .I(\DLX_EXinst__n0017<27>/FROM ),
    .O(DLX_EXinst__n0017[27])
  );
  X_BUF \DLX_EXinst__n0017<27>/YUSED  (
    .I(\DLX_EXinst__n0017<27>/GROM ),
    .O(DLX_EXinst__n0017[25])
  );
  defparam vga_top_vga1__n00094.INIT = 16'hFFFE;
  X_LUT4 vga_top_vga1__n00094 (
    .ADR0(vga_top_vga1_vcounter[5]),
    .ADR1(vga_top_vga1_vcounter[3]),
    .ADR2(vga_top_vga1_vcounter[2]),
    .ADR3(vga_top_vga1_vcounter[4]),
    .O(\CHOICE3412/FROM )
  );
  defparam vga_top_vga1__n0007_SW0.INIT = 16'hFF7F;
  X_LUT4 vga_top_vga1__n0007_SW0 (
    .ADR0(vga_top_vga1_vcounter[1]),
    .ADR1(vga_top_vga1_vcounter[2]),
    .ADR2(vga_top_vga1_vcounter[3]),
    .ADR3(vga_top_vga1_vcounter[0]),
    .O(\CHOICE3412/GROM )
  );
  X_BUF \CHOICE3412/XUSED  (
    .I(\CHOICE3412/FROM ),
    .O(CHOICE3412)
  );
  X_BUF \CHOICE3412/YUSED  (
    .I(\CHOICE3412/GROM ),
    .O(N100333)
  );
  defparam \DLX_IDinst__n0086<1>25 .INIT = 16'hCCDC;
  X_LUT4 \DLX_IDinst__n0086<1>25  (
    .ADR0(DLX_IDinst_N70918),
    .ADR1(CHOICE2584),
    .ADR2(CHOICE2580),
    .ADR3(DLX_IDinst__n0364),
    .O(\DLX_IDinst_branch_address<1>/FROM )
  );
  defparam \DLX_IDinst__n0086<1>31 .INIT = 16'hFF88;
  X_LUT4 \DLX_IDinst__n0086<1>31  (
    .ADR0(DLX_IDinst__n0128[1]),
    .ADR1(N100609),
    .ADR2(VCC),
    .ADR3(CHOICE2585),
    .O(N105224)
  );
  X_BUF \DLX_IDinst_branch_address<1>/XUSED  (
    .I(\DLX_IDinst_branch_address<1>/FROM ),
    .O(CHOICE2585)
  );
  defparam \DLX_IDinst__n0086<4>6 .INIT = 16'hECA0;
  X_LUT4 \DLX_IDinst__n0086<4>6  (
    .ADR0(DLX_IDinst_branch_address[4]),
    .ADR1(DLX_IDinst__n0071),
    .ADR2(DLX_IDinst_N70786),
    .ADR3(DLX_IDinst_EPC[4]),
    .O(\CHOICE2602/FROM )
  );
  defparam \DLX_IDinst__n0086<18>6 .INIT = 16'hEAC0;
  X_LUT4 \DLX_IDinst__n0086<18>6  (
    .ADR0(DLX_IDinst_N70786),
    .ADR1(DLX_IDinst_EPC[18]),
    .ADR2(DLX_IDinst__n0071),
    .ADR3(DLX_IDinst_branch_address[18]),
    .O(\CHOICE2602/GROM )
  );
  X_BUF \CHOICE2602/XUSED  (
    .I(\CHOICE2602/FROM ),
    .O(CHOICE2602)
  );
  X_BUF \CHOICE2602/YUSED  (
    .I(\CHOICE2602/GROM ),
    .O(CHOICE2767)
  );
  defparam \DLX_IDinst__n0086<5>6 .INIT = 16'hECA0;
  X_LUT4 \DLX_IDinst__n0086<5>6  (
    .ADR0(DLX_IDinst_branch_address[5]),
    .ADR1(DLX_IDinst_EPC[5]),
    .ADR2(DLX_IDinst_N70786),
    .ADR3(DLX_IDinst__n0071),
    .O(\CHOICE2613/FROM )
  );
  defparam \DLX_IDinst__n0086<26>6 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst__n0086<26>6  (
    .ADR0(DLX_IDinst_N70786),
    .ADR1(DLX_IDinst_branch_address[26]),
    .ADR2(DLX_IDinst_EPC[26]),
    .ADR3(DLX_IDinst__n0071),
    .O(\CHOICE2613/GROM )
  );
  X_BUF \CHOICE2613/XUSED  (
    .I(\CHOICE2613/FROM ),
    .O(CHOICE2613)
  );
  X_BUF \CHOICE2613/YUSED  (
    .I(\CHOICE2613/GROM ),
    .O(CHOICE2866)
  );
  defparam \DLX_EXinst__n0017<29>1 .INIT = 16'hEAC0;
  X_LUT4 \DLX_EXinst__n0017<29>1  (
    .ADR0(N100440),
    .ADR1(DLX_EXinst__n0030_1),
    .ADR2(DLX_IDinst_reg_out_B[29]),
    .ADR3(\DLX_IDinst_Imm[31] ),
    .O(\DLX_EXinst__n0017<29>/FROM )
  );
  defparam \DLX_EXinst__n0017<26>1 .INIT = 16'hECA0;
  X_LUT4 \DLX_EXinst__n0017<26>1  (
    .ADR0(\DLX_IDinst_Imm[31] ),
    .ADR1(DLX_EXinst__n0030_1),
    .ADR2(N100440),
    .ADR3(DLX_IDinst_reg_out_B[26]),
    .O(\DLX_EXinst__n0017<29>/GROM )
  );
  X_BUF \DLX_EXinst__n0017<29>/XUSED  (
    .I(\DLX_EXinst__n0017<29>/FROM ),
    .O(DLX_EXinst__n0017[29])
  );
  X_BUF \DLX_EXinst__n0017<29>/YUSED  (
    .I(\DLX_EXinst__n0017<29>/GROM ),
    .O(DLX_EXinst__n0017[26])
  );
  defparam DLX_EXinst_Ker6624854_SW0.INIT = 16'h0A00;
  X_LUT4 DLX_EXinst_Ker6624854_SW0 (
    .ADR0(DLX_EXinst_N66112),
    .ADR1(VCC),
    .ADR2(\DLX_IDinst_Imm[31] ),
    .ADR3(DLX_IDinst_IR_opcode_field[1]),
    .O(\N125999/FROM )
  );
  defparam \DLX_EXinst__n0017<19>1 .INIT = 16'hEAC0;
  X_LUT4 \DLX_EXinst__n0017<19>1  (
    .ADR0(\DLX_IDinst_Imm[31] ),
    .ADR1(DLX_EXinst__n0030_1),
    .ADR2(DLX_IDinst_reg_out_B[19]),
    .ADR3(N100440),
    .O(\N125999/GROM )
  );
  X_BUF \N125999/XUSED  (
    .I(\N125999/FROM ),
    .O(N125999)
  );
  X_BUF \N125999/YUSED  (
    .I(\N125999/GROM ),
    .O(DLX_EXinst__n0017[19])
  );
  defparam \DLX_IDinst__n0086<2>25 .INIT = 16'hCCCE;
  X_LUT4 \DLX_IDinst__n0086<2>25  (
    .ADR0(CHOICE2569),
    .ADR1(CHOICE2573),
    .ADR2(DLX_IDinst__n0364),
    .ADR3(DLX_IDinst_N70918),
    .O(\DLX_IDinst_branch_address<2>/FROM )
  );
  defparam \DLX_IDinst__n0086<2>31 .INIT = 16'hFFA0;
  X_LUT4 \DLX_IDinst__n0086<2>31  (
    .ADR0(DLX_IDinst__n0128[2]),
    .ADR1(VCC),
    .ADR2(N100609),
    .ADR3(CHOICE2574),
    .O(N105161)
  );
  X_BUF \DLX_IDinst_branch_address<2>/XUSED  (
    .I(\DLX_IDinst_branch_address<2>/FROM ),
    .O(CHOICE2574)
  );
  defparam DLX_IDinst__n0339116.INIT = 16'h0033;
  X_LUT4 DLX_IDinst__n0339116 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_IR_latched[28]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_IR_latched[30]),
    .O(\CHOICE1410/FROM )
  );
  defparam DLX_IDinst__n0339120.INIT = 16'hD000;
  X_LUT4 DLX_IDinst__n0339120 (
    .ADR0(DLX_IDinst_IR_latched[27]),
    .ADR1(DLX_IDinst_IR_latched[26]),
    .ADR2(DLX_IDinst_IR_latched[31]),
    .ADR3(CHOICE1410),
    .O(\CHOICE1410/GROM )
  );
  X_BUF \CHOICE1410/XUSED  (
    .I(\CHOICE1410/FROM ),
    .O(CHOICE1410)
  );
  X_BUF \CHOICE1410/YUSED  (
    .I(\CHOICE1410/GROM ),
    .O(CHOICE1411)
  );
  defparam \DLX_EXinst__n0006<24>91_SW0 .INIT = 16'hAE0C;
  X_LUT4 \DLX_EXinst__n0006<24>91_SW0  (
    .ADR0(DLX_EXinst__n0077),
    .ADR1(N98127),
    .ADR2(DLX_IDinst_IR_function_field[4]),
    .ADR3(\DLX_IDinst_Imm[8] ),
    .O(\N126597/FROM )
  );
  defparam \DLX_EXinst__n0006<22>100_SW0 .INIT = 16'hF222;
  X_LUT4 \DLX_EXinst__n0006<22>100_SW0  (
    .ADR0(N108101),
    .ADR1(DLX_IDinst_IR_function_field[4]),
    .ADR2(DLX_EXinst__n0077),
    .ADR3(\DLX_IDinst_Imm[6] ),
    .O(\N126597/GROM )
  );
  X_BUF \N126597/XUSED  (
    .I(\N126597/FROM ),
    .O(N126597)
  );
  X_BUF \N126597/YUSED  (
    .I(\N126597/GROM ),
    .O(N126524)
  );
  defparam \DLX_IDinst__n0086<27>20 .INIT = 16'hCC00;
  X_LUT4 \DLX_IDinst__n0086<27>20  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_N70295),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_regA_eff[27]),
    .O(\CHOICE2881/FROM )
  );
  defparam \DLX_IDinst__n0086<3>20 .INIT = 16'hC0C0;
  X_LUT4 \DLX_IDinst__n0086<3>20  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_N70295),
    .ADR2(DLX_IDinst_regA_eff[3]),
    .ADR3(VCC),
    .O(\CHOICE2881/GROM )
  );
  X_BUF \CHOICE2881/XUSED  (
    .I(\CHOICE2881/FROM ),
    .O(CHOICE2881)
  );
  X_BUF \CHOICE2881/YUSED  (
    .I(\CHOICE2881/GROM ),
    .O(CHOICE2595)
  );
  defparam DLX_IDinst__n0339126.INIT = 16'hAFAE;
  X_LUT4 DLX_IDinst__n0339126 (
    .ADR0(CHOICE1411),
    .ADR1(CHOICE1402),
    .ADR2(DLX_IDinst_IR_latched[31]),
    .ADR3(CHOICE1387),
    .O(\N98420/FROM )
  );
  defparam DLX_IDinst__n03471.INIT = 16'hFAF0;
  X_LUT4 DLX_IDinst__n03471 (
    .ADR0(DLX_IDinst_N70663),
    .ADR1(VCC),
    .ADR2(N98806),
    .ADR3(N98420),
    .O(\N98420/GROM )
  );
  X_BUF \N98420/XUSED  (
    .I(\N98420/FROM ),
    .O(N98420)
  );
  X_BUF \N98420/YUSED  (
    .I(\N98420/GROM ),
    .O(DLX_IDinst__n0347)
  );
  defparam DLX_IDinst_Ker703311.INIT = 16'hF3F3;
  X_LUT4 DLX_IDinst_Ker703311 (
    .ADR0(VCC),
    .ADR1(INT_IBUF),
    .ADR2(DLX_IDinst_CLI),
    .ADR3(VCC),
    .O(\DLX_IDinst_N70333/GROM )
  );
  X_BUF \DLX_IDinst_N70333/YUSED  (
    .I(\DLX_IDinst_N70333/GROM ),
    .O(DLX_IDinst_N70333)
  );
  defparam \DLX_IDinst__n0086<3>25 .INIT = 16'hF0F2;
  X_LUT4 \DLX_IDinst__n0086<3>25  (
    .ADR0(CHOICE2591),
    .ADR1(DLX_IDinst_N70918),
    .ADR2(CHOICE2595),
    .ADR3(DLX_IDinst__n0364),
    .O(\DLX_IDinst_branch_address<3>/FROM )
  );
  defparam \DLX_IDinst__n0086<3>31 .INIT = 16'hFF88;
  X_LUT4 \DLX_IDinst__n0086<3>31  (
    .ADR0(N100609),
    .ADR1(DLX_IDinst__n0128[3]),
    .ADR2(VCC),
    .ADR3(CHOICE2596),
    .O(N105287)
  );
  X_BUF \DLX_IDinst_branch_address<3>/XUSED  (
    .I(\DLX_IDinst_branch_address<3>/FROM ),
    .O(CHOICE2596)
  );
  defparam DLX_IDinst_Ker703261.INIT = 16'hF888;
  X_LUT4 DLX_IDinst_Ker703261 (
    .ADR0(DLX_IDinst__n0250),
    .ADR1(DLX_IDinst_N70885),
    .ADR2(DLX_IDinst_IR_latched[30]),
    .ADR3(DLX_IDinst_N70918),
    .O(\DLX_IDinst_N70328/FROM )
  );
  defparam \DLX_IDinst__n0086<31>27_SW0 .INIT = 16'hECA0;
  X_LUT4 \DLX_IDinst__n0086<31>27_SW0  (
    .ADR0(DLX_IDinst_N70072),
    .ADR1(DLX_IDinst_regA_eff[31]),
    .ADR2(DLX_IDinst__n0128[31]),
    .ADR3(DLX_IDinst_N70328),
    .O(\DLX_IDinst_N70328/GROM )
  );
  X_BUF \DLX_IDinst_N70328/XUSED  (
    .I(\DLX_IDinst_N70328/FROM ),
    .O(DLX_IDinst_N70328)
  );
  X_BUF \DLX_IDinst_N70328/YUSED  (
    .I(\DLX_IDinst_N70328/GROM ),
    .O(N127435)
  );
  defparam \DLX_IDinst__n0086<4>25 .INIT = 16'hF1F0;
  X_LUT4 \DLX_IDinst__n0086<4>25  (
    .ADR0(DLX_IDinst_N70918),
    .ADR1(DLX_IDinst__n0364),
    .ADR2(CHOICE2606),
    .ADR3(CHOICE2602),
    .O(\DLX_IDinst_branch_address<4>/FROM )
  );
  defparam \DLX_IDinst__n0086<4>31 .INIT = 16'hFFC0;
  X_LUT4 \DLX_IDinst__n0086<4>31  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst__n0128[4]),
    .ADR2(N100609),
    .ADR3(CHOICE2607),
    .O(N105350)
  );
  X_BUF \DLX_IDinst_branch_address<4>/XUSED  (
    .I(\DLX_IDinst_branch_address<4>/FROM ),
    .O(CHOICE2607)
  );
  defparam DLX_IDinst_Ker69912_SW0.INIT = 16'h7F6F;
  X_LUT4 DLX_IDinst_Ker69912_SW0 (
    .ADR0(DLX_IDinst_IR_latched[26]),
    .ADR1(DLX_IDinst_IR_latched[31]),
    .ADR2(DLX_IDinst__n0387),
    .ADR3(DLX_IDinst__n03641_1),
    .O(\N100688/FROM )
  );
  defparam DLX_IDinst_Ker69912.INIT = 16'h5545;
  X_LUT4 DLX_IDinst_Ker69912 (
    .ADR0(DLX_IDinst__n0151),
    .ADR1(DLX_IDinst__n0331),
    .ADR2(DLX_IDinst_N70673),
    .ADR3(N100688),
    .O(\N100688/GROM )
  );
  X_BUF \N100688/XUSED  (
    .I(\N100688/FROM ),
    .O(N100688)
  );
  X_BUF \N100688/YUSED  (
    .I(\N100688/GROM ),
    .O(DLX_IDinst_N69914)
  );
  defparam \DLX_IDinst__n0086<5>25 .INIT = 16'hCCDC;
  X_LUT4 \DLX_IDinst__n0086<5>25  (
    .ADR0(DLX_IDinst__n0364),
    .ADR1(CHOICE2617),
    .ADR2(CHOICE2613),
    .ADR3(DLX_IDinst_N70918),
    .O(\DLX_IDinst_branch_address<5>/FROM )
  );
  defparam \DLX_IDinst__n0086<5>31 .INIT = 16'hFFC0;
  X_LUT4 \DLX_IDinst__n0086<5>31  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst__n0128[5]),
    .ADR2(N100609),
    .ADR3(CHOICE2618),
    .O(N105413)
  );
  X_BUF \DLX_IDinst_branch_address<5>/XUSED  (
    .I(\DLX_IDinst_branch_address<5>/FROM ),
    .O(CHOICE2618)
  );
  defparam DLX_IDinst_Ker706211.INIT = 16'h00AA;
  X_LUT4 DLX_IDinst_Ker706211 (
    .ADR0(DLX_IDinst_N70909),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_IR_latched[28]),
    .O(\DLX_IDinst_N70623/FROM )
  );
  defparam DLX_IDinst__n00701.INIT = 16'h0800;
  X_LUT4 DLX_IDinst__n00701 (
    .ADR0(DLX_IDinst_IR_latched[30]),
    .ADR1(DLX_IDinst_IR_latched[26]),
    .ADR2(DLX_IDinst_IR_latched[27]),
    .ADR3(DLX_IDinst_N70623),
    .O(\DLX_IDinst_N70623/GROM )
  );
  X_BUF \DLX_IDinst_N70623/XUSED  (
    .I(\DLX_IDinst_N70623/FROM ),
    .O(DLX_IDinst_N70623)
  );
  X_BUF \DLX_IDinst_N70623/YUSED  (
    .I(\DLX_IDinst_N70623/GROM ),
    .O(DLX_IDinst__n0070)
  );
  defparam \DLX_IDinst__n0086<6>25 .INIT = 16'hCCCE;
  X_LUT4 \DLX_IDinst__n0086<6>25  (
    .ADR0(CHOICE2635),
    .ADR1(CHOICE2639),
    .ADR2(DLX_IDinst__n0364),
    .ADR3(DLX_IDinst_N70918),
    .O(\DLX_IDinst_branch_address<6>/FROM )
  );
  defparam \DLX_IDinst__n0086<6>31 .INIT = 16'hFFC0;
  X_LUT4 \DLX_IDinst__n0086<6>31  (
    .ADR0(VCC),
    .ADR1(N100609),
    .ADR2(DLX_IDinst__n0128[6]),
    .ADR3(CHOICE2640),
    .O(N105535)
  );
  X_BUF \DLX_IDinst_branch_address<6>/XUSED  (
    .I(\DLX_IDinst_branch_address<6>/FROM ),
    .O(CHOICE2640)
  );
  defparam \DLX_IDinst__n0086<7>11 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst__n0086<7>11  (
    .ADR0(DLX_IDinst__n0071),
    .ADR1(DLX_IDinst_EPC[7]),
    .ADR2(DLX_IDinst_branch_address[7]),
    .ADR3(DLX_IDinst_N70786),
    .O(\DLX_IDinst_branch_address<7>/FROM )
  );
  defparam \DLX_IDinst__n0086<7>27 .INIT = 16'hAFAE;
  X_LUT4 \DLX_IDinst__n0086<7>27  (
    .ADR0(N127423),
    .ADR1(DLX_IDinst__n0364),
    .ADR2(DLX_IDinst_N70918),
    .ADR3(CHOICE2627),
    .O(N105474)
  );
  X_BUF \DLX_IDinst_branch_address<7>/XUSED  (
    .I(\DLX_IDinst_branch_address<7>/FROM ),
    .O(CHOICE2627)
  );
  defparam DLX_IDinst__n02521.INIT = 16'h0001;
  X_LUT4 DLX_IDinst__n02521 (
    .ADR0(DLX_IDinst_IR_latched[30]),
    .ADR1(DLX_IDinst_IR_latched[27]),
    .ADR2(DLX_IDinst_IR_latched[26]),
    .ADR3(DLX_IDinst_IR_latched[28]),
    .O(\DLX_IDinst__n0252/FROM )
  );
  defparam DLX_IDinst_Ker706331.INIT = 16'h0022;
  X_LUT4 DLX_IDinst_Ker706331 (
    .ADR0(DLX_IDinst_IR_latched[28]),
    .ADR1(DLX_IDinst_IR_latched[27]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_IR_latched[30]),
    .O(\DLX_IDinst__n0252/GROM )
  );
  X_BUF \DLX_IDinst__n0252/XUSED  (
    .I(\DLX_IDinst__n0252/FROM ),
    .O(DLX_IDinst__n0252)
  );
  X_BUF \DLX_IDinst__n0252/YUSED  (
    .I(\DLX_IDinst__n0252/GROM ),
    .O(DLX_IDinst_N70635)
  );
  defparam DLX_IDinst_Ker707141.INIT = 16'h0077;
  X_LUT4 DLX_IDinst_Ker707141 (
    .ADR0(DLX_MEMinst_reg_write_MEM),
    .ADR1(DLX_IDinst__n0315),
    .ADR2(VCC),
    .ADR3(DLX_IDinst__n0004),
    .O(\DLX_IDinst_N70716/FROM )
  );
  defparam \DLX_IDinst_regB_eff<0>1 .INIT = 16'hECA0;
  X_LUT4 \DLX_IDinst_regB_eff<0>1  (
    .ADR0(DLX_RF_data_in[0]),
    .ADR1(DLX_IDinst_reg_out_B_RF[0]),
    .ADR2(DLX_IDinst__n0145),
    .ADR3(DLX_IDinst_N70716),
    .O(\DLX_IDinst_N70716/GROM )
  );
  X_BUF \DLX_IDinst_N70716/XUSED  (
    .I(\DLX_IDinst_N70716/FROM ),
    .O(DLX_IDinst_N70716)
  );
  X_BUF \DLX_IDinst_N70716/YUSED  (
    .I(\DLX_IDinst_N70716/GROM ),
    .O(DLX_IDinst_regB_eff[0])
  );
  defparam \DLX_EXinst__n0006<12>15_SW0 .INIT = 16'h0033;
  X_LUT4 \DLX_EXinst__n0006<12>15_SW0  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[12]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_IR_opcode_field[0]),
    .O(\N127366/FROM )
  );
  defparam \DLX_EXinst__n0006<15>59_SW0 .INIT = 16'h0055;
  X_LUT4 \DLX_EXinst__n0006<15>59_SW0  (
    .ADR0(DLX_IDinst_reg_out_A[15]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_IR_opcode_field[0]),
    .O(\N127366/GROM )
  );
  X_BUF \N127366/XUSED  (
    .I(\N127366/FROM ),
    .O(N127366)
  );
  X_BUF \N127366/YUSED  (
    .I(\N127366/GROM ),
    .O(N127294)
  );
  defparam \DLX_EXinst__n0006<27>36_SW0 .INIT = 16'h0505;
  X_LUT4 \DLX_EXinst__n0006<27>36_SW0  (
    .ADR0(DLX_IDinst_reg_out_A[27]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_IR_opcode_field[0]),
    .ADR3(VCC),
    .O(\N127362/FROM )
  );
  defparam \DLX_EXinst__n0006<16>35_SW0 .INIT = 16'h000F;
  X_LUT4 \DLX_EXinst__n0006<16>35_SW0  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_IR_opcode_field[0]),
    .ADR3(DLX_IDinst_reg_out_A[16]),
    .O(\N127362/GROM )
  );
  X_BUF \N127362/XUSED  (
    .I(\N127362/FROM ),
    .O(N127362)
  );
  X_BUF \N127362/YUSED  (
    .I(\N127362/GROM ),
    .O(N127290)
  );
  defparam \mask<3>_SW0 .INIT = 16'hEAE0;
  X_LUT4 \mask<3>_SW0  (
    .ADR0(DLX_EXinst_ALU_result[0]),
    .ADR1(DLX_EXinst_ALU_result[1]),
    .ADR2(DLX_EXinst_byte),
    .ADR3(DLX_EXinst_word),
    .O(\N90497/FROM )
  );
  defparam \mask<3> .INIT = 16'h00F0;
  X_LUT4 \mask<3>  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(vga_select_6[0]),
    .ADR3(N90497),
    .O(\N90497/GROM )
  );
  X_BUF \N90497/XUSED  (
    .I(\N90497/FROM ),
    .O(N90497)
  );
  X_BUF \N90497/YUSED  (
    .I(\N90497/GROM ),
    .O(mask_3_OBUF)
  );
  defparam DLX_IDinst_Ker6997996.INIT = 16'h0001;
  X_LUT4 DLX_IDinst_Ker6997996 (
    .ADR0(DLX_opcode_of_MEM[0]),
    .ADR1(DLX_opcode_of_MEM[1]),
    .ADR2(DLX_opcode_of_MEM[4]),
    .ADR3(DLX_opcode_of_MEM[2]),
    .O(\CHOICE1479/FROM )
  );
  defparam DLX_IDinst_Ker706611.INIT = 16'h0300;
  X_LUT4 DLX_IDinst_Ker706611 (
    .ADR0(VCC),
    .ADR1(DLX_opcode_of_MEM[1]),
    .ADR2(DLX_opcode_of_MEM[5]),
    .ADR3(DLX_opcode_of_MEM[3]),
    .O(\CHOICE1479/GROM )
  );
  X_BUF \CHOICE1479/XUSED  (
    .I(\CHOICE1479/FROM ),
    .O(CHOICE1479)
  );
  X_BUF \CHOICE1479/YUSED  (
    .I(\CHOICE1479/GROM ),
    .O(DLX_IDinst_N70663)
  );
  defparam DLX_EXinst_Ker6628812.INIT = 16'h0004;
  X_LUT4 DLX_EXinst_Ker6628812 (
    .ADR0(DLX_IDinst_IR_opcode_field[5]),
    .ADR1(DLX_IDinst_IR_opcode_field[3]),
    .ADR2(DLX_IDinst_IR_opcode_field[0]),
    .ADR3(DLX_IDinst_IR_opcode_field[2]),
    .O(\CHOICE1757/FROM )
  );
  defparam DLX_IDinst_Ker706451.INIT = 16'h1100;
  X_LUT4 DLX_IDinst_Ker706451 (
    .ADR0(DLX_IDinst_IR_opcode_field[5]),
    .ADR1(DLX_IDinst_IR_opcode_field[1]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_IR_opcode_field[3]),
    .O(\CHOICE1757/GROM )
  );
  X_BUF \CHOICE1757/XUSED  (
    .I(\CHOICE1757/FROM ),
    .O(CHOICE1757)
  );
  X_BUF \CHOICE1757/YUSED  (
    .I(\CHOICE1757/GROM ),
    .O(DLX_IDinst_N70647)
  );
  defparam \DLX_IDinst_regA_eff<0>1 .INIT = 16'hA3A0;
  X_LUT4 \DLX_IDinst_regA_eff<0>1  (
    .ADR0(DLX_RF_data_in[0]),
    .ADR1(DLX_IDinst__n0002),
    .ADR2(DLX_IDinst__n0144),
    .ADR3(DLX_IDinst_reg_out_A_RF[0]),
    .O(\DLX_IDinst_regA_eff<0>/FROM )
  );
  defparam \DLX_IDinst__n0086<0>20 .INIT = 16'hF000;
  X_LUT4 \DLX_IDinst__n0086<0>20  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_N70295),
    .ADR3(DLX_IDinst_regA_eff[0]),
    .O(\DLX_IDinst_regA_eff<0>/GROM )
  );
  X_BUF \DLX_IDinst_regA_eff<0>/XUSED  (
    .I(\DLX_IDinst_regA_eff<0>/FROM ),
    .O(DLX_IDinst_regA_eff[0])
  );
  X_BUF \DLX_IDinst_regA_eff<0>/YUSED  (
    .I(\DLX_IDinst_regA_eff<0>/GROM ),
    .O(CHOICE2562)
  );
  defparam \DLX_IDinst_regA_eff<1>1 .INIT = 16'hD1C0;
  X_LUT4 \DLX_IDinst_regA_eff<1>1  (
    .ADR0(DLX_IDinst__n0002),
    .ADR1(DLX_IDinst__n0144),
    .ADR2(DLX_RF_data_in[1]),
    .ADR3(DLX_IDinst_reg_out_A_RF[1]),
    .O(\DLX_IDinst_regA_eff<1>/FROM )
  );
  defparam \DLX_IDinst__n0086<1>20 .INIT = 16'hAA00;
  X_LUT4 \DLX_IDinst__n0086<1>20  (
    .ADR0(DLX_IDinst_N70295),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_regA_eff[1]),
    .O(\DLX_IDinst_regA_eff<1>/GROM )
  );
  X_BUF \DLX_IDinst_regA_eff<1>/XUSED  (
    .I(\DLX_IDinst_regA_eff<1>/FROM ),
    .O(DLX_IDinst_regA_eff[1])
  );
  X_BUF \DLX_IDinst_regA_eff<1>/YUSED  (
    .I(\DLX_IDinst_regA_eff<1>/GROM ),
    .O(CHOICE2584)
  );
  defparam DLX_IDinst_Ker706711.INIT = 16'h0010;
  X_LUT4 DLX_IDinst_Ker706711 (
    .ADR0(DLX_IDinst_IR_latched[28]),
    .ADR1(DLX_IDinst_IR_latched[29]),
    .ADR2(DLX_IDinst_IR_latched[30]),
    .ADR3(DLX_IDinst_IR_latched[27]),
    .O(\DLX_IDinst_N70673/FROM )
  );
  defparam DLX_IDinst_Mmux__n0151_Result_SW0.INIT = 16'hC000;
  X_LUT4 DLX_IDinst_Mmux__n0151_Result_SW0 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_IR_latched[31]),
    .ADR2(DLX_IDinst_IR_latched[26]),
    .ADR3(DLX_IDinst_N70673),
    .O(\DLX_IDinst_N70673/GROM )
  );
  X_BUF \DLX_IDinst_N70673/XUSED  (
    .I(\DLX_IDinst_N70673/FROM ),
    .O(DLX_IDinst_N70673)
  );
  X_BUF \DLX_IDinst_N70673/YUSED  (
    .I(\DLX_IDinst_N70673/GROM ),
    .O(N95818)
  );
  defparam \DLX_IDinst__n0086<8>25 .INIT = 16'hCCCE;
  X_LUT4 \DLX_IDinst__n0086<8>25  (
    .ADR0(CHOICE2646),
    .ADR1(CHOICE2650),
    .ADR2(DLX_IDinst__n0364),
    .ADR3(DLX_IDinst_N70918),
    .O(\DLX_IDinst_branch_address<8>/FROM )
  );
  defparam \DLX_IDinst__n0086<8>31 .INIT = 16'hFFA0;
  X_LUT4 \DLX_IDinst__n0086<8>31  (
    .ADR0(N100609),
    .ADR1(VCC),
    .ADR2(DLX_IDinst__n0128[8]),
    .ADR3(CHOICE2651),
    .O(N105598)
  );
  X_BUF \DLX_IDinst_branch_address<8>/XUSED  (
    .I(\DLX_IDinst_branch_address<8>/FROM ),
    .O(CHOICE2651)
  );
  defparam DLX_IDinst_Ker705681.INIT = 16'hFFFC;
  X_LUT4 DLX_IDinst_Ker705681 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_counter[1]),
    .ADR2(DLX_IDinst_intr_slot),
    .ADR3(DLX_IDinst_counter[0]),
    .O(\DLX_IDinst_N70570/FROM )
  );
  defparam DLX_IDinst__n03351.INIT = 16'h0002;
  X_LUT4 DLX_IDinst__n03351 (
    .ADR0(DLX_IDinst_stall),
    .ADR1(DLX_IDinst_delay_slot),
    .ADR2(FREEZE_IBUF),
    .ADR3(DLX_IDinst_N70570),
    .O(\DLX_IDinst_N70570/GROM )
  );
  X_BUF \DLX_IDinst_N70570/XUSED  (
    .I(\DLX_IDinst_N70570/FROM ),
    .O(DLX_IDinst_N70570)
  );
  X_BUF \DLX_IDinst_N70570/YUSED  (
    .I(\DLX_IDinst_N70570/GROM ),
    .O(DLX_IDinst__n0335)
  );
  defparam \DLX_EXinst__n0006<10>42 .INIT = 16'h8A80;
  X_LUT4 \DLX_EXinst__n0006<10>42  (
    .ADR0(DLX_EXinst_N66475),
    .ADR1(DLX_EXinst_N64550),
    .ADR2(DLX_IDinst_IR_function_field[2]),
    .ADR3(DLX_EXinst_N64814),
    .O(\CHOICE4498/FROM )
  );
  defparam \DLX_EXinst__n0006<10>71 .INIT = 16'hFFFA;
  X_LUT4 \DLX_EXinst__n0006<10>71  (
    .ADR0(CHOICE4505),
    .ADR1(VCC),
    .ADR2(CHOICE4504),
    .ADR3(CHOICE4498),
    .O(\CHOICE4498/GROM )
  );
  X_BUF \CHOICE4498/XUSED  (
    .I(\CHOICE4498/FROM ),
    .O(CHOICE4498)
  );
  X_BUF \CHOICE4498/YUSED  (
    .I(\CHOICE4498/GROM ),
    .O(CHOICE4507)
  );
  defparam \DLX_IDinst_regA_eff<2>1 .INIT = 16'hA0E4;
  X_LUT4 \DLX_IDinst_regA_eff<2>1  (
    .ADR0(DLX_IDinst__n0144),
    .ADR1(DLX_IDinst_reg_out_A_RF[2]),
    .ADR2(DLX_RF_data_in[2]),
    .ADR3(DLX_IDinst__n0002),
    .O(\DLX_IDinst_regA_eff<2>/FROM )
  );
  defparam \DLX_IDinst__n0086<2>20 .INIT = 16'hF000;
  X_LUT4 \DLX_IDinst__n0086<2>20  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_N70295),
    .ADR3(DLX_IDinst_regA_eff[2]),
    .O(\DLX_IDinst_regA_eff<2>/GROM )
  );
  X_BUF \DLX_IDinst_regA_eff<2>/XUSED  (
    .I(\DLX_IDinst_regA_eff<2>/FROM ),
    .O(DLX_IDinst_regA_eff[2])
  );
  X_BUF \DLX_IDinst_regA_eff<2>/YUSED  (
    .I(\DLX_IDinst_regA_eff<2>/GROM ),
    .O(CHOICE2573)
  );
  defparam \DLX_EXinst__n0006<14>67 .INIT = 16'hCE00;
  X_LUT4 \DLX_EXinst__n0006<14>67  (
    .ADR0(DLX_EXinst__n0080),
    .ADR1(DLX_EXinst__n0079),
    .ADR2(\DLX_IDinst_Imm[14] ),
    .ADR3(DLX_IDinst_reg_out_A[14]),
    .O(\CHOICE4248/FROM )
  );
  defparam \DLX_EXinst__n0006<11>21 .INIT = 16'hCC08;
  X_LUT4 \DLX_EXinst__n0006<11>21  (
    .ADR0(DLX_EXinst__n0080),
    .ADR1(DLX_IDinst_reg_out_A[11]),
    .ADR2(\DLX_IDinst_Imm[11] ),
    .ADR3(DLX_EXinst__n0079),
    .O(\CHOICE4248/GROM )
  );
  X_BUF \CHOICE4248/XUSED  (
    .I(\CHOICE4248/FROM ),
    .O(CHOICE4248)
  );
  X_BUF \CHOICE4248/YUSED  (
    .I(\CHOICE4248/GROM ),
    .O(CHOICE3922)
  );
  defparam \DLX_IDinst_regA_eff<3>1 .INIT = 16'hAA0C;
  X_LUT4 \DLX_IDinst_regA_eff<3>1  (
    .ADR0(DLX_RF_data_in[3]),
    .ADR1(DLX_IDinst_reg_out_A_RF[3]),
    .ADR2(DLX_IDinst__n0002),
    .ADR3(DLX_IDinst__n0144),
    .O(\DLX_IDinst_regA_eff<3>/FROM )
  );
  defparam DLX_IDinst__n014612.INIT = 16'h0001;
  X_LUT4 DLX_IDinst__n014612 (
    .ADR0(DLX_IDinst_regA_eff[0]),
    .ADR1(DLX_IDinst_regA_eff[2]),
    .ADR2(DLX_IDinst_regA_eff[1]),
    .ADR3(DLX_IDinst_regA_eff[3]),
    .O(\DLX_IDinst_regA_eff<3>/GROM )
  );
  X_BUF \DLX_IDinst_regA_eff<3>/XUSED  (
    .I(\DLX_IDinst_regA_eff<3>/FROM ),
    .O(DLX_IDinst_regA_eff[3])
  );
  X_BUF \DLX_IDinst_regA_eff<3>/YUSED  (
    .I(\DLX_IDinst_regA_eff<3>/GROM ),
    .O(CHOICE3620)
  );
  defparam \DLX_IDinst__n0086<9>25 .INIT = 16'hCDCC;
  X_LUT4 \DLX_IDinst__n0086<9>25  (
    .ADR0(DLX_IDinst_N70918),
    .ADR1(CHOICE2661),
    .ADR2(DLX_IDinst__n0364),
    .ADR3(CHOICE2657),
    .O(\DLX_IDinst_branch_address<9>/FROM )
  );
  defparam \DLX_IDinst__n0086<9>31 .INIT = 16'hFFA0;
  X_LUT4 \DLX_IDinst__n0086<9>31  (
    .ADR0(DLX_IDinst__n0128[9]),
    .ADR1(VCC),
    .ADR2(N100609),
    .ADR3(CHOICE2662),
    .O(N105661)
  );
  X_BUF \DLX_IDinst_branch_address<9>/XUSED  (
    .I(\DLX_IDinst_branch_address<9>/FROM ),
    .O(CHOICE2662)
  );
  defparam DLX_IDinst_Ker709161.INIT = 16'h2000;
  X_LUT4 DLX_IDinst_Ker709161 (
    .ADR0(DLX_IDinst_N70909),
    .ADR1(DLX_IDinst_IR_latched[28]),
    .ADR2(DLX_IDinst_IR_latched[26]),
    .ADR3(DLX_IDinst_IR_latched[27]),
    .O(\DLX_IDinst_rd_addr<0>/FROM )
  );
  defparam \DLX_IDinst__n0107<0>1 .INIT = 16'h0F0A;
  X_LUT4 \DLX_IDinst__n0107<0>1  (
    .ADR0(DLX_IDinst_N70918),
    .ADR1(VCC),
    .ADR2(DLX_IDinst__n0331),
    .ADR3(DLX_IDinst__n0023[0]),
    .O(DLX_IDinst__n0107[0])
  );
  X_BUF \DLX_IDinst_rd_addr<0>/XUSED  (
    .I(\DLX_IDinst_rd_addr<0>/FROM ),
    .O(DLX_IDinst_N70918)
  );
  defparam \DLX_EXinst__n0006<11>42 .INIT = 16'hC088;
  X_LUT4 \DLX_EXinst__n0006<11>42  (
    .ADR0(DLX_EXinst_N65100),
    .ADR1(DLX_EXinst_N66475),
    .ADR2(N97305),
    .ADR3(DLX_IDinst_IR_function_field[2]),
    .O(\CHOICE3928/FROM )
  );
  defparam \DLX_EXinst__n0006<11>71 .INIT = 16'hFFFC;
  X_LUT4 \DLX_EXinst__n0006<11>71  (
    .ADR0(VCC),
    .ADR1(CHOICE3934),
    .ADR2(CHOICE3935),
    .ADR3(CHOICE3928),
    .O(\CHOICE3928/GROM )
  );
  X_BUF \CHOICE3928/XUSED  (
    .I(\CHOICE3928/FROM ),
    .O(CHOICE3928)
  );
  X_BUF \CHOICE3928/YUSED  (
    .I(\CHOICE3928/GROM ),
    .O(CHOICE3937)
  );
  defparam \DLX_IDinst_regA_eff<4>1 .INIT = 16'h88D8;
  X_LUT4 \DLX_IDinst_regA_eff<4>1  (
    .ADR0(DLX_IDinst__n0144),
    .ADR1(DLX_RF_data_in[4]),
    .ADR2(DLX_IDinst_reg_out_A_RF[4]),
    .ADR3(DLX_IDinst__n0002),
    .O(\DLX_IDinst_regA_eff<4>/FROM )
  );
  defparam \DLX_IDinst__n0086<4>20 .INIT = 16'hAA00;
  X_LUT4 \DLX_IDinst__n0086<4>20  (
    .ADR0(DLX_IDinst_N70295),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_regA_eff[4]),
    .O(\DLX_IDinst_regA_eff<4>/GROM )
  );
  X_BUF \DLX_IDinst_regA_eff<4>/XUSED  (
    .I(\DLX_IDinst_regA_eff<4>/FROM ),
    .O(DLX_IDinst_regA_eff[4])
  );
  X_BUF \DLX_IDinst_regA_eff<4>/YUSED  (
    .I(\DLX_IDinst_regA_eff<4>/GROM ),
    .O(CHOICE2606)
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<127>1 .INIT = 16'h0100;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<127>1  (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(DLX_IDinst_reg_out_B[0]),
    .ADR2(DLX_EXinst_N62740),
    .ADR3(DLX_IDinst_reg_out_A[31]),
    .O(\DLX_EXinst_Mshift__n0023_Sh<127>/FROM )
  );
  defparam \DLX_EXinst__n0006<15>172 .INIT = 16'hA820;
  X_LUT4 \DLX_EXinst__n0006<15>172  (
    .ADR0(DLX_EXinst_N66177),
    .ADR1(DLX_IDinst_reg_out_B[5]),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(\DLX_EXinst_Mshift__n0023_Sh[127] ),
    .O(\DLX_EXinst_Mshift__n0023_Sh<127>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0023_Sh<127>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0023_Sh<127>/FROM ),
    .O(\DLX_EXinst_Mshift__n0023_Sh[127] )
  );
  X_BUF \DLX_EXinst_Mshift__n0023_Sh<127>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0023_Sh<127>/GROM ),
    .O(CHOICE4849)
  );
  defparam \DLX_EXinst__n0006<3>120 .INIT = 16'h8000;
  X_LUT4 \DLX_EXinst__n0006<3>120  (
    .ADR0(CHOICE3377),
    .ADR1(CHOICE3408),
    .ADR2(DLX_IDinst_IR_function_field[4]),
    .ADR3(N101537),
    .O(\CHOICE5047/FROM )
  );
  defparam \DLX_EXinst__n0006<11>62 .INIT = 16'h8000;
  X_LUT4 \DLX_EXinst__n0006<11>62  (
    .ADR0(DLX_IDinst_IR_function_field[4]),
    .ADR1(CHOICE3377),
    .ADR2(N101253),
    .ADR3(CHOICE3408),
    .O(\CHOICE5047/GROM )
  );
  X_BUF \CHOICE5047/XUSED  (
    .I(\CHOICE5047/FROM ),
    .O(CHOICE5047)
  );
  X_BUF \CHOICE5047/YUSED  (
    .I(\CHOICE5047/GROM ),
    .O(CHOICE3935)
  );
  defparam \DLX_EXinst__n0006<21>85 .INIT = 16'h8200;
  X_LUT4 \DLX_EXinst__n0006<21>85  (
    .ADR0(\DLX_IDinst_Imm[31] ),
    .ADR1(DLX_IDinst_IR_opcode_field[1]),
    .ADR2(N127370),
    .ADR3(DLX_EXinst_N66105),
    .O(\CHOICE4185/FROM )
  );
  defparam \DLX_EXinst__n0006<12>15 .INIT = 16'h8020;
  X_LUT4 \DLX_EXinst__n0006<12>15  (
    .ADR0(\DLX_IDinst_Imm[12] ),
    .ADR1(N127366),
    .ADR2(DLX_EXinst_N66105),
    .ADR3(DLX_IDinst_IR_opcode_field[1]),
    .O(\CHOICE4185/GROM )
  );
  X_BUF \CHOICE4185/XUSED  (
    .I(\CHOICE4185/FROM ),
    .O(CHOICE4185)
  );
  X_BUF \CHOICE4185/YUSED  (
    .I(\CHOICE4185/GROM ),
    .O(CHOICE3861)
  );
  defparam \DLX_IDinst_regA_eff<5>1 .INIT = 16'hA0E4;
  X_LUT4 \DLX_IDinst_regA_eff<5>1  (
    .ADR0(DLX_IDinst__n0144),
    .ADR1(DLX_IDinst_reg_out_A_RF[5]),
    .ADR2(DLX_RF_data_in[5]),
    .ADR3(DLX_IDinst__n0002),
    .O(\DLX_IDinst_regA_eff<5>/FROM )
  );
  defparam \DLX_IDinst__n0086<5>20 .INIT = 16'hF000;
  X_LUT4 \DLX_IDinst__n0086<5>20  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_N70295),
    .ADR3(DLX_IDinst_regA_eff[5]),
    .O(\DLX_IDinst_regA_eff<5>/GROM )
  );
  X_BUF \DLX_IDinst_regA_eff<5>/XUSED  (
    .I(\DLX_IDinst_regA_eff<5>/FROM ),
    .O(DLX_IDinst_regA_eff[5])
  );
  X_BUF \DLX_IDinst_regA_eff<5>/YUSED  (
    .I(\DLX_IDinst_regA_eff<5>/GROM ),
    .O(CHOICE2617)
  );
  defparam DLX_EXinst_Ker66150_SW0.INIT = 16'hAFAC;
  X_LUT4 DLX_EXinst_Ker66150_SW0 (
    .ADR0(\DLX_EXinst_Mshift__n0027_Sh[0] ),
    .ADR1(CHOICE1006),
    .ADR2(DLX_IDinst_IR_function_field_2_1),
    .ADR3(CHOICE1012),
    .O(\N90656/FROM )
  );
  defparam DLX_EXinst_Ker66150.INIT = 16'h0200;
  X_LUT4 DLX_EXinst_Ker66150 (
    .ADR0(DLX_EXinst__n0081),
    .ADR1(DLX_IDinst_IR_function_field_3_1),
    .ADR2(N109130),
    .ADR3(N90656),
    .O(\N90656/GROM )
  );
  X_BUF \N90656/XUSED  (
    .I(\N90656/FROM ),
    .O(N90656)
  );
  X_BUF \N90656/YUSED  (
    .I(\N90656/GROM ),
    .O(DLX_EXinst_N66152)
  );
  defparam DLX_IDinst_Ker70640122.INIT = 16'h0015;
  X_LUT4 DLX_IDinst_Ker70640122 (
    .ADR0(N126506),
    .ADR1(DLX_IDinst_IR_latched[30]),
    .ADR2(DLX_IDinst_N70918),
    .ADR3(DLX_IDinst__n0071),
    .O(\N109741/FROM )
  );
  defparam \DLX_IDinst_slot_num_FFd3-In15 .INIT = 16'hE0C0;
  X_LUT4 \DLX_IDinst_slot_num_FFd3-In15  (
    .ADR0(DLX_IDinst_N70333),
    .ADR1(FREEZE_IBUF),
    .ADR2(N126589),
    .ADR3(N109741),
    .O(\N109741/GROM )
  );
  X_BUF \N109741/XUSED  (
    .I(\N109741/FROM ),
    .O(N109741)
  );
  X_BUF \N109741/YUSED  (
    .I(\N109741/GROM ),
    .O(CHOICE2508)
  );
  defparam DLX_IDinst_Ker707841.INIT = 16'hF080;
  X_LUT4 DLX_IDinst_Ker707841 (
    .ADR0(DLX_IDinst_N70610),
    .ADR1(DLX_IDinst_N70924),
    .ADR2(DLX_IDinst_N69568),
    .ADR3(DLX_IDinst_N69963),
    .O(\DLX_IDinst_N70786/FROM )
  );
  defparam \DLX_IDinst__n0086<10>6 .INIT = 16'hEAC0;
  X_LUT4 \DLX_IDinst__n0086<10>6  (
    .ADR0(DLX_IDinst_branch_address[10]),
    .ADR1(DLX_IDinst__n0071),
    .ADR2(DLX_IDinst_EPC[10]),
    .ADR3(DLX_IDinst_N70786),
    .O(\DLX_IDinst_N70786/GROM )
  );
  X_BUF \DLX_IDinst_N70786/XUSED  (
    .I(\DLX_IDinst_N70786/FROM ),
    .O(DLX_IDinst_N70786)
  );
  X_BUF \DLX_IDinst_N70786/YUSED  (
    .I(\DLX_IDinst_N70786/GROM ),
    .O(CHOICE2668)
  );
  defparam DLX_IDinst_Ker6995596.INIT = 16'h0001;
  X_LUT4 DLX_IDinst_Ker6995596 (
    .ADR0(DLX_IDinst_IR_opcode_field[2]),
    .ADR1(DLX_IDinst_IR_opcode_field[0]),
    .ADR2(DLX_IDinst_IR_opcode_field[4]),
    .ADR3(DLX_IDinst_IR_opcode_field[1]),
    .O(\CHOICE1444/FROM )
  );
  defparam \DLX_EXinst__n0006<20>18 .INIT = 16'h0080;
  X_LUT4 \DLX_EXinst__n0006<20>18  (
    .ADR0(DLX_IDinst_IR_opcode_field[1]),
    .ADR1(DLX_EXinst_N66112),
    .ADR2(\DLX_EXinst_Mshift__n0028_Sh[52] ),
    .ADR3(DLX_IDinst_IR_opcode_field[0]),
    .O(\CHOICE1444/GROM )
  );
  X_BUF \CHOICE1444/XUSED  (
    .I(\CHOICE1444/FROM ),
    .O(CHOICE1444)
  );
  X_BUF \CHOICE1444/YUSED  (
    .I(\CHOICE1444/GROM ),
    .O(CHOICE4879)
  );
  defparam \DLX_EXinst__n0006<14>18 .INIT = 16'hC0C0;
  X_LUT4 \DLX_EXinst__n0006<14>18  (
    .ADR0(VCC),
    .ADR1(N102270),
    .ADR2(DLX_IDinst_IR_function_field[4]),
    .ADR3(VCC),
    .O(\CHOICE4234/FROM )
  );
  defparam \DLX_EXinst__n0006<12>18 .INIT = 16'hFA00;
  X_LUT4 \DLX_EXinst__n0006<12>18  (
    .ADR0(CHOICE2085),
    .ADR1(VCC),
    .ADR2(CHOICE2081),
    .ADR3(DLX_IDinst_IR_function_field[4]),
    .O(\CHOICE4234/GROM )
  );
  X_BUF \CHOICE4234/XUSED  (
    .I(\CHOICE4234/FROM ),
    .O(CHOICE4234)
  );
  X_BUF \CHOICE4234/YUSED  (
    .I(\CHOICE4234/GROM ),
    .O(CHOICE3862)
  );
  defparam \DLX_EXinst__n0006<21>272_SW0 .INIT = 16'hFAF0;
  X_LUT4 \DLX_EXinst__n0006<21>272_SW0  (
    .ADR0(DLX_EXinst_N66226),
    .ADR1(VCC),
    .ADR2(CHOICE4220),
    .ADR3(CHOICE4206),
    .O(\N126419/FROM )
  );
  defparam \DLX_EXinst__n0006<21>272 .INIT = 16'hF0E0;
  X_LUT4 \DLX_EXinst__n0006<21>272  (
    .ADR0(CHOICE4196),
    .ADR1(CHOICE4211),
    .ADR2(DLX_EXinst__n0030),
    .ADR3(N126419),
    .O(\N126419/GROM )
  );
  X_BUF \N126419/XUSED  (
    .I(\N126419/FROM ),
    .O(N126419)
  );
  X_BUF \N126419/YUSED  (
    .I(\N126419/GROM ),
    .O(CHOICE4223)
  );
  defparam \DLX_EXinst__n0006<27>36 .INIT = 16'h8008;
  X_LUT4 \DLX_EXinst__n0006<27>36  (
    .ADR0(DLX_EXinst_N66105),
    .ADR1(\DLX_IDinst_Imm[31] ),
    .ADR2(DLX_IDinst_IR_opcode_field[1]),
    .ADR3(N127362),
    .O(\CHOICE4621/FROM )
  );
  defparam \DLX_EXinst__n0006<11>59 .INIT = 16'h8008;
  X_LUT4 \DLX_EXinst__n0006<11>59  (
    .ADR0(DLX_EXinst_N66105),
    .ADR1(\DLX_IDinst_Imm[11] ),
    .ADR2(DLX_IDinst_IR_opcode_field[1]),
    .ADR3(N127334),
    .O(\CHOICE4621/GROM )
  );
  X_BUF \CHOICE4621/XUSED  (
    .I(\CHOICE4621/FROM ),
    .O(CHOICE4621)
  );
  X_BUF \CHOICE4621/YUSED  (
    .I(\CHOICE4621/GROM ),
    .O(CHOICE3934)
  );
  defparam \DLX_IDinst_regA_eff<6>1 .INIT = 16'hC0E2;
  X_LUT4 \DLX_IDinst_regA_eff<6>1  (
    .ADR0(DLX_IDinst_reg_out_A_RF[6]),
    .ADR1(DLX_IDinst__n0144),
    .ADR2(DLX_RF_data_in[6]),
    .ADR3(DLX_IDinst__n0002),
    .O(\DLX_IDinst_regA_eff<6>/FROM )
  );
  defparam \DLX_IDinst__n0086<6>20 .INIT = 16'hAA00;
  X_LUT4 \DLX_IDinst__n0086<6>20  (
    .ADR0(DLX_IDinst_N70295),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_regA_eff[6]),
    .O(\DLX_IDinst_regA_eff<6>/GROM )
  );
  X_BUF \DLX_IDinst_regA_eff<6>/XUSED  (
    .I(\DLX_IDinst_regA_eff<6>/FROM ),
    .O(DLX_IDinst_regA_eff[6])
  );
  X_BUF \DLX_IDinst_regA_eff<6>/YUSED  (
    .I(\DLX_IDinst_regA_eff<6>/GROM ),
    .O(CHOICE2639)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_inv_11.INIT = 16'h50F5;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_inv_11 (
    .ADR0(DLX_EXinst_Mcompar__n0063_inst_cy_260),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[31]),
    .ADR3(DLX_IDinst_reg_out_A[31]),
    .O(\DLX_EXinst__n0063/FROM )
  );
  defparam \DLX_EXinst__n0006<0>220 .INIT = 16'hA820;
  X_LUT4 \DLX_EXinst__n0006<0>220  (
    .ADR0(DLX_IDinst_IR_function_field[0]),
    .ADR1(DLX_IDinst_IR_function_field[2]),
    .ADR2(DLX_EXinst__n0055),
    .ADR3(DLX_EXinst__n0063),
    .O(\DLX_EXinst__n0063/GROM )
  );
  X_BUF \DLX_EXinst__n0063/XUSED  (
    .I(\DLX_EXinst__n0063/FROM ),
    .O(DLX_EXinst__n0063)
  );
  X_BUF \DLX_EXinst__n0063/YUSED  (
    .I(\DLX_EXinst__n0063/GROM ),
    .O(CHOICE5899)
  );
  defparam \DLX_EXinst__n0006<4>228_SW0 .INIT = 16'hFACC;
  X_LUT4 \DLX_EXinst__n0006<4>228_SW0  (
    .ADR0(CHOICE4000),
    .ADR1(CHOICE4018),
    .ADR2(CHOICE4004),
    .ADR3(DLX_IDinst_reg_out_B[4]),
    .O(\N126239/FROM )
  );
  defparam \DLX_EXinst__n0006<4>228 .INIT = 16'hFFF8;
  X_LUT4 \DLX_EXinst__n0006<4>228  (
    .ADR0(N101725),
    .ADR1(DLX_EXinst_ALU_result[4]),
    .ADR2(CHOICE4021),
    .ADR3(N126239),
    .O(\N126239/GROM )
  );
  X_BUF \N126239/XUSED  (
    .I(\N126239/FROM ),
    .O(N126239)
  );
  X_BUF \N126239/YUSED  (
    .I(\N126239/GROM ),
    .O(CHOICE4023)
  );
  defparam \DLX_EXinst__n0006<27>10 .INIT = 16'h4000;
  X_LUT4 \DLX_EXinst__n0006<27>10  (
    .ADR0(N109130),
    .ADR1(DLX_EXinst__n0081),
    .ADR2(DLX_IDinst_IR_function_field[4]),
    .ADR3(\DLX_EXinst_Mshift__n0027_Sh[43] ),
    .O(\CHOICE4611/FROM )
  );
  defparam \DLX_EXinst__n0006<20>38 .INIT = 16'hDDDC;
  X_LUT4 \DLX_EXinst__n0006<20>38  (
    .ADR0(N109130),
    .ADR1(N97892),
    .ADR2(CHOICE4879),
    .ADR3(CHOICE4878),
    .O(\CHOICE4611/GROM )
  );
  X_BUF \CHOICE4611/XUSED  (
    .I(\CHOICE4611/FROM ),
    .O(CHOICE4611)
  );
  X_BUF \CHOICE4611/YUSED  (
    .I(\CHOICE4611/GROM ),
    .O(CHOICE4882)
  );
  defparam \DLX_EXinst__n0006<18>42_SW0 .INIT = 16'h0033;
  X_LUT4 \DLX_EXinst__n0006<18>42_SW0  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_IR_opcode_field[0]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[18]),
    .O(\N127354/FROM )
  );
  defparam \DLX_EXinst__n0006<23>85_SW0 .INIT = 16'h0303;
  X_LUT4 \DLX_EXinst__n0006<23>85_SW0  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_IR_opcode_field[0]),
    .ADR2(DLX_IDinst_reg_out_A[23]),
    .ADR3(VCC),
    .O(\N127354/GROM )
  );
  X_BUF \N127354/XUSED  (
    .I(\N127354/FROM ),
    .O(N127354)
  );
  X_BUF \N127354/YUSED  (
    .I(\N127354/GROM ),
    .O(N127400)
  );
  defparam \DLX_EXinst__n0006<12>71 .INIT = 16'hFF54;
  X_LUT4 \DLX_EXinst__n0006<12>71  (
    .ADR0(DLX_IDinst_IR_function_field[4]),
    .ADR1(CHOICE3870),
    .ADR2(CHOICE3869),
    .ADR3(CHOICE3876),
    .O(\CHOICE3877/FROM )
  );
  defparam \DLX_EXinst__n0006<12>98 .INIT = 16'h0F0E;
  X_LUT4 \DLX_EXinst__n0006<12>98  (
    .ADR0(CHOICE3861),
    .ADR1(CHOICE3862),
    .ADR2(DLX_EXinst__n0030),
    .ADR3(CHOICE3877),
    .O(\CHOICE3877/GROM )
  );
  X_BUF \CHOICE3877/XUSED  (
    .I(\CHOICE3877/FROM ),
    .O(CHOICE3877)
  );
  X_BUF \CHOICE3877/YUSED  (
    .I(\CHOICE3877/GROM ),
    .O(CHOICE3879)
  );
  defparam \DLX_EXinst__n0006<26>10 .INIT = 16'h4000;
  X_LUT4 \DLX_EXinst__n0006<26>10  (
    .ADR0(N109130),
    .ADR1(DLX_EXinst__n0081),
    .ADR2(DLX_IDinst_IR_function_field[4]),
    .ADR3(\DLX_EXinst_Mshift__n0027_Sh[42] ),
    .O(\CHOICE4676/FROM )
  );
  defparam \DLX_EXinst__n0006<11>87 .INIT = 16'hFFBA;
  X_LUT4 \DLX_EXinst__n0006<11>87  (
    .ADR0(CHOICE3922),
    .ADR1(N109130),
    .ADR2(CHOICE3917),
    .ADR3(CHOICE3937),
    .O(\CHOICE4676/GROM )
  );
  X_BUF \CHOICE4676/XUSED  (
    .I(\CHOICE4676/FROM ),
    .O(CHOICE4676)
  );
  X_BUF \CHOICE4676/YUSED  (
    .I(\CHOICE4676/GROM ),
    .O(CHOICE3938)
  );
  defparam \DLX_EXinst__n0006<24>76 .INIT = 16'h9000;
  X_LUT4 \DLX_EXinst__n0006<24>76  (
    .ADR0(DLX_IDinst_IR_opcode_field[1]),
    .ADR1(N127358),
    .ADR2(DLX_EXinst_N66105),
    .ADR3(\DLX_IDinst_Imm[31] ),
    .O(\CHOICE3755/FROM )
  );
  defparam \DLX_EXinst__n0006<13>15 .INIT = 16'h9000;
  X_LUT4 \DLX_EXinst__n0006<13>15  (
    .ADR0(N127326),
    .ADR1(DLX_IDinst_IR_opcode_field[1]),
    .ADR2(DLX_EXinst_N66105),
    .ADR3(\DLX_IDinst_Imm[13] ),
    .O(\CHOICE3755/GROM )
  );
  X_BUF \CHOICE3755/XUSED  (
    .I(\CHOICE3755/FROM ),
    .O(CHOICE3755)
  );
  X_BUF \CHOICE3755/YUSED  (
    .I(\CHOICE3755/GROM ),
    .O(CHOICE4293)
  );
  defparam \DLX_IDinst_regA_eff<7>1 .INIT = 16'h88D8;
  X_LUT4 \DLX_IDinst_regA_eff<7>1  (
    .ADR0(DLX_IDinst__n0144),
    .ADR1(DLX_RF_data_in[7]),
    .ADR2(DLX_IDinst_reg_out_A_RF[7]),
    .ADR3(DLX_IDinst__n0002),
    .O(\DLX_IDinst_regA_eff<7>/FROM )
  );
  defparam DLX_IDinst__n014625.INIT = 16'h0001;
  X_LUT4 DLX_IDinst__n014625 (
    .ADR0(DLX_IDinst_regA_eff[5]),
    .ADR1(DLX_IDinst_regA_eff[4]),
    .ADR2(DLX_IDinst_regA_eff[6]),
    .ADR3(DLX_IDinst_regA_eff[7]),
    .O(\DLX_IDinst_regA_eff<7>/GROM )
  );
  X_BUF \DLX_IDinst_regA_eff<7>/XUSED  (
    .I(\DLX_IDinst_regA_eff<7>/FROM ),
    .O(DLX_IDinst_regA_eff[7])
  );
  X_BUF \DLX_IDinst_regA_eff<7>/YUSED  (
    .I(\DLX_IDinst_regA_eff<7>/GROM ),
    .O(CHOICE3627)
  );
  defparam DLX_IDinst__n0122130_SW0.INIT = 16'hCFCE;
  X_LUT4 DLX_IDinst__n0122130_SW0 (
    .ADR0(CHOICE3297),
    .ADR1(CHOICE3317),
    .ADR2(DLX_IDinst__n0364),
    .ADR3(CHOICE3311),
    .O(\DLX_IDinst_delay_slot/FROM )
  );
  defparam DLX_IDinst__n0122130.INIT = 16'h0800;
  X_LUT4 DLX_IDinst__n0122130 (
    .ADR0(N95693),
    .ADR1(N127182),
    .ADR2(DLX_IDinst_intr_slot),
    .ADR3(DLX_EXinst__n0149),
    .O(N109531)
  );
  X_BUF \DLX_IDinst_delay_slot/XUSED  (
    .I(\DLX_IDinst_delay_slot/FROM ),
    .O(N127182)
  );
  defparam \DLX_EXinst__n0006<14>41 .INIT = 16'h8A80;
  X_LUT4 \DLX_EXinst__n0006<14>41  (
    .ADR0(DLX_EXinst_N66202),
    .ADR1(DLX_EXinst_N62826),
    .ADR2(DLX_IDinst_IR_function_field[3]),
    .ADR3(N93331),
    .O(\CHOICE4242/FROM )
  );
  defparam \DLX_EXinst__n0006<13>41 .INIT = 16'hA280;
  X_LUT4 \DLX_EXinst__n0006<13>41  (
    .ADR0(DLX_EXinst_N66202),
    .ADR1(DLX_IDinst_IR_function_field[3]),
    .ADR2(DLX_EXinst_N62821),
    .ADR3(N93279),
    .O(\CHOICE4242/GROM )
  );
  X_BUF \CHOICE4242/XUSED  (
    .I(\CHOICE4242/FROM ),
    .O(CHOICE4242)
  );
  X_BUF \CHOICE4242/YUSED  (
    .I(\CHOICE4242/GROM ),
    .O(CHOICE4302)
  );
  defparam vga_top_vga1_Ker73382_SW0.INIT = 16'hFFBF;
  X_LUT4 vga_top_vga1_Ker73382_SW0 (
    .ADR0(vga_top_vga1_hcounter[8]),
    .ADR1(vga_top_vga1_hcounter[3]),
    .ADR2(vga_top_vga1_hcounter[0]),
    .ADR3(vga_top_vga1_hcounter[9]),
    .O(\N100282/FROM )
  );
  defparam vga_top_vga1_Ker73382.INIT = 16'h0040;
  X_LUT4 vga_top_vga1_Ker73382 (
    .ADR0(vga_top_vga1_vcounter[0]),
    .ADR1(vga_top_vga1_N73389),
    .ADR2(vga_top_vga1_vcounter[1]),
    .ADR3(N100282),
    .O(\N100282/GROM )
  );
  X_BUF \N100282/XUSED  (
    .I(\N100282/FROM ),
    .O(N100282)
  );
  X_BUF \N100282/YUSED  (
    .I(\N100282/GROM ),
    .O(vga_top_vga1_N73384)
  );
  defparam \DLX_EXinst__n0006<25>10 .INIT = 16'h0800;
  X_LUT4 \DLX_EXinst__n0006<25>10  (
    .ADR0(DLX_EXinst__n0081),
    .ADR1(DLX_IDinst_IR_function_field[4]),
    .ADR2(N109130),
    .ADR3(\DLX_EXinst_Mshift__n0027_Sh[41] ),
    .O(\CHOICE4741/FROM )
  );
  defparam \DLX_EXinst__n0006<13>18 .INIT = 16'hCC00;
  X_LUT4 \DLX_EXinst__n0006<13>18  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_IR_function_field[4]),
    .ADR2(VCC),
    .ADR3(N102162),
    .O(\CHOICE4741/GROM )
  );
  X_BUF \CHOICE4741/XUSED  (
    .I(\CHOICE4741/FROM ),
    .O(CHOICE4741)
  );
  X_BUF \CHOICE4741/YUSED  (
    .I(\CHOICE4741/GROM ),
    .O(CHOICE4294)
  );
  defparam \DLX_EXinst__n0006<20>59 .INIT = 16'hFCAA;
  X_LUT4 \DLX_EXinst__n0006<20>59  (
    .ADR0(CHOICE4882),
    .ADR1(DLX_EXinst_N66152),
    .ADR2(DLX_EXinst__n0077),
    .ADR3(DLX_IDinst_IR_function_field[4]),
    .O(\CHOICE4884/FROM )
  );
  defparam \DLX_EXinst__n0006<20>336_SW0 .INIT = 16'h0F0C;
  X_LUT4 \DLX_EXinst__n0006<20>336_SW0  (
    .ADR0(VCC),
    .ADR1(CHOICE4897),
    .ADR2(DLX_EXinst__n0030),
    .ADR3(CHOICE4884),
    .O(\CHOICE4884/GROM )
  );
  X_BUF \CHOICE4884/XUSED  (
    .I(\CHOICE4884/FROM ),
    .O(CHOICE4884)
  );
  X_BUF \CHOICE4884/YUSED  (
    .I(\CHOICE4884/GROM ),
    .O(N127200)
  );
  defparam \DLX_IDinst_regA_eff<8>1 .INIT = 16'hC5C0;
  X_LUT4 \DLX_IDinst_regA_eff<8>1  (
    .ADR0(DLX_IDinst__n0002),
    .ADR1(DLX_MEMinst_RF_data_in[8]),
    .ADR2(DLX_IDinst__n0144),
    .ADR3(DLX_IDinst_reg_out_A_RF[8]),
    .O(\DLX_IDinst_regA_eff<8>/FROM )
  );
  defparam \DLX_IDinst__n0086<8>20 .INIT = 16'hAA00;
  X_LUT4 \DLX_IDinst__n0086<8>20  (
    .ADR0(DLX_IDinst_N70295),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_regA_eff[8]),
    .O(\DLX_IDinst_regA_eff<8>/GROM )
  );
  X_BUF \DLX_IDinst_regA_eff<8>/XUSED  (
    .I(\DLX_IDinst_regA_eff<8>/FROM ),
    .O(DLX_IDinst_regA_eff[8])
  );
  X_BUF \DLX_IDinst_regA_eff<8>/YUSED  (
    .I(\DLX_IDinst_regA_eff<8>/GROM ),
    .O(CHOICE2650)
  );
  defparam \DLX_EXinst__n0006<21>28 .INIT = 16'h0B08;
  X_LUT4 \DLX_EXinst__n0006<21>28  (
    .ADR0(DLX_EXinst_N64062),
    .ADR1(DLX_IDinst_IR_function_field[2]),
    .ADR2(DLX_IDinst_IR_function_field[4]),
    .ADR3(DLX_EXinst_N64304),
    .O(\CHOICE4173/FROM )
  );
  defparam \DLX_EXinst__n0006<21>41 .INIT = 16'h0C04;
  X_LUT4 \DLX_EXinst__n0006<21>41  (
    .ADR0(N127126),
    .ADR1(DLX_EXinst__n0081),
    .ADR2(N109130),
    .ADR3(CHOICE4173),
    .O(\CHOICE4173/GROM )
  );
  X_BUF \CHOICE4173/XUSED  (
    .I(\CHOICE4173/FROM ),
    .O(CHOICE4173)
  );
  X_BUF \CHOICE4173/YUSED  (
    .I(\CHOICE4173/GROM ),
    .O(CHOICE4175)
  );
  defparam \DLX_EXinst__n0006<14>38 .INIT = 16'hC480;
  X_LUT4 \DLX_EXinst__n0006<14>38  (
    .ADR0(DLX_IDinst_IR_function_field[2]),
    .ADR1(DLX_EXinst_N63185),
    .ADR2(DLX_EXinst_N64859),
    .ADR3(DLX_EXinst_N64550),
    .O(\CHOICE4241/FROM )
  );
  defparam \DLX_EXinst__n0006<13>38 .INIT = 16'hC840;
  X_LUT4 \DLX_EXinst__n0006<13>38  (
    .ADR0(DLX_IDinst_IR_function_field[2]),
    .ADR1(DLX_EXinst_N63185),
    .ADR2(DLX_EXinst_N64560),
    .ADR3(DLX_EXinst_N64854),
    .O(\CHOICE4241/GROM )
  );
  X_BUF \CHOICE4241/XUSED  (
    .I(\CHOICE4241/FROM ),
    .O(CHOICE4241)
  );
  X_BUF \CHOICE4241/YUSED  (
    .I(\CHOICE4241/GROM ),
    .O(CHOICE4301)
  );
  defparam \DLX_EXinst__n0006<18>42 .INIT = 16'h8008;
  X_LUT4 \DLX_EXinst__n0006<18>42  (
    .ADR0(\DLX_IDinst_Imm[31] ),
    .ADR1(DLX_EXinst_N66105),
    .ADR2(DLX_IDinst_IR_opcode_field[1]),
    .ADR3(N127354),
    .O(\CHOICE5421/FROM )
  );
  defparam \DLX_EXinst__n0006<14>15 .INIT = 16'h8008;
  X_LUT4 \DLX_EXinst__n0006<14>15  (
    .ADR0(DLX_EXinst_N66105),
    .ADR1(\DLX_IDinst_Imm[14] ),
    .ADR2(N127350),
    .ADR3(DLX_IDinst_IR_opcode_field[1]),
    .O(\CHOICE5421/GROM )
  );
  X_BUF \CHOICE5421/XUSED  (
    .I(\CHOICE5421/FROM ),
    .O(CHOICE5421)
  );
  X_BUF \CHOICE5421/YUSED  (
    .I(\CHOICE5421/GROM ),
    .O(CHOICE4233)
  );
  defparam \DLX_IDinst_regA_eff<9>1 .INIT = 16'hAE04;
  X_LUT4 \DLX_IDinst_regA_eff<9>1  (
    .ADR0(DLX_IDinst__n0144),
    .ADR1(DLX_IDinst_reg_out_A_RF[9]),
    .ADR2(DLX_IDinst__n0002),
    .ADR3(DLX_MEMinst_RF_data_in[9]),
    .O(\DLX_IDinst_regA_eff<9>/FROM )
  );
  defparam \DLX_IDinst__n0086<9>20 .INIT = 16'hF000;
  X_LUT4 \DLX_IDinst__n0086<9>20  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_N70295),
    .ADR3(DLX_IDinst_regA_eff[9]),
    .O(\DLX_IDinst_regA_eff<9>/GROM )
  );
  X_BUF \DLX_IDinst_regA_eff<9>/XUSED  (
    .I(\DLX_IDinst_regA_eff<9>/FROM ),
    .O(DLX_IDinst_regA_eff[9])
  );
  X_BUF \DLX_IDinst_regA_eff<9>/YUSED  (
    .I(\DLX_IDinst_regA_eff<9>/GROM ),
    .O(CHOICE2661)
  );
  defparam DLX_IDinst_Ker709831.INIT = 16'h0001;
  X_LUT4 DLX_IDinst_Ker709831 (
    .ADR0(DLX_IDinst__n0348),
    .ADR1(DLX_IDinst__n0345),
    .ADR2(DLX_IDinst__n0136),
    .ADR3(DLX_IDinst__n0135),
    .O(\DLX_IDinst_N70985/FROM )
  );
  defparam DLX_IDinst__n012249_SW0.INIT = 16'hEEFF;
  X_LUT4 DLX_IDinst__n012249_SW0 (
    .ADR0(DLX_IDinst_IR_latched[30]),
    .ADR1(DLX_IDinst_IR_latched[27]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_N70985),
    .O(\DLX_IDinst_N70985/GROM )
  );
  X_BUF \DLX_IDinst_N70985/XUSED  (
    .I(\DLX_IDinst_N70985/FROM ),
    .O(DLX_IDinst_N70985)
  );
  X_BUF \DLX_IDinst_N70985/YUSED  (
    .I(\DLX_IDinst_N70985/GROM ),
    .O(N126675)
  );
  defparam \DLX_EXinst__n0006<13>71 .INIT = 16'hAAFE;
  X_LUT4 \DLX_EXinst__n0006<13>71  (
    .ADR0(CHOICE4308),
    .ADR1(CHOICE4302),
    .ADR2(CHOICE4301),
    .ADR3(DLX_IDinst_IR_function_field[4]),
    .O(\CHOICE4309/FROM )
  );
  defparam \DLX_EXinst__n0006<13>98 .INIT = 16'h3332;
  X_LUT4 \DLX_EXinst__n0006<13>98  (
    .ADR0(CHOICE4293),
    .ADR1(DLX_EXinst__n0030),
    .ADR2(CHOICE4294),
    .ADR3(CHOICE4309),
    .O(\CHOICE4309/GROM )
  );
  X_BUF \CHOICE4309/XUSED  (
    .I(\CHOICE4309/FROM ),
    .O(CHOICE4309)
  );
  X_BUF \CHOICE4309/YUSED  (
    .I(\CHOICE4309/GROM ),
    .O(CHOICE4311)
  );
  defparam \DLX_EXinst__n0006<26>36 .INIT = 16'h9000;
  X_LUT4 \DLX_EXinst__n0006<26>36  (
    .ADR0(DLX_IDinst_IR_opcode_field[1]),
    .ADR1(N127342),
    .ADR2(DLX_EXinst_N66105),
    .ADR3(\DLX_IDinst_Imm[31] ),
    .O(\CHOICE4686/FROM )
  );
  defparam \DLX_EXinst__n0006<20>96 .INIT = 16'h9000;
  X_LUT4 \DLX_EXinst__n0006<20>96  (
    .ADR0(N127338),
    .ADR1(DLX_IDinst_IR_opcode_field[1]),
    .ADR2(DLX_EXinst_N66105),
    .ADR3(\DLX_IDinst_Imm[31] ),
    .O(\CHOICE4686/GROM )
  );
  X_BUF \CHOICE4686/XUSED  (
    .I(\CHOICE4686/FROM ),
    .O(CHOICE4686)
  );
  X_BUF \CHOICE4686/YUSED  (
    .I(\CHOICE4686/GROM ),
    .O(CHOICE4895)
  );
  defparam \DLX_EXinst__n0006<15>21 .INIT = 16'hF200;
  X_LUT4 \DLX_EXinst__n0006<15>21  (
    .ADR0(DLX_EXinst__n0080),
    .ADR1(\DLX_IDinst_Imm[15] ),
    .ADR2(DLX_EXinst__n0079),
    .ADR3(DLX_IDinst_reg_out_A[15]),
    .O(\CHOICE4811/FROM )
  );
  defparam \DLX_EXinst__n0006<13>67 .INIT = 16'hA2A0;
  X_LUT4 \DLX_EXinst__n0006<13>67  (
    .ADR0(DLX_IDinst_reg_out_A[13]),
    .ADR1(\DLX_IDinst_Imm[13] ),
    .ADR2(DLX_EXinst__n0079),
    .ADR3(DLX_EXinst__n0080),
    .O(\CHOICE4811/GROM )
  );
  X_BUF \CHOICE4811/XUSED  (
    .I(\CHOICE4811/FROM ),
    .O(CHOICE4811)
  );
  X_BUF \CHOICE4811/YUSED  (
    .I(\CHOICE4811/GROM ),
    .O(CHOICE4308)
  );
  defparam \DLX_EXinst__n0006<22>28 .INIT = 16'h5404;
  X_LUT4 \DLX_EXinst__n0006<22>28  (
    .ADR0(DLX_IDinst_IR_function_field[4]),
    .ADR1(DLX_EXinst_N64309),
    .ADR2(DLX_IDinst_IR_function_field[2]),
    .ADR3(DLX_EXinst_N64067),
    .O(\CHOICE4107/FROM )
  );
  defparam \DLX_EXinst__n0006<22>41 .INIT = 16'h4404;
  X_LUT4 \DLX_EXinst__n0006<22>41  (
    .ADR0(N109130),
    .ADR1(DLX_EXinst__n0081),
    .ADR2(N127155),
    .ADR3(CHOICE4107),
    .O(\CHOICE4107/GROM )
  );
  X_BUF \CHOICE4107/XUSED  (
    .I(\CHOICE4107/FROM ),
    .O(CHOICE4107)
  );
  X_BUF \CHOICE4107/YUSED  (
    .I(\CHOICE4107/GROM ),
    .O(CHOICE4109)
  );
  defparam \DLX_EXinst__n0006<29>28 .INIT = 16'hBA10;
  X_LUT4 \DLX_EXinst__n0006<29>28  (
    .ADR0(DLX_IDinst_IR_function_field[3]),
    .ADR1(DLX_EXinst_N63129),
    .ADR2(DLX_IDinst_reg_out_A[29]),
    .ADR3(\DLX_EXinst_Mshift__n0027_Sh[21] ),
    .O(\CHOICE5341/FROM )
  );
  defparam \DLX_EXinst__n0006<30>28 .INIT = 16'hBA10;
  X_LUT4 \DLX_EXinst__n0006<30>28  (
    .ADR0(DLX_IDinst_IR_function_field[3]),
    .ADR1(DLX_EXinst_N63129),
    .ADR2(DLX_IDinst_reg_out_A[30]),
    .ADR3(\DLX_EXinst_Mshift__n0027_Sh[22] ),
    .O(\CHOICE5341/GROM )
  );
  X_BUF \CHOICE5341/XUSED  (
    .I(\CHOICE5341/FROM ),
    .O(CHOICE5341)
  );
  X_BUF \CHOICE5341/YUSED  (
    .I(\CHOICE5341/GROM ),
    .O(CHOICE5264)
  );
  defparam \DLX_EXinst__n0006<14>71 .INIT = 16'hCFCE;
  X_LUT4 \DLX_EXinst__n0006<14>71  (
    .ADR0(CHOICE4242),
    .ADR1(CHOICE4248),
    .ADR2(DLX_IDinst_IR_function_field[4]),
    .ADR3(CHOICE4241),
    .O(\CHOICE4249/FROM )
  );
  defparam \DLX_EXinst__n0006<14>98 .INIT = 16'h3332;
  X_LUT4 \DLX_EXinst__n0006<14>98  (
    .ADR0(CHOICE4234),
    .ADR1(DLX_EXinst__n0030),
    .ADR2(CHOICE4233),
    .ADR3(CHOICE4249),
    .O(\CHOICE4249/GROM )
  );
  X_BUF \CHOICE4249/XUSED  (
    .I(\CHOICE4249/FROM ),
    .O(CHOICE4249)
  );
  X_BUF \CHOICE4249/YUSED  (
    .I(\CHOICE4249/GROM ),
    .O(CHOICE4251)
  );
  defparam DLX_IDlc_master_ctrlID__n0001_SW19.INIT = 16'hFF3F;
  X_LUT4 DLX_IDlc_master_ctrlID__n0001_SW19 (
    .ADR0(VCC),
    .ADR1(DLX_IDlc_master_ctrlID_nro),
    .ADR2(DLX_ackin_ID),
    .ADR3(reset_IBUF_3),
    .O(\CHOICE19/FROM )
  );
  defparam DLX_IDlc_master_ctrlID__n0001_SW111.INIT = 16'hF0FF;
  X_LUT4 DLX_IDlc_master_ctrlID__n0001_SW111 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IDlc_md_outp2),
    .ADR3(CHOICE19),
    .O(\CHOICE19/GROM )
  );
  X_BUF \CHOICE19/XUSED  (
    .I(\CHOICE19/FROM ),
    .O(CHOICE19)
  );
  X_BUF \CHOICE19/YUSED  (
    .I(\CHOICE19/GROM ),
    .O(DLX_ackin_ID)
  );
  defparam DLX_EXlc_md_mda33_a1.INIT = 16'h3300;
  X_LUT4 DLX_EXlc_md_mda33_a1 (
    .ADR0(VCC),
    .ADR1(DLX_EXlc_pd_wint5),
    .ADR2(VCC),
    .ADR3(DLX_EXlc_md_wint32),
    .O(\DLX_EXlc_md_wint33/FROM )
  );
  defparam DLX_EXlc_md_mda1_a1.INIT = 16'h2222;
  X_LUT4 DLX_EXlc_md_mda1_a1 (
    .ADR0(DLX_EXlc_ridp3),
    .ADR1(DLX_EXlc_pd_wint5),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_EXlc_md_wint33/GROM )
  );
  X_BUF \DLX_EXlc_md_wint33/XUSED  (
    .I(\DLX_EXlc_md_wint33/FROM ),
    .O(DLX_EXlc_md_wint33)
  );
  X_BUF \DLX_EXlc_md_wint33/YUSED  (
    .I(\DLX_EXlc_md_wint33/GROM ),
    .O(DLX_EXlc_md_wint1)
  );
  defparam \DLX_EXinst__n0006<4>211 .INIT = 16'hC0C0;
  X_LUT4 \DLX_EXinst__n0006<4>211  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[4]),
    .ADR2(DLX_EXinst_N64448),
    .ADR3(VCC),
    .O(\CHOICE4021/FROM )
  );
  defparam \DLX_EXinst__n0006<31>42 .INIT = 16'hEEFE;
  X_LUT4 \DLX_EXinst__n0006<31>42  (
    .ADR0(DLX_EXinst_N64448),
    .ADR1(CHOICE5753),
    .ADR2(N111221),
    .ADR3(DLX_IDinst_reg_out_B[5]),
    .O(\CHOICE4021/GROM )
  );
  X_BUF \CHOICE4021/XUSED  (
    .I(\CHOICE4021/FROM ),
    .O(CHOICE4021)
  );
  X_BUF \CHOICE4021/YUSED  (
    .I(\CHOICE4021/GROM ),
    .O(CHOICE5754)
  );
  defparam \DLX_EXinst__n0006<15>42 .INIT = 16'hE020;
  X_LUT4 \DLX_EXinst__n0006<15>42  (
    .ADR0(N97305),
    .ADR1(DLX_IDinst_IR_function_field[2]),
    .ADR2(DLX_EXinst_N66475),
    .ADR3(DLX_EXinst_N64849),
    .O(\CHOICE4817/FROM )
  );
  defparam \DLX_EXinst__n0006<15>87 .INIT = 16'hFFEE;
  X_LUT4 \DLX_EXinst__n0006<15>87  (
    .ADR0(CHOICE4823),
    .ADR1(CHOICE4828),
    .ADR2(VCC),
    .ADR3(CHOICE4817),
    .O(\CHOICE4817/GROM )
  );
  X_BUF \CHOICE4817/XUSED  (
    .I(\CHOICE4817/FROM ),
    .O(CHOICE4817)
  );
  X_BUF \CHOICE4817/YUSED  (
    .I(\CHOICE4817/GROM ),
    .O(CHOICE4830)
  );
  defparam DLX_IDinst_Ker709891.INIT = 16'h0050;
  X_LUT4 DLX_IDinst_Ker709891 (
    .ADR0(DLX_IDinst_IR_latched[26]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_N70909),
    .ADR3(DLX_IDinst_IR_latched[28]),
    .O(\DLX_IDinst_N70991/FROM )
  );
  defparam DLX_IDinst_Ker70640111.INIT = 16'hCDDD;
  X_LUT4 DLX_IDinst_Ker70640111 (
    .ADR0(DLX_IDinst_N70918),
    .ADR1(DLX_IDinst_IR_latched[30]),
    .ADR2(DLX_IDinst_IR_latched[27]),
    .ADR3(DLX_IDinst_N70991),
    .O(\DLX_IDinst_N70991/GROM )
  );
  X_BUF \DLX_IDinst_N70991/XUSED  (
    .I(\DLX_IDinst_N70991/FROM ),
    .O(DLX_IDinst_N70991)
  );
  X_BUF \DLX_IDinst_N70991/YUSED  (
    .I(\DLX_IDinst_N70991/GROM ),
    .O(CHOICE3353)
  );
  defparam \DLX_EXinst__n0006<19>309_SW0 .INIT = 16'hFCFA;
  X_LUT4 \DLX_EXinst__n0006<19>309_SW0  (
    .ADR0(DLX_EXinst__n0047),
    .ADR1(DLX_EXinst__n0045),
    .ADR2(DLX_EXinst_N64448),
    .ADR3(DLX_IDinst_reg_out_B[19]),
    .O(\N126482/FROM )
  );
  defparam \DLX_EXinst__n0006<31>36 .INIT = 16'hCCAA;
  X_LUT4 \DLX_EXinst__n0006<31>36  (
    .ADR0(DLX_EXinst__n0047),
    .ADR1(DLX_EXinst__n0045),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[31]),
    .O(\N126482/GROM )
  );
  X_BUF \N126482/XUSED  (
    .I(\N126482/FROM ),
    .O(N126482)
  );
  X_BUF \N126482/YUSED  (
    .I(\N126482/GROM ),
    .O(CHOICE5753)
  );
  defparam \DLX_EXinst__n0006<17>207 .INIT = 16'h2000;
  X_LUT4 \DLX_EXinst__n0006<17>207  (
    .ADR0(DLX_EXinst_N66226),
    .ADR1(DLX_EXinst_N62740),
    .ADR2(DLX_IDinst_reg_out_B[4]),
    .ADR3(\DLX_EXinst_Mshift__n0025_Sh[1] ),
    .O(\CHOICE5617/FROM )
  );
  defparam \DLX_EXinst__n0006<0>204 .INIT = 16'h0008;
  X_LUT4 \DLX_EXinst__n0006<0>204  (
    .ADR0(\DLX_EXinst_Mshift__n0025_Sh[0] ),
    .ADR1(DLX_EXinst_N66226),
    .ADR2(DLX_IDinst_reg_out_B[4]),
    .ADR3(DLX_EXinst_N62740),
    .O(\CHOICE5617/GROM )
  );
  X_BUF \CHOICE5617/XUSED  (
    .I(\CHOICE5617/FROM ),
    .O(CHOICE5617)
  );
  X_BUF \CHOICE5617/YUSED  (
    .I(\CHOICE5617/GROM ),
    .O(CHOICE5891)
  );
  defparam \DLX_EXinst__n0006<23>28 .INIT = 16'h00CA;
  X_LUT4 \DLX_EXinst__n0006<23>28  (
    .ADR0(DLX_EXinst_N64314),
    .ADR1(DLX_EXinst_N64072),
    .ADR2(DLX_IDinst_IR_function_field[2]),
    .ADR3(DLX_IDinst_IR_function_field[4]),
    .O(\CHOICE4041/FROM )
  );
  defparam \DLX_EXinst__n0006<23>41 .INIT = 16'h4404;
  X_LUT4 \DLX_EXinst__n0006<23>41  (
    .ADR0(N109130),
    .ADR1(DLX_EXinst__n0081),
    .ADR2(N127189),
    .ADR3(CHOICE4041),
    .O(\CHOICE4041/GROM )
  );
  X_BUF \CHOICE4041/XUSED  (
    .I(\CHOICE4041/FROM ),
    .O(CHOICE4041)
  );
  X_BUF \CHOICE4041/YUSED  (
    .I(\CHOICE4041/GROM ),
    .O(CHOICE4043)
  );
  defparam DLX_IDinst_Ker7066665_SW0.INIT = 16'hA2F7;
  X_LUT4 DLX_IDinst_Ker7066665_SW0 (
    .ADR0(DLX_IFinst_IR_latched[28]),
    .ADR1(CHOICE3267),
    .ADR2(DLX_IFinst_IR_latched[27]),
    .ADR3(DLX_IFinst_IR_latched[30]),
    .O(\N126054/FROM )
  );
  defparam DLX_IDinst_Ker7066665.INIT = 16'h00CD;
  X_LUT4 DLX_IDinst_Ker7066665 (
    .ADR0(DLX_IDinst__n0075),
    .ADR1(DLX_IDinst__n0004),
    .ADR2(DLX_IDinst__n0078),
    .ADR3(N126054),
    .O(\N126054/GROM )
  );
  X_BUF \N126054/XUSED  (
    .I(\N126054/FROM ),
    .O(N126054)
  );
  X_BUF \N126054/YUSED  (
    .I(\N126054/GROM ),
    .O(CHOICE3274)
  );
  defparam DLX_EXinst_Ker6489279.INIT = 16'h1000;
  X_LUT4 DLX_EXinst_Ker6489279 (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(DLX_IDinst_reg_out_B[0]),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(DLX_IDinst_reg_out_B_2_1),
    .O(\CHOICE2548/FROM )
  );
  defparam \DLX_EXinst__n0006<31>71 .INIT = 16'h4450;
  X_LUT4 \DLX_EXinst__n0006<31>71  (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(DLX_IDinst_reg_out_A[29]),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(DLX_IDinst_reg_out_B[1]),
    .O(\CHOICE2548/GROM )
  );
  X_BUF \CHOICE2548/XUSED  (
    .I(\CHOICE2548/FROM ),
    .O(CHOICE2548)
  );
  X_BUF \CHOICE2548/YUSED  (
    .I(\CHOICE2548/GROM ),
    .O(CHOICE5764)
  );
  defparam \DLX_EXinst__n0006<24>23 .INIT = 16'h0A0C;
  X_LUT4 \DLX_EXinst__n0006<24>23  (
    .ADR0(DLX_EXinst_N64077),
    .ADR1(N97960),
    .ADR2(DLX_IDinst_IR_function_field[4]),
    .ADR3(DLX_IDinst_IR_function_field[2]),
    .O(\CHOICE3743/FROM )
  );
  defparam \DLX_EXinst__n0006<24>36 .INIT = 16'hCC80;
  X_LUT4 \DLX_EXinst__n0006<24>36  (
    .ADR0(\DLX_EXinst_Mshift__n0027_Sh[40] ),
    .ADR1(DLX_EXinst_N66202),
    .ADR2(DLX_IDinst_IR_function_field[4]),
    .ADR3(CHOICE3743),
    .O(\CHOICE3743/GROM )
  );
  X_BUF \CHOICE3743/XUSED  (
    .I(\CHOICE3743/FROM ),
    .O(CHOICE3743)
  );
  X_BUF \CHOICE3743/YUSED  (
    .I(\CHOICE3743/GROM ),
    .O(CHOICE3745)
  );
  defparam DLX_EXlc_ridp31.INIT = 16'h0F0F;
  X_LUT4 DLX_EXlc_ridp31 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_EXlc_pd_wint5),
    .ADR3(VCC),
    .O(\DLX_EXlc_ridp3/FROM )
  );
  defparam DLX_EXlc_md_mda2_a1.INIT = 16'h0C0C;
  X_LUT4 DLX_EXlc_md_mda2_a1 (
    .ADR0(VCC),
    .ADR1(DLX_EXlc_md_wint1),
    .ADR2(DLX_EXlc_pd_wint5),
    .ADR3(VCC),
    .O(\DLX_EXlc_ridp3/GROM )
  );
  X_BUF \DLX_EXlc_ridp3/XUSED  (
    .I(\DLX_EXlc_ridp3/FROM ),
    .O(DLX_EXlc_ridp3)
  );
  X_BUF \DLX_EXlc_ridp3/YUSED  (
    .I(\DLX_EXlc_ridp3/GROM ),
    .O(DLX_EXlc_md_wint2)
  );
  defparam \DLX_EXinst__n0006<0>136 .INIT = 16'hEECC;
  X_LUT4 \DLX_EXinst__n0006<0>136  (
    .ADR0(DLX_EXinst__n0045),
    .ADR1(DLX_EXinst_N64448),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[0]),
    .O(\CHOICE5875/FROM )
  );
  defparam \DLX_EXinst__n0006<0>145 .INIT = 16'hCC40;
  X_LUT4 \DLX_EXinst__n0006<0>145  (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(DLX_IDinst_reg_out_A[0]),
    .ADR2(DLX_EXinst__n0047),
    .ADR3(CHOICE5875),
    .O(\CHOICE5875/GROM )
  );
  X_BUF \CHOICE5875/XUSED  (
    .I(\CHOICE5875/FROM ),
    .O(CHOICE5875)
  );
  X_BUF \CHOICE5875/YUSED  (
    .I(\CHOICE5875/GROM ),
    .O(CHOICE5877)
  );
  defparam \DLX_EXinst__n0006<30>88 .INIT = 16'h8040;
  X_LUT4 \DLX_EXinst__n0006<30>88  (
    .ADR0(N127408),
    .ADR1(\DLX_IDinst_Imm[31] ),
    .ADR2(DLX_EXinst_N66105),
    .ADR3(DLX_IDinst_IR_opcode_field[1]),
    .O(\CHOICE5276/FROM )
  );
  defparam \DLX_EXinst__n0006<30>99 .INIT = 16'hFFEA;
  X_LUT4 \DLX_EXinst__n0006<30>99  (
    .ADR0(N126560),
    .ADR1(\DLX_IDinst_Imm[14] ),
    .ADR2(DLX_EXinst__n0077),
    .ADR3(CHOICE5276),
    .O(\CHOICE5276/GROM )
  );
  X_BUF \CHOICE5276/XUSED  (
    .I(\CHOICE5276/FROM ),
    .O(CHOICE5276)
  );
  X_BUF \CHOICE5276/YUSED  (
    .I(\CHOICE5276/GROM ),
    .O(CHOICE5278)
  );
  defparam DLX_EXinst_Ker6514812.INIT = 16'hA808;
  X_LUT4 DLX_EXinst_Ker6514812 (
    .ADR0(DLX_IDinst_IR_function_field_2_1),
    .ADR1(\DLX_EXinst_Mshift__n0024_Sh[25] ),
    .ADR2(DLX_IDinst_IR_function_field_3_1),
    .ADR3(DLX_IDinst_reg_out_A[31]),
    .O(\CHOICE3085/FROM )
  );
  defparam DLX_EXinst_Ker6511326.INIT = 16'h00E4;
  X_LUT4 DLX_EXinst_Ker6511326 (
    .ADR0(DLX_IDinst_IR_function_field_2_1),
    .ADR1(\DLX_EXinst_Mshift__n0024_Sh[25] ),
    .ADR2(\DLX_EXinst_Mshift__n0024_Sh[29] ),
    .ADR3(\DLX_IDinst_Imm[5] ),
    .O(\CHOICE3085/GROM )
  );
  X_BUF \CHOICE3085/XUSED  (
    .I(\CHOICE3085/FROM ),
    .O(CHOICE3085)
  );
  X_BUF \CHOICE3085/YUSED  (
    .I(\CHOICE3085/GROM ),
    .O(CHOICE1991)
  );
  defparam DLX_IDinst__n03641_1_1176.INIT = 16'hFF02;
  X_LUT4 DLX_IDinst__n03641_1_1176 (
    .ADR0(INT_IBUF),
    .ADR1(DLX_IDinst_delay_slot),
    .ADR2(DLX_IDinst_CLI),
    .ADR3(DLX_IDinst__n0070),
    .O(\DLX_IDinst__n03641_1/FROM )
  );
  defparam DLX_IDinst_Ker708191.INIT = 16'h00B7;
  X_LUT4 DLX_IDinst_Ker708191 (
    .ADR0(DLX_IDinst_IR_latched[30]),
    .ADR1(DLX_IDinst_N70991),
    .ADR2(DLX_IDinst_IR_latched[27]),
    .ADR3(DLX_IDinst__n03641_1),
    .O(\DLX_IDinst__n03641_1/GROM )
  );
  X_BUF \DLX_IDinst__n03641_1/XUSED  (
    .I(\DLX_IDinst__n03641_1/FROM ),
    .O(DLX_IDinst__n03641_1)
  );
  X_BUF \DLX_IDinst__n03641_1/YUSED  (
    .I(\DLX_IDinst__n03641_1/GROM ),
    .O(DLX_IDinst_N70821)
  );
  defparam \DLX_IDinst__n0023<0>1 .INIT = 16'hEA00;
  X_LUT4 \DLX_IDinst__n0023<0>1  (
    .ADR0(DLX_IDinst__n0364),
    .ADR1(DLX_IDinst_N69568),
    .ADR2(N102453),
    .ADR3(DLX_IDinst_jtarget[11]),
    .O(\DLX_IDinst_Imm<11>/FROM )
  );
  defparam DLX_IDinst__n00941.INIT = 16'h1100;
  X_LUT4 DLX_IDinst__n00941 (
    .ADR0(DLX_IDinst_N70918),
    .ADR1(DLX_IDinst__n0331),
    .ADR2(VCC),
    .ADR3(DLX_IDinst__n0023[0]),
    .O(DLX_IDinst__n0094)
  );
  X_BUF \DLX_IDinst_Imm<11>/XUSED  (
    .I(\DLX_IDinst_Imm<11>/FROM ),
    .O(DLX_IDinst__n0023[0])
  );
  defparam \DLX_EXinst__n0006<0>314 .INIT = 16'h0080;
  X_LUT4 \DLX_EXinst__n0006<0>314  (
    .ADR0(DLX_IDinst_IR_function_field[5]),
    .ADR1(DLX_IDinst_IR_function_field[3]),
    .ADR2(CHOICE5915),
    .ADR3(DLX_IDinst_IR_function_field[4]),
    .O(\CHOICE5917/FROM )
  );
  defparam \DLX_EXinst__n0006<0>369_SW0_SW0 .INIT = 16'hFF80;
  X_LUT4 \DLX_EXinst__n0006<0>369_SW0_SW0  (
    .ADR0(N111221),
    .ADR1(DLX_IDinst_reg_out_B[5]),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(CHOICE5917),
    .O(\CHOICE5917/GROM )
  );
  X_BUF \CHOICE5917/XUSED  (
    .I(\CHOICE5917/FROM ),
    .O(CHOICE5917)
  );
  X_BUF \CHOICE5917/YUSED  (
    .I(\CHOICE5917/GROM ),
    .O(N127252)
  );
  defparam DLX_EXinst_Ker6515348.INIT = 16'h5700;
  X_LUT4 DLX_EXinst_Ker6515348 (
    .ADR0(DLX_IDinst_IR_function_field_3_1),
    .ADR1(DLX_IDinst_IR_function_field_1_1),
    .ADR2(DLX_IDinst_IR_function_field_2_1),
    .ADR3(\DLX_IDinst_Imm[5] ),
    .O(\CHOICE3068/FROM )
  );
  defparam DLX_EXinst_Ker6512313.INIT = 16'h2AAA;
  X_LUT4 DLX_EXinst_Ker6512313 (
    .ADR0(\DLX_IDinst_Imm[5] ),
    .ADR1(DLX_IDinst_IR_function_field_1_1),
    .ADR2(DLX_IDinst_IR_function_field_2_1),
    .ADR3(DLX_IDinst_IR_function_field_3_1),
    .O(\CHOICE3068/GROM )
  );
  X_BUF \CHOICE3068/XUSED  (
    .I(\CHOICE3068/FROM ),
    .O(CHOICE3068)
  );
  X_BUF \CHOICE3068/YUSED  (
    .I(\CHOICE3068/GROM ),
    .O(CHOICE1861)
  );
  defparam \DLX_EXinst__n0006<3>117 .INIT = 16'h9000;
  X_LUT4 \DLX_EXinst__n0006<3>117  (
    .ADR0(DLX_IDinst_IR_opcode_field[1]),
    .ADR1(N127346),
    .ADR2(DLX_IDinst_IR_function_field[3]),
    .ADR3(DLX_EXinst_N66105),
    .O(\CHOICE5046/FROM )
  );
  defparam \DLX_EXinst__n0006<15>59 .INIT = 16'h8008;
  X_LUT4 \DLX_EXinst__n0006<15>59  (
    .ADR0(\DLX_IDinst_Imm[15] ),
    .ADR1(DLX_EXinst_N66105),
    .ADR2(DLX_IDinst_IR_opcode_field[1]),
    .ADR3(N127294),
    .O(\CHOICE5046/GROM )
  );
  X_BUF \CHOICE5046/XUSED  (
    .I(\CHOICE5046/FROM ),
    .O(CHOICE5046)
  );
  X_BUF \CHOICE5046/YUSED  (
    .I(\CHOICE5046/GROM ),
    .O(CHOICE4823)
  );
  defparam \DLX_EXinst__n0006<25>36 .INIT = 16'h8200;
  X_LUT4 \DLX_EXinst__n0006<25>36  (
    .ADR0(DLX_EXinst_N66105),
    .ADR1(DLX_IDinst_IR_opcode_field[1]),
    .ADR2(N127330),
    .ADR3(\DLX_IDinst_Imm[31] ),
    .O(\CHOICE4751/FROM )
  );
  defparam \DLX_EXinst__n0006<16>35 .INIT = 16'h8200;
  X_LUT4 \DLX_EXinst__n0006<16>35  (
    .ADR0(\DLX_IDinst_Imm[31] ),
    .ADR1(N127290),
    .ADR2(DLX_IDinst_IR_opcode_field[1]),
    .ADR3(DLX_EXinst_N66105),
    .O(\CHOICE4751/GROM )
  );
  X_BUF \CHOICE4751/XUSED  (
    .I(\CHOICE4751/FROM ),
    .O(CHOICE4751)
  );
  X_BUF \CHOICE4751/YUSED  (
    .I(\CHOICE4751/GROM ),
    .O(CHOICE5107)
  );
  defparam DLX_EXinst_Ker6582521.INIT = 16'h2060;
  X_LUT4 DLX_EXinst_Ker6582521 (
    .ADR0(DLX_EXinst_N62733),
    .ADR1(\DLX_IDinst_Imm[5] ),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(DLX_IDinst_IR_function_field_1_1),
    .O(\CHOICE2060/FROM )
  );
  defparam DLX_EXinst_Ker6510811.INIT = 16'h20A0;
  X_LUT4 DLX_EXinst_Ker6510811 (
    .ADR0(\DLX_IDinst_Imm[5] ),
    .ADR1(DLX_IDinst_IR_function_field_2_1),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(DLX_IDinst_IR_function_field_1_1),
    .O(\CHOICE2060/GROM )
  );
  X_BUF \CHOICE2060/XUSED  (
    .I(\CHOICE2060/FROM ),
    .O(CHOICE2060)
  );
  X_BUF \CHOICE2060/YUSED  (
    .I(\CHOICE2060/GROM ),
    .O(CHOICE1951)
  );
  defparam \DLX_EXinst__n0006<17>42 .INIT = 16'h9000;
  X_LUT4 \DLX_EXinst__n0006<17>42  (
    .ADR0(DLX_IDinst_IR_opcode_field[1]),
    .ADR1(N127322),
    .ADR2(DLX_EXinst_N66105),
    .ADR3(\DLX_IDinst_Imm[31] ),
    .O(\CHOICE5587/FROM )
  );
  defparam \DLX_EXinst__n0006<23>85 .INIT = 16'h9000;
  X_LUT4 \DLX_EXinst__n0006<23>85  (
    .ADR0(N127400),
    .ADR1(DLX_IDinst_IR_opcode_field[1]),
    .ADR2(DLX_EXinst_N66105),
    .ADR3(\DLX_IDinst_Imm[31] ),
    .O(\CHOICE5587/GROM )
  );
  X_BUF \CHOICE5587/XUSED  (
    .I(\CHOICE5587/FROM ),
    .O(CHOICE5587)
  );
  X_BUF \CHOICE5587/YUSED  (
    .I(\CHOICE5587/GROM ),
    .O(CHOICE4053)
  );
  defparam \DLX_IDinst__n0023<1>1 .INIT = 16'hE0A0;
  X_LUT4 \DLX_IDinst__n0023<1>1  (
    .ADR0(DLX_IDinst__n0364),
    .ADR1(N102453),
    .ADR2(DLX_IDinst_jtarget[12]),
    .ADR3(DLX_IDinst_N69568),
    .O(\DLX_IDinst_Imm<12>/FROM )
  );
  defparam DLX_IDinst__n00931.INIT = 16'h0500;
  X_LUT4 DLX_IDinst__n00931 (
    .ADR0(DLX_IDinst_N70918),
    .ADR1(VCC),
    .ADR2(DLX_IDinst__n0331),
    .ADR3(DLX_IDinst__n0023[1]),
    .O(DLX_IDinst__n0093)
  );
  X_BUF \DLX_IDinst_Imm<12>/XUSED  (
    .I(\DLX_IDinst_Imm<12>/FROM ),
    .O(DLX_IDinst__n0023[1])
  );
  defparam \DLX_IDinst__n0030<5>1 .INIT = 16'hCC80;
  X_LUT4 \DLX_IDinst__n0030<5>1  (
    .ADR0(N102453),
    .ADR1(DLX_IDinst_jtarget[5]),
    .ADR2(DLX_IDinst_N69568),
    .ADR3(DLX_IDinst__n0364),
    .O(\DLX_IDinst_Imm<5>/FROM )
  );
  defparam DLX_IDinst__n01001.INIT = 16'h0300;
  X_LUT4 DLX_IDinst__n01001 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst__n0331),
    .ADR2(DLX_IDinst_N70918),
    .ADR3(DLX_IDinst__n0030[5]),
    .O(DLX_IDinst__n0100)
  );
  X_BUF \DLX_IDinst_Imm<5>/XUSED  (
    .I(\DLX_IDinst_Imm<5>/FROM ),
    .O(DLX_IDinst__n0030[5])
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<26>11 .INIT = 16'h88C0;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<26>11  (
    .ADR0(DLX_IDinst_reg_out_A[29]),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(DLX_IDinst_reg_out_A[28]),
    .ADR3(DLX_IDinst_reg_out_B[0]),
    .O(\CHOICE1138/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<25>11 .INIT = 16'hC840;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<25>11  (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(DLX_IDinst_reg_out_B[0]),
    .ADR2(DLX_IDinst_reg_out_A[26]),
    .ADR3(DLX_IDinst_reg_out_A[28]),
    .O(\CHOICE1138/GROM )
  );
  X_BUF \CHOICE1138/XUSED  (
    .I(\CHOICE1138/FROM ),
    .O(CHOICE1138)
  );
  X_BUF \CHOICE1138/YUSED  (
    .I(\CHOICE1138/GROM ),
    .O(CHOICE1306)
  );
  defparam DLX_MEMlc_pd_wint11.INIT = 16'h5555;
  X_LUT4 DLX_MEMlc_pd_wint11 (
    .ADR0(DLX_reqout_EX),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_MEMlc_pd_wint1/FROM )
  );
  defparam DLX_MEMlc_md_mda20_a1.INIT = 16'h00CC;
  X_LUT4 DLX_MEMlc_md_mda20_a1 (
    .ADR0(VCC),
    .ADR1(DLX_MEMlc_md_wint19),
    .ADR2(VCC),
    .ADR3(DLX_MEMlc_pd_wint1),
    .O(\DLX_MEMlc_pd_wint1/GROM )
  );
  X_BUF \DLX_MEMlc_pd_wint1/XUSED  (
    .I(\DLX_MEMlc_pd_wint1/FROM ),
    .O(DLX_MEMlc_pd_wint1)
  );
  X_BUF \DLX_MEMlc_pd_wint1/YUSED  (
    .I(\DLX_MEMlc_pd_wint1/GROM ),
    .O(DLX_MEMlc_md_wint20)
  );
  defparam \DLX_EXinst__n0006<19>199 .INIT = 16'hAA20;
  X_LUT4 \DLX_EXinst__n0006<19>199  (
    .ADR0(DLX_IDinst_reg_out_B[19]),
    .ADR1(DLX_IDinst_reg_out_A[19]),
    .ADR2(DLX_EXinst__n0047),
    .ADR3(DLX_EXinst__n0046),
    .O(\CHOICE4980/FROM )
  );
  defparam \DLX_EXinst__n0006<0>183 .INIT = 16'hDC00;
  X_LUT4 \DLX_EXinst__n0006<0>183  (
    .ADR0(DLX_IDinst_reg_out_A[0]),
    .ADR1(DLX_EXinst__n0046),
    .ADR2(DLX_EXinst__n0047),
    .ADR3(DLX_IDinst_reg_out_B[0]),
    .O(\CHOICE4980/GROM )
  );
  X_BUF \CHOICE4980/XUSED  (
    .I(\CHOICE4980/FROM ),
    .O(CHOICE4980)
  );
  X_BUF \CHOICE4980/YUSED  (
    .I(\CHOICE4980/GROM ),
    .O(CHOICE5883)
  );
  defparam DLX_EXinst_Ker6512333.INIT = 16'h2320;
  X_LUT4 DLX_EXinst_Ker6512333 (
    .ADR0(DLX_EXinst_N62941),
    .ADR1(\DLX_IDinst_Imm[5] ),
    .ADR2(DLX_IDinst_IR_function_field_2_1),
    .ADR3(DLX_EXinst_N64859),
    .O(\CHOICE1868/FROM )
  );
  defparam DLX_EXinst_Ker6512336.INIT = 16'hFFA0;
  X_LUT4 DLX_EXinst_Ker6512336 (
    .ADR0(CHOICE1861),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(CHOICE1868),
    .O(\CHOICE1868/GROM )
  );
  X_BUF \CHOICE1868/XUSED  (
    .I(\CHOICE1868/FROM ),
    .O(CHOICE1868)
  );
  X_BUF \CHOICE1868/YUSED  (
    .I(\CHOICE1868/GROM ),
    .O(N101095)
  );
  defparam DLX_EXlc_md_mda32_a1.INIT = 16'h0F00;
  X_LUT4 DLX_EXlc_md_mda32_a1 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_EXlc_pd_wint5),
    .ADR3(DLX_EXlc_md_wint31),
    .O(\DLX_EXlc_md_wint32/FROM )
  );
  defparam DLX_EXlc_md_mda3_a1.INIT = 16'h0F00;
  X_LUT4 DLX_EXlc_md_mda3_a1 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_EXlc_pd_wint5),
    .ADR3(DLX_EXlc_md_wint2),
    .O(\DLX_EXlc_md_wint32/GROM )
  );
  X_BUF \DLX_EXlc_md_wint32/XUSED  (
    .I(\DLX_EXlc_md_wint32/FROM ),
    .O(DLX_EXlc_md_wint32)
  );
  X_BUF \DLX_EXlc_md_wint32/YUSED  (
    .I(\DLX_EXlc_md_wint32/GROM ),
    .O(DLX_EXlc_md_wint3)
  );
  defparam \DLX_EXinst__n0006<0>512 .INIT = 16'h8400;
  X_LUT4 \DLX_EXinst__n0006<0>512  (
    .ADR0(DLX_IDinst_IR_opcode_field[1]),
    .ADR1(DLX_EXinst_N66105),
    .ADR2(N127310),
    .ADR3(DLX_IDinst_IR_function_field[0]),
    .O(\CHOICE5953/FROM )
  );
  defparam \DLX_EXinst__n0006<0>516 .INIT = 16'hFF88;
  X_LUT4 \DLX_EXinst__n0006<0>516  (
    .ADR0(DLX_EXinst__n0016[0]),
    .ADR1(DLX_EXinst__n0128),
    .ADR2(VCC),
    .ADR3(CHOICE5953),
    .O(\CHOICE5953/GROM )
  );
  X_BUF \CHOICE5953/XUSED  (
    .I(\CHOICE5953/FROM ),
    .O(CHOICE5953)
  );
  X_BUF \CHOICE5953/YUSED  (
    .I(\CHOICE5953/GROM ),
    .O(CHOICE5954)
  );
  defparam DLX_EXinst_Ker6510824.INIT = 16'h0E02;
  X_LUT4 DLX_EXinst_Ker6510824 (
    .ADR0(\DLX_EXinst_Mshift__n0024_Sh[26] ),
    .ADR1(DLX_IDinst_IR_function_field_2_1),
    .ADR2(\DLX_IDinst_Imm[5] ),
    .ADR3(\DLX_EXinst_Mshift__n0024_Sh[30] ),
    .O(\CHOICE1957/FROM )
  );
  defparam \DLX_EXinst__n0006<1>120 .INIT = 16'hC888;
  X_LUT4 \DLX_EXinst__n0006<1>120  (
    .ADR0(CHOICE1911),
    .ADR1(DLX_EXinst_N66060),
    .ADR2(CHOICE1904),
    .ADR3(\DLX_IDinst_Imm[5] ),
    .O(\CHOICE1957/GROM )
  );
  X_BUF \CHOICE1957/XUSED  (
    .I(\CHOICE1957/FROM ),
    .O(CHOICE1957)
  );
  X_BUF \CHOICE1957/YUSED  (
    .I(\CHOICE1957/GROM ),
    .O(CHOICE5684)
  );
  defparam \DLX_IDinst__n0023<2>1 .INIT = 16'hE0C0;
  X_LUT4 \DLX_IDinst__n0023<2>1  (
    .ADR0(N102453),
    .ADR1(DLX_IDinst__n0364),
    .ADR2(DLX_IDinst_jtarget[13]),
    .ADR3(DLX_IDinst_N69568),
    .O(\DLX_IDinst_Imm<13>/FROM )
  );
  defparam DLX_IDinst__n00921.INIT = 16'h0300;
  X_LUT4 DLX_IDinst__n00921 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_N70918),
    .ADR2(DLX_IDinst__n0331),
    .ADR3(DLX_IDinst__n0023[2]),
    .O(DLX_IDinst__n0092)
  );
  X_BUF \DLX_IDinst_Imm<13>/XUSED  (
    .I(\DLX_IDinst_Imm<13>/FROM ),
    .O(DLX_IDinst__n0023[2])
  );
  defparam \DLX_EXinst__n0006<1>203 .INIT = 16'h0C0A;
  X_LUT4 \DLX_EXinst__n0006<1>203  (
    .ADR0(DLX_EXinst_N64864),
    .ADR1(DLX_EXinst_N64255),
    .ADR2(DLX_IDinst_reg_out_B[3]),
    .ADR3(DLX_IDinst_reg_out_B[0]),
    .O(\CHOICE5704/FROM )
  );
  defparam \DLX_EXinst__n0006<1>217 .INIT = 16'h5540;
  X_LUT4 \DLX_EXinst__n0006<1>217  (
    .ADR0(DLX_IDinst_reg_out_B[2]),
    .ADR1(DLX_IDinst_reg_out_B[3]),
    .ADR2(\DLX_EXinst_Mshift__n0023_Sh[9] ),
    .ADR3(CHOICE5704),
    .O(\CHOICE5704/GROM )
  );
  X_BUF \CHOICE5704/XUSED  (
    .I(\CHOICE5704/FROM ),
    .O(CHOICE5704)
  );
  X_BUF \CHOICE5704/YUSED  (
    .I(\CHOICE5704/GROM ),
    .O(CHOICE5706)
  );
  defparam \DLX_EXinst__n0006<22>100 .INIT = 16'hFFEC;
  X_LUT4 \DLX_EXinst__n0006<22>100  (
    .ADR0(DLX_EXinst__n0016[22]),
    .ADR1(N126524),
    .ADR2(DLX_EXinst__n0128),
    .ADR3(CHOICE4119),
    .O(\CHOICE4123/FROM )
  );
  defparam \DLX_EXinst__n0006<24>91 .INIT = 16'hFFEC;
  X_LUT4 \DLX_EXinst__n0006<24>91  (
    .ADR0(DLX_EXinst__n0016[24]),
    .ADR1(N126597),
    .ADR2(DLX_EXinst__n0128),
    .ADR3(CHOICE3755),
    .O(\CHOICE4123/GROM )
  );
  X_BUF \CHOICE4123/XUSED  (
    .I(\CHOICE4123/FROM ),
    .O(CHOICE4123)
  );
  X_BUF \CHOICE4123/YUSED  (
    .I(\CHOICE4123/GROM ),
    .O(CHOICE3759)
  );
  defparam \DLX_EXinst__n0006<25>51 .INIT = 16'hAC00;
  X_LUT4 \DLX_EXinst__n0006<25>51  (
    .ADR0(DLX_EXinst_N64304),
    .ADR1(N97665),
    .ADR2(DLX_IDinst_IR_function_field[2]),
    .ADR3(DLX_EXinst__n0081),
    .O(\CHOICE4758/FROM )
  );
  defparam \DLX_EXinst__n0006<25>75_SW0 .INIT = 16'hFFC0;
  X_LUT4 \DLX_EXinst__n0006<25>75_SW0  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst__n0082),
    .ADR2(\DLX_EXinst_Mshift__n0028_Sh[57] ),
    .ADR3(CHOICE4758),
    .O(\CHOICE4758/GROM )
  );
  X_BUF \CHOICE4758/XUSED  (
    .I(\CHOICE4758/FROM ),
    .O(CHOICE4758)
  );
  X_BUF \CHOICE4758/YUSED  (
    .I(\CHOICE4758/GROM ),
    .O(N126306)
  );
  defparam \DLX_EXinst__n0006<0>277 .INIT = 16'h0202;
  X_LUT4 \DLX_EXinst__n0006<0>277  (
    .ADR0(DLX_IDinst_IR_function_field[1]),
    .ADR1(N126107),
    .ADR2(DLX_IDinst_IR_function_field[2]),
    .ADR3(VCC),
    .O(\CHOICE5914/FROM )
  );
  defparam \DLX_EXinst__n0006<0>284 .INIT = 16'hFF54;
  X_LUT4 \DLX_EXinst__n0006<0>284  (
    .ADR0(DLX_IDinst_IR_function_field[1]),
    .ADR1(CHOICE5905),
    .ADR2(CHOICE5899),
    .ADR3(CHOICE5914),
    .O(\CHOICE5914/GROM )
  );
  X_BUF \CHOICE5914/XUSED  (
    .I(\CHOICE5914/FROM ),
    .O(CHOICE5914)
  );
  X_BUF \CHOICE5914/YUSED  (
    .I(\CHOICE5914/GROM ),
    .O(CHOICE5915)
  );
  defparam DLX_EXinst_Ker6435714.INIT = 16'h2320;
  X_LUT4 DLX_EXinst_Ker6435714 (
    .ADR0(DLX_IDinst_reg_out_A[25]),
    .ADR1(DLX_IDinst_reg_out_B[0]),
    .ADR2(DLX_IDinst_reg_out_B[1]),
    .ADR3(DLX_IDinst_reg_out_A[27]),
    .O(\CHOICE1825/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<25>26 .INIT = 16'h5044;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<25>26  (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(DLX_IDinst_reg_out_A[25]),
    .ADR2(DLX_IDinst_reg_out_A[27]),
    .ADR3(DLX_IDinst_reg_out_B[1]),
    .O(\CHOICE1825/GROM )
  );
  X_BUF \CHOICE1825/XUSED  (
    .I(\CHOICE1825/FROM ),
    .O(CHOICE1825)
  );
  X_BUF \CHOICE1825/YUSED  (
    .I(\CHOICE1825/GROM ),
    .O(CHOICE1312)
  );
  defparam \DLX_IDinst__n0023<3>1 .INIT = 16'hE0C0;
  X_LUT4 \DLX_IDinst__n0023<3>1  (
    .ADR0(N102453),
    .ADR1(DLX_IDinst__n0364),
    .ADR2(DLX_IDinst_jtarget[14]),
    .ADR3(DLX_IDinst_N69568),
    .O(\DLX_IDinst_Imm<14>/FROM )
  );
  defparam DLX_IDinst__n00911.INIT = 16'h1100;
  X_LUT4 DLX_IDinst__n00911 (
    .ADR0(DLX_IDinst__n0331),
    .ADR1(DLX_IDinst_N70918),
    .ADR2(VCC),
    .ADR3(DLX_IDinst__n0023[3]),
    .O(DLX_IDinst__n0091)
  );
  X_BUF \DLX_IDinst_Imm<14>/XUSED  (
    .I(\DLX_IDinst_Imm<14>/FROM ),
    .O(DLX_IDinst__n0023[3])
  );
  defparam \DLX_EXinst__n0006<2>117 .INIT = 16'h9000;
  X_LUT4 \DLX_EXinst__n0006<2>117  (
    .ADR0(DLX_IDinst_IR_opcode_field[1]),
    .ADR1(N127306),
    .ADR2(DLX_EXinst_N66105),
    .ADR3(DLX_IDinst_IR_function_field[2]),
    .O(\CHOICE5517/FROM )
  );
  defparam \DLX_EXinst__n0006<1>117 .INIT = 16'h8040;
  X_LUT4 \DLX_EXinst__n0006<1>117  (
    .ADR0(DLX_IDinst_IR_opcode_field[1]),
    .ADR1(DLX_EXinst_N66105),
    .ADR2(DLX_IDinst_IR_function_field[1]),
    .ADR3(N127314),
    .O(\CHOICE5517/GROM )
  );
  X_BUF \CHOICE5517/XUSED  (
    .I(\CHOICE5517/FROM ),
    .O(CHOICE5517)
  );
  X_BUF \CHOICE5517/YUSED  (
    .I(\CHOICE5517/GROM ),
    .O(CHOICE5683)
  );
  defparam DLX_EXinst_Ker6510860.INIT = 16'hAFAE;
  X_LUT4 DLX_EXinst_Ker6510860 (
    .ADR0(CHOICE1962),
    .ADR1(CHOICE1957),
    .ADR2(DLX_IDinst_IR_function_field_3_1),
    .ADR3(CHOICE1951),
    .O(\N101641/FROM )
  );
  defparam \DLX_EXinst__n0006<10>62 .INIT = 16'h8000;
  X_LUT4 \DLX_EXinst__n0006<10>62  (
    .ADR0(CHOICE3377),
    .ADR1(DLX_IDinst_IR_function_field[4]),
    .ADR2(CHOICE3408),
    .ADR3(N101641),
    .O(\N101641/GROM )
  );
  X_BUF \N101641/XUSED  (
    .I(\N101641/FROM ),
    .O(N101641)
  );
  X_BUF \N101641/YUSED  (
    .I(\N101641/GROM ),
    .O(CHOICE4505)
  );
  defparam DLX_EXinst_Ker6582020.INIT = 16'h0040;
  X_LUT4 DLX_EXinst_Ker6582020 (
    .ADR0(DLX_IDinst_IR_function_field_3_1),
    .ADR1(\DLX_EXinst_Mshift__n0024_Sh[61] ),
    .ADR2(\DLX_IDinst_Imm[5] ),
    .ADR3(DLX_IDinst_IR_function_field_2_1),
    .O(\CHOICE2046/FROM )
  );
  defparam DLX_EXinst_Ker6511813.INIT = 16'hE2AA;
  X_LUT4 DLX_EXinst_Ker6511813 (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(DLX_IDinst_IR_function_field_2_1),
    .ADR2(\DLX_EXinst_Mshift__n0024_Sh[61] ),
    .ADR3(DLX_IDinst_IR_function_field_3_1),
    .O(\CHOICE2046/GROM )
  );
  X_BUF \CHOICE2046/XUSED  (
    .I(\CHOICE2046/FROM ),
    .O(CHOICE2046)
  );
  X_BUF \CHOICE2046/YUSED  (
    .I(\CHOICE2046/GROM ),
    .O(CHOICE1904)
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<25>28 .INIT = 16'hFAFA;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<25>28  (
    .ADR0(CHOICE1306),
    .ADR1(VCC),
    .ADR2(CHOICE1312),
    .ADR3(VCC),
    .O(\DLX_EXinst_Mshift__n0023_Sh<25>/FROM )
  );
  defparam DLX_EXinst_Ker6488227.INIT = 16'h4540;
  X_LUT4 DLX_EXinst_Ker6488227 (
    .ADR0(DLX_IDinst_reg_out_B[5]),
    .ADR1(\DLX_EXinst_Mshift__n0023_Sh[29] ),
    .ADR2(DLX_IDinst_reg_out_B_2_1),
    .ADR3(\DLX_EXinst_Mshift__n0023_Sh[25] ),
    .O(\DLX_EXinst_Mshift__n0023_Sh<25>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0023_Sh<25>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0023_Sh<25>/FROM ),
    .O(\DLX_EXinst_Mshift__n0023_Sh[25] )
  );
  X_BUF \DLX_EXinst_Mshift__n0023_Sh<25>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0023_Sh<25>/GROM ),
    .O(CHOICE3145)
  );
  defparam DLX_EXlc_md_mda29_a1.INIT = 16'h00AA;
  X_LUT4 DLX_EXlc_md_mda29_a1 (
    .ADR0(DLX_EXlc_md_wint28),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_EXlc_pd_wint5),
    .O(\DLX_EXlc_md_wint29/FROM )
  );
  defparam DLX_EXlc_md_mda4_a1.INIT = 16'h00CC;
  X_LUT4 DLX_EXlc_md_mda4_a1 (
    .ADR0(VCC),
    .ADR1(DLX_EXlc_md_wint3),
    .ADR2(VCC),
    .ADR3(DLX_EXlc_pd_wint5),
    .O(\DLX_EXlc_md_wint29/GROM )
  );
  X_BUF \DLX_EXlc_md_wint29/XUSED  (
    .I(\DLX_EXlc_md_wint29/FROM ),
    .O(DLX_EXlc_md_wint29)
  );
  X_BUF \DLX_EXlc_md_wint29/YUSED  (
    .I(\DLX_EXlc_md_wint29/GROM ),
    .O(DLX_EXlc_md_wint4)
  );
  defparam \DLX_EXinst_Mshift__n0026_Sh<24> .INIT = 16'hCCAA;
  X_LUT4 \DLX_EXinst_Mshift__n0026_Sh<24>  (
    .ADR0(DLX_EXinst_N63780),
    .ADR1(N94107),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[0]),
    .O(\DLX_EXinst_Mshift__n0026_Sh<24>/FROM )
  );
  defparam DLX_EXinst_Ker632971.INIT = 16'hFBC8;
  X_LUT4 DLX_EXinst_Ker632971 (
    .ADR0(CHOICE1156),
    .ADR1(DLX_IDinst_reg_out_B_2_1),
    .ADR2(CHOICE1150),
    .ADR3(\DLX_EXinst_Mshift__n0026_Sh[24] ),
    .O(\DLX_EXinst_Mshift__n0026_Sh<24>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0026_Sh<24>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0026_Sh<24>/FROM ),
    .O(\DLX_EXinst_Mshift__n0026_Sh[24] )
  );
  X_BUF \DLX_EXinst_Mshift__n0026_Sh<24>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0026_Sh<24>/GROM ),
    .O(DLX_EXinst_N63299)
  );
  defparam \DLX_EXinst__n0006<1>129 .INIT = 16'hFEFA;
  X_LUT4 \DLX_EXinst__n0006<1>129  (
    .ADR0(CHOICE5684),
    .ADR1(N126571),
    .ADR2(CHOICE5683),
    .ADR3(DLX_EXinst_N66475),
    .O(\CHOICE5686/FROM )
  );
  defparam \DLX_EXinst__n0006<1>160 .INIT = 16'h5554;
  X_LUT4 \DLX_EXinst__n0006<1>160  (
    .ADR0(DLX_EXinst__n0030),
    .ADR1(CHOICE5659),
    .ADR2(CHOICE5663),
    .ADR3(CHOICE5686),
    .O(\CHOICE5686/GROM )
  );
  X_BUF \CHOICE5686/XUSED  (
    .I(\CHOICE5686/FROM ),
    .O(CHOICE5686)
  );
  X_BUF \CHOICE5686/YUSED  (
    .I(\CHOICE5686/GROM ),
    .O(CHOICE5688)
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<29>1 .INIT = 16'hAACC;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<29>1  (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(DLX_EXinst_N62721),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[1]),
    .O(\DLX_EXinst_Mshift__n0023_Sh<29>/FROM )
  );
  defparam DLX_EXinst_Ker6505423.INIT = 16'hA0A0;
  X_LUT4 DLX_EXinst_Ker6505423 (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(VCC),
    .ADR2(CHOICE1771),
    .ADR3(VCC),
    .O(\DLX_EXinst_Mshift__n0023_Sh<29>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0023_Sh<29>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0023_Sh<29>/FROM ),
    .O(\DLX_EXinst_Mshift__n0023_Sh[29] )
  );
  X_BUF \DLX_EXinst_Mshift__n0023_Sh<29>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0023_Sh<29>/GROM ),
    .O(N100490)
  );
  defparam \DLX_EXinst__n0006<0>449 .INIT = 16'h0044;
  X_LUT4 \DLX_EXinst__n0006<0>449  (
    .ADR0(N126092),
    .ADR1(DLX_IDinst_IR_opcode_field[1]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_IR_opcode_field[2]),
    .O(\CHOICE5943/FROM )
  );
  defparam \DLX_EXinst__n0006<0>456 .INIT = 16'hFF54;
  X_LUT4 \DLX_EXinst__n0006<0>456  (
    .ADR0(DLX_IDinst_IR_opcode_field[1]),
    .ADR1(CHOICE5934),
    .ADR2(CHOICE5928),
    .ADR3(CHOICE5943),
    .O(\CHOICE5943/GROM )
  );
  X_BUF \CHOICE5943/XUSED  (
    .I(\CHOICE5943/FROM ),
    .O(CHOICE5943)
  );
  X_BUF \CHOICE5943/YUSED  (
    .I(\CHOICE5943/GROM ),
    .O(CHOICE5944)
  );
  defparam \DLX_IDinst__n0023<4>1 .INIT = 16'hF800;
  X_LUT4 \DLX_IDinst__n0023<4>1  (
    .ADR0(N102453),
    .ADR1(DLX_IDinst_N69568),
    .ADR2(DLX_IDinst__n0364),
    .ADR3(DLX_IDinst_jtarget[15]),
    .O(\DLX_IDinst_Imm<15>/FROM )
  );
  defparam DLX_IDinst__n00901.INIT = 16'h0300;
  X_LUT4 DLX_IDinst__n00901 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_N70918),
    .ADR2(DLX_IDinst__n0331),
    .ADR3(DLX_IDinst__n0023[4]),
    .O(DLX_IDinst__n0090)
  );
  X_BUF \DLX_IDinst_Imm<15>/XUSED  (
    .I(\DLX_IDinst_Imm<15>/FROM ),
    .O(DLX_IDinst__n0023[4])
  );
  defparam DLX_EXinst_Ker6510856.INIT = 16'h3000;
  X_LUT4 DLX_EXinst_Ker6510856 (
    .ADR0(VCC),
    .ADR1(\DLX_IDinst_Imm[5] ),
    .ADR2(DLX_IDinst_IR_function_field_3_1),
    .ADR3(DLX_IDinst_reg_out_A[31]),
    .O(\CHOICE1962/FROM )
  );
  defparam DLX_EXinst_Ker6511364.INIT = 16'hFF0E;
  X_LUT4 DLX_EXinst_Ker6511364 (
    .ADR0(CHOICE1985),
    .ADR1(CHOICE1991),
    .ADR2(DLX_IDinst_IR_function_field_3_1),
    .ADR3(CHOICE1962),
    .O(\CHOICE1962/GROM )
  );
  X_BUF \CHOICE1962/XUSED  (
    .I(\CHOICE1962/FROM ),
    .O(CHOICE1962)
  );
  X_BUF \CHOICE1962/YUSED  (
    .I(\CHOICE1962/GROM ),
    .O(N101839)
  );
  defparam \DLX_EXinst__n0006<1>306 .INIT = 16'h0E0C;
  X_LUT4 \DLX_EXinst__n0006<1>306  (
    .ADR0(DLX_EXinst_N66383),
    .ADR1(CHOICE5722),
    .ADR2(N110935),
    .ADR3(\DLX_EXinst_Mshift__n0026_Sh[49] ),
    .O(\CHOICE5724/FROM )
  );
  defparam \DLX_EXinst__n0006<1>320 .INIT = 16'hFFAA;
  X_LUT4 \DLX_EXinst__n0006<1>320  (
    .ADR0(CHOICE5728),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(CHOICE5724),
    .O(\CHOICE5724/GROM )
  );
  X_BUF \CHOICE5724/XUSED  (
    .I(\CHOICE5724/FROM ),
    .O(CHOICE5724)
  );
  X_BUF \CHOICE5724/YUSED  (
    .I(\CHOICE5724/GROM ),
    .O(CHOICE5729)
  );
  defparam DLX_EXinst_Ker6426225.INIT = 16'h5044;
  X_LUT4 DLX_EXinst_Ker6426225 (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(DLX_EXinst_N64587),
    .ADR2(DLX_EXinst_N63409),
    .ADR3(DLX_IDinst_reg_out_B[3]),
    .O(\CHOICE1036/FROM )
  );
  defparam DLX_EXinst_Ker6426228.INIT = 16'hFFAA;
  X_LUT4 DLX_EXinst_Ker6426228 (
    .ADR0(CHOICE1030),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(CHOICE1036),
    .O(\CHOICE1036/GROM )
  );
  X_BUF \CHOICE1036/XUSED  (
    .I(\CHOICE1036/FROM ),
    .O(CHOICE1036)
  );
  X_BUF \CHOICE1036/YUSED  (
    .I(\CHOICE1036/GROM ),
    .O(N96153)
  );
  defparam \DLX_EXinst__n0006<26>51 .INIT = 16'hD800;
  X_LUT4 \DLX_EXinst__n0006<26>51  (
    .ADR0(DLX_IDinst_IR_function_field[2]),
    .ADR1(DLX_EXinst_N64309),
    .ADR2(N98032),
    .ADR3(DLX_EXinst__n0081),
    .O(\CHOICE4693/FROM )
  );
  defparam \DLX_EXinst__n0006<26>75_SW0 .INIT = 16'hFFA0;
  X_LUT4 \DLX_EXinst__n0006<26>75_SW0  (
    .ADR0(\DLX_EXinst_Mshift__n0028_Sh[58] ),
    .ADR1(VCC),
    .ADR2(DLX_EXinst__n0082),
    .ADR3(CHOICE4693),
    .O(\CHOICE4693/GROM )
  );
  X_BUF \CHOICE4693/XUSED  (
    .I(\CHOICE4693/FROM ),
    .O(CHOICE4693)
  );
  X_BUF \CHOICE4693/YUSED  (
    .I(\CHOICE4693/GROM ),
    .O(N126383)
  );
  defparam \DLX_EXinst__n0006<25>75 .INIT = 16'hF444;
  X_LUT4 \DLX_EXinst__n0006<25>75  (
    .ADR0(N109130),
    .ADR1(N126306),
    .ADR2(N110065),
    .ADR3(N101839),
    .O(\CHOICE4763/FROM )
  );
  defparam \DLX_EXinst__n0006<25>110_SW0 .INIT = 16'hD5C0;
  X_LUT4 \DLX_EXinst__n0006<25>110_SW0  (
    .ADR0(DLX_IDinst_IR_function_field[4]),
    .ADR1(DLX_EXinst__n0077),
    .ADR2(\DLX_IDinst_Imm[9] ),
    .ADR3(CHOICE4763),
    .O(\CHOICE4763/GROM )
  );
  X_BUF \CHOICE4763/XUSED  (
    .I(\CHOICE4763/FROM ),
    .O(CHOICE4763)
  );
  X_BUF \CHOICE4763/YUSED  (
    .I(\CHOICE4763/GROM ),
    .O(N126301)
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<26>25 .INIT = 16'h0C0A;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<26>25  (
    .ADR0(DLX_IDinst_reg_out_A[26]),
    .ADR1(DLX_IDinst_reg_out_A[27]),
    .ADR2(DLX_IDinst_reg_out_B[1]),
    .ADR3(DLX_IDinst_reg_out_B[0]),
    .O(\CHOICE1144/FROM )
  );
  defparam DLX_EXinst_Ker64872113.INIT = 16'h0C08;
  X_LUT4 DLX_EXinst_Ker64872113 (
    .ADR0(CHOICE1138),
    .ADR1(DLX_IDinst_reg_out_B_2_1),
    .ADR2(DLX_IDinst_reg_out_B_3_1),
    .ADR3(CHOICE1144),
    .O(\CHOICE1144/GROM )
  );
  X_BUF \CHOICE1144/XUSED  (
    .I(\CHOICE1144/FROM ),
    .O(CHOICE1144)
  );
  X_BUF \CHOICE1144/YUSED  (
    .I(\CHOICE1144/GROM ),
    .O(CHOICE3208)
  );
  defparam \DLX_EXinst_Mshift__n0026_Sh<50> .INIT = 16'hACAC;
  X_LUT4 \DLX_EXinst_Mshift__n0026_Sh<50>  (
    .ADR0(N94255),
    .ADR1(DLX_EXinst_N64334),
    .ADR2(DLX_IDinst_reg_out_B_2_1),
    .ADR3(VCC),
    .O(\DLX_EXinst_Mshift__n0026_Sh<50>/FROM )
  );
  defparam \DLX_EXinst__n0006<18>302_SW0 .INIT = 16'hFCF0;
  X_LUT4 \DLX_EXinst__n0006<18>302_SW0  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst__n0049),
    .ADR2(CHOICE5471),
    .ADR3(\DLX_EXinst_Mshift__n0026_Sh[50] ),
    .O(\DLX_EXinst_Mshift__n0026_Sh<50>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0026_Sh<50>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0026_Sh<50>/FROM ),
    .O(\DLX_EXinst_Mshift__n0026_Sh[50] )
  );
  X_BUF \DLX_EXinst_Mshift__n0026_Sh<50>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0026_Sh<50>/GROM ),
    .O(N126370)
  );
  defparam \DLX_EXinst__n0006<1>334 .INIT = 16'hFEFC;
  X_LUT4 \DLX_EXinst__n0006<1>334  (
    .ADR0(N101725),
    .ADR1(CHOICE5716),
    .ADR2(CHOICE5729),
    .ADR3(DLX_EXinst_ALU_result[1]),
    .O(\CHOICE5730/FROM )
  );
  defparam \DLX_EXinst__n0006<1>371_SW0 .INIT = 16'hFFF8;
  X_LUT4 \DLX_EXinst__n0006<1>371_SW0  (
    .ADR0(DLX_EXinst__n0114),
    .ADR1(DLX_EXinst__n0016[1]),
    .ADR2(CHOICE5709),
    .ADR3(CHOICE5730),
    .O(\CHOICE5730/GROM )
  );
  X_BUF \CHOICE5730/XUSED  (
    .I(\CHOICE5730/FROM ),
    .O(CHOICE5730)
  );
  X_BUF \CHOICE5730/YUSED  (
    .I(\CHOICE5730/GROM ),
    .O(N127163)
  );
  defparam \DLX_EXinst__n0006<3>117_SW0 .INIT = 16'h0055;
  X_LUT4 \DLX_EXinst__n0006<3>117_SW0  (
    .ADR0(DLX_IDinst_reg_out_A[3]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_IR_opcode_field[0]),
    .O(\N127346/FROM )
  );
  defparam \DLX_EXinst__n0006<0>512_SW0 .INIT = 16'h0055;
  X_LUT4 \DLX_EXinst__n0006<0>512_SW0  (
    .ADR0(DLX_IDinst_reg_out_A[0]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_IR_opcode_field[0]),
    .O(\N127346/GROM )
  );
  X_BUF \N127346/XUSED  (
    .I(\N127346/FROM ),
    .O(N127346)
  );
  X_BUF \N127346/YUSED  (
    .I(\N127346/GROM ),
    .O(N127310)
  );
  defparam DLX_EXinst_Ker6511836.INIT = 16'h0B08;
  X_LUT4 DLX_EXinst_Ker6511836 (
    .ADR0(DLX_EXinst_N62936),
    .ADR1(DLX_IDinst_IR_function_field_2_1),
    .ADR2(\DLX_IDinst_Imm[5] ),
    .ADR3(DLX_EXinst_N64854),
    .O(\CHOICE1911/FROM )
  );
  defparam DLX_EXinst_Ker6511839.INIT = 16'hFFC0;
  X_LUT4 DLX_EXinst_Ker6511839 (
    .ADR0(VCC),
    .ADR1(\DLX_IDinst_Imm[5] ),
    .ADR2(CHOICE1904),
    .ADR3(CHOICE1911),
    .O(\CHOICE1911/GROM )
  );
  X_BUF \CHOICE1911/XUSED  (
    .I(\CHOICE1911/FROM ),
    .O(CHOICE1911)
  );
  X_BUF \CHOICE1911/YUSED  (
    .I(\CHOICE1911/GROM ),
    .O(N101338)
  );
  defparam DLX_EXinst__n012719.INIT = 16'hFFFD;
  X_LUT4 DLX_EXinst__n012719 (
    .ADR0(DLX_IDinst_IR_function_field[0]),
    .ADR1(DLX_IDinst_IR_function_field[3]),
    .ADR2(DLX_IDinst_IR_function_field[2]),
    .ADR3(DLX_IDinst_IR_function_field[1]),
    .O(\CHOICE1972/FROM )
  );
  defparam \DLX_EXinst__n0006<19>14 .INIT = 16'h0020;
  X_LUT4 \DLX_EXinst__n0006<19>14  (
    .ADR0(\DLX_EXinst_Mshift__n0027_Sh[3] ),
    .ADR1(DLX_IDinst_IR_function_field[2]),
    .ADR2(DLX_EXinst_N66087),
    .ADR3(DLX_IDinst_IR_function_field[3]),
    .O(\CHOICE1972/GROM )
  );
  X_BUF \CHOICE1972/XUSED  (
    .I(\CHOICE1972/FROM ),
    .O(CHOICE1972)
  );
  X_BUF \CHOICE1972/YUSED  (
    .I(\CHOICE1972/GROM ),
    .O(CHOICE4944)
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<26>28 .INIT = 16'hFFAA;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<26>28  (
    .ADR0(CHOICE1138),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(CHOICE1144),
    .O(\DLX_EXinst_Mshift__n0023_Sh<26>/FROM )
  );
  defparam DLX_EXinst_Ker6488725.INIT = 16'h0D08;
  X_LUT4 DLX_EXinst_Ker6488725 (
    .ADR0(DLX_IDinst_reg_out_B_2_1),
    .ADR1(\DLX_EXinst_Mshift__n0023_Sh[30] ),
    .ADR2(DLX_IDinst_reg_out_B[5]),
    .ADR3(\DLX_EXinst_Mshift__n0023_Sh[26] ),
    .O(\DLX_EXinst_Mshift__n0023_Sh<26>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0023_Sh<26>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0023_Sh<26>/FROM ),
    .O(\DLX_EXinst_Mshift__n0023_Sh[26] )
  );
  X_BUF \DLX_EXinst_Mshift__n0023_Sh<26>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0023_Sh<26>/GROM ),
    .O(CHOICE3038)
  );
  defparam \DLX_EXinst__n0006<1>271 .INIT = 16'hFF88;
  X_LUT4 \DLX_EXinst__n0006<1>271  (
    .ADR0(DLX_EXinst__n0045),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N64448),
    .O(\CHOICE5714/FROM )
  );
  defparam \DLX_EXinst__n0006<1>280 .INIT = 16'hF040;
  X_LUT4 \DLX_EXinst__n0006<1>280  (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(DLX_EXinst__n0047),
    .ADR2(DLX_IDinst_reg_out_A[1]),
    .ADR3(CHOICE5714),
    .O(\CHOICE5714/GROM )
  );
  X_BUF \CHOICE5714/XUSED  (
    .I(\CHOICE5714/FROM ),
    .O(CHOICE5714)
  );
  X_BUF \CHOICE5714/YUSED  (
    .I(\CHOICE5714/GROM ),
    .O(CHOICE5716)
  );
  defparam DLX_EXinst_Ker6450325.INIT = 16'h00CA;
  X_LUT4 DLX_EXinst_Ker6450325 (
    .ADR0(DLX_EXinst_N64909),
    .ADR1(DLX_EXinst_N62976),
    .ADR2(DLX_IDinst_IR_function_field[0]),
    .ADR3(DLX_IDinst_IR_function_field[3]),
    .O(\CHOICE1276/FROM )
  );
  defparam DLX_EXinst_Ker6450328.INIT = 16'hFFCC;
  X_LUT4 DLX_EXinst_Ker6450328 (
    .ADR0(VCC),
    .ADR1(CHOICE1270),
    .ADR2(VCC),
    .ADR3(CHOICE1276),
    .O(\CHOICE1276/GROM )
  );
  X_BUF \CHOICE1276/XUSED  (
    .I(\CHOICE1276/FROM ),
    .O(CHOICE1276)
  );
  X_BUF \CHOICE1276/YUSED  (
    .I(\CHOICE1276/GROM ),
    .O(N97593)
  );
  defparam \DLX_EXinst__n0006<10>138 .INIT = 16'hA2A0;
  X_LUT4 \DLX_EXinst__n0006<10>138  (
    .ADR0(DLX_IDinst_reg_out_B[10]),
    .ADR1(DLX_IDinst_reg_out_A[10]),
    .ADR2(DLX_EXinst__n0046),
    .ADR3(DLX_EXinst__n0047),
    .O(\CHOICE4520/FROM )
  );
  defparam \DLX_EXinst__n0006<1>319 .INIT = 16'h88C8;
  X_LUT4 \DLX_EXinst__n0006<1>319  (
    .ADR0(DLX_EXinst__n0046),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(DLX_EXinst__n0047),
    .ADR3(DLX_IDinst_reg_out_A[1]),
    .O(\CHOICE4520/GROM )
  );
  X_BUF \CHOICE4520/XUSED  (
    .I(\CHOICE4520/FROM ),
    .O(CHOICE4520)
  );
  X_BUF \CHOICE4520/YUSED  (
    .I(\CHOICE4520/GROM ),
    .O(CHOICE5728)
  );
  defparam DLX_EXlc_md_mda28_a1.INIT = 16'h5500;
  X_LUT4 DLX_EXlc_md_mda28_a1 (
    .ADR0(DLX_EXlc_pd_wint5),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_EXlc_md_wint27),
    .O(\DLX_EXlc_md_wint28/FROM )
  );
  defparam DLX_EXlc_md_mda5_a1.INIT = 16'h4444;
  X_LUT4 DLX_EXlc_md_mda5_a1 (
    .ADR0(DLX_EXlc_pd_wint5),
    .ADR1(DLX_EXlc_md_wint4),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_EXlc_md_wint28/GROM )
  );
  X_BUF \DLX_EXlc_md_wint28/XUSED  (
    .I(\DLX_EXlc_md_wint28/FROM ),
    .O(DLX_EXlc_md_wint28)
  );
  X_BUF \DLX_EXlc_md_wint28/YUSED  (
    .I(\DLX_EXlc_md_wint28/GROM ),
    .O(DLX_EXlc_md_wint5)
  );
  defparam DLX_EXinst_Ker6488711.INIT = 16'h7000;
  X_LUT4 DLX_EXinst_Ker6488711 (
    .ADR0(DLX_IDinst_reg_out_B_2_1),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(DLX_IDinst_reg_out_B[5]),
    .O(\CHOICE3032/FROM )
  );
  defparam \DLX_EXinst__n0006<2>120 .INIT = 16'hE0C0;
  X_LUT4 \DLX_EXinst__n0006<2>120  (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(CHOICE1868),
    .ADR2(DLX_EXinst_N66060),
    .ADR3(CHOICE1861),
    .O(\CHOICE3032/GROM )
  );
  X_BUF \CHOICE3032/XUSED  (
    .I(\CHOICE3032/FROM ),
    .O(CHOICE3032)
  );
  X_BUF \CHOICE3032/YUSED  (
    .I(\CHOICE3032/GROM ),
    .O(CHOICE5518)
  );
  defparam vga_top_vga1_Ker73377_SW0.INIT = 16'hFFFE;
  X_LUT4 vga_top_vga1_Ker73377_SW0 (
    .ADR0(vga_top_vga1_hcounter[12]),
    .ADR1(vga_top_vga1_hcounter[13]),
    .ADR2(vga_top_vga1_hcounter[11]),
    .ADR3(vga_top_vga1_hcounter[10]),
    .O(\N98808/FROM )
  );
  defparam vga_top_vga1_Ker73377.INIT = 16'h0001;
  X_LUT4 vga_top_vga1_Ker73377 (
    .ADR0(vga_top_vga1_hcounter[15]),
    .ADR1(vga_top_vga1_hcounter[14]),
    .ADR2(vga_top_vga1_hcounter[6]),
    .ADR3(N98808),
    .O(\N98808/GROM )
  );
  X_BUF \N98808/XUSED  (
    .I(\N98808/FROM ),
    .O(N98808)
  );
  X_BUF \N98808/YUSED  (
    .I(\N98808/GROM ),
    .O(vga_top_vga1_N73379)
  );
  defparam \DLX_EXinst__n0006<0>729 .INIT = 16'h3332;
  X_LUT4 \DLX_EXinst__n0006<0>729  (
    .ADR0(CHOICE5954),
    .ADR1(DLX_EXinst__n0030),
    .ADR2(N126252),
    .ADR3(CHOICE5983),
    .O(\DLX_EXinst_ALU_result<0>/FROM )
  );
  defparam \DLX_EXinst__n0006<0>753 .INIT = 16'h0504;
  X_LUT4 \DLX_EXinst__n0006<0>753  (
    .ADR0(DLX_IDinst_counter[0]),
    .ADR1(CHOICE5921),
    .ADR2(DLX_IDinst_counter[1]),
    .ADR3(CHOICE5991),
    .O(\DLX_EXinst_ALU_result<0>/GROM )
  );
  X_BUF \DLX_EXinst_ALU_result<0>/XUSED  (
    .I(\DLX_EXinst_ALU_result<0>/FROM ),
    .O(CHOICE5991)
  );
  X_BUF \DLX_EXinst_ALU_result<0>/YUSED  (
    .I(\DLX_EXinst_ALU_result<0>/GROM ),
    .O(N125635)
  );
  defparam DLX_EXinst_Ker6512856_SW0.INIT = 16'hE222;
  X_LUT4 DLX_EXinst_Ker6512856_SW0 (
    .ADR0(DLX_EXinst_N64849),
    .ADR1(DLX_IDinst_IR_function_field_2_1),
    .ADR2(DLX_IDinst_IR_function_field_3_1),
    .ADR3(DLX_IDinst_reg_out_A[31]),
    .O(\N125971/FROM )
  );
  defparam DLX_EXinst_Ker6515312.INIT = 16'hA0C0;
  X_LUT4 DLX_EXinst_Ker6515312 (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(\DLX_EXinst_Mshift__n0024_Sh[26] ),
    .ADR2(DLX_IDinst_IR_function_field_2_1),
    .ADR3(DLX_IDinst_IR_function_field_3_1),
    .O(\N125971/GROM )
  );
  X_BUF \N125971/XUSED  (
    .I(\N125971/FROM ),
    .O(N125971)
  );
  X_BUF \N125971/YUSED  (
    .I(\N125971/GROM ),
    .O(CHOICE3058)
  );
  defparam \DLX_EXinst__n0006<0>674 .INIT = 16'hCE00;
  X_LUT4 \DLX_EXinst__n0006<0>674  (
    .ADR0(DLX_EXinst__n0080),
    .ADR1(DLX_EXinst__n0079),
    .ADR2(DLX_IDinst_IR_function_field[0]),
    .ADR3(DLX_IDinst_reg_out_A[0]),
    .O(\CHOICE5982/FROM )
  );
  defparam \DLX_EXinst__n0006<0>678 .INIT = 16'hFF54;
  X_LUT4 \DLX_EXinst__n0006<0>678  (
    .ADR0(DLX_IDinst_IR_function_field[4]),
    .ADR1(CHOICE5976),
    .ADR2(CHOICE5973),
    .ADR3(CHOICE5982),
    .O(\CHOICE5982/GROM )
  );
  X_BUF \CHOICE5982/XUSED  (
    .I(\CHOICE5982/FROM ),
    .O(CHOICE5982)
  );
  X_BUF \CHOICE5982/YUSED  (
    .I(\CHOICE5982/GROM ),
    .O(CHOICE5983)
  );
  defparam \DLX_EXinst__n0006<1>371 .INIT = 16'hF808;
  X_LUT4 \DLX_EXinst__n0006<1>371  (
    .ADR0(DLX_EXinst__n0016[1]),
    .ADR1(DLX_EXinst__n0128),
    .ADR2(DLX_EXinst__n0030),
    .ADR3(N127163),
    .O(\DLX_EXinst_ALU_result<1>/FROM )
  );
  defparam \DLX_EXinst__n0006<1>411 .INIT = 16'hEEEA;
  X_LUT4 \DLX_EXinst__n0006<1>411  (
    .ADR0(DLX_EXinst_N63689),
    .ADR1(DLX_EXinst__n0149),
    .ADR2(CHOICE5688),
    .ADR3(CHOICE5733),
    .O(\DLX_EXinst_ALU_result<1>/GROM )
  );
  X_BUF \DLX_EXinst_ALU_result<1>/XUSED  (
    .I(\DLX_EXinst_ALU_result<1>/FROM ),
    .O(CHOICE5733)
  );
  X_BUF \DLX_EXinst_ALU_result<1>/YUSED  (
    .I(\DLX_EXinst_ALU_result<1>/GROM ),
    .O(N124056)
  );
  defparam \DLX_EXinst__n0006<5>147 .INIT = 16'hCA00;
  X_LUT4 \DLX_EXinst__n0006<5>147  (
    .ADR0(\DLX_EXinst_Mshift__n0026_Sh[13] ),
    .ADR1(\DLX_EXinst_Mshift__n0026_Sh[17] ),
    .ADR2(DLX_IDinst_reg_out_B[2]),
    .ADR3(DLX_IDinst_reg_out_B[3]),
    .O(\CHOICE4453/FROM )
  );
  defparam \DLX_EXinst__n0006<1>187 .INIT = 16'hD800;
  X_LUT4 \DLX_EXinst__n0006<1>187  (
    .ADR0(DLX_IDinst_reg_out_B[3]),
    .ADR1(\DLX_EXinst_Mshift__n0026_Sh[13] ),
    .ADR2(\DLX_EXinst_Mshift__n0023_Sh[5] ),
    .ADR3(DLX_IDinst_reg_out_B[2]),
    .O(\CHOICE4453/GROM )
  );
  X_BUF \CHOICE4453/XUSED  (
    .I(\CHOICE4453/FROM ),
    .O(CHOICE4453)
  );
  X_BUF \CHOICE4453/YUSED  (
    .I(\CHOICE4453/GROM ),
    .O(CHOICE5696)
  );
  defparam \DLX_EXinst__n0006<26>75 .INIT = 16'hDC50;
  X_LUT4 \DLX_EXinst__n0006<26>75  (
    .ADR0(N109130),
    .ADR1(N110065),
    .ADR2(N126383),
    .ADR3(N101641),
    .O(\CHOICE4698/FROM )
  );
  defparam \DLX_EXinst__n0006<26>110_SW0 .INIT = 16'hB3A0;
  X_LUT4 \DLX_EXinst__n0006<26>110_SW0  (
    .ADR0(\DLX_IDinst_Imm[10] ),
    .ADR1(DLX_IDinst_IR_function_field[4]),
    .ADR2(DLX_EXinst__n0077),
    .ADR3(CHOICE4698),
    .O(\CHOICE4698/GROM )
  );
  X_BUF \CHOICE4698/XUSED  (
    .I(\CHOICE4698/FROM ),
    .O(CHOICE4698)
  );
  X_BUF \CHOICE4698/YUSED  (
    .I(\CHOICE4698/GROM ),
    .O(N126375)
  );
  X_ONE \vga_top_vga1_videoon/LOGIC_ONE_1177  (
    .O(\vga_top_vga1_videoon/LOGIC_ONE )
  );
  defparam DLX_EXinst_Ker6514347.INIT = 16'h0400;
  X_LUT4 DLX_EXinst_Ker6514347 (
    .ADR0(N110935),
    .ADR1(DLX_EXinst_N63299),
    .ADR2(DLX_IDinst_reg_out_B_3_1),
    .ADR3(DLX_EXinst__n0049),
    .O(\CHOICE1379/FROM )
  );
  defparam DLX_EXinst_Ker6514350.INIT = 16'hFFC0;
  X_LUT4 DLX_EXinst_Ker6514350 (
    .ADR0(VCC),
    .ADR1(N127223),
    .ADR2(N111221),
    .ADR3(CHOICE1379),
    .O(\CHOICE1379/GROM )
  );
  X_BUF \CHOICE1379/XUSED  (
    .I(\CHOICE1379/FROM ),
    .O(CHOICE1379)
  );
  X_BUF \CHOICE1379/YUSED  (
    .I(\CHOICE1379/GROM ),
    .O(N98218)
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<28>10 .INIT = 16'h88A0;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<28>10  (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(DLX_IDinst_reg_out_A[31]),
    .ADR2(DLX_IDinst_reg_out_A[29]),
    .ADR3(DLX_IDinst_reg_out_B[1]),
    .O(\CHOICE1150/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0026_Sh<60>1 .INIT = 16'h1110;
  X_LUT4 \DLX_EXinst_Mshift__n0026_Sh<60>1  (
    .ADR0(DLX_IDinst_reg_out_B_3_1),
    .ADR1(DLX_IDinst_reg_out_B_2_1),
    .ADR2(CHOICE1156),
    .ADR3(CHOICE1150),
    .O(\CHOICE1150/GROM )
  );
  X_BUF \CHOICE1150/XUSED  (
    .I(\CHOICE1150/FROM ),
    .O(CHOICE1150)
  );
  X_BUF \CHOICE1150/YUSED  (
    .I(\CHOICE1150/GROM ),
    .O(\DLX_EXinst_Mshift__n0026_Sh[60] )
  );
  defparam DLX_EXinst_Ker6582563.INIT = 16'h0200;
  X_LUT4 DLX_EXinst_Ker6582563 (
    .ADR0(DLX_EXinst_N66507),
    .ADR1(DLX_IDinst_IR_function_field_3_1),
    .ADR2(DLX_IDinst_IR_function_field_2_1),
    .ADR3(\DLX_EXinst_Mshift__n0028_Sh[30] ),
    .O(\CHOICE2069/FROM )
  );
  defparam DLX_EXinst_Ker6515316.INIT = 16'h0B08;
  X_LUT4 DLX_EXinst_Ker6515316 (
    .ADR0(\DLX_EXinst_Mshift__n0024_Sh[30] ),
    .ADR1(DLX_IDinst_IR_function_field_3_1),
    .ADR2(DLX_IDinst_IR_function_field_2_1),
    .ADR3(\DLX_EXinst_Mshift__n0028_Sh[22] ),
    .O(\CHOICE2069/GROM )
  );
  X_BUF \CHOICE2069/XUSED  (
    .I(\CHOICE2069/FROM ),
    .O(CHOICE2069)
  );
  X_BUF \CHOICE2069/YUSED  (
    .I(\CHOICE2069/GROM ),
    .O(CHOICE3060)
  );
  defparam DLX_EXlc_md_mda25_a1.INIT = 16'h4444;
  X_LUT4 DLX_EXlc_md_mda25_a1 (
    .ADR0(DLX_EXlc_pd_wint5),
    .ADR1(DLX_EXlc_md_wint24),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_EXlc_md_wint25/FROM )
  );
  defparam DLX_EXlc_md_mda6_a1.INIT = 16'h5050;
  X_LUT4 DLX_EXlc_md_mda6_a1 (
    .ADR0(DLX_EXlc_pd_wint5),
    .ADR1(VCC),
    .ADR2(DLX_EXlc_md_wint5),
    .ADR3(VCC),
    .O(\DLX_EXlc_md_wint25/GROM )
  );
  X_BUF \DLX_EXlc_md_wint25/XUSED  (
    .I(\DLX_EXlc_md_wint25/FROM ),
    .O(DLX_EXlc_md_wint25)
  );
  X_BUF \DLX_EXlc_md_wint25/YUSED  (
    .I(\DLX_EXlc_md_wint25/GROM ),
    .O(DLX_EXlc_md_wint6)
  );
  defparam \DLX_EXinst__n0006<2>240 .INIT = 16'h5400;
  X_LUT4 \DLX_EXinst__n0006<2>240  (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(CHOICE5540),
    .ADR2(CHOICE5530),
    .ADR3(DLX_EXinst_N62631),
    .O(\CHOICE5542/FROM )
  );
  defparam \DLX_EXinst__n0006<2>255 .INIT = 16'hFF80;
  X_LUT4 \DLX_EXinst__n0006<2>255  (
    .ADR0(N111221),
    .ADR1(N101009),
    .ADR2(DLX_IDinst_reg_out_B[4]),
    .ADR3(CHOICE5542),
    .O(\CHOICE5542/GROM )
  );
  X_BUF \CHOICE5542/XUSED  (
    .I(\CHOICE5542/FROM ),
    .O(CHOICE5542)
  );
  X_BUF \CHOICE5542/YUSED  (
    .I(\CHOICE5542/GROM ),
    .O(CHOICE5543)
  );
  defparam \DLX_EXinst__n0006<22>152 .INIT = 16'h8C88;
  X_LUT4 \DLX_EXinst__n0006<22>152  (
    .ADR0(DLX_EXinst__n0046),
    .ADR1(DLX_IDinst_reg_out_B[22]),
    .ADR2(DLX_IDinst_reg_out_A[22]),
    .ADR3(DLX_EXinst__n0047),
    .O(\CHOICE4130/FROM )
  );
  defparam \DLX_EXinst__n0006<2>320 .INIT = 16'hDC00;
  X_LUT4 \DLX_EXinst__n0006<2>320  (
    .ADR0(DLX_IDinst_reg_out_A[2]),
    .ADR1(DLX_EXinst__n0046),
    .ADR2(DLX_EXinst__n0047),
    .ADR3(DLX_IDinst_reg_out_B[2]),
    .O(\CHOICE4130/GROM )
  );
  X_BUF \CHOICE4130/XUSED  (
    .I(\CHOICE4130/FROM ),
    .O(CHOICE4130)
  );
  X_BUF \CHOICE4130/YUSED  (
    .I(\CHOICE4130/GROM ),
    .O(CHOICE5562)
  );
  defparam \DLX_EXinst__n0006<6>147 .INIT = 16'hB080;
  X_LUT4 \DLX_EXinst__n0006<6>147  (
    .ADR0(\DLX_EXinst_Mshift__n0026_Sh[18] ),
    .ADR1(DLX_IDinst_reg_out_B[2]),
    .ADR2(DLX_IDinst_reg_out_B[3]),
    .ADR3(\DLX_EXinst_Mshift__n0026_Sh[14] ),
    .O(\CHOICE4385/FROM )
  );
  defparam \DLX_EXinst__n0006<1>297 .INIT = 16'h0400;
  X_LUT4 \DLX_EXinst__n0006<1>297  (
    .ADR0(DLX_IDinst_reg_out_B[3]),
    .ADR1(DLX_EXinst_N66535),
    .ADR2(DLX_IDinst_reg_out_B[2]),
    .ADR3(\DLX_EXinst_Mshift__n0025_Sh[1] ),
    .O(\CHOICE4385/GROM )
  );
  X_BUF \CHOICE4385/XUSED  (
    .I(\CHOICE4385/FROM ),
    .O(CHOICE4385)
  );
  X_BUF \CHOICE4385/YUSED  (
    .I(\CHOICE4385/GROM ),
    .O(CHOICE5722)
  );
  defparam \DLX_EXinst__n0006<2>129 .INIT = 16'hFEEE;
  X_LUT4 \DLX_EXinst__n0006<2>129  (
    .ADR0(CHOICE5517),
    .ADR1(CHOICE5518),
    .ADR2(DLX_EXinst_N66475),
    .ADR3(N126297),
    .O(\CHOICE5520/FROM )
  );
  defparam \DLX_EXinst__n0006<2>160 .INIT = 16'h5554;
  X_LUT4 \DLX_EXinst__n0006<2>160  (
    .ADR0(DLX_EXinst__n0030),
    .ADR1(CHOICE5497),
    .ADR2(CHOICE5493),
    .ADR3(CHOICE5520),
    .O(\CHOICE5520/GROM )
  );
  X_BUF \CHOICE5520/XUSED  (
    .I(\CHOICE5520/FROM ),
    .O(CHOICE5520)
  );
  X_BUF \CHOICE5520/YUSED  (
    .I(\CHOICE5520/GROM ),
    .O(CHOICE5522)
  );
  defparam \DLX_EXinst__n0006<0>697 .INIT = 16'hECCC;
  X_LUT4 \DLX_EXinst__n0006<0>697  (
    .ADR0(DLX_IDinst_IR_function_field[4]),
    .ADR1(N126811),
    .ADR2(DLX_EXinst_N63185),
    .ADR3(\DLX_EXinst_Mshift__n0024_Sh[80] ),
    .O(\CHOICE5988/FROM )
  );
  defparam \DLX_EXinst__n0006<0>729_SW0 .INIT = 16'hFF80;
  X_LUT4 \DLX_EXinst__n0006<0>729_SW0  (
    .ADR0(CHOICE5944),
    .ADR1(DLX_EXinst_N66443),
    .ADR2(DLX_IDinst_IR_opcode_field[4]),
    .ADR3(CHOICE5988),
    .O(\CHOICE5988/GROM )
  );
  X_BUF \CHOICE5988/XUSED  (
    .I(\CHOICE5988/FROM ),
    .O(CHOICE5988)
  );
  X_BUF \CHOICE5988/YUSED  (
    .I(\CHOICE5988/GROM ),
    .O(N126252)
  );
  defparam DLX_EXinst_Ker6487712.INIT = 16'hACA0;
  X_LUT4 DLX_EXinst_Ker6487712 (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(\DLX_EXinst_Mshift__n0023_Sh[27] ),
    .ADR2(DLX_IDinst_reg_out_B_3_1),
    .ADR3(DLX_IDinst_reg_out_B_2_1),
    .O(\CHOICE2980/FROM )
  );
  defparam DLX_EXinst_Ker6514350_SW0.INIT = 16'h0AAC;
  X_LUT4 DLX_EXinst_Ker6514350_SW0 (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(DLX_EXinst_N63299),
    .ADR2(DLX_IDinst_reg_out_B_3_1),
    .ADR3(DLX_IDinst_reg_out_B[5]),
    .O(\CHOICE2980/GROM )
  );
  X_BUF \CHOICE2980/XUSED  (
    .I(\CHOICE2980/FROM ),
    .O(CHOICE2980)
  );
  X_BUF \CHOICE2980/YUSED  (
    .I(\CHOICE2980/GROM ),
    .O(N127223)
  );
  defparam \DLX_EXinst__n0006<2>307 .INIT = 16'h5450;
  X_LUT4 \DLX_EXinst__n0006<2>307  (
    .ADR0(N110935),
    .ADR1(DLX_EXinst_N66383),
    .ADR2(CHOICE5556),
    .ADR3(\DLX_EXinst_Mshift__n0026_Sh[50] ),
    .O(\CHOICE5558/FROM )
  );
  defparam \DLX_EXinst__n0006<2>321 .INIT = 16'hFFAA;
  X_LUT4 \DLX_EXinst__n0006<2>321  (
    .ADR0(CHOICE5562),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(CHOICE5558),
    .O(\CHOICE5558/GROM )
  );
  X_BUF \CHOICE5558/XUSED  (
    .I(\CHOICE5558/FROM ),
    .O(CHOICE5558)
  );
  X_BUF \CHOICE5558/YUSED  (
    .I(\CHOICE5558/GROM ),
    .O(CHOICE5563)
  );
  defparam \DLX_EXinst_Mshift__n0024_Sh<25>_SW0 .INIT = 16'hAAF0;
  X_LUT4 \DLX_EXinst_Mshift__n0024_Sh<25>_SW0  (
    .ADR0(DLX_IDinst_reg_out_A[28]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[26]),
    .ADR3(DLX_IDinst_IR_function_field_1_1),
    .O(\N94205/FROM )
  );
  defparam \DLX_EXinst__n0006<28>28 .INIT = 16'hAA30;
  X_LUT4 \DLX_EXinst__n0006<28>28  (
    .ADR0(\DLX_EXinst_Mshift__n0027_Sh[20] ),
    .ADR1(DLX_EXinst_N63129),
    .ADR2(DLX_IDinst_reg_out_A[28]),
    .ADR3(DLX_IDinst_IR_function_field[3]),
    .O(\N94205/GROM )
  );
  X_BUF \N94205/XUSED  (
    .I(\N94205/FROM ),
    .O(N94205)
  );
  X_BUF \N94205/YUSED  (
    .I(\N94205/GROM ),
    .O(CHOICE5189)
  );
  defparam \DLX_EXinst_Mshift__n0026_Sh<30>1 .INIT = 16'h5044;
  X_LUT4 \DLX_EXinst_Mshift__n0026_Sh<30>1  (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(DLX_IDinst_reg_out_A[30]),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(DLX_IDinst_reg_out_B[0]),
    .O(\DLX_EXinst_Mshift__n0026_Sh<30>/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<28>26 .INIT = 16'h4540;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<28>26  (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(DLX_IDinst_reg_out_A[30]),
    .ADR2(DLX_IDinst_reg_out_B[1]),
    .ADR3(DLX_IDinst_reg_out_A[28]),
    .O(\DLX_EXinst_Mshift__n0026_Sh<30>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0026_Sh<30>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0026_Sh<30>/FROM ),
    .O(\DLX_EXinst_Mshift__n0026_Sh[30] )
  );
  X_BUF \DLX_EXinst_Mshift__n0026_Sh<30>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0026_Sh<30>/GROM ),
    .O(CHOICE1156)
  );
  defparam DLX_EXinst_Ker6515349.INIT = 16'h8888;
  X_LUT4 DLX_EXinst_Ker6515349 (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(CHOICE3068),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\CHOICE3069/FROM )
  );
  defparam DLX_EXinst_Ker65153107_SW0.INIT = 16'hFF32;
  X_LUT4 DLX_EXinst_Ker65153107_SW0 (
    .ADR0(CHOICE3060),
    .ADR1(\DLX_IDinst_Imm[5] ),
    .ADR2(CHOICE3058),
    .ADR3(CHOICE3069),
    .O(\CHOICE3069/GROM )
  );
  X_BUF \CHOICE3069/XUSED  (
    .I(\CHOICE3069/FROM ),
    .O(CHOICE3069)
  );
  X_BUF \CHOICE3069/YUSED  (
    .I(\CHOICE3069/GROM ),
    .O(N126469)
  );
  defparam DLX_EXlc_md_mda24_a1.INIT = 16'h00AA;
  X_LUT4 DLX_EXlc_md_mda24_a1 (
    .ADR0(DLX_EXlc_md_wint23),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_EXlc_pd_wint5),
    .O(\DLX_EXlc_md_wint24/FROM )
  );
  defparam DLX_EXlc_md_mda7_a1.INIT = 16'h3030;
  X_LUT4 DLX_EXlc_md_mda7_a1 (
    .ADR0(VCC),
    .ADR1(DLX_EXlc_pd_wint5),
    .ADR2(DLX_EXlc_md_wint6),
    .ADR3(VCC),
    .O(\DLX_EXlc_md_wint24/GROM )
  );
  X_BUF \DLX_EXlc_md_wint24/XUSED  (
    .I(\DLX_EXlc_md_wint24/FROM ),
    .O(DLX_EXlc_md_wint24)
  );
  X_BUF \DLX_EXlc_md_wint24/YUSED  (
    .I(\DLX_EXlc_md_wint24/GROM ),
    .O(DLX_EXlc_md_wint7)
  );
  defparam \DLX_EXinst_Mshift__n0026_Sh<6>1 .INIT = 16'hF5A0;
  X_LUT4 \DLX_EXinst_Mshift__n0026_Sh<6>1  (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N63785),
    .ADR3(DLX_EXinst_N62946),
    .O(\DLX_EXinst_Mshift__n0026_Sh<6>/FROM )
  );
  defparam \DLX_EXinst__n0006<6>161 .INIT = 16'h0D08;
  X_LUT4 \DLX_EXinst__n0006<6>161  (
    .ADR0(DLX_IDinst_reg_out_B[2]),
    .ADR1(\DLX_EXinst_Mshift__n0026_Sh[10] ),
    .ADR2(DLX_IDinst_reg_out_B[3]),
    .ADR3(\DLX_EXinst_Mshift__n0026_Sh[6] ),
    .O(\DLX_EXinst_Mshift__n0026_Sh<6>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0026_Sh<6>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0026_Sh<6>/FROM ),
    .O(\DLX_EXinst_Mshift__n0026_Sh[6] )
  );
  X_BUF \DLX_EXinst_Mshift__n0026_Sh<6>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0026_Sh<6>/GROM ),
    .O(CHOICE4391)
  );
  defparam \DLX_EXinst__n0006<10>213 .INIT = 16'hF888;
  X_LUT4 \DLX_EXinst__n0006<10>213  (
    .ADR0(DLX_EXinst_ALU_result[10]),
    .ADR1(N101725),
    .ADR2(DLX_IDinst_reg_out_B[4]),
    .ADR3(N107934),
    .O(\CHOICE4537/FROM )
  );
  defparam \DLX_EXinst__n0006<2>335 .INIT = 16'hFEEE;
  X_LUT4 \DLX_EXinst__n0006<2>335  (
    .ADR0(CHOICE5550),
    .ADR1(CHOICE5563),
    .ADR2(DLX_EXinst_ALU_result[2]),
    .ADR3(N101725),
    .O(\CHOICE4537/GROM )
  );
  X_BUF \CHOICE4537/XUSED  (
    .I(\CHOICE4537/FROM ),
    .O(CHOICE4537)
  );
  X_BUF \CHOICE4537/YUSED  (
    .I(\CHOICE4537/GROM ),
    .O(CHOICE5564)
  );
  defparam \DLX_EXinst__n0006<2>272 .INIT = 16'hEECC;
  X_LUT4 \DLX_EXinst__n0006<2>272  (
    .ADR0(DLX_IDinst_reg_out_B[2]),
    .ADR1(DLX_EXinst_N64448),
    .ADR2(VCC),
    .ADR3(DLX_EXinst__n0045),
    .O(\CHOICE5548/FROM )
  );
  defparam \DLX_EXinst__n0006<2>281 .INIT = 16'hAA20;
  X_LUT4 \DLX_EXinst__n0006<2>281  (
    .ADR0(DLX_IDinst_reg_out_A[2]),
    .ADR1(DLX_IDinst_reg_out_B[2]),
    .ADR2(DLX_EXinst__n0047),
    .ADR3(CHOICE5548),
    .O(\CHOICE5548/GROM )
  );
  X_BUF \CHOICE5548/XUSED  (
    .I(\CHOICE5548/FROM ),
    .O(CHOICE5548)
  );
  X_BUF \CHOICE5548/YUSED  (
    .I(\CHOICE5548/GROM ),
    .O(CHOICE5550)
  );
  defparam \DLX_EXinst__n0006<30>216 .INIT = 16'h0400;
  X_LUT4 \DLX_EXinst__n0006<30>216  (
    .ADR0(DLX_IDinst_reg_out_B[3]),
    .ADR1(DLX_EXinst_N66392),
    .ADR2(DLX_IDinst_reg_out_B[2]),
    .ADR3(\DLX_EXinst_Mshift__n0026_Sh[30] ),
    .O(\CHOICE5300/FROM )
  );
  defparam \DLX_EXinst__n0006<2>186 .INIT = 16'h8C80;
  X_LUT4 \DLX_EXinst__n0006<2>186  (
    .ADR0(\DLX_EXinst_Mshift__n0026_Sh[14] ),
    .ADR1(DLX_IDinst_reg_out_B[2]),
    .ADR2(DLX_IDinst_reg_out_B[3]),
    .ADR3(\DLX_EXinst_Mshift__n0026_Sh[6] ),
    .O(\CHOICE5300/GROM )
  );
  X_BUF \CHOICE5300/XUSED  (
    .I(\CHOICE5300/FROM ),
    .O(CHOICE5300)
  );
  X_BUF \CHOICE5300/YUSED  (
    .I(\CHOICE5300/GROM ),
    .O(CHOICE5530)
  );
  defparam DLX_EXinst_Ker6540425.INIT = 16'h00D8;
  X_LUT4 DLX_EXinst_Ker6540425 (
    .ADR0(DLX_IDinst_IR_function_field[0]),
    .ADR1(DLX_EXinst_N62811),
    .ADR2(DLX_EXinst_N63309),
    .ADR3(DLX_IDinst_IR_function_field_3_1),
    .O(\CHOICE1349/FROM )
  );
  defparam DLX_EXinst_Ker6540428.INIT = 16'hFFAA;
  X_LUT4 DLX_EXinst_Ker6540428 (
    .ADR0(CHOICE1343),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(CHOICE1349),
    .O(\CHOICE1349/GROM )
  );
  X_BUF \CHOICE1349/XUSED  (
    .I(\CHOICE1349/FROM ),
    .O(CHOICE1349)
  );
  X_BUF \CHOICE1349/YUSED  (
    .I(\CHOICE1349/GROM ),
    .O(N98032)
  );
  defparam DLX_EXinst_Ker6539410.INIT = 16'hC840;
  X_LUT4 DLX_EXinst_Ker6539410 (
    .ADR0(DLX_IDinst_IR_function_field[0]),
    .ADR1(DLX_IDinst_IR_function_field_3_1),
    .ADR2(DLX_EXinst_N62991),
    .ADR3(DLX_EXinst_N63499),
    .O(\CHOICE1102/FROM )
  );
  defparam DLX_EXinst_Ker6541411.INIT = 16'hE400;
  X_LUT4 DLX_EXinst_Ker6541411 (
    .ADR0(DLX_IDinst_IR_function_field[0]),
    .ADR1(DLX_EXinst_N63454),
    .ADR2(DLX_EXinst_N62786),
    .ADR3(DLX_IDinst_IR_function_field_3_1),
    .O(\CHOICE1102/GROM )
  );
  X_BUF \CHOICE1102/XUSED  (
    .I(\CHOICE1102/FROM ),
    .O(CHOICE1102)
  );
  X_BUF \CHOICE1102/YUSED  (
    .I(\CHOICE1102/GROM ),
    .O(CHOICE1331)
  );
  defparam \DLX_EXinst_Mshift__n0026_Sh<21>1 .INIT = 16'hFA0A;
  X_LUT4 \DLX_EXinst_Mshift__n0026_Sh<21>1  (
    .ADR0(DLX_EXinst_N63061),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[0]),
    .ADR3(DLX_EXinst_N63434),
    .O(\DLX_EXinst_Mshift__n0026_Sh<21>/FROM )
  );
  defparam DLX_EXinst_Ker630691.INIT = 16'hCFC0;
  X_LUT4 DLX_EXinst_Ker630691 (
    .ADR0(VCC),
    .ADR1(\DLX_EXinst_Mshift__n0026_Sh[29] ),
    .ADR2(DLX_IDinst_reg_out_B[3]),
    .ADR3(\DLX_EXinst_Mshift__n0026_Sh[21] ),
    .O(\DLX_EXinst_Mshift__n0026_Sh<21>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0026_Sh<21>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0026_Sh<21>/FROM ),
    .O(\DLX_EXinst_Mshift__n0026_Sh[21] )
  );
  X_BUF \DLX_EXinst_Mshift__n0026_Sh<21>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0026_Sh<21>/GROM ),
    .O(DLX_EXinst_N63071)
  );
  defparam DLX_EXlc_md_mda23_a1.INIT = 16'h00AA;
  X_LUT4 DLX_EXlc_md_mda23_a1 (
    .ADR0(DLX_EXlc_md_wint22),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_EXlc_pd_wint5),
    .O(\DLX_EXlc_md_wint23/FROM )
  );
  defparam DLX_EXlc_md_mda8_a1.INIT = 16'h3300;
  X_LUT4 DLX_EXlc_md_mda8_a1 (
    .ADR0(VCC),
    .ADR1(DLX_EXlc_pd_wint5),
    .ADR2(VCC),
    .ADR3(DLX_EXlc_md_wint7),
    .O(\DLX_EXlc_md_wint23/GROM )
  );
  X_BUF \DLX_EXlc_md_wint23/XUSED  (
    .I(\DLX_EXlc_md_wint23/FROM ),
    .O(DLX_EXlc_md_wint23)
  );
  X_BUF \DLX_EXlc_md_wint23/YUSED  (
    .I(\DLX_EXlc_md_wint23/GROM ),
    .O(DLX_EXlc_md_wint8)
  );
  defparam \DLX_EXinst__n0006<28>88 .INIT = 16'h8008;
  X_LUT4 \DLX_EXinst__n0006<28>88  (
    .ADR0(DLX_EXinst_N66105),
    .ADR1(\DLX_IDinst_Imm[31] ),
    .ADR2(N127298),
    .ADR3(DLX_IDinst_IR_opcode_field[1]),
    .O(\CHOICE5201/FROM )
  );
  defparam \DLX_EXinst__n0006<28>99 .INIT = 16'hFFEC;
  X_LUT4 \DLX_EXinst__n0006<28>99  (
    .ADR0(DLX_EXinst__n0077),
    .ADR1(N126636),
    .ADR2(\DLX_IDinst_Imm[12] ),
    .ADR3(CHOICE5201),
    .O(\CHOICE5201/GROM )
  );
  X_BUF \CHOICE5201/XUSED  (
    .I(\CHOICE5201/FROM ),
    .O(CHOICE5201)
  );
  X_BUF \CHOICE5201/YUSED  (
    .I(\CHOICE5201/GROM ),
    .O(CHOICE5203)
  );
  defparam \DLX_EXinst__n0006<3>129 .INIT = 16'hFEFC;
  X_LUT4 \DLX_EXinst__n0006<3>129  (
    .ADR0(N126393),
    .ADR1(CHOICE5046),
    .ADR2(CHOICE5047),
    .ADR3(DLX_EXinst_N66475),
    .O(\CHOICE5049/FROM )
  );
  defparam \DLX_EXinst__n0006<3>160 .INIT = 16'h0F0E;
  X_LUT4 \DLX_EXinst__n0006<3>160  (
    .ADR0(CHOICE5022),
    .ADR1(CHOICE5026),
    .ADR2(DLX_EXinst__n0030),
    .ADR3(CHOICE5049),
    .O(\CHOICE5049/GROM )
  );
  X_BUF \CHOICE5049/XUSED  (
    .I(\CHOICE5049/FROM ),
    .O(CHOICE5049)
  );
  X_BUF \CHOICE5049/YUSED  (
    .I(\CHOICE5049/GROM ),
    .O(CHOICE5051)
  );
  defparam DLX_EXinst_Ker6513856_SW0.INIT = 16'hB830;
  X_LUT4 DLX_EXinst_Ker6513856_SW0 (
    .ADR0(DLX_IDinst_reg_out_B_3_1),
    .ADR1(DLX_IDinst_reg_out_B_2_1),
    .ADR2(DLX_EXinst_N64324),
    .ADR3(DLX_IDinst_reg_out_A[31]),
    .O(\N126006/FROM )
  );
  defparam DLX_EXinst_Ker6513896.INIT = 16'hB080;
  X_LUT4 DLX_EXinst_Ker6513896 (
    .ADR0(DLX_EXinst_N63081),
    .ADR1(DLX_IDinst_reg_out_B_2_1),
    .ADR2(DLX_EXinst_N66494),
    .ADR3(DLX_EXinst_N64324),
    .O(\N126006/GROM )
  );
  X_BUF \N126006/XUSED  (
    .I(\N126006/FROM ),
    .O(N126006)
  );
  X_BUF \N126006/YUSED  (
    .I(\N126006/GROM ),
    .O(CHOICE2971)
  );
  defparam \DLX_EXinst__n0006<3>314 .INIT = 16'hDDDC;
  X_LUT4 \DLX_EXinst__n0006<3>314  (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(CHOICE5085),
    .ADR2(CHOICE5080),
    .ADR3(CHOICE5077),
    .O(\CHOICE5086/FROM )
  );
  defparam \DLX_EXinst__n0006<3>340 .INIT = 16'hF0E0;
  X_LUT4 \DLX_EXinst__n0006<3>340  (
    .ADR0(CHOICE5062),
    .ADR1(CHOICE5058),
    .ADR2(DLX_EXinst__n0030_1),
    .ADR3(CHOICE5086),
    .O(\CHOICE5086/GROM )
  );
  X_BUF \CHOICE5086/XUSED  (
    .I(\CHOICE5086/FROM ),
    .O(CHOICE5086)
  );
  X_BUF \CHOICE5086/YUSED  (
    .I(\CHOICE5086/GROM ),
    .O(CHOICE5088)
  );
  defparam \DLX_EXinst_Mshift__n0026_Sh<22>1 .INIT = 16'hCCF0;
  X_LUT4 \DLX_EXinst_Mshift__n0026_Sh<22>1  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N63066),
    .ADR2(DLX_EXinst_N63434),
    .ADR3(DLX_IDinst_reg_out_B[0]),
    .O(\DLX_EXinst_Mshift__n0026_Sh<22>/FROM )
  );
  defparam DLX_EXinst_Ker64872106.INIT = 16'h3120;
  X_LUT4 DLX_EXinst_Ker64872106 (
    .ADR0(DLX_IDinst_reg_out_B_3_1),
    .ADR1(DLX_IDinst_reg_out_B_2_1),
    .ADR2(\DLX_EXinst_Mshift__n0026_Sh[30] ),
    .ADR3(\DLX_EXinst_Mshift__n0026_Sh[22] ),
    .O(\DLX_EXinst_Mshift__n0026_Sh<22>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0026_Sh<22>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0026_Sh<22>/FROM ),
    .O(\DLX_EXinst_Mshift__n0026_Sh[22] )
  );
  X_BUF \DLX_EXinst_Mshift__n0026_Sh<22>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0026_Sh<22>/GROM ),
    .O(CHOICE3205)
  );
  defparam DLX_IDinst_Ker70070_SW0.INIT = 16'hC0A0;
  X_LUT4 DLX_IDinst_Ker70070_SW0 (
    .ADR0(DLX_IDinst_current_IR[27]),
    .ADR1(DLX_IFinst_IR_latched[27]),
    .ADR2(DLX_IDinst_N70623),
    .ADR3(DLX_EXinst__n0149),
    .O(\N100191/FROM )
  );
  defparam DLX_IDinst_Ker70666115.INIT = 16'h2330;
  X_LUT4 DLX_IDinst_Ker70666115 (
    .ADR0(DLX_IFinst_IR_latched[26]),
    .ADR1(DLX_IFinst_IR_latched[28]),
    .ADR2(DLX_IFinst_IR_latched[30]),
    .ADR3(DLX_IFinst_IR_latched[27]),
    .O(\N100191/GROM )
  );
  X_BUF \N100191/XUSED  (
    .I(\N100191/FROM ),
    .O(N100191)
  );
  X_BUF \N100191/YUSED  (
    .I(\N100191/GROM ),
    .O(CHOICE3283)
  );
  defparam DLX_EXinst_Ker6541425.INIT = 16'h5140;
  X_LUT4 DLX_EXinst_Ker6541425 (
    .ADR0(DLX_IDinst_IR_function_field_3_1),
    .ADR1(DLX_IDinst_IR_function_field[0]),
    .ADR2(DLX_EXinst_N62806),
    .ADR3(DLX_EXinst_N63474),
    .O(\CHOICE1337/FROM )
  );
  defparam DLX_EXinst_Ker6541428.INIT = 16'hFFF0;
  X_LUT4 DLX_EXinst_Ker6541428 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(CHOICE1331),
    .ADR3(CHOICE1337),
    .O(\CHOICE1337/GROM )
  );
  X_BUF \CHOICE1337/XUSED  (
    .I(\CHOICE1337/FROM ),
    .O(CHOICE1337)
  );
  X_BUF \CHOICE1337/YUSED  (
    .I(\CHOICE1337/GROM ),
    .O(N97960)
  );
  defparam DLX_EXinst_Ker6513899.INIT = 16'hFF88;
  X_LUT4 DLX_EXinst_Ker6513899 (
    .ADR0(N111221),
    .ADR1(CHOICE2965),
    .ADR2(VCC),
    .ADR3(CHOICE2971),
    .O(\N107444/FROM )
  );
  defparam \DLX_EXinst__n0006<3>310 .INIT = 16'hECA0;
  X_LUT4 \DLX_EXinst__n0006<3>310  (
    .ADR0(N101725),
    .ADR1(DLX_IDinst_reg_out_B[4]),
    .ADR2(DLX_EXinst_ALU_result[3]),
    .ADR3(N107444),
    .O(\N107444/GROM )
  );
  X_BUF \N107444/XUSED  (
    .I(\N107444/FROM ),
    .O(N107444)
  );
  X_BUF \N107444/YUSED  (
    .I(\N107444/GROM ),
    .O(CHOICE5085)
  );
  defparam DLX_EXinst_Ker66070.INIT = 16'h0010;
  X_LUT4 DLX_EXinst_Ker66070 (
    .ADR0(N90062),
    .ADR1(DLX_IDinst_reg_out_B_3_1),
    .ADR2(DLX_EXinst_N66226),
    .ADR3(DLX_IDinst_reg_out_B[4]),
    .O(\DLX_EXinst_N66072/FROM )
  );
  defparam DLX_EXinst_Ker6516811.INIT = 16'hD800;
  X_LUT4 DLX_EXinst_Ker6516811 (
    .ADR0(DLX_IDinst_reg_out_B_3_1),
    .ADR1(DLX_EXinst_N62876),
    .ADR2(DLX_EXinst_N62896),
    .ADR3(DLX_IDinst_reg_out_B[0]),
    .O(\DLX_EXinst_N66072/GROM )
  );
  X_BUF \DLX_EXinst_N66072/XUSED  (
    .I(\DLX_EXinst_N66072/FROM ),
    .O(DLX_EXinst_N66072)
  );
  X_BUF \DLX_EXinst_N66072/YUSED  (
    .I(\DLX_EXinst_N66072/GROM ),
    .O(CHOICE1174)
  );
  defparam \DLX_EXinst__n0006<14>15_SW0 .INIT = 16'h0303;
  X_LUT4 \DLX_EXinst__n0006<14>15_SW0  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_IR_opcode_field[0]),
    .ADR2(DLX_IDinst_reg_out_A[14]),
    .ADR3(VCC),
    .O(\N127350/FROM )
  );
  defparam \DLX_EXinst__n0006<8>16_SW0 .INIT = 16'h0303;
  X_LUT4 \DLX_EXinst__n0006<8>16_SW0  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_IR_opcode_field[0]),
    .ADR2(DLX_IDinst_reg_out_A[8]),
    .ADR3(VCC),
    .O(\N127350/GROM )
  );
  X_BUF \N127350/XUSED  (
    .I(\N127350/FROM ),
    .O(N127350)
  );
  X_BUF \N127350/YUSED  (
    .I(\N127350/GROM ),
    .O(N127302)
  );
  defparam DLX_EXlc_md_mda22_a1.INIT = 16'h3030;
  X_LUT4 DLX_EXlc_md_mda22_a1 (
    .ADR0(VCC),
    .ADR1(DLX_EXlc_pd_wint5),
    .ADR2(DLX_EXlc_md_wint21),
    .ADR3(VCC),
    .O(\DLX_EXlc_md_wint22/FROM )
  );
  defparam DLX_EXlc_md_mda9_a1.INIT = 16'h0F00;
  X_LUT4 DLX_EXlc_md_mda9_a1 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_EXlc_pd_wint5),
    .ADR3(DLX_EXlc_md_wint8),
    .O(\DLX_EXlc_md_wint22/GROM )
  );
  X_BUF \DLX_EXlc_md_wint22/XUSED  (
    .I(\DLX_EXlc_md_wint22/FROM ),
    .O(DLX_EXlc_md_wint22)
  );
  X_BUF \DLX_EXlc_md_wint22/YUSED  (
    .I(\DLX_EXlc_md_wint22/GROM ),
    .O(DLX_EXlc_md_wint9)
  );
  defparam \DLX_EXinst__n0006<29>88 .INIT = 16'h8040;
  X_LUT4 \DLX_EXinst__n0006<29>88  (
    .ADR0(DLX_IDinst_IR_opcode_field[1]),
    .ADR1(DLX_EXinst_N66105),
    .ADR2(\DLX_IDinst_Imm[31] ),
    .ADR3(N127374),
    .O(\CHOICE5353/FROM )
  );
  defparam \DLX_EXinst__n0006<29>99 .INIT = 16'hFFEA;
  X_LUT4 \DLX_EXinst__n0006<29>99  (
    .ADR0(N126486),
    .ADR1(DLX_EXinst__n0077),
    .ADR2(\DLX_IDinst_Imm[13] ),
    .ADR3(CHOICE5353),
    .O(\CHOICE5353/GROM )
  );
  X_BUF \CHOICE5353/XUSED  (
    .I(\CHOICE5353/FROM ),
    .O(CHOICE5353)
  );
  X_BUF \CHOICE5353/YUSED  (
    .I(\CHOICE5353/GROM ),
    .O(CHOICE5355)
  );
  defparam \DLX_EXinst__n0006<3>352 .INIT = 16'hEEAA;
  X_LUT4 \DLX_EXinst__n0006<3>352  (
    .ADR0(CHOICE5088),
    .ADR1(DLX_EXinst__n0016[3]),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N63836),
    .O(\DLX_EXinst_ALU_result<3>/FROM )
  );
  defparam \DLX_EXinst__n0006<3>393 .INIT = 16'hFCEC;
  X_LUT4 \DLX_EXinst__n0006<3>393  (
    .ADR0(CHOICE5051),
    .ADR1(DLX_EXinst_N63689),
    .ADR2(DLX_EXinst__n0149),
    .ADR3(CHOICE5089),
    .O(\DLX_EXinst_ALU_result<3>/GROM )
  );
  X_BUF \DLX_EXinst_ALU_result<3>/XUSED  (
    .I(\DLX_EXinst_ALU_result<3>/FROM ),
    .O(CHOICE5089)
  );
  X_BUF \DLX_EXinst_ALU_result<3>/YUSED  (
    .I(\DLX_EXinst_ALU_result<3>/GROM ),
    .O(N120114)
  );
  defparam vga_top_vga1__n00084.INIT = 16'h8000;
  X_LUT4 vga_top_vga1__n00084 (
    .ADR0(vga_top_vga1_hcounter[7]),
    .ADR1(vga_top_vga1_hcounter[5]),
    .ADR2(vga_top_vga1_hcounter[1]),
    .ADR3(vga_top_vga1_hcounter[4]),
    .O(\CHOICE3214/FROM )
  );
  defparam vga_top_vga1__n00131.INIT = 16'h8080;
  X_LUT4 vga_top_vga1__n00131 (
    .ADR0(vga_top_vga1__n0037),
    .ADR1(vga_top_vga1_hcounter[0]),
    .ADR2(vga_top_vga1_hcounter[1]),
    .ADR3(VCC),
    .O(\CHOICE3214/GROM )
  );
  X_BUF \CHOICE3214/XUSED  (
    .I(\CHOICE3214/FROM ),
    .O(CHOICE3214)
  );
  X_BUF \CHOICE3214/YUSED  (
    .I(\CHOICE3214/GROM ),
    .O(vga_top_vga1__n0013)
  );
  defparam \DLX_EXinst__n0006<3>178 .INIT = 16'hEECC;
  X_LUT4 \DLX_EXinst__n0006<3>178  (
    .ADR0(DLX_IDinst_reg_out_B[3]),
    .ADR1(DLX_EXinst_N64448),
    .ADR2(VCC),
    .ADR3(DLX_EXinst__n0045),
    .O(\CHOICE5056/FROM )
  );
  defparam \DLX_EXinst__n0006<3>187 .INIT = 16'hCC08;
  X_LUT4 \DLX_EXinst__n0006<3>187  (
    .ADR0(DLX_EXinst__n0047),
    .ADR1(DLX_IDinst_reg_out_A[3]),
    .ADR2(DLX_IDinst_reg_out_B[3]),
    .ADR3(CHOICE5056),
    .O(\CHOICE5056/GROM )
  );
  X_BUF \CHOICE5056/XUSED  (
    .I(\CHOICE5056/FROM ),
    .O(CHOICE5056)
  );
  X_BUF \CHOICE5056/YUSED  (
    .I(\CHOICE5056/GROM ),
    .O(CHOICE5058)
  );
  defparam DLX_IDinst_Ker70666139.INIT = 16'h0032;
  X_LUT4 DLX_IDinst_Ker70666139 (
    .ADR0(CHOICE3283),
    .ADR1(DLX_IFinst_IR_latched[29]),
    .ADR2(CHOICE3275),
    .ADR3(DLX_IFinst_IR_latched[31]),
    .O(\N109350/FROM )
  );
  defparam \DLX_IDinst_slot_num_FFd2-In48 .INIT = 16'hA000;
  X_LUT4 \DLX_IDinst_slot_num_FFd2-In48  (
    .ADR0(DLX_IDinst_slot_num_FFd2),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_delay_slot),
    .ADR3(N109350),
    .O(\N109350/GROM )
  );
  X_BUF \N109350/XUSED  (
    .I(\N109350/FROM ),
    .O(N109350)
  );
  X_BUF \N109350/YUSED  (
    .I(\N109350/GROM ),
    .O(CHOICE2525)
  );
  defparam \DLX_EXinst_Mshift__n0026_Sh<16>1 .INIT = 16'hEE22;
  X_LUT4 \DLX_EXinst_Mshift__n0026_Sh<16>1  (
    .ADR0(DLX_EXinst_N63419),
    .ADR1(DLX_IDinst_reg_out_B[0]),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N63051),
    .O(\DLX_EXinst_Mshift__n0026_Sh<16>/FROM )
  );
  defparam DLX_EXinst_Ker648021.INIT = 16'hEE22;
  X_LUT4 DLX_EXinst_Ker648021 (
    .ADR0(\DLX_EXinst_Mshift__n0023_Sh[8] ),
    .ADR1(DLX_IDinst_reg_out_B_3_1),
    .ADR2(VCC),
    .ADR3(\DLX_EXinst_Mshift__n0026_Sh[16] ),
    .O(\DLX_EXinst_Mshift__n0026_Sh<16>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0026_Sh<16>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0026_Sh<16>/FROM ),
    .O(\DLX_EXinst_Mshift__n0026_Sh[16] )
  );
  X_BUF \DLX_EXinst_Mshift__n0026_Sh<16>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0026_Sh<16>/GROM ),
    .O(DLX_EXinst_N64804)
  );
  defparam \DLX_EXinst__n0006<4>123 .INIT = 16'hFAAA;
  X_LUT4 \DLX_EXinst__n0006<4>123  (
    .ADR0(DLX_EXinst__n0046),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[4]),
    .ADR3(DLX_EXinst__n0045),
    .O(\CHOICE4003/FROM )
  );
  defparam \DLX_EXinst__n0006<4>125 .INIT = 16'hFF20;
  X_LUT4 \DLX_EXinst__n0006<4>125  (
    .ADR0(\DLX_EXinst_Mshift__n0026_Sh[52] ),
    .ADR1(N110935),
    .ADR2(DLX_EXinst__n0049),
    .ADR3(CHOICE4003),
    .O(\CHOICE4003/GROM )
  );
  X_BUF \CHOICE4003/XUSED  (
    .I(\CHOICE4003/FROM ),
    .O(CHOICE4003)
  );
  X_BUF \CHOICE4003/YUSED  (
    .I(\CHOICE4003/GROM ),
    .O(CHOICE4004)
  );
  defparam \DLX_EXinst_Mshift__n0028_Sh<57>1 .INIT = 16'h3022;
  X_LUT4 \DLX_EXinst_Mshift__n0028_Sh<57>1  (
    .ADR0(\DLX_EXinst_Mshift__n0024_Sh[25] ),
    .ADR1(DLX_IDinst_IR_function_field_3_1),
    .ADR2(\DLX_EXinst_Mshift__n0028_Sh[29] ),
    .ADR3(DLX_IDinst_IR_function_field_2_1),
    .O(\DLX_EXinst_Mshift__n0028_Sh<57>/FROM )
  );
  defparam DLX_EXinst_Ker6514897.INIT = 16'h2F20;
  X_LUT4 DLX_EXinst_Ker6514897 (
    .ADR0(\DLX_EXinst_Mshift__n0024_Sh[25] ),
    .ADR1(DLX_IDinst_IR_function_field_3_1),
    .ADR2(DLX_IDinst_IR_function_field_2_1),
    .ADR3(DLX_EXinst_N63021),
    .O(\DLX_EXinst_Mshift__n0028_Sh<57>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0028_Sh<57>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0028_Sh<57>/FROM ),
    .O(\DLX_EXinst_Mshift__n0028_Sh[57] )
  );
  X_BUF \DLX_EXinst_Mshift__n0028_Sh<57>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0028_Sh<57>/GROM ),
    .O(CHOICE3104)
  );
  defparam DLX_EXinst_Ker6516825.INIT = 16'h00AC;
  X_LUT4 DLX_EXinst_Ker6516825 (
    .ADR0(DLX_EXinst_N63379),
    .ADR1(DLX_EXinst_N63274),
    .ADR2(DLX_IDinst_reg_out_B_3_1),
    .ADR3(DLX_IDinst_reg_out_B[0]),
    .O(\CHOICE1180/FROM )
  );
  defparam DLX_EXinst_Ker6516828.INIT = 16'hFFCC;
  X_LUT4 DLX_EXinst_Ker6516828 (
    .ADR0(VCC),
    .ADR1(CHOICE1174),
    .ADR2(VCC),
    .ADR3(CHOICE1180),
    .O(\CHOICE1180/GROM )
  );
  X_BUF \CHOICE1180/XUSED  (
    .I(\CHOICE1180/FROM ),
    .O(CHOICE1180)
  );
  X_BUF \CHOICE1180/YUSED  (
    .I(\CHOICE1180/GROM ),
    .O(N97017)
  );
  defparam DLX_IDinst_Ker697091.INIT = 16'hFF57;
  X_LUT4 DLX_IDinst_Ker697091 (
    .ADR0(DLX_IDinst__n0387),
    .ADR1(DLX_IDinst_N70006),
    .ADR2(DLX_IDinst_N70918),
    .ADR3(DLX_IDinst__n0331),
    .O(\DLX_IDinst_reg_out_B<0>/FROM )
  );
  defparam \DLX_IDinst__n0118<0>1 .INIT = 16'hF000;
  X_LUT4 \DLX_IDinst__n0118<0>1  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_regB_eff[0]),
    .ADR3(DLX_IDinst_N69711),
    .O(DLX_IDinst__n0118[0])
  );
  X_BUF \DLX_IDinst_reg_out_B<0>/XUSED  (
    .I(\DLX_IDinst_reg_out_B<0>/FROM ),
    .O(DLX_IDinst_N69711)
  );
  defparam \DLX_EXinst_Mshift__n0025_Sh<2>_SW0 .INIT = 16'h4477;
  X_LUT4 \DLX_EXinst_Mshift__n0025_Sh<2>_SW0  (
    .ADR0(DLX_IDinst_reg_out_A[0]),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[2]),
    .O(\N94921/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0025_Sh<2> .INIT = 16'h085D;
  X_LUT4 \DLX_EXinst_Mshift__n0025_Sh<2>  (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(DLX_IDinst_reg_out_A[1]),
    .ADR2(DLX_IDinst_reg_out_B[1]),
    .ADR3(N94921),
    .O(\N94921/GROM )
  );
  X_BUF \N94921/XUSED  (
    .I(\N94921/FROM ),
    .O(N94921)
  );
  X_BUF \N94921/YUSED  (
    .I(\N94921/GROM ),
    .O(\DLX_EXinst_Mshift__n0025_Sh[2] )
  );
  defparam \DLX_EXinst__n0006<5>194 .INIT = 16'h2020;
  X_LUT4 \DLX_EXinst__n0006<5>194  (
    .ADR0(DLX_EXinst_N66226),
    .ADR1(DLX_IDinst_reg_out_B[3]),
    .ADR2(DLX_EXinst_N62906),
    .ADR3(VCC),
    .O(\CHOICE4464/FROM )
  );
  defparam \DLX_EXinst__n0006<3>277 .INIT = 16'h0400;
  X_LUT4 \DLX_EXinst__n0006<3>277  (
    .ADR0(DLX_IDinst_reg_out_B[2]),
    .ADR1(\DLX_EXinst_Mshift__n0025_Sh[3] ),
    .ADR2(DLX_IDinst_reg_out_B[3]),
    .ADR3(DLX_EXinst_N66226),
    .O(\CHOICE4464/GROM )
  );
  X_BUF \CHOICE4464/XUSED  (
    .I(\CHOICE4464/FROM ),
    .O(CHOICE4464)
  );
  X_BUF \CHOICE4464/YUSED  (
    .I(\CHOICE4464/GROM ),
    .O(CHOICE5080)
  );
  defparam \DLX_EXinst__n0006<7>199 .INIT = 16'h8C88;
  X_LUT4 \DLX_EXinst__n0006<7>199  (
    .ADR0(DLX_EXinst__n0046),
    .ADR1(DLX_IDinst_reg_out_B[7]),
    .ADR2(DLX_IDinst_reg_out_A[7]),
    .ADR3(DLX_EXinst__n0047),
    .O(\CHOICE3844/FROM )
  );
  defparam \DLX_EXinst__n0006<4>119 .INIT = 16'h8F88;
  X_LUT4 \DLX_EXinst__n0006<4>119  (
    .ADR0(N111221),
    .ADR1(DLX_EXinst_N64500),
    .ADR2(DLX_IDinst_reg_out_A[4]),
    .ADR3(DLX_EXinst__n0047),
    .O(\CHOICE3844/GROM )
  );
  X_BUF \CHOICE3844/XUSED  (
    .I(\CHOICE3844/FROM ),
    .O(CHOICE3844)
  );
  X_BUF \CHOICE3844/YUSED  (
    .I(\CHOICE3844/GROM ),
    .O(CHOICE4000)
  );
  defparam \DLX_EXinst__n0006<17>199 .INIT = 16'hF040;
  X_LUT4 \DLX_EXinst__n0006<17>199  (
    .ADR0(DLX_IDinst_reg_out_A[17]),
    .ADR1(DLX_EXinst__n0047),
    .ADR2(DLX_IDinst_reg_out_B[17]),
    .ADR3(DLX_EXinst__n0046),
    .O(\CHOICE5613/FROM )
  );
  defparam \DLX_EXinst__n0006<3>199 .INIT = 16'hA0A8;
  X_LUT4 \DLX_EXinst__n0006<3>199  (
    .ADR0(DLX_IDinst_reg_out_B[3]),
    .ADR1(DLX_EXinst__n0047),
    .ADR2(DLX_EXinst__n0046),
    .ADR3(DLX_IDinst_reg_out_A[3]),
    .O(\CHOICE5613/GROM )
  );
  X_BUF \CHOICE5613/XUSED  (
    .I(\CHOICE5613/FROM ),
    .O(CHOICE5613)
  );
  X_BUF \CHOICE5613/YUSED  (
    .I(\CHOICE5613/GROM ),
    .O(CHOICE5062)
  );
  defparam DLX_EXinst_Ker6540926.INIT = 16'h5140;
  X_LUT4 DLX_EXinst_Ker6540926 (
    .ADR0(DLX_IDinst_IR_function_field_3_1),
    .ADR1(DLX_IDinst_IR_function_field[0]),
    .ADR2(DLX_EXinst_N63474),
    .ADR3(DLX_EXinst_N62811),
    .O(\CHOICE1288/FROM )
  );
  defparam DLX_EXinst_Ker6540928.INIT = 16'hFFF0;
  X_LUT4 DLX_EXinst_Ker6540928 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(CHOICE1282),
    .ADR3(CHOICE1288),
    .O(\CHOICE1288/GROM )
  );
  X_BUF \CHOICE1288/XUSED  (
    .I(\CHOICE1288/FROM ),
    .O(CHOICE1288)
  );
  X_BUF \CHOICE1288/YUSED  (
    .I(\CHOICE1288/GROM ),
    .O(N97665)
  );
  defparam DLX_EXinst_Ker6630711.INIT = 16'h4000;
  X_LUT4 DLX_EXinst_Ker6630711 (
    .ADR0(DLX_IDinst_IR_function_field[5]),
    .ADR1(DLX_EXinst_N66096),
    .ADR2(DLX_IDinst_IR_function_field_1_1),
    .ADR3(DLX_IDinst_IR_function_field[0]),
    .O(\CHOICE3564/FROM )
  );
  defparam DLX_EXinst_Ker66307161.INIT = 16'h0100;
  X_LUT4 DLX_EXinst_Ker66307161 (
    .ADR0(DLX_IDinst_reg_out_B[31]),
    .ADR1(N126424),
    .ADR2(DLX_IDinst_reg_out_B[30]),
    .ADR3(CHOICE3564),
    .O(\CHOICE3564/GROM )
  );
  X_BUF \CHOICE3564/XUSED  (
    .I(\CHOICE3564/FROM ),
    .O(CHOICE3564)
  );
  X_BUF \CHOICE3564/YUSED  (
    .I(\CHOICE3564/GROM ),
    .O(N111221)
  );
  defparam \DLX_EXinst_Mshift__n0027_Sh<44>25 .INIT = 16'h3202;
  X_LUT4 \DLX_EXinst_Mshift__n0027_Sh<44>25  (
    .ADR0(\DLX_EXinst_Mshift__n0027_Sh[12] ),
    .ADR1(DLX_IDinst_IR_function_field_3_1),
    .ADR2(DLX_IDinst_IR_function_field_2_1),
    .ADR3(\DLX_EXinst_Mshift__n0027_Sh[8] ),
    .O(\CHOICE1048/FROM )
  );
  defparam \DLX_EXinst__n0006<12>41 .INIT = 16'h0A08;
  X_LUT4 \DLX_EXinst__n0006<12>41  (
    .ADR0(DLX_EXinst__n0081),
    .ADR1(CHOICE1042),
    .ADR2(N109130),
    .ADR3(CHOICE1048),
    .O(\CHOICE1048/GROM )
  );
  X_BUF \CHOICE1048/XUSED  (
    .I(\CHOICE1048/FROM ),
    .O(CHOICE1048)
  );
  X_BUF \CHOICE1048/YUSED  (
    .I(\CHOICE1048/GROM ),
    .O(CHOICE3870)
  );
  defparam \DLX_EXinst__n0006<4>252 .INIT = 16'hF888;
  X_LUT4 \DLX_EXinst__n0006<4>252  (
    .ADR0(DLX_EXinst__n0030_1),
    .ADR1(CHOICE4023),
    .ADR2(DLX_EXinst__n0016[4]),
    .ADR3(DLX_EXinst_N63836),
    .O(\DLX_EXinst_ALU_result<4>/FROM )
  );
  defparam \DLX_EXinst__n0006<4>291 .INIT = 16'hFCEC;
  X_LUT4 \DLX_EXinst__n0006<4>291  (
    .ADR0(CHOICE3994),
    .ADR1(DLX_EXinst_N63689),
    .ADR2(DLX_EXinst__n0149),
    .ADR3(CHOICE4025),
    .O(\DLX_EXinst_ALU_result<4>/GROM )
  );
  X_BUF \DLX_EXinst_ALU_result<4>/XUSED  (
    .I(\DLX_EXinst_ALU_result<4>/FROM ),
    .O(CHOICE4025)
  );
  X_BUF \DLX_EXinst_ALU_result<4>/YUSED  (
    .I(\DLX_EXinst_ALU_result<4>/GROM ),
    .O(N113660)
  );
  defparam \DLX_EXinst__n0006<4>180 .INIT = 16'hEAEA;
  X_LUT4 \DLX_EXinst__n0006<4>180  (
    .ADR0(CHOICE4016),
    .ADR1(DLX_EXinst__n0047),
    .ADR2(DLX_IDinst_reg_out_A[4]),
    .ADR3(VCC),
    .O(\CHOICE4017/FROM )
  );
  defparam \DLX_EXinst__n0006<4>189 .INIT = 16'hFF20;
  X_LUT4 \DLX_EXinst__n0006<4>189  (
    .ADR0(DLX_EXinst_N62901),
    .ADR1(DLX_IDinst_reg_out_B[3]),
    .ADR2(DLX_EXinst_N66226),
    .ADR3(CHOICE4017),
    .O(\CHOICE4017/GROM )
  );
  X_BUF \CHOICE4017/XUSED  (
    .I(\CHOICE4017/FROM ),
    .O(CHOICE4017)
  );
  X_BUF \CHOICE4017/YUSED  (
    .I(\CHOICE4017/GROM ),
    .O(CHOICE4018)
  );
  defparam \DLX_EXinst__n0006<28>271 .INIT = 16'hFFA0;
  X_LUT4 \DLX_EXinst__n0006<28>271  (
    .ADR0(DLX_IDinst_reg_out_B[28]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst__n0045),
    .ADR3(DLX_EXinst_N64448),
    .O(\CHOICE5236/FROM )
  );
  defparam DLX_EXinst_Ker6630731.INIT = 16'h0001;
  X_LUT4 DLX_EXinst_Ker6630731 (
    .ADR0(DLX_IDinst_reg_out_B[28]),
    .ADR1(DLX_IDinst_reg_out_B[26]),
    .ADR2(DLX_IDinst_reg_out_B[27]),
    .ADR3(DLX_IDinst_reg_out_B[29]),
    .O(\CHOICE5236/GROM )
  );
  X_BUF \CHOICE5236/XUSED  (
    .I(\CHOICE5236/FROM ),
    .O(CHOICE5236)
  );
  X_BUF \CHOICE5236/YUSED  (
    .I(\CHOICE5236/GROM ),
    .O(CHOICE3572)
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<30>1 .INIT = 16'h4F40;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<30>1  (
    .ADR0(DLX_opcode_of_WB[2]),
    .ADR1(DLX_IDinst_Mmux__n0148__net123),
    .ADR2(DLX_IDinst__n0147),
    .ADR3(DLX_MEMinst_RF_data_in[30]),
    .O(\DLX_IDinst_WB_data_eff<30>/FROM )
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<20>1 .INIT = 16'h30AA;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<20>1  (
    .ADR0(DLX_MEMinst_RF_data_in[20]),
    .ADR1(DLX_opcode_of_WB[2]),
    .ADR2(DLX_IDinst_Mmux__n0148__net123),
    .ADR3(DLX_IDinst__n0147),
    .O(\DLX_IDinst_WB_data_eff<30>/GROM )
  );
  X_BUF \DLX_IDinst_WB_data_eff<30>/XUSED  (
    .I(\DLX_IDinst_WB_data_eff<30>/FROM ),
    .O(DLX_IDinst_WB_data_eff[30])
  );
  X_BUF \DLX_IDinst_WB_data_eff<30>/YUSED  (
    .I(\DLX_IDinst_WB_data_eff<30>/GROM ),
    .O(DLX_IDinst_WB_data_eff[20])
  );
  defparam vga_top_vga1__n00098.INIT = 16'hFFFC;
  X_LUT4 vga_top_vga1__n00098 (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_vcounter[0]),
    .ADR2(vga_top_vga1_vcounter[1]),
    .ADR3(vga_top_vga1_vcounter[8]),
    .O(\CHOICE3415/FROM )
  );
  defparam vga_top_vga1__n000910.INIT = 16'hFFFC;
  X_LUT4 vga_top_vga1__n000910 (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_vcounter[7]),
    .ADR2(vga_top_vga1_vcounter[6]),
    .ADR3(CHOICE3415),
    .O(\CHOICE3415/GROM )
  );
  X_BUF \CHOICE3415/XUSED  (
    .I(\CHOICE3415/FROM ),
    .O(CHOICE3415)
  );
  X_BUF \CHOICE3415/YUSED  (
    .I(\CHOICE3415/GROM ),
    .O(CHOICE3416)
  );
  defparam \DLX_EXinst_Mshift__n0026_Sh<24>_SW0 .INIT = 16'hDD88;
  X_LUT4 \DLX_EXinst_Mshift__n0026_Sh<24>_SW0  (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(DLX_IDinst_reg_out_A[27]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[25]),
    .O(\N94107/FROM )
  );
  defparam DLX_EXinst_Ker6458015.INIT = 16'h0D08;
  X_LUT4 DLX_EXinst_Ker6458015 (
    .ADR0(DLX_IDinst_IR_function_field_1_1),
    .ADR1(DLX_IDinst_reg_out_A[25]),
    .ADR2(DLX_IDinst_IR_function_field[0]),
    .ADR3(DLX_IDinst_reg_out_A[27]),
    .O(\N94107/GROM )
  );
  X_BUF \N94107/XUSED  (
    .I(\N94107/FROM ),
    .O(N94107)
  );
  X_BUF \N94107/YUSED  (
    .I(\N94107/GROM ),
    .O(CHOICE1838)
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<28>1 .INIT = 16'h5D08;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<28>1  (
    .ADR0(DLX_IDinst__n0147),
    .ADR1(DLX_IDinst_Mmux__n0148__net123),
    .ADR2(DLX_opcode_of_WB[2]),
    .ADR3(DLX_MEMinst_RF_data_in[28]),
    .O(\DLX_IDinst_WB_data_eff<28>/FROM )
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<21>1 .INIT = 16'h0CAA;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<21>1  (
    .ADR0(DLX_MEMinst_RF_data_in[21]),
    .ADR1(DLX_IDinst_Mmux__n0148__net123),
    .ADR2(DLX_opcode_of_WB[2]),
    .ADR3(DLX_IDinst__n0147),
    .O(\DLX_IDinst_WB_data_eff<28>/GROM )
  );
  X_BUF \DLX_IDinst_WB_data_eff<28>/XUSED  (
    .I(\DLX_IDinst_WB_data_eff<28>/FROM ),
    .O(DLX_IDinst_WB_data_eff[28])
  );
  X_BUF \DLX_IDinst_WB_data_eff<28>/YUSED  (
    .I(\DLX_IDinst_WB_data_eff<28>/GROM ),
    .O(DLX_IDinst_WB_data_eff[21])
  );
  defparam \DLX_EXinst__n0006<23>152 .INIT = 16'h88A8;
  X_LUT4 \DLX_EXinst__n0006<23>152  (
    .ADR0(DLX_IDinst_reg_out_B[23]),
    .ADR1(DLX_EXinst__n0046),
    .ADR2(DLX_EXinst__n0047),
    .ADR3(DLX_IDinst_reg_out_A[23]),
    .O(\CHOICE4064/FROM )
  );
  defparam DLX_EXinst_Ker6630744.INIT = 16'h0001;
  X_LUT4 DLX_EXinst_Ker6630744 (
    .ADR0(DLX_IDinst_reg_out_B[25]),
    .ADR1(DLX_IDinst_reg_out_B[22]),
    .ADR2(DLX_IDinst_reg_out_B[24]),
    .ADR3(DLX_IDinst_reg_out_B[23]),
    .O(\CHOICE4064/GROM )
  );
  X_BUF \CHOICE4064/XUSED  (
    .I(\CHOICE4064/FROM ),
    .O(CHOICE4064)
  );
  X_BUF \CHOICE4064/YUSED  (
    .I(\CHOICE4064/GROM ),
    .O(CHOICE3579)
  );
  defparam DLX_EXinst_Ker6615544.INIT = 16'hAA80;
  X_LUT4 DLX_EXinst_Ker6615544 (
    .ADR0(N110065),
    .ADR1(CHOICE1321),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(CHOICE1324),
    .O(\N97892/FROM )
  );
  defparam \DLX_EXinst__n0006<4>57_SW0 .INIT = 16'hFFEC;
  X_LUT4 \DLX_EXinst__n0006<4>57_SW0  (
    .ADR0(\DLX_EXinst_Mshift__n0028_Sh[52] ),
    .ADR1(DLX_EXinst__n0079),
    .ADR2(DLX_EXinst_N66507),
    .ADR3(N97892),
    .O(\N97892/GROM )
  );
  X_BUF \N97892/XUSED  (
    .I(\N97892/FROM ),
    .O(N97892)
  );
  X_BUF \N97892/YUSED  (
    .I(\N97892/GROM ),
    .O(N126038)
  );
  defparam \DLX_EXinst__n0006<5>124 .INIT = 16'hEECC;
  X_LUT4 \DLX_EXinst__n0006<5>124  (
    .ADR0(DLX_IDinst_reg_out_B[5]),
    .ADR1(DLX_EXinst_N64448),
    .ADR2(VCC),
    .ADR3(DLX_EXinst__n0045),
    .O(\CHOICE4446/FROM )
  );
  defparam \DLX_EXinst__n0006<5>133 .INIT = 16'hF020;
  X_LUT4 \DLX_EXinst__n0006<5>133  (
    .ADR0(DLX_EXinst__n0047),
    .ADR1(DLX_IDinst_reg_out_B[5]),
    .ADR2(DLX_IDinst_reg_out_A[5]),
    .ADR3(CHOICE4446),
    .O(\CHOICE4446/GROM )
  );
  X_BUF \CHOICE4446/XUSED  (
    .I(\CHOICE4446/FROM ),
    .O(CHOICE4446)
  );
  X_BUF \CHOICE4446/YUSED  (
    .I(\CHOICE4446/GROM ),
    .O(CHOICE4448)
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<27>1 .INIT = 16'h30AA;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<27>1  (
    .ADR0(DLX_MEMinst_RF_data_in[27]),
    .ADR1(DLX_opcode_of_WB[2]),
    .ADR2(DLX_IDinst_Mmux__n0148__net123),
    .ADR3(DLX_IDinst__n0147),
    .O(\DLX_IDinst_WB_data_eff<27>/FROM )
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<22>1 .INIT = 16'h7520;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<22>1  (
    .ADR0(DLX_IDinst__n0147),
    .ADR1(DLX_opcode_of_WB[2]),
    .ADR2(DLX_IDinst_Mmux__n0148__net123),
    .ADR3(DLX_MEMinst_RF_data_in[22]),
    .O(\DLX_IDinst_WB_data_eff<27>/GROM )
  );
  X_BUF \DLX_IDinst_WB_data_eff<27>/XUSED  (
    .I(\DLX_IDinst_WB_data_eff<27>/FROM ),
    .O(DLX_IDinst_WB_data_eff[27])
  );
  X_BUF \DLX_IDinst_WB_data_eff<27>/YUSED  (
    .I(\DLX_IDinst_WB_data_eff<27>/GROM ),
    .O(DLX_IDinst_WB_data_eff[22])
  );
  defparam DLX_EXinst__n003538.INIT = 16'hFFFE;
  X_LUT4 DLX_EXinst__n003538 (
    .ADR0(DLX_IDinst_reg_out_B[17]),
    .ADR1(DLX_IDinst_reg_out_B[18]),
    .ADR2(DLX_IDinst_reg_out_B[16]),
    .ADR3(DLX_IDinst_reg_out_B[19]),
    .O(\CHOICE3547/FROM )
  );
  defparam DLX_EXinst_Ker6630783.INIT = 16'h0001;
  X_LUT4 DLX_EXinst_Ker6630783 (
    .ADR0(DLX_IDinst_reg_out_B[19]),
    .ADR1(DLX_IDinst_reg_out_B[21]),
    .ADR2(DLX_IDinst_reg_out_B[20]),
    .ADR3(DLX_IDinst_reg_out_B[18]),
    .O(\CHOICE3547/GROM )
  );
  X_BUF \CHOICE3547/XUSED  (
    .I(\CHOICE3547/FROM ),
    .O(CHOICE3547)
  );
  X_BUF \CHOICE3547/YUSED  (
    .I(\CHOICE3547/GROM ),
    .O(CHOICE3588)
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<26>1 .INIT = 16'h50D8;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<26>1  (
    .ADR0(DLX_IDinst__n0147),
    .ADR1(DLX_IDinst_Mmux__n0148__net123),
    .ADR2(DLX_MEMinst_RF_data_in[26]),
    .ADR3(DLX_opcode_of_WB[2]),
    .O(\DLX_IDinst_WB_data_eff<26>/FROM )
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<23>1 .INIT = 16'h0CAA;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<23>1  (
    .ADR0(DLX_MEMinst_RF_data_in[23]),
    .ADR1(DLX_IDinst_Mmux__n0148__net123),
    .ADR2(DLX_opcode_of_WB[2]),
    .ADR3(DLX_IDinst__n0147),
    .O(\DLX_IDinst_WB_data_eff<26>/GROM )
  );
  X_BUF \DLX_IDinst_WB_data_eff<26>/XUSED  (
    .I(\DLX_IDinst_WB_data_eff<26>/FROM ),
    .O(DLX_IDinst_WB_data_eff[26])
  );
  X_BUF \DLX_IDinst_WB_data_eff<26>/YUSED  (
    .I(\DLX_IDinst_WB_data_eff<26>/GROM ),
    .O(DLX_IDinst_WB_data_eff[23])
  );
  defparam \DLX_EXinst__n0006<5>252 .INIT = 16'hECA0;
  X_LUT4 \DLX_EXinst__n0006<5>252  (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(DLX_EXinst_ALU_result[5]),
    .ADR2(N108433),
    .ADR3(N101725),
    .O(\CHOICE4475/FROM )
  );
  defparam \DLX_EXinst__n0006<5>276_SW0 .INIT = 16'hFF50;
  X_LUT4 \DLX_EXinst__n0006<5>276_SW0  (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(VCC),
    .ADR2(CHOICE4465),
    .ADR3(CHOICE4475),
    .O(\CHOICE4475/GROM )
  );
  X_BUF \CHOICE4475/XUSED  (
    .I(\CHOICE4475/FROM ),
    .O(CHOICE4475)
  );
  X_BUF \CHOICE4475/YUSED  (
    .I(\CHOICE4475/GROM ),
    .O(N126556)
  );
  defparam \DLX_EXinst__n0006<5>316 .INIT = 16'hD0C0;
  X_LUT4 \DLX_EXinst__n0006<5>316  (
    .ADR0(DLX_EXinst__n0030_1),
    .ADR1(CHOICE4479),
    .ADR2(DLX_EXinst__n0149),
    .ADR3(CHOICE4440),
    .O(\DLX_EXinst_ALU_result<5>/FROM )
  );
  defparam \DLX_EXinst__n0006<5>326 .INIT = 16'hFFF0;
  X_LUT4 \DLX_EXinst__n0006<5>326  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N63689),
    .ADR3(CHOICE4481),
    .O(\DLX_EXinst_ALU_result<5>/GROM )
  );
  X_BUF \DLX_EXinst_ALU_result<5>/XUSED  (
    .I(\DLX_EXinst_ALU_result<5>/FROM ),
    .O(CHOICE4481)
  );
  X_BUF \DLX_EXinst_ALU_result<5>/YUSED  (
    .I(\DLX_EXinst_ALU_result<5>/GROM ),
    .O(N116396)
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<25>1 .INIT = 16'h7250;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<25>1  (
    .ADR0(DLX_IDinst__n0147),
    .ADR1(DLX_opcode_of_WB[2]),
    .ADR2(DLX_MEMinst_RF_data_in[25]),
    .ADR3(DLX_IDinst_Mmux__n0148__net123),
    .O(\DLX_IDinst_WB_data_eff<25>/FROM )
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<24>1 .INIT = 16'h50CC;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<24>1  (
    .ADR0(DLX_opcode_of_WB[2]),
    .ADR1(DLX_MEMinst_RF_data_in[24]),
    .ADR2(DLX_IDinst_Mmux__n0148__net123),
    .ADR3(DLX_IDinst__n0147),
    .O(\DLX_IDinst_WB_data_eff<25>/GROM )
  );
  X_BUF \DLX_IDinst_WB_data_eff<25>/XUSED  (
    .I(\DLX_IDinst_WB_data_eff<25>/FROM ),
    .O(DLX_IDinst_WB_data_eff[25])
  );
  X_BUF \DLX_IDinst_WB_data_eff<25>/YUSED  (
    .I(\DLX_IDinst_WB_data_eff<25>/GROM ),
    .O(DLX_IDinst_WB_data_eff[24])
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<19>1 .INIT = 16'h50CC;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<19>1  (
    .ADR0(DLX_opcode_of_WB[2]),
    .ADR1(DLX_MEMinst_RF_data_in[19]),
    .ADR2(DLX_IDinst_Mmux__n0148__net123),
    .ADR3(DLX_IDinst__n0147),
    .O(\DLX_IDinst_WB_data_eff<19>/FROM )
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<16>1 .INIT = 16'h4F40;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<16>1  (
    .ADR0(DLX_opcode_of_WB[2]),
    .ADR1(DLX_IDinst_Mmux__n0148__net123),
    .ADR2(DLX_IDinst__n0147),
    .ADR3(DLX_MEMinst_RF_data_in[16]),
    .O(\DLX_IDinst_WB_data_eff<19>/GROM )
  );
  X_BUF \DLX_IDinst_WB_data_eff<19>/XUSED  (
    .I(\DLX_IDinst_WB_data_eff<19>/FROM ),
    .O(DLX_IDinst_WB_data_eff[19])
  );
  X_BUF \DLX_IDinst_WB_data_eff<19>/YUSED  (
    .I(\DLX_IDinst_WB_data_eff<19>/GROM ),
    .O(DLX_IDinst_WB_data_eff[16])
  );
  defparam DLX_EXinst__n003550.INIT = 16'hFFFE;
  X_LUT4 DLX_EXinst__n003550 (
    .ADR0(DLX_IDinst_reg_out_B[15]),
    .ADR1(DLX_IDinst_reg_out_B[14]),
    .ADR2(DLX_IDinst_reg_out_B[13]),
    .ADR3(DLX_IDinst_reg_out_B[12]),
    .O(\CHOICE3551/FROM )
  );
  defparam DLX_EXinst_Ker6630796.INIT = 16'h0001;
  X_LUT4 DLX_EXinst_Ker6630796 (
    .ADR0(DLX_IDinst_reg_out_B[16]),
    .ADR1(DLX_IDinst_reg_out_B[17]),
    .ADR2(DLX_IDinst_reg_out_B[14]),
    .ADR3(DLX_IDinst_reg_out_B[15]),
    .O(\CHOICE3551/GROM )
  );
  X_BUF \CHOICE3551/XUSED  (
    .I(\CHOICE3551/FROM ),
    .O(CHOICE3551)
  );
  X_BUF \CHOICE3551/YUSED  (
    .I(\CHOICE3551/GROM ),
    .O(CHOICE3595)
  );
  defparam DLX_EXinst_Ker6538495.INIT = 16'h30AA;
  X_LUT4 DLX_EXinst_Ker6538495 (
    .ADR0(DLX_EXinst_N63031),
    .ADR1(DLX_IDinst_IR_function_field_3_1),
    .ADR2(\DLX_EXinst_Mshift__n0024_Sh[27] ),
    .ADR3(DLX_IDinst_IR_function_field_2_1),
    .O(\CHOICE3024/FROM )
  );
  defparam DLX_EXinst_Ker6538412.INIT = 16'hEA40;
  X_LUT4 DLX_EXinst_Ker6538412 (
    .ADR0(DLX_IDinst_IR_function_field_3_1),
    .ADR1(\DLX_EXinst_Mshift__n0024_Sh[27] ),
    .ADR2(DLX_IDinst_IR_function_field_2_1),
    .ADR3(DLX_IDinst_reg_out_A[31]),
    .O(\CHOICE3024/GROM )
  );
  X_BUF \CHOICE3024/XUSED  (
    .I(\CHOICE3024/FROM ),
    .O(CHOICE3024)
  );
  X_BUF \CHOICE3024/YUSED  (
    .I(\CHOICE3024/GROM ),
    .O(CHOICE3007)
  );
  defparam \DLX_EXinst__n0006<20>96_SW0 .INIT = 16'h0055;
  X_LUT4 \DLX_EXinst__n0006<20>96_SW0  (
    .ADR0(DLX_IDinst_reg_out_A[20]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_IR_opcode_field[0]),
    .O(\N127338/FROM )
  );
  defparam \DLX_EXinst__n0006<25>36_SW0 .INIT = 16'h0505;
  X_LUT4 \DLX_EXinst__n0006<25>36_SW0  (
    .ADR0(DLX_IDinst_IR_opcode_field[0]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[25]),
    .ADR3(VCC),
    .O(\N127338/GROM )
  );
  X_BUF \N127338/XUSED  (
    .I(\N127338/FROM ),
    .O(N127338)
  );
  X_BUF \N127338/YUSED  (
    .I(\N127338/GROM ),
    .O(N127330)
  );
  defparam \DLX_EXinst__n0006<26>36_SW0 .INIT = 16'h1111;
  X_LUT4 \DLX_EXinst__n0006<26>36_SW0  (
    .ADR0(DLX_IDinst_reg_out_A[26]),
    .ADR1(DLX_IDinst_IR_opcode_field[0]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\N127342/FROM )
  );
  defparam \DLX_EXinst__n0006<24>76_SW0 .INIT = 16'h0055;
  X_LUT4 \DLX_EXinst__n0006<24>76_SW0  (
    .ADR0(DLX_IDinst_reg_out_A[24]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_IR_opcode_field[0]),
    .O(\N127342/GROM )
  );
  X_BUF \N127342/XUSED  (
    .I(\N127342/FROM ),
    .O(N127342)
  );
  X_BUF \N127342/YUSED  (
    .I(\N127342/GROM ),
    .O(N127358)
  );
  defparam DLX_IDinst_Ker697791.INIT = 16'hBBFF;
  X_LUT4 DLX_IDinst_Ker697791 (
    .ADR0(DLX_IDinst_IR_latched[30]),
    .ADR1(DLX_IDinst_IR_latched[27]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_N70991),
    .O(\DLX_IDinst_N69781/FROM )
  );
  defparam DLX_IDinst__n0108120.INIT = 16'h0100;
  X_LUT4 DLX_IDinst__n0108120 (
    .ADR0(DLX_IDinst__n0364),
    .ADR1(DLX_IDinst__n0135),
    .ADR2(DLX_IDinst__n0136),
    .ADR3(DLX_IDinst_N69781),
    .O(\DLX_IDinst_N69781/GROM )
  );
  X_BUF \DLX_IDinst_N69781/XUSED  (
    .I(\DLX_IDinst_N69781/FROM ),
    .O(DLX_IDinst_N69781)
  );
  X_BUF \DLX_IDinst_N69781/YUSED  (
    .I(\DLX_IDinst_N69781/GROM ),
    .O(CHOICE3457)
  );
  defparam \DLX_EXinst__n0006<9>210 .INIT = 16'hCE00;
  X_LUT4 \DLX_EXinst__n0006<9>210  (
    .ADR0(DLX_EXinst__n0047),
    .ADR1(DLX_EXinst__n0046),
    .ADR2(DLX_IDinst_reg_out_A[9]),
    .ADR3(DLX_IDinst_reg_out_B[9]),
    .O(\CHOICE4596/FROM )
  );
  defparam \DLX_EXinst__n0006<5>247 .INIT = 16'hB0A0;
  X_LUT4 \DLX_EXinst__n0006<5>247  (
    .ADR0(DLX_EXinst__n0046),
    .ADR1(DLX_IDinst_reg_out_A[5]),
    .ADR2(DLX_IDinst_reg_out_B[5]),
    .ADR3(DLX_EXinst__n0047),
    .O(\CHOICE4596/GROM )
  );
  X_BUF \CHOICE4596/XUSED  (
    .I(\CHOICE4596/FROM ),
    .O(CHOICE4596)
  );
  X_BUF \CHOICE4596/YUSED  (
    .I(\CHOICE4596/GROM ),
    .O(CHOICE4472)
  );
  defparam \DLX_EXinst__n0006<31>306 .INIT = 16'h0E04;
  X_LUT4 \DLX_EXinst__n0006<31>306  (
    .ADR0(DLX_IDinst_IR_function_field[1]),
    .ADR1(DLX_IDinst_reg_out_A[31]),
    .ADR2(DLX_IDinst_IR_function_field[0]),
    .ADR3(DLX_IDinst_reg_out_A[29]),
    .O(\CHOICE5801/FROM )
  );
  defparam DLX_EXinst_Ker6481710.INIT = 16'hA280;
  X_LUT4 DLX_EXinst_Ker6481710 (
    .ADR0(DLX_IDinst_IR_function_field[3]),
    .ADR1(DLX_IDinst_IR_function_field[0]),
    .ADR2(DLX_EXinst_N63011),
    .ADR3(DLX_EXinst_N63514),
    .O(\CHOICE5801/GROM )
  );
  X_BUF \CHOICE5801/XUSED  (
    .I(\CHOICE5801/FROM ),
    .O(CHOICE5801)
  );
  X_BUF \CHOICE5801/YUSED  (
    .I(\CHOICE5801/GROM ),
    .O(CHOICE1210)
  );
  defparam DLX_EXinst_Ker6480726.INIT = 16'h00E2;
  X_LUT4 DLX_EXinst_Ker6480726 (
    .ADR0(DLX_EXinst_N62921),
    .ADR1(DLX_IDinst_IR_function_field[0]),
    .ADR2(DLX_EXinst_N63339),
    .ADR3(DLX_IDinst_IR_function_field[3]),
    .O(\CHOICE1096/FROM )
  );
  defparam DLX_EXinst_Ker6480728.INIT = 16'hFFCC;
  X_LUT4 DLX_EXinst_Ker6480728 (
    .ADR0(VCC),
    .ADR1(CHOICE1090),
    .ADR2(VCC),
    .ADR3(CHOICE1096),
    .O(\CHOICE1096/GROM )
  );
  X_BUF \CHOICE1096/XUSED  (
    .I(\CHOICE1096/FROM ),
    .O(CHOICE1096)
  );
  X_BUF \CHOICE1096/YUSED  (
    .I(\CHOICE1096/GROM ),
    .O(N96513)
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<18>1 .INIT = 16'h30B8;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<18>1  (
    .ADR0(DLX_IDinst_Mmux__n0148__net123),
    .ADR1(DLX_IDinst__n0147),
    .ADR2(DLX_MEMinst_RF_data_in[18]),
    .ADR3(DLX_opcode_of_WB[2]),
    .O(\DLX_IDinst_WB_data_eff<18>/FROM )
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<17>1 .INIT = 16'h7340;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<17>1  (
    .ADR0(DLX_opcode_of_WB[2]),
    .ADR1(DLX_IDinst__n0147),
    .ADR2(DLX_IDinst_Mmux__n0148__net123),
    .ADR3(DLX_MEMinst_RF_data_in[17]),
    .O(\DLX_IDinst_WB_data_eff<18>/GROM )
  );
  X_BUF \DLX_IDinst_WB_data_eff<18>/XUSED  (
    .I(\DLX_IDinst_WB_data_eff<18>/FROM ),
    .O(DLX_IDinst_WB_data_eff[18])
  );
  X_BUF \DLX_IDinst_WB_data_eff<18>/YUSED  (
    .I(\DLX_IDinst_WB_data_eff<18>/GROM ),
    .O(DLX_IDinst_WB_data_eff[17])
  );
  defparam \DLX_EXinst__n0006<1>129_SW0 .INIT = 16'hFBC8;
  X_LUT4 \DLX_EXinst__n0006<1>129_SW0  (
    .ADR0(CHOICE1108),
    .ADR1(DLX_IDinst_IR_function_field[2]),
    .ADR2(CHOICE1102),
    .ADR3(N127444),
    .O(\N126571/FROM )
  );
  defparam DLX_EXinst__n000520.INIT = 16'h0001;
  X_LUT4 DLX_EXinst__n000520 (
    .ADR0(DLX_IDinst_IR_function_field[3]),
    .ADR1(DLX_IDinst_IR_function_field[1]),
    .ADR2(DLX_IDinst_IR_function_field[2]),
    .ADR3(DLX_IDinst_IR_function_field[4]),
    .O(\N126571/GROM )
  );
  X_BUF \N126571/XUSED  (
    .I(\N126571/FROM ),
    .O(N126571)
  );
  X_BUF \N126571/YUSED  (
    .I(\N126571/GROM ),
    .O(CHOICE2008)
  );
  defparam \DLX_EXinst_Mshift__n0027_Sh<2>_SW0 .INIT = 16'h03F3;
  X_LUT4 \DLX_EXinst_Mshift__n0027_Sh<2>_SW0  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[2]),
    .ADR2(DLX_IDinst_IR_function_field_1_1),
    .ADR3(DLX_IDinst_reg_out_A[0]),
    .O(\N94857/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0027_Sh<2> .INIT = 16'h085D;
  X_LUT4 \DLX_EXinst_Mshift__n0027_Sh<2>  (
    .ADR0(DLX_IDinst_IR_function_field_0_1),
    .ADR1(DLX_IDinst_reg_out_A[1]),
    .ADR2(DLX_IDinst_IR_function_field_1_1),
    .ADR3(N94857),
    .O(\N94857/GROM )
  );
  X_BUF \N94857/XUSED  (
    .I(\N94857/FROM ),
    .O(N94857)
  );
  X_BUF \N94857/YUSED  (
    .I(\N94857/GROM ),
    .O(\DLX_EXinst_Mshift__n0027_Sh[2] )
  );
  defparam \DLX_EXinst__n0006<6>124 .INIT = 16'hF8F8;
  X_LUT4 \DLX_EXinst__n0006<6>124  (
    .ADR0(DLX_IDinst_reg_out_B[6]),
    .ADR1(DLX_EXinst__n0045),
    .ADR2(DLX_EXinst_N64448),
    .ADR3(VCC),
    .O(\CHOICE4378/FROM )
  );
  defparam \DLX_EXinst__n0006<6>133 .INIT = 16'hAA08;
  X_LUT4 \DLX_EXinst__n0006<6>133  (
    .ADR0(DLX_IDinst_reg_out_A[6]),
    .ADR1(DLX_EXinst__n0047),
    .ADR2(DLX_IDinst_reg_out_B[6]),
    .ADR3(CHOICE4378),
    .O(\CHOICE4378/GROM )
  );
  X_BUF \CHOICE4378/XUSED  (
    .I(\CHOICE4378/FROM ),
    .O(CHOICE4378)
  );
  X_BUF \CHOICE4378/YUSED  (
    .I(\CHOICE4378/GROM ),
    .O(CHOICE4380)
  );
  defparam \DLX_EXinst__n0006<5>276 .INIT = 16'hF0E0;
  X_LUT4 \DLX_EXinst__n0006<5>276  (
    .ADR0(CHOICE4472),
    .ADR1(CHOICE4448),
    .ADR2(DLX_EXinst__n0030_1),
    .ADR3(N126556),
    .O(\CHOICE4478/FROM )
  );
  defparam \DLX_EXinst__n0006<5>288 .INIT = 16'hFFC0;
  X_LUT4 \DLX_EXinst__n0006<5>288  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst__n0016[5]),
    .ADR2(DLX_EXinst_N63836),
    .ADR3(CHOICE4478),
    .O(\CHOICE4478/GROM )
  );
  X_BUF \CHOICE4478/XUSED  (
    .I(\CHOICE4478/FROM ),
    .O(CHOICE4478)
  );
  X_BUF \CHOICE4478/YUSED  (
    .I(\CHOICE4478/GROM ),
    .O(CHOICE4479)
  );
  defparam \DLX_EXinst__n0006<6>197 .INIT = 16'hFAF8;
  X_LUT4 \DLX_EXinst__n0006<6>197  (
    .ADR0(DLX_EXinst_N62631),
    .ADR1(CHOICE4385),
    .ADR2(CHOICE4396),
    .ADR3(CHOICE4391),
    .O(\CHOICE4397/FROM )
  );
  defparam \DLX_EXinst__n0006<5>197 .INIT = 16'hFAF8;
  X_LUT4 \DLX_EXinst__n0006<5>197  (
    .ADR0(DLX_EXinst_N62631),
    .ADR1(CHOICE4453),
    .ADR2(CHOICE4464),
    .ADR3(CHOICE4459),
    .O(\CHOICE4397/GROM )
  );
  X_BUF \CHOICE4397/XUSED  (
    .I(\CHOICE4397/FROM ),
    .O(CHOICE4397)
  );
  X_BUF \CHOICE4397/YUSED  (
    .I(\CHOICE4397/GROM ),
    .O(CHOICE4465)
  );
  defparam DLX_IDinst_Ker699558.INIT = 16'h0C0C;
  X_LUT4 DLX_IDinst_Ker699558 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_IR_opcode_field[4]),
    .ADR2(DLX_IDinst_IR_opcode_field[5]),
    .ADR3(VCC),
    .O(\CHOICE1417/FROM )
  );
  defparam DLX_IDinst_Ker6995512.INIT = 16'h8A00;
  X_LUT4 DLX_IDinst_Ker6995512 (
    .ADR0(DLX_IDinst_IR_opcode_field[2]),
    .ADR1(DLX_IDinst_IR_opcode_field[1]),
    .ADR2(DLX_IDinst_IR_opcode_field[0]),
    .ADR3(CHOICE1417),
    .O(\CHOICE1417/GROM )
  );
  X_BUF \CHOICE1417/XUSED  (
    .I(\CHOICE1417/FROM ),
    .O(CHOICE1417)
  );
  X_BUF \CHOICE1417/YUSED  (
    .I(\CHOICE1417/GROM ),
    .O(CHOICE1418)
  );
  defparam \DLX_EXinst_Mshift__n0026_Sh<49>1 .INIT = 16'hEE22;
  X_LUT4 \DLX_EXinst_Mshift__n0026_Sh<49>1  (
    .ADR0(DLX_EXinst_N64329),
    .ADR1(DLX_IDinst_reg_out_B_2_1),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N63071),
    .O(\DLX_EXinst_Mshift__n0026_Sh<49>/FROM )
  );
  defparam \DLX_EXinst__n0006<17>302_SW0 .INIT = 16'hFAAA;
  X_LUT4 \DLX_EXinst__n0006<17>302_SW0  (
    .ADR0(CHOICE5637),
    .ADR1(VCC),
    .ADR2(DLX_EXinst__n0049),
    .ADR3(\DLX_EXinst_Mshift__n0026_Sh[49] ),
    .O(\DLX_EXinst_Mshift__n0026_Sh<49>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0026_Sh<49>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0026_Sh<49>/FROM ),
    .O(\DLX_EXinst_Mshift__n0026_Sh[49] )
  );
  X_BUF \DLX_EXinst_Mshift__n0026_Sh<49>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0026_Sh<49>/GROM ),
    .O(N126610)
  );
  defparam DLX_EXinst_Ker6481726.INIT = 16'h00AC;
  X_LUT4 DLX_EXinst_Ker6481726 (
    .ADR0(DLX_EXinst_N62991),
    .ADR1(DLX_EXinst_N63494),
    .ADR2(DLX_IDinst_IR_function_field[0]),
    .ADR3(DLX_IDinst_IR_function_field[3]),
    .O(\CHOICE1216/FROM )
  );
  defparam DLX_EXinst_Ker6481728.INIT = 16'hFFF0;
  X_LUT4 DLX_EXinst_Ker6481728 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(CHOICE1210),
    .ADR3(CHOICE1216),
    .O(\CHOICE1216/GROM )
  );
  X_BUF \CHOICE1216/XUSED  (
    .I(\CHOICE1216/FROM ),
    .O(CHOICE1216)
  );
  X_BUF \CHOICE1216/YUSED  (
    .I(\CHOICE1216/GROM ),
    .O(N97233)
  );
  defparam DLX_EXinst_Ker6624854.INIT = 16'h0400;
  X_LUT4 DLX_EXinst_Ker6624854 (
    .ADR0(\DLX_IDinst_Imm[31] ),
    .ADR1(DLX_IDinst_IR_opcode_field[0]),
    .ADR2(\DLX_IDinst_Imm[6] ),
    .ADR3(N125999),
    .O(\CHOICE3377/FROM )
  );
  defparam DLX_EXinst_Ker66248157.INIT = 16'hCC00;
  X_LUT4 DLX_EXinst_Ker66248157 (
    .ADR0(VCC),
    .ADR1(CHOICE3408),
    .ADR2(VCC),
    .ADR3(CHOICE3377),
    .O(\CHOICE3377/GROM )
  );
  X_BUF \CHOICE3377/XUSED  (
    .I(\CHOICE3377/FROM ),
    .O(CHOICE3377)
  );
  X_BUF \CHOICE3377/YUSED  (
    .I(\CHOICE3377/GROM ),
    .O(N110065)
  );
  defparam \DLX_EXinst__n0006<22>312_SW0 .INIT = 16'h00FE;
  X_LUT4 \DLX_EXinst__n0006<22>312_SW0  (
    .ADR0(CHOICE4109),
    .ADR1(CHOICE4123),
    .ADR2(CHOICE4098),
    .ADR3(DLX_EXinst__n0030),
    .O(\DLX_EXinst_ALU_result<22>/FROM )
  );
  defparam \DLX_EXinst__n0006<22>312 .INIT = 16'hAAA8;
  X_LUT4 \DLX_EXinst__n0006<22>312  (
    .ADR0(DLX_EXinst__n0149),
    .ADR1(N100490),
    .ADR2(CHOICE4157),
    .ADR3(N126478),
    .O(N114452)
  );
  X_BUF \DLX_EXinst_ALU_result<22>/XUSED  (
    .I(\DLX_EXinst_ALU_result<22>/FROM ),
    .O(N126478)
  );
  defparam \DLX_EXinst__n0006<6>315 .INIT = 16'hA0A8;
  X_LUT4 \DLX_EXinst__n0006<6>315  (
    .ADR0(DLX_EXinst__n0149),
    .ADR1(CHOICE4372),
    .ADR2(CHOICE4411),
    .ADR3(DLX_EXinst__n0030_1),
    .O(\DLX_EXinst_ALU_result<6>/FROM )
  );
  defparam \DLX_EXinst__n0006<6>325 .INIT = 16'hFFAA;
  X_LUT4 \DLX_EXinst__n0006<6>325  (
    .ADR0(DLX_EXinst_N63689),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(CHOICE4413),
    .O(\DLX_EXinst_ALU_result<6>/GROM )
  );
  X_BUF \DLX_EXinst_ALU_result<6>/XUSED  (
    .I(\DLX_EXinst_ALU_result<6>/FROM ),
    .O(CHOICE4413)
  );
  X_BUF \DLX_EXinst_ALU_result<6>/YUSED  (
    .I(\DLX_EXinst_ALU_result<6>/GROM ),
    .O(N115984)
  );
  defparam \DLX_EXinst__n0006<6>251 .INIT = 16'hF888;
  X_LUT4 \DLX_EXinst__n0006<6>251  (
    .ADR0(N108909),
    .ADR1(DLX_IDinst_reg_out_B[4]),
    .ADR2(DLX_EXinst_ALU_result[6]),
    .ADR3(N101725),
    .O(\CHOICE4407/FROM )
  );
  defparam \DLX_EXinst__n0006<6>275_SW0 .INIT = 16'hFF50;
  X_LUT4 \DLX_EXinst__n0006<6>275_SW0  (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(VCC),
    .ADR2(CHOICE4397),
    .ADR3(CHOICE4407),
    .O(\CHOICE4407/GROM )
  );
  X_BUF \CHOICE4407/XUSED  (
    .I(\CHOICE4407/FROM ),
    .O(CHOICE4407)
  );
  X_BUF \CHOICE4407/YUSED  (
    .I(\CHOICE4407/GROM ),
    .O(N126614)
  );
  defparam DLX_EXinst_Ker6539426.INIT = 16'h2320;
  X_LUT4 DLX_EXinst_Ker6539426 (
    .ADR0(DLX_EXinst_N63334),
    .ADR1(DLX_IDinst_IR_function_field_3_1),
    .ADR2(DLX_IDinst_IR_function_field[0]),
    .ADR3(DLX_EXinst_N62976),
    .O(\CHOICE1108/FROM )
  );
  defparam DLX_EXinst_Ker6539428.INIT = 16'hFFF0;
  X_LUT4 DLX_EXinst_Ker6539428 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(CHOICE1102),
    .ADR3(CHOICE1108),
    .O(\CHOICE1108/GROM )
  );
  X_BUF \CHOICE1108/XUSED  (
    .I(\CHOICE1108/FROM ),
    .O(CHOICE1108)
  );
  X_BUF \CHOICE1108/YUSED  (
    .I(\CHOICE1108/GROM ),
    .O(N96585)
  );
  defparam \DLX_EXinst__n0006<29>253 .INIT = 16'hA0A8;
  X_LUT4 \DLX_EXinst__n0006<29>253  (
    .ADR0(DLX_IDinst_reg_out_B[29]),
    .ADR1(DLX_EXinst__n0047),
    .ADR2(DLX_EXinst__n0046),
    .ADR3(DLX_IDinst_reg_out_A[29]),
    .O(\CHOICE5383/FROM )
  );
  defparam \DLX_EXinst__n0006<6>246 .INIT = 16'hF400;
  X_LUT4 \DLX_EXinst__n0006<6>246  (
    .ADR0(DLX_IDinst_reg_out_A[6]),
    .ADR1(DLX_EXinst__n0047),
    .ADR2(DLX_EXinst__n0046),
    .ADR3(DLX_IDinst_reg_out_B[6]),
    .O(\CHOICE5383/GROM )
  );
  X_BUF \CHOICE5383/XUSED  (
    .I(\CHOICE5383/FROM ),
    .O(CHOICE5383)
  );
  X_BUF \CHOICE5383/YUSED  (
    .I(\CHOICE5383/GROM ),
    .O(CHOICE4404)
  );
  defparam DLX_EXlc_md_mda21_a1.INIT = 16'h00CC;
  X_LUT4 DLX_EXlc_md_mda21_a1 (
    .ADR0(VCC),
    .ADR1(DLX_EXlc_md_wint20),
    .ADR2(VCC),
    .ADR3(DLX_EXlc_pd_wint5),
    .O(\DLX_EXlc_md_wint21/FROM )
  );
  defparam DLX_EXlc_md_mda10_a1.INIT = 16'h00CC;
  X_LUT4 DLX_EXlc_md_mda10_a1 (
    .ADR0(VCC),
    .ADR1(DLX_EXlc_md_wint9),
    .ADR2(VCC),
    .ADR3(DLX_EXlc_pd_wint5),
    .O(\DLX_EXlc_md_wint21/GROM )
  );
  X_BUF \DLX_EXlc_md_wint21/XUSED  (
    .I(\DLX_EXlc_md_wint21/FROM ),
    .O(DLX_EXlc_md_wint21)
  );
  X_BUF \DLX_EXlc_md_wint21/YUSED  (
    .I(\DLX_EXlc_md_wint21/GROM ),
    .O(DLX_EXlc_md_wint10)
  );
  defparam DLX_EXinst_Ker6482736.INIT = 16'h5140;
  X_LUT4 DLX_EXinst_Ker6482736 (
    .ADR0(DLX_IDinst_reg_out_B[5]),
    .ADR1(DLX_IDinst_reg_out_B_2_1),
    .ADR2(DLX_EXinst_N62966),
    .ADR3(DLX_EXinst_N64329),
    .O(\CHOICE1926/FROM )
  );
  defparam DLX_EXinst_Ker6482739.INIT = 16'hFFC0;
  X_LUT4 DLX_EXinst_Ker6482739 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_B[5]),
    .ADR2(CHOICE1919),
    .ADR3(CHOICE1926),
    .O(\CHOICE1926/GROM )
  );
  X_BUF \CHOICE1926/XUSED  (
    .I(\CHOICE1926/FROM ),
    .O(CHOICE1926)
  );
  X_BUF \CHOICE1926/YUSED  (
    .I(\CHOICE1926/GROM ),
    .O(N101425)
  );
  defparam \DLX_EXinst__n0006<6>275 .INIT = 16'hAAA8;
  X_LUT4 \DLX_EXinst__n0006<6>275  (
    .ADR0(DLX_EXinst__n0030_1),
    .ADR1(N126614),
    .ADR2(CHOICE4380),
    .ADR3(CHOICE4404),
    .O(\CHOICE4410/FROM )
  );
  defparam \DLX_EXinst__n0006<6>287 .INIT = 16'hFFA0;
  X_LUT4 \DLX_EXinst__n0006<6>287  (
    .ADR0(DLX_EXinst__n0016[6]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N63836),
    .ADR3(CHOICE4410),
    .O(\CHOICE4410/GROM )
  );
  X_BUF \CHOICE4410/XUSED  (
    .I(\CHOICE4410/FROM ),
    .O(CHOICE4410)
  );
  X_BUF \CHOICE4410/YUSED  (
    .I(\CHOICE4410/GROM ),
    .O(CHOICE4411)
  );
  defparam \DLX_EXinst__n0006<7>124 .INIT = 16'hFAF0;
  X_LUT4 \DLX_EXinst__n0006<7>124  (
    .ADR0(DLX_EXinst__n0045),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N64448),
    .ADR3(DLX_IDinst_reg_out_B[7]),
    .O(\CHOICE3826/FROM )
  );
  defparam \DLX_EXinst__n0006<7>133 .INIT = 16'hF020;
  X_LUT4 \DLX_EXinst__n0006<7>133  (
    .ADR0(DLX_EXinst__n0047),
    .ADR1(DLX_IDinst_reg_out_B[7]),
    .ADR2(DLX_IDinst_reg_out_A[7]),
    .ADR3(CHOICE3826),
    .O(\CHOICE3826/GROM )
  );
  X_BUF \CHOICE3826/XUSED  (
    .I(\CHOICE3826/FROM ),
    .O(CHOICE3826)
  );
  X_BUF \CHOICE3826/YUSED  (
    .I(\CHOICE3826/GROM ),
    .O(CHOICE3828)
  );
  defparam \DLX_IDinst__n0086<23>20 .INIT = 16'hAA00;
  X_LUT4 \DLX_IDinst__n0086<23>20  (
    .ADR0(DLX_IDinst_N70295),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_regA_eff[23]),
    .O(\CHOICE2815/FROM )
  );
  defparam \DLX_IDinst__n0086<11>20 .INIT = 16'hC0C0;
  X_LUT4 \DLX_IDinst__n0086<11>20  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_N70295),
    .ADR2(DLX_IDinst_regA_eff[11]),
    .ADR3(VCC),
    .O(\CHOICE2815/GROM )
  );
  X_BUF \CHOICE2815/XUSED  (
    .I(\CHOICE2815/FROM ),
    .O(CHOICE2815)
  );
  X_BUF \CHOICE2815/YUSED  (
    .I(\CHOICE2815/GROM ),
    .O(CHOICE2683)
  );
  defparam DLX_EXinst_Ker6488761.INIT = 16'hB080;
  X_LUT4 DLX_EXinst_Ker6488761 (
    .ADR0(\DLX_EXinst_Mshift__n0026_Sh[30] ),
    .ADR1(DLX_IDinst_reg_out_B_2_1),
    .ADR2(DLX_EXinst_N66494),
    .ADR3(\DLX_EXinst_Mshift__n0023_Sh[26] ),
    .O(\CHOICE3045/FROM )
  );
  defparam DLX_EXinst_Ker6488265.INIT = 16'hAC00;
  X_LUT4 DLX_EXinst_Ker6488265 (
    .ADR0(\DLX_EXinst_Mshift__n0026_Sh[29] ),
    .ADR1(\DLX_EXinst_Mshift__n0023_Sh[25] ),
    .ADR2(DLX_IDinst_reg_out_B_2_1),
    .ADR3(DLX_EXinst_N66494),
    .O(\CHOICE3045/GROM )
  );
  X_BUF \CHOICE3045/XUSED  (
    .I(\CHOICE3045/FROM ),
    .O(CHOICE3045)
  );
  X_BUF \CHOICE3045/YUSED  (
    .I(\CHOICE3045/GROM ),
    .O(CHOICE3152)
  );
  defparam \DLX_EXinst__n0006<9>117 .INIT = 16'hFFA0;
  X_LUT4 \DLX_EXinst__n0006<9>117  (
    .ADR0(DLX_IDinst_reg_out_B[9]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst__n0045),
    .ADR3(DLX_EXinst_N64448),
    .O(\CHOICE4576/FROM )
  );
  defparam \DLX_EXinst__n0006<9>126 .INIT = 16'hCC08;
  X_LUT4 \DLX_EXinst__n0006<9>126  (
    .ADR0(DLX_EXinst__n0047),
    .ADR1(DLX_IDinst_reg_out_A[9]),
    .ADR2(DLX_IDinst_reg_out_B[9]),
    .ADR3(CHOICE4576),
    .O(\CHOICE4576/GROM )
  );
  X_BUF \CHOICE4576/XUSED  (
    .I(\CHOICE4576/FROM ),
    .O(CHOICE4576)
  );
  X_BUF \CHOICE4576/YUSED  (
    .I(\CHOICE4576/GROM ),
    .O(CHOICE4578)
  );
  defparam DLX_IFlc_master_ctrlIF__n00021.INIT = 16'hFF30;
  X_LUT4 DLX_IFlc_master_ctrlIF__n00021 (
    .ADR0(VCC),
    .ADR1(DLX_IFlc_slave_ctrlIF_l),
    .ADR2(DLX_IFlc_master_ctrlIF_nro),
    .ADR3(DLX_IFlc_master_ctrlIF_l),
    .O(\DLX_IFlc_master_ctrlIF_nro/FROM )
  );
  defparam DLX_IFlc_slave_ctrlIF__n00021.INIT = 16'h51F3;
  X_LUT4 DLX_IFlc_slave_ctrlIF__n00021 (
    .ADR0(CHOICE25),
    .ADR1(DLX_ackin_ID),
    .ADR2(DLX_reqout_IF),
    .ADR3(DLX_IFlc_master_ctrlIF_nro),
    .O(\DLX_IFlc_master_ctrlIF_nro/GROM )
  );
  X_BUF \DLX_IFlc_master_ctrlIF_nro/XUSED  (
    .I(\DLX_IFlc_master_ctrlIF_nro/FROM ),
    .O(DLX_IFlc_master_ctrlIF_nro)
  );
  X_BUF \DLX_IFlc_master_ctrlIF_nro/YUSED  (
    .I(\DLX_IFlc_master_ctrlIF_nro/GROM ),
    .O(DLX_reqout_IF)
  );
  defparam DLX_IDinst__n01209.INIT = 16'hD000;
  X_LUT4 DLX_IDinst__n01209 (
    .ADR0(DLX_IDinst__n0077),
    .ADR1(DLX_IDinst__n0002),
    .ADR2(DLX_IDinst__n0350),
    .ADR3(DLX_IDinst__n0348),
    .O(\CHOICE3491/FROM )
  );
  defparam DLX_IDinst__n012018.INIT = 16'h3320;
  X_LUT4 DLX_IDinst__n012018 (
    .ADR0(DLX_IDinst__n0347),
    .ADR1(DLX_IDinst__n0136),
    .ADR2(DLX_IDinst__n0345),
    .ADR3(CHOICE3491),
    .O(\CHOICE3491/GROM )
  );
  X_BUF \CHOICE3491/XUSED  (
    .I(\CHOICE3491/FROM ),
    .O(CHOICE3491)
  );
  X_BUF \CHOICE3491/YUSED  (
    .I(\CHOICE3491/GROM ),
    .O(CHOICE3493)
  );
  defparam \DLX_IDinst__n0086<11>25 .INIT = 16'hF1F0;
  X_LUT4 \DLX_IDinst__n0086<11>25  (
    .ADR0(DLX_IDinst_N70918),
    .ADR1(DLX_IDinst__n0364),
    .ADR2(CHOICE2683),
    .ADR3(CHOICE2679),
    .O(\DLX_IDinst_branch_address<11>/FROM )
  );
  defparam \DLX_IDinst__n0086<11>31 .INIT = 16'hFFA0;
  X_LUT4 \DLX_IDinst__n0086<11>31  (
    .ADR0(N100609),
    .ADR1(VCC),
    .ADR2(DLX_IDinst__n0128[11]),
    .ADR3(CHOICE2684),
    .O(N105787)
  );
  X_BUF \DLX_IDinst_branch_address<11>/XUSED  (
    .I(\DLX_IDinst_branch_address<11>/FROM ),
    .O(CHOICE2684)
  );
  defparam DLX_IDinst__n01321.INIT = 16'hFEFF;
  X_LUT4 DLX_IDinst__n01321 (
    .ADR0(DLX_IDinst_IR_latched[31]),
    .ADR1(DLX_IDinst_IR_latched[28]),
    .ADR2(DLX_IDinst_IR_latched[29]),
    .ADR3(DLX_IDinst_IR_latched[27]),
    .O(\DLX_IDinst_mem_to_reg/FROM )
  );
  defparam DLX_IDinst__n0110_1178.INIT = 16'h4000;
  X_LUT4 DLX_IDinst__n0110_1178 (
    .ADR0(N100496),
    .ADR1(DLX_IDinst__n0133),
    .ADR2(DLX_IDinst_N70679),
    .ADR3(DLX_IDinst__n0132),
    .O(DLX_IDinst__n0110)
  );
  X_BUF \DLX_IDinst_mem_to_reg/XUSED  (
    .I(\DLX_IDinst_mem_to_reg/FROM ),
    .O(DLX_IDinst__n0132)
  );
  defparam DLX_EXlc_md_mda36_a1.INIT = 16'h3030;
  X_LUT4 DLX_EXlc_md_mda36_a1 (
    .ADR0(VCC),
    .ADR1(DLX_EXlc_pd_wint5),
    .ADR2(DLX_EXlc_md_wint35),
    .ADR3(VCC),
    .O(\DLX_EXlc_md_wint36/FROM )
  );
  defparam DLX_EXlc_md_mda15_a1.INIT = 16'h2222;
  X_LUT4 DLX_EXlc_md_mda15_a1 (
    .ADR0(DLX_EXlc_md_wint14),
    .ADR1(DLX_EXlc_pd_wint5),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_EXlc_md_wint36/GROM )
  );
  X_BUF \DLX_EXlc_md_wint36/XUSED  (
    .I(\DLX_EXlc_md_wint36/FROM ),
    .O(DLX_EXlc_md_wint36)
  );
  X_BUF \DLX_EXlc_md_wint36/YUSED  (
    .I(\DLX_EXlc_md_wint36/GROM ),
    .O(DLX_EXlc_md_wint15)
  );
  defparam \DLX_EXinst_Mshift__n0027_Sh<0>1 .INIT = 16'h0050;
  X_LUT4 \DLX_EXinst_Mshift__n0027_Sh<0>1  (
    .ADR0(DLX_IDinst_IR_function_field_0_1),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[0]),
    .ADR3(DLX_IDinst_IR_function_field_1_1),
    .O(\DLX_EXinst_Mshift__n0027_Sh<0>/FROM )
  );
  defparam \DLX_EXinst__n0006<16>99 .INIT = 16'hBAAA;
  X_LUT4 \DLX_EXinst__n0006<16>99  (
    .ADR0(CHOICE5125),
    .ADR1(DLX_EXinst_N62733),
    .ADR2(DLX_IDinst_IR_function_field[4]),
    .ADR3(\DLX_EXinst_Mshift__n0027_Sh[0] ),
    .O(\DLX_EXinst_Mshift__n0027_Sh<0>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0027_Sh<0>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0027_Sh<0>/FROM ),
    .O(\DLX_EXinst_Mshift__n0027_Sh[0] )
  );
  X_BUF \DLX_EXinst_Mshift__n0027_Sh<0>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0027_Sh<0>/GROM ),
    .O(CHOICE5126)
  );
  defparam \DLX_EXinst_Mshift__n0027_Sh<41> .INIT = 16'h0A33;
  X_LUT4 \DLX_EXinst_Mshift__n0027_Sh<41>  (
    .ADR0(\DLX_EXinst_Mshift__n0027_Sh[1] ),
    .ADR1(N127149),
    .ADR2(DLX_IDinst_IR_function_field_2_1),
    .ADR3(DLX_IDinst_IR_function_field_3_1),
    .O(\DLX_EXinst_Mshift__n0027_Sh<41>/FROM )
  );
  defparam \DLX_EXinst__n0006<9>6 .INIT = 16'hECA0;
  X_LUT4 \DLX_EXinst__n0006<9>6  (
    .ADR0(DLX_EXinst_N66373),
    .ADR1(DLX_EXinst_N66525),
    .ADR2(\DLX_EXinst_Mshift__n0028_Sh[57] ),
    .ADR3(\DLX_EXinst_Mshift__n0027_Sh[41] ),
    .O(\DLX_EXinst_Mshift__n0027_Sh<41>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0027_Sh<41>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0027_Sh<41>/FROM ),
    .O(\DLX_EXinst_Mshift__n0027_Sh[41] )
  );
  X_BUF \DLX_EXinst_Mshift__n0027_Sh<41>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0027_Sh<41>/GROM ),
    .O(CHOICE4549)
  );
  defparam \DLX_EXinst__n0006<9>162 .INIT = 16'hAA00;
  X_LUT4 \DLX_EXinst__n0006<9>162  (
    .ADR0(\DLX_EXinst_Mshift__n0025_Sh[41] ),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N66226),
    .O(\CHOICE4588/FROM )
  );
  defparam \DLX_EXinst__n0006<9>239_SW0 .INIT = 16'hF5F4;
  X_LUT4 \DLX_EXinst__n0006<9>239_SW0  (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(CHOICE4587),
    .ADR2(CHOICE4599),
    .ADR3(CHOICE4588),
    .O(\CHOICE4588/GROM )
  );
  X_BUF \CHOICE4588/XUSED  (
    .I(\CHOICE4588/FROM ),
    .O(CHOICE4588)
  );
  X_BUF \CHOICE4588/YUSED  (
    .I(\CHOICE4588/GROM ),
    .O(N126457)
  );
  defparam \DLX_EXinst__n0006<18>410_SW0 .INIT = 16'h3332;
  X_LUT4 \DLX_EXinst__n0006<18>410_SW0  (
    .ADR0(CHOICE5408),
    .ADR1(DLX_EXinst__n0030),
    .ADR2(CHOICE5440),
    .ADR3(CHOICE5411),
    .O(\DLX_EXinst_ALU_result<18>/FROM )
  );
  defparam \DLX_EXinst__n0006<18>410 .INIT = 16'hAAA8;
  X_LUT4 \DLX_EXinst__n0006<18>410  (
    .ADR0(DLX_EXinst__n0149),
    .ADR1(N100490),
    .ADR2(CHOICE5482),
    .ADR3(N126358),
    .O(N122511)
  );
  X_BUF \DLX_EXinst_ALU_result<18>/XUSED  (
    .I(\DLX_EXinst_ALU_result<18>/FROM ),
    .O(N126358)
  );
  defparam \DLX_EXinst__n0006<26>306_SW0 .INIT = 16'h3332;
  X_LUT4 \DLX_EXinst__n0006<26>306_SW0  (
    .ADR0(CHOICE4701),
    .ADR1(DLX_EXinst__n0030),
    .ADR2(CHOICE4676),
    .ADR3(CHOICE4675),
    .O(\DLX_EXinst_ALU_result<26>/FROM )
  );
  defparam \DLX_EXinst__n0006<26>306 .INIT = 16'hCCC8;
  X_LUT4 \DLX_EXinst__n0006<26>306  (
    .ADR0(CHOICE4733),
    .ADR1(DLX_EXinst__n0149),
    .ADR2(N100490),
    .ADR3(N126349),
    .O(N117936)
  );
  X_BUF \DLX_EXinst_ALU_result<26>/XUSED  (
    .I(\DLX_EXinst_ALU_result<26>/FROM ),
    .O(N126349)
  );
  defparam DLX_IDinst__n01229.INIT = 16'hFFFE;
  X_LUT4 DLX_IDinst__n01229 (
    .ADR0(DLX_IDinst_IR_latched[27]),
    .ADR1(DLX_IDinst_IR_latched[29]),
    .ADR2(DLX_IDinst_IR_latched[31]),
    .ADR3(DLX_IDinst_IR_latched[28]),
    .O(\CHOICE3295/FROM )
  );
  defparam DLX_IDinst__n012219.INIT = 16'hCCC4;
  X_LUT4 DLX_IDinst__n012219 (
    .ADR0(DLX_IDinst_IR_latched[30]),
    .ADR1(DLX_IDinst_delay_slot),
    .ADR2(DLX_IDinst_IR_latched[26]),
    .ADR3(CHOICE3295),
    .O(\CHOICE3295/GROM )
  );
  X_BUF \CHOICE3295/XUSED  (
    .I(\CHOICE3295/FROM ),
    .O(CHOICE3295)
  );
  X_BUF \CHOICE3295/YUSED  (
    .I(\CHOICE3295/GROM ),
    .O(CHOICE3297)
  );
  defparam \DLX_EXinst_Mshift__n0027_Sh<3>11 .INIT = 16'hC480;
  X_LUT4 \DLX_EXinst_Mshift__n0027_Sh<3>11  (
    .ADR0(DLX_IDinst_IR_function_field_0_1),
    .ADR1(DLX_IDinst_IR_function_field_1_1),
    .ADR2(DLX_IDinst_reg_out_A[0]),
    .ADR3(DLX_IDinst_reg_out_A[1]),
    .O(\CHOICE994/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0027_Sh<1>1 .INIT = 16'h3120;
  X_LUT4 \DLX_EXinst_Mshift__n0027_Sh<1>1  (
    .ADR0(DLX_IDinst_IR_function_field_0_1),
    .ADR1(DLX_IDinst_IR_function_field_1_1),
    .ADR2(DLX_IDinst_reg_out_A[0]),
    .ADR3(DLX_IDinst_reg_out_A[1]),
    .O(\CHOICE994/GROM )
  );
  X_BUF \CHOICE994/XUSED  (
    .I(\CHOICE994/FROM ),
    .O(CHOICE994)
  );
  X_BUF \CHOICE994/YUSED  (
    .I(\CHOICE994/GROM ),
    .O(\DLX_EXinst_Mshift__n0027_Sh[1] )
  );
  defparam DLX_RF_delay_inst_wint41.INIT = 16'h00FF;
  X_LUT4 DLX_RF_delay_inst_wint41 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_RF_delay_inst_wint3),
    .O(\DLX_RF_delay_inst_wint4/GROM )
  );
  X_BUF \DLX_RF_delay_inst_wint4/YUSED  (
    .I(\DLX_RF_delay_inst_wint4/GROM ),
    .O(DLX_RF_delay_inst_wint4)
  );
  defparam DLX_EXinst_Ker6489291.INIT = 16'h2322;
  X_LUT4 DLX_EXinst_Ker6489291 (
    .ADR0(CHOICE2548),
    .ADR1(DLX_IDinst_reg_out_B_3_1),
    .ADR2(DLX_IDinst_reg_out_B_2_1),
    .ADR3(\DLX_EXinst_Mshift__n0023_Sh[27] ),
    .O(\CHOICE2551/FROM )
  );
  defparam DLX_EXinst_Ker64892105.INIT = 16'hEAC0;
  X_LUT4 DLX_EXinst_Ker64892105 (
    .ADR0(DLX_EXinst_N66494),
    .ADR1(N111221),
    .ADR2(CHOICE2542),
    .ADR3(CHOICE2551),
    .O(\CHOICE2551/GROM )
  );
  X_BUF \CHOICE2551/XUSED  (
    .I(\CHOICE2551/FROM ),
    .O(CHOICE2551)
  );
  X_BUF \CHOICE2551/YUSED  (
    .I(\CHOICE2551/GROM ),
    .O(N105035)
  );
  defparam DLX_IDinst__n00711.INIT = 16'h5000;
  X_LUT4 DLX_IDinst__n00711 (
    .ADR0(DLX_IDinst_IR_latched[27]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_IR_latched[30]),
    .ADR3(DLX_IDinst_N70991),
    .O(\DLX_IDinst_CLI/FROM )
  );
  defparam DLX_IDinst__n01241.INIT = 16'hB8BA;
  X_LUT4 DLX_IDinst__n01241 (
    .ADR0(DLX_IDinst_CLI),
    .ADR1(DLX_IDinst_N70918),
    .ADR2(DLX_IDinst__n0364),
    .ADR3(DLX_IDinst__n0071),
    .O(\DLX_IDinst_CLI/GROM )
  );
  X_BUF \DLX_IDinst_CLI/XUSED  (
    .I(\DLX_IDinst_CLI/FROM ),
    .O(DLX_IDinst__n0071)
  );
  X_BUF \DLX_IDinst_CLI/YUSED  (
    .I(\DLX_IDinst_CLI/GROM ),
    .O(DLX_IDinst__n0124)
  );
  defparam DLX_IDinst__n01351.INIT = 16'hAA8A;
  X_LUT4 DLX_IDinst__n01351 (
    .ADR0(DLX_IDinst__n0073),
    .ADR1(DLX_IDinst_regA_index[1]),
    .ADR2(DLX_IDinst_N70658),
    .ADR3(DLX_IDinst_regA_index[0]),
    .O(\DLX_IDinst__n0135/FROM )
  );
  defparam DLX_IDinst_Ker706081.INIT = 16'h000B;
  X_LUT4 DLX_IDinst_Ker706081 (
    .ADR0(DLX_IDinst__n0004),
    .ADR1(DLX_IDinst__n0075),
    .ADR2(DLX_IDinst__n0345),
    .ADR3(DLX_IDinst__n0135),
    .O(\DLX_IDinst__n0135/GROM )
  );
  X_BUF \DLX_IDinst__n0135/XUSED  (
    .I(\DLX_IDinst__n0135/FROM ),
    .O(DLX_IDinst__n0135)
  );
  X_BUF \DLX_IDinst__n0135/YUSED  (
    .I(\DLX_IDinst__n0135/GROM ),
    .O(DLX_IDinst_N70610)
  );
  defparam DLX_RF_delay_inst_wint51.INIT = 16'h0F0F;
  X_LUT4 DLX_RF_delay_inst_wint51 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_RF_delay_inst_wint4),
    .ADR3(VCC),
    .O(\DLX_RF_delay_inst_wint5/GROM )
  );
  X_BUF \DLX_RF_delay_inst_wint5/YUSED  (
    .I(\DLX_RF_delay_inst_wint5/GROM ),
    .O(DLX_RF_delay_inst_wint5)
  );
  defparam \DLX_EXinst__n0006<9>239 .INIT = 16'hAAA8;
  X_LUT4 \DLX_EXinst__n0006<9>239  (
    .ADR0(DLX_EXinst__n0030_1),
    .ADR1(N126457),
    .ADR2(CHOICE4578),
    .ADR3(CHOICE4596),
    .O(\CHOICE4602/FROM )
  );
  defparam \DLX_EXinst__n0006<9>251 .INIT = 16'hFFA0;
  X_LUT4 \DLX_EXinst__n0006<9>251  (
    .ADR0(DLX_EXinst_N63836),
    .ADR1(VCC),
    .ADR2(DLX_EXinst__n0016[9]),
    .ADR3(CHOICE4602),
    .O(\CHOICE4602/GROM )
  );
  X_BUF \CHOICE4602/XUSED  (
    .I(\CHOICE4602/FROM ),
    .O(CHOICE4602)
  );
  X_BUF \CHOICE4602/YUSED  (
    .I(\CHOICE4602/GROM ),
    .O(CHOICE4603)
  );
  defparam DLX_IDinst__n01451.INIT = 16'h5000;
  X_LUT4 DLX_IDinst__n01451 (
    .ADR0(DLX_IDinst__n0004),
    .ADR1(VCC),
    .ADR2(DLX_IDinst__n0315),
    .ADR3(DLX_MEMinst_reg_write_MEM),
    .O(\DLX_IDinst__n0145/FROM )
  );
  defparam DLX_IDinst__n01361.INIT = 16'h5500;
  X_LUT4 DLX_IDinst__n01361 (
    .ADR0(DLX_IDinst__n0004),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst__n0075),
    .O(\DLX_IDinst__n0145/GROM )
  );
  X_BUF \DLX_IDinst__n0145/XUSED  (
    .I(\DLX_IDinst__n0145/FROM ),
    .O(DLX_IDinst__n0145)
  );
  X_BUF \DLX_IDinst__n0145/YUSED  (
    .I(\DLX_IDinst__n0145/GROM ),
    .O(DLX_IDinst__n0136)
  );
  defparam DLX_IDinst__n01441.INIT = 16'h00A0;
  X_LUT4 DLX_IDinst__n01441 (
    .ADR0(DLX_MEMinst_reg_write_MEM),
    .ADR1(VCC),
    .ADR2(DLX_IDinst__n0314),
    .ADR3(DLX_IDinst__n0002),
    .O(\DLX_IDinst__n0144/FROM )
  );
  defparam \DLX_IDinst_regA_eff<30>1 .INIT = 16'hF022;
  X_LUT4 \DLX_IDinst_regA_eff<30>1  (
    .ADR0(DLX_IDinst_reg_out_A_RF[30]),
    .ADR1(DLX_IDinst__n0002),
    .ADR2(DLX_MEMinst_RF_data_in[30]),
    .ADR3(DLX_IDinst__n0144),
    .O(\DLX_IDinst__n0144/GROM )
  );
  X_BUF \DLX_IDinst__n0144/XUSED  (
    .I(\DLX_IDinst__n0144/FROM ),
    .O(DLX_IDinst__n0144)
  );
  X_BUF \DLX_IDinst__n0144/YUSED  (
    .I(\DLX_IDinst__n0144/GROM ),
    .O(DLX_IDinst_regA_eff[30])
  );
  defparam \DLX_IDinst__n0086<12>25 .INIT = 16'hFF02;
  X_LUT4 \DLX_IDinst__n0086<12>25  (
    .ADR0(CHOICE2690),
    .ADR1(DLX_IDinst__n0364),
    .ADR2(DLX_IDinst_N70918),
    .ADR3(CHOICE2694),
    .O(\DLX_IDinst_branch_address<12>/FROM )
  );
  defparam \DLX_IDinst__n0086<12>31 .INIT = 16'hFFC0;
  X_LUT4 \DLX_IDinst__n0086<12>31  (
    .ADR0(VCC),
    .ADR1(N100609),
    .ADR2(DLX_IDinst__n0128[12]),
    .ADR3(CHOICE2695),
    .O(N105850)
  );
  X_BUF \DLX_IDinst_branch_address<12>/XUSED  (
    .I(\DLX_IDinst_branch_address<12>/FROM ),
    .O(CHOICE2695)
  );
  defparam DLX_EXlc_md_mda37_a1.INIT = 16'h0C0C;
  X_LUT4 DLX_EXlc_md_mda37_a1 (
    .ADR0(VCC),
    .ADR1(DLX_EXlc_md_wint36),
    .ADR2(DLX_EXlc_pd_wint5),
    .ADR3(VCC),
    .O(\DLX_EXlc_md_wint37/FROM )
  );
  defparam DLX_EXlc_md_mda16_a1.INIT = 16'h00AA;
  X_LUT4 DLX_EXlc_md_mda16_a1 (
    .ADR0(DLX_EXlc_md_wint15),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_EXlc_pd_wint5),
    .O(\DLX_EXlc_md_wint37/GROM )
  );
  X_BUF \DLX_EXlc_md_wint37/XUSED  (
    .I(\DLX_EXlc_md_wint37/FROM ),
    .O(DLX_EXlc_md_wint37)
  );
  X_BUF \DLX_EXlc_md_wint37/YUSED  (
    .I(\DLX_EXlc_md_wint37/GROM ),
    .O(DLX_EXlc_md_wint16)
  );
  defparam \DLX_IDinst__n0086<20>25 .INIT = 16'hCDCC;
  X_LUT4 \DLX_IDinst__n0086<20>25  (
    .ADR0(DLX_IDinst_N70918),
    .ADR1(CHOICE2782),
    .ADR2(DLX_IDinst__n0364),
    .ADR3(CHOICE2778),
    .O(\DLX_IDinst_branch_address<20>/FROM )
  );
  defparam \DLX_IDinst__n0086<20>31 .INIT = 16'hFFA0;
  X_LUT4 \DLX_IDinst__n0086<20>31  (
    .ADR0(N100609),
    .ADR1(VCC),
    .ADR2(DLX_IDinst__n0128[20]),
    .ADR3(CHOICE2783),
    .O(N106354)
  );
  X_BUF \DLX_IDinst_branch_address<20>/XUSED  (
    .I(\DLX_IDinst_branch_address<20>/FROM ),
    .O(CHOICE2783)
  );
  defparam \DLX_EXinst__n0006<9>280 .INIT = 16'hAE00;
  X_LUT4 \DLX_EXinst__n0006<9>280  (
    .ADR0(CHOICE4603),
    .ADR1(CHOICE4570),
    .ADR2(DLX_EXinst__n0030_1),
    .ADR3(DLX_EXinst__n0149),
    .O(\DLX_EXinst_ALU_result<9>/FROM )
  );
  defparam \DLX_EXinst__n0006<9>290 .INIT = 16'hFFF0;
  X_LUT4 \DLX_EXinst__n0006<9>290  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N63689),
    .ADR3(CHOICE4605),
    .O(\DLX_EXinst_ALU_result<9>/GROM )
  );
  X_BUF \DLX_EXinst_ALU_result<9>/XUSED  (
    .I(\DLX_EXinst_ALU_result<9>/FROM ),
    .O(CHOICE4605)
  );
  X_BUF \DLX_EXinst_ALU_result<9>/YUSED  (
    .I(\DLX_EXinst_ALU_result<9>/GROM ),
    .O(N117154)
  );
  defparam DLX_RF_delay_inst_wint61.INIT = 16'h00FF;
  X_LUT4 DLX_RF_delay_inst_wint61 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_RF_delay_inst_wint5),
    .O(\DLX_RF_delay_inst_wint6/GROM )
  );
  X_BUF \DLX_RF_delay_inst_wint6/YUSED  (
    .I(\DLX_RF_delay_inst_wint6/GROM ),
    .O(DLX_RF_delay_inst_wint6)
  );
  defparam DLX_IDinst_Ker709161_1_1179.INIT = 16'h4000;
  X_LUT4 DLX_IDinst_Ker709161_1_1179 (
    .ADR0(DLX_IDinst_IR_latched[28]),
    .ADR1(DLX_IDinst_N70909),
    .ADR2(DLX_IDinst_IR_latched[27]),
    .ADR3(DLX_IDinst_IR_latched[26]),
    .O(\DLX_IDinst_Ker709161_1/FROM )
  );
  defparam DLX_IDinst_Mmux__n0151_Result.INIT = 16'hAEA2;
  X_LUT4 DLX_IDinst_Mmux__n0151_Result (
    .ADR0(N95818),
    .ADR1(DLX_IDinst__n0387),
    .ADR2(DLX_IDinst__n0331),
    .ADR3(DLX_IDinst_Ker709161_1),
    .O(\DLX_IDinst_Ker709161_1/GROM )
  );
  X_BUF \DLX_IDinst_Ker709161_1/XUSED  (
    .I(\DLX_IDinst_Ker709161_1/FROM ),
    .O(DLX_IDinst_Ker709161_1)
  );
  X_BUF \DLX_IDinst_Ker709161_1/YUSED  (
    .I(\DLX_IDinst_Ker709161_1/GROM ),
    .O(DLX_IDinst__n0151)
  );
  defparam DLX_RF_delay_inst_wint71.INIT = 16'h00FF;
  X_LUT4 DLX_RF_delay_inst_wint71 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_RF_delay_inst_wint6),
    .O(\DLX_RF_delay_inst_wint7/GROM )
  );
  X_BUF \DLX_RF_delay_inst_wint7/YUSED  (
    .I(\DLX_RF_delay_inst_wint7/GROM ),
    .O(DLX_RF_delay_inst_wint7)
  );
  defparam DLX_RF_delay_inst_wint81.INIT = 16'h3333;
  X_LUT4 DLX_RF_delay_inst_wint81 (
    .ADR0(VCC),
    .ADR1(DLX_RF_delay_inst_wint7),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_RF_delay_inst_wint8/GROM )
  );
  X_BUF \DLX_RF_delay_inst_wint8/YUSED  (
    .I(\DLX_RF_delay_inst_wint8/GROM ),
    .O(DLX_RF_delay_inst_wint8)
  );
  defparam DLX_IDinst__n01471.INIT = 16'h0010;
  X_LUT4 DLX_IDinst__n01471 (
    .ADR0(DLX_opcode_of_WB[4]),
    .ADR1(DLX_opcode_of_WB[3]),
    .ADR2(DLX_opcode_of_WB[5]),
    .ADR3(DLX_opcode_of_WB[1]),
    .O(\DLX_IDinst__n0147/FROM )
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<31>1 .INIT = 16'h50CC;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<31>1  (
    .ADR0(DLX_opcode_of_WB[2]),
    .ADR1(DLX_MEMinst_RF_data_in[31]),
    .ADR2(DLX_IDinst_Mmux__n0148__net123),
    .ADR3(DLX_IDinst__n0147),
    .O(\DLX_IDinst__n0147/GROM )
  );
  X_BUF \DLX_IDinst__n0147/XUSED  (
    .I(\DLX_IDinst__n0147/FROM ),
    .O(DLX_IDinst__n0147)
  );
  X_BUF \DLX_IDinst__n0147/YUSED  (
    .I(\DLX_IDinst__n0147/GROM ),
    .O(DLX_IDinst_WB_data_eff[31])
  );
  defparam DLX_IDinst_Ker70883_SW0.INIT = 16'hF6F0;
  X_LUT4 DLX_IDinst_Ker70883_SW0 (
    .ADR0(DLX_IDinst_IR_latched[30]),
    .ADR1(DLX_IDinst_IR_latched[27]),
    .ADR2(DLX_IDinst_N70918),
    .ADR3(DLX_IDinst_N70991),
    .O(\N90255/FROM )
  );
  defparam DLX_IDinst__n01631.INIT = 16'h1100;
  X_LUT4 DLX_IDinst__n01631 (
    .ADR0(DLX_IDinst_IR_latched[30]),
    .ADR1(DLX_IDinst_IR_latched[27]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_N70991),
    .O(\N90255/GROM )
  );
  X_BUF \N90255/XUSED  (
    .I(\N90255/FROM ),
    .O(N90255)
  );
  X_BUF \N90255/YUSED  (
    .I(\N90255/GROM ),
    .O(DLX_IDinst__n0448[1])
  );
  defparam DLX_RF_delay_inst_wint91.INIT = 16'h0F0F;
  X_LUT4 DLX_RF_delay_inst_wint91 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_RF_delay_inst_wint8),
    .ADR3(VCC),
    .O(\DLX_RF_delay_inst_wint9/GROM )
  );
  X_BUF \DLX_RF_delay_inst_wint9/YUSED  (
    .I(\DLX_RF_delay_inst_wint9/GROM ),
    .O(DLX_RF_delay_inst_wint9)
  );
  defparam \DLX_IDinst__n0086<21>25 .INIT = 16'hAABA;
  X_LUT4 \DLX_IDinst__n0086<21>25  (
    .ADR0(CHOICE2804),
    .ADR1(DLX_IDinst__n0364),
    .ADR2(CHOICE2800),
    .ADR3(DLX_IDinst_N70918),
    .O(\DLX_IDinst_branch_address<21>/FROM )
  );
  defparam \DLX_IDinst__n0086<21>31 .INIT = 16'hFFC0;
  X_LUT4 \DLX_IDinst__n0086<21>31  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst__n0128[21]),
    .ADR2(N100609),
    .ADR3(CHOICE2805),
    .O(N106480)
  );
  X_BUF \DLX_IDinst_branch_address<21>/XUSED  (
    .I(\DLX_IDinst_branch_address<21>/FROM ),
    .O(CHOICE2805)
  );
  defparam \DLX_IDinst__n0086<13>25 .INIT = 16'hFF10;
  X_LUT4 \DLX_IDinst__n0086<13>25  (
    .ADR0(DLX_IDinst__n0364),
    .ADR1(DLX_IDinst_N70918),
    .ADR2(CHOICE2701),
    .ADR3(CHOICE2705),
    .O(\DLX_IDinst_branch_address<13>/FROM )
  );
  defparam \DLX_IDinst__n0086<13>31 .INIT = 16'hFFC0;
  X_LUT4 \DLX_IDinst__n0086<13>31  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst__n0128[13]),
    .ADR2(N100609),
    .ADR3(CHOICE2706),
    .O(N105913)
  );
  X_BUF \DLX_IDinst_branch_address<13>/XUSED  (
    .I(\DLX_IDinst_branch_address<13>/FROM ),
    .O(CHOICE2706)
  );
  defparam DLX_IDlc_md_mda33_a1.INIT = 16'h5500;
  X_LUT4 DLX_IDlc_md_mda33_a1 (
    .ADR0(DLX_IDlc_pd_wint1),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDlc_md_wint32),
    .O(\DLX_IDlc_md_wint33/FROM )
  );
  defparam DLX_IDlc_ridp31.INIT = 16'h5555;
  X_LUT4 DLX_IDlc_ridp31 (
    .ADR0(DLX_IDlc_pd_wint1),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IDlc_md_wint33/GROM )
  );
  X_BUF \DLX_IDlc_md_wint33/XUSED  (
    .I(\DLX_IDlc_md_wint33/FROM ),
    .O(DLX_IDlc_md_wint33)
  );
  X_BUF \DLX_IDlc_md_wint33/YUSED  (
    .I(\DLX_IDlc_md_wint33/GROM ),
    .O(DLX_IDlc_ridp3)
  );
  defparam DLX_EXinst_Ker6489726.INIT = 16'h00E4;
  X_LUT4 DLX_EXinst_Ker6489726 (
    .ADR0(DLX_IDinst_reg_out_B_3_1),
    .ADR1(DLX_EXinst_N63785),
    .ADR2(DLX_EXinst_N63046),
    .ADR3(DLX_IDinst_reg_out_B[0]),
    .O(\CHOICE1168/FROM )
  );
  defparam DLX_EXinst_Ker6489728.INIT = 16'hFFF0;
  X_LUT4 DLX_EXinst_Ker6489728 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(CHOICE1162),
    .ADR3(CHOICE1168),
    .O(\CHOICE1168/GROM )
  );
  X_BUF \CHOICE1168/XUSED  (
    .I(\CHOICE1168/FROM ),
    .O(CHOICE1168)
  );
  X_BUF \CHOICE1168/YUSED  (
    .I(\CHOICE1168/GROM ),
    .O(N96945)
  );
  defparam DLX_IDinst_Ker6995577.INIT = 16'h3F7F;
  X_LUT4 DLX_IDinst_Ker6995577 (
    .ADR0(DLX_IDinst_IR_opcode_field[1]),
    .ADR1(DLX_IDinst_IR_opcode_field[2]),
    .ADR2(DLX_IDinst_IR_opcode_field[4]),
    .ADR3(DLX_IDinst_IR_opcode_field[0]),
    .O(\CHOICE1436/FROM )
  );
  defparam DLX_EXinst__n0030_SW0.INIT = 16'hFFEE;
  X_LUT4 DLX_EXinst__n0030_SW0 (
    .ADR0(DLX_IDinst_IR_opcode_field[4]),
    .ADR1(DLX_IDinst_IR_opcode_field[3]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_IR_opcode_field[2]),
    .O(\CHOICE1436/GROM )
  );
  X_BUF \CHOICE1436/XUSED  (
    .I(\CHOICE1436/FROM ),
    .O(CHOICE1436)
  );
  X_BUF \CHOICE1436/YUSED  (
    .I(\CHOICE1436/GROM ),
    .O(N95411)
  );
  defparam DLX_IDinst__n01731.INIT = 16'h0300;
  X_LUT4 DLX_IDinst__n01731 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_slot_num_FFd1),
    .ADR2(DLX_IDinst_slot_num_FFd3),
    .ADR3(DLX_IDinst_slot_num_FFd2),
    .O(\DLX_IDinst__n0173/FROM )
  );
  defparam DLX_IDinst__n0440_SW0.INIT = 16'hF505;
  X_LUT4 DLX_IDinst__n0440_SW0 (
    .ADR0(FREEZE_IBUF),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_delay_slot),
    .ADR3(DLX_IDinst__n0173),
    .O(\DLX_IDinst__n0173/GROM )
  );
  X_BUF \DLX_IDinst__n0173/XUSED  (
    .I(\DLX_IDinst__n0173/FROM ),
    .O(DLX_IDinst__n0173)
  );
  X_BUF \DLX_IDinst__n0173/YUSED  (
    .I(\DLX_IDinst__n0173/GROM ),
    .O(N95693)
  );
  defparam \DLX_IDinst__n0086<19>20 .INIT = 16'hAA00;
  X_LUT4 \DLX_IDinst__n0086<19>20  (
    .ADR0(DLX_IDinst_N70295),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_regA_eff[19]),
    .O(\CHOICE2760/FROM )
  );
  defparam \DLX_IDinst__n0086<30>20 .INIT = 16'hF000;
  X_LUT4 \DLX_IDinst__n0086<30>20  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_N70295),
    .ADR3(DLX_IDinst_regA_eff[30]),
    .O(\CHOICE2760/GROM )
  );
  X_BUF \CHOICE2760/XUSED  (
    .I(\CHOICE2760/FROM ),
    .O(CHOICE2760)
  );
  X_BUF \CHOICE2760/YUSED  (
    .I(\CHOICE2760/GROM ),
    .O(CHOICE2793)
  );
  defparam DLX_EXinst__n000533_SW0.INIT = 16'hCFFF;
  X_LUT4 DLX_EXinst__n000533_SW0 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_IR_function_field[0]),
    .ADR2(CHOICE2008),
    .ADR3(DLX_EXinst__n0030),
    .O(\DLX_EXinst_noop/FROM )
  );
  defparam DLX_EXinst__n000533.INIT = 16'hEEEF;
  X_LUT4 DLX_EXinst__n000533 (
    .ADR0(DLX_IDinst_counter[1]),
    .ADR1(DLX_IDinst_counter[0]),
    .ADR2(DLX_IDinst_IR_function_field[5]),
    .ADR3(N127196),
    .O(N101911)
  );
  X_BUF \DLX_EXinst_noop/XUSED  (
    .I(\DLX_EXinst_noop/FROM ),
    .O(N127196)
  );
  defparam DLX_IDinst__n03501.INIT = 16'hEECC;
  X_LUT4 DLX_IDinst__n03501 (
    .ADR0(N100686),
    .ADR1(N98806),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_N70663),
    .O(\DLX_IDinst__n0350/FROM )
  );
  defparam DLX_IDinst_Ker709221.INIT = 16'h0030;
  X_LUT4 DLX_IDinst_Ker709221 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst__n0004),
    .ADR2(DLX_IDinst__n0078),
    .ADR3(DLX_IDinst__n0350),
    .O(\DLX_IDinst__n0350/GROM )
  );
  X_BUF \DLX_IDinst__n0350/XUSED  (
    .I(\DLX_IDinst__n0350/FROM ),
    .O(DLX_IDinst__n0350)
  );
  X_BUF \DLX_IDinst__n0350/YUSED  (
    .I(\DLX_IDinst__n0350/GROM ),
    .O(DLX_IDinst_N70924)
  );
  defparam DLX_IDinst__n04411.INIT = 16'hFAFF;
  X_LUT4 DLX_IDinst__n04411 (
    .ADR0(DLX_IDinst_stall),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_N70653),
    .ADR3(DLX_IDinst__n0331),
    .O(\DLX_IDinst__n0441/FROM )
  );
  defparam DLX_IDinst__n04221.INIT = 16'hFDF5;
  X_LUT4 DLX_IDinst__n04221 (
    .ADR0(DLX_IDinst_stall),
    .ADR1(DLX_IDinst_delay_slot),
    .ADR2(DLX_IDinst__n0331),
    .ADR3(DLX_IDinst_slot_num_FFd2),
    .O(\DLX_IDinst__n0441/GROM )
  );
  X_BUF \DLX_IDinst__n0441/XUSED  (
    .I(\DLX_IDinst__n0441/FROM ),
    .O(DLX_IDinst__n0441)
  );
  X_BUF \DLX_IDinst__n0441/YUSED  (
    .I(\DLX_IDinst__n0441/GROM ),
    .O(DLX_IDinst__n0422)
  );
  defparam \DLX_EXinst__n0006<0>369_SW0 .INIT = 16'hFFFE;
  X_LUT4 \DLX_EXinst__n0006<0>369_SW0  (
    .ADR0(N127252),
    .ADR1(CHOICE5883),
    .ADR2(CHOICE5877),
    .ADR3(CHOICE5891),
    .O(\N126388/FROM )
  );
  defparam \DLX_EXinst__n0006<0>369 .INIT = 16'hF0E0;
  X_LUT4 \DLX_EXinst__n0006<0>369  (
    .ADR0(CHOICE5871),
    .ADR1(CHOICE5850),
    .ADR2(DLX_EXinst__n0030),
    .ADR3(N126388),
    .O(\N126388/GROM )
  );
  X_BUF \N126388/XUSED  (
    .I(\N126388/FROM ),
    .O(N126388)
  );
  X_BUF \N126388/YUSED  (
    .I(\N126388/GROM ),
    .O(CHOICE5921)
  );
  defparam \DLX_IDinst__n0086<14>25 .INIT = 16'hFF04;
  X_LUT4 \DLX_IDinst__n0086<14>25  (
    .ADR0(DLX_IDinst__n0364),
    .ADR1(CHOICE2712),
    .ADR2(DLX_IDinst_N70918),
    .ADR3(CHOICE2716),
    .O(\DLX_IDinst_branch_address<14>/FROM )
  );
  defparam \DLX_IDinst__n0086<14>31 .INIT = 16'hFF88;
  X_LUT4 \DLX_IDinst__n0086<14>31  (
    .ADR0(DLX_IDinst__n0128[14]),
    .ADR1(N100609),
    .ADR2(VCC),
    .ADR3(CHOICE2717),
    .O(N105976)
  );
  X_BUF \DLX_IDinst_branch_address<14>/XUSED  (
    .I(\DLX_IDinst_branch_address<14>/FROM ),
    .O(CHOICE2717)
  );
  defparam \DLX_IDinst__n0086<22>25 .INIT = 16'hF0F4;
  X_LUT4 \DLX_IDinst__n0086<22>25  (
    .ADR0(DLX_IDinst__n0364),
    .ADR1(CHOICE2822),
    .ADR2(CHOICE2826),
    .ADR3(DLX_IDinst_N70918),
    .O(\DLX_IDinst_branch_address<22>/FROM )
  );
  defparam \DLX_IDinst__n0086<22>31 .INIT = 16'hFFA0;
  X_LUT4 \DLX_IDinst__n0086<22>31  (
    .ADR0(N100609),
    .ADR1(VCC),
    .ADR2(DLX_IDinst__n0128[22]),
    .ADR3(CHOICE2827),
    .O(N106606)
  );
  X_BUF \DLX_IDinst_branch_address<22>/XUSED  (
    .I(\DLX_IDinst_branch_address<22>/FROM ),
    .O(CHOICE2827)
  );
  defparam \DLX_IDinst__n0086<30>25 .INIT = 16'hCCCE;
  X_LUT4 \DLX_IDinst__n0086<30>25  (
    .ADR0(CHOICE2789),
    .ADR1(CHOICE2793),
    .ADR2(DLX_IDinst_N70918),
    .ADR3(DLX_IDinst__n0364),
    .O(\DLX_IDinst_branch_address<30>/FROM )
  );
  defparam \DLX_IDinst__n0086<30>31 .INIT = 16'hFF88;
  X_LUT4 \DLX_IDinst__n0086<30>31  (
    .ADR0(DLX_IDinst__n0128[30]),
    .ADR1(N100609),
    .ADR2(VCC),
    .ADR3(CHOICE2794),
    .O(N106417)
  );
  X_BUF \DLX_IDinst_branch_address<30>/XUSED  (
    .I(\DLX_IDinst_branch_address<30>/FROM ),
    .O(CHOICE2794)
  );
  defparam DLX_IDinst__n03441.INIT = 16'hF8F8;
  X_LUT4 DLX_IDinst__n03441 (
    .ADR0(DLX_IDinst_N70647),
    .ADR1(N100686),
    .ADR2(N98613),
    .ADR3(VCC),
    .O(\DLX_IDinst__n0344/FROM )
  );
  defparam DLX_IDinst__n012022.INIT = 16'h0A00;
  X_LUT4 DLX_IDinst__n012022 (
    .ADR0(DLX_IDinst__n0075),
    .ADR1(VCC),
    .ADR2(DLX_IDinst__n0004),
    .ADR3(DLX_IDinst__n0344),
    .O(\DLX_IDinst__n0344/GROM )
  );
  X_BUF \DLX_IDinst__n0344/XUSED  (
    .I(\DLX_IDinst__n0344/FROM ),
    .O(DLX_IDinst__n0344)
  );
  X_BUF \DLX_IDinst__n0344/YUSED  (
    .I(\DLX_IDinst__n0344/GROM ),
    .O(CHOICE3494)
  );
  defparam DLX_EXlc_md_mda34_a1.INIT = 16'h4444;
  X_LUT4 DLX_EXlc_md_mda34_a1 (
    .ADR0(DLX_EXlc_pd_wint5),
    .ADR1(DLX_EXlc_md_wint33),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_EXlc_md_wint34/FROM )
  );
  defparam DLX_EXlc_md_mda35_a1.INIT = 16'h3300;
  X_LUT4 DLX_EXlc_md_mda35_a1 (
    .ADR0(VCC),
    .ADR1(DLX_EXlc_pd_wint5),
    .ADR2(VCC),
    .ADR3(DLX_EXlc_md_wint34),
    .O(\DLX_EXlc_md_wint34/GROM )
  );
  X_BUF \DLX_EXlc_md_wint34/XUSED  (
    .I(\DLX_EXlc_md_wint34/FROM ),
    .O(DLX_EXlc_md_wint34)
  );
  X_BUF \DLX_EXlc_md_wint34/YUSED  (
    .I(\DLX_EXlc_md_wint34/GROM ),
    .O(DLX_EXlc_md_wint35)
  );
  defparam DLX_EXlc_md_mda26_a1.INIT = 16'h3300;
  X_LUT4 DLX_EXlc_md_mda26_a1 (
    .ADR0(VCC),
    .ADR1(DLX_EXlc_pd_wint5),
    .ADR2(VCC),
    .ADR3(DLX_EXlc_md_wint25),
    .O(\DLX_EXlc_md_wint26/FROM )
  );
  defparam DLX_EXlc_md_mda27_a1.INIT = 16'h3300;
  X_LUT4 DLX_EXlc_md_mda27_a1 (
    .ADR0(VCC),
    .ADR1(DLX_EXlc_pd_wint5),
    .ADR2(VCC),
    .ADR3(DLX_EXlc_md_wint26),
    .O(\DLX_EXlc_md_wint26/GROM )
  );
  X_BUF \DLX_EXlc_md_wint26/XUSED  (
    .I(\DLX_EXlc_md_wint26/FROM ),
    .O(DLX_EXlc_md_wint26)
  );
  X_BUF \DLX_EXlc_md_wint26/YUSED  (
    .I(\DLX_EXlc_md_wint26/GROM ),
    .O(DLX_EXlc_md_wint27)
  );
  defparam \DLX_IDinst__n0086<31>11 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst__n0086<31>11  (
    .ADR0(DLX_IDinst_EPC[31]),
    .ADR1(DLX_IDinst__n0071),
    .ADR2(DLX_IDinst_N70786),
    .ADR3(DLX_IDinst_branch_address[31]),
    .O(\DLX_IDinst_branch_address<31>/FROM )
  );
  defparam \DLX_IDinst__n0086<31>27 .INIT = 16'hAFAE;
  X_LUT4 \DLX_IDinst__n0086<31>27  (
    .ADR0(N127435),
    .ADR1(DLX_IDinst__n0364),
    .ADR2(DLX_IDinst_N70918),
    .ADR3(CHOICE2913),
    .O(N107102)
  );
  X_BUF \DLX_IDinst_branch_address<31>/XUSED  (
    .I(\DLX_IDinst_branch_address<31>/FROM ),
    .O(CHOICE2913)
  );
  defparam \DLX_IDinst__n0117<3>15 .INIT = 16'h0CA0;
  X_LUT4 \DLX_IDinst__n0117<3>15  (
    .ADR0(DLX_IDinst_EPC[3]),
    .ADR1(DLX_IDinst_Cause_Reg[3]),
    .ADR2(DLX_IDinst_regA_index[1]),
    .ADR3(DLX_IDinst_regA_index[0]),
    .O(\CHOICE2182/FROM )
  );
  defparam DLX_IDinst__n03451.INIT = 16'hAA8A;
  X_LUT4 DLX_IDinst__n03451 (
    .ADR0(DLX_IDinst__n0077),
    .ADR1(DLX_IDinst_regA_index[0]),
    .ADR2(DLX_IDinst_N70658),
    .ADR3(DLX_IDinst_regA_index[1]),
    .O(\CHOICE2182/GROM )
  );
  X_BUF \CHOICE2182/XUSED  (
    .I(\CHOICE2182/FROM ),
    .O(CHOICE2182)
  );
  X_BUF \CHOICE2182/YUSED  (
    .I(\CHOICE2182/GROM ),
    .O(DLX_IDinst__n0345)
  );
  defparam \DLX_IDinst__n0086<15>20 .INIT = 16'hCC00;
  X_LUT4 \DLX_IDinst__n0086<15>20  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_regA_eff[15]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_N70295),
    .O(\CHOICE2727/GROM )
  );
  X_BUF \CHOICE2727/YUSED  (
    .I(\CHOICE2727/GROM ),
    .O(CHOICE2727)
  );
  defparam \DLX_EXinst_Mshift__n0027_Sh<7>1 .INIT = 16'hCFC0;
  X_LUT4 \DLX_EXinst_Mshift__n0027_Sh<7>1  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N63479),
    .ADR2(DLX_IDinst_IR_function_field_0_1),
    .ADR3(DLX_EXinst_N62766),
    .O(\DLX_EXinst_Mshift__n0027_Sh<7>/FROM )
  );
  defparam DLX_EXinst_Ker628291.INIT = 16'hFBC8;
  X_LUT4 DLX_EXinst_Ker628291 (
    .ADR0(CHOICE994),
    .ADR1(DLX_IDinst_IR_function_field[2]),
    .ADR2(CHOICE1000),
    .ADR3(\DLX_EXinst_Mshift__n0027_Sh[7] ),
    .O(\DLX_EXinst_Mshift__n0027_Sh<7>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0027_Sh<7>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0027_Sh<7>/FROM ),
    .O(\DLX_EXinst_Mshift__n0027_Sh[7] )
  );
  X_BUF \DLX_EXinst_Mshift__n0027_Sh<7>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0027_Sh<7>/GROM ),
    .O(DLX_EXinst_N62831)
  );
  defparam DLX_IDinst__n00886.INIT = 16'hEA00;
  X_LUT4 DLX_IDinst__n00886 (
    .ADR0(DLX_IDinst__n0250),
    .ADR1(DLX_IDinst_N70635),
    .ADR2(DLX_IDinst__n0377),
    .ADR3(DLX_IDinst_N70909),
    .O(\CHOICE3466/FROM )
  );
  defparam DLX_IDinst__n008827.INIT = 16'hE0C0;
  X_LUT4 DLX_IDinst__n008827 (
    .ADR0(DLX_IDinst_N70985),
    .ADR1(CHOICE3470),
    .ADR2(DLX_IDinst_N69568),
    .ADR3(CHOICE3466),
    .O(\CHOICE3466/GROM )
  );
  X_BUF \CHOICE3466/XUSED  (
    .I(\CHOICE3466/FROM ),
    .O(CHOICE3466)
  );
  X_BUF \CHOICE3466/YUSED  (
    .I(\CHOICE3466/GROM ),
    .O(CHOICE3472)
  );
  defparam DLX_IFlc_ridp31.INIT = 16'h3333;
  X_LUT4 DLX_IFlc_ridp31 (
    .ADR0(VCC),
    .ADR1(DLX_IFlc_ridp2),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IFlc_ridp3/GROM )
  );
  X_BUF \DLX_IFlc_ridp3/YUSED  (
    .I(\DLX_IFlc_ridp3/GROM ),
    .O(DLX_IFlc_ridp3)
  );
  defparam \DLX_IDinst__n0086<23>25 .INIT = 16'hAAAE;
  X_LUT4 \DLX_IDinst__n0086<23>25  (
    .ADR0(CHOICE2815),
    .ADR1(CHOICE2811),
    .ADR2(DLX_IDinst__n0364),
    .ADR3(DLX_IDinst_N70918),
    .O(\DLX_IDinst_branch_address<23>/FROM )
  );
  defparam \DLX_IDinst__n0086<23>31 .INIT = 16'hFF88;
  X_LUT4 \DLX_IDinst__n0086<23>31  (
    .ADR0(DLX_IDinst__n0128[23]),
    .ADR1(N100609),
    .ADR2(VCC),
    .ADR3(CHOICE2816),
    .O(N106543)
  );
  X_BUF \DLX_IDinst_branch_address<23>/XUSED  (
    .I(\DLX_IDinst_branch_address<23>/FROM ),
    .O(CHOICE2816)
  );
  defparam \DLX_IDinst__n0086<15>25 .INIT = 16'hFF04;
  X_LUT4 \DLX_IDinst__n0086<15>25  (
    .ADR0(DLX_IDinst__n0364),
    .ADR1(CHOICE2723),
    .ADR2(DLX_IDinst_N70918),
    .ADR3(CHOICE2727),
    .O(\DLX_IDinst_branch_address<15>/FROM )
  );
  defparam \DLX_IDinst__n0086<15>31 .INIT = 16'hFF88;
  X_LUT4 \DLX_IDinst__n0086<15>31  (
    .ADR0(DLX_IDinst__n0128[15]),
    .ADR1(N100609),
    .ADR2(VCC),
    .ADR3(CHOICE2728),
    .O(N106039)
  );
  X_BUF \DLX_IDinst_branch_address<15>/XUSED  (
    .I(\DLX_IDinst_branch_address<15>/FROM ),
    .O(CHOICE2728)
  );
  defparam DLX_IDinst__n03481.INIT = 16'h5500;
  X_LUT4 DLX_IDinst__n03481 (
    .ADR0(DLX_IDinst__n0004),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst__n0078),
    .O(\DLX_IDinst__n0348/FROM )
  );
  defparam DLX_IDinst_Ker6960415.INIT = 16'h0037;
  X_LUT4 DLX_IDinst_Ker6960415 (
    .ADR0(DLX_IDinst__n0250),
    .ADR1(DLX_IDinst_N70909),
    .ADR2(DLX_IDinst_N70635),
    .ADR3(DLX_IDinst__n0348),
    .O(\DLX_IDinst__n0348/GROM )
  );
  X_BUF \DLX_IDinst__n0348/XUSED  (
    .I(\DLX_IDinst__n0348/FROM ),
    .O(DLX_IDinst__n0348)
  );
  X_BUF \DLX_IDinst__n0348/YUSED  (
    .I(\DLX_IDinst__n0348/GROM ),
    .O(CHOICE2093)
  );
  defparam DLX_IDinst__n03641.INIT = 16'hF0F2;
  X_LUT4 DLX_IDinst__n03641 (
    .ADR0(INT_IBUF),
    .ADR1(DLX_IDinst_CLI),
    .ADR2(DLX_IDinst__n0070),
    .ADR3(DLX_IDinst_delay_slot),
    .O(\DLX_IDinst__n0364/FROM )
  );
  defparam DLX_IDinst__n010875.INIT = 16'hFFA8;
  X_LUT4 DLX_IDinst__n010875 (
    .ADR0(DLX_IDinst_N69781),
    .ADR1(CHOICE3445),
    .ADR2(CHOICE3436),
    .ADR3(DLX_IDinst__n0364),
    .O(\DLX_IDinst__n0364/GROM )
  );
  X_BUF \DLX_IDinst__n0364/XUSED  (
    .I(\DLX_IDinst__n0364/FROM ),
    .O(DLX_IDinst__n0364)
  );
  X_BUF \DLX_IDinst__n0364/YUSED  (
    .I(\DLX_IDinst__n0364/GROM ),
    .O(CHOICE3448)
  );
  defparam \DLX_EXinst_Mshift__n0027_Sh<9>1 .INIT = 16'hEE44;
  X_LUT4 \DLX_EXinst_Mshift__n0027_Sh<9>1  (
    .ADR0(DLX_IDinst_IR_function_field_0_1),
    .ADR1(DLX_EXinst_N62771),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N63484),
    .O(\DLX_EXinst_Mshift__n0027_Sh<9>/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0027_Sh<41>_SW1 .INIT = 16'h101F;
  X_LUT4 \DLX_EXinst_Mshift__n0027_Sh<41>_SW1  (
    .ADR0(CHOICE1024),
    .ADR1(CHOICE1018),
    .ADR2(DLX_IDinst_IR_function_field_2_1),
    .ADR3(\DLX_EXinst_Mshift__n0027_Sh[9] ),
    .O(\DLX_EXinst_Mshift__n0027_Sh<9>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0027_Sh<9>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0027_Sh<9>/FROM ),
    .O(\DLX_EXinst_Mshift__n0027_Sh[9] )
  );
  X_BUF \DLX_EXinst_Mshift__n0027_Sh<9>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0027_Sh<9>/GROM ),
    .O(N127149)
  );
  defparam \DLX_IDinst__n0086<16>25 .INIT = 16'hF0F4;
  X_LUT4 \DLX_IDinst__n0086<16>25  (
    .ADR0(DLX_IDinst_N70918),
    .ADR1(CHOICE2734),
    .ADR2(CHOICE2738),
    .ADR3(DLX_IDinst__n0364),
    .O(\DLX_IDinst_branch_address<16>/FROM )
  );
  defparam \DLX_IDinst__n0086<16>31 .INIT = 16'hFFC0;
  X_LUT4 \DLX_IDinst__n0086<16>31  (
    .ADR0(VCC),
    .ADR1(N100609),
    .ADR2(DLX_IDinst__n0128[16]),
    .ADR3(CHOICE2739),
    .O(N106102)
  );
  X_BUF \DLX_IDinst_branch_address<16>/XUSED  (
    .I(\DLX_IDinst_branch_address<16>/FROM ),
    .O(CHOICE2739)
  );
  defparam \DLX_IDinst__n0086<24>25 .INIT = 16'hF1F0;
  X_LUT4 \DLX_IDinst__n0086<24>25  (
    .ADR0(DLX_IDinst_N70918),
    .ADR1(DLX_IDinst__n0364),
    .ADR2(CHOICE2837),
    .ADR3(CHOICE2833),
    .O(\DLX_IDinst_branch_address<24>/FROM )
  );
  defparam \DLX_IDinst__n0086<24>31 .INIT = 16'hFFA0;
  X_LUT4 \DLX_IDinst__n0086<24>31  (
    .ADR0(N100609),
    .ADR1(VCC),
    .ADR2(DLX_IDinst__n0128[24]),
    .ADR3(CHOICE2838),
    .O(N106669)
  );
  X_BUF \DLX_IDinst_branch_address<24>/XUSED  (
    .I(\DLX_IDinst_branch_address<24>/FROM ),
    .O(CHOICE2838)
  );
  defparam DLX_IDinst_Ker7003710.INIT = 16'hFF08;
  X_LUT4 DLX_IDinst_Ker7003710 (
    .ADR0(DLX_IDinst_N70991),
    .ADR1(DLX_IDinst_IR_latched[27]),
    .ADR2(DLX_IDinst__n03641_1),
    .ADR3(DLX_IDinst_N70918),
    .O(\CHOICE1786/FROM )
  );
  defparam DLX_IDinst__n04561.INIT = 16'h0F08;
  X_LUT4 DLX_IDinst__n04561 (
    .ADR0(DLX_IDinst_IR_latched[27]),
    .ADR1(DLX_IDinst_N70991),
    .ADR2(DLX_IDinst_IR_latched[30]),
    .ADR3(DLX_IDinst_N70918),
    .O(\CHOICE1786/GROM )
  );
  X_BUF \CHOICE1786/XUSED  (
    .I(\CHOICE1786/FROM ),
    .O(CHOICE1786)
  );
  X_BUF \CHOICE1786/YUSED  (
    .I(\CHOICE1786/GROM ),
    .O(DLX_IDinst__n0456)
  );
  defparam DLX_EXlc_pd_wint21.INIT = 16'h0F0F;
  X_LUT4 DLX_EXlc_pd_wint21 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_EXlc_pd_wint1),
    .ADR3(VCC),
    .O(\DLX_EXlc_pd_wint2/GROM )
  );
  X_BUF \DLX_EXlc_pd_wint2/YUSED  (
    .I(\DLX_EXlc_pd_wint2/GROM ),
    .O(DLX_EXlc_pd_wint2)
  );
  defparam DLX_EXinst__n0030_1_1180.INIT = 16'h0001;
  X_LUT4 DLX_EXinst__n0030_1_1180 (
    .ADR0(DLX_IDinst_IR_opcode_field[5]),
    .ADR1(DLX_IDinst_IR_opcode_field[1]),
    .ADR2(DLX_IDinst_IR_opcode_field[0]),
    .ADR3(N95411),
    .O(\DLX_EXinst__n0030_1/FROM )
  );
  defparam DLX_EXinst_Ker66070_SW0.INIT = 16'hF0FF;
  X_LUT4 DLX_EXinst_Ker66070_SW0 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B_2_1),
    .ADR3(DLX_EXinst__n0030_1),
    .O(\DLX_EXinst__n0030_1/GROM )
  );
  X_BUF \DLX_EXinst__n0030_1/XUSED  (
    .I(\DLX_EXinst__n0030_1/FROM ),
    .O(DLX_EXinst__n0030_1)
  );
  X_BUF \DLX_EXinst__n0030_1/YUSED  (
    .I(\DLX_EXinst__n0030_1/GROM ),
    .O(N90062)
  );
  defparam DLX_IDinst_Ker7064058_SW2.INIT = 16'hDF7F;
  X_LUT4 DLX_IDinst_Ker7064058_SW2 (
    .ADR0(DLX_IDinst_IR_latched[28]),
    .ADR1(DLX_IDinst_zflag),
    .ADR2(DLX_IDinst_N70909),
    .ADR3(DLX_IDinst_IR_latched[26]),
    .O(\N127555/FROM )
  );
  defparam DLX_IDinst__n03771.INIT = 16'h2800;
  X_LUT4 DLX_IDinst__n03771 (
    .ADR0(DLX_IDinst_N70635),
    .ADR1(DLX_IDinst_zflag),
    .ADR2(DLX_IDinst_IR_latched[26]),
    .ADR3(DLX_IDinst_N70909),
    .O(\N127555/GROM )
  );
  X_BUF \N127555/XUSED  (
    .I(\N127555/FROM ),
    .O(N127555)
  );
  X_BUF \N127555/YUSED  (
    .I(\N127555/GROM ),
    .O(DLX_IDinst__n0377)
  );
  defparam DLX_EXlc_pd_wint31.INIT = 16'h3333;
  X_LUT4 DLX_EXlc_pd_wint31 (
    .ADR0(VCC),
    .ADR1(DLX_EXlc_pd_wint2),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_EXlc_pd_wint3/GROM )
  );
  X_BUF \DLX_EXlc_pd_wint3/YUSED  (
    .I(\DLX_EXlc_pd_wint3/GROM ),
    .O(DLX_EXlc_pd_wint3)
  );
  defparam DLX_EXlc_pd_wint41.INIT = 16'h3333;
  X_LUT4 DLX_EXlc_pd_wint41 (
    .ADR0(VCC),
    .ADR1(DLX_EXlc_pd_wint3),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_EXlc_pd_wint4/GROM )
  );
  X_BUF \DLX_EXlc_pd_wint4/YUSED  (
    .I(\DLX_EXlc_pd_wint4/GROM ),
    .O(DLX_EXlc_pd_wint4)
  );
  defparam DLX_IDinst__n03871.INIT = 16'h88F8;
  X_LUT4 DLX_IDinst__n03871 (
    .ADR0(DLX_IDinst_slot_num_FFd2),
    .ADR1(DLX_IDinst_delay_slot),
    .ADR2(DLX_EXinst__n0149),
    .ADR3(DLX_IDinst_stall),
    .O(\DLX_IDinst_stall/FROM )
  );
  defparam DLX_IDinst__n0120111.INIT = 16'hF888;
  X_LUT4 DLX_IDinst__n0120111 (
    .ADR0(DLX_IDinst__n0331),
    .ADR1(DLX_IDinst_N70653),
    .ADR2(N126293),
    .ADR3(DLX_IDinst__n0387),
    .O(\DLX_IDinst_stall/GROM )
  );
  X_BUF \DLX_IDinst_stall/XUSED  (
    .I(\DLX_IDinst_stall/FROM ),
    .O(DLX_IDinst__n0387)
  );
  X_BUF \DLX_IDinst_stall/YUSED  (
    .I(\DLX_IDinst_stall/GROM ),
    .O(N110648)
  );
  defparam DLX_EXlc_pd_wint51.INIT = 16'h3333;
  X_LUT4 DLX_EXlc_pd_wint51 (
    .ADR0(VCC),
    .ADR1(DLX_EXlc_pd_wint4),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_EXlc_pd_wint5/FROM )
  );
  defparam DLX_EXlc_md_mda40_a1.INIT = 16'h00CC;
  X_LUT4 DLX_EXlc_md_mda40_a1 (
    .ADR0(VCC),
    .ADR1(DLX_EXlc_md_wint39),
    .ADR2(VCC),
    .ADR3(DLX_EXlc_pd_wint5),
    .O(\DLX_EXlc_pd_wint5/GROM )
  );
  X_BUF \DLX_EXlc_pd_wint5/XUSED  (
    .I(\DLX_EXlc_pd_wint5/FROM ),
    .O(DLX_EXlc_pd_wint5)
  );
  X_BUF \DLX_EXlc_pd_wint5/YUSED  (
    .I(\DLX_EXlc_pd_wint5/GROM ),
    .O(DLX_EXlc_md_wint40)
  );
  defparam \DLX_IDinst__n0086<17>25 .INIT = 16'hCDCC;
  X_LUT4 \DLX_IDinst__n0086<17>25  (
    .ADR0(DLX_IDinst__n0364),
    .ADR1(CHOICE2749),
    .ADR2(DLX_IDinst_N70918),
    .ADR3(CHOICE2745),
    .O(\DLX_IDinst_branch_address<17>/FROM )
  );
  defparam \DLX_IDinst__n0086<17>31 .INIT = 16'hFFA0;
  X_LUT4 \DLX_IDinst__n0086<17>31  (
    .ADR0(N100609),
    .ADR1(VCC),
    .ADR2(DLX_IDinst__n0128[17]),
    .ADR3(CHOICE2750),
    .O(N106165)
  );
  X_BUF \DLX_IDinst_branch_address<17>/XUSED  (
    .I(\DLX_IDinst_branch_address<17>/FROM ),
    .O(CHOICE2750)
  );
  defparam \DLX_IDinst__n0086<25>25 .INIT = 16'hABAA;
  X_LUT4 \DLX_IDinst__n0086<25>25  (
    .ADR0(CHOICE2859),
    .ADR1(DLX_IDinst_N70918),
    .ADR2(DLX_IDinst__n0364),
    .ADR3(CHOICE2855),
    .O(\DLX_IDinst_branch_address<25>/FROM )
  );
  defparam \DLX_IDinst__n0086<25>31 .INIT = 16'hFFA0;
  X_LUT4 \DLX_IDinst__n0086<25>31  (
    .ADR0(N100609),
    .ADR1(VCC),
    .ADR2(DLX_IDinst__n0128[25]),
    .ADR3(CHOICE2860),
    .O(N106789)
  );
  X_BUF \DLX_IDinst_branch_address<25>/XUSED  (
    .I(\DLX_IDinst_branch_address<25>/FROM ),
    .O(CHOICE2860)
  );
  defparam DLX_EXinst_Ker62713.INIT = 16'hEEE2;
  X_LUT4 DLX_EXinst_Ker62713 (
    .ADR0(N94007),
    .ADR1(DLX_IDinst_IR_function_field[3]),
    .ADR2(CHOICE1126),
    .ADR3(CHOICE1132),
    .O(\DLX_EXinst_N62715/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0028_Sh<52>1 .INIT = 16'h2F20;
  X_LUT4 \DLX_EXinst_Mshift__n0028_Sh<52>1  (
    .ADR0(\DLX_EXinst_Mshift__n0028_Sh[24] ),
    .ADR1(DLX_IDinst_IR_function_field_3_1),
    .ADR2(DLX_IDinst_IR_function_field_2_1),
    .ADR3(DLX_EXinst_N62715),
    .O(\DLX_EXinst_N62715/GROM )
  );
  X_BUF \DLX_EXinst_N62715/XUSED  (
    .I(\DLX_EXinst_N62715/FROM ),
    .O(DLX_EXinst_N62715)
  );
  X_BUF \DLX_EXinst_N62715/YUSED  (
    .I(\DLX_EXinst_N62715/GROM ),
    .O(\DLX_EXinst_Mshift__n0028_Sh[52] )
  );
  defparam \DLX_IFinst__n0001<10>_SW0 .INIT = 16'h4477;
  X_LUT4 \DLX_IFinst__n0001<10>_SW0  (
    .ADR0(DLX_IFinst_PC[10]),
    .ADR1(DLX_IFinst__n0000),
    .ADR2(VCC),
    .ADR3(DLX_IFinst__n0015[10]),
    .O(\DLX_IFinst_NPC<10>/FROM )
  );
  defparam \DLX_IFinst__n0001<10> .INIT = 16'hA0AF;
  X_LUT4 \DLX_IFinst__n0001<10>  (
    .ADR0(DLX_IDinst_branch_address[10]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(N92607),
    .O(\DLX_IFinst_NPC<10>/GROM )
  );
  X_BUF \DLX_IFinst_NPC<10>/XUSED  (
    .I(\DLX_IFinst_NPC<10>/FROM ),
    .O(N92607)
  );
  X_BUF \DLX_IFinst_NPC<10>/YUSED  (
    .I(\DLX_IFinst_NPC<10>/GROM ),
    .O(DLX_IFinst__n0001[10])
  );
  defparam \DLX_IDinst__n0086<26>25 .INIT = 16'hF0F2;
  X_LUT4 \DLX_IDinst__n0086<26>25  (
    .ADR0(CHOICE2866),
    .ADR1(DLX_IDinst_N70918),
    .ADR2(CHOICE2870),
    .ADR3(DLX_IDinst__n0364),
    .O(\DLX_IDinst_branch_address<26>/FROM )
  );
  defparam \DLX_IDinst__n0086<26>31 .INIT = 16'hFFC0;
  X_LUT4 \DLX_IDinst__n0086<26>31  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst__n0128[26]),
    .ADR2(N100609),
    .ADR3(CHOICE2871),
    .O(N106852)
  );
  X_BUF \DLX_IDinst_branch_address<26>/XUSED  (
    .I(\DLX_IDinst_branch_address<26>/FROM ),
    .O(CHOICE2871)
  );
  defparam \DLX_IDinst__n0086<18>25 .INIT = 16'hFF10;
  X_LUT4 \DLX_IDinst__n0086<18>25  (
    .ADR0(DLX_IDinst__n0364),
    .ADR1(DLX_IDinst_N70918),
    .ADR2(CHOICE2767),
    .ADR3(CHOICE2771),
    .O(\DLX_IDinst_branch_address<18>/FROM )
  );
  defparam \DLX_IDinst__n0086<18>31 .INIT = 16'hFF88;
  X_LUT4 \DLX_IDinst__n0086<18>31  (
    .ADR0(N100609),
    .ADR1(DLX_IDinst__n0128[18]),
    .ADR2(VCC),
    .ADR3(CHOICE2772),
    .O(N106291)
  );
  X_BUF \DLX_IDinst_branch_address<18>/XUSED  (
    .I(\DLX_IDinst_branch_address<18>/FROM ),
    .O(CHOICE2772)
  );
  defparam DLX_MEMlc_master_ctrlMEM__n0001_SW19.INIT = 16'hFFF3;
  X_LUT4 DLX_MEMlc_master_ctrlMEM__n0001_SW19 (
    .ADR0(VCC),
    .ADR1(DLX_MEMlc_master_ctrlMEM_nro),
    .ADR2(DLX_MEMlc_master_ctrlMEM_l),
    .ADR3(reset_IBUF_1),
    .O(\CHOICE5/FROM )
  );
  defparam DLX_MEMlc_master_ctrlMEM__n0001_SW111.INIT = 16'h3300;
  X_LUT4 DLX_MEMlc_master_ctrlMEM__n0001_SW111 (
    .ADR0(VCC),
    .ADR1(DLX_MEMlc_md_outp2),
    .ADR2(VCC),
    .ADR3(CHOICE5),
    .O(\CHOICE5/GROM )
  );
  X_BUF \CHOICE5/XUSED  (
    .I(\CHOICE5/FROM ),
    .O(CHOICE5)
  );
  X_BUF \CHOICE5/YUSED  (
    .I(\CHOICE5/GROM ),
    .O(DLX_MEMlc_master_ctrlMEM_l)
  );
  defparam DLX_EXlc_md_mda38_a1.INIT = 16'h2222;
  X_LUT4 DLX_EXlc_md_mda38_a1 (
    .ADR0(DLX_EXlc_md_wint37),
    .ADR1(DLX_EXlc_pd_wint5),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_EXlc_md_wint38/GROM )
  );
  X_BUF \DLX_EXlc_md_wint38/YUSED  (
    .I(\DLX_EXlc_md_wint38/GROM ),
    .O(DLX_EXlc_md_wint38)
  );
  defparam DLX_EXinst_Ker62725.INIT = 16'hEEF0;
  X_LUT4 DLX_EXinst_Ker62725 (
    .ADR0(CHOICE1150),
    .ADR1(CHOICE1156),
    .ADR2(N94057),
    .ADR3(DLX_IDinst_reg_out_B[3]),
    .O(\DLX_EXinst_N62727/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0026_Sh<52>1 .INIT = 16'h2F20;
  X_LUT4 \DLX_EXinst_Mshift__n0026_Sh<52>1  (
    .ADR0(\DLX_EXinst_Mshift__n0026_Sh[24] ),
    .ADR1(DLX_IDinst_reg_out_B_3_1),
    .ADR2(DLX_IDinst_reg_out_B_2_1),
    .ADR3(DLX_EXinst_N62727),
    .O(\DLX_EXinst_N62727/GROM )
  );
  X_BUF \DLX_EXinst_N62727/XUSED  (
    .I(\DLX_EXinst_N62727/FROM ),
    .O(DLX_EXinst_N62727)
  );
  X_BUF \DLX_EXinst_N62727/YUSED  (
    .I(\DLX_EXinst_N62727/GROM ),
    .O(\DLX_EXinst_Mshift__n0026_Sh[52] )
  );
  defparam DLX_EXinst_Ker64179.INIT = 16'hAAEA;
  X_LUT4 DLX_EXinst_Ker64179 (
    .ADR0(N95259),
    .ADR1(DLX_IDinst_reg_out_B[0]),
    .ADR2(DLX_EXinst_N66072),
    .ADR3(DLX_IDinst_reg_out_B[1]),
    .O(\DLX_EXinst_N64181/FROM )
  );
  defparam \DLX_EXinst__n0006<29>350 .INIT = 16'hECA0;
  X_LUT4 \DLX_EXinst__n0006<29>350  (
    .ADR0(DLX_IDinst_reg_out_A[27]),
    .ADR1(DLX_IDinst_reg_out_A[28]),
    .ADR2(DLX_EXinst_N63996),
    .ADR3(DLX_EXinst_N64181),
    .O(\DLX_EXinst_N64181/GROM )
  );
  X_BUF \DLX_EXinst_N64181/XUSED  (
    .I(\DLX_EXinst_N64181/FROM ),
    .O(DLX_EXinst_N64181)
  );
  X_BUF \DLX_EXinst_N64181/YUSED  (
    .I(\DLX_EXinst_N64181/GROM ),
    .O(CHOICE5401)
  );
  defparam \DLX_IDinst__n0086<27>25 .INIT = 16'hFF10;
  X_LUT4 \DLX_IDinst__n0086<27>25  (
    .ADR0(DLX_IDinst_N70918),
    .ADR1(DLX_IDinst__n0364),
    .ADR2(CHOICE2877),
    .ADR3(CHOICE2881),
    .O(\DLX_IDinst_branch_address<27>/FROM )
  );
  defparam \DLX_IDinst__n0086<27>31 .INIT = 16'hFFA0;
  X_LUT4 \DLX_IDinst__n0086<27>31  (
    .ADR0(DLX_IDinst__n0128[27]),
    .ADR1(VCC),
    .ADR2(N100609),
    .ADR3(CHOICE2882),
    .O(N106915)
  );
  X_BUF \DLX_IDinst_branch_address<27>/XUSED  (
    .I(\DLX_IDinst_branch_address<27>/FROM ),
    .O(CHOICE2882)
  );
  defparam \DLX_IDinst__n0086<19>25 .INIT = 16'hFF02;
  X_LUT4 \DLX_IDinst__n0086<19>25  (
    .ADR0(CHOICE2756),
    .ADR1(DLX_IDinst__n0364),
    .ADR2(DLX_IDinst_N70918),
    .ADR3(CHOICE2760),
    .O(\DLX_IDinst_branch_address<19>/FROM )
  );
  defparam \DLX_IDinst__n0086<19>31 .INIT = 16'hFFC0;
  X_LUT4 \DLX_IDinst__n0086<19>31  (
    .ADR0(VCC),
    .ADR1(N100609),
    .ADR2(DLX_IDinst__n0128[19]),
    .ADR3(CHOICE2761),
    .O(N106228)
  );
  X_BUF \DLX_IDinst_branch_address<19>/XUSED  (
    .I(\DLX_IDinst_branch_address<19>/FROM ),
    .O(CHOICE2761)
  );
  defparam DLX_EXlc_md_mda39_a1.INIT = 16'h5050;
  X_LUT4 DLX_EXlc_md_mda39_a1 (
    .ADR0(DLX_EXlc_pd_wint5),
    .ADR1(VCC),
    .ADR2(DLX_EXlc_md_wint38),
    .ADR3(VCC),
    .O(\DLX_EXlc_md_wint39/GROM )
  );
  X_BUF \DLX_EXlc_md_wint39/YUSED  (
    .I(\DLX_EXlc_md_wint39/GROM ),
    .O(DLX_EXlc_md_wint39)
  );
  defparam DLX_EXinst_Ker64446.INIT = 16'h0104;
  X_LUT4 DLX_EXinst_Ker64446 (
    .ADR0(N127412),
    .ADR1(DLX_IDinst_IR_function_field[4]),
    .ADR2(DLX_IDinst_IR_function_field[3]),
    .ADR3(DLX_IDinst_IR_function_field_2_1),
    .O(\DLX_EXinst_N64448/FROM )
  );
  defparam \DLX_EXinst__n0006<29>275 .INIT = 16'hFF88;
  X_LUT4 \DLX_EXinst__n0006<29>275  (
    .ADR0(DLX_EXinst__n0045),
    .ADR1(DLX_IDinst_reg_out_B[29]),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N64448),
    .O(\DLX_EXinst_N64448/GROM )
  );
  X_BUF \DLX_EXinst_N64448/XUSED  (
    .I(\DLX_EXinst_N64448/FROM ),
    .O(DLX_EXinst_N64448)
  );
  X_BUF \DLX_EXinst_N64448/YUSED  (
    .I(\DLX_EXinst_N64448/GROM ),
    .O(CHOICE5390)
  );
  defparam \DLX_EXinst__n0006<27>110_SW0 .INIT = 16'hF222;
  X_LUT4 \DLX_EXinst__n0006<27>110_SW0  (
    .ADR0(CHOICE4633),
    .ADR1(DLX_IDinst_IR_function_field[4]),
    .ADR2(\DLX_IDinst_Imm[11] ),
    .ADR3(DLX_EXinst__n0077),
    .O(\N126428/FROM )
  );
  defparam \DLX_EXinst__n0006<27>110 .INIT = 16'hFFEC;
  X_LUT4 \DLX_EXinst__n0006<27>110  (
    .ADR0(DLX_EXinst__n0128),
    .ADR1(CHOICE4621),
    .ADR2(DLX_EXinst__n0016[27]),
    .ADR3(N126428),
    .O(\N126428/GROM )
  );
  X_BUF \N126428/XUSED  (
    .I(\N126428/FROM ),
    .O(N126428)
  );
  X_BUF \N126428/YUSED  (
    .I(\N126428/GROM ),
    .O(CHOICE4636)
  );
  defparam DLX_IDinst_Ker7003722.INIT = 16'h0A00;
  X_LUT4 DLX_IDinst_Ker7003722 (
    .ADR0(DLX_IDinst_N70885),
    .ADR1(VCC),
    .ADR2(DLX_IDinst__n03641_1),
    .ADR3(DLX_IDinst_N70635),
    .O(\CHOICE1790/FROM )
  );
  defparam DLX_IDinst_Ker7003725.INIT = 16'hFF22;
  X_LUT4 DLX_IDinst_Ker7003725 (
    .ADR0(CHOICE1786),
    .ADR1(DLX_IDinst_IR_latched[30]),
    .ADR2(VCC),
    .ADR3(CHOICE1790),
    .O(\CHOICE1790/GROM )
  );
  X_BUF \CHOICE1790/XUSED  (
    .I(\CHOICE1790/FROM ),
    .O(CHOICE1790)
  );
  X_BUF \CHOICE1790/YUSED  (
    .I(\CHOICE1790/GROM ),
    .O(N100609)
  );
  defparam \DLX_IDinst__n0086<28>25 .INIT = 16'hFF04;
  X_LUT4 \DLX_IDinst__n0086<28>25  (
    .ADR0(DLX_IDinst__n0364),
    .ADR1(CHOICE2888),
    .ADR2(DLX_IDinst_N70918),
    .ADR3(CHOICE2892),
    .O(\DLX_IDinst_branch_address<28>/FROM )
  );
  defparam \DLX_IDinst__n0086<28>31 .INIT = 16'hFFA0;
  X_LUT4 \DLX_IDinst__n0086<28>31  (
    .ADR0(N100609),
    .ADR1(VCC),
    .ADR2(DLX_IDinst__n0128[28]),
    .ADR3(CHOICE2893),
    .O(N106978)
  );
  X_BUF \DLX_IDinst_branch_address<28>/XUSED  (
    .I(\DLX_IDinst_branch_address<28>/FROM ),
    .O(CHOICE2893)
  );
  defparam \DLX_EXinst__n0006<31>163_SW0 .INIT = 16'hF0EE;
  X_LUT4 \DLX_EXinst__n0006<31>163_SW0  (
    .ADR0(CHOICE5764),
    .ADR1(CHOICE5769),
    .ADR2(\DLX_EXinst_Mshift__n0025_Sh[23] ),
    .ADR3(DLX_IDinst_reg_out_B[3]),
    .O(\N126169/FROM )
  );
  defparam DLX_EXinst_Ker63908.INIT = 16'hF3C0;
  X_LUT4 DLX_EXinst_Ker63908 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_B[3]),
    .ADR2(\DLX_EXinst_Mshift__n0025_Sh[9] ),
    .ADR3(N93487),
    .O(\N126169/GROM )
  );
  X_BUF \N126169/XUSED  (
    .I(\N126169/FROM ),
    .O(N126169)
  );
  X_BUF \N126169/YUSED  (
    .I(\N126169/GROM ),
    .O(DLX_EXinst_N63910)
  );
  defparam DLX_EXinst_Ker63687.INIT = 16'hA0A3;
  X_LUT4 DLX_EXinst_Ker63687 (
    .ADR0(N101921),
    .ADR1(DLX_IDinst_IR_function_field[4]),
    .ADR2(DLX_EXinst__n0030_1),
    .ADR3(N101919),
    .O(\DLX_EXinst_ALU_result<14>/FROM )
  );
  defparam \DLX_EXinst__n0006<14>277 .INIT = 16'hFFC8;
  X_LUT4 \DLX_EXinst__n0006<14>277  (
    .ADR0(CHOICE4251),
    .ADR1(DLX_EXinst__n0149),
    .ADR2(CHOICE4283),
    .ADR3(DLX_EXinst_N63689),
    .O(\DLX_EXinst_ALU_result<14>/GROM )
  );
  X_BUF \DLX_EXinst_ALU_result<14>/XUSED  (
    .I(\DLX_EXinst_ALU_result<14>/FROM ),
    .O(DLX_EXinst_N63689)
  );
  X_BUF \DLX_EXinst_ALU_result<14>/YUSED  (
    .I(\DLX_EXinst_ALU_result<14>/GROM ),
    .O(N115216)
  );
  defparam DLX_EXinst__n0030_1181.INIT = 16'h0001;
  X_LUT4 DLX_EXinst__n0030_1181 (
    .ADR0(DLX_IDinst_IR_opcode_field[1]),
    .ADR1(N95411),
    .ADR2(DLX_IDinst_IR_opcode_field[0]),
    .ADR3(DLX_IDinst_IR_opcode_field[5]),
    .O(\DLX_EXinst__n0030/FROM )
  );
  defparam \DLX_EXinst__n0006<29>367_SW0 .INIT = 16'hFAFE;
  X_LUT4 \DLX_EXinst__n0006<29>367_SW0  (
    .ADR0(CHOICE5398),
    .ADR1(CHOICE5356),
    .ADR2(CHOICE5401),
    .ADR3(DLX_EXinst__n0030),
    .O(\DLX_EXinst__n0030/GROM )
  );
  X_BUF \DLX_EXinst__n0030/XUSED  (
    .I(\DLX_EXinst__n0030/FROM ),
    .O(DLX_EXinst__n0030)
  );
  X_BUF \DLX_EXinst__n0030/YUSED  (
    .I(\DLX_EXinst__n0030/GROM ),
    .O(N126437)
  );
  defparam \DLX_IDinst__n0086<29>25 .INIT = 16'hAAAE;
  X_LUT4 \DLX_IDinst__n0086<29>25  (
    .ADR0(CHOICE2903),
    .ADR1(CHOICE2899),
    .ADR2(DLX_IDinst__n0364),
    .ADR3(DLX_IDinst_N70918),
    .O(\DLX_IDinst_branch_address<29>/FROM )
  );
  defparam \DLX_IDinst__n0086<29>31 .INIT = 16'hFF88;
  X_LUT4 \DLX_IDinst__n0086<29>31  (
    .ADR0(DLX_IDinst__n0128[29]),
    .ADR1(N100609),
    .ADR2(VCC),
    .ADR3(CHOICE2904),
    .O(N107041)
  );
  X_BUF \DLX_IDinst_branch_address<29>/XUSED  (
    .I(\DLX_IDinst_branch_address<29>/FROM ),
    .O(CHOICE2904)
  );
  defparam DLX_EXinst_Ker66517.INIT = 16'h0001;
  X_LUT4 DLX_EXinst_Ker66517 (
    .ADR0(DLX_IDinst_IR_function_field[4]),
    .ADR1(N127093),
    .ADR2(DLX_IDinst_IR_function_field_3_1),
    .ADR3(DLX_EXinst__n0030_1),
    .O(\DLX_EXinst_N66519/FROM )
  );
  defparam DLX_EXinst_Ker64179_SW0.INIT = 16'h5000;
  X_LUT4 DLX_EXinst_Ker64179_SW0 (
    .ADR0(DLX_IDinst_IR_function_field_1_1),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_IR_function_field[0]),
    .ADR3(DLX_EXinst_N66519),
    .O(\DLX_EXinst_N66519/GROM )
  );
  X_BUF \DLX_EXinst_N66519/XUSED  (
    .I(\DLX_EXinst_N66519/FROM ),
    .O(DLX_EXinst_N66519)
  );
  X_BUF \DLX_EXinst_N66519/YUSED  (
    .I(\DLX_EXinst_N66519/GROM ),
    .O(N95259)
  );
  defparam DLX_EXinst_Ker64917.INIT = 16'hAFA0;
  X_LUT4 DLX_EXinst_Ker64917 (
    .ADR0(\DLX_EXinst_Mshift__n0027_Sh[8] ),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_IR_function_field_3_1),
    .ADR3(N93179),
    .O(\DLX_EXinst_N64919/FROM )
  );
  defparam \DLX_EXinst__n0006<20>16 .INIT = 16'hC808;
  X_LUT4 \DLX_EXinst__n0006<20>16  (
    .ADR0(DLX_EXinst_N64077),
    .ADR1(DLX_EXinst__n0081),
    .ADR2(DLX_IDinst_IR_function_field[2]),
    .ADR3(DLX_EXinst_N64919),
    .O(\DLX_EXinst_N64919/GROM )
  );
  X_BUF \DLX_EXinst_N64919/XUSED  (
    .I(\DLX_EXinst_N64919/FROM ),
    .O(DLX_EXinst_N64919)
  );
  X_BUF \DLX_EXinst_N64919/YUSED  (
    .I(\DLX_EXinst_N64919/GROM ),
    .O(CHOICE4878)
  );
  defparam \DLX_EXinst__n0006<22>272_SW0 .INIT = 16'hEEAA;
  X_LUT4 \DLX_EXinst__n0006<22>272_SW0  (
    .ADR0(CHOICE4154),
    .ADR1(DLX_EXinst_N66226),
    .ADR2(VCC),
    .ADR3(CHOICE4140),
    .O(\N126490/FROM )
  );
  defparam \DLX_EXinst__n0006<22>272 .INIT = 16'hCCC8;
  X_LUT4 \DLX_EXinst__n0006<22>272  (
    .ADR0(CHOICE4145),
    .ADR1(DLX_EXinst__n0030),
    .ADR2(CHOICE4130),
    .ADR3(N126490),
    .O(\N126490/GROM )
  );
  X_BUF \N126490/XUSED  (
    .I(\N126490/FROM ),
    .O(N126490)
  );
  X_BUF \N126490/YUSED  (
    .I(\N126490/GROM ),
    .O(CHOICE4157)
  );
  defparam \DLX_IFinst__n0001<11>_SW0 .INIT = 16'h5353;
  X_LUT4 \DLX_IFinst__n0001<11>_SW0  (
    .ADR0(DLX_IFinst_PC[11]),
    .ADR1(DLX_IFinst__n0015[11]),
    .ADR2(DLX_IFinst__n0000),
    .ADR3(VCC),
    .O(\DLX_IFinst_NPC<11>/FROM )
  );
  defparam \DLX_IFinst__n0001<11> .INIT = 16'h88DD;
  X_LUT4 \DLX_IFinst__n0001<11>  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(DLX_IDinst_branch_address[11]),
    .ADR2(VCC),
    .ADR3(N92503),
    .O(\DLX_IFinst_NPC<11>/GROM )
  );
  X_BUF \DLX_IFinst_NPC<11>/XUSED  (
    .I(\DLX_IFinst_NPC<11>/FROM ),
    .O(N92503)
  );
  X_BUF \DLX_IFinst_NPC<11>/YUSED  (
    .I(\DLX_IFinst_NPC<11>/GROM ),
    .O(DLX_IFinst__n0001[11])
  );
  defparam DLX_EXinst__n0128_1182.INIT = 16'h0E0A;
  X_LUT4 DLX_EXinst__n0128_1182 (
    .ADR0(N89980),
    .ADR1(DLX_EXinst_N63269),
    .ADR2(DLX_IDinst_IR_opcode_field[4]),
    .ADR3(DLX_IDinst_IR_opcode_field[5]),
    .O(\DLX_EXinst__n0128/FROM )
  );
  defparam \DLX_EXinst__n0006<25>110 .INIT = 16'hFEFC;
  X_LUT4 \DLX_EXinst__n0006<25>110  (
    .ADR0(DLX_EXinst__n0016[25]),
    .ADR1(N126301),
    .ADR2(CHOICE4751),
    .ADR3(DLX_EXinst__n0128),
    .O(\DLX_EXinst__n0128/GROM )
  );
  X_BUF \DLX_EXinst__n0128/XUSED  (
    .I(\DLX_EXinst__n0128/FROM ),
    .O(DLX_EXinst__n0128)
  );
  X_BUF \DLX_EXinst__n0128/YUSED  (
    .I(\DLX_EXinst__n0128/GROM ),
    .O(CHOICE4766)
  );
  defparam DLX_IDlc_md_mda32_a1.INIT = 16'h4444;
  X_LUT4 DLX_IDlc_md_mda32_a1 (
    .ADR0(DLX_IDlc_pd_wint1),
    .ADR1(DLX_IDlc_md_wint31),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IDlc_md_wint32/FROM )
  );
  defparam DLX_IDlc_md_mda10_a1.INIT = 16'h00AA;
  X_LUT4 DLX_IDlc_md_mda10_a1 (
    .ADR0(DLX_IDlc_md_wint9),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDlc_pd_wint1),
    .O(\DLX_IDlc_md_wint32/GROM )
  );
  X_BUF \DLX_IDlc_md_wint32/XUSED  (
    .I(\DLX_IDlc_md_wint32/FROM ),
    .O(DLX_IDlc_md_wint32)
  );
  X_BUF \DLX_IDlc_md_wint32/YUSED  (
    .I(\DLX_IDlc_md_wint32/GROM ),
    .O(DLX_IDlc_md_wint10)
  );
  defparam DLX_IDlc_md_mda29_a1.INIT = 16'h4444;
  X_LUT4 DLX_IDlc_md_mda29_a1 (
    .ADR0(DLX_IDlc_pd_wint1),
    .ADR1(DLX_IDlc_md_wint28),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IDlc_md_wint29/FROM )
  );
  defparam DLX_IDlc_md_mda11_a1.INIT = 16'h4444;
  X_LUT4 DLX_IDlc_md_mda11_a1 (
    .ADR0(DLX_IDlc_pd_wint1),
    .ADR1(DLX_IDlc_md_wint10),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IDlc_md_wint29/GROM )
  );
  X_BUF \DLX_IDlc_md_wint29/XUSED  (
    .I(\DLX_IDlc_md_wint29/FROM ),
    .O(DLX_IDlc_md_wint29)
  );
  X_BUF \DLX_IDlc_md_wint29/YUSED  (
    .I(\DLX_IDlc_md_wint29/GROM ),
    .O(DLX_IDlc_md_wint11)
  );
  defparam \DLX_EXinst__n0006<21>222 .INIT = 16'hFCCC;
  X_LUT4 \DLX_EXinst__n0006<21>222  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N64448),
    .ADR2(DLX_IDinst_reg_out_B[21]),
    .ADR3(DLX_EXinst__n0045),
    .O(\CHOICE4217/FROM )
  );
  defparam \DLX_EXinst__n0006<15>210_SW0 .INIT = 16'hFDEC;
  X_LUT4 \DLX_EXinst__n0006<15>210_SW0  (
    .ADR0(DLX_IDinst_reg_out_B[15]),
    .ADR1(DLX_EXinst_N64448),
    .ADR2(DLX_EXinst__n0045),
    .ADR3(DLX_EXinst__n0047),
    .O(\CHOICE4217/GROM )
  );
  X_BUF \CHOICE4217/XUSED  (
    .I(\CHOICE4217/FROM ),
    .O(CHOICE4217)
  );
  X_BUF \CHOICE4217/YUSED  (
    .I(\CHOICE4217/GROM ),
    .O(N126257)
  );
  defparam \DLX_IFinst__n0001<20>_SW0 .INIT = 16'h0F55;
  X_LUT4 \DLX_IFinst__n0001<20>_SW0  (
    .ADR0(DLX_IFinst__n0015[20]),
    .ADR1(VCC),
    .ADR2(DLX_IFinst_PC[20]),
    .ADR3(DLX_IFinst__n0000),
    .O(\DLX_IFinst_NPC<20>/FROM )
  );
  defparam \DLX_IFinst__n0001<20> .INIT = 16'h88DD;
  X_LUT4 \DLX_IFinst__n0001<20>  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(DLX_IDinst_branch_address[20]),
    .ADR2(VCC),
    .ADR3(N92087),
    .O(DLX_IFinst__n0001[20])
  );
  X_BUF \DLX_IFinst_NPC<20>/XUSED  (
    .I(\DLX_IFinst_NPC<20>/FROM ),
    .O(N92087)
  );
  defparam \DLX_IFinst__n0001<12>_SW0 .INIT = 16'h11DD;
  X_LUT4 \DLX_IFinst__n0001<12>_SW0  (
    .ADR0(DLX_IFinst__n0015[12]),
    .ADR1(DLX_IFinst__n0000),
    .ADR2(VCC),
    .ADR3(DLX_IFinst_PC[12]),
    .O(\DLX_IFinst_NPC<12>/FROM )
  );
  defparam \DLX_IFinst__n0001<12> .INIT = 16'hC0CF;
  X_LUT4 \DLX_IFinst__n0001<12>  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_branch_address[12]),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(N92555),
    .O(\DLX_IFinst_NPC<12>/GROM )
  );
  X_BUF \DLX_IFinst_NPC<12>/XUSED  (
    .I(\DLX_IFinst_NPC<12>/FROM ),
    .O(N92555)
  );
  X_BUF \DLX_IFinst_NPC<12>/YUSED  (
    .I(\DLX_IFinst_NPC<12>/GROM ),
    .O(DLX_IFinst__n0001[12])
  );
  defparam DLX_IDlc_md_mda28_a1.INIT = 16'h00AA;
  X_LUT4 DLX_IDlc_md_mda28_a1 (
    .ADR0(DLX_IDlc_md_wint27),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDlc_pd_wint1),
    .O(\DLX_IDlc_md_wint28/FROM )
  );
  defparam DLX_IDlc_md_mda20_a1.INIT = 16'h00AA;
  X_LUT4 DLX_IDlc_md_mda20_a1 (
    .ADR0(DLX_IDlc_md_wint19),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDlc_pd_wint1),
    .O(\DLX_IDlc_md_wint28/GROM )
  );
  X_BUF \DLX_IDlc_md_wint28/XUSED  (
    .I(\DLX_IDlc_md_wint28/FROM ),
    .O(DLX_IDlc_md_wint28)
  );
  X_BUF \DLX_IDlc_md_wint28/YUSED  (
    .I(\DLX_IDlc_md_wint28/GROM ),
    .O(DLX_IDlc_md_wint20)
  );
  defparam DLX_IDlc_md_mda25_a1.INIT = 16'h00AA;
  X_LUT4 DLX_IDlc_md_mda25_a1 (
    .ADR0(DLX_IDlc_md_wint24),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDlc_pd_wint1),
    .O(\DLX_IDlc_md_wint25/FROM )
  );
  defparam DLX_IDlc_md_mda12_a1.INIT = 16'h00CC;
  X_LUT4 DLX_IDlc_md_mda12_a1 (
    .ADR0(VCC),
    .ADR1(DLX_IDlc_md_wint11),
    .ADR2(VCC),
    .ADR3(DLX_IDlc_pd_wint1),
    .O(\DLX_IDlc_md_wint25/GROM )
  );
  X_BUF \DLX_IDlc_md_wint25/XUSED  (
    .I(\DLX_IDlc_md_wint25/FROM ),
    .O(DLX_IDlc_md_wint25)
  );
  X_BUF \DLX_IDlc_md_wint25/YUSED  (
    .I(\DLX_IDlc_md_wint25/GROM ),
    .O(DLX_IDlc_md_wint12)
  );
  defparam clk_DM1.INIT = 16'hFA00;
  X_LUT4 clk_DM1 (
    .ADR0(DLX_EXinst_mem_read_EX),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_mem_write_EX),
    .ADR3(clk_EX_del),
    .O(\clk_DM_OBUF/GROM )
  );
  X_BUF \clk_DM_OBUF/YUSED  (
    .I(\clk_DM_OBUF/GROM ),
    .O(clk_DM_OBUF)
  );
  defparam \DLX_IFinst__n0001<0>_SW0 .INIT = 16'h4477;
  X_LUT4 \DLX_IFinst__n0001<0>_SW0  (
    .ADR0(DLX_IFinst_PC[0]),
    .ADR1(DLX_IFinst__n0000),
    .ADR2(VCC),
    .ADR3(DLX_IFinst_NPC[0]),
    .O(\DLX_IFinst_NPC<0>/FROM )
  );
  defparam \DLX_IFinst__n0001<0> .INIT = 16'hC0F3;
  X_LUT4 \DLX_IFinst__n0001<0>  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(DLX_IDinst_branch_address[0]),
    .ADR3(N91463),
    .O(\DLX_IFinst_NPC<0>/GROM )
  );
  X_BUF \DLX_IFinst_NPC<0>/XUSED  (
    .I(\DLX_IFinst_NPC<0>/FROM ),
    .O(N91463)
  );
  X_BUF \DLX_IFinst_NPC<0>/YUSED  (
    .I(\DLX_IFinst_NPC<0>/GROM ),
    .O(DLX_IFinst__n0001[0])
  );
  defparam DLX_IDlc_md_mda24_a1.INIT = 16'h5050;
  X_LUT4 DLX_IDlc_md_mda24_a1 (
    .ADR0(DLX_IDlc_pd_wint1),
    .ADR1(VCC),
    .ADR2(DLX_IDlc_md_wint23),
    .ADR3(VCC),
    .O(\DLX_IDlc_md_wint24/FROM )
  );
  defparam DLX_IDlc_md_mda21_a1.INIT = 16'h4444;
  X_LUT4 DLX_IDlc_md_mda21_a1 (
    .ADR0(DLX_IDlc_pd_wint1),
    .ADR1(DLX_IDlc_md_wint20),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IDlc_md_wint24/GROM )
  );
  X_BUF \DLX_IDlc_md_wint24/XUSED  (
    .I(\DLX_IDlc_md_wint24/FROM ),
    .O(DLX_IDlc_md_wint24)
  );
  X_BUF \DLX_IDlc_md_wint24/YUSED  (
    .I(\DLX_IDlc_md_wint24/GROM ),
    .O(DLX_IDlc_md_wint21)
  );
  defparam DLX_IDlc_md_mda23_a1.INIT = 16'h4444;
  X_LUT4 DLX_IDlc_md_mda23_a1 (
    .ADR0(DLX_IDlc_pd_wint1),
    .ADR1(DLX_IDlc_md_wint22),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IDlc_md_wint23/FROM )
  );
  defparam DLX_IDlc_md_mda13_a1.INIT = 16'h0C0C;
  X_LUT4 DLX_IDlc_md_mda13_a1 (
    .ADR0(VCC),
    .ADR1(DLX_IDlc_md_wint12),
    .ADR2(DLX_IDlc_pd_wint1),
    .ADR3(VCC),
    .O(\DLX_IDlc_md_wint23/GROM )
  );
  X_BUF \DLX_IDlc_md_wint23/XUSED  (
    .I(\DLX_IDlc_md_wint23/FROM ),
    .O(DLX_IDlc_md_wint23)
  );
  X_BUF \DLX_IDlc_md_wint23/YUSED  (
    .I(\DLX_IDlc_md_wint23/GROM ),
    .O(DLX_IDlc_md_wint13)
  );
  defparam \DLX_EXinst__n0006<0>568_SW0 .INIT = 16'hEE22;
  X_LUT4 \DLX_EXinst__n0006<0>568_SW0  (
    .ADR0(DLX_IDinst_reg_out_A[0]),
    .ADR1(DLX_IDinst_IR_function_field[1]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[2]),
    .O(\N126048/FROM )
  );
  defparam \DLX_EXinst__n0006<0>568 .INIT = 16'h2320;
  X_LUT4 \DLX_EXinst__n0006<0>568  (
    .ADR0(DLX_EXinst_N65135),
    .ADR1(DLX_IDinst_IR_function_field[3]),
    .ADR2(DLX_IDinst_IR_function_field[0]),
    .ADR3(N126048),
    .O(\N126048/GROM )
  );
  X_BUF \N126048/XUSED  (
    .I(\N126048/FROM ),
    .O(N126048)
  );
  X_BUF \N126048/YUSED  (
    .I(\N126048/GROM ),
    .O(CHOICE5969)
  );
  defparam \DLX_IDinst__n0086<8>6 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst__n0086<8>6  (
    .ADR0(DLX_IDinst_N70786),
    .ADR1(DLX_IDinst_branch_address[8]),
    .ADR2(DLX_IDinst_EPC[8]),
    .ADR3(DLX_IDinst__n0071),
    .O(\CHOICE2646/GROM )
  );
  X_BUF \CHOICE2646/YUSED  (
    .I(\CHOICE2646/GROM ),
    .O(CHOICE2646)
  );
  defparam \DLX_IDinst_regA_eff<10>1 .INIT = 16'hC5C0;
  X_LUT4 \DLX_IDinst_regA_eff<10>1  (
    .ADR0(DLX_IDinst__n0002),
    .ADR1(DLX_MEMinst_RF_data_in[10]),
    .ADR2(DLX_IDinst__n0144),
    .ADR3(DLX_IDinst_reg_out_A_RF[10]),
    .O(\DLX_IDinst_regA_eff<10>/FROM )
  );
  defparam \DLX_IDinst__n0086<10>20 .INIT = 16'hAA00;
  X_LUT4 \DLX_IDinst__n0086<10>20  (
    .ADR0(DLX_IDinst_N70295),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_regA_eff[10]),
    .O(\DLX_IDinst_regA_eff<10>/GROM )
  );
  X_BUF \DLX_IDinst_regA_eff<10>/XUSED  (
    .I(\DLX_IDinst_regA_eff<10>/FROM ),
    .O(DLX_IDinst_regA_eff[10])
  );
  X_BUF \DLX_IDinst_regA_eff<10>/YUSED  (
    .I(\DLX_IDinst_regA_eff<10>/GROM ),
    .O(CHOICE2672)
  );
  defparam DLX_IDlc_md_mda30_a1.INIT = 16'h00CC;
  X_LUT4 DLX_IDlc_md_mda30_a1 (
    .ADR0(VCC),
    .ADR1(DLX_IDlc_md_wint29),
    .ADR2(VCC),
    .ADR3(DLX_IDlc_pd_wint1),
    .O(\DLX_IDlc_md_wint30/FROM )
  );
  defparam DLX_IDlc_md_mda31_a1.INIT = 16'h5500;
  X_LUT4 DLX_IDlc_md_mda31_a1 (
    .ADR0(DLX_IDlc_pd_wint1),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDlc_md_wint30),
    .O(\DLX_IDlc_md_wint30/GROM )
  );
  X_BUF \DLX_IDlc_md_wint30/XUSED  (
    .I(\DLX_IDlc_md_wint30/FROM ),
    .O(DLX_IDlc_md_wint30)
  );
  X_BUF \DLX_IDlc_md_wint30/YUSED  (
    .I(\DLX_IDlc_md_wint30/GROM ),
    .O(DLX_IDlc_md_wint31)
  );
  defparam DLX_IDlc_md_mda19_a1.INIT = 16'h2222;
  X_LUT4 DLX_IDlc_md_mda19_a1 (
    .ADR0(DLX_IDlc_md_wint18),
    .ADR1(DLX_IDlc_pd_wint1),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IDlc_md_wint19/FROM )
  );
  defparam DLX_IDlc_md_mda22_a1.INIT = 16'h2222;
  X_LUT4 DLX_IDlc_md_mda22_a1 (
    .ADR0(DLX_IDlc_md_wint21),
    .ADR1(DLX_IDlc_pd_wint1),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IDlc_md_wint19/GROM )
  );
  X_BUF \DLX_IDlc_md_wint19/XUSED  (
    .I(\DLX_IDlc_md_wint19/FROM ),
    .O(DLX_IDlc_md_wint19)
  );
  X_BUF \DLX_IDlc_md_wint19/YUSED  (
    .I(\DLX_IDlc_md_wint19/GROM ),
    .O(DLX_IDlc_md_wint22)
  );
  defparam DLX_IDlc_md_mda18_a1.INIT = 16'h5050;
  X_LUT4 DLX_IDlc_md_mda18_a1 (
    .ADR0(DLX_IDlc_pd_wint1),
    .ADR1(VCC),
    .ADR2(DLX_IDlc_md_wint17),
    .ADR3(VCC),
    .O(\DLX_IDlc_md_wint18/FROM )
  );
  defparam DLX_IDlc_md_mda14_a1.INIT = 16'h0F00;
  X_LUT4 DLX_IDlc_md_mda14_a1 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IDlc_pd_wint1),
    .ADR3(DLX_IDlc_md_wint13),
    .O(\DLX_IDlc_md_wint18/GROM )
  );
  X_BUF \DLX_IDlc_md_wint18/XUSED  (
    .I(\DLX_IDlc_md_wint18/FROM ),
    .O(DLX_IDlc_md_wint18)
  );
  X_BUF \DLX_IDlc_md_wint18/YUSED  (
    .I(\DLX_IDlc_md_wint18/GROM ),
    .O(DLX_IDlc_md_wint14)
  );
  defparam DLX_IFlc_master_ctrlIF__n0001_SW19.INIT = 16'hFCFF;
  X_LUT4 DLX_IFlc_master_ctrlIF__n0001_SW19 (
    .ADR0(VCC),
    .ADR1(reset_IBUF_1),
    .ADR2(DLX_IFlc_master_ctrlIF_l),
    .ADR3(DLX_IFlc_master_ctrlIF_nro),
    .O(\CHOICE32/FROM )
  );
  defparam DLX_IFlc_master_ctrlIF__n0001_SW111.INIT = 16'h5500;
  X_LUT4 DLX_IFlc_master_ctrlIF__n0001_SW111 (
    .ADR0(DLX_IFlc_md_outp2),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(CHOICE32),
    .O(\CHOICE32/GROM )
  );
  X_BUF \CHOICE32/XUSED  (
    .I(\CHOICE32/FROM ),
    .O(CHOICE32)
  );
  X_BUF \CHOICE32/YUSED  (
    .I(\CHOICE32/GROM ),
    .O(DLX_IFlc_master_ctrlIF_l)
  );
  defparam DLX_IDinst_Ker7064013.INIT = 16'h00FA;
  X_LUT4 DLX_IDinst_Ker7064013 (
    .ADR0(DLX_IDinst__n0075),
    .ADR1(VCC),
    .ADR2(DLX_IDinst__n0078),
    .ADR3(DLX_IDinst__n0004),
    .O(\CHOICE3328/FROM )
  );
  defparam DLX_IDinst_Ker7064017.INIT = 16'hFF32;
  X_LUT4 DLX_IDinst_Ker7064017 (
    .ADR0(DLX_IDinst__n0073),
    .ADR1(DLX_IDinst__n0002),
    .ADR2(DLX_IDinst__n0077),
    .ADR3(CHOICE3328),
    .O(\CHOICE3328/GROM )
  );
  X_BUF \CHOICE3328/XUSED  (
    .I(\CHOICE3328/FROM ),
    .O(CHOICE3328)
  );
  X_BUF \CHOICE3328/YUSED  (
    .I(\CHOICE3328/GROM ),
    .O(CHOICE3329)
  );
  defparam \DLX_IDinst_regA_eff<11>1 .INIT = 16'hB1A0;
  X_LUT4 \DLX_IDinst_regA_eff<11>1  (
    .ADR0(DLX_IDinst__n0144),
    .ADR1(DLX_IDinst__n0002),
    .ADR2(DLX_MEMinst_RF_data_in[11]),
    .ADR3(DLX_IDinst_reg_out_A_RF[11]),
    .O(\DLX_IDinst_regA_eff<11>/FROM )
  );
  defparam DLX_IDinst__n014649.INIT = 16'h0001;
  X_LUT4 DLX_IDinst__n014649 (
    .ADR0(DLX_IDinst_regA_eff[10]),
    .ADR1(DLX_IDinst_regA_eff[9]),
    .ADR2(DLX_IDinst_regA_eff[8]),
    .ADR3(DLX_IDinst_regA_eff[11]),
    .O(\DLX_IDinst_regA_eff<11>/GROM )
  );
  X_BUF \DLX_IDinst_regA_eff<11>/XUSED  (
    .I(\DLX_IDinst_regA_eff<11>/FROM ),
    .O(DLX_IDinst_regA_eff[11])
  );
  X_BUF \DLX_IDinst_regA_eff<11>/YUSED  (
    .I(\DLX_IDinst_regA_eff<11>/GROM ),
    .O(CHOICE3635)
  );
  defparam DLX_EXinst_Ker63994_SW0.INIT = 16'hF3FF;
  X_LUT4 DLX_EXinst_Ker63994_SW0 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_IR_function_field_1_1),
    .ADR2(DLX_IDinst_IR_function_field[0]),
    .ADR3(DLX_EXinst_N66519),
    .O(\N95327/FROM )
  );
  defparam DLX_EXinst_Ker63994.INIT = 16'h08FF;
  X_LUT4 DLX_EXinst_Ker63994 (
    .ADR0(DLX_EXinst_N66072),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(DLX_IDinst_reg_out_B[0]),
    .ADR3(N95327),
    .O(\N95327/GROM )
  );
  X_BUF \N95327/XUSED  (
    .I(\N95327/FROM ),
    .O(N95327)
  );
  X_BUF \N95327/YUSED  (
    .I(\N95327/GROM ),
    .O(DLX_EXinst_N63996)
  );
  defparam \DLX_IDinst_regA_eff<12>1 .INIT = 16'h88D8;
  X_LUT4 \DLX_IDinst_regA_eff<12>1  (
    .ADR0(DLX_IDinst__n0144),
    .ADR1(DLX_MEMinst_RF_data_in[12]),
    .ADR2(DLX_IDinst_reg_out_A_RF[12]),
    .ADR3(DLX_IDinst__n0002),
    .O(\DLX_IDinst_regA_eff<12>/FROM )
  );
  defparam \DLX_IDinst__n0086<12>20 .INIT = 16'hF000;
  X_LUT4 \DLX_IDinst__n0086<12>20  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_N70295),
    .ADR3(DLX_IDinst_regA_eff[12]),
    .O(\DLX_IDinst_regA_eff<12>/GROM )
  );
  X_BUF \DLX_IDinst_regA_eff<12>/XUSED  (
    .I(\DLX_IDinst_regA_eff<12>/FROM ),
    .O(DLX_IDinst_regA_eff[12])
  );
  X_BUF \DLX_IDinst_regA_eff<12>/YUSED  (
    .I(\DLX_IDinst_regA_eff<12>/GROM ),
    .O(CHOICE2694)
  );
  defparam \DLX_IDinst_regA_eff<20>1 .INIT = 16'hA3A0;
  X_LUT4 \DLX_IDinst_regA_eff<20>1  (
    .ADR0(DLX_MEMinst_RF_data_in[20]),
    .ADR1(DLX_IDinst__n0002),
    .ADR2(DLX_IDinst__n0144),
    .ADR3(DLX_IDinst_reg_out_A_RF[20]),
    .O(\DLX_IDinst_regA_eff<20>/FROM )
  );
  defparam \DLX_IDinst__n0086<20>20 .INIT = 16'hF000;
  X_LUT4 \DLX_IDinst__n0086<20>20  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_N70295),
    .ADR3(DLX_IDinst_regA_eff[20]),
    .O(\DLX_IDinst_regA_eff<20>/GROM )
  );
  X_BUF \DLX_IDinst_regA_eff<20>/XUSED  (
    .I(\DLX_IDinst_regA_eff<20>/FROM ),
    .O(DLX_IDinst_regA_eff[20])
  );
  X_BUF \DLX_IDinst_regA_eff<20>/YUSED  (
    .I(\DLX_IDinst_regA_eff<20>/GROM ),
    .O(CHOICE2782)
  );
  defparam DLX_IDlc_md_mda17_a1.INIT = 16'h00CC;
  X_LUT4 DLX_IDlc_md_mda17_a1 (
    .ADR0(VCC),
    .ADR1(DLX_IDlc_md_wint16),
    .ADR2(VCC),
    .ADR3(DLX_IDlc_pd_wint1),
    .O(\DLX_IDlc_md_wint17/FROM )
  );
  defparam DLX_IDlc_md_mda15_a1.INIT = 16'h3300;
  X_LUT4 DLX_IDlc_md_mda15_a1 (
    .ADR0(VCC),
    .ADR1(DLX_IDlc_pd_wint1),
    .ADR2(VCC),
    .ADR3(DLX_IDlc_md_wint14),
    .O(\DLX_IDlc_md_wint17/GROM )
  );
  X_BUF \DLX_IDlc_md_wint17/XUSED  (
    .I(\DLX_IDlc_md_wint17/FROM ),
    .O(DLX_IDlc_md_wint17)
  );
  X_BUF \DLX_IDlc_md_wint17/YUSED  (
    .I(\DLX_IDlc_md_wint17/GROM ),
    .O(DLX_IDlc_md_wint15)
  );
  defparam \DLX_EXinst_Mshift__n0027_Sh<10>1 .INIT = 16'hAFA0;
  X_LUT4 \DLX_EXinst_Mshift__n0027_Sh<10>1  (
    .ADR0(DLX_EXinst_N62771),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_IR_function_field_0_1),
    .ADR3(DLX_EXinst_N63439),
    .O(\DLX_EXinst_Mshift__n0027_Sh<10>/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0027_Sh<46>_SW0 .INIT = 16'hFA50;
  X_LUT4 \DLX_EXinst_Mshift__n0027_Sh<46>_SW0  (
    .ADR0(DLX_IDinst_IR_function_field_2_1),
    .ADR1(VCC),
    .ADR2(\DLX_EXinst_Mshift__n0027_Sh[14] ),
    .ADR3(\DLX_EXinst_Mshift__n0027_Sh[10] ),
    .O(\DLX_EXinst_Mshift__n0027_Sh<10>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0027_Sh<10>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0027_Sh<10>/FROM ),
    .O(\DLX_EXinst_Mshift__n0027_Sh[10] )
  );
  X_BUF \DLX_EXinst_Mshift__n0027_Sh<10>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0027_Sh<10>/GROM ),
    .O(N93331)
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<30>1 .INIT = 16'hFE10;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<30>1  (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(DLX_IDinst_reg_out_A[30]),
    .ADR3(DLX_IDinst_reg_out_A[31]),
    .O(\DLX_EXinst_Mshift__n0023_Sh<30>/FROM )
  );
  defparam DLX_EXinst_Ker6509333.INIT = 16'hCDCC;
  X_LUT4 DLX_EXinst_Ker6509333 (
    .ADR0(DLX_IDinst_reg_out_B[5]),
    .ADR1(CHOICE859),
    .ADR2(DLX_EXinst_N62740),
    .ADR3(\DLX_EXinst_Mshift__n0023_Sh[30] ),
    .O(\DLX_EXinst_Mshift__n0023_Sh<30>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0023_Sh<30>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0023_Sh<30>/FROM ),
    .O(\DLX_EXinst_Mshift__n0023_Sh[30] )
  );
  X_BUF \DLX_EXinst_Mshift__n0023_Sh<30>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0023_Sh<30>/GROM ),
    .O(N95120)
  );
  X_INV \DLX_MEMinst_noop/CKINV  (
    .I(DLX_MEMlc_master_ctrlMEM_l),
    .O(\DLX_MEMinst_noop/CKMUXNOT )
  );
  defparam \DLX_IDinst_regA_eff<13>1 .INIT = 16'hA0E4;
  X_LUT4 \DLX_IDinst_regA_eff<13>1  (
    .ADR0(DLX_IDinst__n0144),
    .ADR1(DLX_IDinst_reg_out_A_RF[13]),
    .ADR2(DLX_MEMinst_RF_data_in[13]),
    .ADR3(DLX_IDinst__n0002),
    .O(\DLX_IDinst_regA_eff<13>/FROM )
  );
  defparam \DLX_IDinst__n0086<13>20 .INIT = 16'hCC00;
  X_LUT4 \DLX_IDinst__n0086<13>20  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_N70295),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_regA_eff[13]),
    .O(\DLX_IDinst_regA_eff<13>/GROM )
  );
  X_BUF \DLX_IDinst_regA_eff<13>/XUSED  (
    .I(\DLX_IDinst_regA_eff<13>/FROM ),
    .O(DLX_IDinst_regA_eff[13])
  );
  X_BUF \DLX_IDinst_regA_eff<13>/YUSED  (
    .I(\DLX_IDinst_regA_eff<13>/GROM ),
    .O(CHOICE2705)
  );
  defparam \DLX_IDinst_regA_eff<21>1 .INIT = 16'hCE02;
  X_LUT4 \DLX_IDinst_regA_eff<21>1  (
    .ADR0(DLX_IDinst_reg_out_A_RF[21]),
    .ADR1(DLX_IDinst__n0144),
    .ADR2(DLX_IDinst__n0002),
    .ADR3(DLX_MEMinst_RF_data_in[21]),
    .O(\DLX_IDinst_regA_eff<21>/FROM )
  );
  defparam \DLX_IDinst__n0086<21>20 .INIT = 16'hAA00;
  X_LUT4 \DLX_IDinst__n0086<21>20  (
    .ADR0(DLX_IDinst_N70295),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_regA_eff[21]),
    .O(\DLX_IDinst_regA_eff<21>/GROM )
  );
  X_BUF \DLX_IDinst_regA_eff<21>/XUSED  (
    .I(\DLX_IDinst_regA_eff<21>/FROM ),
    .O(DLX_IDinst_regA_eff[21])
  );
  X_BUF \DLX_IDinst_regA_eff<21>/YUSED  (
    .I(\DLX_IDinst_regA_eff<21>/GROM ),
    .O(CHOICE2804)
  );
  defparam \DLX_IFinst__n0001<13>_SW0 .INIT = 16'h2727;
  X_LUT4 \DLX_IFinst__n0001<13>_SW0  (
    .ADR0(DLX_IFinst__n0000),
    .ADR1(DLX_IFinst_PC[13]),
    .ADR2(DLX_IFinst__n0015[13]),
    .ADR3(VCC),
    .O(\DLX_IFinst_NPC<13>/FROM )
  );
  defparam \DLX_IFinst__n0001<13> .INIT = 16'hA0AF;
  X_LUT4 \DLX_IFinst__n0001<13>  (
    .ADR0(DLX_IDinst_branch_address[13]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(N92451),
    .O(\DLX_IFinst_NPC<13>/GROM )
  );
  X_BUF \DLX_IFinst_NPC<13>/XUSED  (
    .I(\DLX_IFinst_NPC<13>/FROM ),
    .O(N92451)
  );
  X_BUF \DLX_IFinst_NPC<13>/YUSED  (
    .I(\DLX_IFinst_NPC<13>/GROM ),
    .O(DLX_IFinst__n0001[13])
  );
  defparam \DLX_IFinst__n0001<21>_SW0 .INIT = 16'h4747;
  X_LUT4 \DLX_IFinst__n0001<21>_SW0  (
    .ADR0(DLX_IFinst_PC[21]),
    .ADR1(DLX_IFinst__n0000),
    .ADR2(DLX_IFinst__n0015[21]),
    .ADR3(VCC),
    .O(\DLX_IFinst_NPC<21>/FROM )
  );
  defparam \DLX_IFinst__n0001<21> .INIT = 16'hC0CF;
  X_LUT4 \DLX_IFinst__n0001<21>  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_branch_address[21]),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(N91983),
    .O(DLX_IFinst__n0001[21])
  );
  X_BUF \DLX_IFinst_NPC<21>/XUSED  (
    .I(\DLX_IFinst_NPC<21>/FROM ),
    .O(N91983)
  );
  defparam \DLX_IDinst_regA_eff<14>1 .INIT = 16'h8D88;
  X_LUT4 \DLX_IDinst_regA_eff<14>1  (
    .ADR0(DLX_IDinst__n0144),
    .ADR1(DLX_MEMinst_RF_data_in[14]),
    .ADR2(DLX_IDinst__n0002),
    .ADR3(DLX_IDinst_reg_out_A_RF[14]),
    .O(\DLX_IDinst_regA_eff<14>/FROM )
  );
  defparam \DLX_IDinst__n0086<14>20 .INIT = 16'hAA00;
  X_LUT4 \DLX_IDinst__n0086<14>20  (
    .ADR0(DLX_IDinst_N70295),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_regA_eff[14]),
    .O(\DLX_IDinst_regA_eff<14>/GROM )
  );
  X_BUF \DLX_IDinst_regA_eff<14>/XUSED  (
    .I(\DLX_IDinst_regA_eff<14>/FROM ),
    .O(DLX_IDinst_regA_eff[14])
  );
  X_BUF \DLX_IDinst_regA_eff<14>/YUSED  (
    .I(\DLX_IDinst_regA_eff<14>/GROM ),
    .O(CHOICE2716)
  );
  defparam \DLX_IDinst_regA_eff<22>1 .INIT = 16'hA0E4;
  X_LUT4 \DLX_IDinst_regA_eff<22>1  (
    .ADR0(DLX_IDinst__n0144),
    .ADR1(DLX_IDinst_reg_out_A_RF[22]),
    .ADR2(DLX_MEMinst_RF_data_in[22]),
    .ADR3(DLX_IDinst__n0002),
    .O(\DLX_IDinst_regA_eff<22>/FROM )
  );
  defparam \DLX_IDinst__n0086<22>20 .INIT = 16'hF000;
  X_LUT4 \DLX_IDinst__n0086<22>20  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_N70295),
    .ADR3(DLX_IDinst_regA_eff[22]),
    .O(\DLX_IDinst_regA_eff<22>/GROM )
  );
  X_BUF \DLX_IDinst_regA_eff<22>/XUSED  (
    .I(\DLX_IDinst_regA_eff<22>/FROM ),
    .O(DLX_IDinst_regA_eff[22])
  );
  X_BUF \DLX_IDinst_regA_eff<22>/YUSED  (
    .I(\DLX_IDinst_regA_eff<22>/GROM ),
    .O(CHOICE2826)
  );
  defparam DLX_IDinst_Ker7064058.INIT = 16'h3EFE;
  X_LUT4 DLX_IDinst_Ker7064058 (
    .ADR0(N127555),
    .ADR1(DLX_IDinst_IR_latched[27]),
    .ADR2(DLX_IDinst_IR_latched[30]),
    .ADR3(DLX_IDinst_N70991),
    .O(\CHOICE3343/FROM )
  );
  defparam DLX_IDinst_Ker70640122_SW0.INIT = 16'hAFBF;
  X_LUT4 DLX_IDinst_Ker70640122_SW0 (
    .ADR0(DLX_IDinst__n0070),
    .ADR1(CHOICE3329),
    .ADR2(CHOICE3353),
    .ADR3(CHOICE3343),
    .O(\CHOICE3343/GROM )
  );
  X_BUF \CHOICE3343/XUSED  (
    .I(\CHOICE3343/FROM ),
    .O(CHOICE3343)
  );
  X_BUF \CHOICE3343/YUSED  (
    .I(\CHOICE3343/GROM ),
    .O(N126506)
  );
  defparam DLX_IDlc_md_mda9_a1.INIT = 16'h4444;
  X_LUT4 DLX_IDlc_md_mda9_a1 (
    .ADR0(DLX_IDlc_pd_wint1),
    .ADR1(DLX_IDlc_md_wint8),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IDlc_md_wint9/FROM )
  );
  defparam DLX_IDlc_md_mda16_a1.INIT = 16'h00CC;
  X_LUT4 DLX_IDlc_md_mda16_a1 (
    .ADR0(VCC),
    .ADR1(DLX_IDlc_md_wint15),
    .ADR2(VCC),
    .ADR3(DLX_IDlc_pd_wint1),
    .O(\DLX_IDlc_md_wint9/GROM )
  );
  X_BUF \DLX_IDlc_md_wint9/XUSED  (
    .I(\DLX_IDlc_md_wint9/FROM ),
    .O(DLX_IDlc_md_wint9)
  );
  X_BUF \DLX_IDlc_md_wint9/YUSED  (
    .I(\DLX_IDlc_md_wint9/GROM ),
    .O(DLX_IDlc_md_wint16)
  );
  defparam \DLX_EXinst_Mshift__n0027_Sh<12>1 .INIT = 16'hFC30;
  X_LUT4 \DLX_EXinst_Mshift__n0027_Sh<12>1  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_IR_function_field_0_1),
    .ADR2(DLX_EXinst_N63444),
    .ADR3(DLX_EXinst_N62776),
    .O(\DLX_EXinst_Mshift__n0027_Sh<12>/FROM )
  );
  defparam DLX_EXinst_Ker640751.INIT = 16'hFA0A;
  X_LUT4 DLX_EXinst_Ker640751 (
    .ADR0(\DLX_EXinst_Mshift__n0027_Sh[20] ),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_IR_function_field[3]),
    .ADR3(\DLX_EXinst_Mshift__n0027_Sh[12] ),
    .O(\DLX_EXinst_Mshift__n0027_Sh<12>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0027_Sh<12>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0027_Sh<12>/FROM ),
    .O(\DLX_EXinst_Mshift__n0027_Sh[12] )
  );
  X_BUF \DLX_EXinst_Mshift__n0027_Sh<12>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0027_Sh<12>/GROM ),
    .O(DLX_EXinst_N64077)
  );
  defparam \DLX_IDinst_regA_eff<15>1 .INIT = 16'hCC50;
  X_LUT4 \DLX_IDinst_regA_eff<15>1  (
    .ADR0(DLX_IDinst__n0002),
    .ADR1(DLX_MEMinst_RF_data_in[15]),
    .ADR2(DLX_IDinst_reg_out_A_RF[15]),
    .ADR3(DLX_IDinst__n0144),
    .O(\DLX_IDinst_regA_eff<15>/FROM )
  );
  defparam DLX_IDinst__n014662.INIT = 16'h0001;
  X_LUT4 DLX_IDinst__n014662 (
    .ADR0(DLX_IDinst_regA_eff[14]),
    .ADR1(DLX_IDinst_regA_eff[12]),
    .ADR2(DLX_IDinst_regA_eff[13]),
    .ADR3(DLX_IDinst_regA_eff[15]),
    .O(\DLX_IDinst_regA_eff<15>/GROM )
  );
  X_BUF \DLX_IDinst_regA_eff<15>/XUSED  (
    .I(\DLX_IDinst_regA_eff<15>/FROM ),
    .O(DLX_IDinst_regA_eff[15])
  );
  X_BUF \DLX_IDinst_regA_eff<15>/YUSED  (
    .I(\DLX_IDinst_regA_eff<15>/GROM ),
    .O(CHOICE3642)
  );
  defparam \DLX_IDinst_regA_eff<23>1 .INIT = 16'hF044;
  X_LUT4 \DLX_IDinst_regA_eff<23>1  (
    .ADR0(DLX_IDinst__n0002),
    .ADR1(DLX_IDinst_reg_out_A_RF[23]),
    .ADR2(DLX_MEMinst_RF_data_in[23]),
    .ADR3(DLX_IDinst__n0144),
    .O(\DLX_IDinst_regA_eff<23>/FROM )
  );
  defparam DLX_IDinst__n0146115.INIT = 16'h0001;
  X_LUT4 DLX_IDinst__n0146115 (
    .ADR0(DLX_IDinst_regA_eff[21]),
    .ADR1(DLX_IDinst_regA_eff[20]),
    .ADR2(DLX_IDinst_regA_eff[22]),
    .ADR3(DLX_IDinst_regA_eff[23]),
    .O(\DLX_IDinst_regA_eff<23>/GROM )
  );
  X_BUF \DLX_IDinst_regA_eff<23>/XUSED  (
    .I(\DLX_IDinst_regA_eff<23>/FROM ),
    .O(DLX_IDinst_regA_eff[23])
  );
  X_BUF \DLX_IDinst_regA_eff<23>/YUSED  (
    .I(\DLX_IDinst_regA_eff<23>/GROM ),
    .O(CHOICE3658)
  );
  defparam \DLX_IDinst_regA_eff<31>1 .INIT = 16'hDC10;
  X_LUT4 \DLX_IDinst_regA_eff<31>1  (
    .ADR0(DLX_IDinst__n0002),
    .ADR1(DLX_IDinst__n0144),
    .ADR2(DLX_IDinst_reg_out_A_RF[31]),
    .ADR3(DLX_MEMinst_RF_data_in[31]),
    .O(\DLX_IDinst_regA_eff<31>/FROM )
  );
  defparam DLX_IDinst__n0146152.INIT = 16'h0001;
  X_LUT4 DLX_IDinst__n0146152 (
    .ADR0(DLX_IDinst_regA_eff[29]),
    .ADR1(DLX_IDinst_regA_eff[28]),
    .ADR2(DLX_IDinst_regA_eff[30]),
    .ADR3(DLX_IDinst_regA_eff[31]),
    .O(\DLX_IDinst_regA_eff<31>/GROM )
  );
  X_BUF \DLX_IDinst_regA_eff<31>/XUSED  (
    .I(\DLX_IDinst_regA_eff<31>/FROM ),
    .O(DLX_IDinst_regA_eff[31])
  );
  X_BUF \DLX_IDinst_regA_eff<31>/YUSED  (
    .I(\DLX_IDinst_regA_eff<31>/GROM ),
    .O(CHOICE3673)
  );
  defparam \DLX_EXinst_Mshift__n0027_Sh<13>1 .INIT = 16'hEE22;
  X_LUT4 \DLX_EXinst_Mshift__n0027_Sh<13>1  (
    .ADR0(DLX_EXinst_N62781),
    .ADR1(DLX_IDinst_IR_function_field_0_1),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N63444),
    .O(\DLX_EXinst_Mshift__n0027_Sh<13>/FROM )
  );
  defparam DLX_EXinst_Ker643021.INIT = 16'hEE44;
  X_LUT4 DLX_EXinst_Ker643021 (
    .ADR0(DLX_IDinst_IR_function_field[3]),
    .ADR1(\DLX_EXinst_Mshift__n0027_Sh[21] ),
    .ADR2(VCC),
    .ADR3(\DLX_EXinst_Mshift__n0027_Sh[13] ),
    .O(\DLX_EXinst_Mshift__n0027_Sh<13>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0027_Sh<13>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0027_Sh<13>/FROM ),
    .O(\DLX_EXinst_Mshift__n0027_Sh[13] )
  );
  X_BUF \DLX_EXinst_Mshift__n0027_Sh<13>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0027_Sh<13>/GROM ),
    .O(DLX_EXinst_N64304)
  );
  defparam \DLX_IFinst__n0001<1>_SW0 .INIT = 16'h5353;
  X_LUT4 \DLX_IFinst__n0001<1>_SW0  (
    .ADR0(DLX_IFinst_PC[1]),
    .ADR1(DLX_IFinst_NPC[1]),
    .ADR2(DLX_IFinst__n0000),
    .ADR3(VCC),
    .O(\DLX_IFinst_NPC<1>/FROM )
  );
  defparam \DLX_IFinst__n0001<1> .INIT = 16'hC0F3;
  X_LUT4 \DLX_IFinst__n0001<1>  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(DLX_IDinst_branch_address[1]),
    .ADR3(N93075),
    .O(\DLX_IFinst_NPC<1>/GROM )
  );
  X_BUF \DLX_IFinst_NPC<1>/XUSED  (
    .I(\DLX_IFinst_NPC<1>/FROM ),
    .O(N93075)
  );
  X_BUF \DLX_IFinst_NPC<1>/YUSED  (
    .I(\DLX_IFinst_NPC<1>/GROM ),
    .O(DLX_IFinst__n0001[1])
  );
  defparam \DLX_IDinst_regA_eff<16>1 .INIT = 16'hAE04;
  X_LUT4 \DLX_IDinst_regA_eff<16>1  (
    .ADR0(DLX_IDinst__n0144),
    .ADR1(DLX_IDinst_reg_out_A_RF[16]),
    .ADR2(DLX_IDinst__n0002),
    .ADR3(DLX_MEMinst_RF_data_in[16]),
    .O(\DLX_IDinst_regA_eff<16>/FROM )
  );
  defparam \DLX_IDinst__n0086<16>20 .INIT = 16'hF000;
  X_LUT4 \DLX_IDinst__n0086<16>20  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_N70295),
    .ADR3(DLX_IDinst_regA_eff[16]),
    .O(\DLX_IDinst_regA_eff<16>/GROM )
  );
  X_BUF \DLX_IDinst_regA_eff<16>/XUSED  (
    .I(\DLX_IDinst_regA_eff<16>/FROM ),
    .O(DLX_IDinst_regA_eff[16])
  );
  X_BUF \DLX_IDinst_regA_eff<16>/YUSED  (
    .I(\DLX_IDinst_regA_eff<16>/GROM ),
    .O(CHOICE2738)
  );
  defparam \DLX_IDinst_regA_eff<24>1 .INIT = 16'hF404;
  X_LUT4 \DLX_IDinst_regA_eff<24>1  (
    .ADR0(DLX_IDinst__n0002),
    .ADR1(DLX_IDinst_reg_out_A_RF[24]),
    .ADR2(DLX_IDinst__n0144),
    .ADR3(DLX_MEMinst_RF_data_in[24]),
    .O(\DLX_IDinst_regA_eff<24>/FROM )
  );
  defparam \DLX_IDinst__n0086<24>20 .INIT = 16'hAA00;
  X_LUT4 \DLX_IDinst__n0086<24>20  (
    .ADR0(DLX_IDinst_N70295),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_regA_eff[24]),
    .O(\DLX_IDinst_regA_eff<24>/GROM )
  );
  X_BUF \DLX_IDinst_regA_eff<24>/XUSED  (
    .I(\DLX_IDinst_regA_eff<24>/FROM ),
    .O(DLX_IDinst_regA_eff[24])
  );
  X_BUF \DLX_IDinst_regA_eff<24>/YUSED  (
    .I(\DLX_IDinst_regA_eff<24>/GROM ),
    .O(CHOICE2837)
  );
  defparam \DLX_EXinst_Mshift__n0027_Sh<14>1 .INIT = 16'hCACA;
  X_LUT4 \DLX_EXinst_Mshift__n0027_Sh<14>1  (
    .ADR0(DLX_EXinst_N63449),
    .ADR1(DLX_EXinst_N62781),
    .ADR2(DLX_IDinst_IR_function_field_0_1),
    .ADR3(VCC),
    .O(\DLX_EXinst_Mshift__n0027_Sh<14>/FROM )
  );
  defparam DLX_EXinst_Ker643071.INIT = 16'hFC0C;
  X_LUT4 DLX_EXinst_Ker643071 (
    .ADR0(VCC),
    .ADR1(\DLX_EXinst_Mshift__n0027_Sh[22] ),
    .ADR2(DLX_IDinst_IR_function_field[3]),
    .ADR3(\DLX_EXinst_Mshift__n0027_Sh[14] ),
    .O(\DLX_EXinst_Mshift__n0027_Sh<14>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0027_Sh<14>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0027_Sh<14>/FROM ),
    .O(\DLX_EXinst_Mshift__n0027_Sh[14] )
  );
  X_BUF \DLX_EXinst_Mshift__n0027_Sh<14>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0027_Sh<14>/GROM ),
    .O(DLX_EXinst_N64309)
  );
  defparam \DLX_EXinst__n0006<10>117 .INIT = 16'hFFA0;
  X_LUT4 \DLX_EXinst__n0006<10>117  (
    .ADR0(DLX_EXinst__n0045),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[10]),
    .ADR3(DLX_EXinst_N64448),
    .O(\CHOICE4514/FROM )
  );
  defparam \DLX_EXinst__n0006<10>126 .INIT = 16'hAA08;
  X_LUT4 \DLX_EXinst__n0006<10>126  (
    .ADR0(DLX_IDinst_reg_out_A[10]),
    .ADR1(DLX_EXinst__n0047),
    .ADR2(DLX_IDinst_reg_out_B[10]),
    .ADR3(CHOICE4514),
    .O(\CHOICE4514/GROM )
  );
  X_BUF \CHOICE4514/XUSED  (
    .I(\CHOICE4514/FROM ),
    .O(CHOICE4514)
  );
  X_BUF \CHOICE4514/YUSED  (
    .I(\CHOICE4514/GROM ),
    .O(CHOICE4516)
  );
  defparam \DLX_IDinst_regA_eff<17>1 .INIT = 16'h88B8;
  X_LUT4 \DLX_IDinst_regA_eff<17>1  (
    .ADR0(DLX_MEMinst_RF_data_in[17]),
    .ADR1(DLX_IDinst__n0144),
    .ADR2(DLX_IDinst_reg_out_A_RF[17]),
    .ADR3(DLX_IDinst__n0002),
    .O(\DLX_IDinst_regA_eff<17>/FROM )
  );
  defparam \DLX_IDinst__n0086<17>20 .INIT = 16'hF000;
  X_LUT4 \DLX_IDinst__n0086<17>20  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_N70295),
    .ADR3(DLX_IDinst_regA_eff[17]),
    .O(\DLX_IDinst_regA_eff<17>/GROM )
  );
  X_BUF \DLX_IDinst_regA_eff<17>/XUSED  (
    .I(\DLX_IDinst_regA_eff<17>/FROM ),
    .O(DLX_IDinst_regA_eff[17])
  );
  X_BUF \DLX_IDinst_regA_eff<17>/YUSED  (
    .I(\DLX_IDinst_regA_eff<17>/GROM ),
    .O(CHOICE2749)
  );
  defparam \DLX_IDinst_regA_eff<25>1 .INIT = 16'hCC50;
  X_LUT4 \DLX_IDinst_regA_eff<25>1  (
    .ADR0(DLX_IDinst__n0002),
    .ADR1(DLX_MEMinst_RF_data_in[25]),
    .ADR2(DLX_IDinst_reg_out_A_RF[25]),
    .ADR3(DLX_IDinst__n0144),
    .O(\DLX_IDinst_regA_eff<25>/FROM )
  );
  defparam \DLX_IDinst__n0086<25>20 .INIT = 16'hF000;
  X_LUT4 \DLX_IDinst__n0086<25>20  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_N70295),
    .ADR3(DLX_IDinst_regA_eff[25]),
    .O(\DLX_IDinst_regA_eff<25>/GROM )
  );
  X_BUF \DLX_IDinst_regA_eff<25>/XUSED  (
    .I(\DLX_IDinst_regA_eff<25>/FROM ),
    .O(DLX_IDinst_regA_eff[25])
  );
  X_BUF \DLX_IDinst_regA_eff<25>/YUSED  (
    .I(\DLX_IDinst_regA_eff<25>/GROM ),
    .O(CHOICE2859)
  );
  defparam \DLX_IDinst_regA_eff<18>1 .INIT = 16'hA0E4;
  X_LUT4 \DLX_IDinst_regA_eff<18>1  (
    .ADR0(DLX_IDinst__n0144),
    .ADR1(DLX_IDinst_reg_out_A_RF[18]),
    .ADR2(DLX_MEMinst_RF_data_in[18]),
    .ADR3(DLX_IDinst__n0002),
    .O(\DLX_IDinst_regA_eff<18>/FROM )
  );
  defparam \DLX_IDinst__n0086<18>20 .INIT = 16'hF000;
  X_LUT4 \DLX_IDinst__n0086<18>20  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_N70295),
    .ADR3(DLX_IDinst_regA_eff[18]),
    .O(\DLX_IDinst_regA_eff<18>/GROM )
  );
  X_BUF \DLX_IDinst_regA_eff<18>/XUSED  (
    .I(\DLX_IDinst_regA_eff<18>/FROM ),
    .O(DLX_IDinst_regA_eff[18])
  );
  X_BUF \DLX_IDinst_regA_eff<18>/YUSED  (
    .I(\DLX_IDinst_regA_eff<18>/GROM ),
    .O(CHOICE2771)
  );
  defparam \DLX_IDinst_regA_eff<26>1 .INIT = 16'h8D88;
  X_LUT4 \DLX_IDinst_regA_eff<26>1  (
    .ADR0(DLX_IDinst__n0144),
    .ADR1(DLX_MEMinst_RF_data_in[26]),
    .ADR2(DLX_IDinst__n0002),
    .ADR3(DLX_IDinst_reg_out_A_RF[26]),
    .O(\DLX_IDinst_regA_eff<26>/FROM )
  );
  defparam \DLX_IDinst__n0086<26>20 .INIT = 16'hF000;
  X_LUT4 \DLX_IDinst__n0086<26>20  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_N70295),
    .ADR3(DLX_IDinst_regA_eff[26]),
    .O(\DLX_IDinst_regA_eff<26>/GROM )
  );
  X_BUF \DLX_IDinst_regA_eff<26>/XUSED  (
    .I(\DLX_IDinst_regA_eff<26>/FROM ),
    .O(DLX_IDinst_regA_eff[26])
  );
  X_BUF \DLX_IDinst_regA_eff<26>/YUSED  (
    .I(\DLX_IDinst_regA_eff<26>/GROM ),
    .O(CHOICE2870)
  );
  defparam DLX_IDlc_md_mda34_a1.INIT = 16'h00AA;
  X_LUT4 DLX_IDlc_md_mda34_a1 (
    .ADR0(DLX_IDlc_md_wint33),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDlc_pd_wint1),
    .O(\DLX_IDlc_md_wint34/FROM )
  );
  defparam DLX_IDlc_md_mda35_a1.INIT = 16'h5500;
  X_LUT4 DLX_IDlc_md_mda35_a1 (
    .ADR0(DLX_IDlc_pd_wint1),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDlc_md_wint34),
    .O(\DLX_IDlc_md_wint34/GROM )
  );
  X_BUF \DLX_IDlc_md_wint34/XUSED  (
    .I(\DLX_IDlc_md_wint34/FROM ),
    .O(DLX_IDlc_md_wint34)
  );
  X_BUF \DLX_IDlc_md_wint34/YUSED  (
    .I(\DLX_IDlc_md_wint34/GROM ),
    .O(DLX_IDlc_md_wint35)
  );
  defparam DLX_IDlc_md_mda26_a1.INIT = 16'h00AA;
  X_LUT4 DLX_IDlc_md_mda26_a1 (
    .ADR0(DLX_IDlc_md_wint25),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDlc_pd_wint1),
    .O(\DLX_IDlc_md_wint26/FROM )
  );
  defparam DLX_IDlc_md_mda27_a1.INIT = 16'h0F00;
  X_LUT4 DLX_IDlc_md_mda27_a1 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IDlc_pd_wint1),
    .ADR3(DLX_IDlc_md_wint26),
    .O(\DLX_IDlc_md_wint26/GROM )
  );
  X_BUF \DLX_IDlc_md_wint26/XUSED  (
    .I(\DLX_IDlc_md_wint26/FROM ),
    .O(DLX_IDlc_md_wint26)
  );
  X_BUF \DLX_IDlc_md_wint26/YUSED  (
    .I(\DLX_IDlc_md_wint26/GROM ),
    .O(DLX_IDlc_md_wint27)
  );
  defparam \DLX_EXinst__n0006<10>243 .INIT = 16'hAAA8;
  X_LUT4 \DLX_EXinst__n0006<10>243  (
    .ADR0(DLX_EXinst__n0030),
    .ADR1(CHOICE4520),
    .ADR2(CHOICE4538),
    .ADR3(CHOICE4516),
    .O(\CHOICE4540/FROM )
  );
  defparam \DLX_EXinst__n0006<10>255 .INIT = 16'hFF88;
  X_LUT4 \DLX_EXinst__n0006<10>255  (
    .ADR0(DLX_EXinst_N63836),
    .ADR1(DLX_EXinst__n0016[10]),
    .ADR2(VCC),
    .ADR3(CHOICE4540),
    .O(\CHOICE4540/GROM )
  );
  X_BUF \CHOICE4540/XUSED  (
    .I(\CHOICE4540/FROM ),
    .O(CHOICE4540)
  );
  X_BUF \CHOICE4540/YUSED  (
    .I(\CHOICE4540/GROM ),
    .O(CHOICE4541)
  );
  defparam \DLX_IDinst_regA_eff<19>1 .INIT = 16'hCC0A;
  X_LUT4 \DLX_IDinst_regA_eff<19>1  (
    .ADR0(DLX_IDinst_reg_out_A_RF[19]),
    .ADR1(DLX_MEMinst_RF_data_in[19]),
    .ADR2(DLX_IDinst__n0002),
    .ADR3(DLX_IDinst__n0144),
    .O(\DLX_IDinst_regA_eff<19>/FROM )
  );
  defparam DLX_IDinst__n0146102.INIT = 16'h0001;
  X_LUT4 DLX_IDinst__n0146102 (
    .ADR0(DLX_IDinst_regA_eff[17]),
    .ADR1(DLX_IDinst_regA_eff[18]),
    .ADR2(DLX_IDinst_regA_eff[16]),
    .ADR3(DLX_IDinst_regA_eff[19]),
    .O(\DLX_IDinst_regA_eff<19>/GROM )
  );
  X_BUF \DLX_IDinst_regA_eff<19>/XUSED  (
    .I(\DLX_IDinst_regA_eff<19>/FROM ),
    .O(DLX_IDinst_regA_eff[19])
  );
  X_BUF \DLX_IDinst_regA_eff<19>/YUSED  (
    .I(\DLX_IDinst_regA_eff<19>/GROM ),
    .O(CHOICE3651)
  );
  defparam \DLX_IDinst_regA_eff<27>1 .INIT = 16'hA0AC;
  X_LUT4 \DLX_IDinst_regA_eff<27>1  (
    .ADR0(DLX_MEMinst_RF_data_in[27]),
    .ADR1(DLX_IDinst_reg_out_A_RF[27]),
    .ADR2(DLX_IDinst__n0144),
    .ADR3(DLX_IDinst__n0002),
    .O(\DLX_IDinst_regA_eff<27>/FROM )
  );
  defparam DLX_IDinst__n0146139.INIT = 16'h0001;
  X_LUT4 DLX_IDinst__n0146139 (
    .ADR0(DLX_IDinst_regA_eff[25]),
    .ADR1(DLX_IDinst_regA_eff[24]),
    .ADR2(DLX_IDinst_regA_eff[26]),
    .ADR3(DLX_IDinst_regA_eff[27]),
    .O(\DLX_IDinst_regA_eff<27>/GROM )
  );
  X_BUF \DLX_IDinst_regA_eff<27>/XUSED  (
    .I(\DLX_IDinst_regA_eff<27>/FROM ),
    .O(DLX_IDinst_regA_eff[27])
  );
  X_BUF \DLX_IDinst_regA_eff<27>/YUSED  (
    .I(\DLX_IDinst_regA_eff<27>/GROM ),
    .O(CHOICE3666)
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<61>1 .INIT = 16'h50F0;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<61>1  (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(DLX_IDinst_reg_out_B[0]),
    .O(\DLX_EXinst_Mshift__n0023_Sh<61>/FROM )
  );
  defparam DLX_EXinst_Ker6482713.INIT = 16'hEC4C;
  X_LUT4 DLX_EXinst_Ker6482713 (
    .ADR0(DLX_IDinst_reg_out_B_2_1),
    .ADR1(DLX_IDinst_reg_out_A[31]),
    .ADR2(DLX_IDinst_reg_out_B_3_1),
    .ADR3(\DLX_EXinst_Mshift__n0023_Sh[61] ),
    .O(\DLX_EXinst_Mshift__n0023_Sh<61>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0023_Sh<61>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0023_Sh<61>/FROM ),
    .O(\DLX_EXinst_Mshift__n0023_Sh[61] )
  );
  X_BUF \DLX_EXinst_Mshift__n0023_Sh<61>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0023_Sh<61>/GROM ),
    .O(CHOICE1919)
  );
  defparam \DLX_EXinst__n0006<10>184 .INIT = 16'hF000;
  X_LUT4 \DLX_EXinst__n0006<10>184  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(\DLX_EXinst_Mshift__n0025_Sh[42] ),
    .ADR3(DLX_EXinst_N66226),
    .O(\CHOICE4532/FROM )
  );
  defparam \DLX_EXinst__n0006<10>217 .INIT = 16'hCFCE;
  X_LUT4 \DLX_EXinst__n0006<10>217  (
    .ADR0(CHOICE4531),
    .ADR1(CHOICE4537),
    .ADR2(DLX_IDinst_reg_out_B[4]),
    .ADR3(CHOICE4532),
    .O(\CHOICE4532/GROM )
  );
  X_BUF \CHOICE4532/XUSED  (
    .I(\CHOICE4532/FROM ),
    .O(CHOICE4532)
  );
  X_BUF \CHOICE4532/YUSED  (
    .I(\CHOICE4532/GROM ),
    .O(CHOICE4538)
  );
  defparam \DLX_IDinst_regA_eff<28>1 .INIT = 16'hA0AC;
  X_LUT4 \DLX_IDinst_regA_eff<28>1  (
    .ADR0(DLX_MEMinst_RF_data_in[28]),
    .ADR1(DLX_IDinst_reg_out_A_RF[28]),
    .ADR2(DLX_IDinst__n0144),
    .ADR3(DLX_IDinst__n0002),
    .O(\DLX_IDinst_regA_eff<28>/FROM )
  );
  defparam \DLX_IDinst__n0086<28>20 .INIT = 16'hF000;
  X_LUT4 \DLX_IDinst__n0086<28>20  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_N70295),
    .ADR3(DLX_IDinst_regA_eff[28]),
    .O(\DLX_IDinst_regA_eff<28>/GROM )
  );
  X_BUF \DLX_IDinst_regA_eff<28>/XUSED  (
    .I(\DLX_IDinst_regA_eff<28>/FROM ),
    .O(DLX_IDinst_regA_eff[28])
  );
  X_BUF \DLX_IDinst_regA_eff<28>/YUSED  (
    .I(\DLX_IDinst_regA_eff<28>/GROM ),
    .O(CHOICE2892)
  );
  defparam \DLX_EXinst__n0006<19>109_SW0 .INIT = 16'hFF88;
  X_LUT4 \DLX_EXinst__n0006<19>109_SW0  (
    .ADR0(DLX_EXinst__n0082),
    .ADR1(\DLX_EXinst_Mshift__n0028_Sh[51] ),
    .ADR2(VCC),
    .ADR3(CHOICE4965),
    .O(\N126564/FROM )
  );
  defparam \DLX_EXinst__n0006<19>109 .INIT = 16'hD5C0;
  X_LUT4 \DLX_EXinst__n0006<19>109  (
    .ADR0(N109130),
    .ADR1(N101537),
    .ADR2(N110065),
    .ADR3(N126564),
    .O(\N126564/GROM )
  );
  X_BUF \N126564/XUSED  (
    .I(\N126564/FROM ),
    .O(N126564)
  );
  X_BUF \N126564/YUSED  (
    .I(\N126564/GROM ),
    .O(CHOICE4970)
  );
  defparam \DLX_EXinst__n0006<10>283 .INIT = 16'hAA08;
  X_LUT4 \DLX_EXinst__n0006<10>283  (
    .ADR0(DLX_EXinst__n0149),
    .ADR1(CHOICE4508),
    .ADR2(DLX_EXinst__n0030),
    .ADR3(CHOICE4541),
    .O(\DLX_EXinst_ALU_result<10>/FROM )
  );
  defparam \DLX_EXinst__n0006<10>293 .INIT = 16'hFFAA;
  X_LUT4 \DLX_EXinst__n0006<10>293  (
    .ADR0(DLX_EXinst_N63689),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(CHOICE4543),
    .O(\DLX_EXinst_ALU_result<10>/GROM )
  );
  X_BUF \DLX_EXinst_ALU_result<10>/XUSED  (
    .I(\DLX_EXinst_ALU_result<10>/FROM ),
    .O(CHOICE4543)
  );
  X_BUF \DLX_EXinst_ALU_result<10>/YUSED  (
    .I(\DLX_EXinst_ALU_result<10>/GROM ),
    .O(N116776)
  );
  defparam \DLX_EXinst__n0006<11>117 .INIT = 16'hF8F8;
  X_LUT4 \DLX_EXinst__n0006<11>117  (
    .ADR0(DLX_IDinst_reg_out_B[11]),
    .ADR1(DLX_EXinst__n0045),
    .ADR2(DLX_EXinst_N64448),
    .ADR3(VCC),
    .O(\CHOICE3944/FROM )
  );
  defparam \DLX_EXinst__n0006<11>126 .INIT = 16'hF400;
  X_LUT4 \DLX_EXinst__n0006<11>126  (
    .ADR0(DLX_IDinst_reg_out_B[11]),
    .ADR1(DLX_EXinst__n0047),
    .ADR2(CHOICE3944),
    .ADR3(DLX_IDinst_reg_out_A[11]),
    .O(\CHOICE3944/GROM )
  );
  X_BUF \CHOICE3944/XUSED  (
    .I(\CHOICE3944/FROM ),
    .O(CHOICE3944)
  );
  X_BUF \CHOICE3944/YUSED  (
    .I(\CHOICE3944/GROM ),
    .O(CHOICE3946)
  );
  defparam \DLX_IDinst_regA_eff<29>1 .INIT = 16'hA0E4;
  X_LUT4 \DLX_IDinst_regA_eff<29>1  (
    .ADR0(DLX_IDinst__n0144),
    .ADR1(DLX_IDinst_reg_out_A_RF[29]),
    .ADR2(DLX_MEMinst_RF_data_in[29]),
    .ADR3(DLX_IDinst__n0002),
    .O(\DLX_IDinst_regA_eff<29>/FROM )
  );
  defparam \DLX_IDinst__n0086<29>20 .INIT = 16'hAA00;
  X_LUT4 \DLX_IDinst__n0086<29>20  (
    .ADR0(DLX_IDinst_N70295),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_regA_eff[29]),
    .O(\DLX_IDinst_regA_eff<29>/GROM )
  );
  X_BUF \DLX_IDinst_regA_eff<29>/XUSED  (
    .I(\DLX_IDinst_regA_eff<29>/FROM ),
    .O(DLX_IDinst_regA_eff[29])
  );
  X_BUF \DLX_IDinst_regA_eff<29>/YUSED  (
    .I(\DLX_IDinst_regA_eff<29>/GROM ),
    .O(CHOICE2903)
  );
  defparam \DLX_IFinst__n0001<30>_SW0 .INIT = 16'h5353;
  X_LUT4 \DLX_IFinst__n0001<30>_SW0  (
    .ADR0(DLX_IFinst_PC[30]),
    .ADR1(DLX_IFinst__n0015[30]),
    .ADR2(DLX_IFinst__n0000),
    .ADR3(VCC),
    .O(\DLX_IFinst_NPC<30>/FROM )
  );
  defparam \DLX_IFinst__n0001<30> .INIT = 16'hA0AF;
  X_LUT4 \DLX_IFinst__n0001<30>  (
    .ADR0(DLX_IDinst_branch_address[30]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(N91619),
    .O(DLX_IFinst__n0001[30])
  );
  X_BUF \DLX_IFinst_NPC<30>/XUSED  (
    .I(\DLX_IFinst_NPC<30>/FROM ),
    .O(N91619)
  );
  defparam \DLX_IFinst__n0001<14>_SW0 .INIT = 16'h05F5;
  X_LUT4 \DLX_IFinst__n0001<14>_SW0  (
    .ADR0(DLX_IFinst__n0015[14]),
    .ADR1(VCC),
    .ADR2(DLX_IFinst__n0000),
    .ADR3(DLX_IFinst_PC[14]),
    .O(\DLX_IFinst_NPC<14>/FROM )
  );
  defparam \DLX_IFinst__n0001<14> .INIT = 16'hA0AF;
  X_LUT4 \DLX_IFinst__n0001<14>  (
    .ADR0(DLX_IDinst_branch_address[14]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(N92399),
    .O(\DLX_IFinst_NPC<14>/GROM )
  );
  X_BUF \DLX_IFinst_NPC<14>/XUSED  (
    .I(\DLX_IFinst_NPC<14>/FROM ),
    .O(N92399)
  );
  X_BUF \DLX_IFinst_NPC<14>/YUSED  (
    .I(\DLX_IFinst_NPC<14>/GROM ),
    .O(DLX_IFinst__n0001[14])
  );
  defparam \DLX_IFinst__n0001<22>_SW0 .INIT = 16'h5353;
  X_LUT4 \DLX_IFinst__n0001<22>_SW0  (
    .ADR0(DLX_IFinst_PC[22]),
    .ADR1(DLX_IFinst__n0015[22]),
    .ADR2(DLX_IFinst__n0000),
    .ADR3(VCC),
    .O(\DLX_IFinst_NPC<22>/FROM )
  );
  defparam \DLX_IFinst__n0001<22> .INIT = 16'hC0F3;
  X_LUT4 \DLX_IFinst__n0001<22>  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(DLX_IDinst_branch_address[22]),
    .ADR3(N92035),
    .O(DLX_IFinst__n0001[22])
  );
  X_BUF \DLX_IFinst_NPC<22>/XUSED  (
    .I(\DLX_IFinst_NPC<22>/FROM ),
    .O(N92035)
  );
  defparam \DLX_EXinst__n0006<11>214 .INIT = 16'hCCC8;
  X_LUT4 \DLX_EXinst__n0006<11>214  (
    .ADR0(CHOICE3950),
    .ADR1(DLX_EXinst__n0030),
    .ADR2(CHOICE3946),
    .ADR3(CHOICE3964),
    .O(\CHOICE3966/FROM )
  );
  defparam \DLX_EXinst__n0006<11>226 .INIT = 16'hFFC0;
  X_LUT4 \DLX_EXinst__n0006<11>226  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst__n0016[11]),
    .ADR2(DLX_EXinst_N63836),
    .ADR3(CHOICE3966),
    .O(\CHOICE3966/GROM )
  );
  X_BUF \CHOICE3966/XUSED  (
    .I(\CHOICE3966/FROM ),
    .O(CHOICE3966)
  );
  X_BUF \CHOICE3966/YUSED  (
    .I(\CHOICE3966/GROM ),
    .O(CHOICE3967)
  );
  defparam DLX_IDinst__n0108160_SW0.INIT = 16'hFFEC;
  X_LUT4 DLX_IDinst__n0108160_SW0 (
    .ADR0(DLX_IDinst__n0448[1]),
    .ADR1(CHOICE3460),
    .ADR2(CHOICE3448),
    .ADR3(CHOICE3458),
    .O(\DLX_IDinst_reg_dst/FROM )
  );
  defparam DLX_IDinst__n0108160.INIT = 16'h4000;
  X_LUT4 DLX_IDinst__n0108160 (
    .ADR0(DLX_IDinst_intr_slot),
    .ADR1(DLX_EXinst__n0149),
    .ADR2(N95693),
    .ADR3(N126807),
    .O(N110380)
  );
  X_BUF \DLX_IDinst_reg_dst/XUSED  (
    .I(\DLX_IDinst_reg_dst/FROM ),
    .O(N126807)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_inv_01.INIT = 16'h50F5;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_inv_01 (
    .ADR0(DLX_EXinst_Mcompar__n0093_inst_cy_228),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(DLX_IDinst_Imm_31_1),
    .O(\DLX_EXinst__n0093/FROM )
  );
  defparam \DLX_EXinst__n0006<0>407 .INIT = 16'h0E02;
  X_LUT4 \DLX_EXinst__n0006<0>407  (
    .ADR0(DLX_EXinst__n0085),
    .ADR1(DLX_IDinst_IR_opcode_field[2]),
    .ADR2(DLX_IDinst_IR_opcode_field[0]),
    .ADR3(DLX_EXinst__n0093),
    .O(\DLX_EXinst__n0093/GROM )
  );
  X_BUF \DLX_EXinst__n0093/XUSED  (
    .I(\DLX_EXinst__n0093/FROM ),
    .O(DLX_EXinst__n0093)
  );
  X_BUF \DLX_EXinst__n0093/YUSED  (
    .I(\DLX_EXinst__n0093/GROM ),
    .O(CHOICE5934)
  );
  defparam \DLX_EXinst__n0006<27>158 .INIT = 16'hC4C0;
  X_LUT4 \DLX_EXinst__n0006<27>158  (
    .ADR0(DLX_IDinst_reg_out_A[27]),
    .ADR1(DLX_IDinst_reg_out_B[27]),
    .ADR2(DLX_EXinst__n0046),
    .ADR3(DLX_EXinst__n0047),
    .O(\CHOICE4643/FROM )
  );
  defparam \DLX_EXinst__n0006<11>138 .INIT = 16'hF400;
  X_LUT4 \DLX_EXinst__n0006<11>138  (
    .ADR0(DLX_IDinst_reg_out_A[11]),
    .ADR1(DLX_EXinst__n0047),
    .ADR2(DLX_EXinst__n0046),
    .ADR3(DLX_IDinst_reg_out_B[11]),
    .O(\CHOICE4643/GROM )
  );
  X_BUF \CHOICE4643/XUSED  (
    .I(\CHOICE4643/FROM ),
    .O(CHOICE4643)
  );
  X_BUF \CHOICE4643/YUSED  (
    .I(\CHOICE4643/GROM ),
    .O(CHOICE3950)
  );
  defparam DLX_IDlc_md_mda8_a1.INIT = 16'h0A0A;
  X_LUT4 DLX_IDlc_md_mda8_a1 (
    .ADR0(DLX_IDlc_md_wint7),
    .ADR1(VCC),
    .ADR2(DLX_IDlc_pd_wint1),
    .ADR3(VCC),
    .O(\DLX_IDlc_md_wint8/FROM )
  );
  defparam DLX_IDlc_md_mda36_a1.INIT = 16'h5050;
  X_LUT4 DLX_IDlc_md_mda36_a1 (
    .ADR0(DLX_IDlc_pd_wint1),
    .ADR1(VCC),
    .ADR2(DLX_IDlc_md_wint35),
    .ADR3(VCC),
    .O(\DLX_IDlc_md_wint8/GROM )
  );
  X_BUF \DLX_IDlc_md_wint8/XUSED  (
    .I(\DLX_IDlc_md_wint8/FROM ),
    .O(DLX_IDlc_md_wint8)
  );
  X_BUF \DLX_IDlc_md_wint8/YUSED  (
    .I(\DLX_IDlc_md_wint8/GROM ),
    .O(DLX_IDlc_md_wint36)
  );
  defparam \DLX_EXinst__n0006<18>207 .INIT = 16'h2000;
  X_LUT4 \DLX_EXinst__n0006<18>207  (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(DLX_EXinst_N62740),
    .ADR2(\DLX_EXinst_Mshift__n0025_Sh[2] ),
    .ADR3(DLX_EXinst_N66226),
    .O(\CHOICE5451/FROM )
  );
  defparam \DLX_EXinst__n0006<11>164 .INIT = 16'hF000;
  X_LUT4 \DLX_EXinst__n0006<11>164  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(\DLX_EXinst_Mshift__n0025_Sh[43] ),
    .ADR3(DLX_EXinst_N66226),
    .O(\CHOICE5451/GROM )
  );
  X_BUF \CHOICE5451/XUSED  (
    .I(\CHOICE5451/FROM ),
    .O(CHOICE5451)
  );
  X_BUF \CHOICE5451/YUSED  (
    .I(\CHOICE5451/GROM ),
    .O(CHOICE3958)
  );
  defparam \DLX_EXinst__n0006<11>254 .INIT = 16'hCE00;
  X_LUT4 \DLX_EXinst__n0006<11>254  (
    .ADR0(CHOICE3938),
    .ADR1(CHOICE3967),
    .ADR2(DLX_EXinst__n0030),
    .ADR3(DLX_EXinst__n0149),
    .O(\DLX_EXinst_ALU_result<11>/FROM )
  );
  defparam \DLX_EXinst__n0006<11>264 .INIT = 16'hFFF0;
  X_LUT4 \DLX_EXinst__n0006<11>264  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N63689),
    .ADR3(CHOICE3969),
    .O(\DLX_EXinst_ALU_result<11>/GROM )
  );
  X_BUF \DLX_EXinst_ALU_result<11>/XUSED  (
    .I(\DLX_EXinst_ALU_result<11>/FROM ),
    .O(CHOICE3969)
  );
  X_BUF \DLX_EXinst_ALU_result<11>/YUSED  (
    .I(\DLX_EXinst_ALU_result<11>/GROM ),
    .O(N113314)
  );
  defparam \DLX_IFinst__n0001<2>_SW0 .INIT = 16'h33AA;
  X_LUT4 \DLX_IFinst__n0001<2>_SW0  (
    .ADR0(DLX_IFinst_NPC[2]),
    .ADR1(DLX_IFinst_PC[2]),
    .ADR2(VCC),
    .ADR3(DLX_IFinst__n0000),
    .O(\DLX_IFinst_NPC<2>/FROM )
  );
  defparam \DLX_IFinst__n0001<2> .INIT = 16'hA0F5;
  X_LUT4 \DLX_IFinst__n0001<2>  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_branch_address[2]),
    .ADR3(N93023),
    .O(\DLX_IFinst_NPC<2>/GROM )
  );
  X_BUF \DLX_IFinst_NPC<2>/XUSED  (
    .I(\DLX_IFinst_NPC<2>/FROM ),
    .O(N93023)
  );
  X_BUF \DLX_IFinst_NPC<2>/YUSED  (
    .I(\DLX_IFinst_NPC<2>/GROM ),
    .O(DLX_IFinst__n0001[2])
  );
  defparam \DLX_EXinst__n0006<11>185 .INIT = 16'hEAC0;
  X_LUT4 \DLX_EXinst__n0006<11>185  (
    .ADR0(DLX_EXinst_ALU_result[11]),
    .ADR1(DLX_IDinst_reg_out_B[4]),
    .ADR2(N105035),
    .ADR3(N101725),
    .O(\CHOICE3963/FROM )
  );
  defparam \DLX_EXinst__n0006<11>189 .INIT = 16'hFF32;
  X_LUT4 \DLX_EXinst__n0006<11>189  (
    .ADR0(CHOICE3957),
    .ADR1(DLX_IDinst_reg_out_B[4]),
    .ADR2(CHOICE3958),
    .ADR3(CHOICE3963),
    .O(\CHOICE3963/GROM )
  );
  X_BUF \CHOICE3963/XUSED  (
    .I(\CHOICE3963/FROM ),
    .O(CHOICE3963)
  );
  X_BUF \CHOICE3963/YUSED  (
    .I(\CHOICE3963/GROM ),
    .O(CHOICE3964)
  );
  defparam DLX_IDlc_md_mda7_a1.INIT = 16'h0F00;
  X_LUT4 DLX_IDlc_md_mda7_a1 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IDlc_pd_wint1),
    .ADR3(DLX_IDlc_md_wint6),
    .O(\DLX_IDlc_md_wint7/FROM )
  );
  defparam DLX_IDlc_md_mda37_a1.INIT = 16'h0C0C;
  X_LUT4 DLX_IDlc_md_mda37_a1 (
    .ADR0(VCC),
    .ADR1(DLX_IDlc_md_wint36),
    .ADR2(DLX_IDlc_pd_wint1),
    .ADR3(VCC),
    .O(\DLX_IDlc_md_wint7/GROM )
  );
  X_BUF \DLX_IDlc_md_wint7/XUSED  (
    .I(\DLX_IDlc_md_wint7/FROM ),
    .O(DLX_IDlc_md_wint7)
  );
  X_BUF \DLX_IDlc_md_wint7/YUSED  (
    .I(\DLX_IDlc_md_wint7/GROM ),
    .O(DLX_IDlc_md_wint37)
  );
  defparam \DLX_EXinst__n0006<30>335 .INIT = 16'hF888;
  X_LUT4 \DLX_EXinst__n0006<30>335  (
    .ADR0(DLX_EXinst_N63712),
    .ADR1(DLX_IDinst_reg_out_A[27]),
    .ADR2(DLX_EXinst__n0030),
    .ADR3(N126519),
    .O(\CHOICE5321/FROM )
  );
  defparam \DLX_EXinst__n0006<30>367_SW0 .INIT = 16'hFFCE;
  X_LUT4 \DLX_EXinst__n0006<30>367_SW0  (
    .ADR0(CHOICE5279),
    .ADR1(CHOICE5324),
    .ADR2(DLX_EXinst__n0030),
    .ADR3(CHOICE5321),
    .O(\CHOICE5321/GROM )
  );
  X_BUF \CHOICE5321/XUSED  (
    .I(\CHOICE5321/FROM ),
    .O(CHOICE5321)
  );
  X_BUF \CHOICE5321/YUSED  (
    .I(\CHOICE5321/GROM ),
    .O(N126514)
  );
  defparam \DLX_EXinst__n0006<20>310 .INIT = 16'hEECC;
  X_LUT4 \DLX_EXinst__n0006<20>310  (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(CHOICE4934),
    .ADR2(VCC),
    .ADR3(CHOICE1771),
    .O(\DLX_EXinst_ALU_result<20>/FROM )
  );
  defparam \DLX_EXinst__n0006<20>336 .INIT = 16'h0302;
  X_LUT4 \DLX_EXinst__n0006<20>336  (
    .ADR0(N127200),
    .ADR1(DLX_IDinst_counter[1]),
    .ADR2(DLX_IDinst_counter[0]),
    .ADR3(CHOICE4935),
    .O(N119151)
  );
  X_BUF \DLX_EXinst_ALU_result<20>/XUSED  (
    .I(\DLX_EXinst_ALU_result<20>/FROM ),
    .O(CHOICE4935)
  );
  defparam \DLX_EXinst_Mshift__n0027_Sh<3>25 .INIT = 16'h00AC;
  X_LUT4 \DLX_EXinst_Mshift__n0027_Sh<3>25  (
    .ADR0(DLX_IDinst_reg_out_A[2]),
    .ADR1(DLX_IDinst_reg_out_A[3]),
    .ADR2(DLX_IDinst_IR_function_field_0_1),
    .ADR3(DLX_IDinst_IR_function_field_1_1),
    .O(\CHOICE1000/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0027_Sh<3>28 .INIT = 16'hFFCC;
  X_LUT4 \DLX_EXinst_Mshift__n0027_Sh<3>28  (
    .ADR0(VCC),
    .ADR1(CHOICE994),
    .ADR2(VCC),
    .ADR3(CHOICE1000),
    .O(\CHOICE1000/GROM )
  );
  X_BUF \CHOICE1000/XUSED  (
    .I(\CHOICE1000/FROM ),
    .O(CHOICE1000)
  );
  X_BUF \CHOICE1000/YUSED  (
    .I(\CHOICE1000/GROM ),
    .O(\DLX_EXinst_Mshift__n0027_Sh[3] )
  );
  defparam \DLX_EXinst__n0006<18>199 .INIT = 16'hAE00;
  X_LUT4 \DLX_EXinst__n0006<18>199  (
    .ADR0(DLX_EXinst__n0046),
    .ADR1(DLX_EXinst__n0047),
    .ADR2(DLX_IDinst_reg_out_A[18]),
    .ADR3(DLX_IDinst_reg_out_B[18]),
    .O(\CHOICE5447/FROM )
  );
  defparam \DLX_EXinst__n0006<12>119 .INIT = 16'hC0C8;
  X_LUT4 \DLX_EXinst__n0006<12>119  (
    .ADR0(DLX_EXinst__n0047),
    .ADR1(DLX_IDinst_reg_out_B[12]),
    .ADR2(DLX_EXinst__n0046),
    .ADR3(DLX_IDinst_reg_out_A[12]),
    .O(\CHOICE5447/GROM )
  );
  X_BUF \CHOICE5447/XUSED  (
    .I(\CHOICE5447/FROM ),
    .O(CHOICE5447)
  );
  X_BUF \CHOICE5447/YUSED  (
    .I(\CHOICE5447/GROM ),
    .O(CHOICE3884)
  );
  defparam \DLX_IDinst_slot_num_FFd2-In23 .INIT = 16'h0400;
  X_LUT4 \DLX_IDinst_slot_num_FFd2-In23  (
    .ADR0(DLX_IDinst_CLI),
    .ADR1(INT_IBUF),
    .ADR2(DLX_IDinst_delay_slot),
    .ADR3(DLX_IDinst_N70077),
    .O(\CHOICE2521/FROM )
  );
  defparam \DLX_IDinst_slot_num_FFd2-In37 .INIT = 16'h0F08;
  X_LUT4 \DLX_IDinst_slot_num_FFd2-In37  (
    .ADR0(CHOICE2516),
    .ADR1(N109350),
    .ADR2(FREEZE_IBUF),
    .ADR3(CHOICE2521),
    .O(\CHOICE2521/GROM )
  );
  X_BUF \CHOICE2521/XUSED  (
    .I(\CHOICE2521/FROM ),
    .O(CHOICE2521)
  );
  X_BUF \CHOICE2521/YUSED  (
    .I(\CHOICE2521/GROM ),
    .O(CHOICE2523)
  );
  defparam \DLX_EXinst__n0006<20>231 .INIT = 16'h4400;
  X_LUT4 \DLX_EXinst__n0006<20>231  (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(DLX_EXinst__n0049),
    .ADR2(VCC),
    .ADR3(\DLX_EXinst_Mshift__n0026_Sh[52] ),
    .O(\CHOICE4928/FROM )
  );
  defparam \DLX_EXinst__n0006<20>248 .INIT = 16'h0F08;
  X_LUT4 \DLX_EXinst__n0006<20>248  (
    .ADR0(DLX_EXinst__n0048),
    .ADR1(CHOICE4926),
    .ADR2(N110935),
    .ADR3(CHOICE4928),
    .O(\CHOICE4928/GROM )
  );
  X_BUF \CHOICE4928/XUSED  (
    .I(\CHOICE4928/FROM ),
    .O(CHOICE4928)
  );
  X_BUF \CHOICE4928/YUSED  (
    .I(\CHOICE4928/GROM ),
    .O(CHOICE4930)
  );
  defparam \DLX_EXinst__n0006<12>216 .INIT = 16'hF0E0;
  X_LUT4 \DLX_EXinst__n0006<12>216  (
    .ADR0(CHOICE3906),
    .ADR1(CHOICE3889),
    .ADR2(DLX_EXinst__n0030),
    .ADR3(CHOICE3884),
    .O(\CHOICE3908/FROM )
  );
  defparam \DLX_EXinst__n0006<12>228 .INIT = 16'hFFA0;
  X_LUT4 \DLX_EXinst__n0006<12>228  (
    .ADR0(DLX_EXinst_N63836),
    .ADR1(VCC),
    .ADR2(DLX_EXinst__n0016[12]),
    .ADR3(CHOICE3908),
    .O(\CHOICE3908/GROM )
  );
  X_BUF \CHOICE3908/XUSED  (
    .I(\CHOICE3908/FROM ),
    .O(CHOICE3908)
  );
  X_BUF \CHOICE3908/YUSED  (
    .I(\CHOICE3908/GROM ),
    .O(CHOICE3909)
  );
  defparam \DLX_EXinst_Mshift__n0024_Sh<26>26 .INIT = 16'h00CA;
  X_LUT4 \DLX_EXinst_Mshift__n0024_Sh<26>26  (
    .ADR0(DLX_IDinst_reg_out_A[26]),
    .ADR1(DLX_IDinst_reg_out_A[28]),
    .ADR2(DLX_IDinst_IR_function_field_1_1),
    .ADR3(DLX_IDinst_IR_function_field_0_1),
    .O(\CHOICE1120/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0027_Sh<4>11 .INIT = 16'hA088;
  X_LUT4 \DLX_EXinst_Mshift__n0027_Sh<4>11  (
    .ADR0(DLX_IDinst_IR_function_field_1_1),
    .ADR1(DLX_IDinst_reg_out_A[2]),
    .ADR2(DLX_IDinst_reg_out_A[1]),
    .ADR3(DLX_IDinst_IR_function_field_0_1),
    .O(\CHOICE1120/GROM )
  );
  X_BUF \CHOICE1120/XUSED  (
    .I(\CHOICE1120/FROM ),
    .O(CHOICE1120)
  );
  X_BUF \CHOICE1120/YUSED  (
    .I(\CHOICE1120/GROM ),
    .O(CHOICE1006)
  );
  defparam \DLX_EXinst__n0006<20>208 .INIT = 16'h2230;
  X_LUT4 \DLX_EXinst__n0006<20>208  (
    .ADR0(DLX_EXinst_N64914),
    .ADR1(DLX_IDinst_reg_out_B[4]),
    .ADR2(DLX_EXinst_N63925),
    .ADR3(DLX_IDinst_reg_out_B[2]),
    .O(\CHOICE4925/FROM )
  );
  defparam \DLX_EXinst__n0006<20>213 .INIT = 16'hFF40;
  X_LUT4 \DLX_EXinst__n0006<20>213  (
    .ADR0(DLX_IDinst_reg_out_B[3]),
    .ADR1(DLX_IDinst_reg_out_B[4]),
    .ADR2(DLX_EXinst_N62901),
    .ADR3(CHOICE4925),
    .O(\CHOICE4925/GROM )
  );
  X_BUF \CHOICE4925/XUSED  (
    .I(\CHOICE4925/FROM ),
    .O(CHOICE4925)
  );
  X_BUF \CHOICE4925/YUSED  (
    .I(\CHOICE4925/GROM ),
    .O(CHOICE4926)
  );
  defparam DLX_IDlc_md_mda6_a1.INIT = 16'h00AA;
  X_LUT4 DLX_IDlc_md_mda6_a1 (
    .ADR0(DLX_IDlc_md_wint5),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDlc_pd_wint1),
    .O(\DLX_IDlc_md_wint6/FROM )
  );
  defparam DLX_IDlc_md_mda38_a1.INIT = 16'h00CC;
  X_LUT4 DLX_IDlc_md_mda38_a1 (
    .ADR0(VCC),
    .ADR1(DLX_IDlc_md_wint37),
    .ADR2(VCC),
    .ADR3(DLX_IDlc_pd_wint1),
    .O(\DLX_IDlc_md_wint6/GROM )
  );
  X_BUF \DLX_IDlc_md_wint6/XUSED  (
    .I(\DLX_IDlc_md_wint6/FROM ),
    .O(DLX_IDlc_md_wint6)
  );
  X_BUF \DLX_IDlc_md_wint6/YUSED  (
    .I(\DLX_IDlc_md_wint6/GROM ),
    .O(DLX_IDlc_md_wint38)
  );
  defparam \DLX_EXinst__n0006<22>213 .INIT = 16'hF888;
  X_LUT4 \DLX_EXinst__n0006<22>213  (
    .ADR0(DLX_EXinst__n0114),
    .ADR1(DLX_EXinst__n0016[22]),
    .ADR2(N101725),
    .ADR3(DLX_EXinst_ALU_result[22]),
    .O(\CHOICE4145/FROM )
  );
  defparam \DLX_EXinst__n0006<20>170 .INIT = 16'hEAC0;
  X_LUT4 \DLX_EXinst__n0006<20>170  (
    .ADR0(DLX_EXinst_ALU_result[20]),
    .ADR1(DLX_EXinst__n0114),
    .ADR2(DLX_EXinst__n0016[20]),
    .ADR3(N101725),
    .O(\CHOICE4145/GROM )
  );
  X_BUF \CHOICE4145/XUSED  (
    .I(\CHOICE4145/FROM ),
    .O(CHOICE4145)
  );
  X_BUF \CHOICE4145/YUSED  (
    .I(\CHOICE4145/GROM ),
    .O(CHOICE4909)
  );
  defparam \DLX_EXinst__n0006<23>100 .INIT = 16'hFFF8;
  X_LUT4 \DLX_EXinst__n0006<23>100  (
    .ADR0(DLX_EXinst__n0016[23]),
    .ADR1(DLX_EXinst__n0128),
    .ADR2(CHOICE4053),
    .ADR3(N126593),
    .O(\CHOICE4057/FROM )
  );
  defparam \DLX_EXinst__n0006<21>100 .INIT = 16'hFFF8;
  X_LUT4 \DLX_EXinst__n0006<21>100  (
    .ADR0(DLX_EXinst__n0016[21]),
    .ADR1(DLX_EXinst__n0128),
    .ADR2(N126451),
    .ADR3(CHOICE4185),
    .O(\CHOICE4057/GROM )
  );
  X_BUF \CHOICE4057/XUSED  (
    .I(\CHOICE4057/FROM ),
    .O(CHOICE4057)
  );
  X_BUF \CHOICE4057/YUSED  (
    .I(\CHOICE4057/GROM ),
    .O(CHOICE4189)
  );
  defparam \DLX_EXinst__n0006<12>149 .INIT = 16'hEAEA;
  X_LUT4 \DLX_EXinst__n0006<12>149  (
    .ADR0(DLX_EXinst_N64448),
    .ADR1(DLX_EXinst__n0045),
    .ADR2(DLX_IDinst_reg_out_B[12]),
    .ADR3(VCC),
    .O(\CHOICE3895/FROM )
  );
  defparam \DLX_EXinst__n0006<12>158 .INIT = 16'hCC40;
  X_LUT4 \DLX_EXinst__n0006<12>158  (
    .ADR0(DLX_IDinst_reg_out_B[12]),
    .ADR1(DLX_IDinst_reg_out_A[12]),
    .ADR2(DLX_EXinst__n0047),
    .ADR3(CHOICE3895),
    .O(\CHOICE3895/GROM )
  );
  X_BUF \CHOICE3895/XUSED  (
    .I(\CHOICE3895/FROM ),
    .O(CHOICE3895)
  );
  X_BUF \CHOICE3895/YUSED  (
    .I(\CHOICE3895/GROM ),
    .O(CHOICE3897)
  );
  defparam \Mshift__n0000_Sh<32>1 .INIT = 16'h0011;
  X_LUT4 \Mshift__n0000_Sh<32>1  (
    .ADR0(DLX_EXinst_ALU_result[14]),
    .ADR1(DLX_EXinst_ALU_result[13]),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_ALU_result[12]),
    .O(\vga_select_6<0>/FROM )
  );
  defparam \DLX_EXinst__n0006<12>190 .INIT = 16'hFEFA;
  X_LUT4 \DLX_EXinst__n0006<12>190  (
    .ADR0(CHOICE3897),
    .ADR1(N101725),
    .ADR2(CHOICE3905),
    .ADR3(DLX_EXinst_ALU_result[12]),
    .O(\vga_select_6<0>/GROM )
  );
  X_BUF \vga_select_6<0>/XUSED  (
    .I(\vga_select_6<0>/FROM ),
    .O(vga_select_6[0])
  );
  X_BUF \vga_select_6<0>/YUSED  (
    .I(\vga_select_6<0>/GROM ),
    .O(CHOICE3906)
  );
  defparam \DLX_EXinst__n0006<14>119 .INIT = 16'hAE00;
  X_LUT4 \DLX_EXinst__n0006<14>119  (
    .ADR0(DLX_EXinst__n0046),
    .ADR1(DLX_EXinst__n0047),
    .ADR2(DLX_IDinst_reg_out_A[14]),
    .ADR3(DLX_IDinst_reg_out_B[14]),
    .O(\CHOICE4256/FROM )
  );
  defparam \DLX_EXinst__n0006<20>158 .INIT = 16'hA0E0;
  X_LUT4 \DLX_EXinst__n0006<20>158  (
    .ADR0(DLX_EXinst__n0046),
    .ADR1(DLX_EXinst__n0047),
    .ADR2(DLX_IDinst_reg_out_B[20]),
    .ADR3(DLX_IDinst_reg_out_A[20]),
    .O(\CHOICE4256/GROM )
  );
  X_BUF \CHOICE4256/XUSED  (
    .I(\CHOICE4256/FROM ),
    .O(CHOICE4256)
  );
  X_BUF \CHOICE4256/YUSED  (
    .I(\CHOICE4256/GROM ),
    .O(CHOICE4904)
  );
  defparam \DLX_EXinst__n0006<12>175 .INIT = 16'hECA0;
  X_LUT4 \DLX_EXinst__n0006<12>175  (
    .ADR0(DLX_EXinst_N66383),
    .ADR1(DLX_EXinst_N66535),
    .ADR2(\DLX_EXinst_Mshift__n0026_Sh[60] ),
    .ADR3(\DLX_EXinst_Mshift__n0025_Sh[44] ),
    .O(\CHOICE3903/FROM )
  );
  defparam \DLX_EXinst__n0006<12>184 .INIT = 16'hD5C0;
  X_LUT4 \DLX_EXinst__n0006<12>184  (
    .ADR0(N110935),
    .ADR1(N95810),
    .ADR2(DLX_EXinst_N66177),
    .ADR3(CHOICE3903),
    .O(\CHOICE3903/GROM )
  );
  X_BUF \CHOICE3903/XUSED  (
    .I(\CHOICE3903/FROM ),
    .O(CHOICE3903)
  );
  X_BUF \CHOICE3903/YUSED  (
    .I(\CHOICE3903/GROM ),
    .O(CHOICE3905)
  );
  defparam \DLX_EXinst__n0006<20>176 .INIT = 16'hF8F8;
  X_LUT4 \DLX_EXinst__n0006<20>176  (
    .ADR0(DLX_EXinst__n0045),
    .ADR1(DLX_IDinst_reg_out_B[20]),
    .ADR2(DLX_EXinst_N64448),
    .ADR3(VCC),
    .O(\CHOICE4913/FROM )
  );
  defparam \DLX_EXinst__n0006<20>185 .INIT = 16'hF040;
  X_LUT4 \DLX_EXinst__n0006<20>185  (
    .ADR0(DLX_IDinst_reg_out_B[20]),
    .ADR1(DLX_EXinst__n0047),
    .ADR2(DLX_IDinst_reg_out_A[20]),
    .ADR3(CHOICE4913),
    .O(\CHOICE4913/GROM )
  );
  X_BUF \CHOICE4913/XUSED  (
    .I(\CHOICE4913/FROM ),
    .O(CHOICE4913)
  );
  X_BUF \CHOICE4913/YUSED  (
    .I(\CHOICE4913/GROM ),
    .O(CHOICE4915)
  );
  defparam \Mshift__n0000_Sh<37>1 .INIT = 16'h00A0;
  X_LUT4 \Mshift__n0000_Sh<37>1  (
    .ADR0(DLX_EXinst_ALU_result[12]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_ALU_result[14]),
    .ADR3(DLX_EXinst_ALU_result[13]),
    .O(\vga_select_6<5>/FROM )
  );
  defparam \DLX_EXinst__n0006<13>200 .INIT = 16'hFEEE;
  X_LUT4 \DLX_EXinst__n0006<13>200  (
    .ADR0(CHOICE4329),
    .ADR1(CHOICE4339),
    .ADR2(N101725),
    .ADR3(DLX_EXinst_ALU_result[13]),
    .O(\vga_select_6<5>/GROM )
  );
  X_BUF \vga_select_6<5>/XUSED  (
    .I(\vga_select_6<5>/FROM ),
    .O(vga_select_6[5])
  );
  X_BUF \vga_select_6<5>/YUSED  (
    .I(\vga_select_6<5>/GROM ),
    .O(CHOICE4340)
  );
  defparam \DLX_EXinst_Mshift__n0027_Sh<4>28 .INIT = 16'hFFAA;
  X_LUT4 \DLX_EXinst_Mshift__n0027_Sh<4>28  (
    .ADR0(CHOICE1012),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(CHOICE1006),
    .O(\DLX_EXinst_Mshift__n0027_Sh<4>/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0027_Sh<44>11 .INIT = 16'h8A80;
  X_LUT4 \DLX_EXinst_Mshift__n0027_Sh<44>11  (
    .ADR0(DLX_IDinst_IR_function_field_3_1),
    .ADR1(\DLX_EXinst_Mshift__n0027_Sh[0] ),
    .ADR2(DLX_IDinst_IR_function_field_2_1),
    .ADR3(\DLX_EXinst_Mshift__n0027_Sh[4] ),
    .O(\DLX_EXinst_Mshift__n0027_Sh<4>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0027_Sh<4>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0027_Sh<4>/FROM ),
    .O(\DLX_EXinst_Mshift__n0027_Sh[4] )
  );
  X_BUF \DLX_EXinst_Mshift__n0027_Sh<4>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0027_Sh<4>/GROM ),
    .O(CHOICE1042)
  );
  defparam DLX_IDlc_md_mda5_a1.INIT = 16'h2222;
  X_LUT4 DLX_IDlc_md_mda5_a1 (
    .ADR0(DLX_IDlc_md_wint4),
    .ADR1(DLX_IDlc_pd_wint1),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IDlc_md_wint5/FROM )
  );
  defparam DLX_IDlc_md_mda39_a1.INIT = 16'h00CC;
  X_LUT4 DLX_IDlc_md_mda39_a1 (
    .ADR0(VCC),
    .ADR1(DLX_IDlc_md_wint38),
    .ADR2(VCC),
    .ADR3(DLX_IDlc_pd_wint1),
    .O(\DLX_IDlc_md_wint5/GROM )
  );
  X_BUF \DLX_IDlc_md_wint5/XUSED  (
    .I(\DLX_IDlc_md_wint5/FROM ),
    .O(DLX_IDlc_md_wint5)
  );
  X_BUF \DLX_IDlc_md_wint5/YUSED  (
    .I(\DLX_IDlc_md_wint5/GROM ),
    .O(DLX_IDlc_md_wint39)
  );
  defparam \DLX_EXinst__n0006<23>312_SW0 .INIT = 16'h00FE;
  X_LUT4 \DLX_EXinst__n0006<23>312_SW0  (
    .ADR0(CHOICE4043),
    .ADR1(CHOICE4057),
    .ADR2(CHOICE4032),
    .ADR3(DLX_EXinst__n0030),
    .O(\DLX_EXinst_ALU_result<23>/FROM )
  );
  defparam \DLX_EXinst__n0006<23>312 .INIT = 16'hCCC8;
  X_LUT4 \DLX_EXinst__n0006<23>312  (
    .ADR0(CHOICE4091),
    .ADR1(DLX_EXinst__n0149),
    .ADR2(N100490),
    .ADR3(N126538),
    .O(N114054)
  );
  X_BUF \DLX_EXinst_ALU_result<23>/XUSED  (
    .I(\DLX_EXinst_ALU_result<23>/FROM ),
    .O(N126538)
  );
  defparam \DLX_EXinst__n0006<19>288 .INIT = 16'hEAC0;
  X_LUT4 \DLX_EXinst__n0006<19>288  (
    .ADR0(N101725),
    .ADR1(DLX_EXinst__n0016[19]),
    .ADR2(DLX_EXinst__n0114),
    .ADR3(DLX_EXinst_ALU_result[19]),
    .O(\CHOICE4999/FROM )
  );
  defparam \DLX_EXinst__n0006<21>213 .INIT = 16'hF888;
  X_LUT4 \DLX_EXinst__n0006<21>213  (
    .ADR0(DLX_EXinst__n0114),
    .ADR1(DLX_EXinst__n0016[21]),
    .ADR2(DLX_EXinst_ALU_result[21]),
    .ADR3(N101725),
    .O(\CHOICE4999/GROM )
  );
  X_BUF \CHOICE4999/XUSED  (
    .I(\CHOICE4999/FROM ),
    .O(CHOICE4999)
  );
  X_BUF \CHOICE4999/YUSED  (
    .I(\CHOICE4999/GROM ),
    .O(CHOICE4211)
  );
  defparam \DLX_IFinst__n0001<15>_SW0 .INIT = 16'h1B1B;
  X_LUT4 \DLX_IFinst__n0001<15>_SW0  (
    .ADR0(DLX_IFinst__n0000),
    .ADR1(DLX_IFinst__n0015[15]),
    .ADR2(DLX_IFinst_PC[15]),
    .ADR3(VCC),
    .O(\DLX_IFinst_NPC<15>/FROM )
  );
  defparam \DLX_IFinst__n0001<15> .INIT = 16'hA0AF;
  X_LUT4 \DLX_IFinst__n0001<15>  (
    .ADR0(DLX_IDinst_branch_address[15]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(N92347),
    .O(\DLX_IFinst_NPC<15>/GROM )
  );
  X_BUF \DLX_IFinst_NPC<15>/XUSED  (
    .I(\DLX_IFinst_NPC<15>/FROM ),
    .O(N92347)
  );
  X_BUF \DLX_IFinst_NPC<15>/YUSED  (
    .I(\DLX_IFinst_NPC<15>/GROM ),
    .O(DLX_IFinst__n0001[15])
  );
  defparam \DLX_IFinst__n0001<31>_SW0 .INIT = 16'h11DD;
  X_LUT4 \DLX_IFinst__n0001<31>_SW0  (
    .ADR0(DLX_IFinst__n0015[31]),
    .ADR1(DLX_IFinst__n0000),
    .ADR2(VCC),
    .ADR3(DLX_IFinst_PC[31]),
    .O(\DLX_IFinst_NPC<31>/FROM )
  );
  defparam \DLX_IFinst__n0001<31> .INIT = 16'hA0AF;
  X_LUT4 \DLX_IFinst__n0001<31>  (
    .ADR0(DLX_IDinst_branch_address[31]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(N91515),
    .O(DLX_IFinst__n0001[31])
  );
  X_BUF \DLX_IFinst_NPC<31>/XUSED  (
    .I(\DLX_IFinst_NPC<31>/FROM ),
    .O(N91515)
  );
  defparam \DLX_IFinst__n0001<23>_SW0 .INIT = 16'h05F5;
  X_LUT4 \DLX_IFinst__n0001<23>_SW0  (
    .ADR0(DLX_IFinst__n0015[23]),
    .ADR1(VCC),
    .ADR2(DLX_IFinst__n0000),
    .ADR3(DLX_IFinst_PC[23]),
    .O(\DLX_IFinst_NPC<23>/FROM )
  );
  defparam \DLX_IFinst__n0001<23> .INIT = 16'hA0AF;
  X_LUT4 \DLX_IFinst__n0001<23>  (
    .ADR0(DLX_IDinst_branch_address[23]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(N91931),
    .O(DLX_IFinst__n0001[23])
  );
  X_BUF \DLX_IFinst_NPC<23>/XUSED  (
    .I(\DLX_IFinst_NPC<23>/FROM ),
    .O(N91931)
  );
  defparam \DLX_EXinst__n0006<21>231 .INIT = 16'h88C8;
  X_LUT4 \DLX_EXinst__n0006<21>231  (
    .ADR0(CHOICE4217),
    .ADR1(DLX_IDinst_reg_out_A[21]),
    .ADR2(DLX_EXinst__n0047),
    .ADR3(DLX_IDinst_reg_out_B[21]),
    .O(\CHOICE4219/FROM )
  );
  defparam \DLX_EXinst__n0006<21>236 .INIT = 16'hFF50;
  X_LUT4 \DLX_EXinst__n0006<21>236  (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(VCC),
    .ADR2(N108433),
    .ADR3(CHOICE4219),
    .O(\CHOICE4219/GROM )
  );
  X_BUF \CHOICE4219/XUSED  (
    .I(\CHOICE4219/FROM ),
    .O(CHOICE4219)
  );
  X_BUF \CHOICE4219/YUSED  (
    .I(\CHOICE4219/GROM ),
    .O(CHOICE4220)
  );
  defparam \DLX_EXinst_Mshift__n0027_Sh<5>26 .INIT = 16'h0C0A;
  X_LUT4 \DLX_EXinst_Mshift__n0027_Sh<5>26  (
    .ADR0(DLX_IDinst_reg_out_A[5]),
    .ADR1(DLX_IDinst_reg_out_A[3]),
    .ADR2(DLX_IDinst_IR_function_field_0_1),
    .ADR3(DLX_IDinst_IR_function_field_1_1),
    .O(\CHOICE1024/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0027_Sh<5>28 .INIT = 16'hFFCC;
  X_LUT4 \DLX_EXinst_Mshift__n0027_Sh<5>28  (
    .ADR0(VCC),
    .ADR1(CHOICE1018),
    .ADR2(VCC),
    .ADR3(CHOICE1024),
    .O(\CHOICE1024/GROM )
  );
  X_BUF \CHOICE1024/XUSED  (
    .I(\CHOICE1024/FROM ),
    .O(CHOICE1024)
  );
  X_BUF \CHOICE1024/YUSED  (
    .I(\CHOICE1024/GROM ),
    .O(\DLX_EXinst_Mshift__n0027_Sh[5] )
  );
  defparam \DLX_EXinst__n0006<26>158 .INIT = 16'hC0C8;
  X_LUT4 \DLX_EXinst__n0006<26>158  (
    .ADR0(DLX_EXinst__n0047),
    .ADR1(DLX_IDinst_reg_out_B[26]),
    .ADR2(DLX_EXinst__n0046),
    .ADR3(DLX_IDinst_reg_out_A[26]),
    .O(\CHOICE4708/FROM )
  );
  defparam \DLX_EXinst__n0006<13>119 .INIT = 16'hC4C0;
  X_LUT4 \DLX_EXinst__n0006<13>119  (
    .ADR0(DLX_IDinst_reg_out_A[13]),
    .ADR1(DLX_IDinst_reg_out_B[13]),
    .ADR2(DLX_EXinst__n0046),
    .ADR3(DLX_EXinst__n0047),
    .O(\CHOICE4708/GROM )
  );
  X_BUF \CHOICE4708/XUSED  (
    .I(\CHOICE4708/FROM ),
    .O(CHOICE4708)
  );
  X_BUF \CHOICE4708/YUSED  (
    .I(\CHOICE4708/GROM ),
    .O(CHOICE4316)
  );
  defparam DLX_EXlc_master_ctrlEX__n00021.INIT = 16'h50DC;
  X_LUT4 DLX_EXlc_master_ctrlEX__n00021 (
    .ADR0(DLX_EXlc_md_outp2),
    .ADR1(DLX_EXlc_master_ctrlEX_nro),
    .ADR2(CHOICE12),
    .ADR3(DLX_EXlc_slave_ctrlEX_l),
    .O(\DLX_EXlc_master_ctrlEX_nro/FROM )
  );
  defparam DLX_EXlc_master_ctrlEX__n0001_SW19.INIT = 16'hBBFF;
  X_LUT4 DLX_EXlc_master_ctrlEX__n0001_SW19 (
    .ADR0(reset_IBUF),
    .ADR1(DLX_ackin_EX),
    .ADR2(VCC),
    .ADR3(DLX_EXlc_master_ctrlEX_nro),
    .O(\DLX_EXlc_master_ctrlEX_nro/GROM )
  );
  X_BUF \DLX_EXlc_master_ctrlEX_nro/XUSED  (
    .I(\DLX_EXlc_master_ctrlEX_nro/FROM ),
    .O(DLX_EXlc_master_ctrlEX_nro)
  );
  X_BUF \DLX_EXlc_master_ctrlEX_nro/YUSED  (
    .I(\DLX_EXlc_master_ctrlEX_nro/GROM ),
    .O(CHOICE12)
  );
  defparam \DLX_EXinst__n0006<13>226 .INIT = 16'hCCC8;
  X_LUT4 \DLX_EXinst__n0006<13>226  (
    .ADR0(CHOICE4321),
    .ADR1(DLX_EXinst__n0030),
    .ADR2(CHOICE4340),
    .ADR3(CHOICE4316),
    .O(\CHOICE4342/FROM )
  );
  defparam \DLX_EXinst__n0006<13>238 .INIT = 16'hFFC0;
  X_LUT4 \DLX_EXinst__n0006<13>238  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N63836),
    .ADR2(DLX_EXinst__n0016[13]),
    .ADR3(CHOICE4342),
    .O(\CHOICE4342/GROM )
  );
  X_BUF \CHOICE4342/XUSED  (
    .I(\CHOICE4342/FROM ),
    .O(CHOICE4342)
  );
  X_BUF \CHOICE4342/YUSED  (
    .I(\CHOICE4342/GROM ),
    .O(CHOICE4343)
  );
  defparam \DLX_EXinst__n0006<21>171 .INIT = 16'h3202;
  X_LUT4 \DLX_EXinst__n0006<21>171  (
    .ADR0(DLX_EXinst_N64094),
    .ADR1(DLX_IDinst_reg_out_B[4]),
    .ADR2(DLX_IDinst_reg_out_B[2]),
    .ADR3(DLX_EXinst_N63910),
    .O(\CHOICE4205/FROM )
  );
  defparam \DLX_EXinst__n0006<21>177 .INIT = 16'hFF08;
  X_LUT4 \DLX_EXinst__n0006<21>177  (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(DLX_EXinst_N62906),
    .ADR2(DLX_IDinst_reg_out_B[3]),
    .ADR3(CHOICE4205),
    .O(\CHOICE4205/GROM )
  );
  X_BUF \CHOICE4205/XUSED  (
    .I(\CHOICE4205/FROM ),
    .O(CHOICE4205)
  );
  X_BUF \CHOICE4205/YUSED  (
    .I(\CHOICE4205/GROM ),
    .O(CHOICE4206)
  );
  defparam \DLX_EXinst__n0006<13>180 .INIT = 16'hFF08;
  X_LUT4 \DLX_EXinst__n0006<13>180  (
    .ADR0(DLX_EXinst_N66383),
    .ADR1(\DLX_EXinst_Mshift__n0026_Sh[29] ),
    .ADR2(DLX_EXinst_N62740),
    .ADR3(CHOICE4336),
    .O(\CHOICE4337/FROM )
  );
  defparam \DLX_EXinst__n0006<13>192 .INIT = 16'hB3A0;
  X_LUT4 \DLX_EXinst__n0006<13>192  (
    .ADR0(DLX_EXinst_N65090),
    .ADR1(N110935),
    .ADR2(DLX_EXinst_N66177),
    .ADR3(CHOICE4337),
    .O(\CHOICE4337/GROM )
  );
  X_BUF \CHOICE4337/XUSED  (
    .I(\CHOICE4337/FROM ),
    .O(CHOICE4337)
  );
  X_BUF \CHOICE4337/YUSED  (
    .I(\CHOICE4337/GROM ),
    .O(CHOICE4339)
  );
  defparam \DLX_EXinst__n0006<13>149 .INIT = 16'hFCF0;
  X_LUT4 \DLX_EXinst__n0006<13>149  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst__n0045),
    .ADR2(DLX_EXinst_N64448),
    .ADR3(DLX_IDinst_reg_out_B[13]),
    .O(\CHOICE4327/FROM )
  );
  defparam \DLX_EXinst__n0006<13>158 .INIT = 16'hAA20;
  X_LUT4 \DLX_EXinst__n0006<13>158  (
    .ADR0(DLX_IDinst_reg_out_A[13]),
    .ADR1(DLX_IDinst_reg_out_B[13]),
    .ADR2(DLX_EXinst__n0047),
    .ADR3(CHOICE4327),
    .O(\CHOICE4327/GROM )
  );
  X_BUF \CHOICE4327/XUSED  (
    .I(\CHOICE4327/FROM ),
    .O(CHOICE4327)
  );
  X_BUF \CHOICE4327/YUSED  (
    .I(\CHOICE4327/GROM ),
    .O(CHOICE4329)
  );
  defparam \Mshift__n0000_Sh<36>1 .INIT = 16'h0300;
  X_LUT4 \Mshift__n0000_Sh<36>1  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_ALU_result[13]),
    .ADR2(DLX_EXinst_ALU_result[12]),
    .ADR3(DLX_EXinst_ALU_result[14]),
    .O(\vga_select_6<4>/FROM )
  );
  defparam \DLX_EXinst__n0006<14>200 .INIT = 16'hFEEE;
  X_LUT4 \DLX_EXinst__n0006<14>200  (
    .ADR0(CHOICE4269),
    .ADR1(CHOICE4279),
    .ADR2(DLX_EXinst_ALU_result[14]),
    .ADR3(N101725),
    .O(\vga_select_6<4>/GROM )
  );
  X_BUF \vga_select_6<4>/XUSED  (
    .I(\vga_select_6<4>/FROM ),
    .O(vga_select_6[4])
  );
  X_BUF \vga_select_6<4>/YUSED  (
    .I(\vga_select_6<4>/GROM ),
    .O(CHOICE4280)
  );
  defparam \DLX_IFinst__n0001<3>_SW0 .INIT = 16'h11DD;
  X_LUT4 \DLX_IFinst__n0001<3>_SW0  (
    .ADR0(DLX_IFinst__n0015[3]),
    .ADR1(DLX_IFinst__n0000),
    .ADR2(VCC),
    .ADR3(DLX_IFinst_PC[3]),
    .O(\DLX_IFinst_NPC<3>/FROM )
  );
  defparam \DLX_IFinst__n0001<3> .INIT = 16'hC0CF;
  X_LUT4 \DLX_IFinst__n0001<3>  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_branch_address[3]),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(N92971),
    .O(\DLX_IFinst_NPC<3>/GROM )
  );
  X_BUF \DLX_IFinst_NPC<3>/XUSED  (
    .I(\DLX_IFinst_NPC<3>/FROM ),
    .O(N92971)
  );
  X_BUF \DLX_IFinst_NPC<3>/YUSED  (
    .I(\DLX_IFinst_NPC<3>/GROM ),
    .O(DLX_IFinst__n0001[3])
  );
  defparam \DLX_EXinst__n0006<22>236 .INIT = 16'hAAFA;
  X_LUT4 \DLX_EXinst__n0006<22>236  (
    .ADR0(CHOICE4153),
    .ADR1(VCC),
    .ADR2(N108909),
    .ADR3(DLX_IDinst_reg_out_B[4]),
    .O(\CHOICE4154/FROM )
  );
  defparam \DLX_EXinst__n0006<27>240_SW0 .INIT = 16'hA0EC;
  X_LUT4 \DLX_EXinst__n0006<27>240_SW0  (
    .ADR0(N101725),
    .ADR1(N105035),
    .ADR2(DLX_EXinst_ALU_result[27]),
    .ADR3(DLX_IDinst_reg_out_B[4]),
    .O(\CHOICE4154/GROM )
  );
  X_BUF \CHOICE4154/XUSED  (
    .I(\CHOICE4154/FROM ),
    .O(CHOICE4154)
  );
  X_BUF \CHOICE4154/YUSED  (
    .I(\CHOICE4154/GROM ),
    .O(N126411)
  );
  defparam \DLX_EXinst__n0006<22>222 .INIT = 16'hFFC0;
  X_LUT4 \DLX_EXinst__n0006<22>222  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst__n0045),
    .ADR2(DLX_IDinst_reg_out_B[22]),
    .ADR3(DLX_EXinst_N64448),
    .O(\CHOICE4151/FROM )
  );
  defparam \DLX_EXinst__n0006<22>231 .INIT = 16'hF020;
  X_LUT4 \DLX_EXinst__n0006<22>231  (
    .ADR0(DLX_EXinst__n0047),
    .ADR1(DLX_IDinst_reg_out_B[22]),
    .ADR2(DLX_IDinst_reg_out_A[22]),
    .ADR3(CHOICE4151),
    .O(\CHOICE4151/GROM )
  );
  X_BUF \CHOICE4151/XUSED  (
    .I(\CHOICE4151/FROM ),
    .O(CHOICE4151)
  );
  X_BUF \CHOICE4151/YUSED  (
    .I(\CHOICE4151/GROM ),
    .O(CHOICE4153)
  );
  defparam \DLX_IDinst_slot_num_FFd3-In24 .INIT = 16'hFFA8;
  X_LUT4 \DLX_IDinst_slot_num_FFd3-In24  (
    .ADR0(DLX_IDinst_delay_slot),
    .ADR1(DLX_IDinst_slot_num_FFd3),
    .ADR2(DLX_IDinst_slot_num_FFd1),
    .ADR3(CHOICE2508),
    .O(\DLX_IDinst_slot_num_FFd3/FROM )
  );
  defparam \DLX_IDinst_slot_num_FFd3-In33 .INIT = 16'hFF8A;
  X_LUT4 \DLX_IDinst_slot_num_FFd3-In33  (
    .ADR0(DLX_IDinst_N70077),
    .ADR1(DLX_IDinst_intr_slot),
    .ADR2(DLX_EXinst__n0149),
    .ADR3(CHOICE2509),
    .O(\DLX_IDinst_slot_num_FFd3-In )
  );
  X_BUF \DLX_IDinst_slot_num_FFd3/XUSED  (
    .I(\DLX_IDinst_slot_num_FFd3/FROM ),
    .O(CHOICE2509)
  );
  defparam \DLX_EXinst__n0006<0>277_SW0_SW0 .INIT = 16'hAFA0;
  X_LUT4 \DLX_EXinst__n0006<0>277_SW0_SW0  (
    .ADR0(DLX_EXinst_Mcompar__n0059_inst_cy_196),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_IR_function_field[0]),
    .ADR3(DLX_EXinst_Mcompar__n0057_inst_cy_164),
    .O(\N127567/FROM )
  );
  defparam \DLX_EXinst__n0006<0>277_SW0 .INIT = 16'h18DB;
  X_LUT4 \DLX_EXinst__n0006<0>277_SW0  (
    .ADR0(DLX_IDinst_IR_function_field[0]),
    .ADR1(DLX_IDinst_reg_out_A[31]),
    .ADR2(DLX_IDinst_reg_out_B[31]),
    .ADR3(N127567),
    .O(\N127567/GROM )
  );
  X_BUF \N127567/XUSED  (
    .I(\N127567/FROM ),
    .O(N127567)
  );
  X_BUF \N127567/YUSED  (
    .I(\N127567/GROM ),
    .O(N126107)
  );
  defparam \DLX_EXinst__n0006<14>226 .INIT = 16'hFE00;
  X_LUT4 \DLX_EXinst__n0006<14>226  (
    .ADR0(CHOICE4280),
    .ADR1(CHOICE4261),
    .ADR2(CHOICE4256),
    .ADR3(DLX_EXinst__n0030),
    .O(\CHOICE4282/FROM )
  );
  defparam \DLX_EXinst__n0006<14>238 .INIT = 16'hFF88;
  X_LUT4 \DLX_EXinst__n0006<14>238  (
    .ADR0(DLX_EXinst_N63836),
    .ADR1(DLX_EXinst__n0016[14]),
    .ADR2(VCC),
    .ADR3(CHOICE4282),
    .O(\CHOICE4282/GROM )
  );
  X_BUF \CHOICE4282/XUSED  (
    .I(\CHOICE4282/FROM ),
    .O(CHOICE4282)
  );
  X_BUF \CHOICE4282/YUSED  (
    .I(\CHOICE4282/GROM ),
    .O(CHOICE4283)
  );
  defparam \DLX_EXinst__n0006<22>171 .INIT = 16'h00E2;
  X_LUT4 \DLX_EXinst__n0006<22>171  (
    .ADR0(DLX_EXinst_N64099),
    .ADR1(DLX_IDinst_reg_out_B[2]),
    .ADR2(DLX_EXinst_N63915),
    .ADR3(DLX_IDinst_reg_out_B[4]),
    .O(\CHOICE4139/FROM )
  );
  defparam \DLX_EXinst__n0006<22>177 .INIT = 16'hFF20;
  X_LUT4 \DLX_EXinst__n0006<22>177  (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(DLX_IDinst_reg_out_B[3]),
    .ADR2(DLX_EXinst_N62911),
    .ADR3(CHOICE4139),
    .O(\CHOICE4139/GROM )
  );
  X_BUF \CHOICE4139/XUSED  (
    .I(\CHOICE4139/FROM ),
    .O(CHOICE4139)
  );
  X_BUF \CHOICE4139/YUSED  (
    .I(\CHOICE4139/GROM ),
    .O(CHOICE4140)
  );
  defparam \DLX_EXinst__n0006<14>180 .INIT = 16'hF2F0;
  X_LUT4 \DLX_EXinst__n0006<14>180  (
    .ADR0(DLX_EXinst_N66383),
    .ADR1(DLX_EXinst_N62740),
    .ADR2(CHOICE4276),
    .ADR3(\DLX_EXinst_Mshift__n0026_Sh[30] ),
    .O(\CHOICE4277/FROM )
  );
  defparam \DLX_EXinst__n0006<14>192 .INIT = 16'hB3A0;
  X_LUT4 \DLX_EXinst__n0006<14>192  (
    .ADR0(DLX_EXinst_N66177),
    .ADR1(N110935),
    .ADR2(N95120),
    .ADR3(CHOICE4277),
    .O(\CHOICE4277/GROM )
  );
  X_BUF \CHOICE4277/XUSED  (
    .I(\CHOICE4277/FROM ),
    .O(CHOICE4277)
  );
  X_BUF \CHOICE4277/YUSED  (
    .I(\CHOICE4277/GROM ),
    .O(CHOICE4279)
  );
  defparam \DLX_EXinst__n0006<14>149 .INIT = 16'hFF88;
  X_LUT4 \DLX_EXinst__n0006<14>149  (
    .ADR0(DLX_IDinst_reg_out_B[14]),
    .ADR1(DLX_EXinst__n0045),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N64448),
    .O(\CHOICE4267/FROM )
  );
  defparam \DLX_EXinst__n0006<14>158 .INIT = 16'hAA08;
  X_LUT4 \DLX_EXinst__n0006<14>158  (
    .ADR0(DLX_IDinst_reg_out_A[14]),
    .ADR1(DLX_EXinst__n0047),
    .ADR2(DLX_IDinst_reg_out_B[14]),
    .ADR3(CHOICE4267),
    .O(\CHOICE4267/GROM )
  );
  X_BUF \CHOICE4267/XUSED  (
    .I(\CHOICE4267/FROM ),
    .O(CHOICE4267)
  );
  X_BUF \CHOICE4267/YUSED  (
    .I(\CHOICE4267/GROM ),
    .O(CHOICE4269)
  );
  defparam \DLX_EXinst__n0006<28>346 .INIT = 16'hF888;
  X_LUT4 \DLX_EXinst__n0006<28>346  (
    .ADR0(DLX_EXinst_N63996),
    .ADR1(DLX_IDinst_reg_out_A[26]),
    .ADR2(DLX_IDinst_reg_out_A[27]),
    .ADR3(DLX_EXinst_N64181),
    .O(\CHOICE5247/FROM )
  );
  defparam \DLX_EXinst__n0006<30>350 .INIT = 16'hF888;
  X_LUT4 \DLX_EXinst__n0006<30>350  (
    .ADR0(DLX_EXinst_N63996),
    .ADR1(DLX_IDinst_reg_out_A[28]),
    .ADR2(DLX_EXinst_N64181),
    .ADR3(DLX_IDinst_reg_out_A[29]),
    .O(\CHOICE5247/GROM )
  );
  X_BUF \CHOICE5247/XUSED  (
    .I(\CHOICE5247/FROM ),
    .O(CHOICE5247)
  );
  X_BUF \CHOICE5247/YUSED  (
    .I(\CHOICE5247/GROM ),
    .O(CHOICE5324)
  );
  defparam \DLX_EXinst__n0006<15>103 .INIT = 16'hFAFE;
  X_LUT4 \DLX_EXinst__n0006<15>103  (
    .ADR0(CHOICE4830),
    .ADR1(CHOICE4806),
    .ADR2(CHOICE4811),
    .ADR3(N109130),
    .O(\CHOICE4831/GROM )
  );
  X_BUF \CHOICE4831/YUSED  (
    .I(\CHOICE4831/GROM ),
    .O(CHOICE4831)
  );
  defparam \DLX_EXinst__n0006<31>224 .INIT = 16'h3222;
  X_LUT4 \DLX_EXinst__n0006<31>224  (
    .ADR0(N126500),
    .ADR1(N110935),
    .ADR2(\DLX_EXinst_Mshift__n0023_Sh[127] ),
    .ADR3(DLX_EXinst_N66392),
    .O(\CHOICE5784/FROM )
  );
  defparam \DLX_EXinst__n0006<30>257 .INIT = 16'hF3F2;
  X_LUT4 \DLX_EXinst__n0006<30>257  (
    .ADR0(CHOICE5297),
    .ADR1(N110935),
    .ADR2(CHOICE5306),
    .ADR3(CHOICE5300),
    .O(\CHOICE5784/GROM )
  );
  X_BUF \CHOICE5784/XUSED  (
    .I(\CHOICE5784/FROM ),
    .O(CHOICE5784)
  );
  X_BUF \CHOICE5784/YUSED  (
    .I(\CHOICE5784/GROM ),
    .O(CHOICE5307)
  );
  defparam \DLX_EXinst__n0006<30>284 .INIT = 16'h8C88;
  X_LUT4 \DLX_EXinst__n0006<30>284  (
    .ADR0(CHOICE5313),
    .ADR1(DLX_IDinst_reg_out_A[30]),
    .ADR2(DLX_IDinst_reg_out_B[30]),
    .ADR3(DLX_EXinst__n0047),
    .O(\CHOICE5315/FROM )
  );
  defparam \DLX_EXinst__n0006<30>288 .INIT = 16'hFFC0;
  X_LUT4 \DLX_EXinst__n0006<30>288  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_ALU_result[30]),
    .ADR2(N101725),
    .ADR3(CHOICE5315),
    .O(\CHOICE5315/GROM )
  );
  X_BUF \CHOICE5315/XUSED  (
    .I(\CHOICE5315/FROM ),
    .O(CHOICE5315)
  );
  X_BUF \CHOICE5315/YUSED  (
    .I(\CHOICE5315/GROM ),
    .O(CHOICE5316)
  );
  defparam \DLX_EXinst__n0006<15>204 .INIT = 16'hECA0;
  X_LUT4 \DLX_EXinst__n0006<15>204  (
    .ADR0(DLX_EXinst_N66535),
    .ADR1(DLX_EXinst_N66383),
    .ADR2(\DLX_EXinst_Mshift__n0025_Sh[47] ),
    .ADR3(\DLX_EXinst_Mshift__n0023_Sh[127] ),
    .O(\CHOICE4860/FROM )
  );
  defparam \DLX_EXinst__n0006<15>210 .INIT = 16'hB3A0;
  X_LUT4 \DLX_EXinst__n0006<15>210  (
    .ADR0(DLX_IDinst_reg_out_A[15]),
    .ADR1(N110935),
    .ADR2(N126257),
    .ADR3(CHOICE4860),
    .O(\CHOICE4860/GROM )
  );
  X_BUF \CHOICE4860/XUSED  (
    .I(\CHOICE4860/FROM ),
    .O(CHOICE4860)
  );
  X_BUF \CHOICE4860/YUSED  (
    .I(\CHOICE4860/GROM ),
    .O(CHOICE4862)
  );
  defparam \DLX_EXinst__n0006<16>323 .INIT = 16'hFFEC;
  X_LUT4 \DLX_EXinst__n0006<16>323  (
    .ADR0(DLX_EXinst_ALU_result[16]),
    .ADR1(CHOICE5147),
    .ADR2(N101725),
    .ADR3(CHOICE5168),
    .O(\CHOICE5169/FROM )
  );
  defparam \DLX_EXinst__n0006<23>213 .INIT = 16'hECA0;
  X_LUT4 \DLX_EXinst__n0006<23>213  (
    .ADR0(DLX_EXinst__n0016[23]),
    .ADR1(N101725),
    .ADR2(DLX_EXinst__n0114),
    .ADR3(DLX_EXinst_ALU_result[23]),
    .O(\CHOICE5169/GROM )
  );
  X_BUF \CHOICE5169/XUSED  (
    .I(\CHOICE5169/FROM ),
    .O(CHOICE5169)
  );
  X_BUF \CHOICE5169/YUSED  (
    .I(\CHOICE5169/GROM ),
    .O(CHOICE4079)
  );
  defparam \DLX_EXinst__n0006<23>222 .INIT = 16'hFCCC;
  X_LUT4 \DLX_EXinst__n0006<23>222  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N64448),
    .ADR2(DLX_EXinst__n0045),
    .ADR3(DLX_IDinst_reg_out_B[23]),
    .O(\CHOICE4085/FROM )
  );
  defparam \DLX_EXinst__n0006<23>231 .INIT = 16'hAA20;
  X_LUT4 \DLX_EXinst__n0006<23>231  (
    .ADR0(DLX_IDinst_reg_out_A[23]),
    .ADR1(DLX_IDinst_reg_out_B[23]),
    .ADR2(DLX_EXinst__n0047),
    .ADR3(CHOICE4085),
    .O(\CHOICE4085/GROM )
  );
  X_BUF \CHOICE4085/XUSED  (
    .I(\CHOICE4085/FROM ),
    .O(CHOICE4085)
  );
  X_BUF \CHOICE4085/YUSED  (
    .I(\CHOICE4085/GROM ),
    .O(CHOICE4087)
  );
  defparam \DLX_IFinst__n0001<24>_SW0 .INIT = 16'h05F5;
  X_LUT4 \DLX_IFinst__n0001<24>_SW0  (
    .ADR0(DLX_IFinst__n0015[24]),
    .ADR1(VCC),
    .ADR2(DLX_IFinst__n0000),
    .ADR3(DLX_IFinst_PC[24]),
    .O(\DLX_IFinst_NPC<24>/FROM )
  );
  defparam \DLX_IFinst__n0001<24> .INIT = 16'h88BB;
  X_LUT4 \DLX_IFinst__n0001<24>  (
    .ADR0(DLX_IDinst_branch_address[24]),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(VCC),
    .ADR3(N91879),
    .O(DLX_IFinst__n0001[24])
  );
  X_BUF \DLX_IFinst_NPC<24>/XUSED  (
    .I(\DLX_IFinst_NPC<24>/FROM ),
    .O(N91879)
  );
  defparam \DLX_IFinst__n0001<16>_SW0 .INIT = 16'h0C3F;
  X_LUT4 \DLX_IFinst__n0001<16>_SW0  (
    .ADR0(VCC),
    .ADR1(DLX_IFinst__n0000),
    .ADR2(DLX_IFinst_PC[16]),
    .ADR3(DLX_IFinst__n0015[16]),
    .O(\DLX_IFinst_NPC<16>/FROM )
  );
  defparam \DLX_IFinst__n0001<16> .INIT = 16'hA0AF;
  X_LUT4 \DLX_IFinst__n0001<16>  (
    .ADR0(DLX_IDinst_branch_address[16]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(N92243),
    .O(DLX_IFinst__n0001[16])
  );
  X_BUF \DLX_IFinst_NPC<16>/XUSED  (
    .I(\DLX_IFinst_NPC<16>/FROM ),
    .O(N92243)
  );
  defparam \DLX_EXinst__n0006<30>367 .INIT = 16'hFEFC;
  X_LUT4 \DLX_EXinst__n0006<30>367  (
    .ADR0(DLX_EXinst_N63836),
    .ADR1(N126514),
    .ADR2(N100490),
    .ADR3(DLX_EXinst__n0016[30]),
    .O(\DLX_EXinst_ALU_result<30>/FROM )
  );
  defparam \DLX_EXinst__n0006<30>378 .INIT = 16'h1100;
  X_LUT4 \DLX_EXinst__n0006<30>378  (
    .ADR0(DLX_IDinst_counter[0]),
    .ADR1(DLX_IDinst_counter[1]),
    .ADR2(VCC),
    .ADR3(CHOICE5326),
    .O(N121549)
  );
  X_BUF \DLX_EXinst_ALU_result<30>/XUSED  (
    .I(\DLX_EXinst_ALU_result<30>/FROM ),
    .O(CHOICE5326)
  );
  defparam \DLX_EXinst__n0006<0>449_SW0_SW0 .INIT = 16'hBB88;
  X_LUT4 \DLX_EXinst__n0006<0>449_SW0_SW0  (
    .ADR0(DLX_EXinst_Mcompar__n0091_inst_cy_196),
    .ADR1(DLX_IDinst_IR_opcode_field[0]),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_Mcompar__n0089_inst_cy_164),
    .O(\N127563/FROM )
  );
  defparam \DLX_EXinst__n0006<0>449_SW0 .INIT = 16'h18DB;
  X_LUT4 \DLX_EXinst__n0006<0>449_SW0  (
    .ADR0(DLX_IDinst_IR_opcode_field[0]),
    .ADR1(DLX_IDinst_reg_out_A[31]),
    .ADR2(\DLX_IDinst_Imm[31] ),
    .ADR3(N127563),
    .O(\N127563/GROM )
  );
  X_BUF \N127563/XUSED  (
    .I(\N127563/FROM ),
    .O(N127563)
  );
  X_BUF \N127563/YUSED  (
    .I(\N127563/GROM ),
    .O(N126092)
  );
  defparam \DLX_EXinst__n0006<24>141 .INIT = 16'hC4C0;
  X_LUT4 \DLX_EXinst__n0006<24>141  (
    .ADR0(DLX_IDinst_reg_out_A[24]),
    .ADR1(DLX_IDinst_reg_out_B[24]),
    .ADR2(DLX_EXinst__n0046),
    .ADR3(DLX_EXinst__n0047),
    .O(\CHOICE3766/FROM )
  );
  defparam \DLX_EXinst__n0006<15>137 .INIT = 16'hCE00;
  X_LUT4 \DLX_EXinst__n0006<15>137  (
    .ADR0(DLX_EXinst__n0047),
    .ADR1(DLX_EXinst__n0046),
    .ADR2(DLX_IDinst_reg_out_A[15]),
    .ADR3(DLX_IDinst_reg_out_B[15]),
    .O(\CHOICE3766/GROM )
  );
  X_BUF \CHOICE3766/XUSED  (
    .I(\CHOICE3766/FROM ),
    .O(CHOICE3766)
  );
  X_BUF \CHOICE3766/YUSED  (
    .I(\CHOICE3766/GROM ),
    .O(CHOICE4837)
  );
  defparam \DLX_EXinst__n0006<15>250 .INIT = 16'hFE00;
  X_LUT4 \DLX_EXinst__n0006<15>250  (
    .ADR0(CHOICE4863),
    .ADR1(CHOICE4837),
    .ADR2(CHOICE4842),
    .ADR3(DLX_EXinst__n0030),
    .O(\CHOICE4865/FROM )
  );
  defparam \DLX_EXinst__n0006<15>262 .INIT = 16'hFF88;
  X_LUT4 \DLX_EXinst__n0006<15>262  (
    .ADR0(DLX_EXinst_N63836),
    .ADR1(DLX_EXinst__n0016[15]),
    .ADR2(VCC),
    .ADR3(CHOICE4865),
    .O(\CHOICE4865/GROM )
  );
  X_BUF \CHOICE4865/XUSED  (
    .I(\CHOICE4865/FROM ),
    .O(CHOICE4865)
  );
  X_BUF \CHOICE4865/YUSED  (
    .I(\CHOICE4865/GROM ),
    .O(CHOICE4866)
  );
  defparam \DLX_EXinst__n0006<23>171 .INIT = 16'h00D8;
  X_LUT4 \DLX_EXinst__n0006<23>171  (
    .ADR0(DLX_IDinst_reg_out_B[2]),
    .ADR1(DLX_EXinst_N63920),
    .ADR2(DLX_EXinst_N64104),
    .ADR3(DLX_IDinst_reg_out_B[4]),
    .O(\CHOICE4073/FROM )
  );
  defparam \DLX_EXinst__n0006<23>177 .INIT = 16'hFF40;
  X_LUT4 \DLX_EXinst__n0006<23>177  (
    .ADR0(DLX_IDinst_reg_out_B[3]),
    .ADR1(DLX_EXinst_N62916),
    .ADR2(DLX_IDinst_reg_out_B[4]),
    .ADR3(CHOICE4073),
    .O(\CHOICE4073/GROM )
  );
  X_BUF \CHOICE4073/XUSED  (
    .I(\CHOICE4073/FROM ),
    .O(CHOICE4073)
  );
  X_BUF \CHOICE4073/YUSED  (
    .I(\CHOICE4073/GROM ),
    .O(CHOICE4074)
  );
  defparam \DLX_EXinst__n0006<18>149 .INIT = 16'hFEFA;
  X_LUT4 \DLX_EXinst__n0006<18>149  (
    .ADR0(CHOICE5421),
    .ADR1(DLX_EXinst__n0128),
    .ADR2(N126398),
    .ADR3(DLX_EXinst__n0016[18]),
    .O(\CHOICE5440/FROM )
  );
  defparam \DLX_EXinst__n0006<31>500 .INIT = 16'hF888;
  X_LUT4 \DLX_EXinst__n0006<31>500  (
    .ADR0(DLX_EXinst__n0016[31]),
    .ADR1(DLX_EXinst__n0128),
    .ADR2(DLX_EXinst__n0077),
    .ADR3(\DLX_IDinst_Imm[15] ),
    .O(\CHOICE5440/GROM )
  );
  X_BUF \CHOICE5440/XUSED  (
    .I(\CHOICE5440/FROM ),
    .O(CHOICE5440)
  );
  X_BUF \CHOICE5440/YUSED  (
    .I(\CHOICE5440/GROM ),
    .O(CHOICE5828)
  );
  defparam \DLX_EXinst__n0006<31>238 .INIT = 16'hFAF0;
  X_LUT4 \DLX_EXinst__n0006<31>238  (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(VCC),
    .ADR2(CHOICE5784),
    .ADR3(CHOICE5754),
    .O(\CHOICE5785/FROM )
  );
  defparam \DLX_EXinst__n0006<31>277_SW0 .INIT = 16'hFF80;
  X_LUT4 \DLX_EXinst__n0006<31>277_SW0  (
    .ADR0(DLX_EXinst_N66078),
    .ADR1(\DLX_EXinst_Mshift__n0023_Sh[127] ),
    .ADR2(DLX_IDinst_reg_out_B[5]),
    .ADR3(CHOICE5785),
    .O(\CHOICE5785/GROM )
  );
  X_BUF \CHOICE5785/XUSED  (
    .I(\CHOICE5785/FROM ),
    .O(CHOICE5785)
  );
  X_BUF \CHOICE5785/YUSED  (
    .I(\CHOICE5785/GROM ),
    .O(N126495)
  );
  defparam \DLX_IFinst__n0001<4>_SW0 .INIT = 16'h0C3F;
  X_LUT4 \DLX_IFinst__n0001<4>_SW0  (
    .ADR0(VCC),
    .ADR1(DLX_IFinst__n0000),
    .ADR2(DLX_IFinst_PC[4]),
    .ADR3(DLX_IFinst__n0015[4]),
    .O(\DLX_IFinst_NPC<4>/FROM )
  );
  defparam \DLX_IFinst__n0001<4> .INIT = 16'h88DD;
  X_LUT4 \DLX_IFinst__n0001<4>  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(DLX_IDinst_branch_address[4]),
    .ADR2(VCC),
    .ADR3(N92919),
    .O(\DLX_IFinst_NPC<4>/GROM )
  );
  X_BUF \DLX_IFinst_NPC<4>/XUSED  (
    .I(\DLX_IFinst_NPC<4>/FROM ),
    .O(N92919)
  );
  X_BUF \DLX_IFinst_NPC<4>/YUSED  (
    .I(\DLX_IFinst_NPC<4>/GROM ),
    .O(DLX_IFinst__n0001[4])
  );
  defparam \DLX_EXinst__n0006<27>306_SW0 .INIT = 16'h0F0E;
  X_LUT4 \DLX_EXinst__n0006<27>306_SW0  (
    .ADR0(CHOICE4610),
    .ADR1(CHOICE4636),
    .ADR2(DLX_EXinst__n0030),
    .ADR3(CHOICE4611),
    .O(\DLX_EXinst_ALU_result<27>/FROM )
  );
  defparam \DLX_EXinst__n0006<27>306 .INIT = 16'hAAA8;
  X_LUT4 \DLX_EXinst__n0006<27>306  (
    .ADR0(DLX_EXinst__n0149),
    .ADR1(CHOICE4668),
    .ADR2(N100490),
    .ADR3(N126403),
    .O(N117545)
  );
  X_BUF \DLX_EXinst_ALU_result<27>/XUSED  (
    .I(\DLX_EXinst_ALU_result<27>/FROM ),
    .O(N126403)
  );
  defparam \DLX_EXinst__n0006<15>290 .INIT = 16'hAE00;
  X_LUT4 \DLX_EXinst__n0006<15>290  (
    .ADR0(CHOICE4866),
    .ADR1(CHOICE4831),
    .ADR2(DLX_EXinst__n0030),
    .ADR3(DLX_EXinst__n0149),
    .O(\DLX_EXinst_ALU_result<15>/FROM )
  );
  defparam \DLX_EXinst__n0006<15>300 .INIT = 16'hFFAA;
  X_LUT4 \DLX_EXinst__n0006<15>300  (
    .ADR0(DLX_EXinst_N63689),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(CHOICE4868),
    .O(N118737)
  );
  X_BUF \DLX_EXinst_ALU_result<15>/XUSED  (
    .I(\DLX_EXinst_ALU_result<15>/FROM ),
    .O(CHOICE4868)
  );
  X_INV \DLX_MEMinst_reg_dst_out<1>/CKINV  (
    .I(DLX_MEMlc_master_ctrlMEM_l),
    .O(\DLX_MEMinst_reg_dst_out<1>/CKMUXNOT )
  );
  defparam \DLX_EXinst__n0006<31>444 .INIT = 16'h0808;
  X_LUT4 \DLX_EXinst__n0006<31>444  (
    .ADR0(DLX_EXinst__n0082),
    .ADR1(\DLX_EXinst_Mshift__n0024_Sh[127] ),
    .ADR2(DLX_IDinst_IR_function_field[4]),
    .ADR3(VCC),
    .O(\CHOICE5818/FROM )
  );
  defparam \DLX_EXinst__n0006<31>584_SW0 .INIT = 16'hF3F2;
  X_LUT4 \DLX_EXinst__n0006<31>584_SW0  (
    .ADR0(CHOICE5815),
    .ADR1(N109130),
    .ADR2(CHOICE5842),
    .ADR3(CHOICE5818),
    .O(\CHOICE5818/GROM )
  );
  X_BUF \CHOICE5818/XUSED  (
    .I(\CHOICE5818/FROM ),
    .O(CHOICE5818)
  );
  X_BUF \CHOICE5818/YUSED  (
    .I(\CHOICE5818/GROM ),
    .O(N126446)
  );
  defparam \DLX_EXinst__n0006<31>277 .INIT = 16'hF0E0;
  X_LUT4 \DLX_EXinst__n0006<31>277  (
    .ADR0(CHOICE5746),
    .ADR1(CHOICE5740),
    .ADR2(DLX_EXinst__n0030),
    .ADR3(N126495),
    .O(\DLX_EXinst_ALU_result<31>/FROM )
  );
  defparam \DLX_EXinst__n0006<31>610 .INIT = 16'h0504;
  X_LUT4 \DLX_EXinst__n0006<31>610  (
    .ADR0(DLX_IDinst_counter[1]),
    .ADR1(CHOICE5845),
    .ADR2(DLX_IDinst_counter[0]),
    .ADR3(CHOICE5788),
    .O(N124731)
  );
  X_BUF \DLX_EXinst_ALU_result<31>/XUSED  (
    .I(\DLX_EXinst_ALU_result<31>/FROM ),
    .O(CHOICE5788)
  );
  defparam \DLX_EXinst__n0006<16>125 .INIT = 16'hECA0;
  X_LUT4 \DLX_EXinst__n0006<16>125  (
    .ADR0(DLX_EXinst_N66202),
    .ADR1(DLX_IDinst_reg_out_A[16]),
    .ADR2(CHOICE5126),
    .ADR3(N126362),
    .O(\CHOICE5128/GROM )
  );
  X_BUF \CHOICE5128/YUSED  (
    .I(\CHOICE5128/GROM ),
    .O(CHOICE5128)
  );
  X_INV \DLX_MEMinst_reg_dst_out<3>/CKINV  (
    .I(DLX_MEMlc_master_ctrlMEM_l),
    .O(\DLX_MEMinst_reg_dst_out<3>/CKMUXNOT )
  );
  defparam \DLX_EXinst__n0006<24>223 .INIT = 16'hFFEA;
  X_LUT4 \DLX_EXinst__n0006<24>223  (
    .ADR0(CHOICE3785),
    .ADR1(DLX_EXinst__n0114),
    .ADR2(DLX_EXinst__n0016[24]),
    .ADR3(N126546),
    .O(\CHOICE3789/FROM )
  );
  defparam \DLX_EXinst__n0006<24>251 .INIT = 16'hF0E0;
  X_LUT4 \DLX_EXinst__n0006<24>251  (
    .ADR0(CHOICE3766),
    .ADR1(CHOICE3775),
    .ADR2(DLX_EXinst__n0030),
    .ADR3(CHOICE3789),
    .O(\CHOICE3789/GROM )
  );
  X_BUF \CHOICE3789/XUSED  (
    .I(\CHOICE3789/FROM ),
    .O(CHOICE3789)
  );
  X_BUF \CHOICE3789/YUSED  (
    .I(\CHOICE3789/GROM ),
    .O(CHOICE3791)
  );
  defparam \DLX_EXinst__n0006<16>207 .INIT = 16'hFFC0;
  X_LUT4 \DLX_EXinst__n0006<16>207  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_B[16]),
    .ADR2(DLX_EXinst__n0045),
    .ADR3(DLX_EXinst_N64448),
    .O(\CHOICE5145/FROM )
  );
  defparam \DLX_EXinst__n0006<16>216 .INIT = 16'hAA20;
  X_LUT4 \DLX_EXinst__n0006<16>216  (
    .ADR0(DLX_IDinst_reg_out_A[16]),
    .ADR1(DLX_IDinst_reg_out_B[16]),
    .ADR2(DLX_EXinst__n0047),
    .ADR3(CHOICE5145),
    .O(\CHOICE5145/GROM )
  );
  X_BUF \CHOICE5145/XUSED  (
    .I(\CHOICE5145/FROM ),
    .O(CHOICE5145)
  );
  X_BUF \CHOICE5145/YUSED  (
    .I(\CHOICE5145/GROM ),
    .O(CHOICE5147)
  );
  X_INV \DLX_MEMinst_reg_dst_out<4>/CKINV  (
    .I(DLX_MEMlc_master_ctrlMEM_l),
    .O(\DLX_MEMinst_reg_dst_out<4>/CKMUXNOT )
  );
  defparam DLX_MEMlc_slave_ctrlMEM__n00021.INIT = 16'h0031;
  X_LUT4 DLX_MEMlc_slave_ctrlMEM__n00021 (
    .ADR0(DLX_ackin_ID),
    .ADR1(DLX_MEMlc_slave_ctrlMEM_l),
    .ADR2(DLX_reqout_MEM),
    .ADR3(reset_IBUF_1),
    .O(\DLX_reqout_MEM/FROM )
  );
  defparam DLX_cg1_c1.INIT = 16'hFCC0;
  X_LUT4 DLX_cg1_c1 (
    .ADR0(VCC),
    .ADR1(DLX_reqout_IF),
    .ADR2(DLX_reqin_ID),
    .ADR3(DLX_reqout_MEM),
    .O(\DLX_reqout_MEM/GROM )
  );
  X_BUF \DLX_reqout_MEM/XUSED  (
    .I(\DLX_reqout_MEM/FROM ),
    .O(DLX_reqout_MEM)
  );
  X_BUF \DLX_reqout_MEM/YUSED  (
    .I(\DLX_reqout_MEM/GROM ),
    .O(DLX_reqin_ID)
  );
  defparam DLX_MEMlc_md_mda10_a1.INIT = 16'h5500;
  X_LUT4 DLX_MEMlc_md_mda10_a1 (
    .ADR0(DLX_MEMlc_pd_wint1),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_MEMlc_md_wint9),
    .O(\DLX_MEMlc_md_wint10/FROM )
  );
  defparam DLX_MEMlc_md_mda11_a1.INIT = 16'h3300;
  X_LUT4 DLX_MEMlc_md_mda11_a1 (
    .ADR0(VCC),
    .ADR1(DLX_MEMlc_pd_wint1),
    .ADR2(VCC),
    .ADR3(DLX_MEMlc_md_wint10),
    .O(\DLX_MEMlc_md_wint10/GROM )
  );
  X_BUF \DLX_MEMlc_md_wint10/XUSED  (
    .I(\DLX_MEMlc_md_wint10/FROM ),
    .O(DLX_MEMlc_md_wint10)
  );
  X_BUF \DLX_MEMlc_md_wint10/YUSED  (
    .I(\DLX_MEMlc_md_wint10/GROM ),
    .O(DLX_MEMlc_md_wint11)
  );
  defparam \DLX_EXinst__n0006<31>481 .INIT = 16'h4000;
  X_LUT4 \DLX_EXinst__n0006<31>481  (
    .ADR0(DLX_IDinst_IR_function_field[4]),
    .ADR1(\DLX_EXinst_Mshift__n0024_Sh[127] ),
    .ADR2(\DLX_IDinst_Imm[5] ),
    .ADR3(N110065),
    .O(\CHOICE5824/FROM )
  );
  defparam \DLX_EXinst__n0006<31>584 .INIT = 16'h5554;
  X_LUT4 \DLX_EXinst__n0006<31>584  (
    .ADR0(DLX_EXinst__n0030),
    .ADR1(CHOICE5828),
    .ADR2(N126446),
    .ADR3(CHOICE5824),
    .O(\CHOICE5824/GROM )
  );
  X_BUF \CHOICE5824/XUSED  (
    .I(\CHOICE5824/FROM ),
    .O(CHOICE5824)
  );
  X_BUF \CHOICE5824/YUSED  (
    .I(\CHOICE5824/GROM ),
    .O(CHOICE5845)
  );
  defparam \DLX_EXinst__n0006<16>306 .INIT = 16'hEAC0;
  X_LUT4 \DLX_EXinst__n0006<16>306  (
    .ADR0(DLX_EXinst_N66226),
    .ADR1(N126263),
    .ADR2(DLX_IDinst_reg_out_B[16]),
    .ADR3(CHOICE5166),
    .O(\CHOICE5168/GROM )
  );
  X_BUF \CHOICE5168/YUSED  (
    .I(\CHOICE5168/GROM ),
    .O(CHOICE5168)
  );
  defparam vga_top_vga1__n000972_SW0.INIT = 16'hFEFA;
  X_LUT4 vga_top_vga1__n000972_SW0 (
    .ADR0(CHOICE3427),
    .ADR1(vga_top_vga1_N73394),
    .ADR2(vga_top_vga1_helpme),
    .ADR3(CHOICE3425),
    .O(\N126344/FROM )
  );
  defparam vga_top_vga1__n000972.INIT = 16'hFFC8;
  X_LUT4 vga_top_vga1__n000972 (
    .ADR0(CHOICE3412),
    .ADR1(vga_top_vga1_vcounter[9]),
    .ADR2(CHOICE3416),
    .ADR3(N126344),
    .O(\N126344/GROM )
  );
  X_BUF \N126344/XUSED  (
    .I(\N126344/FROM ),
    .O(N126344)
  );
  X_BUF \N126344/YUSED  (
    .I(\N126344/GROM ),
    .O(N110183)
  );
  defparam \DLX_EXinst__n0006<24>155 .INIT = 16'h5044;
  X_LUT4 \DLX_EXinst__n0006<24>155  (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(N97161),
    .ADR2(DLX_EXinst_N63925),
    .ADR3(DLX_IDinst_reg_out_B[2]),
    .O(\CHOICE3773/FROM )
  );
  defparam \DLX_EXinst__n0006<24>168 .INIT = 16'hCC80;
  X_LUT4 \DLX_EXinst__n0006<24>168  (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(DLX_EXinst_N66226),
    .ADR2(\DLX_EXinst_Mshift__n0025_Sh[40] ),
    .ADR3(CHOICE3773),
    .O(\CHOICE3773/GROM )
  );
  X_BUF \CHOICE3773/XUSED  (
    .I(\CHOICE3773/FROM ),
    .O(CHOICE3773)
  );
  X_BUF \CHOICE3773/YUSED  (
    .I(\CHOICE3773/GROM ),
    .O(CHOICE3775)
  );
  defparam \DLX_EXinst__n0006<17>109 .INIT = 16'hCE0A;
  X_LUT4 \DLX_EXinst__n0006<17>109  (
    .ADR0(N126631),
    .ADR1(N110065),
    .ADR2(N109130),
    .ADR3(N101338),
    .O(\CHOICE5603/FROM )
  );
  defparam \DLX_EXinst__n0006<17>149_SW0 .INIT = 16'h8F88;
  X_LUT4 \DLX_EXinst__n0006<17>149_SW0  (
    .ADR0(DLX_IDinst_IR_function_field[1]),
    .ADR1(DLX_EXinst__n0077),
    .ADR2(DLX_IDinst_IR_function_field[4]),
    .ADR3(CHOICE5603),
    .O(\CHOICE5603/GROM )
  );
  X_BUF \CHOICE5603/XUSED  (
    .I(\CHOICE5603/FROM ),
    .O(CHOICE5603)
  );
  X_BUF \CHOICE5603/YUSED  (
    .I(\CHOICE5603/GROM ),
    .O(N126627)
  );
  defparam \DLX_IDinst__n0086<7>27_SW0 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst__n0086<7>27_SW0  (
    .ADR0(DLX_IDinst_N70328),
    .ADR1(DLX_IDinst_regA_eff[7]),
    .ADR2(DLX_IDinst__n0128[7]),
    .ADR3(DLX_IDinst_N70072),
    .O(\N127423/GROM )
  );
  X_BUF \N127423/YUSED  (
    .I(\N127423/GROM ),
    .O(N127423)
  );
  defparam \DLX_IFinst__n0001<17>_SW0 .INIT = 16'h3355;
  X_LUT4 \DLX_IFinst__n0001<17>_SW0  (
    .ADR0(DLX_IFinst__n0015[17]),
    .ADR1(DLX_IFinst_PC[17]),
    .ADR2(VCC),
    .ADR3(DLX_IFinst__n0000),
    .O(\DLX_IFinst_NPC<17>/FROM )
  );
  defparam \DLX_IFinst__n0001<17> .INIT = 16'hA0F5;
  X_LUT4 \DLX_IFinst__n0001<17>  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_branch_address[17]),
    .ADR3(N92295),
    .O(DLX_IFinst__n0001[17])
  );
  X_BUF \DLX_IFinst_NPC<17>/XUSED  (
    .I(\DLX_IFinst_NPC<17>/FROM ),
    .O(N92295)
  );
  defparam DLX_IDinst__n0004_SW0.INIT = 16'hFFF0;
  X_LUT4 DLX_IDinst__n0004_SW0 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_regB_index[1]),
    .ADR3(DLX_IDinst_regB_index[0]),
    .O(\N90373/FROM )
  );
  defparam DLX_IDinst__n0004_1183.INIT = 16'h0001;
  X_LUT4 DLX_IDinst__n0004_1183 (
    .ADR0(DLX_IDinst_regB_index[3]),
    .ADR1(DLX_IDinst_regB_index[2]),
    .ADR2(DLX_IDinst_regB_index[4]),
    .ADR3(N90373),
    .O(\N90373/GROM )
  );
  X_BUF \N90373/XUSED  (
    .I(\N90373/FROM ),
    .O(N90373)
  );
  X_BUF \N90373/YUSED  (
    .I(\N90373/GROM ),
    .O(DLX_IDinst__n0004)
  );
  defparam \DLX_EXinst__n0006<17>302 .INIT = 16'hDC50;
  X_LUT4 \DLX_EXinst__n0006<17>302  (
    .ADR0(N110935),
    .ADR1(N101425),
    .ADR2(N126610),
    .ADR3(N111221),
    .O(\CHOICE5642/FROM )
  );
  defparam \DLX_EXinst__n0006<17>343_SW0 .INIT = 16'hB3A0;
  X_LUT4 \DLX_EXinst__n0006<17>343_SW0  (
    .ADR0(N101725),
    .ADR1(DLX_IDinst_reg_out_B[4]),
    .ADR2(DLX_EXinst_ALU_result[17]),
    .ADR3(CHOICE5642),
    .O(\CHOICE5642/GROM )
  );
  X_BUF \CHOICE5642/XUSED  (
    .I(\CHOICE5642/FROM ),
    .O(CHOICE5642)
  );
  X_BUF \CHOICE5642/YUSED  (
    .I(\CHOICE5642/GROM ),
    .O(N126606)
  );
  defparam \DLX_IFinst__n0001<25>_SW0 .INIT = 16'h2277;
  X_LUT4 \DLX_IFinst__n0001<25>_SW0  (
    .ADR0(DLX_IFinst__n0000),
    .ADR1(DLX_IFinst_PC[25]),
    .ADR2(VCC),
    .ADR3(DLX_IFinst__n0015[25]),
    .O(\DLX_IFinst_NPC<25>/FROM )
  );
  defparam \DLX_IFinst__n0001<25> .INIT = 16'h88BB;
  X_LUT4 \DLX_IFinst__n0001<25>  (
    .ADR0(DLX_IDinst_branch_address[25]),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(VCC),
    .ADR3(N91827),
    .O(DLX_IFinst__n0001[25])
  );
  X_BUF \DLX_IFinst_NPC<25>/XUSED  (
    .I(\DLX_IFinst_NPC<25>/FROM ),
    .O(N91827)
  );
  defparam \DLX_EXinst__n0006<24>199 .INIT = 16'hFFC0;
  X_LUT4 \DLX_EXinst__n0006<24>199  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst__n0045),
    .ADR2(DLX_IDinst_reg_out_B[24]),
    .ADR3(DLX_EXinst_N64448),
    .O(\CHOICE3783/FROM )
  );
  defparam \DLX_EXinst__n0006<24>208 .INIT = 16'hF020;
  X_LUT4 \DLX_EXinst__n0006<24>208  (
    .ADR0(DLX_EXinst__n0047),
    .ADR1(DLX_IDinst_reg_out_B[24]),
    .ADR2(DLX_IDinst_reg_out_A[24]),
    .ADR3(CHOICE3783),
    .O(\CHOICE3783/GROM )
  );
  X_BUF \CHOICE3783/XUSED  (
    .I(\CHOICE3783/FROM ),
    .O(CHOICE3783)
  );
  X_BUF \CHOICE3783/YUSED  (
    .I(\CHOICE3783/GROM ),
    .O(CHOICE3785)
  );
  defparam \DLX_EXinst__n0006<16>375 .INIT = 16'hFF32;
  X_LUT4 \DLX_EXinst__n0006<16>375  (
    .ADR0(CHOICE5100),
    .ADR1(DLX_EXinst__n0030),
    .ADR2(CHOICE5129),
    .ADR3(CHOICE5172),
    .O(\DLX_EXinst_ALU_result<16>/FROM )
  );
  defparam \DLX_EXinst__n0006<16>401 .INIT = 16'hF1F0;
  X_LUT4 \DLX_EXinst__n0006<16>401  (
    .ADR0(DLX_IDinst_counter[0]),
    .ADR1(DLX_IDinst_counter[1]),
    .ADR2(DLX_EXinst_N63689),
    .ADR3(CHOICE5173),
    .O(N120627)
  );
  X_BUF \DLX_EXinst_ALU_result<16>/XUSED  (
    .I(\DLX_EXinst_ALU_result<16>/FROM ),
    .O(CHOICE5173)
  );
  defparam \DLX_EXinst__n0006<25>216 .INIT = 16'hFCCC;
  X_LUT4 \DLX_EXinst__n0006<25>216  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N64448),
    .ADR2(DLX_EXinst__n0045),
    .ADR3(DLX_IDinst_reg_out_B[25]),
    .O(\CHOICE4790/FROM )
  );
  defparam \DLX_EXinst__n0006<25>225 .INIT = 16'hF200;
  X_LUT4 \DLX_EXinst__n0006<25>225  (
    .ADR0(DLX_EXinst__n0047),
    .ADR1(DLX_IDinst_reg_out_B[25]),
    .ADR2(CHOICE4790),
    .ADR3(DLX_IDinst_reg_out_A[25]),
    .O(\CHOICE4790/GROM )
  );
  X_BUF \CHOICE4790/XUSED  (
    .I(\CHOICE4790/FROM ),
    .O(CHOICE4790)
  );
  X_BUF \CHOICE4790/YUSED  (
    .I(\CHOICE4790/GROM ),
    .O(CHOICE4792)
  );
  defparam \Mshift__n0000_Sh<33>1 .INIT = 16'h1100;
  X_LUT4 \Mshift__n0000_Sh<33>1  (
    .ADR0(DLX_EXinst_ALU_result[13]),
    .ADR1(DLX_EXinst_ALU_result[14]),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_ALU_result[12]),
    .O(\vga_select_6<1>/GROM )
  );
  X_BUF \vga_select_6<1>/YUSED  (
    .I(\vga_select_6<1>/GROM ),
    .O(vga_select_6[1])
  );
  defparam \DLX_EXinst__n0006<17>227 .INIT = 16'hEECC;
  X_LUT4 \DLX_EXinst__n0006<17>227  (
    .ADR0(DLX_EXinst__n0045),
    .ADR1(DLX_EXinst_N64448),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[17]),
    .O(\CHOICE5625/FROM )
  );
  defparam \DLX_EXinst__n0006<17>236 .INIT = 16'hAA20;
  X_LUT4 \DLX_EXinst__n0006<17>236  (
    .ADR0(DLX_IDinst_reg_out_A[17]),
    .ADR1(DLX_IDinst_reg_out_B[17]),
    .ADR2(DLX_EXinst__n0047),
    .ADR3(CHOICE5625),
    .O(\CHOICE5625/GROM )
  );
  X_BUF \CHOICE5625/XUSED  (
    .I(\CHOICE5625/FROM ),
    .O(CHOICE5625)
  );
  X_BUF \CHOICE5625/YUSED  (
    .I(\CHOICE5625/GROM ),
    .O(CHOICE5627)
  );
  defparam \DLX_EXinst__n0006<26>110 .INIT = 16'hFEEE;
  X_LUT4 \DLX_EXinst__n0006<26>110  (
    .ADR0(CHOICE4686),
    .ADR1(N126375),
    .ADR2(DLX_EXinst__n0128),
    .ADR3(DLX_EXinst__n0016[26]),
    .O(\CHOICE4701/FROM )
  );
  defparam \DLX_EXinst__n0006<17>149 .INIT = 16'hFFEC;
  X_LUT4 \DLX_EXinst__n0006<17>149  (
    .ADR0(DLX_EXinst__n0128),
    .ADR1(N126627),
    .ADR2(DLX_EXinst__n0016[17]),
    .ADR3(CHOICE5587),
    .O(\CHOICE4701/GROM )
  );
  X_BUF \CHOICE4701/XUSED  (
    .I(\CHOICE4701/FROM ),
    .O(CHOICE4701)
  );
  X_BUF \CHOICE4701/YUSED  (
    .I(\CHOICE4701/GROM ),
    .O(CHOICE5606)
  );
  defparam \Mshift__n0000_Sh<34>1 .INIT = 16'h1010;
  X_LUT4 \Mshift__n0000_Sh<34>1  (
    .ADR0(DLX_EXinst_ALU_result[14]),
    .ADR1(DLX_EXinst_ALU_result[12]),
    .ADR2(DLX_EXinst_ALU_result[13]),
    .ADR3(VCC),
    .O(\vga_select_6<2>/FROM )
  );
  defparam Ker5730284_SW0.INIT = 16'hAA00;
  X_LUT4 Ker5730284_SW0 (
    .ADR0(vram_out_cpu[1]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_select_6[2]),
    .O(\vga_select_6<2>/GROM )
  );
  X_BUF \vga_select_6<2>/XUSED  (
    .I(\vga_select_6<2>/FROM ),
    .O(vga_select_6[2])
  );
  X_BUF \vga_select_6<2>/YUSED  (
    .I(\vga_select_6<2>/GROM ),
    .O(N126029)
  );
  defparam \DLX_EXinst__n0006<25>158 .INIT = 16'hAA08;
  X_LUT4 \DLX_EXinst__n0006<25>158  (
    .ADR0(DLX_IDinst_reg_out_B[25]),
    .ADR1(DLX_EXinst__n0047),
    .ADR2(DLX_IDinst_reg_out_A[25]),
    .ADR3(DLX_EXinst__n0046),
    .O(\CHOICE4773/GROM )
  );
  X_BUF \CHOICE4773/YUSED  (
    .I(\CHOICE4773/GROM ),
    .O(CHOICE4773)
  );
  defparam \DLX_EXinst__n0006<17>343 .INIT = 16'hFFF8;
  X_LUT4 \DLX_EXinst__n0006<17>343  (
    .ADR0(DLX_EXinst__n0114),
    .ADR1(DLX_EXinst__n0016[17]),
    .ADR2(N126606),
    .ADR3(CHOICE5627),
    .O(\CHOICE5646/FROM )
  );
  defparam \DLX_EXinst__n0006<17>371 .INIT = 16'hF0E0;
  X_LUT4 \DLX_EXinst__n0006<17>371  (
    .ADR0(CHOICE5617),
    .ADR1(CHOICE5613),
    .ADR2(DLX_EXinst__n0030),
    .ADR3(CHOICE5646),
    .O(\CHOICE5646/GROM )
  );
  X_BUF \CHOICE5646/XUSED  (
    .I(\CHOICE5646/FROM ),
    .O(CHOICE5646)
  );
  X_BUF \CHOICE5646/YUSED  (
    .I(\CHOICE5646/GROM ),
    .O(CHOICE5648)
  );
  defparam \DLX_IFinst__n0001<5>_SW0 .INIT = 16'h4747;
  X_LUT4 \DLX_IFinst__n0001<5>_SW0  (
    .ADR0(DLX_IFinst_PC[5]),
    .ADR1(DLX_IFinst__n0000),
    .ADR2(DLX_IFinst__n0015[5]),
    .ADR3(VCC),
    .O(\DLX_IFinst_NPC<5>/FROM )
  );
  defparam \DLX_IFinst__n0001<5> .INIT = 16'hAF05;
  X_LUT4 \DLX_IFinst__n0001<5>  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(VCC),
    .ADR2(N92815),
    .ADR3(DLX_IDinst_branch_address[5]),
    .O(\DLX_IFinst_NPC<5>/GROM )
  );
  X_BUF \DLX_IFinst_NPC<5>/XUSED  (
    .I(\DLX_IFinst_NPC<5>/FROM ),
    .O(N92815)
  );
  X_BUF \DLX_IFinst_NPC<5>/YUSED  (
    .I(\DLX_IFinst_NPC<5>/GROM ),
    .O(DLX_IFinst__n0001[5])
  );
  defparam \DLX_EXinst__n0006<25>185 .INIT = 16'hC8C0;
  X_LUT4 \DLX_EXinst__n0006<25>185  (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(DLX_EXinst_N66226),
    .ADR2(CHOICE4780),
    .ADR3(\DLX_EXinst_Mshift__n0025_Sh[41] ),
    .O(\CHOICE4782/FROM )
  );
  defparam \DLX_EXinst__n0006<25>268 .INIT = 16'hCCC8;
  X_LUT4 \DLX_EXinst__n0006<25>268  (
    .ADR0(CHOICE4773),
    .ADR1(DLX_EXinst__n0030),
    .ADR2(CHOICE4796),
    .ADR3(CHOICE4782),
    .O(\CHOICE4782/GROM )
  );
  X_BUF \CHOICE4782/XUSED  (
    .I(\CHOICE4782/FROM ),
    .O(CHOICE4782)
  );
  X_BUF \CHOICE4782/YUSED  (
    .I(\CHOICE4782/GROM ),
    .O(CHOICE4798)
  );
  defparam \Mshift__n0000_Sh<35>1 .INIT = 16'h0C00;
  X_LUT4 \Mshift__n0000_Sh<35>1  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_ALU_result[13]),
    .ADR2(DLX_EXinst_ALU_result[14]),
    .ADR3(DLX_EXinst_ALU_result[12]),
    .O(\vga_select_6<3>/FROM )
  );
  defparam Ker57310_SW0.INIT = 16'hFFFA;
  X_LUT4 Ker57310_SW0 (
    .ADR0(vga_select_6[5]),
    .ADR1(VCC),
    .ADR2(vga_select_6[4]),
    .ADR3(vga_select_6[3]),
    .O(\vga_select_6<3>/GROM )
  );
  X_BUF \vga_select_6<3>/XUSED  (
    .I(\vga_select_6<3>/FROM ),
    .O(vga_select_6[3])
  );
  X_BUF \vga_select_6<3>/YUSED  (
    .I(\vga_select_6<3>/GROM ),
    .O(N95202)
  );
  defparam Ker5730215.INIT = 16'hFD0D;
  X_LUT4 Ker5730215 (
    .ADR0(vga_select_6[5]),
    .ADR1(vram_out_cpu[4]),
    .ADR2(vga_select_6[4]),
    .ADR3(vram_out_cpu[3]),
    .O(\CHOICE2937/FROM )
  );
  defparam Ker5730239.INIT = 16'h0D08;
  X_LUT4 Ker5730239 (
    .ADR0(vga_select_6[3]),
    .ADR1(vram_out_cpu[2]),
    .ADR2(vga_select_6[2]),
    .ADR3(CHOICE2937),
    .O(\CHOICE2937/GROM )
  );
  X_BUF \CHOICE2937/XUSED  (
    .I(\CHOICE2937/FROM ),
    .O(CHOICE2937)
  );
  X_BUF \CHOICE2937/YUSED  (
    .I(\CHOICE2937/GROM ),
    .O(CHOICE2941)
  );
  defparam \DLX_EXinst__n0006<18>109 .INIT = 16'hAE0C;
  X_LUT4 \DLX_EXinst__n0006<18>109  (
    .ADR0(N110065),
    .ADR1(N126407),
    .ADR2(N109130),
    .ADR3(N101095),
    .O(\CHOICE5437/FROM )
  );
  defparam \DLX_EXinst__n0006<18>149_SW0 .INIT = 16'hD5C0;
  X_LUT4 \DLX_EXinst__n0006<18>149_SW0  (
    .ADR0(DLX_IDinst_IR_function_field[4]),
    .ADR1(DLX_EXinst__n0077),
    .ADR2(DLX_IDinst_IR_function_field[2]),
    .ADR3(CHOICE5437),
    .O(\CHOICE5437/GROM )
  );
  X_BUF \CHOICE5437/XUSED  (
    .I(\CHOICE5437/FROM ),
    .O(CHOICE5437)
  );
  X_BUF \CHOICE5437/YUSED  (
    .I(\CHOICE5437/GROM ),
    .O(N126398)
  );
  defparam \DLX_EXinst__n0006<18>302 .INIT = 16'hB3A0;
  X_LUT4 \DLX_EXinst__n0006<18>302  (
    .ADR0(N111221),
    .ADR1(N110935),
    .ADR2(N101009),
    .ADR3(N126370),
    .O(\CHOICE5476/FROM )
  );
  defparam \DLX_EXinst__n0006<18>343_SW0 .INIT = 16'h8F88;
  X_LUT4 \DLX_EXinst__n0006<18>343_SW0  (
    .ADR0(N101725),
    .ADR1(DLX_EXinst_ALU_result[18]),
    .ADR2(DLX_IDinst_reg_out_B[4]),
    .ADR3(CHOICE5476),
    .O(\CHOICE5476/GROM )
  );
  X_BUF \CHOICE5476/XUSED  (
    .I(\CHOICE5476/FROM ),
    .O(CHOICE5476)
  );
  X_BUF \CHOICE5476/YUSED  (
    .I(\CHOICE5476/GROM ),
    .O(N126366)
  );
  defparam \DLX_EXinst__n0006<26>216 .INIT = 16'hF8F8;
  X_LUT4 \DLX_EXinst__n0006<26>216  (
    .ADR0(DLX_IDinst_reg_out_B[26]),
    .ADR1(DLX_EXinst__n0045),
    .ADR2(DLX_EXinst_N64448),
    .ADR3(VCC),
    .O(\CHOICE4725/FROM )
  );
  defparam \DLX_EXinst__n0006<26>225 .INIT = 16'hCC08;
  X_LUT4 \DLX_EXinst__n0006<26>225  (
    .ADR0(DLX_EXinst__n0047),
    .ADR1(DLX_IDinst_reg_out_A[26]),
    .ADR2(DLX_IDinst_reg_out_B[26]),
    .ADR3(CHOICE4725),
    .O(\CHOICE4725/GROM )
  );
  X_BUF \CHOICE4725/XUSED  (
    .I(\CHOICE4725/FROM ),
    .O(CHOICE4725)
  );
  X_BUF \CHOICE4725/YUSED  (
    .I(\CHOICE4725/GROM ),
    .O(CHOICE4727)
  );
  defparam \DLX_EXinst__n0006<26>240 .INIT = 16'hFFEC;
  X_LUT4 \DLX_EXinst__n0006<26>240  (
    .ADR0(DLX_EXinst__n0016[26]),
    .ADR1(N126354),
    .ADR2(DLX_EXinst__n0114),
    .ADR3(CHOICE4727),
    .O(\CHOICE4731/FROM )
  );
  defparam \DLX_EXinst__n0006<26>268 .INIT = 16'hF0E0;
  X_LUT4 \DLX_EXinst__n0006<26>268  (
    .ADR0(CHOICE4708),
    .ADR1(CHOICE4717),
    .ADR2(DLX_EXinst__n0030),
    .ADR3(CHOICE4731),
    .O(\CHOICE4731/GROM )
  );
  X_BUF \CHOICE4731/XUSED  (
    .I(\CHOICE4731/FROM ),
    .O(CHOICE4731)
  );
  X_BUF \CHOICE4731/YUSED  (
    .I(\CHOICE4731/GROM ),
    .O(CHOICE4733)
  );
  defparam DLX_MEMlc_md_mda14_a1.INIT = 16'h0F00;
  X_LUT4 DLX_MEMlc_md_mda14_a1 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_MEMlc_pd_wint1),
    .ADR3(DLX_MEMlc_md_wint13),
    .O(\DLX_MEMlc_md_wint14/FROM )
  );
  defparam DLX_MEMlc_md_mda15_a1.INIT = 16'h3300;
  X_LUT4 DLX_MEMlc_md_mda15_a1 (
    .ADR0(VCC),
    .ADR1(DLX_MEMlc_pd_wint1),
    .ADR2(VCC),
    .ADR3(DLX_MEMlc_md_wint14),
    .O(\DLX_MEMlc_md_wint14/GROM )
  );
  X_BUF \DLX_MEMlc_md_wint14/XUSED  (
    .I(\DLX_MEMlc_md_wint14/FROM ),
    .O(DLX_MEMlc_md_wint14)
  );
  X_BUF \DLX_MEMlc_md_wint14/YUSED  (
    .I(\DLX_MEMlc_md_wint14/GROM ),
    .O(DLX_MEMlc_md_wint15)
  );
  defparam \DLX_EXinst__n0006<18>227 .INIT = 16'hFAF0;
  X_LUT4 \DLX_EXinst__n0006<18>227  (
    .ADR0(DLX_EXinst__n0045),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N64448),
    .ADR3(DLX_IDinst_reg_out_B[18]),
    .O(\CHOICE5459/FROM )
  );
  defparam \DLX_EXinst__n0006<18>236 .INIT = 16'hF040;
  X_LUT4 \DLX_EXinst__n0006<18>236  (
    .ADR0(DLX_IDinst_reg_out_B[18]),
    .ADR1(DLX_EXinst__n0047),
    .ADR2(DLX_IDinst_reg_out_A[18]),
    .ADR3(CHOICE5459),
    .O(\CHOICE5459/GROM )
  );
  X_BUF \CHOICE5459/XUSED  (
    .I(\CHOICE5459/FROM ),
    .O(CHOICE5459)
  );
  X_BUF \CHOICE5459/YUSED  (
    .I(\CHOICE5459/GROM ),
    .O(CHOICE5461)
  );
  defparam \DLX_EXinst__n0006<26>172 .INIT = 16'h0D08;
  X_LUT4 \DLX_EXinst__n0006<26>172  (
    .ADR0(DLX_IDinst_reg_out_B[2]),
    .ADR1(DLX_EXinst_N64099),
    .ADR2(DLX_IDinst_reg_out_B[4]),
    .ADR3(N97017),
    .O(\CHOICE4715/FROM )
  );
  defparam \DLX_EXinst__n0006<26>185 .INIT = 16'hF080;
  X_LUT4 \DLX_EXinst__n0006<26>185  (
    .ADR0(\DLX_EXinst_Mshift__n0025_Sh[42] ),
    .ADR1(DLX_IDinst_reg_out_B[4]),
    .ADR2(DLX_EXinst_N66226),
    .ADR3(CHOICE4715),
    .O(\CHOICE4715/GROM )
  );
  X_BUF \CHOICE4715/XUSED  (
    .I(\CHOICE4715/FROM ),
    .O(CHOICE4715)
  );
  X_BUF \CHOICE4715/YUSED  (
    .I(\CHOICE4715/GROM ),
    .O(CHOICE4717)
  );
  defparam DLX_IDlc_slave_ctrlID__n00021.INIT = 16'h1011;
  X_LUT4 DLX_IDlc_slave_ctrlID__n00021 (
    .ADR0(reset_IBUF_3),
    .ADR1(DLX_IDlc_slave_ctrlID_l),
    .ADR2(DLX_reqout_ID),
    .ADR3(DLX_ackout_ID),
    .O(\DLX_reqout_ID/FROM )
  );
  defparam DLX_EXlc_pd_wint11.INIT = 16'h00FF;
  X_LUT4 DLX_EXlc_pd_wint11 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_reqout_ID),
    .O(\DLX_reqout_ID/GROM )
  );
  X_BUF \DLX_reqout_ID/XUSED  (
    .I(\DLX_reqout_ID/FROM ),
    .O(DLX_reqout_ID)
  );
  X_BUF \DLX_reqout_ID/YUSED  (
    .I(\DLX_reqout_ID/GROM ),
    .O(DLX_EXlc_pd_wint1)
  );
  defparam \vga_top_vga1_redout<1>1 .INIT = 16'h0300;
  X_LUT4 \vga_top_vga1_redout<1>1  (
    .ADR0(VCC),
    .ADR1(vram_out_vga_eff),
    .ADR2(reset_IBUF_1),
    .ADR3(vga_top_vga1_videoon),
    .O(\red_1_OBUF/FROM )
  );
  defparam \vga_top_vga1_blueout<0>1 .INIT = 16'h1100;
  X_LUT4 \vga_top_vga1_blueout<0>1  (
    .ADR0(reset_IBUF_1),
    .ADR1(vram_out_vga_eff),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_videoon),
    .O(\red_1_OBUF/GROM )
  );
  X_BUF \red_1_OBUF/XUSED  (
    .I(\red_1_OBUF/FROM ),
    .O(red_1_OBUF)
  );
  X_BUF \red_1_OBUF/YUSED  (
    .I(\red_1_OBUF/GROM ),
    .O(blue_0_OBUF)
  );
  defparam \DLX_EXinst__n0006<18>343 .INIT = 16'hFEFA;
  X_LUT4 \DLX_EXinst__n0006<18>343  (
    .ADR0(N126366),
    .ADR1(DLX_EXinst__n0016[18]),
    .ADR2(CHOICE5461),
    .ADR3(DLX_EXinst__n0114),
    .O(\CHOICE5480/FROM )
  );
  defparam \DLX_EXinst__n0006<18>371 .INIT = 16'hCCC8;
  X_LUT4 \DLX_EXinst__n0006<18>371  (
    .ADR0(CHOICE5451),
    .ADR1(DLX_EXinst__n0030),
    .ADR2(CHOICE5447),
    .ADR3(CHOICE5480),
    .O(\CHOICE5480/GROM )
  );
  X_BUF \CHOICE5480/XUSED  (
    .I(\CHOICE5480/FROM ),
    .O(CHOICE5480)
  );
  X_BUF \CHOICE5480/YUSED  (
    .I(\CHOICE5480/GROM ),
    .O(CHOICE5482)
  );
  defparam Ker5730284.INIT = 16'hAAFC;
  X_LUT4 Ker5730284 (
    .ADR0(vram_out_cpu[0]),
    .ADR1(N126029),
    .ADR2(CHOICE2941),
    .ADR3(vga_select_6[1]),
    .O(\N107291/FROM )
  );
  defparam \DM_read_data<0>1 .INIT = 16'hDD88;
  X_LUT4 \DM_read_data<0>1  (
    .ADR0(vga_select_6[0]),
    .ADR1(RAM_read_data[0]),
    .ADR2(VCC),
    .ADR3(N107291),
    .O(\N107291/GROM )
  );
  X_BUF \N107291/XUSED  (
    .I(\N107291/FROM ),
    .O(N107291)
  );
  X_BUF \N107291/YUSED  (
    .I(\N107291/GROM ),
    .O(DM_read_data[0])
  );
  defparam \DLX_EXinst_Mshift__n0025_Sh<7> .INIT = 16'hFC0C;
  X_LUT4 \DLX_EXinst_Mshift__n0025_Sh<7>  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N62851),
    .ADR2(DLX_IDinst_reg_out_B[0]),
    .ADR3(N94305),
    .O(\DLX_EXinst_Mshift__n0025_Sh<7>/FROM )
  );
  defparam DLX_EXinst_Ker629141.INIT = 16'hFDA8;
  X_LUT4 DLX_EXinst_Ker629141 (
    .ADR0(DLX_IDinst_reg_out_B_2_1),
    .ADR1(CHOICE1054),
    .ADR2(CHOICE1060),
    .ADR3(\DLX_EXinst_Mshift__n0025_Sh[7] ),
    .O(\DLX_EXinst_Mshift__n0025_Sh<7>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0025_Sh<7>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0025_Sh<7>/FROM ),
    .O(\DLX_EXinst_Mshift__n0025_Sh[7] )
  );
  X_BUF \DLX_EXinst_Mshift__n0025_Sh<7>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0025_Sh<7>/GROM ),
    .O(DLX_EXinst_N62916)
  );
  defparam \DLX_EXinst__n0006<19>149_SW0 .INIT = 16'hF444;
  X_LUT4 \DLX_EXinst__n0006<19>149_SW0  (
    .ADR0(DLX_IDinst_IR_function_field[4]),
    .ADR1(CHOICE4970),
    .ADR2(DLX_IDinst_IR_function_field[3]),
    .ADR3(DLX_EXinst__n0077),
    .O(\N126542/FROM )
  );
  defparam \DLX_EXinst__n0006<19>149 .INIT = 16'hFFEC;
  X_LUT4 \DLX_EXinst__n0006<19>149  (
    .ADR0(DLX_EXinst__n0128),
    .ADR1(CHOICE4954),
    .ADR2(DLX_EXinst__n0016[19]),
    .ADR3(N126542),
    .O(\N126542/GROM )
  );
  X_BUF \N126542/XUSED  (
    .I(\N126542/FROM ),
    .O(N126542)
  );
  X_BUF \N126542/YUSED  (
    .I(\N126542/GROM ),
    .O(CHOICE4973)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_inv_11.INIT = 16'h3F03;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_inv_11 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[31]),
    .ADR2(DLX_EXinst_Mcompar__n0095_inst_cy_260),
    .ADR3(DLX_IDinst_Imm_31_1),
    .O(\DLX_EXinst__n0095/FROM )
  );
  defparam \DLX_EXinst__n0006<0>392 .INIT = 16'hA820;
  X_LUT4 \DLX_EXinst__n0006<0>392  (
    .ADR0(DLX_IDinst_IR_opcode_field[0]),
    .ADR1(DLX_IDinst_IR_opcode_field[2]),
    .ADR2(DLX_EXinst__n0087),
    .ADR3(DLX_EXinst__n0095),
    .O(\DLX_EXinst__n0095/GROM )
  );
  X_BUF \DLX_EXinst__n0095/XUSED  (
    .I(\DLX_EXinst__n0095/FROM ),
    .O(DLX_EXinst__n0095)
  );
  X_BUF \DLX_EXinst__n0095/YUSED  (
    .I(\DLX_EXinst__n0095/GROM ),
    .O(CHOICE5928)
  );
  defparam \DLX_IFinst__n0001<26>_SW0 .INIT = 16'h05AF;
  X_LUT4 \DLX_IFinst__n0001<26>_SW0  (
    .ADR0(DLX_IFinst__n0000),
    .ADR1(VCC),
    .ADR2(DLX_IFinst__n0015[26]),
    .ADR3(DLX_IFinst_PC[26]),
    .O(\DLX_IFinst_NPC<26>/FROM )
  );
  defparam \DLX_IFinst__n0001<26> .INIT = 16'hC0CF;
  X_LUT4 \DLX_IFinst__n0001<26>  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_branch_address[26]),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(N91723),
    .O(DLX_IFinst__n0001[26])
  );
  X_BUF \DLX_IFinst_NPC<26>/XUSED  (
    .I(\DLX_IFinst_NPC<26>/FROM ),
    .O(N91723)
  );
  defparam \DLX_EXinst__n0006<27>75_SW0 .INIT = 16'hEECC;
  X_LUT4 \DLX_EXinst__n0006<27>75_SW0  (
    .ADR0(DLX_EXinst__n0082),
    .ADR1(CHOICE4628),
    .ADR2(VCC),
    .ADR3(\DLX_EXinst_Mshift__n0028_Sh[59] ),
    .O(\N126432/FROM )
  );
  defparam \DLX_EXinst__n0006<27>75 .INIT = 16'h8F88;
  X_LUT4 \DLX_EXinst__n0006<27>75  (
    .ADR0(N101253),
    .ADR1(N110065),
    .ADR2(N109130),
    .ADR3(N126432),
    .O(\N126432/GROM )
  );
  X_BUF \N126432/XUSED  (
    .I(\N126432/FROM ),
    .O(N126432)
  );
  X_BUF \N126432/YUSED  (
    .I(\N126432/GROM ),
    .O(CHOICE4633)
  );
  defparam \DLX_IFinst__n0001<18>_SW0 .INIT = 16'h4477;
  X_LUT4 \DLX_IFinst__n0001<18>_SW0  (
    .ADR0(DLX_IFinst_PC[18]),
    .ADR1(DLX_IFinst__n0000),
    .ADR2(VCC),
    .ADR3(DLX_IFinst__n0015[18]),
    .O(\DLX_IFinst_NPC<18>/FROM )
  );
  defparam \DLX_IFinst__n0001<18> .INIT = 16'hA0AF;
  X_LUT4 \DLX_IFinst__n0001<18>  (
    .ADR0(DLX_IDinst_branch_address[18]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(N92191),
    .O(DLX_IFinst__n0001[18])
  );
  X_BUF \DLX_IFinst_NPC<18>/XUSED  (
    .I(\DLX_IFinst_NPC<18>/FROM ),
    .O(N92191)
  );
  defparam \DLX_EXinst__n0006<27>216 .INIT = 16'hEEAA;
  X_LUT4 \DLX_EXinst__n0006<27>216  (
    .ADR0(DLX_EXinst_N64448),
    .ADR1(DLX_EXinst__n0045),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[27]),
    .O(\CHOICE4660/FROM )
  );
  defparam \DLX_EXinst__n0006<27>225 .INIT = 16'hAA20;
  X_LUT4 \DLX_EXinst__n0006<27>225  (
    .ADR0(DLX_IDinst_reg_out_A[27]),
    .ADR1(DLX_IDinst_reg_out_B[27]),
    .ADR2(DLX_EXinst__n0047),
    .ADR3(CHOICE4660),
    .O(\CHOICE4660/GROM )
  );
  X_BUF \CHOICE4660/XUSED  (
    .I(\CHOICE4660/FROM ),
    .O(CHOICE4660)
  );
  X_BUF \CHOICE4660/YUSED  (
    .I(\CHOICE4660/GROM ),
    .O(CHOICE4662)
  );
  defparam \DLX_EXinst__n0006<27>240 .INIT = 16'hFEFA;
  X_LUT4 \DLX_EXinst__n0006<27>240  (
    .ADR0(N126411),
    .ADR1(DLX_EXinst__n0114),
    .ADR2(CHOICE4662),
    .ADR3(DLX_EXinst__n0016[27]),
    .O(\CHOICE4666/FROM )
  );
  defparam \DLX_EXinst__n0006<27>268 .INIT = 16'hAAA8;
  X_LUT4 \DLX_EXinst__n0006<27>268  (
    .ADR0(DLX_EXinst__n0030),
    .ADR1(CHOICE4643),
    .ADR2(CHOICE4652),
    .ADR3(CHOICE4666),
    .O(\CHOICE4666/GROM )
  );
  X_BUF \CHOICE4666/XUSED  (
    .I(\CHOICE4666/FROM ),
    .O(CHOICE4666)
  );
  X_BUF \CHOICE4666/YUSED  (
    .I(\CHOICE4666/GROM ),
    .O(CHOICE4668)
  );
  defparam DLX_MEMlc_md_mda18_a1.INIT = 16'h0C0C;
  X_LUT4 DLX_MEMlc_md_mda18_a1 (
    .ADR0(VCC),
    .ADR1(DLX_MEMlc_md_wint17),
    .ADR2(DLX_MEMlc_pd_wint1),
    .ADR3(VCC),
    .O(\DLX_MEMlc_md_wint18/FROM )
  );
  defparam DLX_MEMlc_md_mda16_a1.INIT = 16'h0C0C;
  X_LUT4 DLX_MEMlc_md_mda16_a1 (
    .ADR0(VCC),
    .ADR1(DLX_MEMlc_md_wint15),
    .ADR2(DLX_MEMlc_pd_wint1),
    .ADR3(VCC),
    .O(\DLX_MEMlc_md_wint18/GROM )
  );
  X_BUF \DLX_MEMlc_md_wint18/XUSED  (
    .I(\DLX_MEMlc_md_wint18/FROM ),
    .O(DLX_MEMlc_md_wint18)
  );
  X_BUF \DLX_MEMlc_md_wint18/YUSED  (
    .I(\DLX_MEMlc_md_wint18/GROM ),
    .O(DLX_MEMlc_md_wint16)
  );
  defparam \DLX_EXinst__n0006<27>172 .INIT = 16'h4450;
  X_LUT4 \DLX_EXinst__n0006<27>172  (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(DLX_EXinst_N64104),
    .ADR2(N100843),
    .ADR3(DLX_IDinst_reg_out_B[2]),
    .O(\CHOICE4650/FROM )
  );
  defparam \DLX_EXinst__n0006<27>185 .INIT = 16'hCC80;
  X_LUT4 \DLX_EXinst__n0006<27>185  (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(DLX_EXinst_N66226),
    .ADR2(\DLX_EXinst_Mshift__n0025_Sh[43] ),
    .ADR3(CHOICE4650),
    .O(\CHOICE4650/GROM )
  );
  X_BUF \CHOICE4650/XUSED  (
    .I(\CHOICE4650/FROM ),
    .O(CHOICE4650)
  );
  X_BUF \CHOICE4650/YUSED  (
    .I(\CHOICE4650/GROM ),
    .O(CHOICE4652)
  );
  defparam \DLX_EXinst__n0006<19>309 .INIT = 16'hAE0C;
  X_LUT4 \DLX_EXinst__n0006<19>309  (
    .ADR0(N126482),
    .ADR1(N107444),
    .ADR2(DLX_IDinst_reg_out_B[4]),
    .ADR3(DLX_IDinst_reg_out_A[19]),
    .O(\CHOICE5008/GROM )
  );
  X_BUF \CHOICE5008/YUSED  (
    .I(\CHOICE5008/GROM ),
    .O(CHOICE5008)
  );
  defparam DLX_EXinst_Ker65153107.INIT = 16'hECA0;
  X_LUT4 DLX_EXinst_Ker65153107 (
    .ADR0(CHOICE3077),
    .ADR1(N110065),
    .ADR2(DLX_EXinst_N66507),
    .ADR3(N126469),
    .O(\N108101/FROM )
  );
  defparam \DLX_EXinst__n0006<6>93 .INIT = 16'hFEFC;
  X_LUT4 \DLX_EXinst__n0006<6>93  (
    .ADR0(DLX_IDinst_IR_function_field[4]),
    .ADR1(CHOICE4371),
    .ADR2(CHOICE4354),
    .ADR3(N108101),
    .O(\N108101/GROM )
  );
  X_BUF \N108101/XUSED  (
    .I(\N108101/FROM ),
    .O(N108101)
  );
  X_BUF \N108101/YUSED  (
    .I(\N108101/GROM ),
    .O(CHOICE4372)
  );
  defparam DLX_MEMlc_md_mda19_a1.INIT = 16'h2222;
  X_LUT4 DLX_MEMlc_md_mda19_a1 (
    .ADR0(DLX_MEMlc_md_wint18),
    .ADR1(DLX_MEMlc_pd_wint1),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_MEMlc_md_wint19/FROM )
  );
  defparam DLX_MEMlc_md_mda17_a1.INIT = 16'h4444;
  X_LUT4 DLX_MEMlc_md_mda17_a1 (
    .ADR0(DLX_MEMlc_pd_wint1),
    .ADR1(DLX_MEMlc_md_wint16),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_MEMlc_md_wint19/GROM )
  );
  X_BUF \DLX_MEMlc_md_wint19/XUSED  (
    .I(\DLX_MEMlc_md_wint19/FROM ),
    .O(DLX_MEMlc_md_wint19)
  );
  X_BUF \DLX_MEMlc_md_wint19/YUSED  (
    .I(\DLX_MEMlc_md_wint19/GROM ),
    .O(DLX_MEMlc_md_wint17)
  );
  defparam \DLX_IFinst__n0001<6>_SW0 .INIT = 16'h5533;
  X_LUT4 \DLX_IFinst__n0001<6>_SW0  (
    .ADR0(DLX_IFinst_PC[6]),
    .ADR1(DLX_IFinst__n0015[6]),
    .ADR2(VCC),
    .ADR3(DLX_IFinst__n0000),
    .O(\DLX_IFinst_NPC<6>/FROM )
  );
  defparam \DLX_IFinst__n0001<6> .INIT = 16'hC0F3;
  X_LUT4 \DLX_IFinst__n0001<6>  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(DLX_IDinst_branch_address[6]),
    .ADR3(N92867),
    .O(\DLX_IFinst_NPC<6>/GROM )
  );
  X_BUF \DLX_IFinst_NPC<6>/XUSED  (
    .I(\DLX_IFinst_NPC<6>/FROM ),
    .O(N92867)
  );
  X_BUF \DLX_IFinst_NPC<6>/YUSED  (
    .I(\DLX_IFinst_NPC<6>/GROM ),
    .O(DLX_IFinst__n0001[6])
  );
  defparam DLX_IDinst__n0109153_SW0.INIT = 16'hF0F8;
  X_LUT4 DLX_IDinst__n0109153_SW0 (
    .ADR0(DLX_IDinst_N69781),
    .ADR1(CHOICE3526),
    .ADR2(CHOICE3460),
    .ADR3(DLX_IDinst__n0364),
    .O(\DLX_IDinst_reg_write/FROM )
  );
  defparam DLX_IDinst__n0109153.INIT = 16'h4000;
  X_LUT4 DLX_IDinst__n0109153 (
    .ADR0(DLX_IDinst_intr_slot),
    .ADR1(DLX_EXinst__n0149),
    .ADR2(N95693),
    .ADR3(N127167),
    .O(N110803)
  );
  X_BUF \DLX_IDinst_reg_write/XUSED  (
    .I(\DLX_IDinst_reg_write/FROM ),
    .O(N127167)
  );
  defparam DLX_IDlc_pd_wint11.INIT = 16'h5555;
  X_LUT4 DLX_IDlc_pd_wint11 (
    .ADR0(DLX_reqin_ID),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IDlc_pd_wint1/FROM )
  );
  defparam DLX_IDlc_md_mda40_a1.INIT = 16'h00CC;
  X_LUT4 DLX_IDlc_md_mda40_a1 (
    .ADR0(VCC),
    .ADR1(DLX_IDlc_md_wint39),
    .ADR2(VCC),
    .ADR3(DLX_IDlc_pd_wint1),
    .O(\DLX_IDlc_pd_wint1/GROM )
  );
  X_BUF \DLX_IDlc_pd_wint1/XUSED  (
    .I(\DLX_IDlc_pd_wint1/FROM ),
    .O(DLX_IDlc_pd_wint1)
  );
  X_BUF \DLX_IDlc_pd_wint1/YUSED  (
    .I(\DLX_IDlc_pd_wint1/GROM ),
    .O(DLX_IDlc_md_wint40)
  );
  defparam \DLX_IDinst__n0116<0>44_SW0 .INIT = 16'h00EF;
  X_LUT4 \DLX_IDinst__n0116<0>44_SW0  (
    .ADR0(DLX_IDinst_intr_slot),
    .ADR1(DLX_IDinst_counter[1]),
    .ADR2(N95693),
    .ADR3(DLX_IDinst_counter[0]),
    .O(\DLX_IDinst_counter<0>/FROM )
  );
  defparam \DLX_IDinst__n0116<0>44 .INIT = 16'hFF80;
  X_LUT4 \DLX_IDinst__n0116<0>44  (
    .ADR0(CHOICE2927),
    .ADR1(DLX_IDinst_N70679),
    .ADR2(DLX_IDinst_N70821),
    .ADR3(N126820),
    .O(N107173)
  );
  X_BUF \DLX_IDinst_counter<0>/XUSED  (
    .I(\DLX_IDinst_counter<0>/FROM ),
    .O(N126820)
  );
  defparam \DLX_EXinst_Mshift__n0024_Sh<127>1 .INIT = 16'h0002;
  X_LUT4 \DLX_EXinst_Mshift__n0024_Sh<127>1  (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(DLX_EXinst_N62733),
    .ADR2(DLX_IDinst_IR_function_field_1_1),
    .ADR3(DLX_IDinst_IR_function_field_0_1),
    .O(\DLX_EXinst_Mshift__n0024_Sh<127>/FROM )
  );
  defparam \DLX_EXinst__n0006<15>72 .INIT = 16'hC808;
  X_LUT4 \DLX_EXinst__n0006<15>72  (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(DLX_EXinst_N66060),
    .ADR2(\DLX_IDinst_Imm[5] ),
    .ADR3(\DLX_EXinst_Mshift__n0024_Sh[127] ),
    .O(\DLX_EXinst_Mshift__n0024_Sh<127>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0024_Sh<127>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0024_Sh<127>/FROM ),
    .O(\DLX_EXinst_Mshift__n0024_Sh[127] )
  );
  X_BUF \DLX_EXinst_Mshift__n0024_Sh<127>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0024_Sh<127>/GROM ),
    .O(CHOICE4828)
  );
  defparam \DLX_EXinst__n0006<29>257 .INIT = 16'hF3F2;
  X_LUT4 \DLX_EXinst__n0006<29>257  (
    .ADR0(CHOICE5374),
    .ADR1(N110935),
    .ADR2(CHOICE5383),
    .ADR3(CHOICE5377),
    .O(\CHOICE5384/FROM )
  );
  defparam \DLX_EXinst__n0006<28>253 .INIT = 16'hF0FE;
  X_LUT4 \DLX_EXinst__n0006<28>253  (
    .ADR0(CHOICE5222),
    .ADR1(CHOICE5223),
    .ADR2(CHOICE5229),
    .ADR3(N110935),
    .O(\CHOICE5384/GROM )
  );
  X_BUF \CHOICE5384/XUSED  (
    .I(\CHOICE5384/FROM ),
    .O(CHOICE5384)
  );
  X_BUF \CHOICE5384/YUSED  (
    .I(\CHOICE5384/GROM ),
    .O(CHOICE5230)
  );
  defparam \DLX_EXinst__n0006<28>280 .INIT = 16'hF400;
  X_LUT4 \DLX_EXinst__n0006<28>280  (
    .ADR0(DLX_IDinst_reg_out_B[28]),
    .ADR1(DLX_EXinst__n0047),
    .ADR2(CHOICE5236),
    .ADR3(DLX_IDinst_reg_out_A[28]),
    .O(\CHOICE5238/FROM )
  );
  defparam \DLX_EXinst__n0006<28>284 .INIT = 16'hFF88;
  X_LUT4 \DLX_EXinst__n0006<28>284  (
    .ADR0(DLX_EXinst_ALU_result[28]),
    .ADR1(N101725),
    .ADR2(VCC),
    .ADR3(CHOICE5238),
    .O(\CHOICE5238/GROM )
  );
  X_BUF \CHOICE5238/XUSED  (
    .I(\CHOICE5238/FROM ),
    .O(CHOICE5238)
  );
  X_BUF \CHOICE5238/YUSED  (
    .I(\CHOICE5238/GROM ),
    .O(CHOICE5239)
  );
  defparam \DLX_EXinst__n0006<28>363 .INIT = 16'hFFF8;
  X_LUT4 \DLX_EXinst__n0006<28>363  (
    .ADR0(DLX_EXinst_N63836),
    .ADR1(DLX_EXinst__n0016[28]),
    .ADR2(N100490),
    .ADR3(N126576),
    .O(\DLX_EXinst_ALU_result<28>/FROM )
  );
  defparam \DLX_EXinst__n0006<28>374 .INIT = 16'h1100;
  X_LUT4 \DLX_EXinst__n0006<28>374  (
    .ADR0(DLX_IDinst_counter[0]),
    .ADR1(DLX_IDinst_counter[1]),
    .ADR2(VCC),
    .ADR3(CHOICE5249),
    .O(N121082)
  );
  X_BUF \DLX_EXinst_ALU_result<28>/XUSED  (
    .I(\DLX_EXinst_ALU_result<28>/FROM ),
    .O(CHOICE5249)
  );
  defparam \DLX_EXinst__n0006<23>272_SW0 .INIT = 16'hFAF0;
  X_LUT4 \DLX_EXinst__n0006<23>272_SW0  (
    .ADR0(CHOICE4074),
    .ADR1(VCC),
    .ADR2(CHOICE4088),
    .ADR3(DLX_EXinst_N66226),
    .O(\N126551/FROM )
  );
  defparam \DLX_EXinst__n0006<23>272 .INIT = 16'hAAA8;
  X_LUT4 \DLX_EXinst__n0006<23>272  (
    .ADR0(DLX_EXinst__n0030),
    .ADR1(CHOICE4079),
    .ADR2(CHOICE4064),
    .ADR3(N126551),
    .O(\N126551/GROM )
  );
  X_BUF \N126551/XUSED  (
    .I(\N126551/FROM ),
    .O(N126551)
  );
  X_BUF \N126551/YUSED  (
    .I(\N126551/GROM ),
    .O(CHOICE4091)
  );
  defparam \DLX_IFinst__n0001<19>_SW0 .INIT = 16'h03CF;
  X_LUT4 \DLX_IFinst__n0001<19>_SW0  (
    .ADR0(VCC),
    .ADR1(DLX_IFinst__n0000),
    .ADR2(DLX_IFinst__n0015[19]),
    .ADR3(DLX_IFinst_PC[19]),
    .O(\DLX_IFinst_NPC<19>/FROM )
  );
  defparam \DLX_IFinst__n0001<19> .INIT = 16'hA0AF;
  X_LUT4 \DLX_IFinst__n0001<19>  (
    .ADR0(DLX_IDinst_branch_address[19]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(N92139),
    .O(DLX_IFinst__n0001[19])
  );
  X_BUF \DLX_IFinst_NPC<19>/XUSED  (
    .I(\DLX_IFinst_NPC<19>/FROM ),
    .O(N92139)
  );
  defparam \DLX_IFinst__n0001<27>_SW0 .INIT = 16'h3355;
  X_LUT4 \DLX_IFinst__n0001<27>_SW0  (
    .ADR0(DLX_IFinst__n0015[27]),
    .ADR1(DLX_IFinst_PC[27]),
    .ADR2(VCC),
    .ADR3(DLX_IFinst__n0000),
    .O(\DLX_IFinst_NPC<27>/FROM )
  );
  defparam \DLX_IFinst__n0001<27> .INIT = 16'hC0F3;
  X_LUT4 \DLX_IFinst__n0001<27>  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(DLX_IDinst_branch_address[27]),
    .ADR3(N91775),
    .O(DLX_IFinst__n0001[27])
  );
  X_BUF \DLX_IFinst_NPC<27>/XUSED  (
    .I(\DLX_IFinst_NPC<27>/FROM ),
    .O(N91775)
  );
  defparam DLX_EXinst_Ker65148108.INIT = 16'hECA0;
  X_LUT4 DLX_EXinst_Ker65148108 (
    .ADR0(N110065),
    .ADR1(DLX_EXinst_N66507),
    .ADR2(CHOICE3097),
    .ADR3(CHOICE3104),
    .O(\N108266/FROM )
  );
  defparam \DLX_EXinst__n0006<5>93 .INIT = 16'hFEEE;
  X_LUT4 \DLX_EXinst__n0006<5>93  (
    .ADR0(CHOICE4422),
    .ADR1(CHOICE4439),
    .ADR2(DLX_IDinst_IR_function_field[4]),
    .ADR3(N108266),
    .O(\N108266/GROM )
  );
  X_BUF \N108266/XUSED  (
    .I(\N108266/FROM ),
    .O(N108266)
  );
  X_BUF \N108266/YUSED  (
    .I(\N108266/GROM ),
    .O(CHOICE4440)
  );
  defparam DLX_IDinst_N695681.INIT = 16'hC3FF;
  X_LUT4 DLX_IDinst_N695681 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_IR_latched[30]),
    .ADR2(DLX_IDinst_IR_latched[27]),
    .ADR3(DLX_IDinst_N70991),
    .O(\DLX_IDinst_N69568/FROM )
  );
  defparam DLX_IDinst__n0111_SW0.INIT = 16'h0100;
  X_LUT4 DLX_IDinst__n0111_SW0 (
    .ADR0(DLX_IDinst__n0331),
    .ADR1(DLX_IDinst__n0364),
    .ADR2(DLX_IDinst_N70918),
    .ADR3(DLX_IDinst_N69568),
    .O(\DLX_IDinst_N69568/GROM )
  );
  X_BUF \DLX_IDinst_N69568/XUSED  (
    .I(\DLX_IDinst_N69568/FROM ),
    .O(DLX_IDinst_N69568)
  );
  X_BUF \DLX_IDinst_N69568/YUSED  (
    .I(\DLX_IDinst_N69568/GROM ),
    .O(N90322)
  );
  defparam \DLX_EXinst_Mshift__n0024_Sh<26>10 .INIT = 16'hC088;
  X_LUT4 \DLX_EXinst_Mshift__n0024_Sh<26>10  (
    .ADR0(DLX_IDinst_reg_out_A[27]),
    .ADR1(DLX_IDinst_IR_function_field_0_1),
    .ADR2(DLX_IDinst_reg_out_A[29]),
    .ADR3(DLX_IDinst_IR_function_field_1_1),
    .O(\CHOICE1114/FROM )
  );
  defparam \DLX_EXinst__n0006<29>166 .INIT = 16'hF404;
  X_LUT4 \DLX_EXinst__n0006<29>166  (
    .ADR0(DLX_EXinst_N63157),
    .ADR1(DLX_IDinst_reg_out_A[29]),
    .ADR2(DLX_IDinst_reg_out_B[3]),
    .ADR3(\DLX_EXinst_Mshift__n0025_Sh[21] ),
    .O(\CHOICE1114/GROM )
  );
  X_BUF \CHOICE1114/XUSED  (
    .I(\CHOICE1114/FROM ),
    .O(CHOICE1114)
  );
  X_BUF \CHOICE1114/YUSED  (
    .I(\CHOICE1114/GROM ),
    .O(CHOICE5368)
  );
  defparam \DLX_EXinst__n0006<29>335 .INIT = 16'hEAC0;
  X_LUT4 \DLX_EXinst__n0006<29>335  (
    .ADR0(DLX_IDinst_reg_out_A[26]),
    .ADR1(N126442),
    .ADR2(DLX_EXinst__n0030),
    .ADR3(DLX_EXinst_N63712),
    .O(\CHOICE5398/GROM )
  );
  X_BUF \CHOICE5398/YUSED  (
    .I(\CHOICE5398/GROM ),
    .O(CHOICE5398)
  );
  defparam DLX_IDinst_Ker6960440.INIT = 16'h00E0;
  X_LUT4 DLX_IDinst_Ker6960440 (
    .ADR0(DLX_IDinst_N70924),
    .ADR1(CHOICE2093),
    .ADR2(CHOICE2099),
    .ADR3(DLX_IDinst__n0135),
    .O(\CHOICE2100/FROM )
  );
  defparam DLX_IDinst_Ker6960449.INIT = 16'hFFAA;
  X_LUT4 DLX_IDinst_Ker6960449 (
    .ADR0(DLX_IDinst_N69963),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(CHOICE2100),
    .O(\CHOICE2100/GROM )
  );
  X_BUF \CHOICE2100/XUSED  (
    .I(\CHOICE2100/FROM ),
    .O(CHOICE2100)
  );
  X_BUF \CHOICE2100/YUSED  (
    .I(\CHOICE2100/GROM ),
    .O(N102453)
  );
  defparam \DLX_IFinst__n0001<7>_SW0 .INIT = 16'h4747;
  X_LUT4 \DLX_IFinst__n0001<7>_SW0  (
    .ADR0(DLX_IFinst_PC[7]),
    .ADR1(DLX_IFinst__n0000),
    .ADR2(DLX_IFinst__n0015[7]),
    .ADR3(VCC),
    .O(\DLX_IFinst_NPC<7>/FROM )
  );
  defparam \DLX_IFinst__n0001<7> .INIT = 16'hC0F3;
  X_LUT4 \DLX_IFinst__n0001<7>  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(DLX_IDinst_branch_address[7]),
    .ADR3(N92763),
    .O(\DLX_IFinst_NPC<7>/GROM )
  );
  X_BUF \DLX_IFinst_NPC<7>/XUSED  (
    .I(\DLX_IFinst_NPC<7>/FROM ),
    .O(N92763)
  );
  X_BUF \DLX_IFinst_NPC<7>/YUSED  (
    .I(\DLX_IFinst_NPC<7>/GROM ),
    .O(DLX_IFinst__n0001[7])
  );
  defparam \DLX_EXinst_Mshift__n0025_Sh<41>_SW0 .INIT = 16'h0257;
  X_LUT4 \DLX_EXinst_Mshift__n0025_Sh<41>_SW0  (
    .ADR0(DLX_IDinst_reg_out_B_2_1),
    .ADR1(CHOICE1066),
    .ADR2(CHOICE1072),
    .ADR3(\DLX_EXinst_Mshift__n0025_Sh[9] ),
    .O(\N94733/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0025_Sh<41> .INIT = 16'h083B;
  X_LUT4 \DLX_EXinst_Mshift__n0025_Sh<41>  (
    .ADR0(\DLX_EXinst_Mshift__n0025_Sh[1] ),
    .ADR1(DLX_IDinst_reg_out_B_3_1),
    .ADR2(DLX_IDinst_reg_out_B_2_1),
    .ADR3(N94733),
    .O(\N94733/GROM )
  );
  X_BUF \N94733/XUSED  (
    .I(\N94733/FROM ),
    .O(N94733)
  );
  X_BUF \N94733/YUSED  (
    .I(\N94733/GROM ),
    .O(\DLX_EXinst_Mshift__n0025_Sh[41] )
  );
  defparam \DLX_EXinst__n0006<29>284 .INIT = 16'hF200;
  X_LUT4 \DLX_EXinst__n0006<29>284  (
    .ADR0(DLX_EXinst__n0047),
    .ADR1(DLX_IDinst_reg_out_B[29]),
    .ADR2(CHOICE5390),
    .ADR3(DLX_IDinst_reg_out_A[29]),
    .O(\CHOICE5392/FROM )
  );
  defparam \DLX_EXinst__n0006<29>288 .INIT = 16'hFFC0;
  X_LUT4 \DLX_EXinst__n0006<29>288  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_ALU_result[29]),
    .ADR2(N101725),
    .ADR3(CHOICE5392),
    .O(\CHOICE5392/GROM )
  );
  X_BUF \CHOICE5392/XUSED  (
    .I(\CHOICE5392/FROM ),
    .O(CHOICE5392)
  );
  X_BUF \CHOICE5392/YUSED  (
    .I(\CHOICE5392/GROM ),
    .O(CHOICE5393)
  );
  defparam DLX_IDlc_master_ctrlID__n00021.INIT = 16'h7373;
  X_LUT4 DLX_IDlc_master_ctrlID__n00021 (
    .ADR0(DLX_IDlc_slave_ctrlID_l),
    .ADR1(DLX_ackin_ID),
    .ADR2(DLX_IDlc_master_ctrlID_nro),
    .ADR3(VCC),
    .O(\DLX_IDlc_master_ctrlID_nro/GROM )
  );
  X_BUF \DLX_IDlc_master_ctrlID_nro/YUSED  (
    .I(\DLX_IDlc_master_ctrlID_nro/GROM ),
    .O(DLX_IDlc_master_ctrlID_nro)
  );
  defparam \DLX_EXinst__n0006<29>367 .INIT = 16'hFFEC;
  X_LUT4 \DLX_EXinst__n0006<29>367  (
    .ADR0(DLX_EXinst_N63836),
    .ADR1(N126437),
    .ADR2(DLX_EXinst__n0016[29]),
    .ADR3(N100490),
    .O(\DLX_EXinst_ALU_result<29>/FROM )
  );
  defparam \DLX_EXinst__n0006<29>378 .INIT = 16'h1100;
  X_LUT4 \DLX_EXinst__n0006<29>378  (
    .ADR0(DLX_IDinst_counter[0]),
    .ADR1(DLX_IDinst_counter[1]),
    .ADR2(VCC),
    .ADR3(CHOICE5403),
    .O(N122016)
  );
  X_BUF \DLX_EXinst_ALU_result<29>/XUSED  (
    .I(\DLX_EXinst_ALU_result<29>/FROM ),
    .O(CHOICE5403)
  );
  defparam DLX_EXinst__n001880_SW1.INIT = 16'hC8EA;
  X_LUT4 DLX_EXinst__n001880_SW1 (
    .ADR0(DLX_IDinst_IR_opcode_field[1]),
    .ADR1(DLX_IDinst_IR_opcode_field[2]),
    .ADR2(DLX_IDinst_IR_opcode_field[3]),
    .ADR3(DLX_IDinst_IR_opcode_field[0]),
    .O(\N126207/FROM )
  );
  defparam \DLX_EXinst__n0006<13>15_SW0 .INIT = 16'h000F;
  X_LUT4 \DLX_EXinst__n0006<13>15_SW0  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[13]),
    .ADR3(DLX_IDinst_IR_opcode_field[0]),
    .O(\N126207/GROM )
  );
  X_BUF \N126207/XUSED  (
    .I(\N126207/FROM ),
    .O(N126207)
  );
  X_BUF \N126207/YUSED  (
    .I(\N126207/GROM ),
    .O(N127326)
  );
  defparam \DLX_EXinst__n0006<20>107_SW0 .INIT = 16'hC0E0;
  X_LUT4 \DLX_EXinst__n0006<20>107_SW0  (
    .ADR0(DLX_EXinst__n0080),
    .ADR1(DLX_EXinst__n0079),
    .ADR2(DLX_IDinst_reg_out_A[20]),
    .ADR3(\DLX_IDinst_Imm[31] ),
    .O(\N126379/FROM )
  );
  defparam \DLX_EXinst__n0006<20>107 .INIT = 16'hFFEA;
  X_LUT4 \DLX_EXinst__n0006<20>107  (
    .ADR0(CHOICE4895),
    .ADR1(DLX_EXinst__n0016[20]),
    .ADR2(DLX_EXinst__n0128),
    .ADR3(N126379),
    .O(\N126379/GROM )
  );
  X_BUF \N126379/XUSED  (
    .I(\N126379/FROM ),
    .O(N126379)
  );
  X_BUF \N126379/YUSED  (
    .I(\N126379/GROM ),
    .O(CHOICE4897)
  );
  defparam \DLX_IFinst__n0001<28>_SW0 .INIT = 16'h2727;
  X_LUT4 \DLX_IFinst__n0001<28>_SW0  (
    .ADR0(DLX_IFinst__n0000),
    .ADR1(DLX_IFinst_PC[28]),
    .ADR2(DLX_IFinst__n0015[28]),
    .ADR3(VCC),
    .O(\DLX_IFinst_NPC<28>/FROM )
  );
  defparam \DLX_IFinst__n0001<28> .INIT = 16'hA0F5;
  X_LUT4 \DLX_IFinst__n0001<28>  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_branch_address[28]),
    .ADR3(N91671),
    .O(DLX_IFinst__n0001[28])
  );
  X_BUF \DLX_IFinst_NPC<28>/XUSED  (
    .I(\DLX_IFinst_NPC<28>/FROM ),
    .O(N91671)
  );
  defparam DLX_IDinst_Ker6963328.INIT = 16'h00BF;
  X_LUT4 DLX_IDinst_Ker6963328 (
    .ADR0(DLX_IDinst__n0331),
    .ADR1(DLX_IDinst__n0387),
    .ADR2(DLX_IDinst_N70918),
    .ADR3(N127551),
    .O(\CHOICE1880/FROM )
  );
  defparam DLX_IDinst_Ker6963336.INIT = 16'h0100;
  X_LUT4 DLX_IDinst_Ker6963336 (
    .ADR0(DLX_IDinst_regA_index[3]),
    .ADR1(DLX_IDinst_regA_index[4]),
    .ADR2(DLX_IDinst_regA_index[2]),
    .ADR3(CHOICE1880),
    .O(\CHOICE1880/GROM )
  );
  X_BUF \CHOICE1880/XUSED  (
    .I(\CHOICE1880/FROM ),
    .O(CHOICE1880)
  );
  X_BUF \CHOICE1880/YUSED  (
    .I(\CHOICE1880/GROM ),
    .O(N101161)
  );
  defparam \DM_read_data<25>1 .INIT = 16'hFAAA;
  X_LUT4 \DM_read_data<25>1  (
    .ADR0(N57312),
    .ADR1(VCC),
    .ADR2(vga_select_6[0]),
    .ADR3(RAM_read_data[25]),
    .O(\DM_read_data<25>/FROM )
  );
  defparam \DM_read_data<10>1 .INIT = 16'hFAF0;
  X_LUT4 \DM_read_data<10>1  (
    .ADR0(RAM_read_data[10]),
    .ADR1(VCC),
    .ADR2(N57312),
    .ADR3(vga_select_6[0]),
    .O(\DM_read_data<25>/GROM )
  );
  X_BUF \DM_read_data<25>/XUSED  (
    .I(\DM_read_data<25>/FROM ),
    .O(DM_read_data[25])
  );
  X_BUF \DM_read_data<25>/YUSED  (
    .I(\DM_read_data<25>/GROM ),
    .O(DM_read_data[10])
  );
  defparam \DLX_IFinst__n0001<8>_SW0 .INIT = 16'h0F55;
  X_LUT4 \DLX_IFinst__n0001<8>_SW0  (
    .ADR0(DLX_IFinst__n0015[8]),
    .ADR1(VCC),
    .ADR2(DLX_IFinst_PC[8]),
    .ADR3(DLX_IFinst__n0000),
    .O(\DLX_IFinst_NPC<8>/FROM )
  );
  defparam \DLX_IFinst__n0001<8> .INIT = 16'hC0F3;
  X_LUT4 \DLX_IFinst__n0001<8>  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(DLX_IDinst_branch_address[8]),
    .ADR3(N92659),
    .O(\DLX_IFinst_NPC<8>/GROM )
  );
  X_BUF \DLX_IFinst_NPC<8>/XUSED  (
    .I(\DLX_IFinst_NPC<8>/FROM ),
    .O(N92659)
  );
  X_BUF \DLX_IFinst_NPC<8>/YUSED  (
    .I(\DLX_IFinst_NPC<8>/GROM ),
    .O(DLX_IFinst__n0001[8])
  );
  defparam \DLX_EXinst_Mshift__n0025_Sh<42>_SW0 .INIT = 16'h111D;
  X_LUT4 \DLX_EXinst_Mshift__n0025_Sh<42>_SW0  (
    .ADR0(\DLX_EXinst_Mshift__n0025_Sh[10] ),
    .ADR1(DLX_IDinst_reg_out_B_2_1),
    .ADR2(CHOICE1300),
    .ADR3(CHOICE1294),
    .O(\N94673/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0025_Sh<42> .INIT = 16'h083B;
  X_LUT4 \DLX_EXinst_Mshift__n0025_Sh<42>  (
    .ADR0(\DLX_EXinst_Mshift__n0025_Sh[2] ),
    .ADR1(DLX_IDinst_reg_out_B_3_1),
    .ADR2(DLX_IDinst_reg_out_B_2_1),
    .ADR3(N94673),
    .O(\N94673/GROM )
  );
  X_BUF \N94673/XUSED  (
    .I(\N94673/FROM ),
    .O(N94673)
  );
  X_BUF \N94673/YUSED  (
    .I(\N94673/GROM ),
    .O(\DLX_EXinst_Mshift__n0025_Sh[42] )
  );
  defparam \DM_read_data<26>1 .INIT = 16'hFCCC;
  X_LUT4 \DM_read_data<26>1  (
    .ADR0(VCC),
    .ADR1(N57312),
    .ADR2(RAM_read_data[26]),
    .ADR3(vga_select_6[0]),
    .O(\DM_read_data<26>/FROM )
  );
  defparam \DM_read_data<11>1 .INIT = 16'hFFA0;
  X_LUT4 \DM_read_data<11>1  (
    .ADR0(RAM_read_data[11]),
    .ADR1(VCC),
    .ADR2(vga_select_6[0]),
    .ADR3(N57312),
    .O(\DM_read_data<26>/GROM )
  );
  X_BUF \DM_read_data<26>/XUSED  (
    .I(\DM_read_data<26>/FROM ),
    .O(DM_read_data[26])
  );
  X_BUF \DM_read_data<26>/YUSED  (
    .I(\DM_read_data<26>/GROM ),
    .O(DM_read_data[11])
  );
  defparam \DLX_EXinst_Mshift__n0028_Sh<30>1 .INIT = 16'h5410;
  X_LUT4 \DLX_EXinst_Mshift__n0028_Sh<30>1  (
    .ADR0(DLX_IDinst_IR_function_field_1_1),
    .ADR1(DLX_IDinst_IR_function_field_0_1),
    .ADR2(DLX_IDinst_reg_out_A[30]),
    .ADR3(DLX_IDinst_reg_out_A[31]),
    .O(\DLX_EXinst_Mshift__n0028_Sh<30>/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0024_Sh<27>_SW0 .INIT = 16'hB8B8;
  X_LUT4 \DLX_EXinst_Mshift__n0024_Sh<27>_SW0  (
    .ADR0(DLX_IDinst_reg_out_A[28]),
    .ADR1(DLX_IDinst_IR_function_field_0_1),
    .ADR2(DLX_IDinst_reg_out_A[27]),
    .ADR3(VCC),
    .O(\DLX_EXinst_Mshift__n0028_Sh<30>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0028_Sh<30>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0028_Sh<30>/FROM ),
    .O(\DLX_EXinst_Mshift__n0028_Sh[30] )
  );
  X_BUF \DLX_EXinst_Mshift__n0028_Sh<30>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0028_Sh<30>/GROM ),
    .O(N93799)
  );
  defparam \DLX_EXinst__n0006<20>300_SW0 .INIT = 16'hFEEE;
  X_LUT4 \DLX_EXinst__n0006<20>300_SW0  (
    .ADR0(CHOICE4915),
    .ADR1(CHOICE4930),
    .ADR2(DLX_EXinst_N66078),
    .ADR3(DLX_EXinst_N64500),
    .O(\N126620/FROM )
  );
  defparam \DLX_EXinst__n0006<20>300 .INIT = 16'hF0E0;
  X_LUT4 \DLX_EXinst__n0006<20>300  (
    .ADR0(CHOICE4904),
    .ADR1(CHOICE4909),
    .ADR2(DLX_EXinst__n0030),
    .ADR3(N126620),
    .O(\N126620/GROM )
  );
  X_BUF \N126620/XUSED  (
    .I(\N126620/FROM ),
    .O(N126620)
  );
  X_BUF \N126620/YUSED  (
    .I(\N126620/GROM ),
    .O(CHOICE4934)
  );
  defparam \DM_read_data<27>1 .INIT = 16'hFF88;
  X_LUT4 \DM_read_data<27>1  (
    .ADR0(RAM_read_data[27]),
    .ADR1(vga_select_6[0]),
    .ADR2(VCC),
    .ADR3(N57312),
    .O(\DM_read_data<27>/FROM )
  );
  defparam \DM_read_data<12>1 .INIT = 16'hEECC;
  X_LUT4 \DM_read_data<12>1  (
    .ADR0(vga_select_6[0]),
    .ADR1(N57312),
    .ADR2(VCC),
    .ADR3(RAM_read_data[12]),
    .O(\DM_read_data<27>/GROM )
  );
  X_BUF \DM_read_data<27>/XUSED  (
    .I(\DM_read_data<27>/FROM ),
    .O(DM_read_data[27])
  );
  X_BUF \DM_read_data<27>/YUSED  (
    .I(\DM_read_data<27>/GROM ),
    .O(DM_read_data[12])
  );
  defparam \DM_read_data<28>1 .INIT = 16'hFAF0;
  X_LUT4 \DM_read_data<28>1  (
    .ADR0(RAM_read_data[28]),
    .ADR1(VCC),
    .ADR2(N57312),
    .ADR3(vga_select_6[0]),
    .O(\DM_read_data<28>/FROM )
  );
  defparam \DM_read_data<20>1 .INIT = 16'hFFA0;
  X_LUT4 \DM_read_data<20>1  (
    .ADR0(vga_select_6[0]),
    .ADR1(VCC),
    .ADR2(RAM_read_data[20]),
    .ADR3(N57312),
    .O(\DM_read_data<28>/GROM )
  );
  X_BUF \DM_read_data<28>/XUSED  (
    .I(\DM_read_data<28>/FROM ),
    .O(DM_read_data[28])
  );
  X_BUF \DM_read_data<28>/YUSED  (
    .I(\DM_read_data<28>/GROM ),
    .O(DM_read_data[20])
  );
  defparam \DLX_EXinst_Mshift__n0024_Sh<26>28 .INIT = 16'hFFAA;
  X_LUT4 \DLX_EXinst_Mshift__n0024_Sh<26>28  (
    .ADR0(CHOICE1120),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(CHOICE1114),
    .O(\DLX_EXinst_Mshift__n0024_Sh<26>/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0028_Sh<58>1 .INIT = 16'h0B08;
  X_LUT4 \DLX_EXinst_Mshift__n0028_Sh<58>1  (
    .ADR0(\DLX_EXinst_Mshift__n0028_Sh[30] ),
    .ADR1(DLX_IDinst_IR_function_field_2_1),
    .ADR2(DLX_IDinst_IR_function_field_3_1),
    .ADR3(\DLX_EXinst_Mshift__n0024_Sh[26] ),
    .O(\DLX_EXinst_Mshift__n0024_Sh<26>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0024_Sh<26>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0024_Sh<26>/FROM ),
    .O(\DLX_EXinst_Mshift__n0024_Sh[26] )
  );
  X_BUF \DLX_EXinst_Mshift__n0024_Sh<26>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0024_Sh<26>/GROM ),
    .O(\DLX_EXinst_Mshift__n0028_Sh[58] )
  );
  defparam DLX_IDinst__n008921_SW0.INIT = 16'hFFA8;
  X_LUT4 DLX_IDinst__n008921_SW0 (
    .ADR0(DLX_IDinst_N69568),
    .ADR1(CHOICE2100),
    .ADR2(DLX_IDinst_N69963),
    .ADR3(DLX_IDinst__n0364),
    .O(\N126776/GROM )
  );
  X_BUF \N126776/YUSED  (
    .I(\N126776/GROM ),
    .O(N126776)
  );
  defparam \DM_read_data<29>1 .INIT = 16'hFAAA;
  X_LUT4 \DM_read_data<29>1  (
    .ADR0(N57312),
    .ADR1(VCC),
    .ADR2(vga_select_6[0]),
    .ADR3(RAM_read_data[29]),
    .O(\DM_read_data<29>/FROM )
  );
  defparam \DM_read_data<13>1 .INIT = 16'hEEAA;
  X_LUT4 \DM_read_data<13>1  (
    .ADR0(N57312),
    .ADR1(vga_select_6[0]),
    .ADR2(VCC),
    .ADR3(RAM_read_data[13]),
    .O(\DM_read_data<29>/GROM )
  );
  X_BUF \DM_read_data<29>/XUSED  (
    .I(\DM_read_data<29>/FROM ),
    .O(DM_read_data[29])
  );
  X_BUF \DM_read_data<29>/YUSED  (
    .I(\DM_read_data<29>/GROM ),
    .O(DM_read_data[13])
  );
  defparam \DM_read_data<31>1 .INIT = 16'hFF88;
  X_LUT4 \DM_read_data<31>1  (
    .ADR0(vga_select_6[0]),
    .ADR1(RAM_read_data[31]),
    .ADR2(VCC),
    .ADR3(N57312),
    .O(\DM_read_data<31>/FROM )
  );
  defparam \DM_read_data<21>1 .INIT = 16'hFAF0;
  X_LUT4 \DM_read_data<21>1  (
    .ADR0(vga_select_6[0]),
    .ADR1(VCC),
    .ADR2(N57312),
    .ADR3(RAM_read_data[21]),
    .O(\DM_read_data<31>/GROM )
  );
  X_BUF \DM_read_data<31>/XUSED  (
    .I(\DM_read_data<31>/FROM ),
    .O(DM_read_data[31])
  );
  X_BUF \DM_read_data<31>/YUSED  (
    .I(\DM_read_data<31>/GROM ),
    .O(DM_read_data[21])
  );
  defparam \vga_top_vga1_redout<0>1 .INIT = 16'h000A;
  X_LUT4 \vga_top_vga1_redout<0>1  (
    .ADR0(vga_top_vga1_videoon),
    .ADR1(VCC),
    .ADR2(reset_IBUF_1),
    .ADR3(vram_out_vga_eff),
    .O(\red_0_OBUF/GROM )
  );
  X_BUF \red_0_OBUF/YUSED  (
    .I(\red_0_OBUF/GROM ),
    .O(red_0_OBUF)
  );
  defparam \DM_read_data<1>1 .INIT = 16'hFFA0;
  X_LUT4 \DM_read_data<1>1  (
    .ADR0(vga_select_6[0]),
    .ADR1(VCC),
    .ADR2(RAM_read_data[1]),
    .ADR3(N57312),
    .O(\DM_read_data<1>/FROM )
  );
  defparam \DM_read_data<14>1 .INIT = 16'hFF88;
  X_LUT4 \DM_read_data<14>1  (
    .ADR0(vga_select_6[0]),
    .ADR1(RAM_read_data[14]),
    .ADR2(VCC),
    .ADR3(N57312),
    .O(\DM_read_data<1>/GROM )
  );
  X_BUF \DM_read_data<1>/XUSED  (
    .I(\DM_read_data<1>/FROM ),
    .O(DM_read_data[1])
  );
  X_BUF \DM_read_data<1>/YUSED  (
    .I(\DM_read_data<1>/GROM ),
    .O(DM_read_data[14])
  );
  defparam \DM_read_data<2>1 .INIT = 16'hEEAA;
  X_LUT4 \DM_read_data<2>1  (
    .ADR0(N57312),
    .ADR1(vga_select_6[0]),
    .ADR2(VCC),
    .ADR3(RAM_read_data[2]),
    .O(\DM_read_data<2>/FROM )
  );
  defparam \DM_read_data<22>1 .INIT = 16'hEECC;
  X_LUT4 \DM_read_data<22>1  (
    .ADR0(vga_select_6[0]),
    .ADR1(N57312),
    .ADR2(VCC),
    .ADR3(RAM_read_data[22]),
    .O(\DM_read_data<2>/GROM )
  );
  X_BUF \DM_read_data<2>/XUSED  (
    .I(\DM_read_data<2>/FROM ),
    .O(DM_read_data[2])
  );
  X_BUF \DM_read_data<2>/YUSED  (
    .I(\DM_read_data<2>/GROM ),
    .O(DM_read_data[22])
  );
  defparam DLX_IDinst_Ker6974431.INIT = 16'hBA30;
  X_LUT4 DLX_IDinst_Ker6974431 (
    .ADR0(CHOICE2112),
    .ADR1(DLX_IDinst__n0448[1]),
    .ADR2(N126580),
    .ADR3(DLX_IDinst_N70985),
    .O(\N102532/FROM )
  );
  defparam DLX_IDinst__n0112_SW0.INIT = 16'hBFFF;
  X_LUT4 DLX_IDinst__n0112_SW0 (
    .ADR0(DLX_IDinst_IR_latched[30]),
    .ADR1(DLX_IDinst__n0132),
    .ADR2(DLX_IDinst__n0338),
    .ADR3(N102532),
    .O(\N102532/GROM )
  );
  X_BUF \N102532/XUSED  (
    .I(\N102532/FROM ),
    .O(N102532)
  );
  X_BUF \N102532/YUSED  (
    .I(\N102532/GROM ),
    .O(N100243)
  );
  defparam DLX_IDinst_Ker6974423.INIT = 16'h5557;
  X_LUT4 DLX_IDinst_Ker6974423 (
    .ADR0(DLX_IDinst_N70909),
    .ADR1(DLX_IDinst_N70635),
    .ADR2(DLX_IDinst__n0250),
    .ADR3(DLX_IDinst__n0252),
    .O(\CHOICE2112/GROM )
  );
  X_BUF \CHOICE2112/YUSED  (
    .I(\CHOICE2112/GROM ),
    .O(CHOICE2112)
  );
  defparam \DLX_EXinst__n0006<19>347_SW0 .INIT = 16'hFAF0;
  X_LUT4 \DLX_EXinst__n0006<19>347_SW0  (
    .ADR0(DLX_EXinst_N66226),
    .ADR1(VCC),
    .ADR2(CHOICE5008),
    .ADR3(CHOICE4994),
    .O(\N126473/FROM )
  );
  defparam \DLX_EXinst__n0006<19>347 .INIT = 16'hAAA8;
  X_LUT4 \DLX_EXinst__n0006<19>347  (
    .ADR0(DLX_EXinst__n0030),
    .ADR1(CHOICE4980),
    .ADR2(CHOICE4999),
    .ADR3(N126473),
    .O(\N126473/GROM )
  );
  X_BUF \N126473/XUSED  (
    .I(\N126473/FROM ),
    .O(N126473)
  );
  X_BUF \N126473/YUSED  (
    .I(\N126473/GROM ),
    .O(CHOICE5011)
  );
  defparam \DM_read_data<3>1 .INIT = 16'hECEC;
  X_LUT4 \DM_read_data<3>1  (
    .ADR0(vga_select_6[0]),
    .ADR1(N57312),
    .ADR2(RAM_read_data[3]),
    .ADR3(VCC),
    .O(\DM_read_data<3>/FROM )
  );
  defparam \DM_read_data<15>1 .INIT = 16'hFCCC;
  X_LUT4 \DM_read_data<15>1  (
    .ADR0(VCC),
    .ADR1(N57312),
    .ADR2(vga_select_6[0]),
    .ADR3(RAM_read_data[15]),
    .O(\DM_read_data<3>/GROM )
  );
  X_BUF \DM_read_data<3>/XUSED  (
    .I(\DM_read_data<3>/FROM ),
    .O(DM_read_data[3])
  );
  X_BUF \DM_read_data<3>/YUSED  (
    .I(\DM_read_data<3>/GROM ),
    .O(DM_read_data[15])
  );
  defparam \DM_read_data<4>1 .INIT = 16'hFAAA;
  X_LUT4 \DM_read_data<4>1  (
    .ADR0(N57312),
    .ADR1(VCC),
    .ADR2(vga_select_6[0]),
    .ADR3(RAM_read_data[4]),
    .O(\DM_read_data<4>/FROM )
  );
  defparam \DM_read_data<23>1 .INIT = 16'hFFA0;
  X_LUT4 \DM_read_data<23>1  (
    .ADR0(vga_select_6[0]),
    .ADR1(VCC),
    .ADR2(RAM_read_data[23]),
    .ADR3(N57312),
    .O(\DM_read_data<4>/GROM )
  );
  X_BUF \DM_read_data<4>/XUSED  (
    .I(\DM_read_data<4>/FROM ),
    .O(DM_read_data[4])
  );
  X_BUF \DM_read_data<4>/YUSED  (
    .I(\DM_read_data<4>/GROM ),
    .O(DM_read_data[23])
  );
  defparam vga_top_vga1__n000839.INIT = 16'hA200;
  X_LUT4 vga_top_vga1__n000839 (
    .ADR0(CHOICE3224),
    .ADR1(vga_top_vga1_vcounter[9]),
    .ADR2(CHOICE3221),
    .ADR3(vga_top_vga1_hcounter[9]),
    .O(\CHOICE3225/FROM )
  );
  defparam vga_top_vga1__n000846.INIT = 16'hAA00;
  X_LUT4 vga_top_vga1__n000846 (
    .ADR0(CHOICE3214),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(CHOICE3225),
    .O(\CHOICE3225/GROM )
  );
  X_BUF \CHOICE3225/XUSED  (
    .I(\CHOICE3225/FROM ),
    .O(CHOICE3225)
  );
  X_BUF \CHOICE3225/YUSED  (
    .I(\CHOICE3225/GROM ),
    .O(N108996)
  );
  defparam \DLX_EXinst_Mshift__n0024_Sh<30>1 .INIT = 16'hABA8;
  X_LUT4 \DLX_EXinst_Mshift__n0024_Sh<30>1  (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(DLX_IDinst_IR_function_field_0_1),
    .ADR2(DLX_IDinst_IR_function_field_1_1),
    .ADR3(DLX_IDinst_reg_out_A[30]),
    .O(\DLX_EXinst_Mshift__n0024_Sh<30>/FROM )
  );
  defparam DLX_EXinst_Ker6582532.INIT = 16'h0100;
  X_LUT4 DLX_EXinst_Ker6582532 (
    .ADR0(DLX_IDinst_IR_function_field_2_1),
    .ADR1(\DLX_IDinst_Imm[5] ),
    .ADR2(DLX_IDinst_IR_function_field_3_1),
    .ADR3(\DLX_EXinst_Mshift__n0024_Sh[30] ),
    .O(\DLX_EXinst_Mshift__n0024_Sh<30>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0024_Sh<30>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0024_Sh<30>/FROM ),
    .O(\DLX_EXinst_Mshift__n0024_Sh[30] )
  );
  X_BUF \DLX_EXinst_Mshift__n0024_Sh<30>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0024_Sh<30>/GROM ),
    .O(CHOICE2064)
  );
  defparam \DLX_EXinst_Mshift__n0024_Sh<28>25 .INIT = 16'h5404;
  X_LUT4 \DLX_EXinst_Mshift__n0024_Sh<28>25  (
    .ADR0(DLX_IDinst_IR_function_field_1_1),
    .ADR1(DLX_IDinst_reg_out_A[28]),
    .ADR2(DLX_IDinst_IR_function_field_0_1),
    .ADR3(DLX_IDinst_reg_out_A[29]),
    .O(\CHOICE1132/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0024_Sh<28>28 .INIT = 16'hFFCC;
  X_LUT4 \DLX_EXinst_Mshift__n0024_Sh<28>28  (
    .ADR0(VCC),
    .ADR1(CHOICE1126),
    .ADR2(VCC),
    .ADR3(CHOICE1132),
    .O(\CHOICE1132/GROM )
  );
  X_BUF \CHOICE1132/XUSED  (
    .I(\CHOICE1132/FROM ),
    .O(CHOICE1132)
  );
  X_BUF \CHOICE1132/YUSED  (
    .I(\CHOICE1132/GROM ),
    .O(\DLX_EXinst_Mshift__n0024_Sh[28] )
  );
  defparam \DLX_IFinst__n0001<29>_SW0 .INIT = 16'h0F33;
  X_LUT4 \DLX_IFinst__n0001<29>_SW0  (
    .ADR0(VCC),
    .ADR1(DLX_IFinst__n0015[29]),
    .ADR2(DLX_IFinst_PC[29]),
    .ADR3(DLX_IFinst__n0000),
    .O(\DLX_IFinst_NPC<29>/FROM )
  );
  defparam \DLX_IFinst__n0001<29> .INIT = 16'hA0F5;
  X_LUT4 \DLX_IFinst__n0001<29>  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_branch_address[29]),
    .ADR3(N91567),
    .O(DLX_IFinst__n0001[29])
  );
  X_BUF \DLX_IFinst_NPC<29>/XUSED  (
    .I(\DLX_IFinst_NPC<29>/FROM ),
    .O(N91567)
  );
  defparam vga_top_vga1__n000962.INIT = 16'hFFF0;
  X_LUT4 vga_top_vga1__n000962 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(vga_top_vga1__n0030),
    .ADR3(vga_top_vga1__n0029),
    .O(\CHOICE3427/GROM )
  );
  X_BUF \CHOICE3427/YUSED  (
    .I(\CHOICE3427/GROM ),
    .O(CHOICE3427)
  );
  defparam \DM_read_data<5>1 .INIT = 16'hFCF0;
  X_LUT4 \DM_read_data<5>1  (
    .ADR0(VCC),
    .ADR1(RAM_read_data[5]),
    .ADR2(N57312),
    .ADR3(vga_select_6[0]),
    .O(\DM_read_data<5>/FROM )
  );
  defparam \DM_read_data<16>1 .INIT = 16'hFAF0;
  X_LUT4 \DM_read_data<16>1  (
    .ADR0(vga_select_6[0]),
    .ADR1(VCC),
    .ADR2(N57312),
    .ADR3(RAM_read_data[16]),
    .O(\DM_read_data<5>/GROM )
  );
  X_BUF \DM_read_data<5>/XUSED  (
    .I(\DM_read_data<5>/FROM ),
    .O(DM_read_data[5])
  );
  X_BUF \DM_read_data<5>/YUSED  (
    .I(\DM_read_data<5>/GROM ),
    .O(DM_read_data[16])
  );
  defparam \DM_read_data<6>1 .INIT = 16'hECEC;
  X_LUT4 \DM_read_data<6>1  (
    .ADR0(vga_select_6[0]),
    .ADR1(N57312),
    .ADR2(RAM_read_data[6]),
    .ADR3(VCC),
    .O(\DM_read_data<6>/FROM )
  );
  defparam \DM_read_data<24>1 .INIT = 16'hFCCC;
  X_LUT4 \DM_read_data<24>1  (
    .ADR0(VCC),
    .ADR1(N57312),
    .ADR2(vga_select_6[0]),
    .ADR3(RAM_read_data[24]),
    .O(\DM_read_data<6>/GROM )
  );
  X_BUF \DM_read_data<6>/XUSED  (
    .I(\DM_read_data<6>/FROM ),
    .O(DM_read_data[6])
  );
  X_BUF \DM_read_data<6>/YUSED  (
    .I(\DM_read_data<6>/GROM ),
    .O(DM_read_data[24])
  );
  defparam DLX_IDinst_Ker70033_SW0.INIT = 16'h0008;
  X_LUT4 DLX_IDinst_Ker70033_SW0 (
    .ADR0(DLX_IDinst_N70924),
    .ADR1(DLX_IDinst_N70991),
    .ADR2(DLX_IDinst_IR_latched[27]),
    .ADR3(DLX_IDinst_IR_latched[30]),
    .O(\N90291/FROM )
  );
  defparam DLX_IDinst_Ker70033.INIT = 16'hFF20;
  X_LUT4 DLX_IDinst_Ker70033 (
    .ADR0(DLX_IDinst_N70909),
    .ADR1(DLX_IDinst__n0348),
    .ADR2(DLX_IDinst__n0252),
    .ADR3(N90291),
    .O(\N90291/GROM )
  );
  X_BUF \N90291/XUSED  (
    .I(\N90291/FROM ),
    .O(N90291)
  );
  X_BUF \N90291/YUSED  (
    .I(\N90291/GROM ),
    .O(DLX_IDinst_N70035)
  );
  defparam \DM_read_data<7>1 .INIT = 16'hFAAA;
  X_LUT4 \DM_read_data<7>1  (
    .ADR0(N57312),
    .ADR1(VCC),
    .ADR2(vga_select_6[0]),
    .ADR3(RAM_read_data[7]),
    .O(\DM_read_data<7>/FROM )
  );
  defparam \DM_read_data<17>1 .INIT = 16'hFAAA;
  X_LUT4 \DM_read_data<17>1  (
    .ADR0(N57312),
    .ADR1(VCC),
    .ADR2(RAM_read_data[17]),
    .ADR3(vga_select_6[0]),
    .O(\DM_read_data<7>/GROM )
  );
  X_BUF \DM_read_data<7>/XUSED  (
    .I(\DM_read_data<7>/FROM ),
    .O(DM_read_data[7])
  );
  X_BUF \DM_read_data<7>/YUSED  (
    .I(\DM_read_data<7>/GROM ),
    .O(DM_read_data[17])
  );
  X_INV \DLX_MEMinst_reg_write_MEM/CKINV  (
    .I(DLX_MEMlc_master_ctrlMEM_l),
    .O(\DLX_MEMinst_reg_write_MEM/CKMUXNOT )
  );
  defparam DLX_IFlc_slave_ctrlIF__n0001_SW18.INIT = 16'hFEFA;
  X_LUT4 DLX_IFlc_slave_ctrlIF__n0001_SW18 (
    .ADR0(reset_IBUF_1),
    .ADR1(DLX_reqout_IF),
    .ADR2(DLX_IFlc_slave_ctrlIF_l),
    .ADR3(DLX_ackin_ID),
    .O(\CHOICE25/FROM )
  );
  defparam DLX_IFlc_slave_ctrlIF__n0001_SW19.INIT = 16'hAA00;
  X_LUT4 DLX_IFlc_slave_ctrlIF__n0001_SW19 (
    .ADR0(DLX_IFlc_master_ctrlIF_nro),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(CHOICE25),
    .O(\CHOICE25/GROM )
  );
  X_BUF \CHOICE25/XUSED  (
    .I(\CHOICE25/FROM ),
    .O(CHOICE25)
  );
  X_BUF \CHOICE25/YUSED  (
    .I(\CHOICE25/GROM ),
    .O(DLX_IFlc_slave_ctrlIF_l)
  );
  defparam \DLX_EXinst_Mshift__n0028_Sh<21>1 .INIT = 16'hAFA0;
  X_LUT4 \DLX_EXinst_Mshift__n0028_Sh<21>1  (
    .ADR0(DLX_EXinst_N63519),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_IR_function_field_0_1),
    .ADR3(DLX_EXinst_N63011),
    .O(\DLX_EXinst_Mshift__n0028_Sh<21>/FROM )
  );
  defparam DLX_EXinst_Ker630191.INIT = 16'hF3C0;
  X_LUT4 DLX_EXinst_Ker630191 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_IR_function_field[3]),
    .ADR2(\DLX_EXinst_Mshift__n0028_Sh[29] ),
    .ADR3(\DLX_EXinst_Mshift__n0028_Sh[21] ),
    .O(\DLX_EXinst_Mshift__n0028_Sh<21>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0028_Sh<21>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0028_Sh<21>/FROM ),
    .O(\DLX_EXinst_Mshift__n0028_Sh[21] )
  );
  X_BUF \DLX_EXinst_Mshift__n0028_Sh<21>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0028_Sh<21>/GROM ),
    .O(DLX_EXinst_N63021)
  );
  defparam \DM_read_data<8>1 .INIT = 16'hFAAA;
  X_LUT4 \DM_read_data<8>1  (
    .ADR0(N57312),
    .ADR1(VCC),
    .ADR2(RAM_read_data[8]),
    .ADR3(vga_select_6[0]),
    .O(\DM_read_data<8>/FROM )
  );
  defparam \DM_read_data<18>1 .INIT = 16'hFAAA;
  X_LUT4 \DM_read_data<18>1  (
    .ADR0(N57312),
    .ADR1(VCC),
    .ADR2(vga_select_6[0]),
    .ADR3(RAM_read_data[18]),
    .O(\DM_read_data<8>/GROM )
  );
  X_BUF \DM_read_data<8>/XUSED  (
    .I(\DM_read_data<8>/FROM ),
    .O(DM_read_data[8])
  );
  X_BUF \DM_read_data<8>/YUSED  (
    .I(\DM_read_data<8>/GROM ),
    .O(DM_read_data[18])
  );
  defparam \DLX_IFinst__n0001<9>_SW0 .INIT = 16'h330F;
  X_LUT4 \DLX_IFinst__n0001<9>_SW0  (
    .ADR0(VCC),
    .ADR1(DLX_IFinst_PC[9]),
    .ADR2(DLX_IFinst__n0015[9]),
    .ADR3(DLX_IFinst__n0000),
    .O(\DLX_IFinst_NPC<9>/FROM )
  );
  defparam \DLX_IFinst__n0001<9> .INIT = 16'hA0F5;
  X_LUT4 \DLX_IFinst__n0001<9>  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_branch_address[9]),
    .ADR3(N92711),
    .O(\DLX_IFinst_NPC<9>/GROM )
  );
  X_BUF \DLX_IFinst_NPC<9>/XUSED  (
    .I(\DLX_IFinst_NPC<9>/FROM ),
    .O(N92711)
  );
  X_BUF \DLX_IFinst_NPC<9>/YUSED  (
    .I(\DLX_IFinst_NPC<9>/GROM ),
    .O(DLX_IFinst__n0001[9])
  );
  defparam \DLX_EXinst_Mshift__n0028_Sh<22>1 .INIT = 16'hBB88;
  X_LUT4 \DLX_EXinst_Mshift__n0028_Sh<22>1  (
    .ADR0(DLX_EXinst_N63016),
    .ADR1(DLX_IDinst_IR_function_field_0_1),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N63519),
    .O(\DLX_EXinst_Mshift__n0028_Sh<22>/FROM )
  );
  defparam DLX_EXinst_Ker629391.INIT = 16'hAFA0;
  X_LUT4 DLX_EXinst_Ker629391 (
    .ADR0(\DLX_EXinst_Mshift__n0024_Sh[30] ),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_IR_function_field[3]),
    .ADR3(\DLX_EXinst_Mshift__n0028_Sh[22] ),
    .O(\DLX_EXinst_Mshift__n0028_Sh<22>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0028_Sh<22>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0028_Sh<22>/FROM ),
    .O(\DLX_EXinst_Mshift__n0028_Sh[22] )
  );
  X_BUF \DLX_EXinst_Mshift__n0028_Sh<22>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0028_Sh<22>/GROM ),
    .O(DLX_EXinst_N62941)
  );
  defparam \DM_read_data<9>1 .INIT = 16'hFCCC;
  X_LUT4 \DM_read_data<9>1  (
    .ADR0(VCC),
    .ADR1(N57312),
    .ADR2(RAM_read_data[9]),
    .ADR3(vga_select_6[0]),
    .O(\DM_read_data<9>/FROM )
  );
  defparam \DM_read_data<19>1 .INIT = 16'hFCCC;
  X_LUT4 \DM_read_data<19>1  (
    .ADR0(VCC),
    .ADR1(N57312),
    .ADR2(vga_select_6[0]),
    .ADR3(RAM_read_data[19]),
    .O(\DM_read_data<9>/GROM )
  );
  X_BUF \DM_read_data<9>/XUSED  (
    .I(\DM_read_data<9>/FROM ),
    .O(DM_read_data[9])
  );
  X_BUF \DM_read_data<9>/YUSED  (
    .I(\DM_read_data<9>/GROM ),
    .O(DM_read_data[19])
  );
  defparam \DLX_EXinst__n0006<16>125_SW0 .INIT = 16'h2600;
  X_LUT4 \DLX_EXinst__n0006<16>125_SW0  (
    .ADR0(DLX_IDinst_IR_opcode_field[0]),
    .ADR1(DLX_IDinst_IR_opcode_field[1]),
    .ADR2(\DLX_IDinst_Imm[31] ),
    .ADR3(DLX_EXinst_N66105),
    .O(\N126362/GROM )
  );
  X_BUF \N126362/YUSED  (
    .I(\N126362/GROM ),
    .O(N126362)
  );
  defparam \DLX_IDinst__n0117<27>15 .INIT = 16'h2C20;
  X_LUT4 \DLX_IDinst__n0117<27>15  (
    .ADR0(DLX_IDinst_Cause_Reg[27]),
    .ADR1(DLX_IDinst_regA_index[1]),
    .ADR2(DLX_IDinst_regA_index[0]),
    .ADR3(DLX_IDinst_EPC[27]),
    .O(\CHOICE2470/FROM )
  );
  defparam \DLX_IDinst__n0117<10>15 .INIT = 16'h22C0;
  X_LUT4 \DLX_IDinst__n0117<10>15  (
    .ADR0(DLX_IDinst_EPC[10]),
    .ADR1(DLX_IDinst_regA_index[0]),
    .ADR2(DLX_IDinst_Cause_Reg[10]),
    .ADR3(DLX_IDinst_regA_index[1]),
    .O(\CHOICE2470/GROM )
  );
  X_BUF \CHOICE2470/XUSED  (
    .I(\CHOICE2470/FROM ),
    .O(CHOICE2470)
  );
  X_BUF \CHOICE2470/YUSED  (
    .I(\CHOICE2470/GROM ),
    .O(CHOICE2254)
  );
  defparam \DLX_IDinst__n0117<2>15 .INIT = 16'h3808;
  X_LUT4 \DLX_IDinst__n0117<2>15  (
    .ADR0(DLX_IDinst_EPC[2]),
    .ADR1(DLX_IDinst_regA_index[1]),
    .ADR2(DLX_IDinst_regA_index[0]),
    .ADR3(DLX_IDinst_Cause_Reg[2]),
    .O(\CHOICE2158/FROM )
  );
  defparam \DLX_IDinst__n0117<23>15 .INIT = 16'h0CA0;
  X_LUT4 \DLX_IDinst__n0117<23>15  (
    .ADR0(DLX_IDinst_Cause_Reg[23]),
    .ADR1(DLX_IDinst_EPC[23]),
    .ADR2(DLX_IDinst_regA_index[0]),
    .ADR3(DLX_IDinst_regA_index[1]),
    .O(\CHOICE2158/GROM )
  );
  X_BUF \CHOICE2158/XUSED  (
    .I(\CHOICE2158/FROM ),
    .O(CHOICE2158)
  );
  X_BUF \CHOICE2158/YUSED  (
    .I(\CHOICE2158/GROM ),
    .O(CHOICE2410)
  );
  defparam \DLX_IDinst__n0117<31>15 .INIT = 16'h0AC0;
  X_LUT4 \DLX_IDinst__n0117<31>15  (
    .ADR0(DLX_IDinst_EPC[31]),
    .ADR1(DLX_IDinst_Cause_Reg[31]),
    .ADR2(DLX_IDinst_regA_index[0]),
    .ADR3(DLX_IDinst_regA_index[1]),
    .O(\CHOICE2122/FROM )
  );
  defparam \DLX_IDinst__n0117<15>15 .INIT = 16'h0AC0;
  X_LUT4 \DLX_IDinst__n0117<15>15  (
    .ADR0(DLX_IDinst_EPC[15]),
    .ADR1(DLX_IDinst_Cause_Reg[15]),
    .ADR2(DLX_IDinst_regA_index[0]),
    .ADR3(DLX_IDinst_regA_index[1]),
    .O(\CHOICE2122/GROM )
  );
  X_BUF \CHOICE2122/XUSED  (
    .I(\CHOICE2122/FROM ),
    .O(CHOICE2122)
  );
  X_BUF \CHOICE2122/YUSED  (
    .I(\CHOICE2122/GROM ),
    .O(CHOICE2314)
  );
  defparam \DLX_EXinst_Mshift__n0028_Sh<49>1 .INIT = 16'hCCAA;
  X_LUT4 \DLX_EXinst_Mshift__n0028_Sh<49>1  (
    .ADR0(DLX_EXinst_N64854),
    .ADR1(DLX_EXinst_N63021),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_IR_function_field_2_1),
    .O(\DLX_EXinst_Mshift__n0028_Sh<49>/FROM )
  );
  defparam \DLX_EXinst__n0006<17>109_SW0 .INIT = 16'hFCCC;
  X_LUT4 \DLX_EXinst__n0006<17>109_SW0  (
    .ADR0(VCC),
    .ADR1(CHOICE5598),
    .ADR2(DLX_EXinst__n0082),
    .ADR3(\DLX_EXinst_Mshift__n0028_Sh[49] ),
    .O(\DLX_EXinst_Mshift__n0028_Sh<49>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0028_Sh<49>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0028_Sh<49>/FROM ),
    .O(\DLX_EXinst_Mshift__n0028_Sh[49] )
  );
  X_BUF \DLX_EXinst_Mshift__n0028_Sh<49>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0028_Sh<49>/GROM ),
    .O(N126631)
  );
  defparam \DLX_IDinst__n0117<19>15 .INIT = 16'h5808;
  X_LUT4 \DLX_IDinst__n0117<19>15  (
    .ADR0(DLX_IDinst_regA_index[0]),
    .ADR1(DLX_IDinst_Cause_Reg[19]),
    .ADR2(DLX_IDinst_regA_index[1]),
    .ADR3(DLX_IDinst_EPC[19]),
    .O(\CHOICE2362/FROM )
  );
  defparam \DLX_IDinst__n0117<0>15 .INIT = 16'h6240;
  X_LUT4 \DLX_IDinst__n0117<0>15  (
    .ADR0(DLX_IDinst_regA_index[1]),
    .ADR1(DLX_IDinst_regA_index[0]),
    .ADR2(DLX_IDinst_Cause_Reg[0]),
    .ADR3(DLX_IDinst_EPC[0]),
    .O(\CHOICE2362/GROM )
  );
  X_BUF \CHOICE2362/XUSED  (
    .I(\CHOICE2362/FROM ),
    .O(CHOICE2362)
  );
  X_BUF \CHOICE2362/YUSED  (
    .I(\CHOICE2362/GROM ),
    .O(CHOICE2146)
  );
  defparam \DLX_IDinst__n0117<23>29 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst__n0117<23>29  (
    .ADR0(CHOICE2410),
    .ADR1(N101161),
    .ADR2(DLX_IDinst_regA_eff[23]),
    .ADR3(DLX_IDinst_N69914),
    .O(\DLX_IDinst_reg_out_A<23>/FROM )
  );
  defparam \DLX_IDinst__n0117<23>39 .INIT = 16'hFF88;
  X_LUT4 \DLX_IDinst__n0117<23>39  (
    .ADR0(DLX_IDinst__n0310),
    .ADR1(DLX_IFinst_NPC[23]),
    .ADR2(VCC),
    .ADR3(CHOICE2413),
    .O(N104236)
  );
  X_BUF \DLX_IDinst_reg_out_A<23>/XUSED  (
    .I(\DLX_IDinst_reg_out_A<23>/FROM ),
    .O(CHOICE2413)
  );
  defparam \DLX_IDinst__n0117<31>29 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst__n0117<31>29  (
    .ADR0(DLX_IDinst_regA_eff[31]),
    .ADR1(DLX_IDinst_N69914),
    .ADR2(CHOICE2122),
    .ADR3(N101161),
    .O(\DLX_IDinst_reg_out_A<31>/FROM )
  );
  defparam \DLX_IDinst__n0117<31>39 .INIT = 16'hFFC0;
  X_LUT4 \DLX_IDinst__n0117<31>39  (
    .ADR0(VCC),
    .ADR1(DLX_IFinst_NPC[31]),
    .ADR2(DLX_IDinst__n0310),
    .ADR3(CHOICE2125),
    .O(N102604)
  );
  X_BUF \DLX_IDinst_reg_out_A<31>/XUSED  (
    .I(\DLX_IDinst_reg_out_A<31>/FROM ),
    .O(CHOICE2125)
  );
  defparam \DLX_IDinst__n0117<15>29 .INIT = 16'hEAC0;
  X_LUT4 \DLX_IDinst__n0117<15>29  (
    .ADR0(DLX_IDinst_regA_eff[15]),
    .ADR1(CHOICE2314),
    .ADR2(N101161),
    .ADR3(DLX_IDinst_N69914),
    .O(\DLX_IDinst_reg_out_A<15>/FROM )
  );
  defparam \DLX_IDinst__n0117<15>39 .INIT = 16'hFFA0;
  X_LUT4 \DLX_IDinst__n0117<15>39  (
    .ADR0(DLX_IFinst_NPC[15]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst__n0310),
    .ADR3(CHOICE2317),
    .O(N103692)
  );
  X_BUF \DLX_IDinst_reg_out_A<15>/XUSED  (
    .I(\DLX_IDinst_reg_out_A<15>/FROM ),
    .O(CHOICE2317)
  );
  defparam \DLX_IDinst__n0117<0>29 .INIT = 16'hEAC0;
  X_LUT4 \DLX_IDinst__n0117<0>29  (
    .ADR0(CHOICE2146),
    .ADR1(DLX_IDinst_N69914),
    .ADR2(DLX_IDinst_regA_eff[0]),
    .ADR3(N101161),
    .O(\DLX_IDinst_reg_out_A<0>/FROM )
  );
  defparam \DLX_IDinst__n0117<0>39 .INIT = 16'hFFC0;
  X_LUT4 \DLX_IDinst__n0117<0>39  (
    .ADR0(VCC),
    .ADR1(DLX_IFinst_NPC[0]),
    .ADR2(DLX_IDinst__n0310),
    .ADR3(CHOICE2149),
    .O(N102740)
  );
  X_BUF \DLX_IDinst_reg_out_A<0>/XUSED  (
    .I(\DLX_IDinst_reg_out_A<0>/FROM ),
    .O(CHOICE2149)
  );
  defparam \DLX_IDinst__n0117<18>15 .INIT = 16'h5088;
  X_LUT4 \DLX_IDinst__n0117<18>15  (
    .ADR0(DLX_IDinst_regA_index[1]),
    .ADR1(DLX_IDinst_EPC[18]),
    .ADR2(DLX_IDinst_Cause_Reg[18]),
    .ADR3(DLX_IDinst_regA_index[0]),
    .O(\CHOICE2350/FROM )
  );
  defparam \DLX_IDinst__n0117<24>15 .INIT = 16'h44A0;
  X_LUT4 \DLX_IDinst__n0117<24>15  (
    .ADR0(DLX_IDinst_regA_index[1]),
    .ADR1(DLX_IDinst_Cause_Reg[24]),
    .ADR2(DLX_IDinst_EPC[24]),
    .ADR3(DLX_IDinst_regA_index[0]),
    .O(\CHOICE2350/GROM )
  );
  X_BUF \CHOICE2350/XUSED  (
    .I(\CHOICE2350/FROM ),
    .O(CHOICE2350)
  );
  X_BUF \CHOICE2350/YUSED  (
    .I(\CHOICE2350/GROM ),
    .O(CHOICE2434)
  );
  defparam \DLX_IDinst__n0117<28>15 .INIT = 16'h3808;
  X_LUT4 \DLX_IDinst__n0117<28>15  (
    .ADR0(DLX_IDinst_Cause_Reg[28]),
    .ADR1(DLX_IDinst_regA_index[0]),
    .ADR2(DLX_IDinst_regA_index[1]),
    .ADR3(DLX_IDinst_EPC[28]),
    .O(\CHOICE2458/FROM )
  );
  defparam \DLX_IDinst__n0117<1>15 .INIT = 16'h6420;
  X_LUT4 \DLX_IDinst__n0117<1>15  (
    .ADR0(DLX_IDinst_regA_index[1]),
    .ADR1(DLX_IDinst_regA_index[0]),
    .ADR2(DLX_IDinst_EPC[1]),
    .ADR3(DLX_IDinst_Cause_Reg[1]),
    .O(\CHOICE2458/GROM )
  );
  X_BUF \CHOICE2458/XUSED  (
    .I(\CHOICE2458/FROM ),
    .O(CHOICE2458)
  );
  X_BUF \CHOICE2458/YUSED  (
    .I(\CHOICE2458/GROM ),
    .O(CHOICE2134)
  );
  defparam \DLX_IDinst__n0117<24>29 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst__n0117<24>29  (
    .ADR0(DLX_IDinst_regA_eff[24]),
    .ADR1(DLX_IDinst_N69914),
    .ADR2(CHOICE2434),
    .ADR3(N101161),
    .O(\DLX_IDinst_reg_out_A<24>/FROM )
  );
  defparam \DLX_IDinst__n0117<24>39 .INIT = 16'hFFA0;
  X_LUT4 \DLX_IDinst__n0117<24>39  (
    .ADR0(DLX_IFinst_NPC[24]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst__n0310),
    .ADR3(CHOICE2437),
    .O(N104372)
  );
  X_BUF \DLX_IDinst_reg_out_A<24>/XUSED  (
    .I(\DLX_IDinst_reg_out_A<24>/FROM ),
    .O(CHOICE2437)
  );
  defparam \DLX_IDinst__n0117<16>29 .INIT = 16'hECA0;
  X_LUT4 \DLX_IDinst__n0117<16>29  (
    .ADR0(CHOICE2338),
    .ADR1(DLX_IDinst_regA_eff[16]),
    .ADR2(N101161),
    .ADR3(DLX_IDinst_N69914),
    .O(\DLX_IDinst_reg_out_A<16>/FROM )
  );
  defparam \DLX_IDinst__n0117<16>39 .INIT = 16'hFFA0;
  X_LUT4 \DLX_IDinst__n0117<16>39  (
    .ADR0(DLX_IDinst__n0310),
    .ADR1(VCC),
    .ADR2(DLX_IFinst_NPC[16]),
    .ADR3(CHOICE2341),
    .O(N103828)
  );
  X_BUF \DLX_IDinst_reg_out_A<16>/XUSED  (
    .I(\DLX_IDinst_reg_out_A<16>/FROM ),
    .O(CHOICE2341)
  );
  defparam DLX_IDinst_Ker6997925.INIT = 16'h00CC;
  X_LUT4 DLX_IDinst_Ker6997925 (
    .ADR0(VCC),
    .ADR1(DLX_opcode_of_MEM[5]),
    .ADR2(VCC),
    .ADR3(DLX_opcode_of_MEM[4]),
    .O(\CHOICE1459/FROM )
  );
  defparam DLX_IDinst_Ker6997930.INIT = 16'h2F00;
  X_LUT4 DLX_IDinst_Ker6997930 (
    .ADR0(DLX_opcode_of_MEM[0]),
    .ADR1(DLX_opcode_of_MEM[2]),
    .ADR2(DLX_opcode_of_MEM[1]),
    .ADR3(CHOICE1459),
    .O(\CHOICE1459/GROM )
  );
  X_BUF \CHOICE1459/XUSED  (
    .I(\CHOICE1459/FROM ),
    .O(CHOICE1459)
  );
  X_BUF \CHOICE1459/YUSED  (
    .I(\CHOICE1459/GROM ),
    .O(CHOICE1460)
  );
  defparam \DLX_IDinst__n0117<1>29 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst__n0117<1>29  (
    .ADR0(CHOICE2134),
    .ADR1(N101161),
    .ADR2(DLX_IDinst_N69914),
    .ADR3(DLX_IDinst_regA_eff[1]),
    .O(\DLX_IDinst_reg_out_A<1>/FROM )
  );
  defparam \DLX_IDinst__n0117<1>39 .INIT = 16'hFFC0;
  X_LUT4 \DLX_IDinst__n0117<1>39  (
    .ADR0(VCC),
    .ADR1(DLX_IFinst_NPC[1]),
    .ADR2(DLX_IDinst__n0310),
    .ADR3(CHOICE2137),
    .O(N102672)
  );
  X_BUF \DLX_IDinst_reg_out_A<1>/XUSED  (
    .I(\DLX_IDinst_reg_out_A<1>/FROM ),
    .O(CHOICE2137)
  );
  defparam \DLX_EXinst_Mshift__n0025_Sh<45>_SW0 .INIT = 16'h0C3F;
  X_LUT4 \DLX_EXinst_Mshift__n0025_Sh<45>_SW0  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_B_2_1),
    .ADR2(\DLX_EXinst_Mshift__n0025_Sh[9] ),
    .ADR3(\DLX_EXinst_Mshift__n0025_Sh[13] ),
    .O(\N93641/FROM )
  );
  defparam \DLX_EXinst__n0006<13>176 .INIT = 16'hC044;
  X_LUT4 \DLX_EXinst__n0006<13>176  (
    .ADR0(N93641),
    .ADR1(DLX_EXinst_N66535),
    .ADR2(DLX_EXinst_N62906),
    .ADR3(DLX_IDinst_reg_out_B[3]),
    .O(\N93641/GROM )
  );
  X_BUF \N93641/XUSED  (
    .I(\N93641/FROM ),
    .O(N93641)
  );
  X_BUF \N93641/YUSED  (
    .I(\N93641/GROM ),
    .O(CHOICE4336)
  );
  defparam \DLX_IDinst__n0117<17>29 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst__n0117<17>29  (
    .ADR0(N101161),
    .ADR1(CHOICE2326),
    .ADR2(DLX_IDinst_N69914),
    .ADR3(DLX_IDinst_regA_eff[17]),
    .O(\DLX_IDinst_reg_out_A<17>/FROM )
  );
  defparam \DLX_IDinst__n0117<17>39 .INIT = 16'hFF88;
  X_LUT4 \DLX_IDinst__n0117<17>39  (
    .ADR0(DLX_IDinst__n0310),
    .ADR1(DLX_IFinst_NPC[17]),
    .ADR2(VCC),
    .ADR3(CHOICE2329),
    .O(N103760)
  );
  X_BUF \DLX_IDinst_reg_out_A<17>/XUSED  (
    .I(\DLX_IDinst_reg_out_A<17>/FROM ),
    .O(CHOICE2329)
  );
  defparam \DLX_IDinst__n0117<25>29 .INIT = 16'hECA0;
  X_LUT4 \DLX_IDinst__n0117<25>29  (
    .ADR0(DLX_IDinst_N69914),
    .ADR1(CHOICE2422),
    .ADR2(DLX_IDinst_regA_eff[25]),
    .ADR3(N101161),
    .O(\DLX_IDinst_reg_out_A<25>/FROM )
  );
  defparam \DLX_IDinst__n0117<25>39 .INIT = 16'hFFC0;
  X_LUT4 \DLX_IDinst__n0117<25>39  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst__n0310),
    .ADR2(DLX_IFinst_NPC[25]),
    .ADR3(CHOICE2425),
    .O(N104304)
  );
  X_BUF \DLX_IDinst_reg_out_A<25>/XUSED  (
    .I(\DLX_IDinst_reg_out_A<25>/FROM ),
    .O(CHOICE2425)
  );
  defparam \DLX_IDinst__n0117<2>29 .INIT = 16'hEAC0;
  X_LUT4 \DLX_IDinst__n0117<2>29  (
    .ADR0(DLX_IDinst_N69914),
    .ADR1(CHOICE2158),
    .ADR2(N101161),
    .ADR3(DLX_IDinst_regA_eff[2]),
    .O(\DLX_IDinst_reg_out_A<2>/FROM )
  );
  defparam \DLX_IDinst__n0117<2>39 .INIT = 16'hFFA0;
  X_LUT4 \DLX_IDinst__n0117<2>39  (
    .ADR0(DLX_IDinst__n0310),
    .ADR1(VCC),
    .ADR2(DLX_IFinst_NPC[2]),
    .ADR3(CHOICE2161),
    .O(N102808)
  );
  X_BUF \DLX_IDinst_reg_out_A<2>/XUSED  (
    .I(\DLX_IDinst_reg_out_A<2>/FROM ),
    .O(CHOICE2161)
  );
  defparam DLX_IDinst_Ker69979112.INIT = 16'h0E0A;
  X_LUT4 DLX_IDinst_Ker69979112 (
    .ADR0(CHOICE1479),
    .ADR1(DLX_opcode_of_MEM[3]),
    .ADR2(DLX_opcode_of_MEM[5]),
    .ADR3(CHOICE1471),
    .O(\CHOICE1481/FROM )
  );
  defparam DLX_IDinst_Ker69979126.INIT = 16'hFF32;
  X_LUT4 DLX_IDinst_Ker69979126 (
    .ADR0(CHOICE1460),
    .ADR1(DLX_opcode_of_MEM[3]),
    .ADR2(CHOICE1453),
    .ADR3(CHOICE1481),
    .O(\CHOICE1481/GROM )
  );
  X_BUF \CHOICE1481/XUSED  (
    .I(\CHOICE1481/FROM ),
    .O(CHOICE1481)
  );
  X_BUF \CHOICE1481/YUSED  (
    .I(\CHOICE1481/GROM ),
    .O(N98806)
  );
  defparam DLX_IDinst_Ker6997977.INIT = 16'h5F7F;
  X_LUT4 DLX_IDinst_Ker6997977 (
    .ADR0(DLX_opcode_of_MEM[2]),
    .ADR1(DLX_opcode_of_MEM[1]),
    .ADR2(DLX_opcode_of_MEM[4]),
    .ADR3(DLX_opcode_of_MEM[0]),
    .O(\CHOICE1471/GROM )
  );
  X_BUF \CHOICE1471/YUSED  (
    .I(\CHOICE1471/GROM ),
    .O(CHOICE1471)
  );
  defparam \DLX_IDinst__n0117<26>29 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst__n0117<26>29  (
    .ADR0(N101161),
    .ADR1(CHOICE2446),
    .ADR2(DLX_IDinst_regA_eff[26]),
    .ADR3(DLX_IDinst_N69914),
    .O(\DLX_IDinst_reg_out_A<26>/FROM )
  );
  defparam \DLX_IDinst__n0117<26>39 .INIT = 16'hFFA0;
  X_LUT4 \DLX_IDinst__n0117<26>39  (
    .ADR0(DLX_IDinst__n0310),
    .ADR1(VCC),
    .ADR2(DLX_IFinst_NPC[26]),
    .ADR3(CHOICE2449),
    .O(N104440)
  );
  X_BUF \DLX_IDinst_reg_out_A<26>/XUSED  (
    .I(\DLX_IDinst_reg_out_A<26>/FROM ),
    .O(CHOICE2449)
  );
  defparam \DLX_IDinst__n0117<18>29 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst__n0117<18>29  (
    .ADR0(DLX_IDinst_regA_eff[18]),
    .ADR1(DLX_IDinst_N69914),
    .ADR2(CHOICE2350),
    .ADR3(N101161),
    .O(\DLX_IDinst_reg_out_A<18>/FROM )
  );
  defparam \DLX_IDinst__n0117<18>39 .INIT = 16'hFF88;
  X_LUT4 \DLX_IDinst__n0117<18>39  (
    .ADR0(DLX_IFinst_NPC[18]),
    .ADR1(DLX_IDinst__n0310),
    .ADR2(VCC),
    .ADR3(CHOICE2353),
    .O(N103896)
  );
  X_BUF \DLX_IDinst_reg_out_A<18>/XUSED  (
    .I(\DLX_IDinst_reg_out_A<18>/FROM ),
    .O(CHOICE2353)
  );
  defparam \DLX_IDinst__n0117<3>29 .INIT = 16'hECA0;
  X_LUT4 \DLX_IDinst__n0117<3>29  (
    .ADR0(DLX_IDinst_regA_eff[3]),
    .ADR1(N101161),
    .ADR2(DLX_IDinst_N69914),
    .ADR3(CHOICE2182),
    .O(\DLX_IDinst_reg_out_A<3>/FROM )
  );
  defparam \DLX_IDinst__n0117<3>39 .INIT = 16'hFFA0;
  X_LUT4 \DLX_IDinst__n0117<3>39  (
    .ADR0(DLX_IFinst_NPC[3]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst__n0310),
    .ADR3(CHOICE2185),
    .O(N102944)
  );
  X_BUF \DLX_IDinst_reg_out_A<3>/XUSED  (
    .I(\DLX_IDinst_reg_out_A<3>/FROM ),
    .O(CHOICE2185)
  );
  defparam \DLX_IDinst__n0117<27>29 .INIT = 16'hECA0;
  X_LUT4 \DLX_IDinst__n0117<27>29  (
    .ADR0(DLX_IDinst_regA_eff[27]),
    .ADR1(CHOICE2470),
    .ADR2(DLX_IDinst_N69914),
    .ADR3(N101161),
    .O(\DLX_IDinst_reg_out_A<27>/FROM )
  );
  defparam \DLX_IDinst__n0117<27>39 .INIT = 16'hFF88;
  X_LUT4 \DLX_IDinst__n0117<27>39  (
    .ADR0(DLX_IDinst__n0310),
    .ADR1(DLX_IFinst_NPC[27]),
    .ADR2(VCC),
    .ADR3(CHOICE2473),
    .O(N104576)
  );
  X_BUF \DLX_IDinst_reg_out_A<27>/XUSED  (
    .I(\DLX_IDinst_reg_out_A<27>/FROM ),
    .O(CHOICE2473)
  );
  defparam \DLX_IDinst__n0117<19>29 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst__n0117<19>29  (
    .ADR0(DLX_IDinst_regA_eff[19]),
    .ADR1(DLX_IDinst_N69914),
    .ADR2(CHOICE2362),
    .ADR3(N101161),
    .O(\DLX_IDinst_reg_out_A<19>/FROM )
  );
  defparam \DLX_IDinst__n0117<19>39 .INIT = 16'hFFA0;
  X_LUT4 \DLX_IDinst__n0117<19>39  (
    .ADR0(DLX_IFinst_NPC[19]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst__n0310),
    .ADR3(CHOICE2365),
    .O(N103964)
  );
  X_BUF \DLX_IDinst_reg_out_A<19>/XUSED  (
    .I(\DLX_IDinst_reg_out_A<19>/FROM ),
    .O(CHOICE2365)
  );
  defparam \DLX_IDinst__n0117<4>29 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst__n0117<4>29  (
    .ADR0(DLX_IDinst_regA_eff[4]),
    .ADR1(DLX_IDinst_N69914),
    .ADR2(CHOICE2170),
    .ADR3(N101161),
    .O(\DLX_IDinst_reg_out_A<4>/FROM )
  );
  defparam \DLX_IDinst__n0117<4>39 .INIT = 16'hFFC0;
  X_LUT4 \DLX_IDinst__n0117<4>39  (
    .ADR0(VCC),
    .ADR1(DLX_IFinst_NPC[4]),
    .ADR2(DLX_IDinst__n0310),
    .ADR3(CHOICE2173),
    .O(N102876)
  );
  X_BUF \DLX_IDinst_reg_out_A<4>/XUSED  (
    .I(\DLX_IDinst_reg_out_A<4>/FROM ),
    .O(CHOICE2173)
  );
  defparam DLX_IDinst__n0410_SW0.INIT = 16'hEEEE;
  X_LUT4 DLX_IDinst__n0410_SW0 (
    .ADR0(DLX_MEMinst_reg_dst_out[3]),
    .ADR1(DLX_MEMinst_reg_dst_out[2]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\N90186/FROM )
  );
  defparam DLX_IDinst__n0410_1184.INIT = 16'hFFFE;
  X_LUT4 DLX_IDinst__n0410_1184 (
    .ADR0(DLX_MEMinst_reg_dst_out[0]),
    .ADR1(DLX_MEMinst_reg_dst_out[4]),
    .ADR2(DLX_MEMinst_reg_dst_out[1]),
    .ADR3(N90186),
    .O(\N90186/GROM )
  );
  X_BUF \N90186/XUSED  (
    .I(\N90186/FROM ),
    .O(N90186)
  );
  X_BUF \N90186/YUSED  (
    .I(\N90186/GROM ),
    .O(DLX_IDinst__n0410)
  );
  defparam DLX_IFinst_IR_latched_10.INIT = 1'b0;
  X_FF DLX_IFinst_IR_latched_10 (
    .I(DLX_IFinst__n0003[10]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_IR_latched<10>/FFX/RST ),
    .O(DLX_IFinst_IR_latched[10])
  );
  X_OR2 \DLX_IFinst_IR_latched<10>/FFX/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IFinst_IR_latched<10>/FFX/RST )
  );
  defparam DLX_IFinst_IR_latched_11.INIT = 1'b0;
  X_FF DLX_IFinst_IR_latched_11 (
    .I(DLX_IFinst__n0003[11]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_IR_latched<11>/FFX/RST ),
    .O(DLX_IFinst_IR_latched[11])
  );
  X_OR2 \DLX_IFinst_IR_latched<11>/FFX/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IFinst_IR_latched<11>/FFX/RST )
  );
  defparam DLX_IFinst_IR_latched_12.INIT = 1'b0;
  X_FF DLX_IFinst_IR_latched_12 (
    .I(DLX_IFinst__n0003[12]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_IR_latched<12>/FFX/RST ),
    .O(DLX_IFinst_IR_latched[12])
  );
  X_OR2 \DLX_IFinst_IR_latched<12>/FFX/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IFinst_IR_latched<12>/FFX/RST )
  );
  defparam DLX_IFinst_IR_latched_20.INIT = 1'b0;
  X_FF DLX_IFinst_IR_latched_20 (
    .I(DLX_IFinst__n0003[20]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_IR_latched<20>/FFX/RST ),
    .O(DLX_IFinst_IR_latched[20])
  );
  X_OR2 \DLX_IFinst_IR_latched<20>/FFX/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IFinst_IR_latched<20>/FFX/RST )
  );
  defparam DLX_IFinst_IR_latched_13.INIT = 1'b0;
  X_FF DLX_IFinst_IR_latched_13 (
    .I(DLX_IFinst__n0003[13]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_IR_latched<13>/FFX/RST ),
    .O(DLX_IFinst_IR_latched[13])
  );
  X_OR2 \DLX_IFinst_IR_latched<13>/FFX/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IFinst_IR_latched<13>/FFX/RST )
  );
  defparam DLX_IFinst_IR_latched_21.INIT = 1'b0;
  X_FF DLX_IFinst_IR_latched_21 (
    .I(DLX_IFinst__n0003[21]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_IR_latched<21>/FFX/RST ),
    .O(DLX_IFinst_IR_latched[21])
  );
  X_OR2 \DLX_IFinst_IR_latched<21>/FFX/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IFinst_IR_latched<21>/FFX/RST )
  );
  defparam DLX_IFinst_IR_latched_14.INIT = 1'b0;
  X_FF DLX_IFinst_IR_latched_14 (
    .I(DLX_IFinst__n0003[14]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_IR_latched<14>/FFX/RST ),
    .O(DLX_IFinst_IR_latched[14])
  );
  X_OR2 \DLX_IFinst_IR_latched<14>/FFX/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IFinst_IR_latched<14>/FFX/RST )
  );
  defparam DLX_MEMinst_RF_data_in_11.INIT = 1'b0;
  X_FF DLX_MEMinst_RF_data_in_11 (
    .I(DLX_MEMinst__n0000[11]),
    .CE(VCC),
    .CLK(\DLX_MEMinst_RF_data_in<11>/CKMUXNOT ),
    .SET(GND),
    .RST(\DLX_MEMinst_RF_data_in<11>/FFX/RST ),
    .O(DLX_MEMinst_RF_data_in[11])
  );
  X_OR2 \DLX_MEMinst_RF_data_in<11>/FFX/RSTOR  (
    .I0(reset_IBUF_1),
    .I1(GSR),
    .O(\DLX_MEMinst_RF_data_in<11>/FFX/RST )
  );
  defparam DLX_MEMinst_RF_data_in_21.INIT = 1'b0;
  X_FF DLX_MEMinst_RF_data_in_21 (
    .I(DLX_MEMinst__n0000[21]),
    .CE(VCC),
    .CLK(\DLX_MEMinst_RF_data_in<21>/CKMUXNOT ),
    .SET(GND),
    .RST(\DLX_MEMinst_RF_data_in<21>/FFX/RST ),
    .O(DLX_MEMinst_RF_data_in[21])
  );
  X_OR2 \DLX_MEMinst_RF_data_in<21>/FFX/RSTOR  (
    .I0(reset_IBUF_1),
    .I1(GSR),
    .O(\DLX_MEMinst_RF_data_in<21>/FFX/RST )
  );
  defparam DLX_MEMinst_RF_data_in_13.INIT = 1'b0;
  X_FF DLX_MEMinst_RF_data_in_13 (
    .I(DLX_MEMinst__n0000[13]),
    .CE(VCC),
    .CLK(\DLX_MEMinst_RF_data_in<13>/CKMUXNOT ),
    .SET(GND),
    .RST(\DLX_MEMinst_RF_data_in<13>/FFX/RST ),
    .O(DLX_MEMinst_RF_data_in[13])
  );
  X_OR2 \DLX_MEMinst_RF_data_in<13>/FFX/RSTOR  (
    .I0(reset_IBUF_1),
    .I1(GSR),
    .O(\DLX_MEMinst_RF_data_in<13>/FFX/RST )
  );
  defparam DLX_MEMinst_RF_data_in_31.INIT = 1'b0;
  X_FF DLX_MEMinst_RF_data_in_31 (
    .I(DLX_MEMinst__n0000[31]),
    .CE(VCC),
    .CLK(\DLX_MEMinst_RF_data_in<31>/CKMUXNOT ),
    .SET(GND),
    .RST(\DLX_MEMinst_RF_data_in<31>/FFX/RST ),
    .O(DLX_MEMinst_RF_data_in[31])
  );
  X_OR2 \DLX_MEMinst_RF_data_in<31>/FFX/RSTOR  (
    .I0(reset_IBUF_1),
    .I1(GSR),
    .O(\DLX_MEMinst_RF_data_in<31>/FFX/RST )
  );
  defparam DLX_MEMinst_RF_data_in_23.INIT = 1'b0;
  X_FF DLX_MEMinst_RF_data_in_23 (
    .I(DLX_MEMinst__n0000[23]),
    .CE(VCC),
    .CLK(\DLX_MEMinst_RF_data_in<23>/CKMUXNOT ),
    .SET(GND),
    .RST(\DLX_MEMinst_RF_data_in<23>/FFX/RST ),
    .O(DLX_MEMinst_RF_data_in[23])
  );
  X_OR2 \DLX_MEMinst_RF_data_in<23>/FFX/RSTOR  (
    .I0(reset_IBUF_1),
    .I1(GSR),
    .O(\DLX_MEMinst_RF_data_in<23>/FFX/RST )
  );
  defparam DLX_EXinst_reg_dst_out_4.INIT = 1'b0;
  X_FF DLX_EXinst_reg_dst_out_4 (
    .I(DLX_EXinst__n0008[4]),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_reg_dst_out<4>/FFY/RST ),
    .O(DLX_EXinst_reg_dst_out[4])
  );
  X_OR2 \DLX_EXinst_reg_dst_out<4>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_reg_dst_out<4>/FFY/RST )
  );
  defparam DLX_IDinst_reg_out_B_11.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_B_11 (
    .I(DLX_IDinst__n0118[11]),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_B<11>/FFX/RST ),
    .O(DLX_IDinst_reg_out_B[11])
  );
  X_OR2 \DLX_IDinst_reg_out_B<11>/FFX/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_B<11>/FFX/RST )
  );
  defparam DLX_IDinst_reg_out_B_21.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_B_21 (
    .I(DLX_IDinst__n0118[21]),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_B<21>/FFX/RST ),
    .O(DLX_IDinst_reg_out_B[21])
  );
  X_OR2 \DLX_IDinst_reg_out_B<21>/FFX/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_B<21>/FFX/RST )
  );
  defparam DLX_IDinst_reg_out_B_12.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_B_12 (
    .I(DLX_IDinst__n0118[12]),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_B<13>/FFY/RST ),
    .O(DLX_IDinst_reg_out_B[12])
  );
  X_OR2 \DLX_IDinst_reg_out_B<13>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_B<13>/FFY/RST )
  );
  defparam DLX_IDinst_reg_out_B_13.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_B_13 (
    .I(DLX_IDinst__n0118[13]),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_B<13>/FFX/RST ),
    .O(DLX_IDinst_reg_out_B[13])
  );
  X_OR2 \DLX_IDinst_reg_out_B<13>/FFX/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_B<13>/FFX/RST )
  );
  defparam DLX_IDinst_reg_out_B_30.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_B_30 (
    .I(DLX_IDinst__n0118[30]),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_B<31>/FFY/RST ),
    .O(DLX_IDinst_reg_out_B[30])
  );
  X_OR2 \DLX_IDinst_reg_out_B<31>/FFY/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_B<31>/FFY/RST )
  );
  defparam DLX_IDinst_reg_out_B_31.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_B_31 (
    .I(DLX_IDinst__n0118[31]),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_B<31>/FFX/RST ),
    .O(DLX_IDinst_reg_out_B[31])
  );
  X_OR2 \DLX_IDinst_reg_out_B<31>/FFX/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_B<31>/FFX/RST )
  );
  defparam DLX_IDinst_reg_out_B_22.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_B_22 (
    .I(DLX_IDinst__n0118[22]),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_B<23>/FFY/RST ),
    .O(DLX_IDinst_reg_out_B[22])
  );
  X_OR2 \DLX_IDinst_reg_out_B<23>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_B<23>/FFY/RST )
  );
  defparam DLX_IDinst_reg_out_B_23.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_B_23 (
    .I(DLX_IDinst__n0118[23]),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_B<23>/FFX/RST ),
    .O(DLX_IDinst_reg_out_B[23])
  );
  X_OR2 \DLX_IDinst_reg_out_B<23>/FFX/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_B<23>/FFX/RST )
  );
  defparam DLX_IDinst_reg_out_B_14.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_B_14 (
    .I(DLX_IDinst__n0118[14]),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_B<15>/FFY/RST ),
    .O(DLX_IDinst_reg_out_B[14])
  );
  X_OR2 \DLX_IDinst_reg_out_B<15>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_B<15>/FFY/RST )
  );
  defparam DLX_IFinst_IR_latched_0.INIT = 1'b0;
  X_FF DLX_IFinst_IR_latched_0 (
    .I(DLX_IFinst__n0003[0]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_IR_latched<0>/FFX/RST ),
    .O(DLX_IFinst_IR_latched[0])
  );
  X_OR2 \DLX_IFinst_IR_latched<0>/FFX/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IFinst_IR_latched<0>/FFX/RST )
  );
  defparam DLX_IFinst_IR_latched_1.INIT = 1'b0;
  X_FF DLX_IFinst_IR_latched_1 (
    .I(DLX_IFinst__n0003[1]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_IR_latched<1>/FFX/RST ),
    .O(DLX_IFinst_IR_latched[1])
  );
  X_OR2 \DLX_IFinst_IR_latched<1>/FFX/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IFinst_IR_latched<1>/FFX/RST )
  );
  defparam DLX_IFinst_IR_latched_2.INIT = 1'b0;
  X_FF DLX_IFinst_IR_latched_2 (
    .I(DLX_IFinst__n0003[2]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_IR_latched<2>/FFX/RST ),
    .O(DLX_IFinst_IR_latched[2])
  );
  X_OR2 \DLX_IFinst_IR_latched<2>/FFX/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IFinst_IR_latched<2>/FFX/RST )
  );
  defparam DLX_IFinst_IR_latched_3.INIT = 1'b0;
  X_FF DLX_IFinst_IR_latched_3 (
    .I(DLX_IFinst__n0003[3]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_IR_latched<3>/FFX/RST ),
    .O(DLX_IFinst_IR_latched[3])
  );
  X_OR2 \DLX_IFinst_IR_latched<3>/FFX/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IFinst_IR_latched<3>/FFX/RST )
  );
  defparam DLX_IFinst_IR_latched_4.INIT = 1'b0;
  X_FF DLX_IFinst_IR_latched_4 (
    .I(DLX_IFinst__n0003[4]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_IR_latched<4>/FFX/RST ),
    .O(DLX_IFinst_IR_latched[4])
  );
  X_OR2 \DLX_IFinst_IR_latched<4>/FFX/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IFinst_IR_latched<4>/FFX/RST )
  );
  defparam DLX_IFinst_IR_latched_5.INIT = 1'b0;
  X_FF DLX_IFinst_IR_latched_5 (
    .I(DLX_IFinst__n0003[5]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_IR_latched<5>/FFX/RST ),
    .O(DLX_IFinst_IR_latched[5])
  );
  X_OR2 \DLX_IFinst_IR_latched<5>/FFX/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IFinst_IR_latched<5>/FFX/RST )
  );
  defparam DLX_IFinst_IR_latched_6.INIT = 1'b0;
  X_FF DLX_IFinst_IR_latched_6 (
    .I(DLX_IFinst__n0003[6]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_IR_latched<6>/FFX/RST ),
    .O(DLX_IFinst_IR_latched[6])
  );
  X_OR2 \DLX_IFinst_IR_latched<6>/FFX/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IFinst_IR_latched<6>/FFX/RST )
  );
  defparam DLX_IFinst_IR_latched_30.INIT = 1'b0;
  X_FF DLX_IFinst_IR_latched_30 (
    .I(DLX_IFinst__n0003[30]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_IR_latched<30>/FFX/RST ),
    .O(DLX_IFinst_IR_latched[30])
  );
  X_OR2 \DLX_IFinst_IR_latched<30>/FFX/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IFinst_IR_latched<30>/FFX/RST )
  );
  defparam DLX_IFinst_IR_latched_22.INIT = 1'b0;
  X_FF DLX_IFinst_IR_latched_22 (
    .I(DLX_IFinst__n0003[22]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_IR_latched<22>/FFX/RST ),
    .O(DLX_IFinst_IR_latched[22])
  );
  X_OR2 \DLX_IFinst_IR_latched<22>/FFX/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IFinst_IR_latched<22>/FFX/RST )
  );
  defparam DLX_IFinst_IR_latched_23.INIT = 1'b0;
  X_FF DLX_IFinst_IR_latched_23 (
    .I(DLX_IFinst__n0003[23]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_IR_latched<23>/FFX/RST ),
    .O(DLX_IFinst_IR_latched[23])
  );
  X_OR2 \DLX_IFinst_IR_latched<23>/FFX/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IFinst_IR_latched<23>/FFX/RST )
  );
  defparam DLX_IFinst_IR_latched_31.INIT = 1'b0;
  X_FF DLX_IFinst_IR_latched_31 (
    .I(DLX_IFinst__n0003[31]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_IR_latched<31>/FFX/RST ),
    .O(DLX_IFinst_IR_latched[31])
  );
  X_OR2 \DLX_IFinst_IR_latched<31>/FFX/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IFinst_IR_latched<31>/FFX/RST )
  );
  defparam DLX_IFinst_IR_latched_15.INIT = 1'b0;
  X_FF DLX_IFinst_IR_latched_15 (
    .I(DLX_IFinst__n0003[15]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_IR_latched<15>/FFX/RST ),
    .O(DLX_IFinst_IR_latched[15])
  );
  X_OR2 \DLX_IFinst_IR_latched<15>/FFX/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IFinst_IR_latched<15>/FFX/RST )
  );
  defparam DLX_IFinst_IR_latched_16.INIT = 1'b0;
  X_FF DLX_IFinst_IR_latched_16 (
    .I(DLX_IFinst__n0003[16]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_IR_latched<16>/FFX/RST ),
    .O(DLX_IFinst_IR_latched[16])
  );
  X_OR2 \DLX_IFinst_IR_latched<16>/FFX/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IFinst_IR_latched<16>/FFX/RST )
  );
  defparam DLX_IFinst_IR_latched_24.INIT = 1'b0;
  X_FF DLX_IFinst_IR_latched_24 (
    .I(DLX_IFinst__n0003[24]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_IR_latched<24>/FFX/RST ),
    .O(DLX_IFinst_IR_latched[24])
  );
  X_OR2 \DLX_IFinst_IR_latched<24>/FFX/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IFinst_IR_latched<24>/FFX/RST )
  );
  defparam DLX_IFinst_IR_latched_25.INIT = 1'b0;
  X_FF DLX_IFinst_IR_latched_25 (
    .I(DLX_IFinst__n0003[25]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_IR_latched<25>/FFX/RST ),
    .O(DLX_IFinst_IR_latched[25])
  );
  X_OR2 \DLX_IFinst_IR_latched<25>/FFX/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IFinst_IR_latched<25>/FFX/RST )
  );
  defparam DLX_IFinst_IR_latched_17.INIT = 1'b0;
  X_FF DLX_IFinst_IR_latched_17 (
    .I(DLX_IFinst__n0003[17]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_IR_latched<17>/FFX/RST ),
    .O(DLX_IFinst_IR_latched[17])
  );
  X_OR2 \DLX_IFinst_IR_latched<17>/FFX/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IFinst_IR_latched<17>/FFX/RST )
  );
  defparam DLX_IFinst_IR_latched_26.INIT = 1'b0;
  X_FF DLX_IFinst_IR_latched_26 (
    .I(DLX_IFinst__n0003[26]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_IR_latched<26>/FFX/RST ),
    .O(DLX_IFinst_IR_latched[26])
  );
  X_OR2 \DLX_IFinst_IR_latched<26>/FFX/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IFinst_IR_latched<26>/FFX/RST )
  );
  defparam DLX_IFinst_IR_latched_18.INIT = 1'b0;
  X_FF DLX_IFinst_IR_latched_18 (
    .I(DLX_IFinst__n0003[18]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_IR_latched<18>/FFX/RST ),
    .O(DLX_IFinst_IR_latched[18])
  );
  X_OR2 \DLX_IFinst_IR_latched<18>/FFX/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IFinst_IR_latched<18>/FFX/RST )
  );
  defparam DLX_IFinst_IR_latched_27.INIT = 1'b0;
  X_FF DLX_IFinst_IR_latched_27 (
    .I(DLX_IFinst__n0003[27]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_IR_latched<27>/FFX/RST ),
    .O(DLX_IFinst_IR_latched[27])
  );
  X_OR2 \DLX_IFinst_IR_latched<27>/FFX/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IFinst_IR_latched<27>/FFX/RST )
  );
  defparam DLX_IFinst_IR_latched_19.INIT = 1'b0;
  X_FF DLX_IFinst_IR_latched_19 (
    .I(DLX_IFinst__n0003[19]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_IR_latched<19>/FFX/RST ),
    .O(DLX_IFinst_IR_latched[19])
  );
  X_OR2 \DLX_IFinst_IR_latched<19>/FFX/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IFinst_IR_latched<19>/FFX/RST )
  );
  defparam DLX_IFinst_IR_latched_28.INIT = 1'b0;
  X_FF DLX_IFinst_IR_latched_28 (
    .I(DLX_IFinst__n0003[28]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_IR_latched<28>/FFX/RST ),
    .O(DLX_IFinst_IR_latched[28])
  );
  X_OR2 \DLX_IFinst_IR_latched<28>/FFX/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IFinst_IR_latched<28>/FFX/RST )
  );
  defparam DLX_IFinst_IR_latched_29.INIT = 1'b0;
  X_FF DLX_IFinst_IR_latched_29 (
    .I(DLX_IFinst__n0003[29]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_IR_latched<29>/FFX/RST ),
    .O(DLX_IFinst_IR_latched[29])
  );
  X_OR2 \DLX_IFinst_IR_latched<29>/FFX/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IFinst_IR_latched<29>/FFX/RST )
  );
  defparam DLX_IFinst_IR_latched_7.INIT = 1'b0;
  X_FF DLX_IFinst_IR_latched_7 (
    .I(DLX_IFinst__n0003[7]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_IR_latched<7>/FFX/RST ),
    .O(DLX_IFinst_IR_latched[7])
  );
  X_OR2 \DLX_IFinst_IR_latched<7>/FFX/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IFinst_IR_latched<7>/FFX/RST )
  );
  defparam DLX_IFinst_IR_latched_8.INIT = 1'b0;
  X_FF DLX_IFinst_IR_latched_8 (
    .I(DLX_IFinst__n0003[8]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_IR_latched<8>/FFX/RST ),
    .O(DLX_IFinst_IR_latched[8])
  );
  X_OR2 \DLX_IFinst_IR_latched<8>/FFX/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IFinst_IR_latched<8>/FFX/RST )
  );
  defparam DLX_IFinst_IR_latched_9.INIT = 1'b0;
  X_FF DLX_IFinst_IR_latched_9 (
    .I(DLX_IFinst__n0003[9]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_IR_latched<9>/FFX/RST ),
    .O(DLX_IFinst_IR_latched[9])
  );
  X_OR2 \DLX_IFinst_IR_latched<9>/FFX/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IFinst_IR_latched<9>/FFX/RST )
  );
  defparam DLX_reg_dst_of_MEM_4.INIT = 1'b0;
  X_SFF DLX_reg_dst_of_MEM_4 (
    .I(DLX_reg_dst_of_EX[4]),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_reg_dst_of_MEM[4])
  );
  defparam DLX_IFinst_PC_0.INIT = 1'b0;
  X_FF DLX_IFinst_PC_0 (
    .I(DLX_IFinst_NPC[0]),
    .CE(DLX_IFinst_PC_N3535),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_PC<1>/FFY/RST ),
    .O(DLX_IFinst_PC[0])
  );
  X_OR2 \DLX_IFinst_PC<1>/FFY/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_PC<1>/FFY/RST )
  );
  defparam DLX_EXinst_ALU_result_19.INIT = 1'b0;
  X_FF DLX_EXinst_ALU_result_19 (
    .I(N119626),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_ALU_result<19>/FFY/RST ),
    .O(DLX_EXinst_ALU_result[19])
  );
  X_OR2 \DLX_EXinst_ALU_result<19>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_ALU_result<19>/FFY/RST )
  );
  defparam DLX_IDinst_reg_out_A_8.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_A_8 (
    .I(N103216),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_A<8>/FFY/RST ),
    .O(DLX_IDinst_reg_out_A[8])
  );
  X_OR2 \DLX_IDinst_reg_out_A<8>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_A<8>/FFY/RST )
  );
  defparam DLX_IDinst_reg_out_A_9.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_A_9 (
    .I(N103284),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_A<9>/FFY/RST ),
    .O(DLX_IDinst_reg_out_A[9])
  );
  X_OR2 \DLX_IDinst_reg_out_A<9>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_A<9>/FFY/RST )
  );
  defparam DLX_IDinst_IR_opcode_field_1.INIT = 1'b0;
  X_FF DLX_IDinst_IR_opcode_field_1 (
    .I(DLX_IDinst__n0113[1]),
    .CE(DLX_IDinst__n0422),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_IR_opcode_field<1>/FFY/RST ),
    .O(DLX_IDinst_IR_opcode_field[1])
  );
  X_OR2 \DLX_IDinst_IR_opcode_field<1>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_IR_opcode_field<1>/FFY/RST )
  );
  defparam vga_top_vga1_vcounter_4.INIT = 1'b0;
  X_SFF vga_top_vga1_vcounter_4 (
    .I(vga_top_vga1_vcounter__n0000[4]),
    .CE(N108996),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0007),
    .O(vga_top_vga1_vcounter[4])
  );
  defparam vga_top_vga1_vcounter_6.INIT = 1'b0;
  X_SFF vga_top_vga1_vcounter_6 (
    .I(vga_top_vga1_vcounter__n0000[6]),
    .CE(N108996),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0007),
    .O(vga_top_vga1_vcounter[6])
  );
  defparam vga_top_vga1_vcounter_9.INIT = 1'b0;
  X_SFF vga_top_vga1_vcounter_9 (
    .I(vga_top_vga1_vcounter__n0000[9]),
    .CE(N108996),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0007),
    .O(vga_top_vga1_vcounter[9])
  );
  defparam vga_top_vga1_hcounter_3.INIT = 1'b0;
  X_SFF vga_top_vga1_hcounter_3 (
    .I(vga_top_vga1_hcounter__n0000[3]),
    .CE(VCC),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0006),
    .O(vga_top_vga1_hcounter[3])
  );
  defparam vga_top_vga1_vcounter_8.INIT = 1'b0;
  X_SFF vga_top_vga1_vcounter_8 (
    .I(vga_top_vga1_vcounter__n0000[8]),
    .CE(N108996),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0007),
    .O(vga_top_vga1_vcounter[8])
  );
  defparam vga_top_vga1_hcounter_1.INIT = 1'b0;
  X_SFF vga_top_vga1_hcounter_1 (
    .I(vga_top_vga1_hcounter__n0000[1]),
    .CE(VCC),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0006),
    .O(vga_top_vga1_hcounter[1])
  );
  defparam vga_top_vga1_hcounter_0.INIT = 1'b0;
  X_SFF vga_top_vga1_hcounter_0 (
    .I(vga_top_vga1_hcounter_Madd__n0000_inst_lut2_19),
    .CE(VCC),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0006),
    .O(vga_top_vga1_hcounter[0])
  );
  defparam vga_top_vga1_hcounter_2.INIT = 1'b0;
  X_SFF vga_top_vga1_hcounter_2 (
    .I(vga_top_vga1_hcounter__n0000[2]),
    .CE(VCC),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0006),
    .O(vga_top_vga1_hcounter[2])
  );
  defparam vga_top_vga1_hcounter_5.INIT = 1'b0;
  X_SFF vga_top_vga1_hcounter_5 (
    .I(vga_top_vga1_hcounter__n0000[5]),
    .CE(VCC),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0006),
    .O(vga_top_vga1_hcounter[5])
  );
  defparam vga_top_vga1_hcounter_9.INIT = 1'b0;
  X_SFF vga_top_vga1_hcounter_9 (
    .I(vga_top_vga1_hcounter__n0000[9]),
    .CE(VCC),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0006),
    .O(vga_top_vga1_hcounter[9])
  );
  defparam vga_top_vga1_hcounter_4.INIT = 1'b0;
  X_SFF vga_top_vga1_hcounter_4 (
    .I(vga_top_vga1_hcounter__n0000[4]),
    .CE(VCC),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0006),
    .O(vga_top_vga1_hcounter[4])
  );
  defparam vga_top_vga1_hcounter_7.INIT = 1'b0;
  X_SFF vga_top_vga1_hcounter_7 (
    .I(vga_top_vga1_hcounter__n0000[7]),
    .CE(VCC),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0006),
    .O(vga_top_vga1_hcounter[7])
  );
  defparam vga_top_vga1_hcounter_6.INIT = 1'b0;
  X_SFF vga_top_vga1_hcounter_6 (
    .I(vga_top_vga1_hcounter__n0000[6]),
    .CE(VCC),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0006),
    .O(vga_top_vga1_hcounter[6])
  );
  defparam vga_top_vga1_hcounter_8.INIT = 1'b0;
  X_SFF vga_top_vga1_hcounter_8 (
    .I(vga_top_vga1_hcounter__n0000[8]),
    .CE(VCC),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0006),
    .O(vga_top_vga1_hcounter[8])
  );
  defparam vga_top_vga1_hcounter_11.INIT = 1'b0;
  X_SFF vga_top_vga1_hcounter_11 (
    .I(vga_top_vga1_hcounter__n0000[11]),
    .CE(VCC),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0006),
    .O(vga_top_vga1_hcounter[11])
  );
  defparam vga_top_vga1_hcounter_15.INIT = 1'b0;
  X_SFF vga_top_vga1_hcounter_15 (
    .I(vga_top_vga1_hcounter__n0000[15]),
    .CE(VCC),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0006),
    .O(vga_top_vga1_hcounter[15])
  );
  defparam vga_top_vga1_hcounter_10.INIT = 1'b0;
  X_SFF vga_top_vga1_hcounter_10 (
    .I(vga_top_vga1_hcounter__n0000[10]),
    .CE(VCC),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0006),
    .O(vga_top_vga1_hcounter[10])
  );
  defparam vga_top_vga1_hcounter_13.INIT = 1'b0;
  X_SFF vga_top_vga1_hcounter_13 (
    .I(vga_top_vga1_hcounter__n0000[13]),
    .CE(VCC),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0006),
    .O(vga_top_vga1_hcounter[13])
  );
  defparam vga_top_vga1_hcounter_12.INIT = 1'b0;
  X_SFF vga_top_vga1_hcounter_12 (
    .I(vga_top_vga1_hcounter__n0000[12]),
    .CE(VCC),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0006),
    .O(vga_top_vga1_hcounter[12])
  );
  defparam vga_top_vga1_hcounter_14.INIT = 1'b0;
  X_SFF vga_top_vga1_hcounter_14 (
    .I(vga_top_vga1_hcounter__n0000[14]),
    .CE(VCC),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0006),
    .O(vga_top_vga1_hcounter[14])
  );
  defparam DLX_IDinst_Imm_11.INIT = 1'b0;
  X_FF DLX_IDinst_Imm_11 (
    .I(DLX_IDinst__n0094),
    .CE(DLX_IDinst__n0422),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_Imm<11>/FFY/RST ),
    .O(\DLX_IDinst_Imm[11] )
  );
  X_OR2 \DLX_IDinst_Imm<11>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_Imm<11>/FFY/RST )
  );
  defparam DLX_IDinst_delay_slot_1185.INIT = 1'b0;
  X_FF DLX_IDinst_delay_slot_1185 (
    .I(N109531),
    .CE(DLX_IDinst__n0442),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_delay_slot/FFY/RST ),
    .O(DLX_IDinst_delay_slot)
  );
  X_OR2 \DLX_IDinst_delay_slot/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_delay_slot/FFY/RST )
  );
  defparam vga_top_vga1_gridvcounter_1.INIT = 1'b0;
  X_SFF vga_top_vga1_gridvcounter_1 (
    .I(vga_top_vga1_gridvcounter__n0000[1]),
    .CE(vga_top_vga1_N73384),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0014),
    .O(vga_top_vga1_gridvcounter[1])
  );
  defparam vga_top_vga1_gridvcounter_3.INIT = 1'b0;
  X_SFF vga_top_vga1_gridvcounter_3 (
    .I(vga_top_vga1_gridvcounter__n0000[3]),
    .CE(vga_top_vga1_N73384),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0014),
    .O(vga_top_vga1_gridvcounter[3])
  );
  defparam vga_top_vga1_gridvcounter_0.INIT = 1'b0;
  X_SFF vga_top_vga1_gridvcounter_0 (
    .I(vga_top_vga1_gridvcounter_Madd__n0000_inst_lut2_0),
    .CE(vga_top_vga1_N73384),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0014),
    .O(vga_top_vga1_gridvcounter[0])
  );
  defparam vga_top_vga1_gridvcounter_5.INIT = 1'b0;
  X_SFF vga_top_vga1_gridvcounter_5 (
    .I(vga_top_vga1_gridvcounter__n0000[5]),
    .CE(vga_top_vga1_N73384),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0014),
    .O(vga_top_vga1_gridvcounter[5])
  );
  defparam vga_top_vga1_gridvcounter_2.INIT = 1'b0;
  X_SFF vga_top_vga1_gridvcounter_2 (
    .I(vga_top_vga1_gridvcounter__n0000[2]),
    .CE(vga_top_vga1_N73384),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0014),
    .O(vga_top_vga1_gridvcounter[2])
  );
  defparam vga_top_vga1_gridvcounter_4.INIT = 1'b0;
  X_SFF vga_top_vga1_gridvcounter_4 (
    .I(vga_top_vga1_gridvcounter__n0000[4]),
    .CE(vga_top_vga1_N73384),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0014),
    .O(vga_top_vga1_gridvcounter[4])
  );
  defparam vga_top_vga1_gridvcounter_7.INIT = 1'b0;
  X_SFF vga_top_vga1_gridvcounter_7 (
    .I(vga_top_vga1_gridvcounter__n0000[7]),
    .CE(vga_top_vga1_N73384),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0014),
    .O(vga_top_vga1_gridvcounter[7])
  );
  defparam vga_top_vga1_gridvcounter_8.INIT = 1'b0;
  X_SFF vga_top_vga1_gridvcounter_8 (
    .I(vga_top_vga1_gridvcounter__n0000[8]),
    .CE(vga_top_vga1_N73384),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0014),
    .O(vga_top_vga1_gridvcounter[8])
  );
  defparam vga_top_vga1_gridvcounter_6.INIT = 1'b0;
  X_SFF vga_top_vga1_gridvcounter_6 (
    .I(vga_top_vga1_gridvcounter__n0000[6]),
    .CE(vga_top_vga1_N73384),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0014),
    .O(vga_top_vga1_gridvcounter[6])
  );
  defparam DLX_EXinst_reg_out_B_EX_30.INIT = 1'b0;
  X_FF DLX_EXinst_reg_out_B_EX_30 (
    .I(DLX_EXinst__n0007[30]),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_reg_out_B_EX<30>/FFY/RST ),
    .O(DLX_EXinst_reg_out_B_EX[30])
  );
  X_OR2 \DLX_EXinst_reg_out_B_EX<30>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_reg_out_B_EX<30>/FFY/RST )
  );
  defparam DLX_MEMinst_RF_data_in_15.INIT = 1'b0;
  X_FF DLX_MEMinst_RF_data_in_15 (
    .I(DLX_MEMinst__n0000[15]),
    .CE(VCC),
    .CLK(\DLX_MEMinst_RF_data_in<15>/CKMUXNOT ),
    .SET(GND),
    .RST(\DLX_MEMinst_RF_data_in<15>/FFX/RST ),
    .O(DLX_MEMinst_RF_data_in[15])
  );
  X_OR2 \DLX_MEMinst_RF_data_in<15>/FFX/RSTOR  (
    .I0(reset_IBUF_1),
    .I1(GSR),
    .O(\DLX_MEMinst_RF_data_in<15>/FFX/RST )
  );
  defparam DLX_MEMinst_RF_data_in_25.INIT = 1'b0;
  X_FF DLX_MEMinst_RF_data_in_25 (
    .I(DLX_MEMinst__n0000[25]),
    .CE(VCC),
    .CLK(\DLX_MEMinst_RF_data_in<25>/CKMUXNOT ),
    .SET(GND),
    .RST(\DLX_MEMinst_RF_data_in<25>/FFX/RST ),
    .O(DLX_MEMinst_RF_data_in[25])
  );
  X_OR2 \DLX_MEMinst_RF_data_in<25>/FFX/RSTOR  (
    .I0(reset_IBUF_1),
    .I1(GSR),
    .O(\DLX_MEMinst_RF_data_in<25>/FFX/RST )
  );
  defparam DLX_MEMinst_RF_data_in_17.INIT = 1'b0;
  X_FF DLX_MEMinst_RF_data_in_17 (
    .I(DLX_MEMinst__n0000[17]),
    .CE(VCC),
    .CLK(\DLX_MEMinst_RF_data_in<17>/CKMUXNOT ),
    .SET(GND),
    .RST(\DLX_MEMinst_RF_data_in<17>/FFX/RST ),
    .O(DLX_MEMinst_RF_data_in[17])
  );
  X_OR2 \DLX_MEMinst_RF_data_in<17>/FFX/RSTOR  (
    .I0(reset_IBUF_1),
    .I1(GSR),
    .O(\DLX_MEMinst_RF_data_in<17>/FFX/RST )
  );
  defparam DLX_MEMinst_RF_data_in_27.INIT = 1'b0;
  X_FF DLX_MEMinst_RF_data_in_27 (
    .I(DLX_MEMinst__n0000[27]),
    .CE(VCC),
    .CLK(\DLX_MEMinst_RF_data_in<27>/CKMUXNOT ),
    .SET(GND),
    .RST(\DLX_MEMinst_RF_data_in<27>/FFX/RST ),
    .O(DLX_MEMinst_RF_data_in[27])
  );
  X_OR2 \DLX_MEMinst_RF_data_in<27>/FFX/RSTOR  (
    .I0(reset_IBUF_1),
    .I1(GSR),
    .O(\DLX_MEMinst_RF_data_in<27>/FFX/RST )
  );
  defparam vga_top_vga1_gridhcounter_1.INIT = 1'b0;
  X_SFF vga_top_vga1_gridhcounter_1 (
    .I(vga_top_vga1_gridhcounter__n0000[1]),
    .CE(vga_top_vga1__n0013),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0012),
    .O(vga_top_vga1_gridhcounter[1])
  );
  defparam vga_top_vga1_gridhcounter_3.INIT = 1'b0;
  X_SFF vga_top_vga1_gridhcounter_3 (
    .I(vga_top_vga1_gridhcounter__n0000[3]),
    .CE(vga_top_vga1__n0013),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0012),
    .O(vga_top_vga1_gridhcounter[3])
  );
  defparam DLX_EXinst_mem_to_reg_EX_1186.INIT = 1'b0;
  X_FF DLX_EXinst_mem_to_reg_EX_1186 (
    .I(DLX_EXinst__n0010),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_mem_to_reg_EX/FFX/RST ),
    .O(DLX_EXinst_mem_to_reg_EX)
  );
  X_OR2 \DLX_EXinst_mem_to_reg_EX/FFX/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_mem_to_reg_EX/FFX/RST )
  );
  defparam DLX_IDinst_EPC_9.INIT = 1'b0;
  X_FF DLX_IDinst_EPC_9 (
    .I(DLX_IDinst__n0123[9]),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_EPC<9>/FFX/RST ),
    .O(DLX_IDinst_EPC[9])
  );
  X_OR2 \DLX_IDinst_EPC<9>/FFX/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_EPC<9>/FFX/RST )
  );
  defparam DLX_IDinst_reg_out_B_2_1_1187.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_B_2_1_1187 (
    .I(\DLX_IDinst_reg_out_B_2_1/GROM ),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_B_2_1/FFY/RST ),
    .O(DLX_IDinst_reg_out_B_2_1)
  );
  X_OR2 \DLX_IDinst_reg_out_B_2_1/FFY/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_B_2_1/FFY/RST )
  );
  defparam DLX_IDinst_reg_out_B_3_1_1188.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_B_3_1_1188 (
    .I(\DLX_IDinst_reg_out_B<3>/GROM ),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_B<3>/FFY/RST ),
    .O(DLX_IDinst_reg_out_B_3_1)
  );
  X_OR2 \DLX_IDinst_reg_out_B<3>/FFY/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_B<3>/FFY/RST )
  );
  defparam DLX_EXinst_ALU_result_12.INIT = 1'b0;
  X_FF DLX_EXinst_ALU_result_12 (
    .I(\DLX_EXinst_ALU_result<13>/GROM ),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_ALU_result<13>/FFY/RST ),
    .O(DLX_EXinst_ALU_result[12])
  );
  X_OR2 \DLX_EXinst_ALU_result<13>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_ALU_result<13>/FFY/RST )
  );
  defparam DLX_IDinst_reg_out_B_3.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_B_3 (
    .I(DLX_IDinst__n0118[3]),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_B<3>/FFX/RST ),
    .O(DLX_IDinst_reg_out_B[3])
  );
  X_OR2 \DLX_IDinst_reg_out_B<3>/FFX/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_B<3>/FFX/RST )
  );
  defparam DLX_EXinst_ALU_result_13.INIT = 1'b0;
  X_FF DLX_EXinst_ALU_result_13 (
    .I(\DLX_EXinst_ALU_result<13>/FROM ),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_ALU_result<13>/FFX/RST ),
    .O(DLX_EXinst_ALU_result[13])
  );
  X_OR2 \DLX_EXinst_ALU_result<13>/FFX/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_ALU_result<13>/FFX/RST )
  );
  defparam DLX_IDinst_current_IR_7.INIT = 1'b0;
  X_FF DLX_IDinst_current_IR_7 (
    .I(\DLX_IDinst_current_IR<7>/FROM ),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_current_IR<7>/FFX/RST ),
    .O(DLX_IDinst_current_IR[7])
  );
  X_OR2 \DLX_IDinst_current_IR<7>/FFX/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_current_IR<7>/FFX/RST )
  );
  defparam DLX_IDinst_EPC_0.INIT = 1'b0;
  X_FF DLX_IDinst_EPC_0 (
    .I(DLX_IDinst__n0123[0]),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_EPC<1>/FFY/RST ),
    .O(DLX_IDinst_EPC[0])
  );
  X_OR2 \DLX_IDinst_EPC<1>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_EPC<1>/FFY/RST )
  );
  defparam DLX_IDinst_current_IR_9.INIT = 1'b0;
  X_FF DLX_IDinst_current_IR_9 (
    .I(\DLX_IDinst_current_IR<9>/FROM ),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_current_IR<9>/FFX/RST ),
    .O(DLX_IDinst_current_IR[9])
  );
  X_OR2 \DLX_IDinst_current_IR<9>/FFX/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_current_IR<9>/FFX/RST )
  );
  defparam DLX_IDinst_EPC_1.INIT = 1'b0;
  X_FF DLX_IDinst_EPC_1 (
    .I(DLX_IDinst__n0123[1]),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_EPC<1>/FFX/RST ),
    .O(DLX_IDinst_EPC[1])
  );
  X_OR2 \DLX_IDinst_EPC<1>/FFX/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_EPC<1>/FFX/RST )
  );
  defparam DLX_IDinst_EPC_2.INIT = 1'b0;
  X_FF DLX_IDinst_EPC_2 (
    .I(DLX_IDinst__n0123[2]),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_EPC<3>/FFY/RST ),
    .O(DLX_IDinst_EPC[2])
  );
  X_OR2 \DLX_IDinst_EPC<3>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_EPC<3>/FFY/RST )
  );
  defparam DLX_IDinst_EPC_3.INIT = 1'b0;
  X_FF DLX_IDinst_EPC_3 (
    .I(DLX_IDinst__n0123[3]),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_EPC<3>/FFX/RST ),
    .O(DLX_IDinst_EPC[3])
  );
  X_OR2 \DLX_IDinst_EPC<3>/FFX/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_EPC<3>/FFX/RST )
  );
  defparam DLX_IDinst_EPC_4.INIT = 1'b0;
  X_FF DLX_IDinst_EPC_4 (
    .I(DLX_IDinst__n0123[4]),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_EPC<5>/FFY/RST ),
    .O(DLX_IDinst_EPC[4])
  );
  X_OR2 \DLX_IDinst_EPC<5>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_EPC<5>/FFY/RST )
  );
  defparam DLX_IDinst_EPC_5.INIT = 1'b0;
  X_FF DLX_IDinst_EPC_5 (
    .I(DLX_IDinst__n0123[5]),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_EPC<5>/FFX/RST ),
    .O(DLX_IDinst_EPC[5])
  );
  X_OR2 \DLX_IDinst_EPC<5>/FFX/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_EPC<5>/FFX/RST )
  );
  defparam DLX_IDinst_EPC_6.INIT = 1'b0;
  X_FF DLX_IDinst_EPC_6 (
    .I(DLX_IDinst__n0123[6]),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_EPC<7>/FFY/RST ),
    .O(DLX_IDinst_EPC[6])
  );
  X_OR2 \DLX_IDinst_EPC<7>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_EPC<7>/FFY/RST )
  );
  defparam DLX_IDinst_EPC_7.INIT = 1'b0;
  X_FF DLX_IDinst_EPC_7 (
    .I(DLX_IDinst__n0123[7]),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_EPC<7>/FFX/RST ),
    .O(DLX_IDinst_EPC[7])
  );
  X_OR2 \DLX_IDinst_EPC<7>/FFX/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_EPC<7>/FFX/RST )
  );
  defparam DLX_IDinst_EPC_8.INIT = 1'b0;
  X_FF DLX_IDinst_EPC_8 (
    .I(DLX_IDinst__n0123[8]),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_EPC<9>/FFY/RST ),
    .O(DLX_IDinst_EPC[8])
  );
  X_OR2 \DLX_IDinst_EPC<9>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_EPC<9>/FFY/RST )
  );
  defparam vga_top_vga1_gridhcounter_0.INIT = 1'b0;
  X_SFF vga_top_vga1_gridhcounter_0 (
    .I(vga_top_vga1_gridhcounter_Madd__n0000_inst_lut2_0),
    .CE(vga_top_vga1__n0013),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0012),
    .O(vga_top_vga1_gridhcounter[0])
  );
  defparam vga_top_vga1_gridhcounter_5.INIT = 1'b0;
  X_SFF vga_top_vga1_gridhcounter_5 (
    .I(vga_top_vga1_gridhcounter__n0000[5]),
    .CE(vga_top_vga1__n0013),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0012),
    .O(vga_top_vga1_gridhcounter[5])
  );
  defparam vga_top_vga1_gridhcounter_2.INIT = 1'b0;
  X_SFF vga_top_vga1_gridhcounter_2 (
    .I(vga_top_vga1_gridhcounter__n0000[2]),
    .CE(vga_top_vga1__n0013),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0012),
    .O(vga_top_vga1_gridhcounter[2])
  );
  defparam vga_top_vga1_gridhcounter_4.INIT = 1'b0;
  X_SFF vga_top_vga1_gridhcounter_4 (
    .I(vga_top_vga1_gridhcounter__n0000[4]),
    .CE(vga_top_vga1__n0013),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0012),
    .O(vga_top_vga1_gridhcounter[4])
  );
  defparam vga_top_vga1_gridhcounter_7.INIT = 1'b0;
  X_SFF vga_top_vga1_gridhcounter_7 (
    .I(vga_top_vga1_gridhcounter__n0000[7]),
    .CE(vga_top_vga1__n0013),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0012),
    .O(vga_top_vga1_gridhcounter[7])
  );
  defparam vga_top_vga1_gridhcounter_8.INIT = 1'b0;
  X_SFF vga_top_vga1_gridhcounter_8 (
    .I(vga_top_vga1_gridhcounter__n0000[8]),
    .CE(vga_top_vga1__n0013),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0012),
    .O(vga_top_vga1_gridhcounter[8])
  );
  defparam vga_top_vga1_gridhcounter_6.INIT = 1'b0;
  X_SFF vga_top_vga1_gridhcounter_6 (
    .I(vga_top_vga1_gridhcounter__n0000[6]),
    .CE(vga_top_vga1__n0013),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0012),
    .O(vga_top_vga1_gridhcounter[6])
  );
  defparam DLX_IDinst_current_IR_0.INIT = 1'b0;
  X_FF DLX_IDinst_current_IR_0 (
    .I(\DLX_IDinst_current_IR<1>/GROM ),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_current_IR<1>/FFY/RST ),
    .O(DLX_IDinst_current_IR[0])
  );
  X_OR2 \DLX_IDinst_current_IR<1>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_current_IR<1>/FFY/RST )
  );
  defparam DLX_IDinst_current_IR_2.INIT = 1'b0;
  X_FF DLX_IDinst_current_IR_2 (
    .I(\DLX_IDinst_current_IR<3>/GROM ),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_current_IR<3>/FFY/RST ),
    .O(DLX_IDinst_current_IR[2])
  );
  X_OR2 \DLX_IDinst_current_IR<3>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_current_IR<3>/FFY/RST )
  );
  defparam DLX_IDinst_current_IR_1.INIT = 1'b0;
  X_FF DLX_IDinst_current_IR_1 (
    .I(\DLX_IDinst_current_IR<1>/FROM ),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_current_IR<1>/FFX/RST ),
    .O(DLX_IDinst_current_IR[1])
  );
  X_OR2 \DLX_IDinst_current_IR<1>/FFX/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_current_IR<1>/FFX/RST )
  );
  defparam DLX_IDinst_current_IR_4.INIT = 1'b0;
  X_FF DLX_IDinst_current_IR_4 (
    .I(\DLX_IDinst_current_IR<5>/GROM ),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_current_IR<5>/FFY/RST ),
    .O(DLX_IDinst_current_IR[4])
  );
  X_OR2 \DLX_IDinst_current_IR<5>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_current_IR<5>/FFY/RST )
  );
  defparam DLX_IDinst_current_IR_3.INIT = 1'b0;
  X_FF DLX_IDinst_current_IR_3 (
    .I(\DLX_IDinst_current_IR<3>/FROM ),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_current_IR<3>/FFX/RST ),
    .O(DLX_IDinst_current_IR[3])
  );
  X_OR2 \DLX_IDinst_current_IR<3>/FFX/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_current_IR<3>/FFX/RST )
  );
  defparam DLX_IDinst_current_IR_6.INIT = 1'b0;
  X_FF DLX_IDinst_current_IR_6 (
    .I(\DLX_IDinst_current_IR<7>/GROM ),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_current_IR<7>/FFY/RST ),
    .O(DLX_IDinst_current_IR[6])
  );
  X_OR2 \DLX_IDinst_current_IR<7>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_current_IR<7>/FFY/RST )
  );
  defparam DLX_IDinst_current_IR_5.INIT = 1'b0;
  X_FF DLX_IDinst_current_IR_5 (
    .I(\DLX_IDinst_current_IR<5>/FROM ),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_current_IR<5>/FFX/RST ),
    .O(DLX_IDinst_current_IR[5])
  );
  X_OR2 \DLX_IDinst_current_IR<5>/FFX/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_current_IR<5>/FFX/RST )
  );
  defparam DLX_IDinst_current_IR_8.INIT = 1'b0;
  X_FF DLX_IDinst_current_IR_8 (
    .I(\DLX_IDinst_current_IR<9>/GROM ),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_current_IR<9>/FFY/RST ),
    .O(DLX_IDinst_current_IR[8])
  );
  X_OR2 \DLX_IDinst_current_IR<9>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_current_IR<9>/FFY/RST )
  );
  defparam DLX_IDinst_slot_num_FFd1_1189.INIT = 1'b0;
  X_FF DLX_IDinst_slot_num_FFd1_1189 (
    .I(\DLX_IDinst_slot_num_FFd1-In ),
    .CE(DLX_IDinst__n0420),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_slot_num_FFd1/FFY/RST ),
    .O(DLX_IDinst_slot_num_FFd1)
  );
  X_OR2 \DLX_IDinst_slot_num_FFd1/FFY/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IDinst_slot_num_FFd1/FFY/RST )
  );
  defparam DLX_reg_dst_of_MEM_3.INIT = 1'b0;
  X_SFF DLX_reg_dst_of_MEM_3 (
    .I(\DLX_reg_dst_of_MEM<3>/FROM ),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_reg_dst_of_MEM[3])
  );
  defparam DLX_IDinst_Cause_Reg_0.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_0 (
    .I(DLX_IDinst__n0127[0]),
    .CE(DLX_IDinst__n0085),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<1>/FFY/RST ),
    .O(DLX_IDinst_Cause_Reg[0])
  );
  X_BUF \DLX_IDinst_Cause_Reg<1>/FFY/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<1>/FFY/RST )
  );
  defparam DLX_EXinst_mem_write_EX_1190.INIT = 1'b0;
  X_FF DLX_EXinst_mem_write_EX_1190 (
    .I(\DLX_EXinst_reg_write_EX/GROM ),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_reg_write_EX/FFY/RST ),
    .O(DLX_EXinst_mem_write_EX)
  );
  X_OR2 \DLX_EXinst_reg_write_EX/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_reg_write_EX/FFY/RST )
  );
  defparam DLX_IDinst_Cause_Reg_2.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_2 (
    .I(DLX_IDinst__n0127[2]),
    .CE(DLX_IDinst__n0085),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<3>/FFY/RST ),
    .O(DLX_IDinst_Cause_Reg[2])
  );
  X_BUF \DLX_IDinst_Cause_Reg<3>/FFY/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<3>/FFY/RST )
  );
  defparam DLX_EXinst_reg_write_EX_1191.INIT = 1'b0;
  X_FF DLX_EXinst_reg_write_EX_1191 (
    .I(DLX_EXinst__n0009),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_reg_write_EX/FFX/RST ),
    .O(DLX_EXinst_reg_write_EX)
  );
  X_OR2 \DLX_EXinst_reg_write_EX/FFX/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_reg_write_EX/FFX/RST )
  );
  defparam DLX_IDinst_Cause_Reg_1.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_1 (
    .I(DLX_IDinst__n0127[1]),
    .CE(DLX_IDinst__n0085),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<1>/FFX/RST ),
    .O(DLX_IDinst_Cause_Reg[1])
  );
  X_BUF \DLX_IDinst_Cause_Reg<1>/FFX/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<1>/FFX/RST )
  );
  defparam DLX_IDinst_Cause_Reg_3.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_3 (
    .I(DLX_IDinst__n0127[3]),
    .CE(DLX_IDinst__n0085),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<3>/FFX/RST ),
    .O(DLX_IDinst_Cause_Reg[3])
  );
  X_BUF \DLX_IDinst_Cause_Reg<3>/FFX/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<3>/FFX/RST )
  );
  defparam DLX_IDinst_Cause_Reg_4.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_4 (
    .I(DLX_IDinst__n0127[4]),
    .CE(DLX_IDinst__n0085),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<5>/FFY/RST ),
    .O(DLX_IDinst_Cause_Reg[4])
  );
  X_BUF \DLX_IDinst_Cause_Reg<5>/FFY/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<5>/FFY/RST )
  );
  defparam DLX_IDinst_Cause_Reg_5.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_5 (
    .I(DLX_IDinst__n0127[5]),
    .CE(DLX_IDinst__n0085),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<5>/FFX/RST ),
    .O(DLX_IDinst_Cause_Reg[5])
  );
  X_BUF \DLX_IDinst_Cause_Reg<5>/FFX/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<5>/FFX/RST )
  );
  defparam DLX_IDinst_Cause_Reg_6.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_6 (
    .I(DLX_IDinst__n0127[6]),
    .CE(DLX_IDinst__n0085),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<7>/FFY/RST ),
    .O(DLX_IDinst_Cause_Reg[6])
  );
  X_BUF \DLX_IDinst_Cause_Reg<7>/FFY/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<7>/FFY/RST )
  );
  defparam DLX_IDinst_EPC_11.INIT = 1'b0;
  X_FF DLX_IDinst_EPC_11 (
    .I(DLX_IDinst__n0123[11]),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_EPC<11>/FFX/RST ),
    .O(DLX_IDinst_EPC[11])
  );
  X_OR2 \DLX_IDinst_EPC<11>/FFX/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_EPC<11>/FFX/RST )
  );
  defparam DLX_IDinst_EPC_13.INIT = 1'b0;
  X_FF DLX_IDinst_EPC_13 (
    .I(DLX_IDinst__n0123[13]),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_EPC<13>/FFX/RST ),
    .O(DLX_IDinst_EPC[13])
  );
  X_OR2 \DLX_IDinst_EPC<13>/FFX/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_EPC<13>/FFX/RST )
  );
  defparam DLX_IDinst_EPC_20.INIT = 1'b0;
  X_FF DLX_IDinst_EPC_20 (
    .I(DLX_IDinst__n0123[20]),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_EPC<21>/FFY/RST ),
    .O(DLX_IDinst_EPC[20])
  );
  X_OR2 \DLX_IDinst_EPC<21>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_EPC<21>/FFY/RST )
  );
  defparam DLX_IDinst_EPC_21.INIT = 1'b0;
  X_FF DLX_IDinst_EPC_21 (
    .I(DLX_IDinst__n0123[21]),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_EPC<21>/FFX/RST ),
    .O(DLX_IDinst_EPC[21])
  );
  X_OR2 \DLX_IDinst_EPC<21>/FFX/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_EPC<21>/FFX/RST )
  );
  defparam DLX_IDinst_EPC_14.INIT = 1'b0;
  X_FF DLX_IDinst_EPC_14 (
    .I(DLX_IDinst__n0123[14]),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_EPC<15>/FFY/RST ),
    .O(DLX_IDinst_EPC[14])
  );
  X_OR2 \DLX_IDinst_EPC<15>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_EPC<15>/FFY/RST )
  );
  defparam DLX_IDinst_EPC_15.INIT = 1'b0;
  X_FF DLX_IDinst_EPC_15 (
    .I(DLX_IDinst__n0123[15]),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_EPC<15>/FFX/RST ),
    .O(DLX_IDinst_EPC[15])
  );
  X_OR2 \DLX_IDinst_EPC<15>/FFX/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_EPC<15>/FFX/RST )
  );
  defparam DLX_IDinst_EPC_22.INIT = 1'b0;
  X_FF DLX_IDinst_EPC_22 (
    .I(DLX_IDinst__n0123[22]),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_EPC<23>/FFY/RST ),
    .O(DLX_IDinst_EPC[22])
  );
  X_OR2 \DLX_IDinst_EPC<23>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_EPC<23>/FFY/RST )
  );
  defparam DLX_IDinst_EPC_23.INIT = 1'b0;
  X_FF DLX_IDinst_EPC_23 (
    .I(DLX_IDinst__n0123[23]),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_EPC<23>/FFX/RST ),
    .O(DLX_IDinst_EPC[23])
  );
  X_OR2 \DLX_IDinst_EPC<23>/FFX/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_EPC<23>/FFX/RST )
  );
  defparam DLX_IDinst_EPC_24.INIT = 1'b0;
  X_FF DLX_IDinst_EPC_24 (
    .I(DLX_IDinst__n0123[24]),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_EPC<25>/FFY/RST ),
    .O(DLX_IDinst_EPC[24])
  );
  X_OR2 \DLX_IDinst_EPC<25>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_EPC<25>/FFY/RST )
  );
  defparam DLX_IDinst_EPC_30.INIT = 1'b0;
  X_FF DLX_IDinst_EPC_30 (
    .I(DLX_IDinst__n0123[30]),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_EPC<31>/FFY/RST ),
    .O(DLX_IDinst_EPC[30])
  );
  X_OR2 \DLX_IDinst_EPC<31>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_EPC<31>/FFY/RST )
  );
  defparam DLX_IDinst_EPC_31.INIT = 1'b0;
  X_FF DLX_IDinst_EPC_31 (
    .I(DLX_IDinst__n0123[31]),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_EPC<31>/FFX/RST ),
    .O(DLX_IDinst_EPC[31])
  );
  X_OR2 \DLX_IDinst_EPC<31>/FFX/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_EPC<31>/FFX/RST )
  );
  defparam DLX_IDinst_EPC_16.INIT = 1'b0;
  X_FF DLX_IDinst_EPC_16 (
    .I(DLX_IDinst__n0123[16]),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_EPC<17>/FFY/RST ),
    .O(DLX_IDinst_EPC[16])
  );
  X_OR2 \DLX_IDinst_EPC<17>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_EPC<17>/FFY/RST )
  );
  defparam DLX_MEMinst_RF_data_in_19.INIT = 1'b0;
  X_FF DLX_MEMinst_RF_data_in_19 (
    .I(DLX_MEMinst__n0000[19]),
    .CE(VCC),
    .CLK(\DLX_MEMinst_RF_data_in<19>/CKMUXNOT ),
    .SET(GND),
    .RST(\DLX_MEMinst_RF_data_in<19>/FFX/RST ),
    .O(DLX_MEMinst_RF_data_in[19])
  );
  X_OR2 \DLX_MEMinst_RF_data_in<19>/FFX/RSTOR  (
    .I0(reset_IBUF_1),
    .I1(GSR),
    .O(\DLX_MEMinst_RF_data_in<19>/FFX/RST )
  );
  defparam DLX_MEMinst_RF_data_in_29.INIT = 1'b0;
  X_FF DLX_MEMinst_RF_data_in_29 (
    .I(DLX_MEMinst__n0000[29]),
    .CE(VCC),
    .CLK(\DLX_MEMinst_RF_data_in<29>/CKMUXNOT ),
    .SET(GND),
    .RST(\DLX_MEMinst_RF_data_in<29>/FFX/RST ),
    .O(DLX_MEMinst_RF_data_in[29])
  );
  X_OR2 \DLX_MEMinst_RF_data_in<29>/FFX/RSTOR  (
    .I0(reset_IBUF_1),
    .I1(GSR),
    .O(\DLX_MEMinst_RF_data_in<29>/FFX/RST )
  );
  defparam DLX_IDinst_current_IR_20.INIT = 1'b0;
  X_FF DLX_IDinst_current_IR_20 (
    .I(\DLX_IDinst_current_IR<20>/GROM ),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_current_IR<20>/FFY/RST ),
    .O(DLX_IDinst_current_IR[20])
  );
  X_OR2 \DLX_IDinst_current_IR<20>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_current_IR<20>/FFY/RST )
  );
  defparam DLX_IDinst_current_IR_11.INIT = 1'b0;
  X_FF DLX_IDinst_current_IR_11 (
    .I(\DLX_IDinst_current_IR<11>/FROM ),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_current_IR<11>/FFX/RST ),
    .O(DLX_IDinst_current_IR[11])
  );
  X_OR2 \DLX_IDinst_current_IR<11>/FFX/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_current_IR<11>/FFX/RST )
  );
  defparam DLX_IDinst_current_IR_14.INIT = 1'b0;
  X_FF DLX_IDinst_current_IR_14 (
    .I(\DLX_IDinst_current_IR<15>/GROM ),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_current_IR<15>/FFY/RST ),
    .O(DLX_IDinst_current_IR[14])
  );
  X_OR2 \DLX_IDinst_current_IR<15>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_current_IR<15>/FFY/RST )
  );
  defparam DLX_IDinst_current_IR_12.INIT = 1'b0;
  X_FF DLX_IDinst_current_IR_12 (
    .I(\DLX_IDinst_current_IR<13>/GROM ),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_current_IR<13>/FFY/RST ),
    .O(DLX_IDinst_current_IR[12])
  );
  X_OR2 \DLX_IDinst_current_IR<13>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_current_IR<13>/FFY/RST )
  );
  defparam DLX_IDinst_current_IR_13.INIT = 1'b0;
  X_FF DLX_IDinst_current_IR_13 (
    .I(\DLX_IDinst_current_IR<13>/FROM ),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_current_IR<13>/FFX/RST ),
    .O(DLX_IDinst_current_IR[13])
  );
  X_OR2 \DLX_IDinst_current_IR<13>/FFX/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_current_IR<13>/FFX/RST )
  );
  defparam DLX_IDinst_current_IR_21.INIT = 1'b0;
  X_FF DLX_IDinst_current_IR_21 (
    .I(\DLX_IDinst_current_IR<21>/FROM ),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_current_IR<21>/FFX/RST ),
    .O(DLX_IDinst_current_IR[21])
  );
  X_OR2 \DLX_IDinst_current_IR<21>/FFX/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_current_IR<21>/FFX/RST )
  );
  defparam DLX_IDinst_current_IR_17.INIT = 1'b0;
  X_FF DLX_IDinst_current_IR_17 (
    .I(\DLX_IDinst_current_IR<17>/FROM ),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_current_IR<17>/FFX/RST ),
    .O(DLX_IDinst_current_IR[17])
  );
  X_OR2 \DLX_IDinst_current_IR<17>/FFX/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_current_IR<17>/FFX/RST )
  );
  defparam DLX_IDinst_current_IR_26.INIT = 1'b0;
  X_FF DLX_IDinst_current_IR_26 (
    .I(\DLX_IDinst_current_IR<26>/FROM ),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_current_IR<26>/FFX/RST ),
    .O(DLX_IDinst_current_IR[26])
  );
  X_OR2 \DLX_IDinst_current_IR<26>/FFX/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_current_IR<26>/FFX/RST )
  );
  defparam DLX_IDinst_current_IR_18.INIT = 1'b0;
  X_FF DLX_IDinst_current_IR_18 (
    .I(\DLX_IDinst_current_IR<19>/GROM ),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_current_IR<19>/FFY/RST ),
    .O(DLX_IDinst_current_IR[18])
  );
  X_OR2 \DLX_IDinst_current_IR<19>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_current_IR<19>/FFY/RST )
  );
  defparam DLX_IDinst_current_IR_19.INIT = 1'b0;
  X_FF DLX_IDinst_current_IR_19 (
    .I(\DLX_IDinst_current_IR<19>/FROM ),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_current_IR<19>/FFX/RST ),
    .O(DLX_IDinst_current_IR[19])
  );
  X_OR2 \DLX_IDinst_current_IR<19>/FFX/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_current_IR<19>/FFX/RST )
  );
  defparam DLX_IDinst_current_IR_27.INIT = 1'b0;
  X_FF DLX_IDinst_current_IR_27 (
    .I(\DLX_IDinst_current_IR<27>/FROM ),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_current_IR<27>/FFX/RST ),
    .O(DLX_IDinst_current_IR[27])
  );
  X_OR2 \DLX_IDinst_current_IR<27>/FFX/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_current_IR<27>/FFX/RST )
  );
  defparam DLX_IDinst_current_IR_28.INIT = 1'b0;
  X_FF DLX_IDinst_current_IR_28 (
    .I(\DLX_IDinst_current_IR<28>/FROM ),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_current_IR<28>/FFX/RST ),
    .O(DLX_IDinst_current_IR[28])
  );
  X_OR2 \DLX_IDinst_current_IR<28>/FFX/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_current_IR<28>/FFX/RST )
  );
  defparam DLX_IDinst_current_IR_29.INIT = 1'b0;
  X_FF DLX_IDinst_current_IR_29 (
    .I(\DLX_IDinst_current_IR<29>/FROM ),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_current_IR<29>/FFX/RST ),
    .O(DLX_IDinst_current_IR[29])
  );
  X_OR2 \DLX_IDinst_current_IR<29>/FFX/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_current_IR<29>/FFX/RST )
  );
  defparam DLX_IDinst_EPC_10.INIT = 1'b0;
  X_FF DLX_IDinst_EPC_10 (
    .I(DLX_IDinst__n0123[10]),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_EPC<11>/FFY/RST ),
    .O(DLX_IDinst_EPC[10])
  );
  X_OR2 \DLX_IDinst_EPC<11>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_EPC<11>/FFY/RST )
  );
  defparam DLX_IDinst_EPC_12.INIT = 1'b0;
  X_FF DLX_IDinst_EPC_12 (
    .I(DLX_IDinst__n0123[12]),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_EPC<13>/FFY/RST ),
    .O(DLX_IDinst_EPC[12])
  );
  X_OR2 \DLX_IDinst_EPC<13>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_EPC<13>/FFY/RST )
  );
  defparam DLX_IDinst_current_IR_22.INIT = 1'b0;
  X_FF DLX_IDinst_current_IR_22 (
    .I(\DLX_IDinst_current_IR<23>/GROM ),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_current_IR<23>/FFY/RST ),
    .O(DLX_IDinst_current_IR[22])
  );
  X_OR2 \DLX_IDinst_current_IR<23>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_current_IR<23>/FFY/RST )
  );
  defparam DLX_IDinst_current_IR_15.INIT = 1'b0;
  X_FF DLX_IDinst_current_IR_15 (
    .I(\DLX_IDinst_current_IR<15>/FROM ),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_current_IR<15>/FFX/RST ),
    .O(DLX_IDinst_current_IR[15])
  );
  X_OR2 \DLX_IDinst_current_IR<15>/FFX/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_current_IR<15>/FFX/RST )
  );
  defparam DLX_IDinst_current_IR_23.INIT = 1'b0;
  X_FF DLX_IDinst_current_IR_23 (
    .I(\DLX_IDinst_current_IR<23>/FROM ),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_current_IR<23>/FFX/RST ),
    .O(DLX_IDinst_current_IR[23])
  );
  X_OR2 \DLX_IDinst_current_IR<23>/FFX/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_current_IR<23>/FFX/RST )
  );
  defparam DLX_IDinst_current_IR_30.INIT = 1'b0;
  X_FF DLX_IDinst_current_IR_30 (
    .I(\DLX_IDinst_current_IR<30>/FROM ),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_current_IR<30>/FFX/RST ),
    .O(DLX_IDinst_current_IR[30])
  );
  X_OR2 \DLX_IDinst_current_IR<30>/FFX/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_current_IR<30>/FFX/RST )
  );
  defparam DLX_IDinst_current_IR_31.INIT = 1'b0;
  X_FF DLX_IDinst_current_IR_31 (
    .I(\DLX_IDinst_current_IR<31>/FROM ),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_current_IR<31>/FFX/RST ),
    .O(DLX_IDinst_current_IR[31])
  );
  X_OR2 \DLX_IDinst_current_IR<31>/FFX/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_current_IR<31>/FFX/RST )
  );
  defparam DLX_IDinst_current_IR_24.INIT = 1'b0;
  X_FF DLX_IDinst_current_IR_24 (
    .I(\DLX_IDinst_current_IR<24>/FROM ),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_current_IR<24>/FFX/RST ),
    .O(DLX_IDinst_current_IR[24])
  );
  X_OR2 \DLX_IDinst_current_IR<24>/FFX/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_current_IR<24>/FFX/RST )
  );
  defparam DLX_IDinst_current_IR_16.INIT = 1'b0;
  X_FF DLX_IDinst_current_IR_16 (
    .I(\DLX_IDinst_current_IR<17>/GROM ),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_current_IR<17>/FFY/RST ),
    .O(DLX_IDinst_current_IR[16])
  );
  X_OR2 \DLX_IDinst_current_IR<17>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_current_IR<17>/FFY/RST )
  );
  defparam DLX_IDinst_current_IR_25.INIT = 1'b0;
  X_FF DLX_IDinst_current_IR_25 (
    .I(\DLX_IDinst_current_IR<25>/GROM ),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_current_IR<25>/FFY/RST ),
    .O(DLX_IDinst_current_IR[25])
  );
  X_OR2 \DLX_IDinst_current_IR<25>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_current_IR<25>/FFY/RST )
  );
  defparam DLX_IDinst_Cause_Reg_7.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_7 (
    .I(DLX_IDinst__n0127[7]),
    .CE(DLX_IDinst__n0085),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<7>/FFX/RST ),
    .O(DLX_IDinst_Cause_Reg[7])
  );
  X_BUF \DLX_IDinst_Cause_Reg<7>/FFX/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<7>/FFX/RST )
  );
  defparam DLX_IDinst_Cause_Reg_8.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_8 (
    .I(DLX_IDinst__n0127[8]),
    .CE(DLX_IDinst__n0085),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<9>/FFY/RST ),
    .O(DLX_IDinst_Cause_Reg[8])
  );
  X_BUF \DLX_IDinst_Cause_Reg<9>/FFY/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<9>/FFY/RST )
  );
  defparam DLX_IDinst_Cause_Reg_9.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_9 (
    .I(DLX_IDinst__n0127[9]),
    .CE(DLX_IDinst__n0085),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<9>/FFX/RST ),
    .O(DLX_IDinst_Cause_Reg[9])
  );
  X_BUF \DLX_IDinst_Cause_Reg<9>/FFX/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<9>/FFX/RST )
  );
  defparam DLX_EXinst_reg_out_B_EX_10.INIT = 1'b0;
  X_FF DLX_EXinst_reg_out_B_EX_10 (
    .I(DLX_EXinst__n0007[10]),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_reg_out_B_EX<11>/FFY/RST ),
    .O(DLX_EXinst_reg_out_B_EX[10])
  );
  X_OR2 \DLX_EXinst_reg_out_B_EX<11>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_reg_out_B_EX<11>/FFY/RST )
  );
  defparam DLX_EXinst_reg_out_B_EX_11.INIT = 1'b0;
  X_FF DLX_EXinst_reg_out_B_EX_11 (
    .I(DLX_EXinst__n0007[11]),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_reg_out_B_EX<11>/FFX/RST ),
    .O(DLX_EXinst_reg_out_B_EX[11])
  );
  X_OR2 \DLX_EXinst_reg_out_B_EX<11>/FFX/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_reg_out_B_EX<11>/FFX/RST )
  );
  defparam DLX_IDinst_IR_function_field_0_1_1192.INIT = 1'b0;
  X_FF DLX_IDinst_IR_function_field_0_1_1192 (
    .I(\DLX_IDinst_IR_function_field<0>/GROM ),
    .CE(DLX_IDinst__n0422),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_IR_function_field<0>/FFY/RST ),
    .O(DLX_IDinst_IR_function_field_0_1)
  );
  X_OR2 \DLX_IDinst_IR_function_field<0>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_IR_function_field<0>/FFY/RST )
  );
  defparam DLX_EXinst_reg_out_B_EX_12.INIT = 1'b0;
  X_FF DLX_EXinst_reg_out_B_EX_12 (
    .I(DLX_EXinst__n0007[12]),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_reg_out_B_EX<13>/FFY/RST ),
    .O(DLX_EXinst_reg_out_B_EX[12])
  );
  X_OR2 \DLX_EXinst_reg_out_B_EX<13>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_reg_out_B_EX<13>/FFY/RST )
  );
  defparam DLX_EXinst_reg_out_B_EX_13.INIT = 1'b0;
  X_FF DLX_EXinst_reg_out_B_EX_13 (
    .I(DLX_EXinst__n0007[13]),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_reg_out_B_EX<13>/FFX/RST ),
    .O(DLX_EXinst_reg_out_B_EX[13])
  );
  X_OR2 \DLX_EXinst_reg_out_B_EX<13>/FFX/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_reg_out_B_EX<13>/FFX/RST )
  );
  defparam DLX_IDinst_IR_function_field_0.INIT = 1'b0;
  X_FF DLX_IDinst_IR_function_field_0 (
    .I(DLX_IDinst__n0105),
    .CE(DLX_IDinst__n0422),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_IR_function_field<0>/FFX/RST ),
    .O(DLX_IDinst_IR_function_field[0])
  );
  X_OR2 \DLX_IDinst_IR_function_field<0>/FFX/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_IR_function_field<0>/FFX/RST )
  );
  defparam DLX_EXinst_reg_out_B_EX_20.INIT = 1'b0;
  X_FF DLX_EXinst_reg_out_B_EX_20 (
    .I(DLX_EXinst__n0007[20]),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_reg_out_B_EX<21>/FFY/RST ),
    .O(DLX_EXinst_reg_out_B_EX[20])
  );
  X_OR2 \DLX_EXinst_reg_out_B_EX<21>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_reg_out_B_EX<21>/FFY/RST )
  );
  defparam DLX_EXinst_reg_out_B_EX_22.INIT = 1'b0;
  X_FF DLX_EXinst_reg_out_B_EX_22 (
    .I(DLX_EXinst__n0007[22]),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_reg_out_B_EX<23>/FFY/RST ),
    .O(DLX_EXinst_reg_out_B_EX[22])
  );
  X_OR2 \DLX_EXinst_reg_out_B_EX<23>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_reg_out_B_EX<23>/FFY/RST )
  );
  defparam DLX_EXinst_reg_out_B_EX_21.INIT = 1'b0;
  X_FF DLX_EXinst_reg_out_B_EX_21 (
    .I(DLX_EXinst__n0007[21]),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_reg_out_B_EX<21>/FFX/RST ),
    .O(DLX_EXinst_reg_out_B_EX[21])
  );
  X_OR2 \DLX_EXinst_reg_out_B_EX<21>/FFX/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_reg_out_B_EX<21>/FFX/RST )
  );
  defparam DLX_IDinst_EPC_17.INIT = 1'b0;
  X_FF DLX_IDinst_EPC_17 (
    .I(DLX_IDinst__n0123[17]),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_EPC<17>/FFX/RST ),
    .O(DLX_IDinst_EPC[17])
  );
  X_OR2 \DLX_IDinst_EPC<17>/FFX/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_EPC<17>/FFX/RST )
  );
  defparam DLX_IDinst_EPC_25.INIT = 1'b0;
  X_FF DLX_IDinst_EPC_25 (
    .I(DLX_IDinst__n0123[25]),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_EPC<25>/FFX/RST ),
    .O(DLX_IDinst_EPC[25])
  );
  X_OR2 \DLX_IDinst_EPC<25>/FFX/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_EPC<25>/FFX/RST )
  );
  defparam DLX_IDinst_EPC_18.INIT = 1'b0;
  X_FF DLX_IDinst_EPC_18 (
    .I(DLX_IDinst__n0123[18]),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_EPC<19>/FFY/RST ),
    .O(DLX_IDinst_EPC[18])
  );
  X_OR2 \DLX_IDinst_EPC<19>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_EPC<19>/FFY/RST )
  );
  defparam DLX_IDinst_EPC_19.INIT = 1'b0;
  X_FF DLX_IDinst_EPC_19 (
    .I(DLX_IDinst__n0123[19]),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_EPC<19>/FFX/RST ),
    .O(DLX_IDinst_EPC[19])
  );
  X_OR2 \DLX_IDinst_EPC<19>/FFX/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_EPC<19>/FFX/RST )
  );
  defparam DLX_IDinst_EPC_26.INIT = 1'b0;
  X_FF DLX_IDinst_EPC_26 (
    .I(DLX_IDinst__n0123[26]),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_EPC<27>/FFY/RST ),
    .O(DLX_IDinst_EPC[26])
  );
  X_OR2 \DLX_IDinst_EPC<27>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_EPC<27>/FFY/RST )
  );
  defparam DLX_IDinst_EPC_27.INIT = 1'b0;
  X_FF DLX_IDinst_EPC_27 (
    .I(DLX_IDinst__n0123[27]),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_EPC<27>/FFX/RST ),
    .O(DLX_IDinst_EPC[27])
  );
  X_OR2 \DLX_IDinst_EPC<27>/FFX/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_EPC<27>/FFX/RST )
  );
  defparam DLX_IDinst_EPC_28.INIT = 1'b0;
  X_FF DLX_IDinst_EPC_28 (
    .I(DLX_IDinst__n0123[28]),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_EPC<29>/FFY/RST ),
    .O(DLX_IDinst_EPC[28])
  );
  X_OR2 \DLX_IDinst_EPC<29>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_EPC<29>/FFY/RST )
  );
  defparam DLX_IDinst_EPC_29.INIT = 1'b0;
  X_FF DLX_IDinst_EPC_29 (
    .I(DLX_IDinst__n0123[29]),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_EPC<29>/FFX/RST ),
    .O(DLX_IDinst_EPC[29])
  );
  X_OR2 \DLX_IDinst_EPC<29>/FFX/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_EPC<29>/FFX/RST )
  );
  defparam DLX_reg_dst_of_MEM_0.INIT = 1'b0;
  X_SFF DLX_reg_dst_of_MEM_0 (
    .I(\DLX_reg_dst_of_MEM<1>/GROM ),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_reg_dst_of_MEM[0])
  );
  defparam DLX_IDinst_counter_1.INIT = 1'b0;
  X_FF DLX_IDinst_counter_1 (
    .I(DLX_IDinst__n0116[1]),
    .CE(DLX_IDinst__n0440),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_counter<1>/FFY/RST ),
    .O(DLX_IDinst_counter[1])
  );
  X_OR2 \DLX_IDinst_counter<1>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_counter<1>/FFY/RST )
  );
  defparam DLX_reg_dst_of_MEM_2.INIT = 1'b0;
  X_SFF DLX_reg_dst_of_MEM_2 (
    .I(\DLX_reg_dst_of_MEM<3>/GROM ),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_reg_dst_of_MEM[2])
  );
  defparam DLX_reg_dst_of_MEM_1.INIT = 1'b0;
  X_SFF DLX_reg_dst_of_MEM_1 (
    .I(\DLX_reg_dst_of_MEM<1>/FROM ),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_reg_dst_of_MEM[1])
  );
  defparam DLX_EXinst_reg_out_B_EX_19.INIT = 1'b0;
  X_FF DLX_EXinst_reg_out_B_EX_19 (
    .I(DLX_EXinst__n0007[19]),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_reg_out_B_EX<19>/FFX/RST ),
    .O(DLX_EXinst_reg_out_B_EX[19])
  );
  X_OR2 \DLX_EXinst_reg_out_B_EX<19>/FFX/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_reg_out_B_EX<19>/FFX/RST )
  );
  defparam DLX_EXinst_reg_out_B_EX_26.INIT = 1'b0;
  X_FF DLX_EXinst_reg_out_B_EX_26 (
    .I(DLX_EXinst__n0007[26]),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_reg_out_B_EX<27>/FFY/RST ),
    .O(DLX_EXinst_reg_out_B_EX[26])
  );
  X_OR2 \DLX_EXinst_reg_out_B_EX<27>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_reg_out_B_EX<27>/FFY/RST )
  );
  defparam DLX_EXinst_reg_out_B_EX_27.INIT = 1'b0;
  X_FF DLX_EXinst_reg_out_B_EX_27 (
    .I(DLX_EXinst__n0007[27]),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_reg_out_B_EX<27>/FFX/RST ),
    .O(DLX_EXinst_reg_out_B_EX[27])
  );
  X_OR2 \DLX_EXinst_reg_out_B_EX<27>/FFX/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_reg_out_B_EX<27>/FFX/RST )
  );
  defparam DLX_IDinst_IR_function_field_2_1_1193.INIT = 1'b0;
  X_FF DLX_IDinst_IR_function_field_2_1_1193 (
    .I(\DLX_IDinst_IR_function_field<2>/GROM ),
    .CE(DLX_IDinst__n0422),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_IR_function_field<2>/FFY/RST ),
    .O(DLX_IDinst_IR_function_field_2_1)
  );
  X_OR2 \DLX_IDinst_IR_function_field<2>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_IR_function_field<2>/FFY/RST )
  );
  defparam DLX_EXinst_reg_out_B_EX_28.INIT = 1'b0;
  X_FF DLX_EXinst_reg_out_B_EX_28 (
    .I(DLX_EXinst__n0007[28]),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_reg_out_B_EX<29>/FFY/RST ),
    .O(DLX_EXinst_reg_out_B_EX[28])
  );
  X_OR2 \DLX_EXinst_reg_out_B_EX<29>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_reg_out_B_EX<29>/FFY/RST )
  );
  defparam DLX_EXinst_reg_out_B_EX_29.INIT = 1'b0;
  X_FF DLX_EXinst_reg_out_B_EX_29 (
    .I(DLX_EXinst__n0007[29]),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_reg_out_B_EX<29>/FFX/RST ),
    .O(DLX_EXinst_reg_out_B_EX[29])
  );
  X_OR2 \DLX_EXinst_reg_out_B_EX<29>/FFX/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_reg_out_B_EX<29>/FFX/RST )
  );
  defparam DLX_IDinst_IR_function_field_2.INIT = 1'b0;
  X_FF DLX_IDinst_IR_function_field_2 (
    .I(DLX_IDinst__n0103),
    .CE(DLX_IDinst__n0422),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_IR_function_field<2>/FFX/RST ),
    .O(DLX_IDinst_IR_function_field[2])
  );
  X_OR2 \DLX_IDinst_IR_function_field<2>/FFX/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_IR_function_field<2>/FFX/RST )
  );
  defparam DLX_IDinst_IR_function_field_3_1_1194.INIT = 1'b0;
  X_FF DLX_IDinst_IR_function_field_3_1_1194 (
    .I(\DLX_IDinst_IR_function_field<3>/GROM ),
    .CE(DLX_IDinst__n0422),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_IR_function_field<3>/FFY/RST ),
    .O(DLX_IDinst_IR_function_field_3_1)
  );
  X_OR2 \DLX_IDinst_IR_function_field<3>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_IR_function_field<3>/FFY/RST )
  );
  defparam DLX_IDinst_reg_out_B_20.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_B_20 (
    .I(DLX_IDinst__n0118[20]),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_B<21>/FFY/RST ),
    .O(DLX_IDinst_reg_out_B[20])
  );
  X_OR2 \DLX_IDinst_reg_out_B<21>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_B<21>/FFY/RST )
  );
  defparam DLX_IDinst_reg_out_B_10.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_B_10 (
    .I(DLX_IDinst__n0118[10]),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_B<11>/FFY/RST ),
    .O(DLX_IDinst_reg_out_B[10])
  );
  X_OR2 \DLX_IDinst_reg_out_B<11>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_B<11>/FFY/RST )
  );
  defparam DLX_IDinst_IR_function_field_3.INIT = 1'b0;
  X_FF DLX_IDinst_IR_function_field_3 (
    .I(DLX_IDinst__n0102),
    .CE(DLX_IDinst__n0422),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_IR_function_field<3>/FFX/RST ),
    .O(DLX_IDinst_IR_function_field[3])
  );
  X_OR2 \DLX_IDinst_IR_function_field<3>/FFX/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_IR_function_field<3>/FFX/RST )
  );
  defparam DLX_EXinst_reg_out_B_EX_23.INIT = 1'b0;
  X_FF DLX_EXinst_reg_out_B_EX_23 (
    .I(DLX_EXinst__n0007[23]),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_reg_out_B_EX<23>/FFX/RST ),
    .O(DLX_EXinst_reg_out_B_EX[23])
  );
  X_OR2 \DLX_EXinst_reg_out_B_EX<23>/FFX/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_reg_out_B_EX<23>/FFX/RST )
  );
  defparam DLX_EXinst_reg_out_B_EX_14.INIT = 1'b0;
  X_FF DLX_EXinst_reg_out_B_EX_14 (
    .I(DLX_EXinst__n0007[14]),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_reg_out_B_EX<14>/FFY/RST ),
    .O(DLX_EXinst_reg_out_B_EX[14])
  );
  X_OR2 \DLX_EXinst_reg_out_B_EX<14>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_reg_out_B_EX<14>/FFY/RST )
  );
  defparam DLX_EXinst_reg_out_B_EX_25.INIT = 1'b0;
  X_FF DLX_EXinst_reg_out_B_EX_25 (
    .I(DLX_EXinst__n0007[25]),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_reg_out_B_EX<25>/FFX/RST ),
    .O(DLX_EXinst_reg_out_B_EX[25])
  );
  X_OR2 \DLX_EXinst_reg_out_B_EX<25>/FFX/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_reg_out_B_EX<25>/FFX/RST )
  );
  defparam DLX_IDinst_IR_function_field_1_1_1195.INIT = 1'b0;
  X_FF DLX_IDinst_IR_function_field_1_1_1195 (
    .I(\DLX_IDinst_IR_function_field<1>/GROM ),
    .CE(DLX_IDinst__n0422),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_IR_function_field<1>/FFY/RST ),
    .O(DLX_IDinst_IR_function_field_1_1)
  );
  X_OR2 \DLX_IDinst_IR_function_field<1>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_IR_function_field<1>/FFY/RST )
  );
  defparam DLX_EXinst_reg_out_B_EX_24.INIT = 1'b0;
  X_FF DLX_EXinst_reg_out_B_EX_24 (
    .I(DLX_EXinst__n0007[24]),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_reg_out_B_EX<25>/FFY/RST ),
    .O(DLX_EXinst_reg_out_B_EX[24])
  );
  X_OR2 \DLX_EXinst_reg_out_B_EX<25>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_reg_out_B_EX<25>/FFY/RST )
  );
  defparam DLX_IDinst_IR_function_field_1.INIT = 1'b0;
  X_FF DLX_IDinst_IR_function_field_1 (
    .I(DLX_IDinst__n0104),
    .CE(DLX_IDinst__n0422),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_IR_function_field<1>/FFX/RST ),
    .O(DLX_IDinst_IR_function_field[1])
  );
  X_OR2 \DLX_IDinst_IR_function_field<1>/FFX/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_IR_function_field<1>/FFX/RST )
  );
  defparam DLX_EXinst_reg_out_B_EX_16.INIT = 1'b0;
  X_FF DLX_EXinst_reg_out_B_EX_16 (
    .I(DLX_EXinst__n0007[16]),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_reg_out_B_EX<17>/FFY/RST ),
    .O(DLX_EXinst_reg_out_B_EX[16])
  );
  X_OR2 \DLX_EXinst_reg_out_B_EX<17>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_reg_out_B_EX<17>/FFY/RST )
  );
  defparam DLX_EXinst_reg_out_B_EX_17.INIT = 1'b0;
  X_FF DLX_EXinst_reg_out_B_EX_17 (
    .I(DLX_EXinst__n0007[17]),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_reg_out_B_EX<17>/FFX/RST ),
    .O(DLX_EXinst_reg_out_B_EX[17])
  );
  X_OR2 \DLX_EXinst_reg_out_B_EX<17>/FFX/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_reg_out_B_EX<17>/FFX/RST )
  );
  defparam DLX_EXinst_reg_out_B_EX_18.INIT = 1'b0;
  X_FF DLX_EXinst_reg_out_B_EX_18 (
    .I(DLX_EXinst__n0007[18]),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_reg_out_B_EX<19>/FFY/RST ),
    .O(DLX_EXinst_reg_out_B_EX[18])
  );
  X_OR2 \DLX_EXinst_reg_out_B_EX<19>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_reg_out_B_EX<19>/FFY/RST )
  );
  defparam DLX_IDinst_reg_out_B_29.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_B_29 (
    .I(DLX_IDinst__n0118[29]),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_B<29>/FFX/RST ),
    .O(DLX_IDinst_reg_out_B[29])
  );
  X_OR2 \DLX_IDinst_reg_out_B<29>/FFX/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_B<29>/FFX/RST )
  );
  defparam DLX_IDinst_Imm_7.INIT = 1'b0;
  X_FF DLX_IDinst_Imm_7 (
    .I(DLX_IDinst__n0098),
    .CE(DLX_IDinst__n0422),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_Imm<8>/FFY/RST ),
    .O(\DLX_IDinst_Imm[7] )
  );
  X_OR2 \DLX_IDinst_Imm<8>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_Imm<8>/FFY/RST )
  );
  defparam DLX_EXinst_ALU_result_2.INIT = 1'b0;
  X_FF DLX_EXinst_ALU_result_2 (
    .I(\DLX_EXinst_ALU_result<2>/GROM ),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_ALU_result<2>/FFY/RST ),
    .O(DLX_EXinst_ALU_result[2])
  );
  X_OR2 \DLX_EXinst_ALU_result<2>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_ALU_result<2>/FFY/RST )
  );
  defparam DLX_IDinst_Imm_6.INIT = 1'b0;
  X_FF DLX_IDinst_Imm_6 (
    .I(DLX_IDinst__n0099),
    .CE(DLX_IDinst__n0422),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_IR_opcode_field<2>/FFY/RST ),
    .O(\DLX_IDinst_Imm[6] )
  );
  X_OR2 \DLX_IDinst_IR_opcode_field<2>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_IR_opcode_field<2>/FFY/RST )
  );
  defparam DLX_IDinst_IR_opcode_field_2.INIT = 1'b0;
  X_FF DLX_IDinst_IR_opcode_field_2 (
    .I(DLX_IDinst__n0113[2]),
    .CE(DLX_IDinst__n0422),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_IR_opcode_field<2>/FFX/RST ),
    .O(DLX_IDinst_IR_opcode_field[2])
  );
  X_OR2 \DLX_IDinst_IR_opcode_field<2>/FFX/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_IR_opcode_field<2>/FFX/RST )
  );
  defparam DLX_MEMinst_RF_data_in_1.INIT = 1'b0;
  X_FF DLX_MEMinst_RF_data_in_1 (
    .I(DLX_MEMinst__n0000[1]),
    .CE(VCC),
    .CLK(\DLX_RF_data_in<1>/CKMUXNOT ),
    .SET(GND),
    .RST(\DLX_RF_data_in<1>/FFX/RST ),
    .O(DLX_RF_data_in[1])
  );
  X_OR2 \DLX_RF_data_in<1>/FFX/RSTOR  (
    .I0(reset_IBUF_1),
    .I1(GSR),
    .O(\DLX_RF_data_in<1>/FFX/RST )
  );
  defparam DLX_IDinst_Imm_8.INIT = 1'b0;
  X_FF DLX_IDinst_Imm_8 (
    .I(DLX_IDinst__n0097),
    .CE(DLX_IDinst__n0422),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_Imm<8>/FFX/RST ),
    .O(\DLX_IDinst_Imm[8] )
  );
  X_OR2 \DLX_IDinst_Imm<8>/FFX/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_Imm<8>/FFX/RST )
  );
  defparam DLX_MEMinst_RF_data_in_2.INIT = 1'b0;
  X_FF DLX_MEMinst_RF_data_in_2 (
    .I(DLX_MEMinst__n0000[2]),
    .CE(VCC),
    .CLK(\DLX_RF_data_in<3>/CKMUXNOT ),
    .SET(GND),
    .RST(\DLX_RF_data_in<3>/FFY/RST ),
    .O(DLX_RF_data_in[2])
  );
  X_OR2 \DLX_RF_data_in<3>/FFY/RSTOR  (
    .I0(reset_IBUF_1),
    .I1(GSR),
    .O(\DLX_RF_data_in<3>/FFY/RST )
  );
  defparam DLX_MEMinst_RF_data_in_0.INIT = 1'b0;
  X_FF DLX_MEMinst_RF_data_in_0 (
    .I(DLX_MEMinst__n0000[0]),
    .CE(VCC),
    .CLK(\DLX_RF_data_in<1>/CKMUXNOT ),
    .SET(GND),
    .RST(\DLX_RF_data_in<1>/FFY/RST ),
    .O(DLX_RF_data_in[0])
  );
  X_OR2 \DLX_RF_data_in<1>/FFY/RSTOR  (
    .I0(reset_IBUF_1),
    .I1(GSR),
    .O(\DLX_RF_data_in<1>/FFY/RST )
  );
  defparam DLX_IDinst_Imm_9.INIT = 1'b0;
  X_FF DLX_IDinst_Imm_9 (
    .I(DLX_IDinst__n0096),
    .CE(DLX_IDinst__n0422),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_Imm<10>/FFY/RST ),
    .O(\DLX_IDinst_Imm[9] )
  );
  X_OR2 \DLX_IDinst_Imm<10>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_Imm<10>/FFY/RST )
  );
  defparam DLX_IDinst_reg_out_B_15.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_B_15 (
    .I(DLX_IDinst__n0118[15]),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_B<15>/FFX/RST ),
    .O(DLX_IDinst_reg_out_B[15])
  );
  X_OR2 \DLX_IDinst_reg_out_B<15>/FFX/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_B<15>/FFX/RST )
  );
  defparam DLX_IDinst_reg_out_B_24.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_B_24 (
    .I(DLX_IDinst__n0118[24]),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_B<25>/FFY/RST ),
    .O(DLX_IDinst_reg_out_B[24])
  );
  X_OR2 \DLX_IDinst_reg_out_B<25>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_B<25>/FFY/RST )
  );
  defparam DLX_IDinst_reg_out_B_25.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_B_25 (
    .I(DLX_IDinst__n0118[25]),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_B<25>/FFX/RST ),
    .O(DLX_IDinst_reg_out_B[25])
  );
  X_OR2 \DLX_IDinst_reg_out_B<25>/FFX/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_B<25>/FFX/RST )
  );
  defparam DLX_IDinst_reg_out_B_16.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_B_16 (
    .I(DLX_IDinst__n0118[16]),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_B<17>/FFY/RST ),
    .O(DLX_IDinst_reg_out_B[16])
  );
  X_OR2 \DLX_IDinst_reg_out_B<17>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_B<17>/FFY/RST )
  );
  defparam DLX_IDinst_reg_out_B_17.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_B_17 (
    .I(DLX_IDinst__n0118[17]),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_B<17>/FFX/RST ),
    .O(DLX_IDinst_reg_out_B[17])
  );
  X_OR2 \DLX_IDinst_reg_out_B<17>/FFX/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_B<17>/FFX/RST )
  );
  defparam DLX_IDinst_reg_out_B_26.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_B_26 (
    .I(DLX_IDinst__n0118[26]),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_B<27>/FFY/RST ),
    .O(DLX_IDinst_reg_out_B[26])
  );
  X_OR2 \DLX_IDinst_reg_out_B<27>/FFY/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_B<27>/FFY/RST )
  );
  defparam DLX_IDinst_reg_out_B_27.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_B_27 (
    .I(DLX_IDinst__n0118[27]),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_B<27>/FFX/RST ),
    .O(DLX_IDinst_reg_out_B[27])
  );
  X_OR2 \DLX_IDinst_reg_out_B<27>/FFX/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_B<27>/FFX/RST )
  );
  defparam DLX_IDinst_reg_out_B_18.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_B_18 (
    .I(DLX_IDinst__n0118[18]),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_B<19>/FFY/RST ),
    .O(DLX_IDinst_reg_out_B[18])
  );
  X_OR2 \DLX_IDinst_reg_out_B<19>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_B<19>/FFY/RST )
  );
  defparam DLX_IDinst_reg_out_B_28.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_B_28 (
    .I(DLX_IDinst__n0118[28]),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_B<29>/FFY/RST ),
    .O(DLX_IDinst_reg_out_B[28])
  );
  X_OR2 \DLX_IDinst_reg_out_B<29>/FFY/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_B<29>/FFY/RST )
  );
  defparam DLX_IDinst_reg_out_B_19.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_B_19 (
    .I(DLX_IDinst__n0118[19]),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_B<19>/FFX/RST ),
    .O(DLX_IDinst_reg_out_B[19])
  );
  X_OR2 \DLX_IDinst_reg_out_B<19>/FFX/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_B<19>/FFX/RST )
  );
  defparam DLX_IDinst_Imm_10.INIT = 1'b0;
  X_FF DLX_IDinst_Imm_10 (
    .I(DLX_IDinst__n0095),
    .CE(DLX_IDinst__n0422),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_Imm<10>/FFX/RST ),
    .O(\DLX_IDinst_Imm[10] )
  );
  X_OR2 \DLX_IDinst_Imm<10>/FFX/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_Imm<10>/FFX/RST )
  );
  defparam DLX_MEMinst_RF_data_in_3.INIT = 1'b0;
  X_FF DLX_MEMinst_RF_data_in_3 (
    .I(DLX_MEMinst__n0000[3]),
    .CE(VCC),
    .CLK(\DLX_RF_data_in<3>/CKMUXNOT ),
    .SET(GND),
    .RST(\DLX_RF_data_in<3>/FFX/RST ),
    .O(DLX_RF_data_in[3])
  );
  X_OR2 \DLX_RF_data_in<3>/FFX/RSTOR  (
    .I0(reset_IBUF_1),
    .I1(GSR),
    .O(\DLX_RF_data_in<3>/FFX/RST )
  );
  defparam DLX_MEMinst_RF_data_in_4.INIT = 1'b0;
  X_FF DLX_MEMinst_RF_data_in_4 (
    .I(DLX_MEMinst__n0000[4]),
    .CE(VCC),
    .CLK(\DLX_RF_data_in<5>/CKMUXNOT ),
    .SET(GND),
    .RST(\DLX_RF_data_in<5>/FFY/RST ),
    .O(DLX_RF_data_in[4])
  );
  X_OR2 \DLX_RF_data_in<5>/FFY/RSTOR  (
    .I0(reset_IBUF_1),
    .I1(GSR),
    .O(\DLX_RF_data_in<5>/FFY/RST )
  );
  defparam DLX_MEMinst_RF_data_in_5.INIT = 1'b0;
  X_FF DLX_MEMinst_RF_data_in_5 (
    .I(DLX_MEMinst__n0000[5]),
    .CE(VCC),
    .CLK(\DLX_RF_data_in<5>/CKMUXNOT ),
    .SET(GND),
    .RST(\DLX_RF_data_in<5>/FFX/RST ),
    .O(DLX_RF_data_in[5])
  );
  X_OR2 \DLX_RF_data_in<5>/FFX/RSTOR  (
    .I0(reset_IBUF_1),
    .I1(GSR),
    .O(\DLX_RF_data_in<5>/FFX/RST )
  );
  defparam DLX_MEMinst_RF_data_in_6.INIT = 1'b0;
  X_FF DLX_MEMinst_RF_data_in_6 (
    .I(DLX_MEMinst__n0000[6]),
    .CE(VCC),
    .CLK(\DLX_RF_data_in<7>/CKMUXNOT ),
    .SET(GND),
    .RST(\DLX_RF_data_in<7>/FFY/RST ),
    .O(DLX_RF_data_in[6])
  );
  X_OR2 \DLX_RF_data_in<7>/FFY/RSTOR  (
    .I0(reset_IBUF_1),
    .I1(GSR),
    .O(\DLX_RF_data_in<7>/FFY/RST )
  );
  defparam DLX_MEMinst_RF_data_in_7.INIT = 1'b0;
  X_FF DLX_MEMinst_RF_data_in_7 (
    .I(DLX_MEMinst__n0000[7]),
    .CE(VCC),
    .CLK(\DLX_RF_data_in<7>/CKMUXNOT ),
    .SET(GND),
    .RST(\DLX_RF_data_in<7>/FFX/RST ),
    .O(DLX_RF_data_in[7])
  );
  X_OR2 \DLX_RF_data_in<7>/FFX/RSTOR  (
    .I0(reset_IBUF_1),
    .I1(GSR),
    .O(\DLX_RF_data_in<7>/FFX/RST )
  );
  defparam DLX_MEMinst_RF_data_in_8.INIT = 1'b0;
  X_FF DLX_MEMinst_RF_data_in_8 (
    .I(DLX_MEMinst__n0000[8]),
    .CE(VCC),
    .CLK(\DLX_MEMinst_RF_data_in<9>/CKMUXNOT ),
    .SET(GND),
    .RST(\DLX_MEMinst_RF_data_in<9>/FFY/RST ),
    .O(DLX_MEMinst_RF_data_in[8])
  );
  X_OR2 \DLX_MEMinst_RF_data_in<9>/FFY/RSTOR  (
    .I0(reset_IBUF_1),
    .I1(GSR),
    .O(\DLX_MEMinst_RF_data_in<9>/FFY/RST )
  );
  defparam DLX_MEMinst_RF_data_in_9.INIT = 1'b0;
  X_FF DLX_MEMinst_RF_data_in_9 (
    .I(DLX_MEMinst__n0000[9]),
    .CE(VCC),
    .CLK(\DLX_MEMinst_RF_data_in<9>/CKMUXNOT ),
    .SET(GND),
    .RST(\DLX_MEMinst_RF_data_in<9>/FFX/RST ),
    .O(DLX_MEMinst_RF_data_in[9])
  );
  X_OR2 \DLX_MEMinst_RF_data_in<9>/FFX/RSTOR  (
    .I0(reset_IBUF_1),
    .I1(GSR),
    .O(\DLX_MEMinst_RF_data_in<9>/FFX/RST )
  );
  defparam DLX_EXinst_byte_1196.INIT = 1'b0;
  X_FF DLX_EXinst_byte_1196 (
    .I(DLX_EXinst__n0014),
    .CE(DLX_EXinst__n0149),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_word/FFY/RST ),
    .O(DLX_EXinst_byte)
  );
  X_OR2 \DLX_EXinst_word/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_word/FFY/RST )
  );
  defparam DLX_IDinst_reg_out_B_5.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_B_5 (
    .I(DLX_IDinst__n0118[5]),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_B<5>/FFX/RST ),
    .O(DLX_IDinst_reg_out_B[5])
  );
  X_OR2 \DLX_IDinst_reg_out_B<5>/FFX/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_B<5>/FFX/RST )
  );
  defparam DLX_IDinst_reg_out_B_6.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_B_6 (
    .I(DLX_IDinst__n0118[6]),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_B<7>/FFY/RST ),
    .O(DLX_IDinst_reg_out_B[6])
  );
  X_OR2 \DLX_IDinst_reg_out_B<7>/FFY/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_B<7>/FFY/RST )
  );
  defparam DLX_IDinst_reg_out_B_7.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_B_7 (
    .I(DLX_IDinst__n0118[7]),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_B<7>/FFX/RST ),
    .O(DLX_IDinst_reg_out_B[7])
  );
  X_OR2 \DLX_IDinst_reg_out_B<7>/FFX/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_B<7>/FFX/RST )
  );
  defparam DLX_IDinst_reg_out_B_8.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_B_8 (
    .I(DLX_IDinst__n0118[8]),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_B<9>/FFY/RST ),
    .O(DLX_IDinst_reg_out_B[8])
  );
  X_OR2 \DLX_IDinst_reg_out_B<9>/FFY/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_B<9>/FFY/RST )
  );
  defparam DLX_IDinst_reg_out_B_9.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_B_9 (
    .I(DLX_IDinst__n0118[9]),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_B<9>/FFX/RST ),
    .O(DLX_IDinst_reg_out_B[9])
  );
  X_OR2 \DLX_IDinst_reg_out_B<9>/FFX/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_B<9>/FFX/RST )
  );
  defparam DLX_IDinst_rt_addr_1.INIT = 1'b0;
  X_FF DLX_IDinst_rt_addr_1 (
    .I(DLX_IDinst__n0106[1]),
    .CE(DLX_IDinst__n0422),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_rt_addr<1>/FFY/RST ),
    .O(DLX_IDinst_rt_addr[1])
  );
  X_OR2 \DLX_IDinst_rt_addr<1>/FFY/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IDinst_rt_addr<1>/FFY/RST )
  );
  defparam DLX_IDinst_rt_addr_3.INIT = 1'b0;
  X_FF DLX_IDinst_rt_addr_3 (
    .I(DLX_IDinst__n0106[3]),
    .CE(DLX_IDinst__n0422),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_rt_addr<3>/FFX/RST ),
    .O(DLX_IDinst_rt_addr[3])
  );
  X_OR2 \DLX_IDinst_rt_addr<3>/FFX/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IDinst_rt_addr<3>/FFX/RST )
  );
  defparam DLX_IDinst_rt_addr_2.INIT = 1'b0;
  X_FF DLX_IDinst_rt_addr_2 (
    .I(DLX_IDinst__n0106[2]),
    .CE(DLX_IDinst__n0422),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_rt_addr<3>/FFY/RST ),
    .O(DLX_IDinst_rt_addr[2])
  );
  X_OR2 \DLX_IDinst_rt_addr<3>/FFY/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IDinst_rt_addr<3>/FFY/RST )
  );
  defparam DLX_IDinst_mem_read_1197.INIT = 1'b0;
  X_FF DLX_IDinst_mem_read_1197 (
    .I(DLX_IDinst__n0111),
    .CE(DLX_IDinst__n0422),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_mem_read/FFY/RST ),
    .O(DLX_IDinst_mem_read)
  );
  X_OR2 \DLX_IDinst_mem_read/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_mem_read/FFY/RST )
  );
  defparam DLX_IDinst_IR_opcode_field_5.INIT = 1'b0;
  X_FF DLX_IDinst_IR_opcode_field_5 (
    .I(DLX_IDinst__n0113[5]),
    .CE(DLX_IDinst__n0422),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_IR_opcode_field<5>/FFX/RST ),
    .O(DLX_IDinst_IR_opcode_field[5])
  );
  X_OR2 \DLX_IDinst_IR_opcode_field<5>/FFX/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_IR_opcode_field<5>/FFX/RST )
  );
  defparam DLX_EXinst_word_1198.INIT = 1'b0;
  X_FF DLX_EXinst_word_1198 (
    .I(DLX_EXinst__n0015),
    .CE(DLX_EXinst__n0149),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_word/FFX/RST ),
    .O(DLX_EXinst_word)
  );
  X_OR2 \DLX_EXinst_word/FFX/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_word/FFX/RST )
  );
  defparam DLX_IFinst_stalled_1199.INIT = 1'b0;
  X_FF DLX_IFinst_stalled_1199 (
    .I(\DLX_IFinst_stalled/GROM ),
    .CE(\DLX_IFinst_stalled/CEMUXNOT ),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_stalled/FFY/RST ),
    .O(DLX_IFinst_stalled)
  );
  X_OR2 \DLX_IFinst_stalled/FFY/RSTOR  (
    .I0(reset_IBUF_1),
    .I1(GSR),
    .O(\DLX_IFinst_stalled/FFY/RST )
  );
  defparam DLX_IDinst_rd_addr_3.INIT = 1'b0;
  X_FF DLX_IDinst_rd_addr_3 (
    .I(DLX_IDinst__n0107[3]),
    .CE(DLX_IDinst__n0422),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_rd_addr<3>/FFX/RST ),
    .O(DLX_IDinst_rd_addr[3])
  );
  X_OR2 \DLX_IDinst_rd_addr<3>/FFX/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_rd_addr<3>/FFX/RST )
  );
  defparam DLX_IDinst_rd_addr_1.INIT = 1'b0;
  X_FF DLX_IDinst_rd_addr_1 (
    .I(DLX_IDinst__n0107[1]),
    .CE(DLX_IDinst__n0422),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_rd_addr<4>/FFY/RST ),
    .O(DLX_IDinst_rd_addr[1])
  );
  X_OR2 \DLX_IDinst_rd_addr<4>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_rd_addr<4>/FFY/RST )
  );
  defparam DLX_IDinst_rd_addr_4.INIT = 1'b0;
  X_FF DLX_IDinst_rd_addr_4 (
    .I(DLX_IDinst__n0107[4]),
    .CE(DLX_IDinst__n0422),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_rd_addr<4>/FFX/RST ),
    .O(DLX_IDinst_rd_addr[4])
  );
  X_OR2 \DLX_IDinst_rd_addr<4>/FFX/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_rd_addr<4>/FFX/RST )
  );
  defparam DLX_IDinst_rd_addr_2.INIT = 1'b0;
  X_FF DLX_IDinst_rd_addr_2 (
    .I(DLX_IDinst__n0107[2]),
    .CE(DLX_IDinst__n0422),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_rd_addr<3>/FFY/RST ),
    .O(DLX_IDinst_rd_addr[2])
  );
  X_OR2 \DLX_IDinst_rd_addr<3>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_rd_addr<3>/FFY/RST )
  );
  defparam DLX_IDinst_reg_out_B_4.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_B_4 (
    .I(DLX_IDinst__n0118[4]),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_B<5>/FFY/RST ),
    .O(DLX_IDinst_reg_out_B[4])
  );
  X_OR2 \DLX_IDinst_reg_out_B<5>/FFY/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_B<5>/FFY/RST )
  );
  defparam DLX_IDinst_reg_out_B_1.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_B_1 (
    .I(DLX_IDinst__n0118[1]),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_B<1>/FFY/RST ),
    .O(DLX_IDinst_reg_out_B[1])
  );
  X_OR2 \DLX_IDinst_reg_out_B<1>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_B<1>/FFY/RST )
  );
  defparam DLX_IDinst_Cause_Reg_10.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_10 (
    .I(DLX_IDinst__n0127[10]),
    .CE(DLX_IDinst__n0085),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<11>/FFY/RST ),
    .O(DLX_IDinst_Cause_Reg[10])
  );
  X_BUF \DLX_IDinst_Cause_Reg<11>/FFY/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<11>/FFY/RST )
  );
  defparam DLX_IDinst_Cause_Reg_11.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_11 (
    .I(DLX_IDinst__n0127[11]),
    .CE(DLX_IDinst__n0085),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<11>/FFX/RST ),
    .O(DLX_IDinst_Cause_Reg[11])
  );
  X_BUF \DLX_IDinst_Cause_Reg<11>/FFX/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<11>/FFX/RST )
  );
  defparam DLX_IDinst_Cause_Reg_12.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_12 (
    .I(DLX_IDinst__n0127[12]),
    .CE(DLX_IDinst__n0085),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<13>/FFY/RST ),
    .O(DLX_IDinst_Cause_Reg[12])
  );
  X_BUF \DLX_IDinst_Cause_Reg<13>/FFY/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<13>/FFY/RST )
  );
  defparam DLX_IDinst_Cause_Reg_13.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_13 (
    .I(DLX_IDinst__n0127[13]),
    .CE(DLX_IDinst__n0085),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<13>/FFX/RST ),
    .O(DLX_IDinst_Cause_Reg[13])
  );
  X_BUF \DLX_IDinst_Cause_Reg<13>/FFX/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<13>/FFX/RST )
  );
  defparam DLX_IDinst_Cause_Reg_20.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_20 (
    .I(DLX_IDinst__n0127[20]),
    .CE(DLX_IDinst__n0085),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<21>/FFY/RST ),
    .O(DLX_IDinst_Cause_Reg[20])
  );
  X_BUF \DLX_IDinst_Cause_Reg<21>/FFY/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<21>/FFY/RST )
  );
  defparam DLX_IDinst_Cause_Reg_21.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_21 (
    .I(DLX_IDinst__n0127[21]),
    .CE(DLX_IDinst__n0085),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<21>/FFX/RST ),
    .O(DLX_IDinst_Cause_Reg[21])
  );
  X_BUF \DLX_IDinst_Cause_Reg<21>/FFX/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<21>/FFX/RST )
  );
  defparam DLX_IDinst_mem_write_1200.INIT = 1'b0;
  X_FF DLX_IDinst_mem_write_1200 (
    .I(DLX_IDinst__n0112),
    .CE(DLX_IDinst__n0422),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_mem_write/FFY/RST ),
    .O(DLX_IDinst_mem_write)
  );
  X_OR2 \DLX_IDinst_mem_write/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_mem_write/FFY/RST )
  );
  defparam DLX_IDinst_Cause_Reg_14.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_14 (
    .I(DLX_IDinst__n0127[14]),
    .CE(DLX_IDinst__n0085),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<15>/FFY/RST ),
    .O(DLX_IDinst_Cause_Reg[14])
  );
  X_BUF \DLX_IDinst_Cause_Reg<15>/FFY/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<15>/FFY/RST )
  );
  defparam DLX_IDinst_Cause_Reg_15.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_15 (
    .I(DLX_IDinst__n0127[15]),
    .CE(DLX_IDinst__n0085),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<15>/FFX/RST ),
    .O(DLX_IDinst_Cause_Reg[15])
  );
  X_BUF \DLX_IDinst_Cause_Reg<15>/FFX/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<15>/FFX/RST )
  );
  defparam DLX_IDinst_Cause_Reg_22.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_22 (
    .I(DLX_IDinst__n0127[22]),
    .CE(DLX_IDinst__n0085),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<23>/FFY/RST ),
    .O(DLX_IDinst_Cause_Reg[22])
  );
  X_BUF \DLX_IDinst_Cause_Reg<23>/FFY/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<23>/FFY/RST )
  );
  defparam DLX_IDinst_Cause_Reg_23.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_23 (
    .I(DLX_IDinst__n0127[23]),
    .CE(DLX_IDinst__n0085),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<23>/FFX/RST ),
    .O(DLX_IDinst_Cause_Reg[23])
  );
  X_BUF \DLX_IDinst_Cause_Reg<23>/FFX/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<23>/FFX/RST )
  );
  defparam DLX_IDinst_Cause_Reg_30.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_30 (
    .I(DLX_IDinst__n0127[30]),
    .CE(DLX_IDinst__n0085),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<31>/FFY/RST ),
    .O(DLX_IDinst_Cause_Reg[30])
  );
  X_BUF \DLX_IDinst_Cause_Reg<31>/FFY/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<31>/FFY/RST )
  );
  defparam DLX_IDinst_Cause_Reg_31.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_31 (
    .I(DLX_IDinst__n0127[31]),
    .CE(DLX_IDinst__n0085),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<31>/FFX/RST ),
    .O(DLX_IDinst_Cause_Reg[31])
  );
  X_BUF \DLX_IDinst_Cause_Reg<31>/FFX/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<31>/FFX/RST )
  );
  defparam DLX_IDinst_Cause_Reg_16.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_16 (
    .I(DLX_IDinst__n0127[16]),
    .CE(DLX_IDinst__n0085),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<17>/FFY/RST ),
    .O(DLX_IDinst_Cause_Reg[16])
  );
  X_BUF \DLX_IDinst_Cause_Reg<17>/FFY/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<17>/FFY/RST )
  );
  defparam DLX_IDinst_Cause_Reg_17.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_17 (
    .I(DLX_IDinst__n0127[17]),
    .CE(DLX_IDinst__n0085),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<17>/FFX/RST ),
    .O(DLX_IDinst_Cause_Reg[17])
  );
  X_BUF \DLX_IDinst_Cause_Reg<17>/FFX/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<17>/FFX/RST )
  );
  defparam DLX_IDinst_Cause_Reg_24.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_24 (
    .I(DLX_IDinst__n0127[24]),
    .CE(DLX_IDinst__n0085),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<25>/FFY/RST ),
    .O(DLX_IDinst_Cause_Reg[24])
  );
  X_BUF \DLX_IDinst_Cause_Reg<25>/FFY/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<25>/FFY/RST )
  );
  defparam DLX_IDinst_Cause_Reg_25.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_25 (
    .I(DLX_IDinst__n0127[25]),
    .CE(DLX_IDinst__n0085),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<25>/FFX/RST ),
    .O(DLX_IDinst_Cause_Reg[25])
  );
  X_BUF \DLX_IDinst_Cause_Reg<25>/FFX/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<25>/FFX/RST )
  );
  defparam DLX_IDinst_Cause_Reg_18.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_18 (
    .I(DLX_IDinst__n0127[18]),
    .CE(DLX_IDinst__n0085),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<19>/FFY/RST ),
    .O(DLX_IDinst_Cause_Reg[18])
  );
  X_BUF \DLX_IDinst_Cause_Reg<19>/FFY/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<19>/FFY/RST )
  );
  defparam DLX_IDinst_Cause_Reg_19.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_19 (
    .I(DLX_IDinst__n0127[19]),
    .CE(DLX_IDinst__n0085),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<19>/FFX/RST ),
    .O(DLX_IDinst_Cause_Reg[19])
  );
  X_BUF \DLX_IDinst_Cause_Reg<19>/FFX/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<19>/FFX/RST )
  );
  defparam DLX_IDinst_Cause_Reg_26.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_26 (
    .I(DLX_IDinst__n0127[26]),
    .CE(DLX_IDinst__n0085),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<27>/FFY/RST ),
    .O(DLX_IDinst_Cause_Reg[26])
  );
  X_BUF \DLX_IDinst_Cause_Reg<27>/FFY/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<27>/FFY/RST )
  );
  defparam DLX_IDinst_Cause_Reg_27.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_27 (
    .I(DLX_IDinst__n0127[27]),
    .CE(DLX_IDinst__n0085),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<27>/FFX/RST ),
    .O(DLX_IDinst_Cause_Reg[27])
  );
  X_BUF \DLX_IDinst_Cause_Reg<27>/FFX/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<27>/FFX/RST )
  );
  defparam DLX_IDinst_Cause_Reg_28.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_28 (
    .I(DLX_IDinst__n0127[28]),
    .CE(DLX_IDinst__n0085),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<29>/FFY/RST ),
    .O(DLX_IDinst_Cause_Reg[28])
  );
  X_BUF \DLX_IDinst_Cause_Reg<29>/FFY/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<29>/FFY/RST )
  );
  defparam DLX_EXinst_reg_out_B_EX_5.INIT = 1'b0;
  X_FF DLX_EXinst_reg_out_B_EX_5 (
    .I(DLX_EXinst__n0007[5]),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_reg_out_B_EX<5>/FFX/RST ),
    .O(DLX_EXinst_reg_out_B_EX[5])
  );
  X_OR2 \DLX_EXinst_reg_out_B_EX<5>/FFX/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_reg_out_B_EX<5>/FFX/RST )
  );
  defparam DLX_EXinst_reg_out_B_EX_2.INIT = 1'b0;
  X_FF DLX_EXinst_reg_out_B_EX_2 (
    .I(DLX_EXinst__n0007[2]),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_reg_out_B_EX<3>/FFY/RST ),
    .O(DLX_EXinst_reg_out_B_EX[2])
  );
  X_OR2 \DLX_EXinst_reg_out_B_EX<3>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_reg_out_B_EX<3>/FFY/RST )
  );
  defparam DLX_IDinst_Cause_Reg_29.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_29 (
    .I(DLX_IDinst__n0127[29]),
    .CE(DLX_IDinst__n0085),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<29>/FFX/RST ),
    .O(DLX_IDinst_Cause_Reg[29])
  );
  X_BUF \DLX_IDinst_Cause_Reg<29>/FFX/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<29>/FFX/RST )
  );
  defparam DLX_EXinst_reg_out_B_EX_0.INIT = 1'b0;
  X_FF DLX_EXinst_reg_out_B_EX_0 (
    .I(\DLX_EXinst_reg_out_B_EX<1>/GROM ),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_reg_out_B_EX<1>/FFY/RST ),
    .O(DLX_EXinst_reg_out_B_EX[0])
  );
  X_OR2 \DLX_EXinst_reg_out_B_EX<1>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_reg_out_B_EX<1>/FFY/RST )
  );
  defparam DLX_EXinst_reg_out_B_EX_1.INIT = 1'b0;
  X_FF DLX_EXinst_reg_out_B_EX_1 (
    .I(DLX_EXinst__n0007[1]),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_reg_out_B_EX<1>/FFX/RST ),
    .O(DLX_EXinst_reg_out_B_EX[1])
  );
  X_OR2 \DLX_EXinst_reg_out_B_EX<1>/FFX/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_reg_out_B_EX<1>/FFX/RST )
  );
  defparam DLX_EXinst_reg_out_B_EX_3.INIT = 1'b0;
  X_FF DLX_EXinst_reg_out_B_EX_3 (
    .I(DLX_EXinst__n0007[3]),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_reg_out_B_EX<3>/FFX/RST ),
    .O(DLX_EXinst_reg_out_B_EX[3])
  );
  X_OR2 \DLX_EXinst_reg_out_B_EX<3>/FFX/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_reg_out_B_EX<3>/FFX/RST )
  );
  defparam DLX_EXinst_reg_out_B_EX_4.INIT = 1'b0;
  X_FF DLX_EXinst_reg_out_B_EX_4 (
    .I(DLX_EXinst__n0007[4]),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_reg_out_B_EX<5>/FFY/RST ),
    .O(DLX_EXinst_reg_out_B_EX[4])
  );
  X_OR2 \DLX_EXinst_reg_out_B_EX<5>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_reg_out_B_EX<5>/FFY/RST )
  );
  defparam DLX_EXinst_reg_out_B_EX_7.INIT = 1'b0;
  X_FF DLX_EXinst_reg_out_B_EX_7 (
    .I(DLX_EXinst__n0007[7]),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_reg_out_B_EX<7>/FFX/RST ),
    .O(DLX_EXinst_reg_out_B_EX[7])
  );
  X_OR2 \DLX_EXinst_reg_out_B_EX<7>/FFX/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_reg_out_B_EX<7>/FFX/RST )
  );
  defparam DLX_EXinst_reg_out_B_EX_6.INIT = 1'b0;
  X_FF DLX_EXinst_reg_out_B_EX_6 (
    .I(DLX_EXinst__n0007[6]),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_reg_out_B_EX<7>/FFY/RST ),
    .O(DLX_EXinst_reg_out_B_EX[6])
  );
  X_OR2 \DLX_EXinst_reg_out_B_EX<7>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_reg_out_B_EX<7>/FFY/RST )
  );
  defparam DLX_EXinst_reg_out_B_EX_8.INIT = 1'b0;
  X_FF DLX_EXinst_reg_out_B_EX_8 (
    .I(DLX_EXinst__n0007[8]),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_reg_out_B_EX<9>/FFY/RST ),
    .O(DLX_EXinst_reg_out_B_EX[8])
  );
  X_OR2 \DLX_EXinst_reg_out_B_EX<9>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_reg_out_B_EX<9>/FFY/RST )
  );
  defparam DLX_EXinst_reg_dst_out_0.INIT = 1'b0;
  X_FF DLX_EXinst_reg_dst_out_0 (
    .I(DLX_EXinst__n0008[0]),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_reg_dst_out<1>/FFY/RST ),
    .O(DLX_EXinst_reg_dst_out[0])
  );
  X_OR2 \DLX_EXinst_reg_dst_out<1>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_reg_dst_out<1>/FFY/RST )
  );
  defparam DLX_opcode_of_WB_0.INIT = 1'b0;
  X_SFF DLX_opcode_of_WB_0 (
    .I(DLX_opcode_of_MEM[0]),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_opcode_of_WB[0])
  );
  defparam DLX_opcode_of_WB_1.INIT = 1'b0;
  X_SFF DLX_opcode_of_WB_1 (
    .I(DLX_opcode_of_MEM[1]),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_opcode_of_WB[1])
  );
  defparam DLX_IDinst_reg_out_A_29.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_A_29 (
    .I(N104644),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_A<29>/FFY/RST ),
    .O(DLX_IDinst_reg_out_A[29])
  );
  X_OR2 \DLX_IDinst_reg_out_A<29>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_A<29>/FFY/RST )
  );
  defparam DLX_opcode_of_WB_2.INIT = 1'b0;
  X_SFF DLX_opcode_of_WB_2 (
    .I(DLX_opcode_of_MEM[2]),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_opcode_of_WB[2])
  );
  defparam DLX_opcode_of_WB_3.INIT = 1'b0;
  X_SFF DLX_opcode_of_WB_3 (
    .I(DLX_opcode_of_MEM[3]),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_opcode_of_WB[3])
  );
  defparam DLX_EXinst_reg_out_B_EX_9.INIT = 1'b0;
  X_FF DLX_EXinst_reg_out_B_EX_9 (
    .I(DLX_EXinst__n0007[9]),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_reg_out_B_EX<9>/FFX/RST ),
    .O(DLX_EXinst_reg_out_B_EX[9])
  );
  X_OR2 \DLX_EXinst_reg_out_B_EX<9>/FFX/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_reg_out_B_EX<9>/FFX/RST )
  );
  defparam DLX_EXinst_reg_dst_out_1.INIT = 1'b0;
  X_FF DLX_EXinst_reg_dst_out_1 (
    .I(DLX_EXinst__n0008[1]),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_reg_dst_out<1>/FFX/RST ),
    .O(DLX_EXinst_reg_dst_out[1])
  );
  X_OR2 \DLX_EXinst_reg_dst_out<1>/FFX/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_reg_dst_out<1>/FFX/RST )
  );
  defparam DLX_EXinst_reg_dst_out_3.INIT = 1'b0;
  X_FF DLX_EXinst_reg_dst_out_3 (
    .I(DLX_EXinst__n0008[3]),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_reg_dst_out<3>/FFX/RST ),
    .O(DLX_EXinst_reg_dst_out[3])
  );
  X_OR2 \DLX_EXinst_reg_dst_out<3>/FFX/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_reg_dst_out<3>/FFX/RST )
  );
  defparam DLX_IDinst_IR_function_field_5.INIT = 1'b0;
  X_FF DLX_IDinst_IR_function_field_5 (
    .I(DLX_IDinst__n0114[5]),
    .CE(DLX_IDinst__n0422),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_IR_function_field<5>/FFX/RST ),
    .O(DLX_IDinst_IR_function_field[5])
  );
  X_OR2 \DLX_IDinst_IR_function_field<5>/FFX/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_IR_function_field<5>/FFX/RST )
  );
  defparam DLX_IDinst_reg_out_A_28.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_A_28 (
    .I(N104508),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_A<28>/FFY/RST ),
    .O(DLX_IDinst_reg_out_A[28])
  );
  X_OR2 \DLX_IDinst_reg_out_A<28>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_A<28>/FFY/RST )
  );
  defparam DLX_IDinst_reg_out_A_5.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_A_5 (
    .I(N103012),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_A<5>/FFY/RST ),
    .O(DLX_IDinst_reg_out_A[5])
  );
  X_OR2 \DLX_IDinst_reg_out_A<5>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_A<5>/FFY/RST )
  );
  defparam DLX_opcode_of_WB_4.INIT = 1'b0;
  X_SFF DLX_opcode_of_WB_4 (
    .I(DLX_opcode_of_MEM[4]),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_opcode_of_WB[4])
  );
  defparam DLX_opcode_of_WB_5.INIT = 1'b0;
  X_SFF DLX_opcode_of_WB_5 (
    .I(DLX_opcode_of_MEM[5]),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_opcode_of_WB[5])
  );
  defparam DLX_IDinst_reg_out_A_7.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_A_7 (
    .I(N103080),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_A<7>/FFY/RST ),
    .O(DLX_IDinst_reg_out_A[7])
  );
  X_OR2 \DLX_IDinst_reg_out_A<7>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_A<7>/FFY/RST )
  );
  defparam DLX_IDinst_IR_opcode_field_3.INIT = 1'b0;
  X_FF DLX_IDinst_IR_opcode_field_3 (
    .I(DLX_IDinst__n0113[3]),
    .CE(DLX_IDinst__n0422),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_IR_opcode_field<3>/FFY/RST ),
    .O(DLX_IDinst_IR_opcode_field[3])
  );
  X_OR2 \DLX_IDinst_IR_opcode_field<3>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_IR_opcode_field<3>/FFY/RST )
  );
  defparam DLX_IFinst_PC_2.INIT = 1'b0;
  X_FF DLX_IFinst_PC_2 (
    .I(DLX_IFinst_NPC[2]),
    .CE(DLX_IFinst_PC_N3535),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_PC<3>/FFY/RST ),
    .O(DLX_IFinst_PC[2])
  );
  X_OR2 \DLX_IFinst_PC<3>/FFY/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_PC<3>/FFY/RST )
  );
  defparam DLX_IFinst_PC_1.INIT = 1'b0;
  X_FF DLX_IFinst_PC_1 (
    .I(DLX_IFinst_NPC[1]),
    .CE(DLX_IFinst_PC_N3535),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_PC<1>/FFX/RST ),
    .O(DLX_IFinst_PC[1])
  );
  X_OR2 \DLX_IFinst_PC<1>/FFX/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_PC<1>/FFX/RST )
  );
  defparam DLX_IFinst_PC_4.INIT = 1'b0;
  X_FF DLX_IFinst_PC_4 (
    .I(DLX_IFinst_NPC[4]),
    .CE(DLX_IFinst_PC_N3535),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_PC<5>/FFY/RST ),
    .O(DLX_IFinst_PC[4])
  );
  X_OR2 \DLX_IFinst_PC<5>/FFY/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_PC<5>/FFY/RST )
  );
  defparam DLX_IFinst_PC_3.INIT = 1'b0;
  X_FF DLX_IFinst_PC_3 (
    .I(DLX_IFinst_NPC[3]),
    .CE(DLX_IFinst_PC_N3535),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_PC<3>/FFX/RST ),
    .O(DLX_IFinst_PC[3])
  );
  X_OR2 \DLX_IFinst_PC<3>/FFX/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_PC<3>/FFX/RST )
  );
  defparam DLX_IFinst_PC_6.INIT = 1'b0;
  X_FF DLX_IFinst_PC_6 (
    .I(DLX_IFinst_NPC[6]),
    .CE(DLX_IFinst_PC_N3535),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_PC<7>/FFY/RST ),
    .O(DLX_IFinst_PC[6])
  );
  X_OR2 \DLX_IFinst_PC<7>/FFY/RSTOR  (
    .I0(reset_IBUF_1),
    .I1(GSR),
    .O(\DLX_IFinst_PC<7>/FFY/RST )
  );
  defparam DLX_IFinst_PC_5.INIT = 1'b0;
  X_FF DLX_IFinst_PC_5 (
    .I(DLX_IFinst_NPC[5]),
    .CE(DLX_IFinst_PC_N3535),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_PC<5>/FFX/RST ),
    .O(DLX_IFinst_PC[5])
  );
  X_OR2 \DLX_IFinst_PC<5>/FFX/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_PC<5>/FFX/RST )
  );
  defparam DLX_IFinst_PC_7.INIT = 1'b0;
  X_FF DLX_IFinst_PC_7 (
    .I(DLX_IFinst_NPC[7]),
    .CE(DLX_IFinst_PC_N3535),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_PC<7>/FFX/RST ),
    .O(DLX_IFinst_PC[7])
  );
  X_OR2 \DLX_IFinst_PC<7>/FFX/RSTOR  (
    .I0(reset_IBUF_1),
    .I1(GSR),
    .O(\DLX_IFinst_PC<7>/FFX/RST )
  );
  defparam DLX_IFinst_PC_9.INIT = 1'b0;
  X_FF DLX_IFinst_PC_9 (
    .I(DLX_IFinst_NPC[9]),
    .CE(DLX_IFinst_PC_N3535),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_PC<9>/FFX/RST ),
    .O(DLX_IFinst_PC[9])
  );
  X_OR2 \DLX_IFinst_PC<9>/FFX/RSTOR  (
    .I0(reset_IBUF_1),
    .I1(GSR),
    .O(\DLX_IFinst_PC<9>/FFX/RST )
  );
  defparam DLX_IDinst_Imm_31.INIT = 1'b0;
  X_FF DLX_IDinst_Imm_31 (
    .I(\DLX_IDinst_Imm_31_1/GROM ),
    .CE(DLX_IDinst__n0422),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_Imm_31_1/FFY/RST ),
    .O(\DLX_IDinst_Imm[31] )
  );
  X_OR2 \DLX_IDinst_Imm_31_1/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_Imm_31_1/FFY/RST )
  );
  defparam DLX_IDinst_Imm_31_1_1201.INIT = 1'b0;
  X_FF DLX_IDinst_Imm_31_1_1201 (
    .I(N106726),
    .CE(DLX_IDinst__n0422),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_Imm_31_1/FFX/RST ),
    .O(DLX_IDinst_Imm_31_1)
  );
  X_OR2 \DLX_IDinst_Imm_31_1/FFX/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_Imm_31_1/FFX/RST )
  );
  defparam DLX_IDinst_branch_sig_1202.INIT = 1'b0;
  X_FF DLX_IDinst_branch_sig_1202 (
    .I(\DLX_IDinst_branch_sig/GROM ),
    .CE(DLX_IDinst__n0422),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_branch_sig/FFY/RST ),
    .O(DLX_IDinst_branch_sig)
  );
  X_OR2 \DLX_IDinst_branch_sig/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_branch_sig/FFY/RST )
  );
  defparam DLX_EXinst_ALU_result_24.INIT = 1'b0;
  X_FF DLX_EXinst_ALU_result_24 (
    .I(N112254),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_ALU_result<24>/FFY/RST ),
    .O(DLX_EXinst_ALU_result[24])
  );
  X_OR2 \DLX_EXinst_ALU_result<24>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_ALU_result<24>/FFY/RST )
  );
  defparam vga_top_vga1_helpcounter_1.INIT = 1'b0;
  X_SFF vga_top_vga1_helpcounter_1 (
    .I(vga_top_vga1_helpcounter__n0000[1]),
    .CE(VCC),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(vga_top_vga1__n0052),
    .SRST(reset_IBUF_1),
    .O(vga_top_vga1_helpcounter[1])
  );
  defparam vga_top_vga1_helpcounter_0.INIT = 1'b0;
  X_SFF vga_top_vga1_helpcounter_0 (
    .I(\vga_top_vga1_helpcounter<0>/BXMUXNOT ),
    .CE(VCC),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(vga_top_vga1__n0052),
    .SRST(reset_IBUF_1),
    .O(vga_top_vga1_helpcounter[0])
  );
  defparam DLX_EXinst_ALU_result_21.INIT = 1'b0;
  X_FF DLX_EXinst_ALU_result_21 (
    .I(N114850),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_ALU_result<21>/FFY/RST ),
    .O(DLX_EXinst_ALU_result[21])
  );
  X_OR2 \DLX_EXinst_ALU_result<21>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_ALU_result<21>/FFY/RST )
  );
  defparam DLX_MEMinst_noop_1203.INIT = 1'b1;
  X_FF DLX_MEMinst_noop_1203 (
    .I(DLX_EXinst_noop),
    .CE(VCC),
    .CLK(\DLX_MEMinst_noop/CKMUXNOT ),
    .SET(\DLX_MEMinst_noop/FFY/SET ),
    .RST(GND),
    .O(DLX_MEMinst_noop)
  );
  X_OR2 \DLX_MEMinst_noop/FFY/SETOR  (
    .I0(GSR),
    .I1(reset_IBUF_1),
    .O(\DLX_MEMinst_noop/FFY/SET )
  );
  defparam DLX_IFinst_NPC_13.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_13 (
    .I(\DLX_IFinst_NPC<13>/GROM ),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_NPC<13>/FFY/RST ),
    .O(DLX_IFinst_NPC[13])
  );
  X_OR2 \DLX_IFinst_NPC<13>/FFY/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_NPC<13>/FFY/RST )
  );
  defparam DLX_IFinst_NPC_21.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_21 (
    .I(DLX_IFinst__n0001[21]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_NPC<21>/FFY/RST ),
    .O(DLX_IFinst_NPC[21])
  );
  X_OR2 \DLX_IFinst_NPC<21>/FFY/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_NPC<21>/FFY/RST )
  );
  defparam DLX_IDinst_rt_addr_0.INIT = 1'b0;
  X_FF DLX_IDinst_rt_addr_0 (
    .I(DLX_IDinst__n0106[0]),
    .CE(DLX_IDinst__n0422),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_rt_addr<0>/FFY/RST ),
    .O(DLX_IDinst_rt_addr[0])
  );
  X_OR2 \DLX_IDinst_rt_addr<0>/FFY/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IDinst_rt_addr<0>/FFY/RST )
  );
  defparam DLX_IDinst_IR_opcode_field_4.INIT = 1'b0;
  X_FF DLX_IDinst_IR_opcode_field_4 (
    .I(DLX_IDinst__n0113[4]),
    .CE(DLX_IDinst__n0422),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_IR_opcode_field<4>/FFY/RST ),
    .O(DLX_IDinst_IR_opcode_field[4])
  );
  X_OR2 \DLX_IDinst_IR_opcode_field<4>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_IR_opcode_field<4>/FFY/RST )
  );
  defparam DLX_EXinst_ALU_result_0.INIT = 1'b0;
  X_FF DLX_EXinst_ALU_result_0 (
    .I(\DLX_EXinst_ALU_result<0>/GROM ),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_ALU_result<0>/FFY/RST ),
    .O(DLX_EXinst_ALU_result[0])
  );
  X_OR2 \DLX_EXinst_ALU_result<0>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_ALU_result<0>/FFY/RST )
  );
  defparam DLX_EXinst_ALU_result_1.INIT = 1'b0;
  X_FF DLX_EXinst_ALU_result_1 (
    .I(\DLX_EXinst_ALU_result<1>/GROM ),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_ALU_result<1>/FFY/RST ),
    .O(DLX_EXinst_ALU_result[1])
  );
  X_OR2 \DLX_EXinst_ALU_result<1>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_ALU_result<1>/FFY/RST )
  );
  defparam DLX_EXinst_reg_out_B_EX_15.INIT = 1'b0;
  X_FF DLX_EXinst_reg_out_B_EX_15 (
    .I(DLX_EXinst__n0007[15]),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_reg_out_B_EX<15>/FFY/RST ),
    .O(DLX_EXinst_reg_out_B_EX[15])
  );
  X_OR2 \DLX_EXinst_reg_out_B_EX<15>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_reg_out_B_EX<15>/FFY/RST )
  );
  defparam DLX_IFinst_IR_previous_10.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_10 (
    .I(DLX_IFinst_IR_latched[10]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[10])
  );
  defparam DLX_IFinst_IR_previous_11.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_11 (
    .I(DLX_IFinst_IR_latched[11]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[11])
  );
  defparam DLX_IFinst_IR_previous_12.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_12 (
    .I(DLX_IFinst_IR_latched[12]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[12])
  );
  defparam DLX_IFinst_IR_previous_20.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_20 (
    .I(DLX_IFinst_IR_latched[20]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[20])
  );
  defparam DLX_EXinst_reg_out_B_EX_31.INIT = 1'b0;
  X_FF DLX_EXinst_reg_out_B_EX_31 (
    .I(DLX_EXinst__n0007[31]),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_reg_out_B_EX<31>/FFY/RST ),
    .O(DLX_EXinst_reg_out_B_EX[31])
  );
  X_OR2 \DLX_EXinst_reg_out_B_EX<31>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_reg_out_B_EX<31>/FFY/RST )
  );
  defparam DLX_IFinst_IR_previous_21.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_21 (
    .I(DLX_IFinst_IR_latched[21]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[21])
  );
  defparam DLX_IFinst_IR_previous_13.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_13 (
    .I(DLX_IFinst_IR_latched[13]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[13])
  );
  defparam DLX_IFinst_IR_previous_22.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_22 (
    .I(DLX_IFinst_IR_latched[22]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[22])
  );
  defparam DLX_IFinst_IR_previous_23.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_23 (
    .I(DLX_IFinst_IR_latched[23]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[23])
  );
  defparam DLX_IFinst_IR_previous_15.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_15 (
    .I(DLX_IFinst_IR_latched[15]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[15])
  );
  defparam DLX_IFinst_IR_previous_14.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_14 (
    .I(DLX_IFinst_IR_latched[14]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[14])
  );
  defparam DLX_IFinst_IR_previous_31.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_31 (
    .I(DLX_IFinst_IR_latched[31]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[31])
  );
  defparam DLX_IFinst_IR_previous_30.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_30 (
    .I(DLX_IFinst_IR_latched[30]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[30])
  );
  defparam DLX_IFinst_IR_previous_24.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_24 (
    .I(DLX_IFinst_IR_latched[24]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[24])
  );
  defparam DLX_IFinst_IR_previous_25.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_25 (
    .I(DLX_IFinst_IR_latched[25]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[25])
  );
  defparam DLX_IFinst_IR_previous_17.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_17 (
    .I(DLX_IFinst_IR_latched[17]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[17])
  );
  defparam DLX_IFinst_IR_previous_16.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_16 (
    .I(DLX_IFinst_IR_latched[16]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[16])
  );
  defparam DLX_IFinst_PC_10.INIT = 1'b0;
  X_FF DLX_IFinst_PC_10 (
    .I(DLX_IFinst_NPC[10]),
    .CE(DLX_IFinst_PC_N3535),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_PC<11>/FFY/RST ),
    .O(DLX_IFinst_PC[10])
  );
  X_OR2 \DLX_IFinst_PC<11>/FFY/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_PC<11>/FFY/RST )
  );
  defparam DLX_IDinst_branch_address_0.INIT = 1'b0;
  X_FF DLX_IDinst_branch_address_0 (
    .I(N105098),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_branch_address<0>/FFY/RST ),
    .O(DLX_IDinst_branch_address[0])
  );
  X_OR2 \DLX_IDinst_branch_address<0>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_IDinst_branch_address<0>/FFY/RST )
  );
  defparam DLX_EXinst_ALU_result_17.INIT = 1'b0;
  X_FF DLX_EXinst_ALU_result_17 (
    .I(N123529),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_ALU_result<17>/FFY/RST ),
    .O(DLX_EXinst_ALU_result[17])
  );
  X_OR2 \DLX_EXinst_ALU_result<17>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_ALU_result<17>/FFY/RST )
  );
  defparam DLX_EXinst_ALU_result_25.INIT = 1'b0;
  X_FF DLX_EXinst_ALU_result_25 (
    .I(N118327),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_ALU_result<25>/FFY/RST ),
    .O(DLX_EXinst_ALU_result[25])
  );
  X_OR2 \DLX_EXinst_ALU_result<25>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_ALU_result<25>/FFY/RST )
  );
  defparam DLX_IFinst_PC_11.INIT = 1'b0;
  X_FF DLX_IFinst_PC_11 (
    .I(DLX_IFinst_NPC[11]),
    .CE(DLX_IFinst_PC_N3535),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_PC<11>/FFX/RST ),
    .O(DLX_IFinst_PC[11])
  );
  X_OR2 \DLX_IFinst_PC<11>/FFX/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_PC<11>/FFX/RST )
  );
  defparam DLX_IFinst_IR_previous_18.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_18 (
    .I(DLX_IFinst_IR_latched[18]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[18])
  );
  defparam DLX_IFinst_PC_20.INIT = 1'b0;
  X_FF DLX_IFinst_PC_20 (
    .I(DLX_IFinst_NPC[20]),
    .CE(DLX_IFinst_PC_N3535),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_PC<21>/FFY/RST ),
    .O(DLX_IFinst_PC[20])
  );
  X_OR2 \DLX_IFinst_PC<21>/FFY/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_PC<21>/FFY/RST )
  );
  defparam DLX_IFinst_IR_previous_19.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_19 (
    .I(DLX_IFinst_IR_latched[19]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[19])
  );
  defparam DLX_IFinst_IR_previous_27.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_27 (
    .I(DLX_IFinst_IR_latched[27]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[27])
  );
  defparam DLX_IFinst_IR_previous_26.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_26 (
    .I(DLX_IFinst_IR_latched[26]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[26])
  );
  defparam DLX_IFinst_PC_21.INIT = 1'b0;
  X_FF DLX_IFinst_PC_21 (
    .I(DLX_IFinst_NPC[21]),
    .CE(DLX_IFinst_PC_N3535),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_PC<21>/FFX/RST ),
    .O(DLX_IFinst_PC[21])
  );
  X_OR2 \DLX_IFinst_PC<21>/FFX/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_PC<21>/FFX/RST )
  );
  defparam DLX_IFinst_PC_13.INIT = 1'b0;
  X_FF DLX_IFinst_PC_13 (
    .I(DLX_IFinst_NPC[13]),
    .CE(DLX_IFinst_PC_N3535),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_PC<13>/FFX/RST ),
    .O(DLX_IFinst_PC[13])
  );
  X_OR2 \DLX_IFinst_PC<13>/FFX/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_PC<13>/FFX/RST )
  );
  defparam DLX_IFinst_IR_previous_29.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_29 (
    .I(DLX_IFinst_IR_latched[29]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[29])
  );
  defparam DLX_IFinst_PC_31.INIT = 1'b0;
  X_FF DLX_IFinst_PC_31 (
    .I(DLX_IFinst_NPC[31]),
    .CE(DLX_IFinst_PC_N3535),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_PC<31>/FFX/RST ),
    .O(DLX_IFinst_PC[31])
  );
  X_OR2 \DLX_IFinst_PC<31>/FFX/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_PC<31>/FFX/RST )
  );
  defparam DLX_IFinst_PC_30.INIT = 1'b0;
  X_FF DLX_IFinst_PC_30 (
    .I(DLX_IFinst_NPC[30]),
    .CE(DLX_IFinst_PC_N3535),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_PC<31>/FFY/RST ),
    .O(DLX_IFinst_PC[30])
  );
  X_OR2 \DLX_IFinst_PC<31>/FFY/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_PC<31>/FFY/RST )
  );
  defparam DLX_IFinst_PC_23.INIT = 1'b0;
  X_FF DLX_IFinst_PC_23 (
    .I(DLX_IFinst_NPC[23]),
    .CE(DLX_IFinst_PC_N3535),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_PC<23>/FFX/RST ),
    .O(DLX_IFinst_PC[23])
  );
  X_OR2 \DLX_IFinst_PC<23>/FFX/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_PC<23>/FFX/RST )
  );
  defparam DLX_IFinst_PC_15.INIT = 1'b0;
  X_FF DLX_IFinst_PC_15 (
    .I(DLX_IFinst_NPC[15]),
    .CE(DLX_IFinst_PC_N3535),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_PC<15>/FFX/RST ),
    .O(DLX_IFinst_PC[15])
  );
  X_OR2 \DLX_IFinst_PC<15>/FFX/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_PC<15>/FFX/RST )
  );
  defparam DLX_IFinst_PC_24.INIT = 1'b0;
  X_FF DLX_IFinst_PC_24 (
    .I(DLX_IFinst_NPC[24]),
    .CE(DLX_IFinst_PC_N3535),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_PC<25>/FFY/RST ),
    .O(DLX_IFinst_PC[24])
  );
  X_OR2 \DLX_IFinst_PC<25>/FFY/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_PC<25>/FFY/RST )
  );
  defparam DLX_IFinst_PC_25.INIT = 1'b0;
  X_FF DLX_IFinst_PC_25 (
    .I(DLX_IFinst_NPC[25]),
    .CE(DLX_IFinst_PC_N3535),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_PC<25>/FFX/RST ),
    .O(DLX_IFinst_PC[25])
  );
  X_OR2 \DLX_IFinst_PC<25>/FFX/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_PC<25>/FFX/RST )
  );
  defparam DLX_IDinst_slot_num_FFd2_1204.INIT = 1'b0;
  X_FF DLX_IDinst_slot_num_FFd2_1204 (
    .I(\DLX_IDinst_slot_num_FFd2-In ),
    .CE(DLX_IDinst__n0420),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_slot_num_FFd2/FFY/RST ),
    .O(DLX_IDinst_slot_num_FFd2)
  );
  X_OR2 \DLX_IDinst_slot_num_FFd2/FFY/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IDinst_slot_num_FFd2/FFY/RST )
  );
  defparam DLX_IFinst_PC_17.INIT = 1'b0;
  X_FF DLX_IFinst_PC_17 (
    .I(DLX_IFinst_NPC[17]),
    .CE(DLX_IFinst_PC_N3535),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_PC<17>/FFX/RST ),
    .O(DLX_IFinst_PC[17])
  );
  X_OR2 \DLX_IFinst_PC<17>/FFX/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_PC<17>/FFX/RST )
  );
  defparam DLX_IFinst_PC_26.INIT = 1'b0;
  X_FF DLX_IFinst_PC_26 (
    .I(DLX_IFinst_NPC[26]),
    .CE(DLX_IFinst_PC_N3535),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_PC<27>/FFY/RST ),
    .O(DLX_IFinst_PC[26])
  );
  X_OR2 \DLX_IFinst_PC<27>/FFY/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_PC<27>/FFY/RST )
  );
  defparam DLX_IFinst_PC_27.INIT = 1'b0;
  X_FF DLX_IFinst_PC_27 (
    .I(DLX_IFinst_NPC[27]),
    .CE(DLX_IFinst_PC_N3535),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_PC<27>/FFX/RST ),
    .O(DLX_IFinst_PC[27])
  );
  X_OR2 \DLX_IFinst_PC<27>/FFX/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_PC<27>/FFX/RST )
  );
  defparam DLX_IFinst_PC_19.INIT = 1'b0;
  X_FF DLX_IFinst_PC_19 (
    .I(DLX_IFinst_NPC[19]),
    .CE(DLX_IFinst_PC_N3535),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_PC<19>/FFX/RST ),
    .O(DLX_IFinst_PC[19])
  );
  X_OR2 \DLX_IFinst_PC<19>/FFX/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_PC<19>/FFX/RST )
  );
  defparam DLX_IFinst_PC_28.INIT = 1'b0;
  X_FF DLX_IFinst_PC_28 (
    .I(DLX_IFinst_NPC[28]),
    .CE(DLX_IFinst_PC_N3535),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_PC<29>/FFY/RST ),
    .O(DLX_IFinst_PC[28])
  );
  X_OR2 \DLX_IFinst_PC<29>/FFY/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_PC<29>/FFY/RST )
  );
  defparam DLX_IFinst_PC_29.INIT = 1'b0;
  X_FF DLX_IFinst_PC_29 (
    .I(DLX_IFinst_NPC[29]),
    .CE(DLX_IFinst_PC_N3535),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_PC<29>/FFX/RST ),
    .O(DLX_IFinst_PC[29])
  );
  X_OR2 \DLX_IFinst_PC<29>/FFX/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_PC<29>/FFX/RST )
  );
  defparam DLX_IDinst_branch_address_1.INIT = 1'b0;
  X_FF DLX_IDinst_branch_address_1 (
    .I(N105224),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_branch_address<1>/FFY/RST ),
    .O(DLX_IDinst_branch_address[1])
  );
  X_OR2 \DLX_IDinst_branch_address<1>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_IDinst_branch_address<1>/FFY/RST )
  );
  defparam vga_top_vga1_clockcounter_FFd1_1205.INIT = 1'b0;
  X_SFF vga_top_vga1_clockcounter_FFd1_1205 (
    .I(vga_top_vga1_clockcounter_FFd2),
    .CE(VCC),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(vga_top_vga1_clockcounter_FFd1)
  );
  defparam vga_top_vga1_clockcounter_FFd2_1206.INIT = 1'b1;
  X_SFF vga_top_vga1_clockcounter_FFd2_1206 (
    .I(vga_top_vga1_clockcounter_FFd1),
    .CE(VCC),
    .CLK(clkdiv_vga),
    .SET(GSR),
    .RST(GND),
    .SSET(reset_IBUF_1),
    .SRST(GND),
    .O(vga_top_vga1_clockcounter_FFd2)
  );
  defparam DLX_IDinst_branch_address_2.INIT = 1'b0;
  X_FF DLX_IDinst_branch_address_2 (
    .I(N105161),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_branch_address<2>/FFY/RST ),
    .O(DLX_IDinst_branch_address[2])
  );
  X_OR2 \DLX_IDinst_branch_address<2>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_branch_address<2>/FFY/RST )
  );
  defparam DLX_IDinst_branch_address_3.INIT = 1'b0;
  X_FF DLX_IDinst_branch_address_3 (
    .I(N105287),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_branch_address<3>/FFY/RST ),
    .O(DLX_IDinst_branch_address[3])
  );
  X_OR2 \DLX_IDinst_branch_address<3>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_branch_address<3>/FFY/RST )
  );
  defparam DLX_IDinst_branch_address_4.INIT = 1'b0;
  X_FF DLX_IDinst_branch_address_4 (
    .I(N105350),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_branch_address<4>/FFY/RST ),
    .O(DLX_IDinst_branch_address[4])
  );
  X_OR2 \DLX_IDinst_branch_address<4>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_branch_address<4>/FFY/RST )
  );
  defparam DLX_IDinst_branch_address_5.INIT = 1'b0;
  X_FF DLX_IDinst_branch_address_5 (
    .I(N105413),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_branch_address<5>/FFY/RST ),
    .O(DLX_IDinst_branch_address[5])
  );
  X_OR2 \DLX_IDinst_branch_address<5>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_branch_address<5>/FFY/RST )
  );
  defparam DLX_IDinst_branch_address_6.INIT = 1'b0;
  X_FF DLX_IDinst_branch_address_6 (
    .I(N105535),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_branch_address<6>/FFY/RST ),
    .O(DLX_IDinst_branch_address[6])
  );
  X_OR2 \DLX_IDinst_branch_address<6>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_branch_address<6>/FFY/RST )
  );
  defparam DLX_IDinst_branch_address_7.INIT = 1'b0;
  X_FF DLX_IDinst_branch_address_7 (
    .I(N105474),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_branch_address<7>/FFY/RST ),
    .O(DLX_IDinst_branch_address[7])
  );
  X_OR2 \DLX_IDinst_branch_address<7>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_branch_address<7>/FFY/RST )
  );
  defparam DLX_IDinst_branch_address_8.INIT = 1'b0;
  X_FF DLX_IDinst_branch_address_8 (
    .I(N105598),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_branch_address<8>/FFY/RST ),
    .O(DLX_IDinst_branch_address[8])
  );
  X_OR2 \DLX_IDinst_branch_address<8>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_branch_address<8>/FFY/RST )
  );
  defparam DLX_IDinst_rd_addr_0.INIT = 1'b0;
  X_FF DLX_IDinst_rd_addr_0 (
    .I(DLX_IDinst__n0107[0]),
    .CE(DLX_IDinst__n0422),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_rd_addr<0>/FFY/RST ),
    .O(DLX_IDinst_rd_addr[0])
  );
  X_OR2 \DLX_IDinst_rd_addr<0>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_rd_addr<0>/FFY/RST )
  );
  defparam DLX_IDinst_branch_address_9.INIT = 1'b0;
  X_FF DLX_IDinst_branch_address_9 (
    .I(N105661),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_branch_address<9>/FFY/RST ),
    .O(DLX_IDinst_branch_address[9])
  );
  X_OR2 \DLX_IDinst_branch_address<9>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_branch_address<9>/FFY/RST )
  );
  defparam DLX_IDinst_Imm_12.INIT = 1'b0;
  X_FF DLX_IDinst_Imm_12 (
    .I(DLX_IDinst__n0093),
    .CE(DLX_IDinst__n0422),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_Imm<12>/FFY/RST ),
    .O(\DLX_IDinst_Imm[12] )
  );
  X_OR2 \DLX_IDinst_Imm<12>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_Imm<12>/FFY/RST )
  );
  defparam DLX_IDinst_Imm_5.INIT = 1'b0;
  X_FF DLX_IDinst_Imm_5 (
    .I(DLX_IDinst__n0100),
    .CE(DLX_IDinst__n0422),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_Imm<5>/FFY/RST ),
    .O(\DLX_IDinst_Imm[5] )
  );
  X_OR2 \DLX_IDinst_Imm<5>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_Imm<5>/FFY/RST )
  );
  defparam DLX_IDinst_Imm_13.INIT = 1'b0;
  X_FF DLX_IDinst_Imm_13 (
    .I(DLX_IDinst__n0092),
    .CE(DLX_IDinst__n0422),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_Imm<13>/FFY/RST ),
    .O(\DLX_IDinst_Imm[13] )
  );
  X_OR2 \DLX_IDinst_Imm<13>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_Imm<13>/FFY/RST )
  );
  defparam DLX_IDinst_Imm_14.INIT = 1'b0;
  X_FF DLX_IDinst_Imm_14 (
    .I(DLX_IDinst__n0091),
    .CE(DLX_IDinst__n0422),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_Imm<14>/FFY/RST ),
    .O(\DLX_IDinst_Imm[14] )
  );
  X_OR2 \DLX_IDinst_Imm<14>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_Imm<14>/FFY/RST )
  );
  defparam DLX_IDinst_Imm_15.INIT = 1'b0;
  X_FF DLX_IDinst_Imm_15 (
    .I(DLX_IDinst__n0090),
    .CE(DLX_IDinst__n0422),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_Imm<15>/FFY/RST ),
    .O(\DLX_IDinst_Imm[15] )
  );
  X_OR2 \DLX_IDinst_Imm<15>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_Imm<15>/FFY/RST )
  );
  defparam vga_top_vga1_videoon_1207.INIT = 1'b0;
  X_SFF vga_top_vga1_videoon_1207 (
    .I(\vga_top_vga1_videoon/LOGIC_ONE ),
    .CE(VCC),
    .CLK(clkdiv_vga),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(N110183),
    .O(vga_top_vga1_videoon)
  );
  defparam DLX_EXinst_ALU_result_3.INIT = 1'b0;
  X_FF DLX_EXinst_ALU_result_3 (
    .I(\DLX_EXinst_ALU_result<3>/GROM ),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_ALU_result<3>/FFY/RST ),
    .O(DLX_EXinst_ALU_result[3])
  );
  X_OR2 \DLX_EXinst_ALU_result<3>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_ALU_result<3>/FFY/RST )
  );
  defparam DLX_IDinst_reg_out_B_0.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_B_0 (
    .I(DLX_IDinst__n0118[0]),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_B<0>/FFY/RST ),
    .O(DLX_IDinst_reg_out_B[0])
  );
  X_OR2 \DLX_IDinst_reg_out_B<0>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_B<0>/FFY/RST )
  );
  defparam DLX_EXinst_ALU_result_4.INIT = 1'b0;
  X_FF DLX_EXinst_ALU_result_4 (
    .I(\DLX_EXinst_ALU_result<4>/GROM ),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_ALU_result<4>/FFY/RST ),
    .O(DLX_EXinst_ALU_result[4])
  );
  X_OR2 \DLX_EXinst_ALU_result<4>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_ALU_result<4>/FFY/RST )
  );
  defparam DLX_EXinst_ALU_result_5.INIT = 1'b0;
  X_FF DLX_EXinst_ALU_result_5 (
    .I(\DLX_EXinst_ALU_result<5>/GROM ),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_ALU_result<5>/FFY/RST ),
    .O(DLX_EXinst_ALU_result[5])
  );
  X_OR2 \DLX_EXinst_ALU_result<5>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_ALU_result<5>/FFY/RST )
  );
  defparam DLX_EXinst_ALU_result_22.INIT = 1'b0;
  X_FF DLX_EXinst_ALU_result_22 (
    .I(N114452),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_ALU_result<22>/FFY/RST ),
    .O(DLX_EXinst_ALU_result[22])
  );
  X_OR2 \DLX_EXinst_ALU_result<22>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_ALU_result<22>/FFY/RST )
  );
  defparam DLX_EXinst_ALU_result_6.INIT = 1'b0;
  X_FF DLX_EXinst_ALU_result_6 (
    .I(\DLX_EXinst_ALU_result<6>/GROM ),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_ALU_result<6>/FFY/RST ),
    .O(DLX_EXinst_ALU_result[6])
  );
  X_OR2 \DLX_EXinst_ALU_result<6>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_ALU_result<6>/FFY/RST )
  );
  defparam DLX_EXinst_ALU_result_7.INIT = 1'b0;
  X_FF DLX_EXinst_ALU_result_7 (
    .I(\DLX_EXinst_ALU_result<7>/GROM ),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_ALU_result<7>/FFY/RST ),
    .O(DLX_EXinst_ALU_result[7])
  );
  X_OR2 \DLX_EXinst_ALU_result<7>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_ALU_result<7>/FFY/RST )
  );
  defparam DLX_IDinst_branch_address_11.INIT = 1'b0;
  X_FF DLX_IDinst_branch_address_11 (
    .I(N105787),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_branch_address<11>/FFY/RST ),
    .O(DLX_IDinst_branch_address[11])
  );
  X_OR2 \DLX_IDinst_branch_address<11>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_IDinst_branch_address<11>/FFY/RST )
  );
  defparam DLX_IDinst_mem_to_reg_1208.INIT = 1'b0;
  X_FF DLX_IDinst_mem_to_reg_1208 (
    .I(DLX_IDinst__n0110),
    .CE(DLX_IDinst__n0422),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_mem_to_reg/FFY/RST ),
    .O(DLX_IDinst_mem_to_reg)
  );
  X_OR2 \DLX_IDinst_mem_to_reg/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_mem_to_reg/FFY/RST )
  );
  defparam DLX_IDinst_branch_address_10.INIT = 1'b0;
  X_FF DLX_IDinst_branch_address_10 (
    .I(N105724),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_branch_address<10>/FFY/RST ),
    .O(DLX_IDinst_branch_address[10])
  );
  X_OR2 \DLX_IDinst_branch_address<10>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_IDinst_branch_address<10>/FFY/RST )
  );
  defparam DLX_EXinst_ALU_result_8.INIT = 1'b0;
  X_FF DLX_EXinst_ALU_result_8 (
    .I(\DLX_EXinst_ALU_result<8>/GROM ),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_ALU_result<8>/FFY/RST ),
    .O(DLX_EXinst_ALU_result[8])
  );
  X_OR2 \DLX_EXinst_ALU_result<8>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_ALU_result<8>/FFY/RST )
  );
  defparam DLX_IDinst_branch_address_12.INIT = 1'b0;
  X_FF DLX_IDinst_branch_address_12 (
    .I(N105850),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_branch_address<12>/FFY/RST ),
    .O(DLX_IDinst_branch_address[12])
  );
  X_OR2 \DLX_IDinst_branch_address<12>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_IDinst_branch_address<12>/FFY/RST )
  );
  defparam DLX_IDinst_branch_address_20.INIT = 1'b0;
  X_FF DLX_IDinst_branch_address_20 (
    .I(N106354),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_branch_address<20>/FFY/RST ),
    .O(DLX_IDinst_branch_address[20])
  );
  X_OR2 \DLX_IDinst_branch_address<20>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_branch_address<20>/FFY/RST )
  );
  defparam DLX_EXinst_ALU_result_9.INIT = 1'b0;
  X_FF DLX_EXinst_ALU_result_9 (
    .I(\DLX_EXinst_ALU_result<9>/GROM ),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_ALU_result<9>/FFY/RST ),
    .O(DLX_EXinst_ALU_result[9])
  );
  X_OR2 \DLX_EXinst_ALU_result<9>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_ALU_result<9>/FFY/RST )
  );
  defparam DLX_EXinst_ALU_result_18.INIT = 1'b0;
  X_FF DLX_EXinst_ALU_result_18 (
    .I(N122511),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_ALU_result<18>/FFY/RST ),
    .O(DLX_EXinst_ALU_result[18])
  );
  X_OR2 \DLX_EXinst_ALU_result<18>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_ALU_result<18>/FFY/RST )
  );
  defparam DLX_EXinst_ALU_result_26.INIT = 1'b0;
  X_FF DLX_EXinst_ALU_result_26 (
    .I(N117936),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_ALU_result<26>/FFY/RST ),
    .O(DLX_EXinst_ALU_result[26])
  );
  X_OR2 \DLX_EXinst_ALU_result<26>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_ALU_result<26>/FFY/RST )
  );
  defparam DLX_IDinst_CLI_1209.INIT = 1'b0;
  X_FF DLX_IDinst_CLI_1209 (
    .I(\DLX_IDinst_CLI/GROM ),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_CLI/FFY/RST ),
    .O(DLX_IDinst_CLI)
  );
  X_OR2 \DLX_IDinst_CLI/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_CLI/FFY/RST )
  );
  defparam DLX_EXinst_noop_1210.INIT = 1'b1;
  X_FF DLX_EXinst_noop_1210 (
    .I(N101911),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(\DLX_EXinst_noop/FFY/SET ),
    .RST(GND),
    .O(DLX_EXinst_noop)
  );
  X_OR2 \DLX_EXinst_noop/FFY/SETOR  (
    .I0(GSR),
    .I1(reset_IBUF),
    .O(\DLX_EXinst_noop/FFY/SET )
  );
  defparam DLX_IDinst_branch_address_14.INIT = 1'b0;
  X_FF DLX_IDinst_branch_address_14 (
    .I(N105976),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_branch_address<14>/FFY/RST ),
    .O(DLX_IDinst_branch_address[14])
  );
  X_OR2 \DLX_IDinst_branch_address<14>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_IDinst_branch_address<14>/FFY/RST )
  );
  defparam DLX_IDinst_branch_address_30.INIT = 1'b0;
  X_FF DLX_IDinst_branch_address_30 (
    .I(N106417),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_branch_address<30>/FFY/RST ),
    .O(DLX_IDinst_branch_address[30])
  );
  X_OR2 \DLX_IDinst_branch_address<30>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_branch_address<30>/FFY/RST )
  );
  defparam DLX_IDinst_branch_address_22.INIT = 1'b0;
  X_FF DLX_IDinst_branch_address_22 (
    .I(N106606),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_branch_address<22>/FFY/RST ),
    .O(DLX_IDinst_branch_address[22])
  );
  X_OR2 \DLX_IDinst_branch_address<22>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_branch_address<22>/FFY/RST )
  );
  defparam DLX_IDinst_branch_address_21.INIT = 1'b0;
  X_FF DLX_IDinst_branch_address_21 (
    .I(N106480),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_branch_address<21>/FFY/RST ),
    .O(DLX_IDinst_branch_address[21])
  );
  X_OR2 \DLX_IDinst_branch_address<21>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_branch_address<21>/FFY/RST )
  );
  defparam DLX_IDinst_branch_address_13.INIT = 1'b0;
  X_FF DLX_IDinst_branch_address_13 (
    .I(N105913),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_branch_address<13>/FFY/RST ),
    .O(DLX_IDinst_branch_address[13])
  );
  X_OR2 \DLX_IDinst_branch_address<13>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_IDinst_branch_address<13>/FFY/RST )
  );
  defparam DLX_IDinst_stall_1211.INIT = 1'b0;
  X_FF DLX_IDinst_stall_1211 (
    .I(\DLX_IDinst_stall/GROM ),
    .CE(DLX_IDinst__n0441),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_stall/FFY/RST ),
    .O(DLX_IDinst_stall)
  );
  X_OR2 \DLX_IDinst_stall/FFY/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IDinst_stall/FFY/RST )
  );
  defparam DLX_IDinst_branch_address_17.INIT = 1'b0;
  X_FF DLX_IDinst_branch_address_17 (
    .I(N106165),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_branch_address<17>/FFY/RST ),
    .O(DLX_IDinst_branch_address[17])
  );
  X_OR2 \DLX_IDinst_branch_address<17>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_branch_address<17>/FFY/RST )
  );
  defparam DLX_IDinst_branch_address_25.INIT = 1'b0;
  X_FF DLX_IDinst_branch_address_25 (
    .I(N106789),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_branch_address<25>/FFY/RST ),
    .O(DLX_IDinst_branch_address[25])
  );
  X_OR2 \DLX_IDinst_branch_address<25>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_branch_address<25>/FFY/RST )
  );
  defparam DLX_IFinst_NPC_10.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_10 (
    .I(\DLX_IFinst_NPC<10>/GROM ),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_NPC<10>/FFY/RST ),
    .O(DLX_IFinst_NPC[10])
  );
  X_OR2 \DLX_IFinst_NPC<10>/FFY/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_NPC<10>/FFY/RST )
  );
  defparam DLX_IDinst_branch_address_31.INIT = 1'b0;
  X_FF DLX_IDinst_branch_address_31 (
    .I(N107102),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_branch_address<31>/FFY/RST ),
    .O(DLX_IDinst_branch_address[31])
  );
  X_OR2 \DLX_IDinst_branch_address<31>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_branch_address<31>/FFY/RST )
  );
  defparam DLX_IFinst_NPC_20.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_20 (
    .I(DLX_IFinst__n0001[20]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_NPC<20>/FFY/RST ),
    .O(DLX_IFinst_NPC[20])
  );
  X_OR2 \DLX_IFinst_NPC<20>/FFY/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_NPC<20>/FFY/RST )
  );
  defparam DLX_IFinst_NPC_12.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_12 (
    .I(\DLX_IFinst_NPC<12>/GROM ),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_NPC<12>/FFY/RST ),
    .O(DLX_IFinst_NPC[12])
  );
  X_OR2 \DLX_IFinst_NPC<12>/FFY/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_NPC<12>/FFY/RST )
  );
  defparam DLX_IFinst_NPC_0.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_0 (
    .I(\DLX_IFinst_NPC<0>/GROM ),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_NPC<0>/FFY/RST ),
    .O(DLX_IFinst_NPC[0])
  );
  X_OR2 \DLX_IFinst_NPC<0>/FFY/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_NPC<0>/FFY/RST )
  );
  defparam DLX_IDinst_branch_address_23.INIT = 1'b0;
  X_FF DLX_IDinst_branch_address_23 (
    .I(N106543),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_branch_address<23>/FFY/RST ),
    .O(DLX_IDinst_branch_address[23])
  );
  X_OR2 \DLX_IDinst_branch_address<23>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_branch_address<23>/FFY/RST )
  );
  defparam DLX_IDinst_branch_address_15.INIT = 1'b0;
  X_FF DLX_IDinst_branch_address_15 (
    .I(N106039),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_branch_address<15>/FFY/RST ),
    .O(DLX_IDinst_branch_address[15])
  );
  X_OR2 \DLX_IDinst_branch_address<15>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_branch_address<15>/FFY/RST )
  );
  defparam DLX_IDinst_branch_address_16.INIT = 1'b0;
  X_FF DLX_IDinst_branch_address_16 (
    .I(N106102),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_branch_address<16>/FFY/RST ),
    .O(DLX_IDinst_branch_address[16])
  );
  X_OR2 \DLX_IDinst_branch_address<16>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_branch_address<16>/FFY/RST )
  );
  defparam DLX_IDinst_branch_address_24.INIT = 1'b0;
  X_FF DLX_IDinst_branch_address_24 (
    .I(N106669),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_branch_address<24>/FFY/RST ),
    .O(DLX_IDinst_branch_address[24])
  );
  X_OR2 \DLX_IDinst_branch_address<24>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_branch_address<24>/FFY/RST )
  );
  defparam DLX_IDinst_branch_address_26.INIT = 1'b0;
  X_FF DLX_IDinst_branch_address_26 (
    .I(N106852),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_branch_address<26>/FFY/RST ),
    .O(DLX_IDinst_branch_address[26])
  );
  X_OR2 \DLX_IDinst_branch_address<26>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_branch_address<26>/FFY/RST )
  );
  defparam DLX_IDinst_branch_address_18.INIT = 1'b0;
  X_FF DLX_IDinst_branch_address_18 (
    .I(N106291),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_branch_address<18>/FFY/RST ),
    .O(DLX_IDinst_branch_address[18])
  );
  X_OR2 \DLX_IDinst_branch_address<18>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_branch_address<18>/FFY/RST )
  );
  defparam DLX_IDinst_branch_address_27.INIT = 1'b0;
  X_FF DLX_IDinst_branch_address_27 (
    .I(N106915),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_branch_address<27>/FFY/RST ),
    .O(DLX_IDinst_branch_address[27])
  );
  X_OR2 \DLX_IDinst_branch_address<27>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_branch_address<27>/FFY/RST )
  );
  defparam DLX_IDinst_branch_address_19.INIT = 1'b0;
  X_FF DLX_IDinst_branch_address_19 (
    .I(N106228),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_branch_address<19>/FFY/RST ),
    .O(DLX_IDinst_branch_address[19])
  );
  X_OR2 \DLX_IDinst_branch_address<19>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_branch_address<19>/FFY/RST )
  );
  defparam DLX_IDinst_branch_address_28.INIT = 1'b0;
  X_FF DLX_IDinst_branch_address_28 (
    .I(N106978),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_branch_address<28>/FFY/RST ),
    .O(DLX_IDinst_branch_address[28])
  );
  X_OR2 \DLX_IDinst_branch_address<28>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_branch_address<28>/FFY/RST )
  );
  defparam DLX_EXinst_ALU_result_14.INIT = 1'b0;
  X_FF DLX_EXinst_ALU_result_14 (
    .I(\DLX_EXinst_ALU_result<14>/GROM ),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_ALU_result<14>/FFY/RST ),
    .O(DLX_EXinst_ALU_result[14])
  );
  X_OR2 \DLX_EXinst_ALU_result<14>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_ALU_result<14>/FFY/RST )
  );
  defparam DLX_IDinst_branch_address_29.INIT = 1'b0;
  X_FF DLX_IDinst_branch_address_29 (
    .I(N107041),
    .CE(DLX_IDinst__n0421),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_branch_address<29>/FFY/RST ),
    .O(DLX_IDinst_branch_address[29])
  );
  X_OR2 \DLX_IDinst_branch_address<29>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_branch_address<29>/FFY/RST )
  );
  defparam DLX_IFinst_IR_previous_0.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_0 (
    .I(DLX_IFinst_IR_latched[0]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[0])
  );
  defparam DLX_IFinst_IR_previous_1.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_1 (
    .I(DLX_IFinst_IR_latched[1]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[1])
  );
  defparam DLX_IFinst_NPC_11.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_11 (
    .I(\DLX_IFinst_NPC<11>/GROM ),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_NPC<11>/FFY/RST ),
    .O(DLX_IFinst_NPC[11])
  );
  X_OR2 \DLX_IFinst_NPC<11>/FFY/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_NPC<11>/FFY/RST )
  );
  defparam DLX_IFinst_IR_previous_2.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_2 (
    .I(DLX_IFinst_IR_latched[2]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[2])
  );
  defparam DLX_IFinst_IR_previous_4.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_4 (
    .I(DLX_IFinst_IR_latched[4]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[4])
  );
  defparam DLX_IFinst_IR_previous_3.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_3 (
    .I(DLX_IFinst_IR_latched[3]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[3])
  );
  defparam DLX_IFinst_IR_previous_5.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_5 (
    .I(DLX_IFinst_IR_latched[5]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[5])
  );
  defparam DLX_IFinst_IR_previous_7.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_7 (
    .I(DLX_IFinst_IR_latched[7]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[7])
  );
  defparam DLX_IFinst_IR_previous_6.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_6 (
    .I(DLX_IFinst_IR_latched[6]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[6])
  );
  defparam DLX_IFinst_IR_previous_9.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_9 (
    .I(DLX_IFinst_IR_latched[9]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[9])
  );
  defparam DLX_IFinst_IR_previous_8.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_8 (
    .I(DLX_IFinst_IR_latched[8]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[8])
  );
  defparam DLX_IFinst_NPC_1.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_1 (
    .I(\DLX_IFinst_NPC<1>/GROM ),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_NPC<1>/FFY/RST ),
    .O(DLX_IFinst_NPC[1])
  );
  X_OR2 \DLX_IFinst_NPC<1>/FFY/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_NPC<1>/FFY/RST )
  );
  defparam DLX_IFinst_NPC_4.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_4 (
    .I(\DLX_IFinst_NPC<4>/GROM ),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_NPC<4>/FFY/RST ),
    .O(DLX_IFinst_NPC[4])
  );
  X_OR2 \DLX_IFinst_NPC<4>/FFY/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_NPC<4>/FFY/RST )
  );
  defparam DLX_EXinst_ALU_result_27.INIT = 1'b0;
  X_FF DLX_EXinst_ALU_result_27 (
    .I(N117545),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_ALU_result<27>/FFY/RST ),
    .O(DLX_EXinst_ALU_result[27])
  );
  X_OR2 \DLX_EXinst_ALU_result<27>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_ALU_result<27>/FFY/RST )
  );
  defparam DLX_EXinst_ALU_result_15.INIT = 1'b0;
  X_FF DLX_EXinst_ALU_result_15 (
    .I(N118737),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_ALU_result<15>/FFY/RST ),
    .O(DLX_EXinst_ALU_result[15])
  );
  X_OR2 \DLX_EXinst_ALU_result<15>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_ALU_result<15>/FFY/RST )
  );
  defparam DLX_MEMinst_reg_dst_out_0.INIT = 1'b0;
  X_FF DLX_MEMinst_reg_dst_out_0 (
    .I(DLX_EXinst_reg_dst_out[0]),
    .CE(VCC),
    .CLK(\DLX_MEMinst_reg_dst_out<1>/CKMUXNOT ),
    .SET(GND),
    .RST(\DLX_MEMinst_reg_dst_out<1>/FFY/RST ),
    .O(DLX_MEMinst_reg_dst_out[0])
  );
  X_OR2 \DLX_MEMinst_reg_dst_out<1>/FFY/RSTOR  (
    .I0(reset_IBUF_1),
    .I1(GSR),
    .O(\DLX_MEMinst_reg_dst_out<1>/FFY/RST )
  );
  defparam DLX_MEMinst_reg_dst_out_1.INIT = 1'b0;
  X_FF DLX_MEMinst_reg_dst_out_1 (
    .I(DLX_EXinst_reg_dst_out[1]),
    .CE(VCC),
    .CLK(\DLX_MEMinst_reg_dst_out<1>/CKMUXNOT ),
    .SET(GND),
    .RST(\DLX_MEMinst_reg_dst_out<1>/FFX/RST ),
    .O(DLX_MEMinst_reg_dst_out[1])
  );
  X_OR2 \DLX_MEMinst_reg_dst_out<1>/FFX/RSTOR  (
    .I0(reset_IBUF_1),
    .I1(GSR),
    .O(\DLX_MEMinst_reg_dst_out<1>/FFX/RST )
  );
  defparam DLX_EXinst_ALU_result_31.INIT = 1'b0;
  X_FF DLX_EXinst_ALU_result_31 (
    .I(N124731),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_ALU_result<31>/FFY/RST ),
    .O(DLX_EXinst_ALU_result[31])
  );
  X_OR2 \DLX_EXinst_ALU_result<31>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_ALU_result<31>/FFY/RST )
  );
  defparam DLX_EXinst_ALU_result_10.INIT = 1'b0;
  X_FF DLX_EXinst_ALU_result_10 (
    .I(\DLX_EXinst_ALU_result<10>/GROM ),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_ALU_result<10>/FFY/RST ),
    .O(DLX_EXinst_ALU_result[10])
  );
  X_OR2 \DLX_EXinst_ALU_result<10>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_ALU_result<10>/FFY/RST )
  );
  defparam DLX_IFinst_NPC_30.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_30 (
    .I(DLX_IFinst__n0001[30]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_NPC<30>/FFY/RST ),
    .O(DLX_IFinst_NPC[30])
  );
  X_OR2 \DLX_IFinst_NPC<30>/FFY/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_NPC<30>/FFY/RST )
  );
  defparam DLX_IFinst_NPC_14.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_14 (
    .I(\DLX_IFinst_NPC<14>/GROM ),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_NPC<14>/FFY/RST ),
    .O(DLX_IFinst_NPC[14])
  );
  X_OR2 \DLX_IFinst_NPC<14>/FFY/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_NPC<14>/FFY/RST )
  );
  defparam DLX_IFinst_NPC_22.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_22 (
    .I(DLX_IFinst__n0001[22]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_NPC<22>/FFY/RST ),
    .O(DLX_IFinst_NPC[22])
  );
  X_OR2 \DLX_IFinst_NPC<22>/FFY/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_NPC<22>/FFY/RST )
  );
  defparam DLX_IDinst_reg_dst_1212.INIT = 1'b0;
  X_FF DLX_IDinst_reg_dst_1212 (
    .I(N110380),
    .CE(DLX_IDinst__n0422),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_dst/FFY/RST ),
    .O(DLX_IDinst_reg_dst)
  );
  X_OR2 \DLX_IDinst_reg_dst/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_dst/FFY/RST )
  );
  defparam DLX_EXinst_ALU_result_11.INIT = 1'b0;
  X_FF DLX_EXinst_ALU_result_11 (
    .I(\DLX_EXinst_ALU_result<11>/GROM ),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_ALU_result<11>/FFY/RST ),
    .O(DLX_EXinst_ALU_result[11])
  );
  X_OR2 \DLX_EXinst_ALU_result<11>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_ALU_result<11>/FFY/RST )
  );
  defparam DLX_IFinst_NPC_2.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_2 (
    .I(\DLX_IFinst_NPC<2>/GROM ),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_NPC<2>/FFY/RST ),
    .O(DLX_IFinst_NPC[2])
  );
  X_OR2 \DLX_IFinst_NPC<2>/FFY/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_NPC<2>/FFY/RST )
  );
  defparam DLX_EXinst_ALU_result_20.INIT = 1'b0;
  X_FF DLX_EXinst_ALU_result_20 (
    .I(N119151),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_ALU_result<20>/FFY/RST ),
    .O(DLX_EXinst_ALU_result[20])
  );
  X_OR2 \DLX_EXinst_ALU_result<20>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_ALU_result<20>/FFY/RST )
  );
  defparam DLX_EXinst_ALU_result_23.INIT = 1'b0;
  X_FF DLX_EXinst_ALU_result_23 (
    .I(N114054),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_ALU_result<23>/FFY/RST ),
    .O(DLX_EXinst_ALU_result[23])
  );
  X_OR2 \DLX_EXinst_ALU_result<23>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_ALU_result<23>/FFY/RST )
  );
  defparam DLX_IFinst_NPC_15.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_15 (
    .I(\DLX_IFinst_NPC<15>/GROM ),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_NPC<15>/FFY/RST ),
    .O(DLX_IFinst_NPC[15])
  );
  X_OR2 \DLX_IFinst_NPC<15>/FFY/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_NPC<15>/FFY/RST )
  );
  defparam DLX_IFinst_NPC_31.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_31 (
    .I(DLX_IFinst__n0001[31]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_NPC<31>/FFY/RST ),
    .O(DLX_IFinst_NPC[31])
  );
  X_OR2 \DLX_IFinst_NPC<31>/FFY/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_NPC<31>/FFY/RST )
  );
  defparam DLX_IFinst_NPC_23.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_23 (
    .I(DLX_IFinst__n0001[23]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_NPC<23>/FFY/RST ),
    .O(DLX_IFinst_NPC[23])
  );
  X_OR2 \DLX_IFinst_NPC<23>/FFY/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_NPC<23>/FFY/RST )
  );
  defparam DLX_IFinst_NPC_3.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_3 (
    .I(\DLX_IFinst_NPC<3>/GROM ),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_NPC<3>/FFY/RST ),
    .O(DLX_IFinst_NPC[3])
  );
  X_OR2 \DLX_IFinst_NPC<3>/FFY/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_NPC<3>/FFY/RST )
  );
  defparam DLX_MEMinst_reg_dst_out_2.INIT = 1'b0;
  X_FF DLX_MEMinst_reg_dst_out_2 (
    .I(DLX_EXinst_reg_dst_out[2]),
    .CE(VCC),
    .CLK(\DLX_MEMinst_reg_dst_out<3>/CKMUXNOT ),
    .SET(GND),
    .RST(\DLX_MEMinst_reg_dst_out<3>/FFY/RST ),
    .O(DLX_MEMinst_reg_dst_out[2])
  );
  X_OR2 \DLX_MEMinst_reg_dst_out<3>/FFY/RSTOR  (
    .I0(reset_IBUF_1),
    .I1(GSR),
    .O(\DLX_MEMinst_reg_dst_out<3>/FFY/RST )
  );
  defparam DLX_MEMinst_reg_dst_out_3.INIT = 1'b0;
  X_FF DLX_MEMinst_reg_dst_out_3 (
    .I(DLX_EXinst_reg_dst_out[3]),
    .CE(VCC),
    .CLK(\DLX_MEMinst_reg_dst_out<3>/CKMUXNOT ),
    .SET(GND),
    .RST(\DLX_MEMinst_reg_dst_out<3>/FFX/RST ),
    .O(DLX_MEMinst_reg_dst_out[3])
  );
  X_OR2 \DLX_MEMinst_reg_dst_out<3>/FFX/RSTOR  (
    .I0(reset_IBUF_1),
    .I1(GSR),
    .O(\DLX_MEMinst_reg_dst_out<3>/FFX/RST )
  );
  defparam DLX_MEMinst_reg_dst_out_4.INIT = 1'b0;
  X_FF DLX_MEMinst_reg_dst_out_4 (
    .I(DLX_EXinst_reg_dst_out[4]),
    .CE(VCC),
    .CLK(\DLX_MEMinst_reg_dst_out<4>/CKMUXNOT ),
    .SET(GND),
    .RST(\DLX_MEMinst_reg_dst_out<4>/FFY/RST ),
    .O(DLX_MEMinst_reg_dst_out[4])
  );
  X_OR2 \DLX_MEMinst_reg_dst_out<4>/FFY/RSTOR  (
    .I0(reset_IBUF_1),
    .I1(GSR),
    .O(\DLX_MEMinst_reg_dst_out<4>/FFY/RST )
  );
  defparam DLX_IDinst_slot_num_FFd3_1213.INIT = 1'b1;
  X_FF DLX_IDinst_slot_num_FFd3_1213 (
    .I(\DLX_IDinst_slot_num_FFd3-In ),
    .CE(DLX_IDinst__n0420),
    .CLK(DLX_clk_ID),
    .SET(\DLX_IDinst_slot_num_FFd3/FFY/SET ),
    .RST(GND),
    .O(DLX_IDinst_slot_num_FFd3)
  );
  X_OR2 \DLX_IDinst_slot_num_FFd3/FFY/SETOR  (
    .I0(GSR),
    .I1(reset_IBUF_3),
    .O(\DLX_IDinst_slot_num_FFd3/FFY/SET )
  );
  defparam DLX_IDinst_reg_out_B_2.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_B_2 (
    .I(DLX_IDinst__n0118[2]),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_B<2>/FFY/RST ),
    .O(DLX_IDinst_reg_out_B[2])
  );
  X_OR2 \DLX_IDinst_reg_out_B<2>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_B<2>/FFY/RST )
  );
  defparam DLX_IFinst_NPC_24.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_24 (
    .I(DLX_IFinst__n0001[24]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_NPC<24>/FFY/RST ),
    .O(DLX_IFinst_NPC[24])
  );
  X_OR2 \DLX_IFinst_NPC<24>/FFY/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_NPC<24>/FFY/RST )
  );
  defparam DLX_IFinst_NPC_16.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_16 (
    .I(DLX_IFinst__n0001[16]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_NPC<16>/FFY/RST ),
    .O(DLX_IFinst_NPC[16])
  );
  X_OR2 \DLX_IFinst_NPC<16>/FFY/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_NPC<16>/FFY/RST )
  );
  defparam DLX_EXinst_ALU_result_30.INIT = 1'b0;
  X_FF DLX_EXinst_ALU_result_30 (
    .I(N121549),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_ALU_result<30>/FFY/RST ),
    .O(DLX_EXinst_ALU_result[30])
  );
  X_OR2 \DLX_EXinst_ALU_result<30>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_ALU_result<30>/FFY/RST )
  );
  defparam DLX_IFinst_NPC_26.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_26 (
    .I(DLX_IFinst__n0001[26]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_NPC<26>/FFY/RST ),
    .O(DLX_IFinst_NPC[26])
  );
  X_OR2 \DLX_IFinst_NPC<26>/FFY/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_NPC<26>/FFY/RST )
  );
  defparam DLX_IFinst_NPC_18.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_18 (
    .I(DLX_IFinst__n0001[18]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_NPC<18>/FFY/RST ),
    .O(DLX_IFinst_NPC[18])
  );
  X_OR2 \DLX_IFinst_NPC<18>/FFY/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_NPC<18>/FFY/RST )
  );
  defparam DLX_IFinst_NPC_17.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_17 (
    .I(DLX_IFinst__n0001[17]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_NPC<17>/FFY/RST ),
    .O(DLX_IFinst_NPC[17])
  );
  X_OR2 \DLX_IFinst_NPC<17>/FFY/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_NPC<17>/FFY/RST )
  );
  defparam DLX_IFinst_NPC_25.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_25 (
    .I(DLX_IFinst__n0001[25]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_NPC<25>/FFY/RST ),
    .O(DLX_IFinst_NPC[25])
  );
  X_OR2 \DLX_IFinst_NPC<25>/FFY/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_NPC<25>/FFY/RST )
  );
  defparam DLX_EXinst_ALU_result_16.INIT = 1'b0;
  X_FF DLX_EXinst_ALU_result_16 (
    .I(N120627),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_ALU_result<16>/FFY/RST ),
    .O(DLX_EXinst_ALU_result[16])
  );
  X_OR2 \DLX_EXinst_ALU_result<16>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_ALU_result<16>/FFY/RST )
  );
  defparam DLX_IDinst_reg_out_A_21.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_A_21 (
    .I(N104168),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_A<21>/FFY/RST ),
    .O(DLX_IDinst_reg_out_A[21])
  );
  X_OR2 \DLX_IDinst_reg_out_A<21>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_A<21>/FFY/RST )
  );
  defparam DLX_IDinst_reg_out_A_13.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_A_13 (
    .I(N103556),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_A<13>/FFY/RST ),
    .O(DLX_IDinst_reg_out_A[13])
  );
  X_OR2 \DLX_IDinst_reg_out_A<13>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_A<13>/FFY/RST )
  );
  defparam DLX_IFinst_NPC_5.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_5 (
    .I(\DLX_IFinst_NPC<5>/GROM ),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_NPC<5>/FFY/RST ),
    .O(DLX_IFinst_NPC[5])
  );
  X_OR2 \DLX_IFinst_NPC<5>/FFY/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_NPC<5>/FFY/RST )
  );
  defparam DLX_IFinst_NPC_6.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_6 (
    .I(\DLX_IFinst_NPC<6>/GROM ),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_NPC<6>/FFY/RST ),
    .O(DLX_IFinst_NPC[6])
  );
  X_OR2 \DLX_IFinst_NPC<6>/FFY/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_NPC<6>/FFY/RST )
  );
  defparam DLX_IDinst_reg_write_1214.INIT = 1'b0;
  X_FF DLX_IDinst_reg_write_1214 (
    .I(N110803),
    .CE(DLX_IDinst__n0422),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_write/FFY/RST ),
    .O(DLX_IDinst_reg_write)
  );
  X_OR2 \DLX_IDinst_reg_write/FFY/RSTOR  (
    .I0(reset_IBUF_3),
    .I1(GSR),
    .O(\DLX_IDinst_reg_write/FFY/RST )
  );
  defparam DLX_IDinst_counter_0.INIT = 1'b0;
  X_FF DLX_IDinst_counter_0 (
    .I(N107173),
    .CE(DLX_IDinst__n0440),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_counter<0>/FFY/RST ),
    .O(DLX_IDinst_counter[0])
  );
  X_OR2 \DLX_IDinst_counter<0>/FFY/RSTOR  (
    .I0(reset_IBUF_5),
    .I1(GSR),
    .O(\DLX_IDinst_counter<0>/FFY/RST )
  );
  defparam DLX_EXinst_ALU_result_28.INIT = 1'b0;
  X_FF DLX_EXinst_ALU_result_28 (
    .I(N121082),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_ALU_result<28>/FFY/RST ),
    .O(DLX_EXinst_ALU_result[28])
  );
  X_OR2 \DLX_EXinst_ALU_result<28>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_ALU_result<28>/FFY/RST )
  );
  defparam DLX_IFinst_NPC_19.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_19 (
    .I(DLX_IFinst__n0001[19]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_NPC<19>/FFY/RST ),
    .O(DLX_IFinst_NPC[19])
  );
  X_OR2 \DLX_IFinst_NPC<19>/FFY/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_NPC<19>/FFY/RST )
  );
  defparam DLX_IFinst_NPC_27.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_27 (
    .I(DLX_IFinst__n0001[27]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_NPC<27>/FFY/RST ),
    .O(DLX_IFinst_NPC[27])
  );
  X_OR2 \DLX_IFinst_NPC<27>/FFY/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_NPC<27>/FFY/RST )
  );
  defparam DLX_IFinst_NPC_7.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_7 (
    .I(\DLX_IFinst_NPC<7>/GROM ),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_NPC<7>/FFY/RST ),
    .O(DLX_IFinst_NPC[7])
  );
  X_OR2 \DLX_IFinst_NPC<7>/FFY/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_NPC<7>/FFY/RST )
  );
  defparam DLX_EXinst_ALU_result_29.INIT = 1'b0;
  X_FF DLX_EXinst_ALU_result_29 (
    .I(N122016),
    .CE(VCC),
    .CLK(DLX_clk_EX),
    .SET(GND),
    .RST(\DLX_EXinst_ALU_result<29>/FFY/RST ),
    .O(DLX_EXinst_ALU_result[29])
  );
  X_OR2 \DLX_EXinst_ALU_result<29>/FFY/RSTOR  (
    .I0(reset_IBUF),
    .I1(GSR),
    .O(\DLX_EXinst_ALU_result<29>/FFY/RST )
  );
  defparam DLX_IFinst_NPC_28.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_28 (
    .I(DLX_IFinst__n0001[28]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_NPC<28>/FFY/RST ),
    .O(DLX_IFinst_NPC[28])
  );
  X_OR2 \DLX_IFinst_NPC<28>/FFY/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_NPC<28>/FFY/RST )
  );
  defparam DLX_IFinst_NPC_8.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_8 (
    .I(\DLX_IFinst_NPC<8>/GROM ),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_NPC<8>/FFY/RST ),
    .O(DLX_IFinst_NPC[8])
  );
  X_OR2 \DLX_IFinst_NPC<8>/FFY/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_NPC<8>/FFY/RST )
  );
  defparam DLX_IFinst_NPC_29.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_29 (
    .I(DLX_IFinst__n0001[29]),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_NPC<29>/FFY/RST ),
    .O(DLX_IFinst_NPC[29])
  );
  X_OR2 \DLX_IFinst_NPC<29>/FFY/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_NPC<29>/FFY/RST )
  );
  defparam DLX_IDinst_reg_out_A_11.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_A_11 (
    .I(N103488),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_A<11>/FFY/RST ),
    .O(DLX_IDinst_reg_out_A[11])
  );
  X_OR2 \DLX_IDinst_reg_out_A<11>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_A<11>/FFY/RST )
  );
  defparam DLX_IDinst_reg_out_A_12.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_A_12 (
    .I(N103420),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_A<12>/FFY/RST ),
    .O(DLX_IDinst_reg_out_A[12])
  );
  X_OR2 \DLX_IDinst_reg_out_A<12>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_A<12>/FFY/RST )
  );
  defparam DLX_IDinst_reg_out_A_20.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_A_20 (
    .I(N104032),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_A<20>/FFY/RST ),
    .O(DLX_IDinst_reg_out_A[20])
  );
  X_OR2 \DLX_IDinst_reg_out_A<20>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_A<20>/FFY/RST )
  );
  defparam DLX_MEMinst_reg_write_MEM_1215.INIT = 1'b0;
  X_FF DLX_MEMinst_reg_write_MEM_1215 (
    .I(DLX_EXinst_reg_write_EX),
    .CE(VCC),
    .CLK(\DLX_MEMinst_reg_write_MEM/CKMUXNOT ),
    .SET(GND),
    .RST(\DLX_MEMinst_reg_write_MEM/FFY/RST ),
    .O(DLX_MEMinst_reg_write_MEM)
  );
  X_OR2 \DLX_MEMinst_reg_write_MEM/FFY/RSTOR  (
    .I0(reset_IBUF_1),
    .I1(GSR),
    .O(\DLX_MEMinst_reg_write_MEM/FFY/RST )
  );
  defparam DLX_IFinst_NPC_9.INIT = 1'b0;
  X_FF DLX_IFinst_NPC_9 (
    .I(\DLX_IFinst_NPC<9>/GROM ),
    .CE(VCC),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(\DLX_IFinst_NPC<9>/FFY/RST ),
    .O(DLX_IFinst_NPC[9])
  );
  X_OR2 \DLX_IFinst_NPC<9>/FFY/RSTOR  (
    .I0(reset_IBUF_2),
    .I1(GSR),
    .O(\DLX_IFinst_NPC<9>/FFY/RST )
  );
  defparam DLX_IDinst_reg_out_A_10.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_A_10 (
    .I(N103352),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_A<10>/FFY/RST ),
    .O(DLX_IDinst_reg_out_A[10])
  );
  X_OR2 \DLX_IDinst_reg_out_A<10>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_A<10>/FFY/RST )
  );
  defparam DLX_IFinst_IR_curr_10.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_10 (
    .I(IR[10]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[10])
  );
  defparam DLX_IFinst_IR_curr_11.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_11 (
    .I(IR[11]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[11])
  );
  defparam DLX_IFinst_IR_curr_1.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_1 (
    .I(IR[1]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[1])
  );
  defparam DLX_IFinst_IR_curr_0.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_0 (
    .I(IR[0]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[0])
  );
  defparam DLX_IFinst_IR_curr_21.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_21 (
    .I(IR[21]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[21])
  );
  defparam DLX_IFinst_IR_curr_20.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_20 (
    .I(IR[20]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[20])
  );
  defparam DLX_IFinst_IR_curr_13.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_13 (
    .I(IR[13]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[13])
  );
  defparam DLX_IFinst_IR_curr_12.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_12 (
    .I(IR[12]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[12])
  );
  defparam DLX_IFinst_IR_curr_3.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_3 (
    .I(IR[3]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[3])
  );
  defparam DLX_IFinst_IR_curr_2.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_2 (
    .I(IR[2]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[2])
  );
  defparam DLX_opcode_of_MEM_0.INIT = 1'b0;
  X_SFF DLX_opcode_of_MEM_0 (
    .I(DLX_IDinst_IR_opcode_field[0]),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_opcode_of_MEM[0])
  );
  defparam DLX_opcode_of_MEM_1.INIT = 1'b0;
  X_SFF DLX_opcode_of_MEM_1 (
    .I(DLX_IDinst_IR_opcode_field[1]),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_opcode_of_MEM[1])
  );
  defparam DLX_IFinst_IR_curr_31.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_31 (
    .I(IR_MSB_7_OBUF),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[31])
  );
  defparam DLX_IFinst_IR_curr_30.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_30 (
    .I(IR_MSB_6_OBUF),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[30])
  );
  defparam DLX_IFinst_IR_curr_23.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_23 (
    .I(IR[23]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[23])
  );
  defparam DLX_IFinst_IR_curr_22.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_22 (
    .I(IR[22]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[22])
  );
  defparam DLX_IFinst_IR_curr_15.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_15 (
    .I(IR[15]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[15])
  );
  defparam DLX_IFinst_IR_curr_14.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_14 (
    .I(IR[14]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[14])
  );
  defparam DLX_IDinst_reg_out_A_14.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_A_14 (
    .I(N103624),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_A<14>/FFY/RST ),
    .O(DLX_IDinst_reg_out_A[14])
  );
  X_OR2 \DLX_IDinst_reg_out_A<14>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_A<14>/FFY/RST )
  );
  defparam DLX_IFinst_IR_curr_5.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_5 (
    .I(IR[5]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[5])
  );
  defparam DLX_IFinst_IR_curr_4.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_4 (
    .I(IR[4]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[4])
  );
  defparam DLX_opcode_of_MEM_2.INIT = 1'b0;
  X_SFF DLX_opcode_of_MEM_2 (
    .I(DLX_IDinst_IR_opcode_field[2]),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_opcode_of_MEM[2])
  );
  defparam DLX_opcode_of_MEM_3.INIT = 1'b0;
  X_SFF DLX_opcode_of_MEM_3 (
    .I(DLX_IDinst_IR_opcode_field[3]),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_opcode_of_MEM[3])
  );
  defparam DLX_IDinst_reg_out_A_22.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_A_22 (
    .I(N104100),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_A<22>/FFY/RST ),
    .O(DLX_IDinst_reg_out_A[22])
  );
  X_OR2 \DLX_IDinst_reg_out_A<22>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_A<22>/FFY/RST )
  );
  defparam DLX_IDinst_reg_out_A_30.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_A_30 (
    .I(N104712),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_A<30>/FFY/RST ),
    .O(DLX_IDinst_reg_out_A[30])
  );
  X_OR2 \DLX_IDinst_reg_out_A<30>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_A<30>/FFY/RST )
  );
  defparam DLX_IFinst_IR_curr_24.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_24 (
    .I(IR_MSB_0_OBUF),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[24])
  );
  defparam DLX_IFinst_IR_curr_25.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_25 (
    .I(IR_MSB_1_OBUF),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[25])
  );
  defparam DLX_IFinst_IR_curr_17.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_17 (
    .I(IR[17]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[17])
  );
  defparam DLX_IFinst_IR_curr_16.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_16 (
    .I(IR[16]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[16])
  );
  defparam DLX_IFinst_IR_curr_7.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_7 (
    .I(IR[7]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[7])
  );
  defparam DLX_IFinst_IR_curr_6.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_6 (
    .I(IR[6]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[6])
  );
  defparam DLX_opcode_of_MEM_4.INIT = 1'b0;
  X_SFF DLX_opcode_of_MEM_4 (
    .I(DLX_IDinst_IR_opcode_field[4]),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_opcode_of_MEM[4])
  );
  defparam DLX_opcode_of_MEM_5.INIT = 1'b0;
  X_SFF DLX_opcode_of_MEM_5 (
    .I(DLX_IDinst_IR_opcode_field[5]),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_opcode_of_MEM[5])
  );
  defparam DLX_IFinst_IR_curr_26.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_26 (
    .I(IR_MSB_2_OBUF),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[26])
  );
  defparam DLX_IFinst_IR_curr_27.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_27 (
    .I(IR_MSB_3_OBUF),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[27])
  );
  defparam DLX_IFinst_IR_curr_19.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_19 (
    .I(IR[19]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[19])
  );
  defparam DLX_IFinst_IR_curr_18.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_18 (
    .I(IR[18]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[18])
  );
  defparam DLX_IFinst_IR_curr_9.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_9 (
    .I(IR[9]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[9])
  );
  defparam DLX_IFinst_IR_curr_8.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_8 (
    .I(IR[8]),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[8])
  );
  defparam DLX_IFinst_IR_curr_29.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_29 (
    .I(IR_MSB_5_OBUF),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[29])
  );
  defparam DLX_IFinst_IR_curr_28.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_28 (
    .I(IR_MSB_4_OBUF),
    .CE(DLX_IFinst_IR_curr_N3638),
    .CLK(DLX_clk_IF),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[28])
  );
  defparam DLX_IDinst_reg_out_A_23.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_A_23 (
    .I(N104236),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_A<23>/FFY/RST ),
    .O(DLX_IDinst_reg_out_A[23])
  );
  X_OR2 \DLX_IDinst_reg_out_A<23>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_A<23>/FFY/RST )
  );
  defparam DLX_IDinst_reg_out_A_31.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_A_31 (
    .I(N102604),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_A<31>/FFY/RST ),
    .O(DLX_IDinst_reg_out_A[31])
  );
  X_OR2 \DLX_IDinst_reg_out_A<31>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_A<31>/FFY/RST )
  );
  defparam DLX_IDinst_reg_out_A_15.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_A_15 (
    .I(N103692),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_A<15>/FFY/RST ),
    .O(DLX_IDinst_reg_out_A[15])
  );
  X_OR2 \DLX_IDinst_reg_out_A<15>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_A<15>/FFY/RST )
  );
  defparam DLX_IDinst_reg_out_A_0.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_A_0 (
    .I(N102740),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_A<0>/FFY/RST ),
    .O(DLX_IDinst_reg_out_A[0])
  );
  X_OR2 \DLX_IDinst_reg_out_A<0>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_A<0>/FFY/RST )
  );
  defparam DLX_IDinst_reg_out_A_24.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_A_24 (
    .I(N104372),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_A<24>/FFY/RST ),
    .O(DLX_IDinst_reg_out_A[24])
  );
  X_OR2 \DLX_IDinst_reg_out_A<24>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_A<24>/FFY/RST )
  );
  defparam DLX_IDinst_reg_out_A_16.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_A_16 (
    .I(N103828),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_A<16>/FFY/RST ),
    .O(DLX_IDinst_reg_out_A[16])
  );
  X_OR2 \DLX_IDinst_reg_out_A<16>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_A<16>/FFY/RST )
  );
  defparam DLX_IDinst_reg_out_A_1.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_A_1 (
    .I(N102672),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_A<1>/FFY/RST ),
    .O(DLX_IDinst_reg_out_A[1])
  );
  X_OR2 \DLX_IDinst_reg_out_A<1>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_A<1>/FFY/RST )
  );
  defparam DLX_IDinst_reg_out_A_17.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_A_17 (
    .I(N103760),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_A<17>/FFY/RST ),
    .O(DLX_IDinst_reg_out_A[17])
  );
  X_OR2 \DLX_IDinst_reg_out_A<17>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_A<17>/FFY/RST )
  );
  defparam DLX_IDinst_reg_out_A_25.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_A_25 (
    .I(N104304),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_A<25>/FFY/RST ),
    .O(DLX_IDinst_reg_out_A[25])
  );
  X_OR2 \DLX_IDinst_reg_out_A<25>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_A<25>/FFY/RST )
  );
  defparam DLX_IDinst_reg_out_A_2.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_A_2 (
    .I(N102808),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_A<2>/FFY/RST ),
    .O(DLX_IDinst_reg_out_A[2])
  );
  X_OR2 \DLX_IDinst_reg_out_A<2>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_A<2>/FFY/RST )
  );
  defparam DLX_IDinst_reg_out_A_26.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_A_26 (
    .I(N104440),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_A<26>/FFY/RST ),
    .O(DLX_IDinst_reg_out_A[26])
  );
  X_OR2 \DLX_IDinst_reg_out_A<26>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_A<26>/FFY/RST )
  );
  defparam DLX_IDinst_reg_out_A_18.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_A_18 (
    .I(N103896),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_A<18>/FFY/RST ),
    .O(DLX_IDinst_reg_out_A[18])
  );
  X_OR2 \DLX_IDinst_reg_out_A<18>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_A<18>/FFY/RST )
  );
  defparam DLX_IDinst_reg_out_A_3.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_A_3 (
    .I(N102944),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_A<3>/FFY/RST ),
    .O(DLX_IDinst_reg_out_A[3])
  );
  X_OR2 \DLX_IDinst_reg_out_A<3>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_A<3>/FFY/RST )
  );
  defparam DLX_IDinst_reg_out_A_27.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_A_27 (
    .I(N104576),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_A<27>/FFY/RST ),
    .O(DLX_IDinst_reg_out_A[27])
  );
  X_OR2 \DLX_IDinst_reg_out_A<27>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_A<27>/FFY/RST )
  );
  defparam DLX_IDinst_reg_out_A_19.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_A_19 (
    .I(N103964),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_A<19>/FFY/RST ),
    .O(DLX_IDinst_reg_out_A[19])
  );
  X_OR2 \DLX_IDinst_reg_out_A<19>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_A<19>/FFY/RST )
  );
  defparam DLX_IDinst_reg_out_A_4.INIT = 1'b0;
  X_FF DLX_IDinst_reg_out_A_4 (
    .I(N102876),
    .CE(VCC),
    .CLK(DLX_clk_ID),
    .SET(GND),
    .RST(\DLX_IDinst_reg_out_A<4>/FFY/RST ),
    .O(DLX_IDinst_reg_out_A[4])
  );
  X_OR2 \DLX_IDinst_reg_out_A<4>/FFY/RSTOR  (
    .I0(reset_IBUF_4),
    .I1(GSR),
    .O(\DLX_IDinst_reg_out_A<4>/FFY/RST )
  );
  X_IPAD \clk_vga/PAD  (
    .PAD(clk_vga)
  );
  X_CKBUF \clk_vga/BUF  (
    .I(clk_vga),
    .O(clkbuf)
  );
  X_CKBUF \DLX_clkbuf2/BUF  (
    .I(DLX_ackin_ID),
    .O(DLX_clk_ID)
  );
  X_CKBUF \DLX_clkbuf3/BUF  (
    .I(DLX_ackin_EX),
    .O(DLX_clk_EX)
  );
  X_CKBUF \clkbuf2/BUF  (
    .I(clk0),
    .O(clk0buf)
  );
  X_CKBUF \clkbuf3/BUF  (
    .I(clkdivub),
    .O(clkdiv_vga)
  );
  defparam \PWR_VCC_0/F .INIT = 16'hFFFF;
  X_LUT4 \PWR_VCC_0/F  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\PWR_VCC_0/FROM )
  );
  defparam \PWR_VCC_0/G .INIT = 16'h0000;
  X_LUT4 \PWR_VCC_0/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\PWR_VCC_0/GROM )
  );
  X_BUF \PWR_VCC_0/XUSED  (
    .I(\PWR_VCC_0/FROM ),
    .O(GLOBAL_LOGIC1)
  );
  X_BUF \PWR_VCC_0/YUSED  (
    .I(\PWR_VCC_0/GROM ),
    .O(GLOBAL_LOGIC0_10)
  );
  defparam \PWR_VCC_1/F .INIT = 16'hFFFF;
  X_LUT4 \PWR_VCC_1/F  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\PWR_VCC_1/FROM )
  );
  defparam \PWR_VCC_1/G .INIT = 16'h0000;
  X_LUT4 \PWR_VCC_1/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\PWR_VCC_1/GROM )
  );
  X_BUF \PWR_VCC_1/XUSED  (
    .I(\PWR_VCC_1/FROM ),
    .O(GLOBAL_LOGIC1_0)
  );
  X_BUF \PWR_VCC_1/YUSED  (
    .I(\PWR_VCC_1/GROM ),
    .O(GLOBAL_LOGIC0_8)
  );
  defparam \PWR_VCC_2/F .INIT = 16'hFFFF;
  X_LUT4 \PWR_VCC_2/F  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\PWR_VCC_2/FROM )
  );
  defparam \PWR_VCC_2/G .INIT = 16'h0000;
  X_LUT4 \PWR_VCC_2/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\PWR_VCC_2/GROM )
  );
  X_BUF \PWR_VCC_2/XUSED  (
    .I(\PWR_VCC_2/FROM ),
    .O(GLOBAL_LOGIC1_1)
  );
  X_BUF \PWR_VCC_2/YUSED  (
    .I(\PWR_VCC_2/GROM ),
    .O(GLOBAL_LOGIC0_7)
  );
  defparam \PWR_VCC_3/F .INIT = 16'hFFFF;
  X_LUT4 \PWR_VCC_3/F  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\PWR_VCC_3/FROM )
  );
  defparam \PWR_VCC_3/G .INIT = 16'h0000;
  X_LUT4 \PWR_VCC_3/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\PWR_VCC_3/GROM )
  );
  X_BUF \PWR_VCC_3/XUSED  (
    .I(\PWR_VCC_3/FROM ),
    .O(GLOBAL_LOGIC1_2)
  );
  X_BUF \PWR_VCC_3/YUSED  (
    .I(\PWR_VCC_3/GROM ),
    .O(GLOBAL_LOGIC0_6)
  );
  defparam \PWR_VCC_4/F .INIT = 16'hFFFF;
  X_LUT4 \PWR_VCC_4/F  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\PWR_VCC_4/FROM )
  );
  defparam \PWR_VCC_4/G .INIT = 16'h0000;
  X_LUT4 \PWR_VCC_4/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\PWR_VCC_4/GROM )
  );
  X_BUF \PWR_VCC_4/XUSED  (
    .I(\PWR_VCC_4/FROM ),
    .O(GLOBAL_LOGIC1_3)
  );
  X_BUF \PWR_VCC_4/YUSED  (
    .I(\PWR_VCC_4/GROM ),
    .O(GLOBAL_LOGIC0_5)
  );
  defparam \PWR_GND_0/G .INIT = 16'h0000;
  X_LUT4 \PWR_GND_0/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\PWR_GND_0/GROM )
  );
  X_BUF \PWR_GND_0/YUSED  (
    .I(\PWR_GND_0/GROM ),
    .O(GLOBAL_LOGIC0)
  );
  defparam \PWR_GND_1/G .INIT = 16'h0000;
  X_LUT4 \PWR_GND_1/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\PWR_GND_1/GROM )
  );
  X_BUF \PWR_GND_1/YUSED  (
    .I(\PWR_GND_1/GROM ),
    .O(GLOBAL_LOGIC0_0)
  );
  defparam \PWR_GND_2/G .INIT = 16'h0000;
  X_LUT4 \PWR_GND_2/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\PWR_GND_2/GROM )
  );
  X_BUF \PWR_GND_2/YUSED  (
    .I(\PWR_GND_2/GROM ),
    .O(GLOBAL_LOGIC0_1)
  );
  defparam \PWR_GND_3/G .INIT = 16'h0000;
  X_LUT4 \PWR_GND_3/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\PWR_GND_3/GROM )
  );
  X_BUF \PWR_GND_3/YUSED  (
    .I(\PWR_GND_3/GROM ),
    .O(GLOBAL_LOGIC0_2)
  );
  defparam \PWR_GND_4/G .INIT = 16'h0000;
  X_LUT4 \PWR_GND_4/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\PWR_GND_4/GROM )
  );
  X_BUF \PWR_GND_4/YUSED  (
    .I(\PWR_GND_4/GROM ),
    .O(GLOBAL_LOGIC0_3)
  );
  defparam \PWR_GND_5/G .INIT = 16'h0000;
  X_LUT4 \PWR_GND_5/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\PWR_GND_5/GROM )
  );
  X_BUF \PWR_GND_5/YUSED  (
    .I(\PWR_GND_5/GROM ),
    .O(GLOBAL_LOGIC0_4)
  );
  defparam \PWR_GND_6/G .INIT = 16'h0000;
  X_LUT4 \PWR_GND_6/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\PWR_GND_6/GROM )
  );
  X_BUF \PWR_GND_6/YUSED  (
    .I(\PWR_GND_6/GROM ),
    .O(GLOBAL_LOGIC0_9)
  );
  X_ONE NlwBlock_DLX_top_VCC (
    .O(VCC)
  );
  X_ZERO NlwBlock_DLX_top_GND (
    .O(GND)
  );
endmodule

