// Xilinx Verilog netlist produced by netgen application (version G.26)
// Command      : -intstyle ise -s 7 -pcf DLX_top.pcf -ngm DLX_top.ngm -w -ofmt verilog -sim DLX_top.ncd DLX_top_timesim.v 
// Input file   : DLX_top.ncd
// Output file  : DLX_top_timesim.v
// Design name  : DLX_top
// # of Modules : 1
// Xilinx       : /usr/local/vlsi/Xilinx-ISE-6.1
// Device       : 2s200epq208-7 (PRODUCTION 1.17 2003-11-04)

// This verilog netlist is a simulation model and uses simulation 
// primitives which may not represent the true implementation of the 
// device, however the netlist is functionally correct and should not 
// be modified. This file cannot be synthesized and should only be used 
// with supported simulation tools.

`timescale 1 ns/1 ps

module DLX_top (
  stall, branch_sig, hsync, DM_write, DM_write_data_0, DM_read, PIPEEMPTY, vsync, CLI, INT, FREEZE, reset, clk, DM_addr_eff, mask, red, NPC_eff, 
IR_MSB, green, blue
);
  output stall;
  output branch_sig;
  output hsync;
  output DM_write;
  output DM_write_data_0;
  output DM_read;
  output PIPEEMPTY;
  output vsync;
  output CLI;
  input INT;
  input FREEZE;
  input reset;
  input clk;
  output [14 : 0] DM_addr_eff;
  output [3 : 0] mask;
  output [1 : 0] red;
  output [15 : 0] NPC_eff;
  output [7 : 0] IR_MSB;
  output [2 : 0] green;
  output [2 : 0] blue;
  wire DLX_IDinst__n0600;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_971;
  wire clkdiv;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_973;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_583;
  wire DLX_IDinst_RegFile_24_28;
  wire DLX_IDinst_RegFile_25_28;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_584;
  wire DLX_IDinst_RegFile_26_28;
  wire DLX_IDinst_RegFile_27_28;
  wire reset_IBUF_8;
  wire DLX_IDinst__n0602;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_331;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_333;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_55;
  wire \DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ;
  wire DLX_IDinst_RegFile_24_20;
  wire DLX_IDinst_RegFile_25_20;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_56;
  wire DLX_IDinst_RegFile_26_20;
  wire DLX_IDinst_RegFile_27_20;
  wire reset_IBUF_7;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_203;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_205;
  wire \DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ;
  wire DLX_IDinst_RegFile_24_12;
  wire DLX_IDinst_RegFile_25_12;
  wire DLX_IDinst_RegFile_26_12;
  wire DLX_IDinst_RegFile_27_12;
  wire DLX_IDinst__n0584;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_983;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_985;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_579;
  wire \DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ;
  wire DLX_IDinst_RegFile_16_29;
  wire DLX_IDinst_RegFile_17_29;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_580;
  wire DLX_IDinst_RegFile_18_29;
  wire DLX_IDinst_RegFile_19_29;
  wire reset_IBUF_11;
  wire DLX_IDinst__n0586;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_343;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_345;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_51;
  wire DLX_IDinst_RegFile_16_21;
  wire DLX_IDinst_RegFile_17_21;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_52;
  wire DLX_IDinst_RegFile_18_21;
  wire DLX_IDinst_RegFile_19_21;
  wire reset_IBUF_10;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_215;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_217;
  wire \DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ;
  wire DLX_IDinst_RegFile_16_13;
  wire DLX_IDinst_RegFile_17_13;
  wire DLX_IDinst_RegFile_18_13;
  wire DLX_IDinst_RegFile_19_13;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_987;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_989;
  wire DLX_IDinst_RegFile_24_29;
  wire DLX_IDinst_RegFile_25_29;
  wire DLX_IDinst_RegFile_26_29;
  wire DLX_IDinst_RegFile_27_29;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_347;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_349;
  wire DLX_IDinst_RegFile_24_21;
  wire DLX_IDinst_RegFile_25_21;
  wire DLX_IDinst_RegFile_26_21;
  wire DLX_IDinst_RegFile_27_21;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_219;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_221;
  wire DLX_IDinst_RegFile_24_13;
  wire DLX_IDinst_RegFile_25_13;
  wire DLX_IDinst_RegFile_26_13;
  wire DLX_IDinst_RegFile_27_13;
  wire vga_top_vga1__n0029;
  wire vga_top_vga1__n0030;
  wire CHOICE3470;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_999;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_1001;
  wire DLX_IDinst_RegFile_16_30;
  wire DLX_IDinst_RegFile_17_30;
  wire DLX_IDinst_RegFile_18_30;
  wire DLX_IDinst_RegFile_19_30;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_359;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_361;
  wire DLX_IDinst_RegFile_16_22;
  wire DLX_IDinst_RegFile_17_22;
  wire DLX_IDinst_RegFile_18_22;
  wire DLX_IDinst_RegFile_19_22;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_231;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_233;
  wire DLX_IDinst_RegFile_16_14;
  wire DLX_IDinst_RegFile_17_14;
  wire DLX_IDinst_RegFile_18_14;
  wire DLX_IDinst_RegFile_19_14;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_1003;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_1005;
  wire DLX_IDinst_RegFile_24_30;
  wire DLX_IDinst_RegFile_25_30;
  wire DLX_IDinst_RegFile_26_30;
  wire DLX_IDinst_RegFile_27_30;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_363;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_365;
  wire DLX_IDinst_RegFile_24_22;
  wire DLX_IDinst_RegFile_25_22;
  wire DLX_IDinst_RegFile_26_22;
  wire DLX_IDinst_RegFile_27_22;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_235;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_237;
  wire DLX_IDinst_RegFile_24_14;
  wire DLX_IDinst_RegFile_25_14;
  wire DLX_IDinst_RegFile_26_14;
  wire DLX_IDinst_RegFile_27_14;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_375;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_377;
  wire DLX_IDinst_RegFile_16_23;
  wire DLX_IDinst_RegFile_17_23;
  wire DLX_IDinst_RegFile_18_23;
  wire DLX_IDinst_RegFile_19_23;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_247;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_249;
  wire DLX_IDinst_RegFile_16_15;
  wire DLX_IDinst_RegFile_17_15;
  wire DLX_IDinst_RegFile_18_15;
  wire DLX_IDinst_RegFile_19_15;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_891;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_893;
  wire \DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ;
  wire DLX_IDinst_RegFile_24_23;
  wire DLX_IDinst_RegFile_25_23;
  wire DLX_IDinst_RegFile_26_23;
  wire DLX_IDinst_RegFile_27_23;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_251;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_253;
  wire DLX_IDinst_RegFile_24_15;
  wire DLX_IDinst_RegFile_25_15;
  wire DLX_IDinst_RegFile_26_15;
  wire DLX_IDinst_RegFile_27_15;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_1015;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_1017;
  wire DLX_IDinst_RegFile_16_31;
  wire DLX_IDinst_RegFile_17_31;
  wire DLX_IDinst_RegFile_18_31;
  wire DLX_IDinst_RegFile_19_31;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_1019;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_1021;
  wire DLX_IDinst_RegFile_24_31;
  wire DLX_IDinst_RegFile_25_31;
  wire DLX_IDinst_RegFile_26_31;
  wire DLX_IDinst_RegFile_27_31;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_391;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_393;
  wire \DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ;
  wire DLX_IDinst_RegFile_16_24;
  wire DLX_IDinst_RegFile_17_24;
  wire DLX_IDinst_RegFile_18_24;
  wire DLX_IDinst_RegFile_19_24;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_263;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_265;
  wire DLX_IDinst_RegFile_16_16;
  wire DLX_IDinst_RegFile_17_16;
  wire DLX_IDinst_RegFile_18_16;
  wire DLX_IDinst_RegFile_19_16;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_395;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_397;
  wire DLX_IDinst_RegFile_24_24;
  wire DLX_IDinst_RegFile_25_24;
  wire DLX_IDinst_RegFile_26_24;
  wire DLX_IDinst_RegFile_27_24;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_267;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_269;
  wire DLX_IDinst_RegFile_24_16;
  wire DLX_IDinst_RegFile_25_16;
  wire DLX_IDinst_RegFile_26_16;
  wire DLX_IDinst_RegFile_27_16;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_407;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_409;
  wire DLX_IDinst_RegFile_16_25;
  wire DLX_IDinst_RegFile_17_25;
  wire DLX_IDinst_RegFile_18_25;
  wire DLX_IDinst_RegFile_19_25;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_279;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_281;
  wire DLX_IDinst_RegFile_16_17;
  wire DLX_IDinst_RegFile_17_17;
  wire DLX_IDinst_RegFile_18_17;
  wire DLX_IDinst_RegFile_19_17;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_411;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_413;
  wire DLX_IDinst_RegFile_24_25;
  wire DLX_IDinst_RegFile_25_25;
  wire DLX_IDinst_RegFile_26_25;
  wire DLX_IDinst_RegFile_27_25;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_283;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_285;
  wire DLX_IDinst_RegFile_24_17;
  wire DLX_IDinst_RegFile_25_17;
  wire DLX_IDinst_RegFile_26_17;
  wire DLX_IDinst_RegFile_27_17;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_423;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_425;
  wire DLX_IDinst_RegFile_16_26;
  wire DLX_IDinst_RegFile_17_26;
  wire DLX_IDinst_RegFile_18_26;
  wire DLX_IDinst_RegFile_19_26;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_295;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_297;
  wire DLX_IDinst_RegFile_16_18;
  wire DLX_IDinst_RegFile_17_18;
  wire DLX_IDinst_RegFile_18_18;
  wire DLX_IDinst_RegFile_19_18;
  wire DLX_IDinst__n0588;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_167;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_169;
  wire DLX_IDinst_RegFile_16_10;
  wire DLX_IDinst_RegFile_17_10;
  wire DLX_IDinst_RegFile_18_10;
  wire DLX_IDinst_RegFile_19_10;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_427;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_429;
  wire DLX_IDinst_RegFile_24_26;
  wire DLX_IDinst_RegFile_25_26;
  wire DLX_IDinst_RegFile_26_26;
  wire DLX_IDinst_RegFile_27_26;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_299;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_301;
  wire DLX_IDinst_RegFile_24_18;
  wire DLX_IDinst_RegFile_25_18;
  wire DLX_IDinst_RegFile_26_18;
  wire DLX_IDinst_RegFile_27_18;
  wire DLX_IDinst__n0604;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_171;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_173;
  wire DLX_IDinst_RegFile_24_10;
  wire DLX_IDinst_RegFile_25_10;
  wire DLX_IDinst_RegFile_26_10;
  wire DLX_IDinst_RegFile_27_10;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_951;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_953;
  wire DLX_IDinst_RegFile_16_27;
  wire DLX_IDinst_RegFile_17_27;
  wire DLX_IDinst_RegFile_18_27;
  wire DLX_IDinst_RegFile_19_27;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_311;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_313;
  wire DLX_IDinst_RegFile_16_19;
  wire DLX_IDinst_RegFile_17_19;
  wire DLX_IDinst_RegFile_18_19;
  wire DLX_IDinst_RegFile_19_19;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_183;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_185;
  wire DLX_IDinst_RegFile_16_11;
  wire DLX_IDinst_RegFile_17_11;
  wire DLX_IDinst_RegFile_18_11;
  wire DLX_IDinst_RegFile_19_11;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_955;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_957;
  wire DLX_IDinst_RegFile_24_27;
  wire DLX_IDinst_RegFile_25_27;
  wire DLX_IDinst_RegFile_26_27;
  wire DLX_IDinst_RegFile_27_27;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_315;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_317;
  wire DLX_IDinst_RegFile_24_19;
  wire DLX_IDinst_RegFile_25_19;
  wire DLX_IDinst_RegFile_26_19;
  wire DLX_IDinst_RegFile_27_19;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_187;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_189;
  wire DLX_IDinst_RegFile_24_11;
  wire DLX_IDinst_RegFile_25_11;
  wire DLX_IDinst_RegFile_26_11;
  wire DLX_IDinst_RegFile_27_11;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_967;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_969;
  wire DLX_IDinst_RegFile_16_28;
  wire DLX_IDinst_RegFile_17_28;
  wire DLX_IDinst_RegFile_18_28;
  wire DLX_IDinst_RegFile_19_28;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_327;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_329;
  wire DLX_IDinst_RegFile_16_20;
  wire DLX_IDinst_RegFile_17_20;
  wire DLX_IDinst_RegFile_18_20;
  wire DLX_IDinst_RegFile_19_20;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_199;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_201;
  wire DLX_IDinst_RegFile_16_12;
  wire DLX_IDinst_RegFile_17_12;
  wire DLX_IDinst_RegFile_18_12;
  wire DLX_IDinst_RegFile_19_12;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_459;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_461;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_843;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_845;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_715;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_717;
  wire \DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_471;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_473;
  wire \DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_855;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_857;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_727;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_729;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_475;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_477;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_859;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_861;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_731;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_733;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_487;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_489;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_871;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_873;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_743;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_745;
  wire \DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_491;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_493;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_875;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_877;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_747;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_749;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_887;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_889;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_759;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_761;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_763;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_765;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_503;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_505;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_507;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_509;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_903;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_905;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_775;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_777;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_907;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_909;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_779;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_781;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_919;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_921;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_791;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_793;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_795;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_797;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_935;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_937;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_807;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_809;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_939;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_941;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_811;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_813;
  wire DLX_IDinst__n0606;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_57;
  wire DLX_IDinst_RegFile_28_10;
  wire DLX_IDinst_RegFile_29_10;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_58;
  wire DLX_IDinst_RegFile_30_10;
  wire DLX_IDinst_RegFile_31_10;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_439;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_441;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_823;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_825;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_443;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_445;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_827;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_829;
  wire DLX_IDinst_RegFile_28_11;
  wire DLX_IDinst_RegFile_29_11;
  wire DLX_IDinst_RegFile_30_11;
  wire DLX_IDinst_RegFile_31_11;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_455;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_457;
  wire DLX_IDinst_RegFile_28_20;
  wire DLX_IDinst_RegFile_29_20;
  wire DLX_IDinst_RegFile_30_20;
  wire DLX_IDinst_RegFile_31_20;
  wire DLX_IDinst_RegFile_28_12;
  wire DLX_IDinst_RegFile_29_12;
  wire DLX_IDinst_RegFile_30_12;
  wire DLX_IDinst_RegFile_31_12;
  wire DLX_IDinst_RegFile_28_21;
  wire DLX_IDinst_RegFile_29_21;
  wire DLX_IDinst_RegFile_30_21;
  wire DLX_IDinst_RegFile_31_21;
  wire DLX_IDinst_RegFile_28_13;
  wire DLX_IDinst_RegFile_29_13;
  wire DLX_IDinst_RegFile_30_13;
  wire DLX_IDinst_RegFile_31_13;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_585;
  wire DLX_IDinst_RegFile_28_30;
  wire DLX_IDinst_RegFile_29_30;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_586;
  wire DLX_IDinst_RegFile_30_30;
  wire DLX_IDinst_RegFile_31_30;
  wire DLX_IDinst_RegFile_28_22;
  wire DLX_IDinst_RegFile_29_22;
  wire DLX_IDinst_RegFile_30_22;
  wire DLX_IDinst_RegFile_31_22;
  wire DLX_IDinst_RegFile_28_14;
  wire DLX_IDinst_RegFile_29_14;
  wire DLX_IDinst_RegFile_30_14;
  wire DLX_IDinst_RegFile_31_14;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_381;
  wire DLX_IDinst_RegFile_28_23;
  wire DLX_IDinst_RegFile_29_23;
  wire DLX_IDinst_RegFile_30_23;
  wire DLX_IDinst_RegFile_31_23;
  wire DLX_IDinst_RegFile_28_15;
  wire DLX_IDinst_RegFile_29_15;
  wire DLX_IDinst_RegFile_30_15;
  wire DLX_IDinst_RegFile_31_15;
  wire DLX_IDinst_RegFile_28_31;
  wire DLX_IDinst_RegFile_29_31;
  wire DLX_IDinst_RegFile_30_31;
  wire DLX_IDinst_RegFile_31_31;
  wire DLX_IDinst_RegFile_28_24;
  wire DLX_IDinst_RegFile_29_24;
  wire DLX_IDinst_RegFile_30_24;
  wire DLX_IDinst_RegFile_31_24;
  wire DLX_IDinst_RegFile_28_16;
  wire DLX_IDinst_RegFile_29_16;
  wire DLX_IDinst_RegFile_30_16;
  wire DLX_IDinst_RegFile_31_16;
  wire DLX_IDinst_RegFile_28_25;
  wire DLX_IDinst_RegFile_29_25;
  wire DLX_IDinst_RegFile_30_25;
  wire DLX_IDinst_RegFile_31_25;
  wire DLX_IDinst_RegFile_28_17;
  wire DLX_IDinst_RegFile_29_17;
  wire DLX_IDinst_RegFile_30_17;
  wire DLX_IDinst_RegFile_31_17;
  wire DLX_IDinst_RegFile_28_26;
  wire DLX_IDinst_RegFile_29_26;
  wire DLX_IDinst_RegFile_30_26;
  wire DLX_IDinst_RegFile_31_26;
  wire DLX_IDinst_RegFile_28_18;
  wire DLX_IDinst_RegFile_29_18;
  wire DLX_IDinst_RegFile_30_18;
  wire DLX_IDinst_RegFile_31_18;
  wire DLX_IDinst__n0608;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_685;
  wire DLX_IDinst_RegFile_28_27;
  wire DLX_IDinst_RegFile_29_27;
  wire DLX_IDinst_RegFile_30_27;
  wire DLX_IDinst_RegFile_31_27;
  wire DLX_IDinst_RegFile_28_19;
  wire DLX_IDinst_RegFile_29_19;
  wire DLX_IDinst_RegFile_30_19;
  wire DLX_IDinst_RegFile_31_19;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_701;
  wire DLX_IDinst_RegFile_28_28;
  wire DLX_IDinst_RegFile_29_28;
  wire DLX_IDinst_RegFile_30_28;
  wire DLX_IDinst_RegFile_31_28;
  wire reset_IBUF_6;
  wire DLX_IDinst_RegFile_28_29;
  wire DLX_IDinst_RegFile_29_29;
  wire DLX_IDinst_RegFile_30_29;
  wire DLX_IDinst_RegFile_31_29;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_925;
  wire \DLX_IDinst_Imm[4] ;
  wire \DLX_IDinst_Imm[2] ;
  wire \DLX_IDinst_Imm[3] ;
  wire \DLX_IDinst_Imm[1] ;
  wire DLX_EXinst__n0127;
  wire CHOICE2089;
  wire CHOICE3008;
  wire CHOICE3010;
  wire CHOICE3575;
  wire CHOICE3576;
  wire \DLX_IDinst_Imm[14] ;
  wire \DLX_IDinst_Imm[13] ;
  wire \DLX_IDinst_Imm[12] ;
  wire \DLX_IDinst_Imm[11] ;
  wire \DLX_IDinst_Imm[15] ;
  wire CHOICE3442;
  wire CHOICE3272;
  wire DLX_IFinst_IR_curr_N3087;
  wire reset_IBUF_2;
  wire CHOICE3639;
  wire CHOICE3587;
  wire DLX_IDinst__n0552;
  wire \DLX_IDinst_Imm[10] ;
  wire \DLX_IDinst_Imm[9] ;
  wire \DLX_IDinst_Imm[8] ;
  wire \DLX_IDinst_Imm[31] ;
  wire CHOICE3275;
  wire N163162;
  wire DLX_IDinst_RegFile_1_28;
  wire \DLX_IDinst_Imm[7] ;
  wire \DLX_IDinst_Imm[6] ;
  wire \DLX_IDinst_Imm[5] ;
  wire DLX_EXinst_N76041;
  wire N146478;
  wire DLX_EXinst__n0006;
  wire DLX_EXinst_N76441;
  wire CHOICE3631;
  wire CHOICE3583;
  wire DLX_IDinst_RegFile_1_29;
  wire CHOICE3590;
  wire N163386;
  wire DLX_EXinst__n0081;
  wire CHOICE3570;
  wire CHOICE3592;
  wire DLX_EXinst_N76421;
  wire DLX_IDinst__n0594;
  wire N138371;
  wire N148609;
  wire N163696;
  wire N148323;
  wire reset_IBUF_9;
  wire CHOICE5342;
  wire DLX_IDinst_RegFile_22_20;
  wire \DLX_IDinst_Imm[0] ;
  wire N163298;
  wire CHOICE1311;
  wire CHOICE1313;
  wire CHOICE1299;
  wire N134884;
  wire DLX_IDinst__n0116;
  wire DLX_IDinst_N108165;
  wire N139656;
  wire N132373;
  wire DLX_IDinst__n0453;
  wire DLX_IDinst_N108456;
  wire DLX_IDinst__n0115;
  wire DLX_IDinst_slot_num_FFd4;
  wire DLX_IDinst_delay_slot;
  wire DLX_IDinst_intr_slot;
  wire DLX_IDinst_slot_num_FFd1;
  wire DLX_EXinst__n0144;
  wire DLX_IDinst_slot_num_FFd2;
  wire DLX_IDinst_slot_num_FFd3;
  wire N163469;
  wire CHOICE2993;
  wire DLX_IDinst_N107033;
  wire N164150;
  wire DLX_IDinst_N107405;
  wire N127652;
  wire N132324;
  wire DLX_IDinst_Ker1084541_1;
  wire CHOICE2119;
  wire N127400;
  wire DLX_IDinst_Imm_0_1;
  wire DLX_IDinst__n0554;
  wire N163132;
  wire CHOICE3000;
  wire DLX_IDinst_RegFile_2_6;
  wire DLX_EXinst_byte;
  wire DLX_EXinst_word;
  wire N164178;
  wire mask_1_OBUF;
  wire DLX_IFinst_PC_N3087;
  wire reset_IBUF_1;
  wire DLX_IDinst_Imm_1_1;
  wire DLX_IDinst_Imm_2_1;
  wire \DLX_EXinst_Mshift__n0020_Sh[30] ;
  wire \DLX_EXinst_Mshift__n0020_Sh[26] ;
  wire CHOICE1865;
  wire \DLX_EXinst_Mshift__n0020_Sh[61] ;
  wire CHOICE1915;
  wire DLX_EXinst_N72791;
  wire DLX_EXinst_N72815;
  wire \DLX_EXinst_Mshift__n0020_Sh[29] ;
  wire CHOICE2017;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_572;
  wire DLX_IDinst_RegFile_2_19;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_581;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_582;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_573;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_578;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_574;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_577;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_575;
  wire \DLX_IDinst_Cause_Reg[31] ;
  wire CHOICE3230;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_576;
  wire DLX_IDinst_RegFile_2_27;
  wire DLX_IDinst_Imm_3_1;
  wire DLX_EXinst_N73379;
  wire DLX_EXinst_N76382;
  wire \DLX_EXinst_Mshift__n0020_Sh[88] ;
  wire CHOICE5185;
  wire DLX_IDinst__n0530;
  wire FREEZE_IBUF;
  wire N146700;
  wire DLX_IDinst_N108100;
  wire CHOICE2131;
  wire CHOICE2128;
  wire CHOICE2136;
  wire reset_IBUF_3;
  wire DLX_IDinst__n0580;
  wire vga_top_vga1_videoon;
  wire vram_out_vga_eff;
  wire blue_2_OBUF;
  wire green_0_OBUF;
  wire DLX_IDinst_RegFile_15_16;
  wire DLX_IDinst_Imm_31_1;
  wire DLX_EXinst_Mcompar__n0067_inst_cy_228;
  wire DLX_EXinst_Mcompar__n0067_inst_cy_229;
  wire DLX_EXinst__n0059;
  wire CHOICE5958;
  wire DLX_IDinst_RegFile_26_5;
  wire CHOICE2981;
  wire N164719;
  wire CHOICE2984;
  wire blue_0_OBUF;
  wire green_2_OBUF;
  wire DLX_IDinst_RegFile_2_21;
  wire DLX_MEMinst_noop;
  wire DLX_EXinst_noop;
  wire N139488;
  wire PIPEEMPTY_OBUF;
  wire DLX_EXinst_N73464;
  wire DLX_EXinst_N72938;
  wire \DLX_EXinst_Mshift__n0021_Sh[14] ;
  wire \DLX_EXinst_Mshift__n0021_Sh[10] ;
  wire N130311;
  wire DLX_IDinst_RegFile_2_13;
  wire DLX_EXinst_N72943;
  wire \DLX_EXinst_Mshift__n0021_Sh[15] ;
  wire \DLX_EXinst_Mshift__n0021_Sh[11] ;
  wire N130415;
  wire DLX_IDinst_RegFile_1_1;
  wire DLX_IDinst__n0572;
  wire DLX_EXinst_N73499;
  wire DLX_EXinst_N72973;
  wire \DLX_EXinst_Mshift__n0021_Sh[20] ;
  wire \DLX_EXinst_Mshift__n0021_Sh[24] ;
  wire reset_IBUF_13;
  wire CHOICE5667;
  wire DLX_IDinst_RegFile_11_21;
  wire DLX_EXinst_N73479;
  wire DLX_EXinst_N72953;
  wire \DLX_EXinst_Mshift__n0021_Sh[16] ;
  wire DLX_EXinst_N75377;
  wire DLX_IDinst_RegFile_2_22;
  wire DLX_EXinst_N72963;
  wire DLX_EXinst_N73484;
  wire CHOICE1727;
  wire \DLX_EXinst_Mshift__n0021_Sh[19] ;
  wire N137282;
  wire DLX_IDinst_RegFile_15_5;
  wire DLX_EXinst_N73519;
  wire DLX_EXinst_N73128;
  wire CHOICE1791;
  wire \DLX_EXinst_Mshift__n0022_Sh[12] ;
  wire N137680;
  wire \DLX_EXinst_Mshift__n0022_Sh[30] ;
  wire \DLX_EXinst_Mshift__n0022_Sh[58] ;
  wire DLX_EXinst_N73544;
  wire DLX_EXinst_N73153;
  wire \DLX_EXinst_Mshift__n0022_Sh[22] ;
  wire DLX_EXinst_N73163;
  wire DLX_IDinst_RegFile_2_23;
  wire DLX_EXinst_N73897;
  wire DLX_EXinst_N73211;
  wire \DLX_EXinst_Mshift__n0022_Sh[23] ;
  wire DLX_EXinst_N73168;
  wire DLX_IDinst_RegFile_2_15;
  wire DLX_IDinst__n0550;
  wire DLX_EXinst_N73529;
  wire DLX_EXinst_N73138;
  wire \DLX_EXinst_Mshift__n0022_Sh[8] ;
  wire \DLX_EXinst_Mshift__n0022_Sh[16] ;
  wire DLX_EXinst_N74946;
  wire DLX_IDinst_RegFile_0_12;
  wire DLX_IDinst__n0596;
  wire DLX_EXinst_N73534;
  wire \DLX_EXinst_Mshift__n0022_Sh[17] ;
  wire \DLX_EXinst_Mshift__n0020_Sh[25] ;
  wire DLX_EXinst_N74981;
  wire DLX_IDinst_RegFile_23_30;
  wire DLX_EXinst_N74986;
  wire CHOICE5220;
  wire DLX_EXinst__n0056;
  wire \DLX_EXinst_Mshift__n0022_Sh[50] ;
  wire N163424;
  wire DLX_IDinst_RegFile_2_24;
  wire DLX_EXinst_N73143;
  wire \DLX_EXinst_Mshift__n0022_Sh[18] ;
  wire DLX_IDinst_RegFile_2_16;
  wire DLX_IDinst__n0582;
  wire DLX_EXinst_N75352;
  wire CHOICE5299;
  wire \DLX_EXinst_Mshift__n0022_Sh[51] ;
  wire N163558;
  wire \DLX_EXinst_Mshift__n0022_Sh[29] ;
  wire CHOICE5076;
  wire \DLX_EXinst_Mshift__n0022_Sh[57] ;
  wire N163610;
  wire DLX_IDinst_RegFile_2_17;
  wire DLX_EXinst_N73158;
  wire CHOICE5378;
  wire \DLX_EXinst_Mshift__n0022_Sh[49] ;
  wire N163635;
  wire DLX_IDinst_RegFile_22_6;
  wire DLX_IDinst_branch_sig;
  wire DLX_IDinst_N108152;
  wire DLX_IDinst_N108465;
  wire CHOICE3348;
  wire N163562;
  wire DLX_IDinst_RegFile_1_23;
  wire DLX_EXinst_N76124;
  wire \DLX_EXinst_Mshift__n0020_Sh[127] ;
  wire CHOICE4308;
  wire DLX_EXinst_N73594;
  wire DLX_EXinst_N72888;
  wire \DLX_EXinst_Mshift__n0023_Sh[20] ;
  wire \DLX_EXinst_Mshift__n0023_Sh[24] ;
  wire CHOICE5617;
  wire DLX_IDinst_RegFile_11_24;
  wire DLX_IDinst__n0562;
  wire DLX_EXinst_N73574;
  wire DLX_EXinst_N72868;
  wire DLX_IDinst_reg_out_B_2_1;
  wire \DLX_EXinst_Mshift__n0023_Sh[16] ;
  wire reset_IBUF_4;
  wire DLX_EXinst_N75006;
  wire DLX_IDinst_RegFile_6_6;
  wire DLX_EXinst_N72878;
  wire DLX_EXinst_N73579;
  wire CHOICE1765;
  wire \DLX_EXinst_Mshift__n0023_Sh[19] ;
  wire N137518;
  wire DLX_EXinst__n0036;
  wire DLX_EXinst_N76501;
  wire DLX_IDinst_RegFile_15_9;
  wire DLX_IDinst__n0175;
  wire DLX_IDinst_N107837;
  wire CHOICE2235;
  wire \DLX_IDinst_regA_eff[10] ;
  wire DLX_IDinst_RegFile_1_26;
  wire N130927;
  wire CHOICE2246;
  wire \DLX_IDinst_regA_eff[11] ;
  wire DLX_IDinst_RegFile_26_2;
  wire \DLX_EXinst_Mshift__n0023_Sh[6] ;
  wire \DLX_EXinst_Mshift__n0023_Sh[2] ;
  wire DLX_EXinst_N72908;
  wire DLX_IDinst_RegFile_22_13;
  wire DLX_IDinst__n0610;
  wire CHOICE2257;
  wire \DLX_IDinst_regA_eff[12] ;
  wire DLX_IDinst__n0556;
  wire \DLX_IDinst_regA_eff[17] ;
  wire \DLX_IDinst_regA_eff[18] ;
  wire \DLX_IDinst_regA_eff[19] ;
  wire \DLX_IDinst_regA_eff[20] ;
  wire reset_IBUF_5;
  wire CHOICE4240;
  wire DLX_IDinst_RegFile_3_13;
  wire N163790;
  wire DLX_IDinst_RegFile_3_21;
  wire CHOICE2268;
  wire \DLX_IDinst_regA_eff[13] ;
  wire DLX_IDinst_RegFile_2_29;
  wire CHOICE2368;
  wire \DLX_IDinst_regA_eff[21] ;
  wire DLX_IDinst_RegFile_23_23;
  wire DLX_IDinst_reg_out_B_3_1;
  wire DLX_EXinst_N75964;
  wire DLX_IDinst_RegFile_3_22;
  wire CHOICE2279;
  wire \DLX_IDinst_regA_eff[14] ;
  wire DLX_IDinst_RegFile_23_17;
  wire CHOICE2379;
  wire \DLX_IDinst_regA_eff[22] ;
  wire DLX_IDinst_RegFile_18_4;
  wire CHOICE2390;
  wire \DLX_IDinst_regA_eff[30] ;
  wire DLX_IDinst_RegFile_3_15;
  wire DLX_EXinst_N76034;
  wire CHOICE2290;
  wire \DLX_IDinst_regA_eff[15] ;
  wire DLX_IDinst_RegFile_3_31;
  wire CHOICE2467;
  wire \DLX_IDinst_regA_eff[23] ;
  wire DLX_IDinst_RegFile_29_7;
  wire DLX_IDinst_RegFile_1_0;
  wire \DLX_IDinst_regA_eff[16] ;
  wire CHOICE4233;
  wire DLX_IDinst_RegFile_3_24;
  wire \DLX_IDinst_regA_eff[24] ;
  wire CHOICE4248;
  wire DLX_IDinst_RegFile_3_17;
  wire DLX_IDinst_RegFile_3_25;
  wire CHOICE2324;
  wire CHOICE2445;
  wire \DLX_IDinst_regA_eff[25] ;
  wire CHOICE5771;
  wire CHOICE5871;
  wire CHOICE2335;
  wire CHOICE2434;
  wire \DLX_IDinst_regA_eff[26] ;
  wire CHOICE2346;
  wire DLX_EXinst_N76463;
  wire \DLX_EXinst_Mshift__n0021_Sh[2] ;
  wire \DLX_EXinst_Mshift__n0021_Sh[1] ;
  wire CHOICE5511;
  wire CHOICE5690;
  wire \DLX_IDinst_regA_eff[27] ;
  wire \DLX_IDinst_regA_eff[28] ;
  wire CHOICE4255;
  wire CHOICE2401;
  wire \DLX_IDinst_regA_eff[29] ;
  wire \DLX_EXinst_Mshift__n0021_Sh[3] ;
  wire DLX_EXinst_N76285;
  wire CHOICE5435;
  wire CHOICE5437;
  wire vga_top_vga1_N112941;
  wire vga_top_vga1_helpme;
  wire N164108;
  wire vga_top_vga1__n0011;
  wire vga_top_vga1_N112904;
  wire vga_top_vga1_N112946;
  wire N127166;
  wire vga_top_vga1__n0012;
  wire \DLX_EXinst_Mshift__n0024_Sh[30] ;
  wire \DLX_EXinst_Mshift__n0019_Sh[26] ;
  wire \DLX_EXinst_Mshift__n0024_Sh[58] ;
  wire \DLX_EXinst_Mshift__n0024_Sh[31] ;
  wire \DLX_EXinst_Mshift__n0019_Sh[27] ;
  wire \DLX_EXinst_Mshift__n0024_Sh[59] ;
  wire DLX_EXinst_N74976;
  wire DLX_EXinst_N73103;
  wire CHOICE5337;
  wire \DLX_EXinst_Mshift__n0024_Sh[51] ;
  wire vga_top_vga1_N112936;
  wire N132499;
  wire vga_top_vga1__n0006;
  wire vga_top_vga1_N112910;
  wire N136799;
  wire vga_top_vga1__n0007;
  wire \DLX_EXinst_Mshift__n0024_Sh[29] ;
  wire \DLX_EXinst_Mshift__n0019_Sh[25] ;
  wire CHOICE2040;
  wire \DLX_EXinst_Mshift__n0024_Sh[57] ;
  wire DLX_EXinst_N74726;
  wire DLX_EXinst_N73093;
  wire CHOICE5416;
  wire \DLX_EXinst_Mshift__n0024_Sh[49] ;
  wire N163598;
  wire DLX_IDinst_RegFile_3_20;
  wire N130569;
  wire \DLX_EXinst_Mshift__n0019_Sh[22] ;
  wire DLX_EXinst_N74441;
  wire N131027;
  wire N164125;
  wire mask_0_OBUF;
  wire DLX_EXinst_N73267;
  wire DLX_EXinst_N76412;
  wire N132037;
  wire N131955;
  wire DLX_IDinst_RegFile_18_1;
  wire N164115;
  wire mask_3_OBUF;
  wire CHOICE1346;
  wire N132091;
  wire DLX_EXinst_reg_write_EX;
  wire DLX_MEMinst_reg_write_MEM;
  wire DLX_IDinst_N108538;
  wire DLX_IDinst__n0578;
  wire DLX_EXinst_N73345;
  wire N126741;
  wire reset_IBUF_12;
  wire DLX_EXinst__n0109;
  wire DLX_IDinst_RegFile_14_23;
  wire DLX_EXinst_N76490;
  wire CHOICE5824;
  wire N132064;
  wire DLX_IDinst_N108496;
  wire CHOICE3352;
  wire CHOICE3359;
  wire CHOICE3361;
  wire N146990;
  wire N163128;
  wire CHOICE2301;
  wire N140698;
  wire N164702;
  wire CHOICE2303;
  wire DLX_IDinst__n0570;
  wire DLX_IDinst_RegFile_10_6;
  wire N163842;
  wire CHOICE3328;
  wire DLX_IDinst__n0462;
  wire CHOICE3335;
  wire CHOICE3337;
  wire DLX_IDinst_RegFile_11_2;
  wire DLX_IDinst__n0167;
  wire DLX_IDinst__n0433;
  wire DLX_IDinst__n0436;
  wire DLX_IDinst__n0434;
  wire DLX_IDinst__n0166;
  wire CHOICE3508;
  wire CHOICE3515;
  wire N163554;
  wire DLX_IDinst__n0437;
  wire DLX_IDinst__n0439;
  wire DLX_IDinst_N108443;
  wire CHOICE3552;
  wire CHOICE3547;
  wire CHOICE3553;
  wire DLX_IDinst_N108264;
  wire DLX_IDinst_N108244;
  wire N164734;
  wire N163836;
  wire DLX_EXinst_N72710;
  wire N136586;
  wire DLX_EXinst_N74347;
  wire DLX_IDinst_N107572;
  wire DLX_IDinst__n0100;
  wire DLX_IDinst__n0382;
  wire CHOICE3524;
  wire CHOICE3526;
  wire N137212;
  wire N138903;
  wire DLX_IDinst_N108238;
  wire N135079;
  wire CHOICE2911;
  wire CHOICE3490;
  wire DLX_IDinst_RegFile_1_5;
  wire DLX_IDinst_N108476;
  wire N127043;
  wire DLX_IDinst__n0427;
  wire DLX_IDinst__n0164;
  wire DLX_IDinst_zflag;
  wire DLX_IDinst_N108221;
  wire N163831;
  wire DLX_IDinst_RegFile_22_11;
  wire DLX_IDinst__n0614;
  wire CHOICE3487;
  wire CHOICE3495;
  wire DLX_IDinst__n0637;
  wire CHOICE3493;
  wire N147786;
  wire DLX_IDinst_stall;
  wire CHOICE3624;
  wire CHOICE3647;
  wire CHOICE3600;
  wire CHOICE3616;
  wire N163733;
  wire N163574;
  wire CHOICE4196;
  wire IR_MSB_4_OBUF;
  wire N163724;
  wire CHOICE4202;
  wire CHOICE1971;
  wire CHOICE1987;
  wire CHOICE1989;
  wire \DLX_IDinst_regA_eff[3] ;
  wire CHOICE4208;
  wire \DLX_IDinst_regA_eff[1] ;
  wire CHOICE4209;
  wire N131907;
  wire DLX_EXinst__n0083;
  wire DLX_IDinst_reg_dst;
  wire CHOICE1338;
  wire N164077;
  wire CHOICE2873;
  wire DLX_IDinst__n0387;
  wire reset_IBUF_14;
  wire DLX_IDinst_N107105;
  wire CHOICE2148;
  wire IR_MSB_5_OBUF;
  wire CHOICE2159;
  wire \DLX_IDinst_regA_eff[2] ;
  wire CHOICE2170;
  wire DLX_IDinst__n0098;
  wire N127094;
  wire DLX_IDinst__n0176;
  wire DLX_IDinst_N107173;
  wire CHOICE2181;
  wire \DLX_IDinst_regA_eff[4] ;
  wire N147200;
  wire DLX_IDinst__n0376;
  wire N132648;
  wire DLX_IDinst_N108233;
  wire CHOICE2192;
  wire \DLX_IDinst_regA_eff[5] ;
  wire N163652;
  wire \DLX_IDinst_regA_eff[7] ;
  wire \DLX_IDinst_regA_eff[8] ;
  wire CHOICE4217;
  wire DLX_IDinst_RegFile_3_19;
  wire CHOICE2224;
  wire \DLX_IDinst_regA_eff[9] ;
  wire N137086;
  wire CHOICE3193;
  wire DLX_EXinst__n0054;
  wire DLX_EXinst__n0053;
  wire CHOICE5058;
  wire CHOICE4479;
  wire \DLX_EXinst_Mshift__n0021_Sh[41] ;
  wire \DLX_EXinst_Mshift__n0021_Sh[42] ;
  wire CHOICE4534;
  wire CHOICE4474;
  wire DLX_IDinst_RegFile_2_5;
  wire DLX_EXinst_N76011;
  wire CHOICE4490;
  wire N147520;
  wire N138037;
  wire N138143;
  wire CHOICE5713;
  wire CHOICE4493;
  wire CHOICE4924;
  wire CHOICE4419;
  wire DLX_EXinst__n0051;
  wire CHOICE4430;
  wire N138713;
  wire N137774;
  wire CHOICE5458;
  wire CHOICE4433;
  wire DLX_EXinst__n0052;
  wire CHOICE4659;
  wire CHOICE4653;
  wire CHOICE4661;
  wire N163174;
  wire CHOICE4669;
  wire CHOICE4676;
  wire N163473;
  wire CHOICE4699;
  wire CHOICE929;
  wire CHOICE4700;
  wire DLX_IDinst_RegFile_3_1;
  wire N163606;
  wire CHOICE3793;
  wire DLX_EXinst_N74051;
  wire DLX_EXinst__n0080;
  wire CHOICE4688;
  wire \DLX_EXinst_Mshift__n0024_Sh[52] ;
  wire N163485;
  wire CHOICE4647;
  wire CHOICE4634;
  wire CHOICE4663;
  wire DLX_EXinst_N74701;
  wire DLX_EXinst_N74706;
  wire DLX_EXinst_N74971;
  wire CHOICE3692;
  wire CHOICE3802;
  wire DLX_IDinst_RegFile_3_27;
  wire DLX_EXinst_N76318;
  wire DLX_EXinst_N72983;
  wire DLX_EXinst_N74223;
  wire CHOICE3803;
  wire DLX_EXinst__n0079;
  wire DLX_EXinst_N74245;
  wire DLX_EXinst__n0077;
  wire DLX_EXinst__n0078;
  wire N163481;
  wire DLX_EXinst_N74966;
  wire CHOICE4693;
  wire CHOICE4696;
  wire CHOICE3809;
  wire CHOICE3810;
  wire CHOICE4172;
  wire N139405;
  wire N139100;
  wire CHOICE3685;
  wire CHOICE3740;
  wire CHOICE3969;
  wire CHOICE3738;
  wire CHOICE4179;
  wire CHOICE4157;
  wire DLX_IDinst_RegFile_3_10;
  wire N133984;
  wire DLX_EXinst_N74941;
  wire DLX_EXinst_N74711;
  wire CHOICE3859;
  wire CHOICE3747;
  wire CHOICE4721;
  wire CHOICE4729;
  wire CHOICE4730;
  wire N145073;
  wire DLX_EXinst_N76268;
  wire CHOICE4181;
  wire DLX_EXinst_N72993;
  wire N130363;
  wire DLX_EXinst_N72988;
  wire CHOICE3693;
  wire CHOICE3748;
  wire CHOICE3754;
  wire CHOICE3755;
  wire CHOICE4153;
  wire N163639;
  wire CHOICE4184;
  wire CHOICE5400;
  wire CHOICE4107;
  wire DLX_EXinst_N73959;
  wire CHOICE4879;
  wire CHOICE4734;
  wire DLX_IDinst__n0564;
  wire CHOICE3910;
  wire CHOICE3683;
  wire DLX_IDinst_RegFile_7_4;
  wire CHOICE4114;
  wire CHOICE4092;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_259;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_260;
  wire CHOICE4741;
  wire N163672;
  wire CHOICE4760;
  wire CHOICE4754;
  wire CHOICE4762;
  wire CHOICE4763;
  wire DLX_IDinst_RegFile_1_9;
  wire DLX_EXinst_N73794;
  wire DLX_EXinst_N74130;
  wire CHOICE4918;
  wire CHOICE4770;
  wire N145644;
  wire CHOICE4102;
  wire CHOICE4116;
  wire N163321;
  wire CHOICE4764;
  wire CHOICE4766;
  wire CHOICE4731;
  wire CHOICE4771;
  wire CHOICE3699;
  wire CHOICE3700;
  wire \DLX_EXinst_Mshift__n0023_Sh[23] ;
  wire CHOICE5791;
  wire CHOICE5797;
  wire CHOICE5796;
  wire CHOICE4088;
  wire CHOICE4119;
  wire \DLX_EXinst_Mshift__n0019_Sh[11] ;
  wire DLX_EXinst_N73239;
  wire \DLX_EXinst_Mshift__n0023_Sh[22] ;
  wire CHOICE5474;
  wire CHOICE4748;
  wire CHOICE5096;
  wire CHOICE4042;
  wire N163518;
  wire CHOICE4294;
  wire CHOICE4049;
  wire CHOICE4027;
  wire DLX_IDinst_RegFile_15_7;
  wire N126777;
  wire CHOICE5441;
  wire CHOICE4312;
  wire DLX_EXinst_N73287;
  wire CHOICE4914;
  wire \DLX_EXinst_Mshift__n0023_Sh[47] ;
  wire CHOICE5801;
  wire CHOICE5805;
  wire CHOICE5807;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_163;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_164;
  wire CHOICE5829;
  wire N134488;
  wire DLX_EXinst_N74951;
  wire DLX_EXinst_N75139;
  wire CHOICE3977;
  wire CHOICE4301;
  wire CHOICE1661;
  wire N136886;
  wire CHOICE4316;
  wire N145258;
  wire DLX_EXinst_N75983;
  wire CHOICE4051;
  wire DLX_IDinst_RegFile_3_11;
  wire \DLX_EXinst_Mshift__n0019_Sh[127] ;
  wire N164729;
  wire CHOICE4587;
  wire CHOICE4589;
  wire CHOICE4023;
  wire N163390;
  wire CHOICE4054;
  wire \DLX_EXinst_Mshift__n0023_Sh[12] ;
  wire CHOICE3043;
  wire CHOICE5618;
  wire DLX_IDinst_RegFile_22_8;
  wire CHOICE5861;
  wire CHOICE4574;
  wire DLX_EXinst_N76338;
  wire CHOICE4579;
  wire CHOICE4591;
  wire CHOICE4592;
  wire CHOICE4594;
  wire DLX_EXinst_N76473;
  wire CHOICE4624;
  wire \DLX_EXinst_Mshift__n0020_Sh[80] ;
  wire CHOICE4545;
  wire CHOICE4625;
  wire CHOICE5846;
  wire CHOICE5841;
  wire DLX_IDinst_RegFile_23_8;
  wire \DLX_EXinst_Mshift__n0021_Sh[0] ;
  wire \DLX_EXinst_Mshift__n0021_Sh[8] ;
  wire CHOICE4608;
  wire N131375;
  wire CHOICE4609;
  wire CHOICE4614;
  wire CHOICE4626;
  wire \DLX_EXinst_Mshift__n0023_Sh[40] ;
  wire CHOICE5622;
  wire CHOICE5628;
  wire CHOICE5630;
  wire CHOICE4140;
  wire CHOICE5850;
  wire DLX_IDinst_RegFile_7_3;
  wire DLX_EXinst__n0055;
  wire CHOICE5671;
  wire CHOICE5677;
  wire CHOICE5679;
  wire CHOICE4850;
  wire N163631;
  wire CHOICE5383;
  wire CHOICE5385;
  wire CHOICE5639;
  wire DLX_IDinst_RegFile_22_16;
  wire \DLX_EXinst_Mshift__n0020_Sh[28] ;
  wire \DLX_EXinst_Mshift__n0022_Sh[24] ;
  wire \DLX_EXinst_Mshift__n0021_Sh[12] ;
  wire N164155;
  wire CHOICE5668;
  wire CHOICE5634;
  wire N163716;
  wire CHOICE5648;
  wire CHOICE5681;
  wire N163522;
  wire CHOICE5091;
  wire CHOICE5113;
  wire CHOICE5116;
  wire \DLX_EXinst_Mshift__n0023_Sh[41] ;
  wire DLX_EXinst_N75973;
  wire N163514;
  wire DLX_IDinst_RegFile_2_7;
  wire N137608;
  wire N163420;
  wire CHOICE5225;
  wire CHOICE5227;
  wire CHOICE5087;
  wire CHOICE5119;
  wire N163593;
  wire CHOICE5393;
  wire CHOICE5389;
  wire N163584;
  wire CHOICE5427;
  wire CHOICE4962;
  wire CHOICE5242;
  wire N137859;
  wire CHOICE5421;
  wire CHOICE5424;
  wire CHOICE5321;
  wire CHOICE5029;
  wire CHOICE5764;
  wire CHOICE5024;
  wire DLX_IDinst_RegFile_3_4;
  wire CHOICE5046;
  wire CHOICE5049;
  wire \DLX_EXinst_Mshift__n0023_Sh[42] ;
  wire N163660;
  wire CHOICE5304;
  wire CHOICE5305;
  wire CHOICE5020;
  wire CHOICE5052;
  wire N163294;
  wire CHOICE5235;
  wire CHOICE5231;
  wire N163290;
  wire CHOICE5269;
  wire N137372;
  wire N163302;
  wire CHOICE5263;
  wire CHOICE5266;
  wire N163338;
  wire CHOICE5278;
  wire CHOICE5307;
  wire CHOICE5275;
  wire CHOICE5310;
  wire N163684;
  wire DLX_EXinst_N72822;
  wire CHOICE5345;
  wire \DLX_EXinst_Mshift__n0023_Sh[3] ;
  wire N163676;
  wire N163412;
  wire CHOICE4957;
  wire CHOICE4979;
  wire CHOICE4982;
  wire \DLX_EXinst_Mshift__n0023_Sh[43] ;
  wire N163399;
  wire N130467;
  wire CHOICE4896;
  wire CHOICE4908;
  wire CHOICE4902;
  wire CHOICE4910;
  wire CHOICE4911;
  wire CHOICE4953;
  wire CHOICE4985;
  wire CHOICE5314;
  wire CHOICE5348;
  wire CHOICE4792;
  wire CHOICE4800;
  wire CHOICE4801;
  wire CHOICE4912;
  wire CHOICE4876;
  wire CHOICE4919;
  wire DLX_EXinst_N73389;
  wire DLX_EXinst_N73043;
  wire \DLX_EXinst_Mshift__n0019_Sh[12] ;
  wire CHOICE1749;
  wire N163136;
  wire N137448;
  wire CHOICE3939;
  wire CHOICE4805;
  wire DLX_EXinst_N73063;
  wire DLX_EXinst_N73414;
  wire \DLX_EXinst_Mshift__n0019_Sh[21] ;
  wire DLX_IDinst_RegFile_1_17;
  wire CHOICE3711;
  wire CHOICE4812;
  wire \DLX_EXinst_Mshift__n0019_Sh[30] ;
  wire CHOICE1883;
  wire CHOICE4831;
  wire CHOICE4825;
  wire CHOICE4833;
  wire CHOICE4834;
  wire CHOICE4835;
  wire CHOICE4837;
  wire CHOICE4841;
  wire CHOICE4802;
  wire CHOICE4842;
  wire \DLX_EXinst_Mshift__n0019_Sh[10] ;
  wire \DLX_EXinst_Mshift__n0023_Sh[21] ;
  wire CHOICE5550;
  wire CHOICE4819;
  wire DLX_EXinst_N73399;
  wire DLX_EXinst_N73053;
  wire \DLX_EXinst_Mshift__n0019_Sh[8] ;
  wire \DLX_EXinst_Mshift__n0019_Sh[16] ;
  wire DLX_EXinst_N74691;
  wire CHOICE3451;
  wire N163148;
  wire DLX_EXinst_N73404;
  wire \DLX_EXinst_Mshift__n0019_Sh[17] ;
  wire DLX_EXinst_N73058;
  wire \DLX_EXinst_Mshift__n0019_Sh[18] ;
  wire DLX_EXinst_N74731;
  wire DLX_EXinst_N73409;
  wire \DLX_EXinst_Mshift__n0019_Sh[19] ;
  wire \DLX_EXinst_Mshift__n0019_Sh[61] ;
  wire CHOICE1933;
  wire DLX_EXinst_N72803;
  wire \DLX_EXinst_Mshift__n0019_Sh[29] ;
  wire CHOICE2032;
  wire DLX_EXinst_N73369;
  wire DLX_EXinst_N76388;
  wire \DLX_EXinst_Mshift__n0019_Sh[88] ;
  wire CHOICE5146;
  wire DLX_IDinst_RegFile_0_0;
  wire DLX_IDinst_RegFile_0_1;
  wire DLX_IDinst_RegFile_0_2;
  wire red_1_OBUF;
  wire red_0_OBUF;
  wire DLX_IDinst_RegFile_0_4;
  wire DLX_IDinst_RegFile_1_2;
  wire DLX_IDinst_RegFile_1_3;
  wire DLX_IDinst__n0558;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_1;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_3;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_45;
  wire DLX_IDinst_RegFile_4_0;
  wire DLX_IDinst_RegFile_5_0;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_46;
  wire DLX_IDinst_RegFile_6_0;
  wire DLX_IDinst_RegFile_7_0;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_17;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_19;
  wire DLX_IDinst_RegFile_4_1;
  wire DLX_IDinst_RegFile_5_1;
  wire DLX_IDinst_RegFile_6_1;
  wire DLX_IDinst_RegFile_7_1;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_33;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_35;
  wire DLX_IDinst_RegFile_4_2;
  wire DLX_IDinst_RegFile_5_2;
  wire DLX_IDinst_RegFile_6_2;
  wire DLX_IDinst_RegFile_7_2;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_49;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_51;
  wire DLX_IDinst_RegFile_4_3;
  wire DLX_IDinst_RegFile_5_3;
  wire DLX_IDinst_RegFile_6_3;
  wire DLX_IDinst_RegFile_3_7;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_65;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_67;
  wire DLX_IDinst_RegFile_4_4;
  wire DLX_IDinst_RegFile_5_4;
  wire DLX_IDinst_RegFile_6_4;
  wire CHOICE3293;
  wire N163314;
  wire DLX_IDinst__n0102;
  wire DLX_IDinst__n0105;
  wire DLX_IDinst__n0381;
  wire CHOICE3300;
  wire DLX_IDinst_RegFile_3_8;
  wire DLX_IDinst__n0560;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_513;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_515;
  wire DLX_IFinst__n0000;
  wire N128287;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_81;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_83;
  wire DLX_IDinst_RegFile_4_5;
  wire DLX_IDinst_RegFile_5_5;
  wire DLX_IDinst_RegFile_6_5;
  wire DLX_IDinst_RegFile_7_5;
  wire DLX_IDinst_RegFile_3_9;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_529;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_531;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_97;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_99;
  wire DLX_IDinst_RegFile_4_6;
  wire DLX_IDinst_RegFile_5_6;
  wire DLX_IDinst_RegFile_7_6;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_545;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_547;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_113;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_115;
  wire DLX_IDinst_RegFile_4_7;
  wire DLX_IDinst_RegFile_5_7;
  wire DLX_IDinst_RegFile_6_7;
  wire DLX_IDinst_RegFile_7_7;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_561;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_563;
  wire \DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_129;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_131;
  wire DLX_IDinst_RegFile_4_8;
  wire DLX_IDinst_RegFile_5_8;
  wire DLX_IDinst_RegFile_6_8;
  wire DLX_IDinst_RegFile_7_8;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_577;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_579;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_145;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_147;
  wire DLX_IDinst_RegFile_4_9;
  wire DLX_IDinst_RegFile_5_9;
  wire DLX_IDinst_RegFile_6_9;
  wire DLX_IDinst_RegFile_7_9;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_593;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_595;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_609;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_611;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_625;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_627;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_641;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_643;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_657;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_659;
  wire DLX_IDinst__n0566;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_5;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_47;
  wire DLX_IDinst_RegFile_8_0;
  wire DLX_IDinst_RegFile_9_0;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_48;
  wire DLX_IDinst_RegFile_10_0;
  wire DLX_IDinst_RegFile_11_0;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_21;
  wire DLX_IDinst_RegFile_8_1;
  wire DLX_IDinst_RegFile_9_1;
  wire DLX_IDinst_RegFile_10_1;
  wire DLX_IDinst_RegFile_11_1;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_37;
  wire DLX_IDinst_RegFile_8_2;
  wire DLX_IDinst_RegFile_9_2;
  wire DLX_IDinst_RegFile_10_2;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_53;
  wire DLX_IDinst_RegFile_8_3;
  wire DLX_IDinst_RegFile_9_3;
  wire DLX_IDinst_RegFile_10_3;
  wire DLX_IDinst_RegFile_11_3;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_69;
  wire DLX_IDinst_RegFile_8_4;
  wire DLX_IDinst_RegFile_9_4;
  wire DLX_IDinst_RegFile_10_4;
  wire DLX_IDinst_RegFile_11_4;
  wire DLX_IDinst__n0568;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_517;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_85;
  wire DLX_IDinst_RegFile_8_5;
  wire DLX_IDinst_RegFile_9_5;
  wire DLX_IDinst_RegFile_10_5;
  wire DLX_IDinst_RegFile_11_5;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_533;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_101;
  wire DLX_IDinst_RegFile_8_6;
  wire DLX_IDinst_RegFile_9_6;
  wire DLX_IDinst_RegFile_11_6;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_549;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_117;
  wire DLX_IDinst_RegFile_8_7;
  wire DLX_IDinst_RegFile_9_7;
  wire DLX_IDinst_RegFile_10_7;
  wire DLX_IDinst_RegFile_11_7;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_565;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_133;
  wire DLX_IDinst_RegFile_8_8;
  wire DLX_IDinst_RegFile_9_8;
  wire DLX_IDinst_RegFile_10_8;
  wire DLX_IDinst_RegFile_11_8;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_581;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_149;
  wire DLX_IDinst_RegFile_8_9;
  wire DLX_IDinst_RegFile_9_9;
  wire DLX_IDinst_RegFile_10_9;
  wire DLX_IDinst_RegFile_11_9;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_597;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_613;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_629;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_645;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_661;
  wire N129899;
  wire N129847;
  wire N164184;
  wire mask_2_OBUF;
  wire N129795;
  wire N129743;
  wire N129691;
  wire N129639;
  wire N129587;
  wire N129535;
  wire N129483;
  wire N136960;
  wire DLX_IDinst_RegFile_11_10;
  wire DLX_IDinst_RegFile_11_14;
  wire DLX_IDinst_RegFile_11_26;
  wire DLX_IDinst_RegFile_11_28;
  wire DLX_IDinst_RegFile_2_0;
  wire CHOICE3995;
  wire CHOICE5196;
  wire CHOICE4125;
  wire CHOICE4708;
  wire CHOICE4060;
  wire N131631;
  wire CHOICE5881;
  wire N164636;
  wire CHOICE5886;
  wire DLX_IDinst_RegFile_6_23;
  wire CHOICE5585;
  wire DLX_IDinst_RegFile_6_16;
  wire CHOICE3827;
  wire CHOICE3830;
  wire CHOICE3841;
  wire CHOICE3821;
  wire CHOICE3838;
  wire N164583;
  wire N163226;
  wire CHOICE5513;
  wire CHOICE5692;
  wire DLX_IDinst_RegFile_6_19;
  wire CHOICE4779;
  wire CHOICE5354;
  wire CHOICE3133;
  wire CHOICE5890;
  wire CHOICE4992;
  wire CHOICE5017;
  wire CHOICE4991;
  wire CHOICE4539;
  wire CHOICE5696;
  wire \DLX_EXinst_Mshift__n0022_Sh[11] ;
  wire \DLX_EXinst_Mshift__n0022_Sh[9] ;
  wire CHOICE5447;
  wire CHOICE5702;
  wire CHOICE5170;
  wire N131693;
  wire CHOICE5517;
  wire CHOICE5455;
  wire CHOICE5710;
  wire \DLX_EXinst_Mshift__n0021_Sh[22] ;
  wire \DLX_EXinst_Mshift__n0022_Sh[10] ;
  wire CHOICE4716;
  wire CHOICE5523;
  wire N163668;
  wire CHOICE5715;
  wire CHOICE5717;
  wire N163704;
  wire CHOICE5531;
  wire N163931;
  wire CHOICE4328;
  wire CHOICE4329;
  wire CHOICE4330;
  wire CHOICE4332;
  wire CHOICE5186;
  wire CHOICE5534;
  wire CHOICE2058;
  wire CHOICE5526;
  wire CHOICE5536;
  wire CHOICE5538;
  wire DLX_EXinst_N74451;
  wire N133480;
  wire DLX_EXinst_N74696;
  wire CHOICE3718;
  wire CHOICE3945;
  wire N163542;
  wire CHOICE5460;
  wire CHOICE5462;
  wire CHOICE4519;
  wire CHOICE3880;
  wire DLX_EXinst_N72903;
  wire CHOICE3889;
  wire CHOICE3948;
  wire DLX_EXinst_N74686;
  wire N133408;
  wire DLX_EXinst_N74681;
  wire CHOICE4273;
  wire CHOICE3886;
  wire CHOICE5127;
  wire CHOICE3956;
  wire CHOICE5139;
  wire DLX_EXinst_N74446;
  wire DLX_EXinst_N74721;
  wire N133552;
  wire DLX_EXinst_N74991;
  wire CHOICE3773;
  wire CHOICE5724;
  wire CHOICE3897;
  wire DLX_EXinst_N72913;
  wire DLX_EXinst_N76479;
  wire CHOICE5729;
  wire DLX_EXinst_N76457;
  wire CHOICE5732;
  wire CHOICE5132;
  wire CHOICE3656;
  wire CHOICE4263;
  wire CHOICE4505;
  wire CHOICE5477;
  wire CHOICE4510;
  wire vga_top_vga1__n0052;
  wire vga_top_vga1__n0033;
  wire vga_top_vga1__n0034;
  wire vga_top_vga1__n0010;
  wire N138249;
  wire CHOICE4459;
  wire CHOICE4465;
  wire N163728;
  wire CHOICE4467;
  wire DLX_EXinst_N76431;
  wire N164228;
  wire N163979;
  wire CHOICE4405;
  wire N137952;
  wire CHOICE4399;
  wire N163286;
  wire CHOICE4407;
  wire reset_IBUF;
  wire DLX_IDinst__n0617;
  wire \DLX_IDinst_Cause_Reg[0] ;
  wire CHOICE3249;
  wire \DLX_IDinst_Cause_Reg[1] ;
  wire N134590;
  wire N163614;
  wire CHOICE2903;
  wire \DLX_IDinst_Cause_Reg[2] ;
  wire N163720;
  wire CHOICE2888;
  wire \DLX_IDinst_Cause_Reg[3] ;
  wire N163437;
  wire CHOICE2483;
  wire \DLX_IDinst_Cause_Reg[4] ;
  wire N163334;
  wire CHOICE2498;
  wire \DLX_IDinst_Cause_Reg[5] ;
  wire N163365;
  wire CHOICE2513;
  wire \DLX_IDinst_Cause_Reg[7] ;
  wire N163712;
  wire CHOICE2528;
  wire \DLX_IDinst_Cause_Reg[8] ;
  wire N163403;
  wire CHOICE2543;
  wire \DLX_IDinst_Cause_Reg[9] ;
  wire N163570;
  wire CHOICE2558;
  wire CHOICE5181;
  wire N163282;
  wire CHOICE1994;
  wire CHOICE3343;
  wire DLX_IDinst__n0615;
  wire CHOICE3323;
  wire CHOICE3344;
  wire N163460;
  wire DLX_IDinst_N108503;
  wire CHOICE3527;
  wire N163190;
  wire CHOICE3558;
  wire DLX_IDinst__n0163;
  wire N163120;
  wire DLX_IDinst_N107223;
  wire CHOICE3565;
  wire DLX_IDinst_reg_write;
  wire CHOICE4224;
  wire CHOICE4225;
  wire CHOICE4256;
  wire N163546;
  wire N127137;
  wire CHOICE5901;
  wire CHOICE5908;
  wire N164591;
  wire CHOICE5896;
  wire N163416;
  wire CHOICE5945;
  wire N129431;
  wire DLX_IDinst_N108305;
  wire CHOICE2430;
  wire DLX_EXinst_Mcompar__n0065_inst_cy_196;
  wire N164614;
  wire N164612;
  wire DLX_IDinst_N107452;
  wire DLX_IDinst__n0106;
  wire N163258;
  wire DLX_IDinst_CLI;
  wire INT_IBUF;
  wire N163222;
  wire DLX_IDinst_N107623;
  wire CHOICE1689;
  wire N163838;
  wire DLX_IDinst_N108249;
  wire DLX_IDinst__n0391;
  wire DLX_IDinst_N108517;
  wire N129379;
  wire DLX_IDinst_N108552;
  wire CHOICE5747;
  wire \DLX_EXinst_Mshift__n0023_Sh[1] ;
  wire N164200;
  wire CHOICE5749;
  wire CHOICE1319;
  wire CHOICE1320;
  wire DLX_IDinst__n0311;
  wire DLX_IDinst_N108574;
  wire DLX_IDinst_N107870;
  wire DLX_IDinst_N108559;
  wire N128911;
  wire N129327;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_196;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_164;
  wire N164620;
  wire N164618;
  wire N128859;
  wire N129275;
  wire CHOICE2231;
  wire CHOICE2236;
  wire N137082;
  wire CHOICE2242;
  wire CHOICE2247;
  wire CHOICE2423;
  wire CHOICE2357;
  wire DLX_IDinst_RegFile_2_12;
  wire CHOICE2353;
  wire CHOICE2358;
  wire CHOICE2253;
  wire CHOICE2258;
  wire CHOICE2264;
  wire CHOICE2269;
  wire CHOICE2364;
  wire CHOICE2369;
  wire N128391;
  wire N129223;
  wire N128807;
  wire CHOICE2375;
  wire CHOICE2380;
  wire CHOICE2275;
  wire CHOICE2280;
  wire CHOICE2386;
  wire CHOICE2391;
  wire CHOICE2286;
  wire CHOICE2291;
  wire CHOICE2463;
  wire CHOICE2468;
  wire CHOICE3164;
  wire CHOICE2313;
  wire DLX_IDinst_N107609;
  wire CHOICE3173;
  wire CHOICE3178;
  wire CHOICE2213;
  wire CHOICE2456;
  wire CHOICE1926;
  wire N163953;
  wire DLX_IDinst_RegFile_3_29;
  wire CHOICE6016;
  wire DLX_EXinst_N76312;
  wire CHOICE5968;
  wire CHOICE6013;
  wire CHOICE5978;
  wire CHOICE6009;
  wire N163238;
  wire DLX_EXinst_ALU_result_0_1;
  wire CHOICE2309;
  wire CHOICE2314;
  wire CHOICE2452;
  wire CHOICE2457;
  wire CHOICE2441;
  wire CHOICE2446;
  wire CHOICE2320;
  wire CHOICE2325;
  wire N128339;
  wire N129171;
  wire N128703;
  wire CHOICE2435;
  wire CHOICE2331;
  wire CHOICE2336;
  wire CHOICE2342;
  wire CHOICE2347;
  wire CHOICE2419;
  wire CHOICE2424;
  wire CHOICE2412;
  wire CHOICE2408;
  wire CHOICE2413;
  wire CHOICE2397;
  wire CHOICE2402;
  wire N128755;
  wire N129119;
  wire CHOICE5009;
  wire N163250;
  wire CHOICE5014;
  wire DLX_IDinst_RegFile_0_7;
  wire N128651;
  wire N129067;
  wire N128599;
  wire N129015;
  wire DLX_EXinst_N73599;
  wire N130725;
  wire N128547;
  wire N128963;
  wire CHOICE5568;
  wire N164082;
  wire CHOICE5570;
  wire N128495;
  wire N128443;
  wire CHOICE3959;
  wire N164596;
  wire N163182;
  wire CHOICE4266;
  wire CHOICE5492;
  wire N164138;
  wire CHOICE5494;
  wire DLX_IDinst__n0574;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_7;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_49;
  wire DLX_IDinst_RegFile_12_0;
  wire DLX_IDinst_RegFile_13_0;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_50;
  wire DLX_IDinst_RegFile_14_0;
  wire DLX_IDinst_RegFile_15_0;
  wire DLX_IDinst__n0590;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_9;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_11;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_53;
  wire DLX_IDinst_RegFile_20_0;
  wire DLX_IDinst_RegFile_21_0;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_54;
  wire DLX_IDinst_RegFile_22_0;
  wire DLX_IDinst_RegFile_23_0;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_23;
  wire DLX_IDinst_RegFile_12_1;
  wire DLX_IDinst_RegFile_13_1;
  wire DLX_IDinst_RegFile_14_1;
  wire DLX_IDinst_RegFile_15_1;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_25;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_27;
  wire DLX_IDinst_RegFile_20_1;
  wire DLX_IDinst_RegFile_21_1;
  wire DLX_IDinst_RegFile_22_1;
  wire DLX_IDinst_RegFile_23_1;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_39;
  wire DLX_IDinst_RegFile_12_2;
  wire DLX_IDinst_RegFile_13_2;
  wire DLX_IDinst_RegFile_14_2;
  wire DLX_IDinst_RegFile_15_2;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_41;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_43;
  wire DLX_IDinst_RegFile_20_2;
  wire DLX_IDinst_RegFile_21_2;
  wire DLX_IDinst_RegFile_22_2;
  wire DLX_IDinst_RegFile_23_2;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_55;
  wire DLX_IDinst_RegFile_12_3;
  wire DLX_IDinst_RegFile_13_3;
  wire DLX_IDinst_RegFile_14_3;
  wire DLX_IDinst_RegFile_15_3;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_57;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_59;
  wire DLX_IDinst_RegFile_20_3;
  wire DLX_IDinst_RegFile_21_3;
  wire DLX_IDinst_RegFile_22_3;
  wire DLX_IDinst_RegFile_23_3;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_71;
  wire DLX_IDinst_RegFile_12_4;
  wire DLX_IDinst_RegFile_13_4;
  wire DLX_IDinst_RegFile_14_4;
  wire DLX_IDinst_RegFile_15_4;
  wire DLX_IDinst__n0576;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_519;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_73;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_75;
  wire DLX_IDinst_RegFile_20_4;
  wire DLX_IDinst_RegFile_21_4;
  wire DLX_IDinst_RegFile_22_4;
  wire DLX_IDinst_RegFile_23_4;
  wire DLX_IDinst__n0592;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_521;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_523;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_87;
  wire DLX_IDinst_RegFile_12_5;
  wire DLX_IDinst_RegFile_13_5;
  wire DLX_IDinst_RegFile_14_5;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_535;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_89;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_91;
  wire DLX_IDinst_RegFile_20_5;
  wire DLX_IDinst_RegFile_21_5;
  wire DLX_IDinst_RegFile_22_5;
  wire DLX_IDinst_RegFile_23_5;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_537;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_539;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_103;
  wire DLX_IDinst_RegFile_12_6;
  wire DLX_IDinst_RegFile_13_6;
  wire DLX_IDinst_RegFile_14_6;
  wire DLX_IDinst_RegFile_15_6;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_551;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_105;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_107;
  wire DLX_IDinst_RegFile_20_6;
  wire DLX_IDinst_RegFile_21_6;
  wire DLX_IDinst_RegFile_23_6;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_553;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_555;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_119;
  wire DLX_IDinst_RegFile_12_7;
  wire DLX_IDinst_RegFile_13_7;
  wire DLX_IDinst_RegFile_14_7;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_567;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_121;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_123;
  wire DLX_IDinst_RegFile_20_7;
  wire DLX_IDinst_RegFile_21_7;
  wire DLX_IDinst_RegFile_22_7;
  wire DLX_IDinst_RegFile_23_7;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_569;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_571;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_135;
  wire DLX_IDinst_RegFile_12_8;
  wire DLX_IDinst_RegFile_13_8;
  wire DLX_IDinst_RegFile_14_8;
  wire DLX_IDinst_RegFile_15_8;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_583;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_137;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_139;
  wire DLX_IDinst_RegFile_20_8;
  wire DLX_IDinst_RegFile_21_8;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_585;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_587;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_13;
  wire DLX_IDinst_RegFile_28_0;
  wire DLX_IDinst_RegFile_29_0;
  wire DLX_IDinst_RegFile_30_0;
  wire DLX_IDinst_RegFile_31_0;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_151;
  wire DLX_IDinst_RegFile_12_9;
  wire DLX_IDinst_RegFile_13_9;
  wire DLX_IDinst_RegFile_14_9;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_599;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_153;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_155;
  wire DLX_IDinst_RegFile_20_9;
  wire DLX_IDinst_RegFile_21_9;
  wire DLX_IDinst_RegFile_22_9;
  wire DLX_IDinst_RegFile_23_9;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_601;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_603;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_29;
  wire DLX_IDinst_RegFile_28_1;
  wire DLX_IDinst_RegFile_29_1;
  wire DLX_IDinst_RegFile_30_1;
  wire DLX_IDinst_RegFile_31_1;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_615;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_617;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_619;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_45;
  wire DLX_IDinst_RegFile_28_2;
  wire DLX_IDinst_RegFile_29_2;
  wire DLX_IDinst_RegFile_30_2;
  wire DLX_IDinst_RegFile_31_2;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_631;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_633;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_635;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_61;
  wire DLX_IDinst_RegFile_28_3;
  wire DLX_IDinst_RegFile_29_3;
  wire DLX_IDinst_RegFile_30_3;
  wire DLX_IDinst_RegFile_31_3;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_647;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_649;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_651;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_77;
  wire DLX_IDinst_RegFile_28_4;
  wire DLX_IDinst_RegFile_29_4;
  wire DLX_IDinst_RegFile_30_4;
  wire DLX_IDinst_RegFile_31_4;
  wire DLX_IDinst__n0612;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_525;
  wire vga_top_vga1__n0037;
  wire N136748;
  wire vga_top_vga1__n0013;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_663;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_665;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_667;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_93;
  wire DLX_IDinst_RegFile_28_5;
  wire DLX_IDinst_RegFile_29_5;
  wire DLX_IDinst_RegFile_30_5;
  wire DLX_IDinst_RegFile_31_5;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_541;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_109;
  wire DLX_IDinst_RegFile_28_6;
  wire DLX_IDinst_RegFile_29_6;
  wire DLX_IDinst_RegFile_30_6;
  wire DLX_IDinst_RegFile_31_6;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_557;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_125;
  wire DLX_IDinst_RegFile_28_7;
  wire DLX_IDinst_RegFile_30_7;
  wire DLX_IDinst_RegFile_31_7;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_573;
  wire DLX_IDinst_RegFile_16_0;
  wire DLX_IDinst_RegFile_17_0;
  wire DLX_IDinst_RegFile_18_0;
  wire DLX_IDinst_RegFile_19_0;
  wire DLX_IDinst__n0598;
  wire DLX_IDinst_RegFile_24_0;
  wire DLX_IDinst_RegFile_25_0;
  wire DLX_IDinst_RegFile_26_0;
  wire DLX_IDinst_RegFile_27_0;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_141;
  wire DLX_IDinst_RegFile_28_8;
  wire DLX_IDinst_RegFile_29_8;
  wire DLX_IDinst_RegFile_30_8;
  wire DLX_IDinst_RegFile_31_8;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_589;
  wire DLX_IDinst_RegFile_16_1;
  wire DLX_IDinst_RegFile_17_1;
  wire DLX_IDinst_RegFile_19_1;
  wire DLX_IDinst_RegFile_24_1;
  wire DLX_IDinst_RegFile_25_1;
  wire DLX_IDinst_RegFile_26_1;
  wire DLX_IDinst_RegFile_27_1;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_157;
  wire DLX_IDinst_RegFile_28_9;
  wire DLX_IDinst_RegFile_29_9;
  wire DLX_IDinst_RegFile_30_9;
  wire DLX_IDinst_RegFile_31_9;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_605;
  wire DLX_IDinst_RegFile_16_2;
  wire DLX_IDinst_RegFile_17_2;
  wire DLX_IDinst_RegFile_18_2;
  wire DLX_IDinst_RegFile_19_2;
  wire DLX_IDinst_RegFile_24_2;
  wire DLX_IDinst_RegFile_25_2;
  wire DLX_IDinst_RegFile_27_2;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_621;
  wire DLX_IDinst_RegFile_16_3;
  wire DLX_IDinst_RegFile_17_3;
  wire DLX_IDinst_RegFile_18_3;
  wire DLX_IDinst_RegFile_19_3;
  wire DLX_IDinst_RegFile_24_3;
  wire DLX_IDinst_RegFile_25_3;
  wire DLX_IDinst_RegFile_26_3;
  wire DLX_IDinst_RegFile_27_3;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_637;
  wire DLX_IDinst_RegFile_16_4;
  wire DLX_IDinst_RegFile_17_4;
  wire DLX_IDinst_RegFile_19_4;
  wire DLX_IDinst_RegFile_24_4;
  wire DLX_IDinst_RegFile_25_4;
  wire DLX_IDinst_RegFile_26_4;
  wire DLX_IDinst_RegFile_27_4;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_653;
  wire DLX_IDinst_RegFile_16_5;
  wire DLX_IDinst_RegFile_17_5;
  wire DLX_IDinst_RegFile_18_5;
  wire DLX_IDinst_RegFile_19_5;
  wire DLX_IDinst_RegFile_24_5;
  wire DLX_IDinst_RegFile_25_5;
  wire DLX_IDinst_RegFile_27_5;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_669;
  wire CHOICE3139;
  wire DLX_IDinst_RegFile_16_6;
  wire DLX_IDinst_RegFile_17_6;
  wire DLX_IDinst_RegFile_18_6;
  wire DLX_IDinst_RegFile_19_6;
  wire DLX_IDinst_RegFile_24_6;
  wire DLX_IDinst_RegFile_25_6;
  wire DLX_IDinst_RegFile_26_6;
  wire DLX_IDinst_RegFile_27_6;
  wire DLX_IDinst_RegFile_16_7;
  wire DLX_IDinst_RegFile_17_7;
  wire DLX_IDinst_RegFile_18_7;
  wire DLX_IDinst_RegFile_19_7;
  wire DLX_IDinst_RegFile_24_7;
  wire DLX_IDinst_RegFile_25_7;
  wire DLX_IDinst_RegFile_26_7;
  wire DLX_IDinst_RegFile_27_7;
  wire CHOICE3455;
  wire DLX_IDinst_RegFile_16_8;
  wire DLX_IDinst_RegFile_17_8;
  wire DLX_IDinst_RegFile_18_8;
  wire DLX_IDinst_RegFile_19_8;
  wire DLX_IDinst_RegFile_24_8;
  wire DLX_IDinst_RegFile_25_8;
  wire DLX_IDinst_RegFile_26_8;
  wire DLX_IDinst_RegFile_27_8;
  wire CHOICE3251;
  wire CHOICE3232;
  wire DLX_IDinst_RegFile_16_9;
  wire DLX_IDinst_RegFile_17_9;
  wire DLX_IDinst_RegFile_18_9;
  wire DLX_IDinst_RegFile_19_9;
  wire DLX_IDinst_RegFile_24_9;
  wire DLX_IDinst_RegFile_25_9;
  wire DLX_IDinst_RegFile_26_9;
  wire DLX_IDinst_RegFile_27_9;
  wire vga_top_vga1_clockcounter_FFd1;
  wire CHOICE3458;
  wire CHOICE3459;
  wire CHOICE1944;
  wire CHOICE4342;
  wire DLX_EXinst_N72898;
  wire N163432;
  wire CHOICE4347;
  wire CHOICE6002;
  wire CHOICE4942;
  wire \DLX_EXinst_Mshift__n0022_Sh[59] ;
  wire N163530;
  wire DLX_IDinst_RegFile_2_14;
  wire DLX_EXinst_N76002;
  wire CHOICE4037;
  wire CHOICE5779;
  wire CHOICE4886;
  wire CHOICE4341;
  wire DLX_IDinst_RegFile_0_21;
  wire DLX_IDinst_RegFile_0_11;
  wire DLX_IDinst_RegFile_0_13;
  wire DLX_IDinst_RegFile_0_30;
  wire DLX_IDinst_RegFile_0_22;
  wire DLX_IDinst_RegFile_0_14;
  wire DLX_IDinst_RegFile_0_31;
  wire DLX_IDinst_RegFile_0_23;
  wire DLX_IDinst_RegFile_0_15;
  wire DLX_IDinst_RegFile_0_24;
  wire DLX_IDinst_RegFile_0_16;
  wire DLX_IDinst_RegFile_0_25;
  wire DLX_IDinst_RegFile_0_17;
  wire DLX_IDinst_RegFile_1_10;
  wire DLX_IDinst_RegFile_0_26;
  wire DLX_IDinst_RegFile_0_18;
  wire DLX_IDinst_RegFile_1_11;
  wire DLX_IDinst_RegFile_0_27;
  wire DLX_IDinst_RegFile_0_19;
  wire DLX_IDinst_RegFile_1_12;
  wire DLX_IDinst_RegFile_0_28;
  wire DLX_IDinst_RegFile_1_20;
  wire DLX_IDinst_RegFile_1_13;
  wire DLX_IDinst_RegFile_0_29;
  wire DLX_IDinst_RegFile_1_21;
  wire DLX_IDinst_RegFile_1_14;
  wire DLX_IDinst_RegFile_1_30;
  wire DLX_IDinst_RegFile_1_22;
  wire DLX_IDinst_RegFile_1_31;
  wire DLX_IDinst_RegFile_1_15;
  wire DLX_IDinst_RegFile_1_16;
  wire DLX_IDinst_RegFile_1_25;
  wire DLX_IDinst_RegFile_2_10;
  wire DLX_IDinst_RegFile_1_18;
  wire DLX_IDinst_RegFile_1_27;
  wire DLX_IDinst_RegFile_2_11;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_161;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_163;
  wire DLX_IDinst_RegFile_4_10;
  wire DLX_IDinst_RegFile_5_10;
  wire DLX_IDinst_RegFile_6_10;
  wire DLX_IDinst_RegFile_7_10;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_177;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_179;
  wire DLX_IDinst_RegFile_4_11;
  wire DLX_IDinst_RegFile_5_11;
  wire DLX_IDinst_RegFile_6_11;
  wire DLX_IDinst_RegFile_7_11;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_193;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_195;
  wire DLX_IDinst_RegFile_4_12;
  wire DLX_IDinst_RegFile_5_12;
  wire DLX_IDinst_RegFile_6_12;
  wire DLX_IDinst_RegFile_7_12;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_321;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_323;
  wire DLX_IDinst_RegFile_4_20;
  wire DLX_IDinst_RegFile_5_20;
  wire DLX_IDinst_RegFile_6_20;
  wire DLX_IDinst_RegFile_7_20;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_209;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_211;
  wire DLX_IDinst_RegFile_4_13;
  wire DLX_IDinst_RegFile_5_13;
  wire DLX_IDinst_RegFile_6_13;
  wire DLX_IDinst_RegFile_7_13;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_337;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_339;
  wire DLX_IDinst_RegFile_4_21;
  wire DLX_IDinst_RegFile_5_21;
  wire DLX_IDinst_RegFile_6_21;
  wire DLX_IDinst_RegFile_7_21;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_225;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_227;
  wire DLX_IDinst_RegFile_4_14;
  wire DLX_IDinst_RegFile_5_14;
  wire DLX_IDinst_RegFile_6_14;
  wire DLX_IDinst_RegFile_7_14;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_353;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_355;
  wire DLX_IDinst_RegFile_4_22;
  wire DLX_IDinst_RegFile_5_22;
  wire DLX_IDinst_RegFile_6_22;
  wire DLX_IDinst_RegFile_7_22;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_993;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_995;
  wire DLX_IDinst_RegFile_4_30;
  wire DLX_IDinst_RegFile_5_30;
  wire DLX_IDinst_RegFile_6_30;
  wire DLX_IDinst_RegFile_7_30;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_1009;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_1011;
  wire DLX_IDinst_RegFile_4_31;
  wire DLX_IDinst_RegFile_5_31;
  wire DLX_IDinst_RegFile_6_31;
  wire DLX_IDinst_RegFile_7_31;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_241;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_243;
  wire DLX_IDinst_RegFile_4_15;
  wire DLX_IDinst_RegFile_5_15;
  wire DLX_IDinst_RegFile_6_15;
  wire DLX_IDinst_RegFile_7_15;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_369;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_371;
  wire DLX_IDinst_RegFile_4_23;
  wire DLX_IDinst_RegFile_5_23;
  wire DLX_IDinst_RegFile_7_23;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_257;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_259;
  wire DLX_IDinst_RegFile_4_16;
  wire DLX_IDinst_RegFile_5_16;
  wire DLX_IDinst_RegFile_7_16;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_385;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_387;
  wire DLX_IDinst_RegFile_4_24;
  wire DLX_IDinst_RegFile_5_24;
  wire DLX_IDinst_RegFile_6_24;
  wire DLX_IDinst_RegFile_7_24;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_273;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_275;
  wire DLX_IDinst_RegFile_4_17;
  wire DLX_IDinst_RegFile_5_17;
  wire DLX_IDinst_RegFile_6_17;
  wire DLX_IDinst_RegFile_7_17;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_401;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_403;
  wire DLX_IDinst_RegFile_4_25;
  wire DLX_IDinst_RegFile_5_25;
  wire DLX_IDinst_RegFile_6_25;
  wire DLX_IDinst_RegFile_7_25;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_289;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_291;
  wire DLX_IDinst_RegFile_4_18;
  wire DLX_IDinst_RegFile_5_18;
  wire DLX_IDinst_RegFile_6_18;
  wire DLX_IDinst_RegFile_7_18;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_417;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_419;
  wire DLX_IDinst_RegFile_4_26;
  wire DLX_IDinst_RegFile_5_26;
  wire DLX_IDinst_RegFile_6_26;
  wire DLX_IDinst_RegFile_7_26;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_673;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_675;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_305;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_307;
  wire DLX_IDinst_RegFile_4_19;
  wire DLX_IDinst_RegFile_5_19;
  wire DLX_IDinst_RegFile_7_19;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_433;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_435;
  wire DLX_IDinst_RegFile_4_27;
  wire DLX_IDinst_RegFile_5_27;
  wire DLX_IDinst_RegFile_6_27;
  wire DLX_IDinst_RegFile_7_27;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_689;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_691;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_961;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_963;
  wire DLX_IDinst_RegFile_4_28;
  wire DLX_IDinst_RegFile_5_28;
  wire DLX_IDinst_RegFile_6_28;
  wire DLX_IDinst_RegFile_7_28;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_833;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_835;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_705;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_707;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_977;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_979;
  wire DLX_IDinst_RegFile_4_29;
  wire DLX_IDinst_RegFile_5_29;
  wire DLX_IDinst_RegFile_6_29;
  wire DLX_IDinst_RegFile_7_29;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_849;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_851;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_721;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_723;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_481;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_483;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_865;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_867;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_737;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_739;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_497;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_499;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_881;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_883;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_753;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_755;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_897;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_899;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_769;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_771;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_913;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_915;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_785;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_787;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_929;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_931;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_801;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_803;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_945;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_947;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_817;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_819;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_449;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_451;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_165;
  wire DLX_IDinst_RegFile_8_10;
  wire DLX_IDinst_RegFile_9_10;
  wire DLX_IDinst_RegFile_10_10;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_181;
  wire DLX_IDinst_RegFile_8_11;
  wire DLX_IDinst_RegFile_9_11;
  wire DLX_IDinst_RegFile_10_11;
  wire DLX_IDinst_RegFile_11_11;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_325;
  wire DLX_IDinst_RegFile_8_20;
  wire DLX_IDinst_RegFile_9_20;
  wire DLX_IDinst_RegFile_10_20;
  wire DLX_IDinst_RegFile_11_20;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_197;
  wire DLX_IDinst_RegFile_8_12;
  wire DLX_IDinst_RegFile_9_12;
  wire DLX_IDinst_RegFile_10_12;
  wire DLX_IDinst_RegFile_11_12;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_341;
  wire DLX_IDinst_RegFile_8_21;
  wire DLX_IDinst_RegFile_9_21;
  wire DLX_IDinst_RegFile_10_21;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_213;
  wire DLX_IDinst_RegFile_8_13;
  wire DLX_IDinst_RegFile_9_13;
  wire DLX_IDinst_RegFile_10_13;
  wire DLX_IDinst_RegFile_11_13;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_997;
  wire DLX_IDinst_RegFile_8_30;
  wire DLX_IDinst_RegFile_9_30;
  wire DLX_IDinst_RegFile_10_30;
  wire DLX_IDinst_RegFile_11_30;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_357;
  wire DLX_IDinst_RegFile_8_22;
  wire DLX_IDinst_RegFile_9_22;
  wire DLX_IDinst_RegFile_10_22;
  wire DLX_IDinst_RegFile_11_22;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_229;
  wire DLX_IDinst_RegFile_8_14;
  wire DLX_IDinst_RegFile_9_14;
  wire DLX_IDinst_RegFile_10_14;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_373;
  wire DLX_IDinst_RegFile_8_23;
  wire DLX_IDinst_RegFile_9_23;
  wire DLX_IDinst_RegFile_10_23;
  wire DLX_IDinst_RegFile_11_23;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_245;
  wire DLX_IDinst_RegFile_8_15;
  wire DLX_IDinst_RegFile_9_15;
  wire DLX_IDinst_RegFile_10_15;
  wire DLX_IDinst_RegFile_11_15;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_1013;
  wire DLX_IDinst_RegFile_8_31;
  wire DLX_IDinst_RegFile_9_31;
  wire DLX_IDinst_RegFile_10_31;
  wire DLX_IDinst_RegFile_11_31;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_389;
  wire DLX_IDinst_RegFile_8_24;
  wire DLX_IDinst_RegFile_9_24;
  wire DLX_IDinst_RegFile_10_24;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_261;
  wire DLX_IDinst_RegFile_8_16;
  wire DLX_IDinst_RegFile_9_16;
  wire DLX_IDinst_RegFile_10_16;
  wire DLX_IDinst_RegFile_11_16;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_405;
  wire DLX_IDinst_RegFile_8_25;
  wire DLX_IDinst_RegFile_9_25;
  wire DLX_IDinst_RegFile_10_25;
  wire DLX_IDinst_RegFile_11_25;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_277;
  wire DLX_IDinst_RegFile_8_17;
  wire DLX_IDinst_RegFile_9_17;
  wire DLX_IDinst_RegFile_10_17;
  wire DLX_IDinst_RegFile_11_17;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_421;
  wire DLX_IDinst_RegFile_8_26;
  wire DLX_IDinst_RegFile_9_26;
  wire DLX_IDinst_RegFile_10_26;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_293;
  wire DLX_IDinst_RegFile_8_18;
  wire DLX_IDinst_RegFile_9_18;
  wire DLX_IDinst_RegFile_10_18;
  wire DLX_IDinst_RegFile_11_18;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_677;
  wire \DLX_EXinst_Mshift__n0022_Sh[52] ;
  wire CHOICE4371;
  wire N163827;
  wire CHOICE4373;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_437;
  wire DLX_IDinst_RegFile_8_27;
  wire DLX_IDinst_RegFile_9_27;
  wire DLX_IDinst_RegFile_10_27;
  wire DLX_IDinst_RegFile_11_27;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_309;
  wire DLX_IDinst_RegFile_8_19;
  wire DLX_IDinst_RegFile_9_19;
  wire DLX_IDinst_RegFile_10_19;
  wire DLX_IDinst_RegFile_11_19;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_693;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_965;
  wire DLX_IDinst_RegFile_8_28;
  wire DLX_IDinst_RegFile_9_28;
  wire DLX_IDinst_RegFile_10_28;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_837;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_709;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_981;
  wire DLX_IDinst_RegFile_8_29;
  wire DLX_IDinst_RegFile_9_29;
  wire DLX_IDinst_RegFile_10_29;
  wire DLX_IDinst_RegFile_11_29;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_853;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_725;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_485;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_869;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_885;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_757;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_501;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_901;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_773;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_917;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_789;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_933;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_805;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_949;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_821;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_453;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_467;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_469;
  wire N136625;
  wire vga_top_vga1_N112926;
  wire DLX_IDinst__n0161;
  wire CHOICE246;
  wire DLX_IDinst_RegFile_3_28;
  wire CHOICE254;
  wire N163210;
  wire \DLX_EXinst_Mshift__n0021_Sh[9] ;
  wire \DLX_EXinst_Mshift__n0021_Sh[5] ;
  wire N131439;
  wire N130261;
  wire DLX_EXinst_N73998;
  wire N131503;
  wire DLX_IDinst_RegFile_0_10;
  wire N164562;
  wire DLX_IDinst_RegFile_2_1;
  wire N130209;
  wire \DLX_EXinst_Mshift__n0021_Sh[13] ;
  wire DLX_EXinst_N73993;
  wire DLX_IDinst_RegFile_0_20;
  wire CHOICE3468;
  wire N163708;
  wire N147636;
  wire CHOICE3113;
  wire CHOICE3130;
  wire N163618;
  wire CHOICE3900;
  wire CHOICE3036;
  wire \DLX_EXinst_Mshift__n0019_Sh[23] ;
  wire CHOICE3052;
  wire CHOICE3072;
  wire DLX_IDinst_RegFile_2_2;
  wire CHOICE3065;
  wire CHOICE2945;
  wire CHOICE2938;
  wire N144481;
  wire CHOICE4084;
  wire CHOICE3646;
  wire DLX_IDinst_RegFile_2_3;
  wire CHOICE2972;
  wire CHOICE2965;
  wire N144646;
  wire CHOICE4149;
  wire CHOICE3449;
  wire \DLX_EXinst_Mshift__n0020_Sh[27] ;
  wire CHOICE2953;
  wire CHOICE3101;
  wire DLX_IDinst_RegFile_2_4;
  wire CHOICE3094;
  wire N145443;
  wire CHOICE4019;
  wire N162801;
  wire N162807;
  wire CHOICE3321;
  wire N136696;
  wire DLX_IDinst__n0104;
  wire DLX_IDinst_RegFile_15_31;
  wire DLX_IDinst__n0367;
  wire DLX_IDinst_RegFile_15_18;
  wire DLX_IDinst__n0368;
  wire CHOICE2118;
  wire DLX_IDinst_RegFile_15_19;
  wire DLX_IDinst_N108531;
  wire DLX_IDinst__n0097;
  wire CHOICE2103;
  wire N139563;
  wire DLX_IDinst_N108254;
  wire N135272;
  wire IR_MSB_6_OBUF;
  wire DLX_IDinst_N108545;
  wire DLX_IDinst_N108510;
  wire DLX_IDinst_N108524;
  wire DLX_IDinst_RegFile_0_3;
  wire N162863;
  wire CHOICE3396;
  wire DLX_IDinst__n0635;
  wire DLX_IDinst_RegFile_0_5;
  wire IR_MSB_2_OBUF;
  wire CHOICE4445;
  wire CHOICE4390;
  wire CHOICE4450;
  wire CHOICE4385;
  wire CHOICE3782;
  wire CHOICE3766;
  wire DLX_EXinst_N75154;
  wire N163526;
  wire CHOICE4642;
  wire CHOICE3774;
  wire CHOICE3784;
  wire CHOICE3785;
  wire N130157;
  wire N130051;
  wire CHOICE4274;
  wire CHOICE3719;
  wire CHOICE5154;
  wire N163538;
  wire CHOICE5156;
  wire CHOICE3727;
  wire DLX_IDinst_RegFile_1_24;
  wire CHOICE3729;
  wire CHOICE3730;
  wire \DLX_EXinst_Mshift__n0023_Sh[5] ;
  wire CHOICE3663;
  wire N130001;
  wire \DLX_EXinst_Mshift__n0023_Sh[10] ;
  wire N130105;
  wire DLX_EXinst_N73853;
  wire CHOICE3664;
  wire CHOICE4929;
  wire CHOICE4075;
  wire DLX_IDinst_RegFile_3_2;
  wire CHOICE5469;
  wire CHOICE3672;
  wire DLX_IDinst_RegFile_3_3;
  wire CHOICE3674;
  wire CHOICE3675;
  wire CHOICE5063;
  wire CHOICE4010;
  wire CHOICE5545;
  wire CHOICE2049;
  wire CHOICE5909;
  wire DLX_IDinst_RegFile_2_8;
  wire \DLX_EXinst_Mshift__n0023_Sh[0] ;
  wire CHOICE5915;
  wire CHOICE4282;
  wire CHOICE4284;
  wire CHOICE4285;
  wire CHOICE4287;
  wire CHOICE1830;
  wire CHOICE5598;
  wire CHOICE5939;
  wire CHOICE5941;
  wire DLX_IDinst_RegFile_3_5;
  wire CHOICE5203;
  wire CHOICE5361;
  wire CHOICE5741;
  wire N163648;
  wire DLX_EXinst_mem_to_reg_EX;
  wire CHOICE5603;
  wire CHOICE5952;
  wire CHOICE5967;
  wire CHOICE5608;
  wire CHOICE5631;
  wire DLX_IDinst_RegFile_2_9;
  wire CHOICE5976;
  wire N138481;
  wire CHOICE5081;
  wire CHOICE5083;
  wire CHOICE5929;
  wire CHOICE5923;
  wire CHOICE5938;
  wire \DLX_EXinst_Mshift__n0019_Sh[9] ;
  wire CHOICE5999;
  wire CHOICE6008;
  wire CHOICE5751;
  wire N164573;
  wire CHOICE5993;
  wire CHOICE5994;
  wire DLX_EXinst_N74625;
  wire CHOICE5503;
  wire CHOICE5758;
  wire CHOICE3912;
  wire CHOICE5015;
  wire N163242;
  wire CHOICE5562;
  wire N163394;
  wire CHOICE4947;
  wire CHOICE4949;
  wire CHOICE5553;
  wire CHOICE5572;
  wire N164587;
  wire \DLX_EXinst_Mshift__n0021_Sh[21] ;
  wire CHOICE4787;
  wire CHOICE4861;
  wire CHOICE5486;
  wire N163493;
  wire CHOICE5496;
  wire N164601;
  wire CHOICE4362;
  wire CHOICE4375;
  wire CHOICE4377;
  wire CHOICE4360;
  wire CHOICE4361;
  wire N162850;
  wire CHOICE4378;
  wire DLX_EXinst_ALU_result_4_1;
  wire CHOICE1859;
  wire CHOICE3971;
  wire CHOICE3921;
  wire CHOICE3980;
  wire CHOICE3986;
  wire CHOICE3987;
  wire N134056;
  wire DLX_EXinst_N74936;
  wire CHOICE3918;
  wire DLX_IDinst_RegFile_14_31;
  wire CHOICE3927;
  wire CHOICE3928;
  wire CHOICE3851;
  wire CHOICE3853;
  wire DLX_EXinst_N72998;
  wire DLX_EXinst_N73018;
  wire CHOICE3862;
  wire CHOICE3377;
  wire DLX_IDinst_RegFile_22_17;
  wire CHOICE3868;
  wire CHOICE3869;
  wire \DLX_EXinst_Mshift__n0021_Sh[40] ;
  wire CHOICE5165;
  wire CHOICE4552;
  wire CHOICE4553;
  wire DLX_IDinst_RegFile_14_18;
  wire CHOICE4554;
  wire CHOICE4555;
  wire N163489;
  wire CHOICE5188;
  wire N164119;
  wire DLX_IDinst_RegFile_23_10;
  wire DLX_IDinst_RegFile_14_27;
  wire DLX_IDinst_RegFile_22_19;
  wire N163156;
  wire N163158;
  wire N144912;
  wire CHOICE1669;
  wire DLX_IDinst_RegFile_15_17;
  wire N163688;
  wire CHOICE4495;
  wire DLX_IFinst_stalled;
  wire DLX_IDinst__n0313;
  wire N127012;
  wire N130977;
  wire N163230;
  wire CHOICE4435;
  wire \DLX_EXinst_Mshift__n0022_Sh[19] ;
  wire N163664;
  wire CHOICE2723;
  wire vga_top_vga1_N112921;
  wire N132456;
  wire vga_top_vga1__n0014;
  wire DLX_IDinst_RegFile_23_27;
  wire CHOICE2112;
  wire \DLX_EXinst_Mshift__n0021_Sh[4] ;
  wire \DLX_EXinst_Mshift__n0021_Sh[6] ;
  wire N163442;
  wire CHOICE2738;
  wire DLX_EXinst_N73509;
  wire DLX_EXinst_N72933;
  wire DLX_IDinst_Mmux__n0162__net105;
  wire CHOICE2188;
  wire CHOICE2177;
  wire CHOICE3171;
  wire CHOICE3156;
  wire CHOICE2166;
  wire CHOICE2220;
  wire CHOICE2155;
  wire CHOICE4135;
  wire N163680;
  wire N163700;
  wire CHOICE2753;
  wire N163325;
  wire CHOICE4573;
  wire CHOICE3146;
  wire CHOICE3149;
  wire N163510;
  wire CHOICE2768;
  wire DLX_EXinst_N72848;
  wire \DLX_EXinst_Mshift__n0023_Sh[7] ;
  wire DLX_EXinst_N73604;
  wire \DLX_EXinst_Mshift__n0023_Sh[8] ;
  wire DLX_EXinst_N73023;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_261;
  wire DLX_EXinst__n0087;
  wire CHOICE4167;
  wire CHOICE3165;
  wire CHOICE2144;
  wire CHOICE2149;
  wire CHOICE2160;
  wire CHOICE4070;
  wire N163278;
  wire CHOICE5258;
  wire \DLX_EXinst_Mshift__n0024_Sh[50] ;
  wire CHOICE2171;
  wire CHOICE2182;
  wire N163447;
  wire CHOICE2663;
  wire N163262;
  wire CHOICE2783;
  wire CHOICE2193;
  wire CHOICE3185;
  wire CHOICE3194;
  wire CHOICE2200;
  wire CHOICE2203;
  wire CHOICE2209;
  wire CHOICE2214;
  wire CHOICE2225;
  wire N163622;
  wire CHOICE2798;
  wire N163588;
  wire CHOICE2678;
  wire DLX_IDinst__n0549;
  wire CHOICE2918;
  wire CHOICE2919;
  wire CHOICE4005;
  wire N163456;
  wire CHOICE4302;
  wire N163477;
  wire CHOICE4314;
  wire N163465;
  wire CHOICE2813;
  wire N163452;
  wire CHOICE2708;
  wire N131077;
  wire \DLX_IDinst_Cause_Reg[10] ;
  wire N163578;
  wire CHOICE2573;
  wire \DLX_IDinst_Cause_Reg[11] ;
  wire N163234;
  wire CHOICE2588;
  wire \DLX_IDinst_Cause_Reg[12] ;
  wire N163361;
  wire CHOICE2603;
  wire \DLX_IDinst_Cause_Reg[13] ;
  wire N163566;
  wire CHOICE2618;
  wire \DLX_IDinst_Cause_Reg[14] ;
  wire N163382;
  wire CHOICE2633;
  wire \DLX_IDinst_Cause_Reg[15] ;
  wire N163329;
  wire CHOICE2648;
  wire N163254;
  wire CHOICE2828;
  wire DLX_EXinst_N73068;
  wire N163737;
  wire CHOICE2693;
  wire N163550;
  wire CHOICE5811;
  wire N163178;
  wire CHOICE3062;
  wire N163643;
  wire CHOICE2843;
  wire \DLX_EXinst_Mshift__n0022_Sh[21] ;
  wire \DLX_EXinst_Mshift__n0021_Sh[23] ;
  wire DLX_EXinst_N73013;
  wire N163186;
  wire DLX_EXinst_N73424;
  wire CHOICE1899;
  wire CHOICE1907;
  wire CHOICE1921;
  wire CHOICE1955;
  wire CHOICE1963;
  wire CHOICE3121;
  wire CHOICE3122;
  wire CHOICE3026;
  wire DLX_IDinst_Mcompar__n0368_inst_cy_263;
  wire CHOICE1870;
  wire CHOICE2053;
  wire CHOICE2035;
  wire DLX_EXinst_N72809;
  wire N164172;
  wire \DLX_EXinst_Mshift__n0019_Sh[28] ;
  wire CHOICE1280;
  wire N139189;
  wire CHOICE1670;
  wire CHOICE2926;
  wire DLX_EXinst_N72746;
  wire CHOICE3608;
  wire CHOICE3615;
  wire CHOICE1276;
  wire N134683;
  wire DLX_IDinst_mem_write;
  wire DLX_EXinst_mem_write_EX;
  wire N139297;
  wire CHOICE3081;
  wire N163140;
  wire CHOICE3091;
  wire CHOICE1291;
  wire CHOICE1295;
  wire CHOICE3795;
  wire CHOICE2020;
  wire CHOICE2071;
  wire DLX_EXinst_N73549;
  wire CHOICE2067;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_43;
  wire CHOICE2025;
  wire CHOICE2076;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_44;
  wire CHOICE1877;
  wire N163506;
  wire CHOICE2858;
  wire CHOICE1888;
  wire CHOICE1939;
  wire N138591;
  wire CHOICE5838;
  wire CHOICE5864;
  wire N163497;
  wire N163246;
  wire N163124;
  wire N126925;
  wire CHOICE1327;
  wire CHOICE1348;
  wire blue_1_OBUF;
  wire green_1_OBUF;
  wire CHOICE5108;
  wire N163534;
  wire DLX_EXinst_N75993;
  wire N163602;
  wire N163627;
  wire CHOICE5041;
  wire N163692;
  wire CHOICE2198;
  wire N162854;
  wire DLX_EXinst_N74136;
  wire N163270;
  wire DLX_EXinst_ALU_result_1_1;
  wire vga_top_vga1_N112931;
  wire N163407;
  wire CHOICE4974;
  wire N163428;
  wire N164207;
  wire CHOICE4525;
  wire N163656;
  wire CHOICE4527;
  wire \DLX_EXinst_Mshift__n0021_Sh[43] ;
  wire N163501;
  wire DLX_EXinst_N73113;
  wire DLX_EXinst_N73429;
  wire DLX_EXinst_N73033;
  wire DLX_EXinst_N73514;
  wire DLX_EXinst_N73123;
  wire DLX_EXinst_N74003;
  wire DLX_EXinst_N73108;
  wire DLX_EXinst_N73028;
  wire DLX_EXinst_N73524;
  wire DLX_EXinst_N73133;
  wire N130825;
  wire DLX_EXinst_N73554;
  wire DLX_EXinst_N73118;
  wire DLX_EXinst_N73384;
  wire DLX_EXinst_N73038;
  wire \DLX_EXinst_Mshift__n0019_Sh[20] ;
  wire DLX_EXinst_N73394;
  wire DLX_EXinst_N73048;
  wire \DLX_EXinst_Mshift__n0023_Sh[13] ;
  wire N133048;
  wire DLX_EXinst_N74024;
  wire DLX_EXinst_N72978;
  wire \DLX_EXinst_Mshift__n0023_Sh[15] ;
  wire DLX_EXinst_N74034;
  wire N130519;
  wire DLX_EXinst_N73083;
  wire DLX_EXinst_N73539;
  wire DLX_EXinst_N73148;
  wire \DLX_EXinst_Mshift__n0022_Sh[20] ;
  wire \DLX_EXinst_Mshift__n0023_Sh[14] ;
  wire N133120;
  wire DLX_EXinst_N74029;
  wire DLX_EXinst_N74206;
  wire CHOICE4866;
  wire CHOICE4874;
  wire N164579;
  wire DLX_EXinst_N73088;
  wire DLX_EXinst_N73354;
  wire DLX_EXinst_N72853;
  wire \DLX_EXinst_Mshift__n0023_Sh[9] ;
  wire N130773;
  wire DLX_EXinst_N73374;
  wire \DLX_EXinst_Mshift__n0019_Sh[24] ;
  wire N130875;
  wire DLX_EXinst_N73474;
  wire DLX_EXinst_N76047;
  wire DLX_EXinst_N72863;
  wire DLX_EXinst_N73564;
  wire N133768;
  wire DLX_EXinst_N74196;
  wire DLX_EXinst_N73559;
  wire DLX_EXinst_N72948;
  wire DLX_EXinst_N73469;
  wire DLX_EXinst_N73494;
  wire DLX_EXinst_N72873;
  wire N129951;
  wire N130621;
  wire DLX_EXinst_N73569;
  wire DLX_EXinst_N72958;
  wire DLX_EXinst_N72858;
  wire \DLX_EXinst_Mshift__n0023_Sh[11] ;
  wire DLX_EXinst_N72883;
  wire DLX_EXinst_N73584;
  wire DLX_EXinst_N72968;
  wire DLX_EXinst_N73489;
  wire N134128;
  wire DLX_EXinst_N74201;
  wire DLX_EXinst_N73589;
  wire DLX_EXinst_N72893;
  wire DLX_EXinst_N72797;
  wire \DLX_EXinst_Mshift__n0023_Sh[4] ;
  wire DLX_EXinst_N73848;
  wire DLX_EXinst_N73858;
  wire N162810;
  wire CHOICE4558;
  wire DLX_EXinst_ALU_result_9_1;
  wire CHOICE4414;
  wire DLX_EXinst_N76496;
  wire N131996;
  wire N164607;
  wire N163198;
  wire CHOICE3211;
  wire CHOICE3213;
  wire CHOICE3373;
  wire CHOICE3386;
  wire CHOICE3301;
  wire DLX_EXinst_Mcompar__n0069_inst_cy_260;
  wire DLX_EXinst_Mcompar__n0069_inst_cy_261;
  wire DLX_EXinst__n0061;
  wire CHOICE1326;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_228;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_229;
  wire DLX_EXinst__n0085;
  wire CHOICE1693;
  wire N162841;
  wire CHOICE5579;
  wire N163266;
  wire DLX_EXinst_ALU_result_2_1;
  wire N132148;
  wire N132422;
  wire N136962;
  wire DLX_IDinst_mem_to_reg;
  wire N164089;
  wire DLX_EXinst_N72765;
  wire N132193;
  wire DLX_IDinst__n0616;
  wire DLX_IDinst_RegFile_0_8;
  wire N164094;
  wire DLX_IDinst_RegFile_0_9;
  wire N132252;
  wire N162860;
  wire N163274;
  wire DLX_EXinst_ALU_result_3_1;
  wire N131191;
  wire N131255;
  wire N131315;
  wire \DLX_EXinst_Mshift__n0021_Sh[7] ;
  wire CHOICE1354;
  wire CHOICE1355;
  wire CHOICE1361;
  wire CHOICE1362;
  wire CHOICE1373;
  wire CHOICE1381;
  wire CHOICE1383;
  wire DLX_IDinst__n0153;
  wire \clk/new_buffer ;
  wire DLX_EXinst_ALU_result_10_1;
  wire DLX_EXinst_ALU_result_11_1;
  wire DLX_EXinst_ALU_result_12_1;
  wire DLX_EXinst_ALU_result_13_1;
  wire DLX_EXinst_ALU_result_14_1;
  wire DLX_EXinst_ALU_result_5_1;
  wire DLX_EXinst_ALU_result_6_1;
  wire DLX_EXinst_ALU_result_7_1;
  wire DLX_EXinst_ALU_result_8_1;
  wire DLX_IDinst_mem_read;
  wire IR_MSB_0_OBUF;
  wire IR_MSB_1_OBUF;
  wire IR_MSB_3_OBUF;
  wire IR_MSB_7_OBUF;
  wire clk0;
  wire clk0buf;
  wire clkdivub;
  wire vga_top_vga1_Madd_addressout_inst_lut2_331;
  wire CHOICE5191;
  wire CHOICE4498;
  wire CHOICE4438;
  wire CHOICE3813;
  wire CHOICE3758;
  wire DLX_IDinst_RegFile_3_12;
  wire CHOICE3703;
  wire DLX_IDinst_RegFile_2_31;
  wire DLX_IDinst_RegFile_1_4;
  wire DLX_IDinst_RegFile_2_20;
  wire DLX_IDinst_RegFile_2_28;
  wire DLX_IDinst_RegFile_14_21;
  wire DLX_IDinst_RegFile_14_10;
  wire DLX_IDinst_RegFile_14_22;
  wire Mmux__COND_2__net2;
  wire DLX_IDinst_RegFile_22_14;
  wire N145733;
  wire vga_top_vga1_vcounter_Madd__n0000_inst_cy_10;
  wire GLOBAL_LOGIC1;
  wire GLOBAL_LOGIC0;
  wire vga_top_vga1_vcounter_Madd__n0000_inst_cy_12;
  wire vga_top_vga1_vcounter_Madd__n0000_inst_cy_14;
  wire vga_top_vga1_vcounter_Madd__n0000_inst_cy_16;
  wire DLX_EXinst_Mcompar__n0059_inst_cy_103;
  wire DLX_EXinst_Mcompar__n0059_inst_cy_105;
  wire DLX_EXinst_Mcompar__n0059_inst_cy_107;
  wire DLX_EXinst_Mcompar__n0059_inst_cy_109;
  wire DLX_EXinst_Mcompar__n0059_inst_cy_111;
  wire DLX_EXinst_Mcompar__n0059_inst_cy_113;
  wire DLX_IDinst_RegFile_14_12;
  wire DLX_EXinst_Mcompar__n0059_inst_cy_115;
  wire DLX_EXinst_Mcompar__n0067_inst_cy_199;
  wire DLX_EXinst_Mcompar__n0067_inst_cy_201;
  wire DLX_EXinst_Mcompar__n0067_inst_cy_203;
  wire DLX_EXinst_Mcompar__n0067_inst_cy_205;
  wire DLX_IDinst_RegFile_14_17;
  wire DLX_EXinst_Mcompar__n0067_inst_cy_207;
  wire DLX_EXinst_Mcompar__n0067_inst_cy_209;
  wire DLX_EXinst_Mcompar__n0067_inst_cy_211;
  wire DLX_EXinst_Mcompar__n0067_inst_cy_213;
  wire DLX_EXinst_Mcompar__n0067_inst_cy_215;
  wire DLX_EXinst_Mcompar__n0067_inst_cy_217;
  wire DLX_EXinst_Mcompar__n0067_inst_cy_219;
  wire DLX_EXinst_Mcompar__n0067_inst_cy_221;
  wire DLX_IDinst_RegFile_22_26;
  wire DLX_EXinst_Mcompar__n0067_inst_cy_223;
  wire DLX_EXinst_Mcompar__n0067_inst_cy_225;
  wire DLX_EXinst_Mcompar__n0067_inst_cy_227;
  wire vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_1;
  wire vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_3;
  wire vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_5;
  wire vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_7;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_167;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_169;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_171;
  wire DLX_IDinst_RegFile_22_30;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_173;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_175;
  wire DLX_IDinst_RegFile_1_6;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_177;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_179;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_181;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_183;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_185;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_187;
  wire DLX_IDinst_RegFile_22_23;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_189;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_191;
  wire DLX_IDinst_RegFile_15_11;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_193;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_195;
  wire DLX_IDinst_RegFile_3_6;
  wire DLX_IDinst_Msub__n0157_inst_cy_266;
  wire DLX_IDinst_Madd__n0158_inst_lut2_230;
  wire DLX_IDinst_RegFile_23_21;
  wire DLX_IDinst_Msub__n0157_inst_cy_268;
  wire DLX_IDinst_Msub__n0157_inst_cy_270;
  wire DLX_IDinst_Msub__n0157_inst_cy_272;
  wire DLX_IDinst_Msub__n0157_inst_cy_274;
  wire DLX_IDinst_Msub__n0157_inst_cy_276;
  wire DLX_IDinst_RegFile_15_20;
  wire DLX_IDinst_Msub__n0157_inst_cy_278;
  wire DLX_IDinst_Msub__n0157_inst_cy_280;
  wire DLX_IDinst_RegFile_14_16;
  wire DLX_IDinst_Msub__n0157_inst_cy_282;
  wire DLX_IDinst_Msub__n0157_inst_cy_284;
  wire DLX_IDinst_RegFile_23_12;
  wire DLX_IDinst_Msub__n0157_inst_cy_286;
  wire DLX_IDinst_Msub__n0157_inst_cy_288;
  wire DLX_IDinst_Msub__n0157_inst_cy_290;
  wire DLX_IDinst_Msub__n0157_inst_cy_292;
  wire DLX_IDinst_RegFile_1_7;
  wire DLX_IDinst_Msub__n0157_inst_cy_294;
  wire vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_1;
  wire vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_3;
  wire vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_5;
  wire vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_7;
  wire vga_top_vga1_hcounter_Madd__n0000_inst_cy_20;
  wire vga_top_vga1_hcounter_Madd__n0000_inst_cy_22;
  wire vga_top_vga1_hcounter_Madd__n0000_inst_cy_24;
  wire vga_top_vga1_hcounter_Madd__n0000_inst_cy_26;
  wire vga_top_vga1_hcounter_Madd__n0000_inst_cy_28;
  wire vga_top_vga1_hcounter_Madd__n0000_inst_cy_30;
  wire vga_top_vga1_hcounter_Madd__n0000_inst_cy_32;
  wire vga_top_vga1_Mmult__n0043_inst_cy_437;
  wire vga_top_vga1_Mmult__n0043_inst_lut2_317;
  wire vga_top_vga1_Mmult__n0043_inst_cy_439;
  wire vga_top_vga1_Mmult__n0043_inst_lut2_318;
  wire vga_top_vga1_Mmult__n0043_inst_lut2_319;
  wire DLX_IDinst_RegFile_3_14;
  wire vga_top_vga1_Mmult__n0043_inst_cy_441;
  wire vga_top_vga1_Mmult__n0043_inst_lut2_320;
  wire vga_top_vga1_Mmult__n0043_inst_lut2_321;
  wire vga_top_vga1_Mmult__n0043_inst_lut2_322;
  wire vga_top_vga1_Mmult__n0043_inst_lut2_323;
  wire vga_top_vga1_Mcompar__n0034_inst_cy_329;
  wire vga_top_vga1_Mcompar__n0034_inst_cy_331;
  wire vga_top_vga1_Mcompar__n0034_inst_cy_333;
  wire vga_top_vga1_Mcompar__n0034_inst_cy_335;
  wire vga_top_vga1_Mcompar__n0034_inst_cy_337;
  wire DLX_IDinst_RegFile_14_29;
  wire DLX_IDinst_RegFile_0_6;
  wire DLX_IDinst_RegFile_1_8;
  wire DLX_IDinst_RegFile_2_18;
  wire DLX_IDinst_RegFile_3_18;
  wire DLX_IDinst_RegFile_12_18;
  wire DLX_IDinst_RegFile_13_18;
  wire DLX_IDinst_RegFile_1_19;
  wire DLX_IDinst_RegFile_2_25;
  wire DLX_IDinst_RegFile_2_26;
  wire DLX_IDinst_RegFile_3_26;
  wire DLX_IDinst_RegFile_3_16;
  wire DLX_IDinst_RegFile_3_23;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_379;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_465;
  wire DLX_IDinst_RegFile_2_30;
  wire DLX_IDinst_RegFile_3_30;
  wire DLX_IDinst_RegFile_3_0;
  wire \DLX_IDinst_Cause_Reg[6] ;
  wire DLX_EXinst_Mcompar__n0065_inst_cy_167;
  wire DLX_EXinst_Mcompar__n0065_inst_cy_169;
  wire DLX_EXinst_Mcompar__n0065_inst_cy_171;
  wire DLX_EXinst_Mcompar__n0065_inst_cy_173;
  wire DLX_EXinst_Mcompar__n0065_inst_cy_175;
  wire DLX_EXinst_Mcompar__n0065_inst_cy_177;
  wire DLX_EXinst_Mcompar__n0065_inst_cy_179;
  wire DLX_EXinst_Mcompar__n0065_inst_cy_181;
  wire DLX_IDinst_RegFile_22_28;
  wire DLX_EXinst_Mcompar__n0065_inst_cy_183;
  wire DLX_EXinst_Mcompar__n0065_inst_cy_185;
  wire DLX_EXinst_Mcompar__n0065_inst_cy_187;
  wire DLX_EXinst_Mcompar__n0065_inst_cy_189;
  wire DLX_EXinst_Mcompar__n0065_inst_cy_191;
  wire DLX_EXinst_Mcompar__n0065_inst_cy_193;
  wire DLX_EXinst_Mcompar__n0065_inst_cy_195;
  wire vga_top_vga1_Mcompar__n0029_inst_cy_371;
  wire DLX_IDinst_RegFile_15_13;
  wire vga_top_vga1_Mcompar__n0029_inst_cy_373;
  wire vga_top_vga1_Mcompar__n0029_inst_cy_375;
  wire vga_top_vga1_Mcompar__n0037_inst_cy_472;
  wire vga_top_vga1_Mcompar__n0037_inst_cy_474;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_135;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_137;
  wire DLX_IDinst_RegFile_15_22;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_139;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_141;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_143;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_145;
  wire DLX_IDinst_RegFile_23_14;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_147;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_149;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_151;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_153;
  wire DLX_IDinst_RegFile_15_23;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_155;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_157;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_159;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_161;
  wire vga_top_vga1_Mcompar__n0030_inst_cy_355;
  wire vga_top_vga1_Mcompar__n0030_inst_cy_357;
  wire vga_top_vga1_Mcompar__n0030_inst_cy_359;
  wire vga_top_vga1_Mcompar__n0030_inst_cy_361;
  wire vga_top_vga1_Mcompar__n0030_inst_cy_363;
  wire vga_top_vga1_Mcompar__n0030_inst_cy_365;
  wire vga_top_vga1_Mcompar__n0030_inst_cy_367;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_135;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_137;
  wire DLX_IDinst_RegFile_23_16;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_139;
  wire vga_top_vga1_clockcounter_FFd2;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_141;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_143;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_145;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_147;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_149;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_151;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_153;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_155;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_157;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_159;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_161;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_163;
  wire DLX_IDinst_Mcompar__n0104_inst_cy_263;
  wire DLX_EXinst_Mcompar__n0061_inst_cy_119;
  wire DLX_EXinst_Mcompar__n0061_inst_cy_121;
  wire DLX_EXinst_Mcompar__n0061_inst_cy_123;
  wire DLX_EXinst_Mcompar__n0061_inst_cy_125;
  wire DLX_EXinst_Mcompar__n0061_inst_cy_127;
  wire DLX_EXinst_Mcompar__n0061_inst_cy_129;
  wire DLX_IDinst_RegFile_23_26;
  wire DLX_EXinst_Mcompar__n0061_inst_cy_131;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_571;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_741;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_923;
  wire DLX_EXinst_Maddsub__n0012_inst_cy_71;
  wire DLX_EXinst_Maddsub__n0012_inst_cy_73;
  wire DLX_EXinst_Maddsub__n0012_inst_cy_75;
  wire DLX_EXinst_Maddsub__n0012_inst_cy_77;
  wire DLX_EXinst_Maddsub__n0012_inst_cy_79;
  wire DLX_EXinst_Maddsub__n0012_inst_cy_81;
  wire DLX_EXinst_Maddsub__n0012_inst_cy_83;
  wire DLX_EXinst_Maddsub__n0012_inst_cy_85;
  wire DLX_EXinst_Maddsub__n0012_inst_cy_87;
  wire DLX_EXinst_Maddsub__n0012_inst_cy_89;
  wire DLX_EXinst_Maddsub__n0012_inst_cy_91;
  wire DLX_EXinst_Maddsub__n0012_inst_cy_93;
  wire DLX_EXinst_Maddsub__n0012_inst_cy_95;
  wire DLX_EXinst_Maddsub__n0012_inst_cy_97;
  wire DLX_EXinst_Maddsub__n0012_inst_cy_99;
  wire DLX_EXinst_Mcompar__n0087_inst_cy_119;
  wire DLX_EXinst_Mcompar__n0087_inst_cy_121;
  wire DLX_EXinst_Mcompar__n0087_inst_cy_123;
  wire DLX_EXinst_Mcompar__n0087_inst_cy_125;
  wire DLX_EXinst_Mcompar__n0087_inst_cy_127;
  wire DLX_EXinst_Mcompar__n0087_inst_cy_129;
  wire DLX_EXinst_Mcompar__n0087_inst_cy_131;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_231;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_233;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_235;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_237;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_239;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_241;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_243;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_245;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_247;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_249;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_251;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_253;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_255;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_257;
  wire DLX_IDinst_Madd__n0158_inst_cy_298;
  wire DLX_IDinst_Madd__n0158_inst_cy_300;
  wire DLX_IDinst_Madd__n0158_inst_cy_302;
  wire DLX_IDinst_Madd__n0158_inst_cy_304;
  wire DLX_IDinst_Madd__n0158_inst_cy_306;
  wire DLX_IDinst_Madd__n0158_inst_cy_308;
  wire DLX_IDinst_Madd__n0158_inst_cy_310;
  wire DLX_IDinst_Madd__n0158_inst_cy_312;
  wire DLX_IDinst_Madd__n0158_inst_cy_314;
  wire DLX_IDinst_Madd__n0158_inst_cy_316;
  wire DLX_IDinst_Madd__n0158_inst_cy_318;
  wire DLX_IDinst_Madd__n0158_inst_cy_320;
  wire DLX_IDinst_Madd__n0158_inst_cy_322;
  wire DLX_IDinst_Madd__n0158_inst_cy_324;
  wire DLX_IDinst_Madd__n0158_inst_cy_326;
  wire DLX_IDinst_Mcompar__n0102_inst_cy_263;
  wire vga_top_vga1_Mcompar__n0033_inst_cy_341;
  wire vga_top_vga1_Mcompar__n0033_inst_cy_343;
  wire vga_top_vga1_Mcompar__n0033_inst_cy_345;
  wire vga_top_vga1_Mcompar__n0033_inst_cy_347;
  wire vga_top_vga1_Mcompar__n0033_inst_cy_349;
  wire vga_top_vga1_Mcompar__n0033_inst_cy_351;
  wire vga_top_vga1_Madd_addressout_inst_cy_463;
  wire vga_top_vga1_Madd_addressout_inst_cy_465;
  wire vga_top_vga1_Madd_addressout_inst_cy_467;
  wire vga_top_vga1_Madd_addressout_inst_cy_469;
  wire DLX_IFinst_Madd__n0005_inst_cy_41;
  wire DLX_IFinst_Madd__n0005_inst_cy_43;
  wire DLX_IFinst_Madd__n0005_inst_cy_45;
  wire DLX_IFinst_Madd__n0005_inst_cy_47;
  wire DLX_IFinst_Madd__n0005_inst_cy_49;
  wire DLX_IFinst_Madd__n0005_inst_cy_51;
  wire DLX_IFinst_Madd__n0005_inst_cy_53;
  wire DLX_IFinst_Madd__n0005_inst_cy_55;
  wire DLX_IFinst_Madd__n0005_inst_cy_57;
  wire DLX_IFinst_Madd__n0005_inst_cy_59;
  wire DLX_IFinst_Madd__n0005_inst_cy_61;
  wire DLX_IFinst_Madd__n0005_inst_cy_63;
  wire DLX_IFinst_Madd__n0005_inst_cy_65;
  wire DLX_IFinst_Madd__n0005_inst_cy_67;
  wire DLX_EXinst_Mcompar__n0085_inst_cy_103;
  wire DLX_EXinst_Mcompar__n0085_inst_cy_105;
  wire DLX_EXinst_Mcompar__n0085_inst_cy_107;
  wire DLX_EXinst_Mcompar__n0085_inst_cy_109;
  wire DLX_EXinst_Mcompar__n0085_inst_cy_111;
  wire DLX_EXinst_Mcompar__n0085_inst_cy_113;
  wire DLX_EXinst_Mcompar__n0085_inst_cy_115;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_199;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_201;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_203;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_205;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_207;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_209;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_211;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_213;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_215;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_217;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_219;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_221;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_223;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_225;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_227;
  wire DLX_EXinst_Mcompar__n0069_inst_cy_231;
  wire DLX_EXinst_Mcompar__n0069_inst_cy_233;
  wire DLX_EXinst_Mcompar__n0069_inst_cy_235;
  wire DLX_EXinst_Mcompar__n0069_inst_cy_237;
  wire DLX_EXinst_Mcompar__n0069_inst_cy_239;
  wire DLX_EXinst_Mcompar__n0069_inst_cy_241;
  wire DLX_EXinst_Mcompar__n0069_inst_cy_243;
  wire DLX_EXinst_Mcompar__n0069_inst_cy_245;
  wire DLX_EXinst_Mcompar__n0069_inst_cy_247;
  wire DLX_EXinst_Mcompar__n0069_inst_cy_249;
  wire DLX_EXinst_Mcompar__n0069_inst_cy_251;
  wire DLX_EXinst_Mcompar__n0069_inst_cy_253;
  wire DLX_EXinst_Mcompar__n0069_inst_cy_255;
  wire DLX_EXinst_Mcompar__n0069_inst_cy_257;
  wire DLX_EXinst_Mcompar__n0069_inst_cy_259;
  wire DLX_IDinst_Mcompar__n0100_inst_cy_263;
  wire DLX_IDinst_Mcompar__n0105_inst_cy_263;
  wire DLX_IDinst_Mcompar__n0367_inst_cy_263;
  wire N162867;
  wire N162828;
  wire N162832;
  wire N162857;
  wire N162813;
  wire N162844;
  wire DLX_IDinst_RegFile_12_10;
  wire DLX_IDinst_RegFile_13_10;
  wire DLX_IDinst_RegFile_15_10;
  wire DLX_IDinst_RegFile_20_10;
  wire DLX_IDinst_RegFile_21_10;
  wire DLX_IDinst_RegFile_22_10;
  wire DLX_IDinst_RegFile_12_11;
  wire DLX_IDinst_RegFile_13_11;
  wire DLX_IDinst_RegFile_14_11;
  wire DLX_IDinst_RegFile_20_11;
  wire DLX_IDinst_RegFile_21_11;
  wire DLX_IDinst_RegFile_23_11;
  wire DLX_IDinst_RegFile_12_20;
  wire DLX_IDinst_RegFile_13_20;
  wire DLX_IDinst_RegFile_14_20;
  wire DLX_IDinst_RegFile_12_12;
  wire DLX_IDinst_RegFile_13_12;
  wire DLX_IDinst_RegFile_15_12;
  wire DLX_IDinst_RegFile_20_20;
  wire DLX_IDinst_RegFile_21_20;
  wire DLX_IDinst_RegFile_23_20;
  wire DLX_IDinst_RegFile_20_12;
  wire DLX_IDinst_RegFile_21_12;
  wire DLX_IDinst_RegFile_22_12;
  wire DLX_IDinst_RegFile_12_21;
  wire DLX_IDinst_RegFile_13_21;
  wire DLX_IDinst_RegFile_15_21;
  wire DLX_IDinst_RegFile_12_13;
  wire DLX_IDinst_RegFile_13_13;
  wire DLX_IDinst_RegFile_14_13;
  wire DLX_IDinst_RegFile_20_21;
  wire DLX_IDinst_RegFile_21_21;
  wire DLX_IDinst_RegFile_22_21;
  wire DLX_IDinst_RegFile_20_13;
  wire DLX_IDinst_RegFile_21_13;
  wire DLX_IDinst_RegFile_23_13;
  wire DLX_IDinst_RegFile_12_30;
  wire DLX_IDinst_RegFile_13_30;
  wire DLX_IDinst_RegFile_14_30;
  wire DLX_IDinst_RegFile_15_30;
  wire DLX_IDinst_RegFile_12_22;
  wire DLX_IDinst_RegFile_13_22;
  wire DLX_IDinst_RegFile_12_14;
  wire DLX_IDinst_RegFile_13_14;
  wire DLX_IDinst_RegFile_14_14;
  wire DLX_IDinst_RegFile_15_14;
  wire DLX_IDinst_RegFile_20_30;
  wire DLX_IDinst_RegFile_21_30;
  wire DLX_IDinst_RegFile_20_22;
  wire DLX_IDinst_RegFile_21_22;
  wire DLX_IDinst_RegFile_22_22;
  wire DLX_IDinst_RegFile_23_22;
  wire DLX_IDinst_RegFile_20_14;
  wire DLX_IDinst_RegFile_21_14;
  wire DLX_IDinst_RegFile_12_23;
  wire DLX_IDinst_RegFile_13_23;
  wire DLX_IDinst_RegFile_12_15;
  wire DLX_IDinst_RegFile_13_15;
  wire DLX_IDinst_RegFile_14_15;
  wire DLX_IDinst_RegFile_15_15;
  wire DLX_IDinst_RegFile_20_23;
  wire DLX_IDinst_RegFile_21_23;
  wire DLX_IDinst_RegFile_20_15;
  wire DLX_IDinst_RegFile_21_15;
  wire DLX_IDinst_RegFile_22_15;
  wire DLX_IDinst_RegFile_23_15;
  wire DLX_IDinst_RegFile_12_31;
  wire DLX_IDinst_RegFile_13_31;
  wire DLX_IDinst_RegFile_20_31;
  wire DLX_IDinst_RegFile_21_31;
  wire DLX_IDinst_RegFile_22_31;
  wire DLX_IDinst_RegFile_23_31;
  wire DLX_IDinst_RegFile_12_24;
  wire DLX_IDinst_RegFile_13_24;
  wire DLX_IDinst_RegFile_14_24;
  wire DLX_IDinst_RegFile_15_24;
  wire DLX_IDinst_RegFile_12_16;
  wire DLX_IDinst_RegFile_13_16;
  wire DLX_IDinst_RegFile_20_24;
  wire DLX_IDinst_RegFile_21_24;
  wire DLX_IDinst_RegFile_22_24;
  wire DLX_IDinst_RegFile_23_24;
  wire DLX_IDinst_RegFile_20_16;
  wire DLX_IDinst_RegFile_21_16;
  wire DLX_IDinst_RegFile_12_25;
  wire DLX_IDinst_RegFile_13_25;
  wire DLX_IDinst_RegFile_14_25;
  wire DLX_IDinst_RegFile_15_25;
  wire DLX_IDinst_RegFile_12_17;
  wire DLX_IDinst_RegFile_13_17;
  wire DLX_IDinst_RegFile_20_25;
  wire DLX_IDinst_RegFile_21_25;
  wire DLX_IDinst_RegFile_22_25;
  wire DLX_IDinst_RegFile_23_25;
  wire DLX_IDinst_RegFile_20_17;
  wire DLX_IDinst_RegFile_21_17;
  wire DLX_IDinst_RegFile_12_26;
  wire DLX_IDinst_RegFile_13_26;
  wire DLX_IDinst_RegFile_14_26;
  wire DLX_IDinst_RegFile_15_26;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_679;
  wire DLX_IDinst_RegFile_20_26;
  wire DLX_IDinst_RegFile_21_26;
  wire DLX_IDinst_RegFile_20_18;
  wire DLX_IDinst_RegFile_21_18;
  wire DLX_IDinst_RegFile_22_18;
  wire DLX_IDinst_RegFile_23_18;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_681;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_683;
  wire DLX_IDinst_RegFile_12_27;
  wire DLX_IDinst_RegFile_13_27;
  wire DLX_IDinst_RegFile_15_27;
  wire DLX_IDinst_RegFile_12_19;
  wire DLX_IDinst_RegFile_13_19;
  wire DLX_IDinst_RegFile_14_19;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_695;
  wire DLX_IDinst_RegFile_20_27;
  wire DLX_IDinst_RegFile_21_27;
  wire DLX_IDinst_RegFile_22_27;
  wire DLX_IDinst_RegFile_20_19;
  wire DLX_IDinst_RegFile_21_19;
  wire DLX_IDinst_RegFile_23_19;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_697;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_699;
  wire DLX_IDinst_RegFile_12_28;
  wire DLX_IDinst_RegFile_13_28;
  wire DLX_IDinst_RegFile_14_28;
  wire DLX_IDinst_RegFile_15_28;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_839;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_711;
  wire DLX_IDinst_RegFile_20_28;
  wire DLX_IDinst_RegFile_21_28;
  wire DLX_IDinst_RegFile_23_28;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_841;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_713;
  wire DLX_IDinst_RegFile_12_29;
  wire DLX_IDinst_RegFile_13_29;
  wire DLX_IDinst_RegFile_15_29;
  wire DLX_IDinst_RegFile_20_29;
  wire DLX_IDinst_RegFile_21_29;
  wire DLX_IDinst_RegFile_22_29;
  wire DLX_IDinst_RegFile_23_29;
  wire CHOICE3150;
  wire GSR = glbl.GSR;
  wire GTS = glbl.GTS;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1047;
  wire \DLX_IDinst_RegFile_25_28/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1048;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_972;
  wire \DLX_IDinst_RegFile_25_28/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_25_28/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_391;
  wire \DLX_IDinst_RegFile_26_20/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_392;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_332;
  wire \DLX_IDinst_RegFile_26_20/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_26_20/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_263;
  wire \DLX_IDinst_RegFile_26_12/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_264;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_204;
  wire \DLX_IDinst_RegFile_26_12/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_26_12/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1059;
  wire \DLX_IDinst_RegFile_17_29/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1060;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_984;
  wire \DLX_IDinst_RegFile_17_29/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_17_29/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_403;
  wire \DLX_IDinst_RegFile_18_21/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_404;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_344;
  wire \DLX_IDinst_RegFile_18_21/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_18_21/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_275;
  wire \DLX_IDinst_RegFile_18_13/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_276;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_216;
  wire \DLX_IDinst_RegFile_18_13/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_18_13/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1063;
  wire \DLX_IDinst_RegFile_25_29/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1064;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_988;
  wire \DLX_IDinst_RegFile_25_29/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_25_29/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_407;
  wire \DLX_IDinst_RegFile_26_21/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_408;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_348;
  wire \DLX_IDinst_RegFile_26_21/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_26_21/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_279;
  wire \DLX_IDinst_RegFile_26_13/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_280;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_220;
  wire \DLX_IDinst_RegFile_26_13/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_26_13/CYINIT ;
  wire \CHOICE3470/GROM ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1075;
  wire \DLX_IDinst_RegFile_18_30/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1076;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_1000;
  wire \DLX_IDinst_RegFile_18_30/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_18_30/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_419;
  wire \DLX_IDinst_RegFile_18_22/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_420;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_360;
  wire \DLX_IDinst_RegFile_18_22/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_18_22/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_291;
  wire \DLX_IDinst_RegFile_18_14/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_292;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_232;
  wire \DLX_IDinst_RegFile_18_14/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_18_14/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1079;
  wire \DLX_IDinst_RegFile_26_30/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1080;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_1004;
  wire \DLX_IDinst_RegFile_26_30/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_26_30/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_423;
  wire \DLX_IDinst_RegFile_26_22/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_424;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_364;
  wire \DLX_IDinst_RegFile_26_22/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_26_22/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_295;
  wire \DLX_IDinst_RegFile_26_14/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_296;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_236;
  wire \DLX_IDinst_RegFile_26_14/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_26_14/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_435;
  wire \DLX_IDinst_RegFile_18_23/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_436;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_376;
  wire \DLX_IDinst_RegFile_18_23/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_18_23/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_307;
  wire \DLX_IDinst_RegFile_18_15/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_308;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_248;
  wire \DLX_IDinst_RegFile_18_15/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_18_15/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_967;
  wire \DLX_IDinst_RegFile_26_23/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_968;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_892;
  wire \DLX_IDinst_RegFile_26_23/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_26_23/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_311;
  wire \DLX_IDinst_RegFile_26_15/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_312;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_252;
  wire \DLX_IDinst_RegFile_26_15/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_26_15/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1091;
  wire \DLX_IDinst_RegFile_18_31/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1092;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_1016;
  wire \DLX_IDinst_RegFile_18_31/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_18_31/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1095;
  wire \DLX_IDinst_RegFile_26_31/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1096;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_1020;
  wire \DLX_IDinst_RegFile_26_31/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_26_31/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_451;
  wire \DLX_IDinst_RegFile_18_24/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_452;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_392;
  wire \DLX_IDinst_RegFile_18_24/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_18_24/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_323;
  wire \DLX_IDinst_RegFile_18_16/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_324;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_264;
  wire \DLX_IDinst_RegFile_18_16/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_18_16/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_455;
  wire \DLX_IDinst_RegFile_26_24/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_456;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_396;
  wire \DLX_IDinst_RegFile_26_24/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_26_24/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_327;
  wire \DLX_IDinst_RegFile_26_16/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_328;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_268;
  wire \DLX_IDinst_RegFile_26_16/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_26_16/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_467;
  wire \DLX_IDinst_RegFile_18_25/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_468;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_408;
  wire \DLX_IDinst_RegFile_18_25/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_18_25/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_339;
  wire \DLX_IDinst_RegFile_18_17/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_340;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_280;
  wire \DLX_IDinst_RegFile_18_17/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_18_17/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_471;
  wire \DLX_IDinst_RegFile_26_25/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_472;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_412;
  wire \DLX_IDinst_RegFile_26_25/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_26_25/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_343;
  wire \DLX_IDinst_RegFile_26_17/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_344;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_284;
  wire \DLX_IDinst_RegFile_26_17/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_26_17/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_483;
  wire \DLX_IDinst_RegFile_18_26/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_484;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_424;
  wire \DLX_IDinst_RegFile_18_26/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_18_26/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_355;
  wire \DLX_IDinst_RegFile_18_18/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_356;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_296;
  wire \DLX_IDinst_RegFile_18_18/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_18_18/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_227;
  wire \DLX_IDinst_RegFile_19_10/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_228;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_168;
  wire \DLX_IDinst_RegFile_19_10/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_19_10/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_487;
  wire \DLX_IDinst_RegFile_26_26/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_488;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_428;
  wire \DLX_IDinst_RegFile_26_26/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_26_26/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_359;
  wire \DLX_IDinst_RegFile_26_18/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_360;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_300;
  wire \DLX_IDinst_RegFile_26_18/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_26_18/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_231;
  wire \DLX_IDinst_RegFile_27_10/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_232;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_172;
  wire \DLX_IDinst_RegFile_27_10/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_27_10/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1027;
  wire \DLX_IDinst_RegFile_18_27/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1028;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_952;
  wire \DLX_IDinst_RegFile_18_27/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_18_27/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_371;
  wire \DLX_IDinst_RegFile_18_19/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_372;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_312;
  wire \DLX_IDinst_RegFile_18_19/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_18_19/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_243;
  wire \DLX_IDinst_RegFile_19_11/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_244;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_184;
  wire \DLX_IDinst_RegFile_19_11/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_19_11/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1031;
  wire \DLX_IDinst_RegFile_26_27/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1032;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_956;
  wire \DLX_IDinst_RegFile_26_27/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_26_27/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_375;
  wire \DLX_IDinst_RegFile_26_19/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_376;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_316;
  wire \DLX_IDinst_RegFile_26_19/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_26_19/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_247;
  wire \DLX_IDinst_RegFile_27_11/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_248;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_188;
  wire \DLX_IDinst_RegFile_27_11/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_27_11/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1043;
  wire \DLX_IDinst_RegFile_18_28/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1044;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_968;
  wire \DLX_IDinst_RegFile_18_28/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_18_28/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_387;
  wire \DLX_IDinst_RegFile_19_20/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_388;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_328;
  wire \DLX_IDinst_RegFile_19_20/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_19_20/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_259;
  wire \DLX_IDinst_RegFile_19_12/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_260;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_200;
  wire \DLX_IDinst_RegFile_19_12/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_19_12/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_519;
  wire \DLX_IDinst_RegFile_26_28/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_520;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_460;
  wire \DLX_IDinst_RegFile_26_28/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_26_28/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_919;
  wire \DLX_IDinst_RegFile_27_20/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_920;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_844;
  wire \DLX_IDinst_RegFile_27_20/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_27_20/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_791;
  wire \DLX_IDinst_RegFile_27_12/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_792;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_716;
  wire \DLX_IDinst_RegFile_27_12/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_27_12/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_531;
  wire \DLX_IDinst_RegFile_18_29/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_532;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_472;
  wire \DLX_IDinst_RegFile_18_29/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_18_29/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_931;
  wire \DLX_IDinst_RegFile_19_21/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_932;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_856;
  wire \DLX_IDinst_RegFile_19_21/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_19_21/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_803;
  wire \DLX_IDinst_RegFile_19_13/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_804;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_728;
  wire \DLX_IDinst_RegFile_19_13/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_19_13/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_535;
  wire \DLX_IDinst_RegFile_26_29/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_536;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_476;
  wire \DLX_IDinst_RegFile_26_29/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_26_29/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_935;
  wire \DLX_IDinst_RegFile_27_21/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_936;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_860;
  wire \DLX_IDinst_RegFile_27_21/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_27_21/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_807;
  wire \DLX_IDinst_RegFile_27_13/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_808;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_732;
  wire \DLX_IDinst_RegFile_27_13/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_27_13/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_547;
  wire \DLX_IDinst_RegFile_19_30/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_548;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_488;
  wire \DLX_IDinst_RegFile_19_30/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_19_30/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_947;
  wire \DLX_IDinst_RegFile_19_22/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_948;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_872;
  wire \DLX_IDinst_RegFile_19_22/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_19_22/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_819;
  wire \DLX_IDinst_RegFile_19_14/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_820;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_744;
  wire \DLX_IDinst_RegFile_19_14/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_19_14/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_551;
  wire \DLX_IDinst_RegFile_27_30/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_552;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_492;
  wire \DLX_IDinst_RegFile_27_30/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_27_30/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_951;
  wire \DLX_IDinst_RegFile_27_22/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_952;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_876;
  wire \DLX_IDinst_RegFile_27_22/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_27_22/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_823;
  wire \DLX_IDinst_RegFile_27_14/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_824;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_748;
  wire \DLX_IDinst_RegFile_27_14/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_27_14/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_963;
  wire \DLX_IDinst_RegFile_19_23/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_964;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_888;
  wire \DLX_IDinst_RegFile_19_23/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_19_23/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_835;
  wire \DLX_IDinst_RegFile_19_15/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_836;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_760;
  wire \DLX_IDinst_RegFile_19_15/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_19_15/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_839;
  wire \DLX_IDinst_RegFile_27_15/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_840;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_764;
  wire \DLX_IDinst_RegFile_27_15/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_27_15/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_563;
  wire \DLX_IDinst_RegFile_19_31/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_564;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_504;
  wire \DLX_IDinst_RegFile_19_31/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_19_31/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_567;
  wire \DLX_IDinst_RegFile_27_31/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_568;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_508;
  wire \DLX_IDinst_RegFile_27_31/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_27_31/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_979;
  wire \DLX_IDinst_RegFile_19_24/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_980;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_904;
  wire \DLX_IDinst_RegFile_19_24/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_19_24/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_851;
  wire \DLX_IDinst_RegFile_19_16/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_852;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_776;
  wire \DLX_IDinst_RegFile_19_16/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_19_16/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_983;
  wire \DLX_IDinst_RegFile_27_24/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_984;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_908;
  wire \DLX_IDinst_RegFile_27_24/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_27_24/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_855;
  wire \DLX_IDinst_RegFile_27_16/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_856;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_780;
  wire \DLX_IDinst_RegFile_27_16/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_27_16/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_995;
  wire \DLX_IDinst_RegFile_19_25/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_996;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_920;
  wire \DLX_IDinst_RegFile_19_25/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_19_25/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_867;
  wire \DLX_IDinst_RegFile_19_17/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_868;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_792;
  wire \DLX_IDinst_RegFile_19_17/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_19_17/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_871;
  wire \DLX_IDinst_RegFile_27_17/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_872;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_796;
  wire \DLX_IDinst_RegFile_27_17/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_27_17/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1011;
  wire \DLX_IDinst_RegFile_19_26/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1012;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_936;
  wire \DLX_IDinst_RegFile_19_26/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_19_26/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_883;
  wire \DLX_IDinst_RegFile_19_18/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_884;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_808;
  wire \DLX_IDinst_RegFile_19_18/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_19_18/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1015;
  wire \DLX_IDinst_RegFile_27_26/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1016;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_940;
  wire \DLX_IDinst_RegFile_27_26/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_27_26/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_887;
  wire \DLX_IDinst_RegFile_27_18/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_888;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_812;
  wire \DLX_IDinst_RegFile_27_18/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_27_18/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_233;
  wire \DLX_IDinst_RegFile_28_10/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_234;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_174;
  wire \DLX_IDinst_RegFile_28_10/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_28_10/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_499;
  wire \DLX_IDinst_RegFile_19_27/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_500;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_440;
  wire \DLX_IDinst_RegFile_19_27/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_19_27/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_899;
  wire \DLX_IDinst_RegFile_19_19/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_900;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_824;
  wire \DLX_IDinst_RegFile_19_19/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_19_19/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_503;
  wire \DLX_IDinst_RegFile_27_27/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_504;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_444;
  wire \DLX_IDinst_RegFile_27_27/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_27_27/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_903;
  wire \DLX_IDinst_RegFile_27_19/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_904;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_828;
  wire \DLX_IDinst_RegFile_27_19/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_27_19/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_249;
  wire \DLX_IDinst_RegFile_28_11/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_250;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_190;
  wire \DLX_IDinst_RegFile_28_11/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_28_11/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_515;
  wire \DLX_IDinst_RegFile_19_28/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_516;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_456;
  wire \DLX_IDinst_RegFile_19_28/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_19_28/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_393;
  wire \DLX_IDinst_RegFile_28_20/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_394;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_334;
  wire \DLX_IDinst_RegFile_28_20/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_28_20/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_265;
  wire \DLX_IDinst_RegFile_28_12/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_266;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_206;
  wire \DLX_IDinst_RegFile_28_12/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_28_12/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_409;
  wire \DLX_IDinst_RegFile_28_21/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_410;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_350;
  wire \DLX_IDinst_RegFile_28_21/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_28_21/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_281;
  wire \DLX_IDinst_RegFile_28_13/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_282;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_222;
  wire \DLX_IDinst_RegFile_28_13/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_28_13/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1081;
  wire \DLX_IDinst_RegFile_28_30/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1082;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_1006;
  wire \DLX_IDinst_RegFile_28_30/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_28_30/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_425;
  wire \DLX_IDinst_RegFile_28_22/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_426;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_366;
  wire \DLX_IDinst_RegFile_28_22/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_28_22/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_297;
  wire \DLX_IDinst_RegFile_28_14/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_298;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_238;
  wire \DLX_IDinst_RegFile_28_14/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_28_14/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_441;
  wire \DLX_IDinst_RegFile_28_23/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_442;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_382;
  wire \DLX_IDinst_RegFile_28_23/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_28_23/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_313;
  wire \DLX_IDinst_RegFile_28_15/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_314;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_254;
  wire \DLX_IDinst_RegFile_28_15/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_28_15/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1097;
  wire \DLX_IDinst_RegFile_28_31/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1098;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_1022;
  wire \DLX_IDinst_RegFile_28_31/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_28_31/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_457;
  wire \DLX_IDinst_RegFile_28_24/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_458;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_398;
  wire \DLX_IDinst_RegFile_28_24/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_28_24/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_329;
  wire \DLX_IDinst_RegFile_28_16/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_330;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_270;
  wire \DLX_IDinst_RegFile_28_16/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_28_16/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_473;
  wire \DLX_IDinst_RegFile_28_25/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_474;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_414;
  wire \DLX_IDinst_RegFile_28_25/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_28_25/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_345;
  wire \DLX_IDinst_RegFile_28_17/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_346;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_286;
  wire \DLX_IDinst_RegFile_28_17/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_28_17/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_489;
  wire \DLX_IDinst_RegFile_28_26/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_490;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_430;
  wire \DLX_IDinst_RegFile_28_26/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_28_26/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_361;
  wire \DLX_IDinst_RegFile_28_18/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_362;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_302;
  wire \DLX_IDinst_RegFile_28_18/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_28_18/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_761;
  wire \DLX_IDinst_RegFile_29_10/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_762;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_686;
  wire \DLX_IDinst_RegFile_29_10/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_29_10/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_505;
  wire \DLX_IDinst_RegFile_28_27/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_506;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_446;
  wire \DLX_IDinst_RegFile_28_27/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_28_27/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_377;
  wire \DLX_IDinst_RegFile_28_19/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_378;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_318;
  wire \DLX_IDinst_RegFile_28_19/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_28_19/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_777;
  wire \DLX_IDinst_RegFile_29_11/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_778;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_702;
  wire \DLX_IDinst_RegFile_29_11/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_29_11/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1049;
  wire \DLX_IDinst_RegFile_28_28/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1050;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_974;
  wire \DLX_IDinst_RegFile_28_28/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_28_28/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_921;
  wire \DLX_IDinst_RegFile_29_20/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_922;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_846;
  wire \DLX_IDinst_RegFile_29_20/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_29_20/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_793;
  wire \DLX_IDinst_RegFile_29_12/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_794;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_718;
  wire \DLX_IDinst_RegFile_29_12/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_29_12/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1065;
  wire \DLX_IDinst_RegFile_28_29/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1066;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_990;
  wire \DLX_IDinst_RegFile_28_29/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_28_29/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_937;
  wire \DLX_IDinst_RegFile_29_21/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_938;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_862;
  wire \DLX_IDinst_RegFile_29_21/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_29_21/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_809;
  wire \DLX_IDinst_RegFile_29_13/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_810;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_734;
  wire \DLX_IDinst_RegFile_29_13/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_29_13/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_553;
  wire \DLX_IDinst_RegFile_29_30/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_554;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_494;
  wire \DLX_IDinst_RegFile_29_30/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_29_30/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_953;
  wire \DLX_IDinst_RegFile_29_22/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_954;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_878;
  wire \DLX_IDinst_RegFile_29_22/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_29_22/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_825;
  wire \DLX_IDinst_RegFile_29_14/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_826;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_750;
  wire \DLX_IDinst_RegFile_29_14/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_29_14/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_969;
  wire \DLX_IDinst_RegFile_29_23/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_970;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_894;
  wire \DLX_IDinst_RegFile_29_23/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_29_23/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_841;
  wire \DLX_IDinst_RegFile_29_15/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_842;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_766;
  wire \DLX_IDinst_RegFile_29_15/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_29_15/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_569;
  wire \DLX_IDinst_RegFile_29_31/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_570;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_510;
  wire \DLX_IDinst_RegFile_29_31/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_29_31/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_985;
  wire \DLX_IDinst_RegFile_29_24/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_986;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_910;
  wire \DLX_IDinst_RegFile_29_24/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_29_24/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_857;
  wire \DLX_IDinst_RegFile_29_16/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_858;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_782;
  wire \DLX_IDinst_RegFile_29_16/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_29_16/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1001;
  wire \DLX_IDinst_RegFile_29_25/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1002;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_926;
  wire \DLX_IDinst_RegFile_29_25/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_29_25/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_873;
  wire \DLX_IDinst_RegFile_29_17/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_874;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_798;
  wire \DLX_IDinst_RegFile_29_17/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_29_17/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1017;
  wire \DLX_IDinst_RegFile_29_26/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1018;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_942;
  wire \DLX_IDinst_RegFile_29_26/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_29_26/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_889;
  wire \DLX_IDinst_RegFile_29_18/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_890;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_814;
  wire \DLX_IDinst_RegFile_29_18/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_29_18/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1033;
  wire \DLX_IDinst_RegFile_29_27/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1034;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_958;
  wire \DLX_IDinst_RegFile_29_27/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_29_27/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_905;
  wire \DLX_IDinst_RegFile_29_19/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_906;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_830;
  wire \DLX_IDinst_RegFile_29_19/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_29_19/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_521;
  wire \DLX_IDinst_RegFile_29_28/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_522;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_462;
  wire \DLX_IDinst_RegFile_29_28/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_29_28/CYINIT ;
  wire \DLX_EXinst__n0127/FROM ;
  wire \DLX_EXinst__n0127/GROM ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_537;
  wire \DLX_IDinst_RegFile_29_29/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_538;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_478;
  wire \DLX_IDinst_RegFile_29_29/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_29_29/CYINIT ;
  wire \CHOICE3008/FROM ;
  wire \CHOICE3008/GROM ;
  wire \CHOICE3575/FROM ;
  wire \CHOICE3575/GROM ;
  wire \CHOICE3442/FROM ;
  wire \CHOICE3442/GROM ;
  wire \DLX_IFinst_IR_previous<26>/FROM ;
  wire \DLX_IFinst_IR_previous<26>/GROM ;
  wire \DLX_IDinst_RegFile_1_28/FROM ;
  wire \DLX_IDinst_RegFile_1_28/GROM ;
  wire \DLX_EXinst_reg_out_B_EX<4>/FROM ;
  wire \DLX_EXinst_reg_out_B_EX<4>/GROM ;
  wire \DLX_IDinst_RegFile_1_29/FROM ;
  wire \DLX_IDinst_RegFile_1_29/GROM ;
  wire \CHOICE3590/FROM ;
  wire \CHOICE3590/GROM ;
  wire \CHOICE3592/FROM ;
  wire \CHOICE3592/GROM ;
  wire \DLX_IDinst_RegFile_22_20/FROM ;
  wire \DLX_IDinst_RegFile_22_20/GROM ;
  wire \N163298/FROM ;
  wire \N163298/GROM ;
  wire \CHOICE1313/FROM ;
  wire \CHOICE1313/GROM ;
  wire \DLX_IDinst_IR_opcode_field<1>/FROM ;
  wire \N163469/FROM ;
  wire \N163469/GROM ;
  wire \DLX_IDinst_IR_opcode_field<3>/FROM ;
  wire \DLX_IDinst_IR_opcode_field<4>/FROM ;
  wire \DLX_IDinst_Imm<0>/FROM ;
  wire \DLX_IDinst_Imm<0>/GROM ;
  wire \DLX_IDinst_RegFile_2_6/FROM ;
  wire \DLX_IDinst_RegFile_2_6/GROM ;
  wire \N164178/FROM ;
  wire \N164178/GROM ;
  wire \DLX_EXinst_Mshift__n0020_Sh<30>/FROM ;
  wire \DLX_EXinst_Mshift__n0020_Sh<30>/GROM ;
  wire \DLX_EXinst_Mshift__n0020_Sh<61>/FROM ;
  wire \DLX_EXinst_Mshift__n0020_Sh<61>/GROM ;
  wire \DLX_EXinst_Mshift__n0020_Sh<29>/FROM ;
  wire \DLX_EXinst_Mshift__n0020_Sh<29>/GROM ;
  wire \CHOICE4693/FROM ;
  wire \CHOICE4693/GROM ;
  wire \CHOICE3809/FROM ;
  wire \CHOICE3809/GROM ;
  wire \CHOICE4172/FROM ;
  wire \CHOICE4172/GROM ;
  wire \CHOICE3685/FROM ;
  wire \CHOICE3685/GROM ;
  wire \CHOICE3969/FROM ;
  wire \CHOICE3969/GROM ;
  wire \DLX_IDinst_RegFile_3_10/FROM ;
  wire \DLX_IDinst_RegFile_3_10/GROM ;
  wire \CHOICE3859/FROM ;
  wire \CHOICE3859/GROM ;
  wire \CHOICE4730/GROM ;
  wire \DLX_EXinst_N76268/FROM ;
  wire \DLX_EXinst_N76268/GROM ;
  wire \CHOICE3693/FROM ;
  wire \CHOICE3693/GROM ;
  wire \CHOICE3754/FROM ;
  wire \CHOICE3754/GROM ;
  wire \DLX_EXinst_ALU_result<21>/FROM ;
  wire CHOICE4185;
  wire \CHOICE5400/FROM ;
  wire \CHOICE5400/GROM ;
  wire \CHOICE4879/FROM ;
  wire \CHOICE4879/GROM ;
  wire \DLX_IDinst_RegFile_7_4/FROM ;
  wire \DLX_IDinst_RegFile_7_4/GROM ;
  wire \CHOICE4114/FROM ;
  wire \CHOICE4114/GROM ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_196;
  wire \CHOICE4741/CYMUXF ;
  wire \CHOICE4741/GROM ;
  wire \CHOICE4741/CYINIT ;
  wire \N163672/FROM ;
  wire \N163672/GROM ;
  wire \DLX_IDinst_RegFile_1_9/FROM ;
  wire \DLX_IDinst_RegFile_1_9/GROM ;
  wire \CHOICE4918/FROM ;
  wire \CHOICE4918/GROM ;
  wire \CHOICE4116/FROM ;
  wire \CHOICE4116/GROM ;
  wire \DLX_EXinst_ALU_result<30>/FROM ;
  wire N162838;
  wire \CHOICE3699/FROM ;
  wire \CHOICE3699/GROM ;
  wire \CHOICE5797/FROM ;
  wire \CHOICE5797/GROM ;
  wire \DLX_EXinst_ALU_result<22>/FROM ;
  wire CHOICE4120;
  wire \CHOICE5474/FROM ;
  wire \CHOICE5474/GROM ;
  wire \CHOICE5096/FROM ;
  wire \CHOICE5096/GROM ;
  wire \N163518/FROM ;
  wire \N163518/GROM ;
  wire \DLX_IDinst_RegFile_15_7/FROM ;
  wire \DLX_IDinst_RegFile_15_7/GROM ;
  wire \N126777/FROM ;
  wire \N126777/GROM ;
  wire \CHOICE5441/FROM ;
  wire \CHOICE5441/GROM ;
  wire \CHOICE4914/FROM ;
  wire \CHOICE4914/GROM ;
  wire \CHOICE5801/FROM ;
  wire \CHOICE5801/GROM ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_100;
  wire \CHOICE5829/CYMUXF ;
  wire \CHOICE5829/GROM ;
  wire \CHOICE5829/CYINIT ;
  wire \CHOICE3977/FROM ;
  wire \CHOICE3977/GROM ;
  wire \N136886/FROM ;
  wire \N136886/GROM ;
  wire \DLX_IDinst_RegFile_3_11/FROM ;
  wire \DLX_IDinst_RegFile_3_11/GROM ;
  wire \N164729/FROM ;
  wire \N164729/GROM ;
  wire \CHOICE4587/FROM ;
  wire \CHOICE4587/GROM ;
  wire \DLX_EXinst_ALU_result<23>/FROM ;
  wire CHOICE4055;
  wire \DLX_IDinst_RegFile_22_8/FROM ;
  wire \DLX_IDinst_RegFile_22_8/GROM ;
  wire \DLX_EXinst_N76124/FROM ;
  wire \DLX_EXinst_N76124/GROM ;
  wire \CHOICE4592/FROM ;
  wire \CHOICE4592/GROM ;
  wire \CHOICE4545/FROM ;
  wire \CHOICE4545/GROM ;
  wire \DLX_IFinst_IR_previous<20>/FROM ;
  wire \DLX_IFinst_IR_previous<20>/GROM ;
  wire \DLX_IDinst_RegFile_2_19/FROM ;
  wire \DLX_IDinst_RegFile_2_19/GROM ;
  wire \DLX_IDinst_Mmux__COND_5_inst_lut4_584/FROM ;
  wire \DLX_IDinst_Mmux__COND_5_inst_lut4_584/GROM ;
  wire \DLX_IDinst_Mmux__COND_5_inst_lut4_582/FROM ;
  wire \DLX_IDinst_Mmux__COND_5_inst_lut4_582/GROM ;
  wire \DLX_IDinst_Mmux__COND_5_inst_lut4_578/FROM ;
  wire \DLX_IDinst_Mmux__COND_5_inst_lut4_578/GROM ;
  wire \DLX_IFinst_IR_previous<16>/FROM ;
  wire \DLX_IFinst_IR_previous<16>/GROM ;
  wire \DLX_IDinst_RegFile_2_27/FROM ;
  wire \DLX_IDinst_RegFile_2_27/GROM ;
  wire \DLX_IDinst_RegFile_18_11/FROM ;
  wire \DLX_IDinst_RegFile_18_11/GROM ;
  wire \DLX_IDinst_slot_num_FFd2/FROM ;
  wire \DLX_IDinst_slot_num_FFd2-In ;
  wire \DLX_IDinst_RegFile_15_16/FROM ;
  wire \DLX_IDinst_RegFile_15_16/GROM ;
  wire \DLX_IDinst_RegFile_26_5/FROM ;
  wire \DLX_IDinst_RegFile_26_5/GROM ;
  wire \DLX_IDinst_slot_num_FFd3-In ;
  wire \DLX_IDinst_slot_num_FFd3/GROM ;
  wire \DLX_IDinst_slot_num_FFd4/FROM ;
  wire \DLX_IDinst_slot_num_FFd4-In ;
  wire \DLX_IDinst_RegFile_2_21/FROM ;
  wire \DLX_IDinst_RegFile_2_21/GROM ;
  wire \DLX_EXinst_noop/FROM ;
  wire \DLX_EXinst_noop/GROM ;
  wire \DLX_EXinst_noop/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_2_13/FROM ;
  wire \DLX_IDinst_RegFile_2_13/GROM ;
  wire \DLX_IDinst_RegFile_1_1/FROM ;
  wire \DLX_IDinst_RegFile_1_1/GROM ;
  wire \DLX_IDinst_RegFile_11_21/FROM ;
  wire \DLX_IDinst_RegFile_11_21/GROM ;
  wire \DLX_IDinst_RegFile_2_22/FROM ;
  wire \DLX_IDinst_RegFile_2_22/GROM ;
  wire \DLX_IDinst_RegFile_15_5/FROM ;
  wire \DLX_IDinst_RegFile_15_5/GROM ;
  wire \DLX_IFinst_IR_previous<13>/FROM ;
  wire \DLX_IFinst_IR_previous<13>/GROM ;
  wire \DLX_EXinst_reg_out_B_EX<7>/FROM ;
  wire \DLX_EXinst_reg_out_B_EX<7>/GROM ;
  wire \DLX_IDinst_RegFile_2_23/FROM ;
  wire \DLX_IDinst_RegFile_2_23/GROM ;
  wire \DLX_IDinst_RegFile_2_15/FROM ;
  wire \DLX_IDinst_RegFile_2_15/GROM ;
  wire \DLX_IDinst_RegFile_0_12/FROM ;
  wire \DLX_IDinst_RegFile_0_12/GROM ;
  wire \DLX_IDinst_RegFile_23_30/FROM ;
  wire \DLX_IDinst_RegFile_23_30/GROM ;
  wire \DLX_IDinst_RegFile_2_24/FROM ;
  wire \DLX_IDinst_RegFile_2_24/GROM ;
  wire \DLX_IDinst_RegFile_2_16/FROM ;
  wire \DLX_IDinst_RegFile_2_16/GROM ;
  wire \DLX_IDinst_RegFile_16_15/FROM ;
  wire \DLX_IDinst_RegFile_16_15/GROM ;
  wire \DLX_IDinst_RegFile_2_17/FROM ;
  wire \DLX_IDinst_RegFile_2_17/GROM ;
  wire \DLX_IDinst_RegFile_22_6/FROM ;
  wire \DLX_IDinst_RegFile_22_6/GROM ;
  wire \DLX_IDinst_RegFile_1_23/FROM ;
  wire \DLX_IDinst_RegFile_1_23/GROM ;
  wire \DLX_MEMinst_opcode_of_WB<5>/FROM ;
  wire \DLX_MEMinst_opcode_of_WB<5>/GROM ;
  wire \DLX_IDinst_RegFile_11_24/FROM ;
  wire \DLX_IDinst_RegFile_11_24/GROM ;
  wire \DLX_IDinst_RegFile_6_6/FROM ;
  wire \DLX_IDinst_RegFile_6_6/GROM ;
  wire \DLX_IFinst_PC<28>/FROM ;
  wire \DLX_IFinst_PC<28>/GROM ;
  wire \DLX_IDinst_RegFile_15_9/FROM ;
  wire \DLX_IDinst_RegFile_15_9/GROM ;
  wire \DLX_IDinst_RegFile_1_26/FROM ;
  wire \DLX_IDinst_RegFile_1_26/GROM ;
  wire \DLX_IFinst_IR_previous<6>/FROM ;
  wire \DLX_IFinst_IR_previous<6>/GROM ;
  wire \DLX_IDinst_RegFile_26_2/FROM ;
  wire \DLX_IDinst_RegFile_26_2/GROM ;
  wire \DLX_IDinst_RegFile_22_13/FROM ;
  wire \DLX_IDinst_RegFile_22_13/GROM ;
  wire \DLX_IDinst_RegFile_30_23/FROM ;
  wire \DLX_IDinst_RegFile_30_23/GROM ;
  wire \DLX_IDinst_RegFile_3_13/FROM ;
  wire \DLX_IDinst_RegFile_3_13/GROM ;
  wire \DLX_IDinst_RegFile_3_21/FROM ;
  wire \DLX_IDinst_RegFile_3_21/GROM ;
  wire \DLX_IDinst_RegFile_2_29/FROM ;
  wire \DLX_IDinst_RegFile_2_29/GROM ;
  wire \DLX_IDinst_RegFile_23_23/FROM ;
  wire \DLX_IDinst_RegFile_23_23/GROM ;
  wire \DLX_IDinst_RegFile_3_22/FROM ;
  wire \DLX_IDinst_RegFile_3_22/GROM ;
  wire \DLX_IDinst_RegFile_23_17/FROM ;
  wire \DLX_IDinst_RegFile_23_17/GROM ;
  wire \DLX_IDinst_RegFile_18_4/FROM ;
  wire \DLX_IDinst_RegFile_18_4/GROM ;
  wire \DLX_IDinst_RegFile_3_15/FROM ;
  wire \DLX_IDinst_RegFile_3_15/GROM ;
  wire \DLX_IDinst_RegFile_17_18/FROM ;
  wire \DLX_IDinst_RegFile_17_18/GROM ;
  wire \DLX_IDinst_RegFile_3_31/FROM ;
  wire \DLX_IDinst_RegFile_3_31/GROM ;
  wire \DLX_IDinst_RegFile_29_7/FROM ;
  wire \DLX_IDinst_RegFile_29_7/GROM ;
  wire \DLX_IDinst_RegFile_1_0/FROM ;
  wire \DLX_IDinst_RegFile_1_0/GROM ;
  wire \DLX_IDinst_RegFile_3_24/FROM ;
  wire \DLX_IDinst_RegFile_3_24/GROM ;
  wire \DLX_IDinst_RegFile_3_17/FROM ;
  wire \DLX_IDinst_RegFile_3_17/GROM ;
  wire \DLX_IDinst_RegFile_3_25/FROM ;
  wire \DLX_IDinst_RegFile_3_25/GROM ;
  wire \CHOICE2324/FROM ;
  wire \CHOICE2324/GROM ;
  wire \CHOICE2445/FROM ;
  wire \CHOICE2445/GROM ;
  wire \DLX_EXinst__n0013<10>/FROM ;
  wire \DLX_EXinst__n0013<10>/GROM ;
  wire \CHOICE5771/FROM ;
  wire \CHOICE5771/GROM ;
  wire \CHOICE2335/FROM ;
  wire \CHOICE2335/GROM ;
  wire \CHOICE2434/FROM ;
  wire \CHOICE2434/GROM ;
  wire \CHOICE2346/FROM ;
  wire \CHOICE2346/GROM ;
  wire \CHOICE5511/FROM ;
  wire \CHOICE5511/GROM ;
  wire \DLX_IDinst_regA_eff<28>/FROM ;
  wire \DLX_IDinst_regA_eff<28>/GROM ;
  wire \CHOICE2401/FROM ;
  wire \CHOICE2401/GROM ;
  wire \CHOICE5435/FROM ;
  wire \CHOICE5435/GROM ;
  wire \N164108/FROM ;
  wire \N164108/GROM ;
  wire \N127166/FROM ;
  wire \N127166/GROM ;
  wire \DLX_EXinst_Mshift__n0024_Sh<30>/FROM ;
  wire \DLX_EXinst_Mshift__n0024_Sh<30>/GROM ;
  wire \DLX_EXinst_Mshift__n0024_Sh<31>/FROM ;
  wire \DLX_EXinst_Mshift__n0024_Sh<31>/GROM ;
  wire \DLX_EXinst_Mshift__n0024_Sh<51>/FROM ;
  wire \DLX_EXinst_Mshift__n0024_Sh<51>/GROM ;
  wire \N132499/FROM ;
  wire \N132499/GROM ;
  wire \N136799/FROM ;
  wire \N136799/GROM ;
  wire \CHOICE2040/FROM ;
  wire \CHOICE2040/GROM ;
  wire \DLX_IDinst_RegFile_3_20/FROM ;
  wire \DLX_IDinst_RegFile_3_20/GROM ;
  wire \DLX_EXinst_N74441/FROM ;
  wire \DLX_EXinst_N74441/GROM ;
  wire \N164125/FROM ;
  wire \N164125/GROM ;
  wire \DLX_IDinst_RegFile_18_1/FROM ;
  wire \DLX_IDinst_RegFile_18_1/GROM ;
  wire \N164115/FROM ;
  wire \N164115/GROM ;
  wire \DLX_IFinst_IR_previous<19>/FROM ;
  wire \DLX_IFinst_IR_previous<19>/GROM ;
  wire \DLX_MEMinst_reg_write_MEM/FROM ;
  wire \DLX_MEMinst_reg_write_MEM/GROM ;
  wire \DLX_IDinst_RegFile_14_23/FROM ;
  wire \DLX_IDinst_RegFile_14_23/GROM ;
  wire \CHOICE5824/FROM ;
  wire \CHOICE5824/GROM ;
  wire \DLX_IDinst_branch_sig/FROM ;
  wire \DLX_IDinst_branch_sig/GROM ;
  wire \N163128/FROM ;
  wire \N163128/GROM ;
  wire \DLX_IDinst_Imm<31>/FROM ;
  wire \DLX_IDinst_Imm<31>/GROM ;
  wire \DLX_IDinst_RegFile_10_6/FROM ;
  wire \DLX_IDinst_RegFile_10_6/GROM ;
  wire \N163842/FROM ;
  wire \N163842/GROM ;
  wire \DLX_IDinst_RegFile_11_2/FROM ;
  wire \DLX_IDinst_RegFile_11_2/GROM ;
  wire \CHOICE3508/FROM ;
  wire \CHOICE3508/GROM ;
  wire \CHOICE3547/FROM ;
  wire \CHOICE3547/GROM ;
  wire \N164734/FROM ;
  wire \N164734/GROM ;
  wire \N136586/FROM ;
  wire \N136586/GROM ;
  wire \CHOICE3524/FROM ;
  wire \CHOICE3524/GROM ;
  wire \DLX_IDinst_RegFile_1_5/FROM ;
  wire \DLX_IDinst_RegFile_1_5/GROM ;
  wire \DLX_IDinst__n0164/FROM ;
  wire \DLX_IDinst__n0164/GROM ;
  wire \DLX_IDinst_RegFile_22_11/FROM ;
  wire \DLX_IDinst_RegFile_22_11/GROM ;
  wire \DLX_IDinst_stall/FROM ;
  wire \DLX_IDinst_stall/GROM ;
  wire \N163733/FROM ;
  wire \N163733/GROM ;
  wire \N163574/FROM ;
  wire \N163574/GROM ;
  wire \DLX_IFinst_IR_curr<28>/FROM ;
  wire \DLX_IFinst_IR_curr<28>/GROM ;
  wire \CHOICE1971/FROM ;
  wire \CHOICE1971/GROM ;
  wire \CHOICE4208/FROM ;
  wire \CHOICE4208/GROM ;
  wire \N131907/FROM ;
  wire \N131907/GROM ;
  wire \CHOICE1338/FROM ;
  wire \CHOICE1338/GROM ;
  wire N162964;
  wire \DLX_IDinst_reg_out_A<30>/GROM ;
  wire \CHOICE2148/FROM ;
  wire \CHOICE2148/GROM ;
  wire \DLX_IFinst_IR_curr<29>/FROM ;
  wire \DLX_IFinst_IR_curr<29>/GROM ;
  wire \CHOICE2170/FROM ;
  wire \CHOICE2170/GROM ;
  wire \DLX_IDinst_reg_out_B<0>/FROM ;
  wire \CHOICE2181/FROM ;
  wire \CHOICE2181/GROM ;
  wire \DLX_IDinst_slot_num_FFd1-In ;
  wire \DLX_IDinst_slot_num_FFd1/GROM ;
  wire \CHOICE2192/FROM ;
  wire \CHOICE2192/GROM ;
  wire \N163652/FROM ;
  wire \N163652/GROM ;
  wire \DLX_IDinst_RegFile_3_19/FROM ;
  wire \DLX_IDinst_RegFile_3_19/GROM ;
  wire \CHOICE2224/FROM ;
  wire \CHOICE2224/GROM ;
  wire \DLX_IDinst_N107837/FROM ;
  wire \DLX_IDinst_N107837/GROM ;
  wire \CHOICE5058/FROM ;
  wire \CHOICE5058/GROM ;
  wire \DLX_IDinst_RegFile_2_5/FROM ;
  wire \DLX_IDinst_RegFile_2_5/GROM ;
  wire \DLX_EXinst__n0054/FROM ;
  wire \DLX_EXinst__n0054/GROM ;
  wire \CHOICE5713/FROM ;
  wire \CHOICE5713/GROM ;
  wire \CHOICE4924/FROM ;
  wire \CHOICE4924/GROM ;
  wire \DLX_IDinst_RegFile_27_25/FROM ;
  wire \DLX_IDinst_RegFile_27_25/GROM ;
  wire \CHOICE5458/FROM ;
  wire \CHOICE5458/GROM ;
  wire \DLX_EXinst__n0052/FROM ;
  wire \DLX_EXinst__n0052/GROM ;
  wire \CHOICE4661/FROM ;
  wire \CHOICE4661/GROM ;
  wire \DLX_IDinst_RegFile_3_1/FROM ;
  wire \DLX_IDinst_RegFile_3_1/GROM ;
  wire \N163606/FROM ;
  wire \N163606/GROM ;
  wire \CHOICE4688/FROM ;
  wire \CHOICE4688/GROM ;
  wire \DLX_EXinst_ALU_result<20>/FROM ;
  wire N162820;
  wire \DLX_IDinst_RegFile_3_27/FROM ;
  wire \DLX_IDinst_RegFile_3_27/GROM ;
  wire \CHOICE4634/FROM ;
  wire \CHOICE4634/GROM ;
  wire \N163481/FROM ;
  wire \N163481/GROM ;
  wire \DLX_IDinst_RegFile_23_8/FROM ;
  wire \DLX_IDinst_RegFile_23_8/GROM ;
  wire \N131375/FROM ;
  wire \N131375/GROM ;
  wire \DLX_EXinst_ALU_result<16>/FROM ;
  wire CHOICE4629;
  wire \CHOICE5622/FROM ;
  wire \CHOICE5622/GROM ;
  wire \DLX_IDinst_RegFile_7_3/FROM ;
  wire \DLX_IDinst_RegFile_7_3/GROM ;
  wire \CHOICE5677/FROM ;
  wire \CHOICE5677/GROM ;
  wire \CHOICE4850/FROM ;
  wire \CHOICE4850/GROM ;
  wire \CHOICE5383/FROM ;
  wire \CHOICE5383/GROM ;
  wire \DLX_IDinst_RegFile_22_16/FROM ;
  wire \DLX_IDinst_RegFile_22_16/GROM ;
  wire \N164155/FROM ;
  wire \N164155/GROM ;
  wire \DLX_EXinst_ALU_result<24>/FROM ;
  wire CHOICE5683;
  wire \N163522/FROM ;
  wire \N163522/GROM ;
  wire \DLX_IDinst_RegFile_2_7/FROM ;
  wire \DLX_IDinst_RegFile_2_7/GROM ;
  wire \CHOICE5225/FROM ;
  wire \CHOICE5225/GROM ;
  wire \DLX_EXinst_ALU_result<25>/FROM ;
  wire CHOICE5120;
  wire \N163593/FROM ;
  wire \N163593/GROM ;
  wire \DLX_EXinst_ALU_result<17>/FROM ;
  wire CHOICE5428;
  wire \CHOICE4962/FROM ;
  wire \CHOICE4962/GROM ;
  wire \CHOICE5421/FROM ;
  wire \CHOICE5421/GROM ;
  wire \CHOICE5321/FROM ;
  wire \CHOICE5321/GROM ;
  wire \DLX_IDinst_RegFile_3_4/FROM ;
  wire \DLX_IDinst_RegFile_3_4/GROM ;
  wire \CHOICE5049/FROM ;
  wire \CHOICE5049/GROM ;
  wire \CHOICE5304/FROM ;
  wire \CHOICE5304/GROM ;
  wire \DLX_EXinst_ALU_result<26>/FROM ;
  wire CHOICE5053;
  wire \N163294/FROM ;
  wire \N163294/GROM ;
  wire \DLX_EXinst_ALU_result<18>/FROM ;
  wire CHOICE5270;
  wire \CHOICE5263/FROM ;
  wire \CHOICE5263/GROM ;
  wire \CHOICE5307/FROM ;
  wire \CHOICE5307/GROM ;
  wire \CHOICE5345/FROM ;
  wire \CHOICE5345/GROM ;
  wire \N163412/FROM ;
  wire \N163412/GROM ;
  wire \CHOICE4982/FROM ;
  wire \CHOICE4982/GROM ;
  wire \N130467/FROM ;
  wire \N130467/GROM ;
  wire \CHOICE4910/FROM ;
  wire \CHOICE4910/GROM ;
  wire \DLX_EXinst_ALU_result<27>/FROM ;
  wire CHOICE4986;
  wire \DLX_EXinst_ALU_result<19>/FROM ;
  wire CHOICE5349;
  wire \N163684/FROM ;
  wire \N163684/GROM ;
  wire \CHOICE4801/GROM ;
  wire \DLX_EXinst_ALU_result<28>/FROM ;
  wire N162804;
  wire \DLX_EXinst_Mshift__n0019_Sh<12>/FROM ;
  wire \DLX_EXinst_Mshift__n0019_Sh<12>/GROM ;
  wire \CHOICE3939/FROM ;
  wire \CHOICE3939/GROM ;
  wire \DLX_EXinst_N76382/FROM ;
  wire \DLX_EXinst_N76382/GROM ;
  wire \DLX_IDinst_RegFile_1_17/FROM ;
  wire \DLX_IDinst_RegFile_1_17/GROM ;
  wire \CHOICE3711/FROM ;
  wire \CHOICE3711/GROM ;
  wire \DLX_EXinst_Mshift__n0019_Sh<30>/FROM ;
  wire \DLX_EXinst_Mshift__n0019_Sh<30>/GROM ;
  wire \CHOICE4833/FROM ;
  wire \CHOICE4833/GROM ;
  wire \DLX_EXinst_ALU_result<29>/FROM ;
  wire N162835;
  wire \CHOICE5550/FROM ;
  wire \CHOICE5550/GROM ;
  wire \DLX_EXinst_Mshift__n0019_Sh<16>/FROM ;
  wire \DLX_EXinst_Mshift__n0019_Sh<16>/GROM ;
  wire \N163148/FROM ;
  wire \N163148/GROM ;
  wire \DLX_IDinst_RegFile_27_29/FROM ;
  wire \DLX_IDinst_RegFile_27_29/GROM ;
  wire \DLX_EXinst_Mshift__n0019_Sh<18>/FROM ;
  wire \DLX_EXinst_Mshift__n0019_Sh<18>/GROM ;
  wire \DLX_EXinst_Mshift__n0019_Sh<19>/FROM ;
  wire \DLX_EXinst_Mshift__n0019_Sh<19>/GROM ;
  wire \DLX_EXinst_Mshift__n0019_Sh<61>/FROM ;
  wire \DLX_EXinst_Mshift__n0019_Sh<61>/GROM ;
  wire \DLX_IDinst_EPC<6>/FROM ;
  wire \DLX_IDinst_EPC<6>/GROM ;
  wire \DLX_EXinst__n0036/FROM ;
  wire \DLX_EXinst__n0036/GROM ;
  wire \DLX_EXinst_Mshift__n0019_Sh<88>/FROM ;
  wire \DLX_EXinst_Mshift__n0019_Sh<88>/GROM ;
  wire \red_1_OBUF/FROM ;
  wire \red_1_OBUF/GROM ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_61;
  wire \DLX_IDinst_RegFile_4_0/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_62;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_2;
  wire \DLX_IDinst_RegFile_4_0/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_4_0/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_77;
  wire \DLX_IDinst_RegFile_4_1/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_78;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_18;
  wire \DLX_IDinst_RegFile_4_1/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_4_1/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_93;
  wire \DLX_IDinst_RegFile_4_2/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_94;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_34;
  wire \DLX_IDinst_RegFile_4_2/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_4_2/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_109;
  wire \DLX_IDinst_RegFile_4_3/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_110;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_50;
  wire \DLX_IDinst_RegFile_4_3/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_4_3/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_125;
  wire \DLX_IDinst_RegFile_4_4/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_126;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_66;
  wire \DLX_IDinst_RegFile_4_4/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_4_4/CYINIT ;
  wire \DLX_IFinst_IR_previous<30>/FROM ;
  wire \DLX_IFinst_IR_previous<30>/GROM ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_589;
  wire \DLX_IDinst_RegFile_5_0/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_590;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_514;
  wire \DLX_IDinst_RegFile_5_0/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_5_0/CYINIT ;
  wire \DLX_IFinst_NPC<0>/FROM ;
  wire \DLX_IFinst_NPC<0>/GROM ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_141;
  wire \DLX_IDinst_RegFile_4_5/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_142;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_82;
  wire \DLX_IDinst_RegFile_4_5/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_4_5/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_605;
  wire \DLX_IDinst_RegFile_5_1/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_606;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_530;
  wire \DLX_IDinst_RegFile_5_1/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_5_1/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_157;
  wire \DLX_IDinst_RegFile_4_6/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_158;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_98;
  wire \DLX_IDinst_RegFile_4_6/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_4_6/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_621;
  wire \DLX_IDinst_RegFile_5_2/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_622;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_546;
  wire \DLX_IDinst_RegFile_5_2/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_5_2/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_173;
  wire \DLX_IDinst_RegFile_4_7/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_174;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_114;
  wire \DLX_IDinst_RegFile_4_7/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_4_7/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_637;
  wire \DLX_IDinst_RegFile_5_3/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_638;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_562;
  wire \DLX_IDinst_RegFile_5_3/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_5_3/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_189;
  wire \DLX_IDinst_RegFile_4_8/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_190;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_130;
  wire \DLX_IDinst_RegFile_4_8/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_4_8/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_653;
  wire \DLX_IDinst_RegFile_5_4/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_654;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_578;
  wire \DLX_IDinst_RegFile_5_4/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_5_4/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_205;
  wire \DLX_IDinst_RegFile_4_9/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_206;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_146;
  wire \DLX_IDinst_RegFile_4_9/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_4_9/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_669;
  wire \DLX_IDinst_RegFile_5_5/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_670;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_594;
  wire \DLX_IDinst_RegFile_5_5/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_5_5/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_685;
  wire \DLX_IDinst_RegFile_5_6/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_686;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_610;
  wire \DLX_IDinst_RegFile_5_6/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_5_6/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_701;
  wire \DLX_IDinst_RegFile_5_7/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_702;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_626;
  wire \DLX_IDinst_RegFile_5_7/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_5_7/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_717;
  wire \DLX_IDinst_RegFile_5_8/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_718;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_642;
  wire \DLX_IDinst_RegFile_5_8/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_5_8/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_733;
  wire \DLX_IDinst_RegFile_5_9/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_734;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_658;
  wire \DLX_IDinst_RegFile_5_9/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_5_9/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_63;
  wire \DLX_IDinst_RegFile_8_0/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_64;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_4;
  wire \DLX_IDinst_RegFile_8_0/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_8_0/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_79;
  wire \DLX_IDinst_RegFile_8_1/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_80;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_20;
  wire \DLX_IDinst_RegFile_8_1/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_8_1/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_95;
  wire \DLX_IDinst_RegFile_8_2/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_96;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_36;
  wire \DLX_IDinst_RegFile_8_2/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_8_2/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_111;
  wire \DLX_IDinst_RegFile_8_3/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_112;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_52;
  wire \DLX_IDinst_RegFile_8_3/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_8_3/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_127;
  wire \DLX_IDinst_RegFile_8_4/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_128;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_68;
  wire \DLX_IDinst_RegFile_8_4/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_8_4/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_591;
  wire \DLX_IDinst_RegFile_9_0/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_592;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_516;
  wire \DLX_IDinst_RegFile_9_0/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_9_0/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_143;
  wire \DLX_IDinst_RegFile_8_5/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_144;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_84;
  wire \DLX_IDinst_RegFile_8_5/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_8_5/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_607;
  wire \DLX_IDinst_RegFile_9_1/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_608;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_532;
  wire \DLX_IDinst_RegFile_9_1/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_9_1/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_159;
  wire \DLX_IDinst_RegFile_8_6/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_160;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_100;
  wire \DLX_IDinst_RegFile_8_6/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_8_6/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_623;
  wire \DLX_IDinst_RegFile_9_2/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_624;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_548;
  wire \DLX_IDinst_RegFile_9_2/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_9_2/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_175;
  wire \DLX_IDinst_RegFile_8_7/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_176;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_116;
  wire \DLX_IDinst_RegFile_8_7/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_8_7/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_639;
  wire \DLX_IDinst_RegFile_9_3/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_640;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_564;
  wire \DLX_IDinst_RegFile_9_3/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_9_3/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_191;
  wire \DLX_IDinst_RegFile_8_8/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_192;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_132;
  wire \DLX_IDinst_RegFile_8_8/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_8_8/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_655;
  wire \DLX_IDinst_RegFile_9_4/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_656;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_580;
  wire \DLX_IDinst_RegFile_9_4/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_9_4/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_207;
  wire \DLX_IDinst_RegFile_8_9/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_208;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_148;
  wire \DLX_IDinst_RegFile_8_9/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_8_9/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_671;
  wire \DLX_IDinst_RegFile_9_5/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_672;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_596;
  wire \DLX_IDinst_RegFile_9_5/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_9_5/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_687;
  wire \DLX_IDinst_RegFile_9_6/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_688;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_612;
  wire \DLX_IDinst_RegFile_9_6/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_9_6/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_703;
  wire \DLX_IDinst_RegFile_9_7/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_704;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_628;
  wire \DLX_IDinst_RegFile_9_7/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_9_7/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_719;
  wire \DLX_IDinst_RegFile_9_8/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_720;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_644;
  wire \DLX_IDinst_RegFile_9_8/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_9_8/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_735;
  wire \DLX_IDinst_RegFile_9_9/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_736;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_660;
  wire \DLX_IDinst_RegFile_9_9/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_9_9/CYINIT ;
  wire \DLX_IFinst_NPC<1>/FROM ;
  wire \DLX_IFinst_NPC<1>/GROM ;
  wire \DLX_IFinst_NPC<2>/FROM ;
  wire \DLX_IFinst_NPC<2>/GROM ;
  wire \N164184/FROM ;
  wire \N164184/GROM ;
  wire \DLX_IFinst_NPC<3>/FROM ;
  wire \DLX_IFinst_NPC<3>/GROM ;
  wire \DLX_IFinst_NPC<4>/FROM ;
  wire \DLX_IFinst_NPC<4>/GROM ;
  wire \DLX_IFinst_NPC<5>/FROM ;
  wire \DLX_IFinst_NPC<5>/GROM ;
  wire \DLX_IFinst_NPC<6>/FROM ;
  wire \DLX_IFinst_NPC<6>/GROM ;
  wire \DLX_IFinst_NPC<7>/FROM ;
  wire \DLX_IFinst_NPC<7>/GROM ;
  wire \DLX_IFinst_NPC<8>/FROM ;
  wire \DLX_IFinst_NPC<8>/GROM ;
  wire \DLX_IFinst_NPC<9>/FROM ;
  wire \DLX_IFinst_NPC<9>/GROM ;
  wire \DLX_IFinst_IR_curr<7>/FROM ;
  wire \DLX_IFinst_IR_curr<7>/GROM ;
  wire \DLX_IDinst_RegFile_11_10/FROM ;
  wire \DLX_IDinst_RegFile_11_10/GROM ;
  wire \DLX_IDinst_RegFile_11_14/FROM ;
  wire \DLX_IDinst_RegFile_11_14/GROM ;
  wire \DLX_IDinst_RegFile_11_26/FROM ;
  wire \DLX_IDinst_RegFile_11_26/GROM ;
  wire \DLX_IDinst_RegFile_11_28/FROM ;
  wire \DLX_IDinst_RegFile_11_28/GROM ;
  wire \DLX_IDinst_RegFile_7_2/FROM ;
  wire \DLX_IDinst_RegFile_7_2/GROM ;
  wire \DLX_IDinst_RegFile_2_0/FROM ;
  wire \DLX_IDinst_RegFile_2_0/GROM ;
  wire \DLX_IDinst_EPC<2>/FROM ;
  wire \DLX_IDinst_EPC<2>/GROM ;
  wire \DLX_IDinst_EPC<3>/FROM ;
  wire \DLX_IDinst_EPC<3>/GROM ;
  wire \DLX_IDinst_EPC<4>/FROM ;
  wire \DLX_IDinst_EPC<4>/GROM ;
  wire \DLX_IDinst_EPC<5>/FROM ;
  wire \DLX_IDinst_EPC<5>/GROM ;
  wire \DLX_IFinst_PC<10>/FROM ;
  wire \DLX_IFinst_PC<10>/GROM ;
  wire \DLX_IDinst_RegFile_11_4/FROM ;
  wire \DLX_IDinst_RegFile_11_4/GROM ;
  wire \DLX_IDinst_RegFile_6_23/FROM ;
  wire \DLX_IDinst_RegFile_6_23/GROM ;
  wire \DLX_IDinst_RegFile_6_16/FROM ;
  wire \DLX_IDinst_RegFile_6_16/GROM ;
  wire \N164583/FROM ;
  wire \N164583/GROM ;
  wire \DLX_IDinst_RegFile_6_19/FROM ;
  wire \DLX_IDinst_RegFile_6_19/GROM ;
  wire \CHOICE4779/FROM ;
  wire \CHOICE4779/GROM ;
  wire \CHOICE3133/FROM ;
  wire \CHOICE3133/GROM ;
  wire \CHOICE4991/FROM ;
  wire \CHOICE4991/GROM ;
  wire \CHOICE4539/FROM ;
  wire \CHOICE4539/GROM ;
  wire \CHOICE5447/FROM ;
  wire \CHOICE5447/GROM ;
  wire \CHOICE5170/FROM ;
  wire \CHOICE5170/GROM ;
  wire \N131693/FROM ;
  wire \N131693/GROM ;
  wire \CHOICE5455/FROM ;
  wire \CHOICE5455/GROM ;
  wire \CHOICE4716/FROM ;
  wire \CHOICE4716/GROM ;
  wire \CHOICE5715/FROM ;
  wire \CHOICE5715/GROM ;
  wire \N163704/FROM ;
  wire \N163704/GROM ;
  wire \N163931/FROM ;
  wire \N163931/GROM ;
  wire \CHOICE4330/FROM ;
  wire \CHOICE4330/GROM ;
  wire \CHOICE5186/FROM ;
  wire \CHOICE5186/GROM ;
  wire \CHOICE2058/FROM ;
  wire \CHOICE2058/GROM ;
  wire \CHOICE5536/FROM ;
  wire \CHOICE5536/GROM ;
  wire \CHOICE3718/FROM ;
  wire \CHOICE3718/GROM ;
  wire \CHOICE5460/FROM ;
  wire \CHOICE5460/GROM ;
  wire \CHOICE4519/FROM ;
  wire \CHOICE4519/GROM ;
  wire \CHOICE3889/FROM ;
  wire \CHOICE3889/GROM ;
  wire \CHOICE4273/FROM ;
  wire \CHOICE4273/GROM ;
  wire \CHOICE5127/FROM ;
  wire \CHOICE5127/GROM ;
  wire \CHOICE5139/FROM ;
  wire \CHOICE5139/GROM ;
  wire \CHOICE3773/FROM ;
  wire \CHOICE3773/GROM ;
  wire \CHOICE5724/FROM ;
  wire \CHOICE5724/GROM ;
  wire \DLX_EXinst_N76479/FROM ;
  wire \DLX_EXinst_N76479/GROM ;
  wire \CHOICE5732/FROM ;
  wire \CHOICE5732/GROM ;
  wire \CHOICE3656/FROM ;
  wire \CHOICE3656/GROM ;
  wire \CHOICE4263/FROM ;
  wire \CHOICE4263/GROM ;
  wire \CHOICE5477/FROM ;
  wire \CHOICE5477/GROM ;
  wire \vga_top_vga1_helpme/GROM ;
  wire \vga_top_vga1_helpme/LOGIC_ZERO ;
  wire \N163728/FROM ;
  wire \N163728/GROM ;
  wire \N164228/FROM ;
  wire \N164228/GROM ;
  wire \N163979/FROM ;
  wire \N163979/GROM ;
  wire \N163286/FROM ;
  wire \N163286/GROM ;
  wire \reset_IBUF_14/FROM ;
  wire \reset_IBUF_14/GROM ;
  wire \reset_IBUF_13/FROM ;
  wire \reset_IBUF_13/GROM ;
  wire \reset_IBUF_9/FROM ;
  wire \reset_IBUF_9/GROM ;
  wire \DLX_IDinst_Cause_Reg<0>/GROM ;
  wire \DLX_IDinst_Cause_Reg<1>/FROM ;
  wire \DLX_IDinst_Cause_Reg<1>/GROM ;
  wire \DLX_IDinst_Cause_Reg<2>/FROM ;
  wire \DLX_IDinst_Cause_Reg<2>/GROM ;
  wire \DLX_IDinst_Cause_Reg<3>/FROM ;
  wire \DLX_IDinst_Cause_Reg<3>/GROM ;
  wire \DLX_IDinst_Cause_Reg<4>/FROM ;
  wire \DLX_IDinst_Cause_Reg<4>/GROM ;
  wire \DLX_IDinst_Cause_Reg<5>/FROM ;
  wire \DLX_IDinst_Cause_Reg<5>/GROM ;
  wire \DLX_IDinst_Cause_Reg<7>/FROM ;
  wire \DLX_IDinst_Cause_Reg<7>/GROM ;
  wire \DLX_IDinst_Cause_Reg<8>/FROM ;
  wire \DLX_IDinst_Cause_Reg<8>/GROM ;
  wire \DLX_IDinst_Cause_Reg<9>/FROM ;
  wire \DLX_IDinst_Cause_Reg<9>/GROM ;
  wire \CHOICE5181/FROM ;
  wire \CHOICE5181/GROM ;
  wire \CHOICE1994/FROM ;
  wire \CHOICE1994/GROM ;
  wire \DLX_IDinst_delay_slot/FROM ;
  wire N146881;
  wire \N163420/FROM ;
  wire \N163420/GROM ;
  wire \DLX_IDinst_reg_dst/FROM ;
  wire N147993;
  wire \CHOICE3558/FROM ;
  wire \CHOICE3558/GROM ;
  wire \DLX_IDinst_reg_write/FROM ;
  wire N148197;
  wire \CHOICE4224/FROM ;
  wire \CHOICE4224/GROM ;
  wire \CHOICE4256/FROM ;
  wire \CHOICE4256/GROM ;
  wire \DLX_IDinst_zflag/FROM ;
  wire \DLX_IDinst_zflag/GROM ;
  wire \N138903/FROM ;
  wire \N138903/GROM ;
  wire \DLX_IDinst_N107223/FROM ;
  wire \DLX_IDinst_N107223/GROM ;
  wire \N163416/FROM ;
  wire \N163416/GROM ;
  wire \DLX_IFinst_NPC<10>/FROM ;
  wire \DLX_IFinst_NPC<10>/GROM ;
  wire \DLX_IDinst_N108305/FROM ;
  wire \DLX_IDinst_N108305/GROM ;
  wire \N164614/FROM ;
  wire \N164614/GROM ;
  wire \DLX_IDinst_N108244/FROM ;
  wire \DLX_IDinst_N108244/GROM ;
  wire \DLX_IDinst_N107452/FROM ;
  wire \DLX_IDinst_N107452/GROM ;
  wire \DLX_IDinst_N108221/FROM ;
  wire \DLX_IDinst_N108221/GROM ;
  wire \DLX_IDinst_N108165/FROM ;
  wire \DLX_IDinst_N108165/GROM ;
  wire \DLX_IDinst_N108238/FROM ;
  wire \DLX_IDinst_N108238/GROM ;
  wire \N163258/GROM ;
  wire \DLX_IDinst_N107623/FROM ;
  wire \DLX_IDinst_N107623/GROM ;
  wire \DLX_IDinst_N108503/FROM ;
  wire \DLX_IDinst_N108503/GROM ;
  wire \DLX_IDinst_N108264/FROM ;
  wire \DLX_IDinst_N108264/GROM ;
  wire \DLX_IDinst_N108249/FROM ;
  wire \DLX_IDinst_N108249/GROM ;
  wire \DLX_IDinst_N108100/FROM ;
  wire \DLX_IDinst_N108100/GROM ;
  wire \DLX_IDinst_N108517/FROM ;
  wire \DLX_IDinst_N108517/GROM ;
  wire \DLX_IFinst_NPC<11>/FROM ;
  wire \DLX_IFinst_NPC<11>/GROM ;
  wire \DLX_IDinst_N108552/FROM ;
  wire \DLX_IDinst_N108552/GROM ;
  wire \N164200/FROM ;
  wire \N164200/GROM ;
  wire \CHOICE1319/FROM ;
  wire \CHOICE1319/GROM ;
  wire \DLX_IDinst_N108574/FROM ;
  wire \DLX_IDinst_N108574/GROM ;
  wire \DLX_IDinst_N108559/FROM ;
  wire \DLX_IDinst_N108559/GROM ;
  wire \DLX_IFinst_NPC<20>/FROM ;
  wire \DLX_IFinst_NPC<12>/FROM ;
  wire \DLX_IFinst_NPC<12>/GROM ;
  wire \N164620/FROM ;
  wire \N164620/GROM ;
  wire \DLX_IFinst_NPC<21>/FROM ;
  wire \DLX_IFinst_NPC<13>/FROM ;
  wire \DLX_IFinst_NPC<13>/GROM ;
  wire \DLX_IDinst_branch_address<10>/FROM ;
  wire N140319;
  wire \DLX_IDinst_branch_address<11>/FROM ;
  wire N140382;
  wire \DLX_IDinst_RegFile_2_12/FROM ;
  wire \DLX_IDinst_RegFile_2_12/GROM ;
  wire \DLX_IDinst_branch_address<20>/FROM ;
  wire N141013;
  wire \DLX_IDinst_branch_address<12>/FROM ;
  wire N140445;
  wire \DLX_IDinst_branch_address<13>/FROM ;
  wire N140508;
  wire \DLX_IDinst_branch_address<21>/FROM ;
  wire N141076;
  wire \DLX_IFinst_NPC<30>/FROM ;
  wire \DLX_IFinst_NPC<14>/FROM ;
  wire \DLX_IFinst_NPC<14>/GROM ;
  wire \DLX_IFinst_NPC<22>/FROM ;
  wire \DLX_IDinst_branch_address<22>/FROM ;
  wire N141139;
  wire \DLX_IDinst_branch_address<14>/FROM ;
  wire N140571;
  wire \DLX_IDinst_branch_address<30>/FROM ;
  wire N141202;
  wire \DLX_IDinst_branch_address<15>/FROM ;
  wire N140634;
  wire \DLX_IDinst_branch_address<23>/FROM ;
  wire N141643;
  wire \CHOICE3164/FROM ;
  wire \CHOICE3164/GROM ;
  wire \DLX_IDinst_branch_address<31>/FROM ;
  wire N145908;
  wire \CHOICE2213/FROM ;
  wire \CHOICE2213/GROM ;
  wire \DLX_IDinst_RegFile_3_29/FROM ;
  wire \DLX_IDinst_RegFile_3_29/GROM ;
  wire \DLX_EXinst_ALU_result<0>/FROM ;
  wire \DLX_EXinst_ALU_result<0>/GROM ;
  wire \DLX_IDinst_branch_address<16>/FROM ;
  wire N140761;
  wire \DLX_IDinst_branch_address<24>/FROM ;
  wire N141580;
  wire \DLX_IDinst_branch_address<25>/FROM ;
  wire N141517;
  wire \DLX_IDinst_branch_address<17>/FROM ;
  wire N140824;
  wire \DLX_IFinst_NPC<31>/FROM ;
  wire \DLX_IFinst_NPC<15>/FROM ;
  wire \DLX_IFinst_NPC<15>/GROM ;
  wire \DLX_IFinst_NPC<23>/FROM ;
  wire \DLX_IDinst_branch_address<26>/FROM ;
  wire N141454;
  wire \DLX_IDinst_branch_address<18>/FROM ;
  wire N140887;
  wire \DLX_IDinst_branch_address<19>/FROM ;
  wire N140950;
  wire \DLX_IDinst_branch_address<27>/FROM ;
  wire N141391;
  wire \DLX_IDinst_reg_out_B<28>/GROM ;
  wire \DLX_IDinst_branch_address<28>/FROM ;
  wire N141328;
  wire \DLX_IDinst_branch_address<29>/FROM ;
  wire N141265;
  wire \DLX_IFinst_NPC<24>/FROM ;
  wire \DLX_IFinst_NPC<16>/FROM ;
  wire \DLX_IDinst_RegFile_0_7/FROM ;
  wire \DLX_IDinst_RegFile_0_7/GROM ;
  wire \DLX_IFinst_NPC<25>/FROM ;
  wire \DLX_IFinst_NPC<17>/FROM ;
  wire \DLX_IFinst_NPC<26>/FROM ;
  wire \DLX_IFinst_NPC<18>/FROM ;
  wire \DLX_EXinst_N73599/FROM ;
  wire \DLX_EXinst_N73599/GROM ;
  wire \DLX_IFinst_NPC<27>/FROM ;
  wire \DLX_IFinst_NPC<19>/FROM ;
  wire \DLX_MEMinst_opcode_of_WB<2>/FROM ;
  wire \DLX_MEMinst_opcode_of_WB<2>/GROM ;
  wire \DLX_IFinst_NPC<28>/FROM ;
  wire \DLX_IFinst_NPC<29>/FROM ;
  wire \N164596/FROM ;
  wire \N164596/GROM ;
  wire \DLX_EXinst_Mshift__n0019_Sh<127>/FROM ;
  wire \DLX_EXinst_Mshift__n0019_Sh<127>/GROM ;
  wire \N164138/FROM ;
  wire \N164138/GROM ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_65;
  wire \DLX_IDinst_RegFile_12_0/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_66;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_6;
  wire \DLX_IDinst_RegFile_12_0/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_12_0/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_69;
  wire \DLX_IDinst_RegFile_20_0/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_70;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_10;
  wire \DLX_IDinst_RegFile_20_0/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_20_0/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_81;
  wire \DLX_IDinst_RegFile_12_1/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_82;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_22;
  wire \DLX_IDinst_RegFile_12_1/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_12_1/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_85;
  wire \DLX_IDinst_RegFile_20_1/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_86;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_26;
  wire \DLX_IDinst_RegFile_20_1/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_20_1/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_97;
  wire \DLX_IDinst_RegFile_12_2/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_98;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_38;
  wire \DLX_IDinst_RegFile_12_2/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_12_2/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_101;
  wire \DLX_IDinst_RegFile_20_2/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_102;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_42;
  wire \DLX_IDinst_RegFile_20_2/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_20_2/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_113;
  wire \DLX_IDinst_RegFile_12_3/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_114;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_54;
  wire \DLX_IDinst_RegFile_12_3/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_12_3/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_117;
  wire \DLX_IDinst_RegFile_20_3/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_118;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_58;
  wire \DLX_IDinst_RegFile_20_3/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_20_3/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_129;
  wire \DLX_IDinst_RegFile_12_4/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_130;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_70;
  wire \DLX_IDinst_RegFile_12_4/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_12_4/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_593;
  wire \DLX_IDinst_RegFile_13_0/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_594;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_518;
  wire \DLX_IDinst_RegFile_13_0/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_13_0/CYINIT ;
  wire \DLX_IDinst_rd_addr<3>/FROM ;
  wire \DLX_IDinst_rd_addr<4>/FROM ;
  wire \N163428/FROM ;
  wire \N163428/GROM ;
  wire \N164207/FROM ;
  wire \N164207/GROM ;
  wire \N163656/FROM ;
  wire \N163656/GROM ;
  wire \N163501/FROM ;
  wire \N163501/GROM ;
  wire \DLX_IDinst_Mmux_IR_latched_Result<21>1_5/FROM ;
  wire \DLX_IDinst_Mmux_IR_latched_Result<21>1_5/GROM ;
  wire \DLX_IDinst_Mmux_IR_latched_Result<21>1_4/FROM ;
  wire \DLX_IDinst_Mmux_IR_latched_Result<21>1_4/GROM ;
  wire \DLX_IDinst_current_IR<21>/FROM ;
  wire \DLX_IDinst_current_IR<21>/GROM ;
  wire \DLX_EXinst_N72938/FROM ;
  wire \DLX_EXinst_N72938/GROM ;
  wire \DLX_EXinst_N73033/FROM ;
  wire \DLX_EXinst_N73033/GROM ;
  wire \DLX_EXinst_N73123/FROM ;
  wire \DLX_EXinst_N73123/GROM ;
  wire \DLX_EXinst_N72868/FROM ;
  wire \DLX_EXinst_N72868/GROM ;
  wire \DLX_EXinst_N74003/GROM ;
  wire \DLX_EXinst_N72933/FROM ;
  wire \DLX_EXinst_N72933/GROM ;
  wire \DLX_EXinst_N72848/FROM ;
  wire \DLX_EXinst_N72848/GROM ;
  wire \DLX_EXinst_N73133/FROM ;
  wire \DLX_EXinst_N73133/GROM ;
  wire \DLX_EXinst_N73138/FROM ;
  wire \DLX_EXinst_N73138/GROM ;
  wire \DLX_EXinst_N73118/FROM ;
  wire \DLX_EXinst_N73118/GROM ;
  wire \DLX_EXinst_N73038/FROM ;
  wire \DLX_EXinst_N73038/GROM ;
  wire \DLX_EXinst_N72973/FROM ;
  wire \DLX_EXinst_N72973/GROM ;
  wire \DLX_EXinst_N73063/FROM ;
  wire \DLX_EXinst_N73063/GROM ;
  wire \DLX_EXinst_N72953/FROM ;
  wire \DLX_EXinst_N72953/GROM ;
  wire \DLX_EXinst_N73048/FROM ;
  wire \DLX_EXinst_N73048/GROM ;
  wire \DLX_EXinst_N74024/FROM ;
  wire \DLX_EXinst_N74024/GROM ;
  wire \DLX_EXinst_N72978/FROM ;
  wire \DLX_EXinst_N72978/GROM ;
  wire \DLX_EXinst_N74034/FROM ;
  wire \DLX_EXinst_N74034/GROM ;
  wire \DLX_EXinst_N73211/FROM ;
  wire \DLX_EXinst_N73211/GROM ;
  wire \DLX_EXinst_N74451/FROM ;
  wire \DLX_EXinst_N74451/GROM ;
  wire \DLX_EXinst_N73148/FROM ;
  wire \DLX_EXinst_N73148/GROM ;
  wire \DLX_EXinst_N73068/FROM ;
  wire \DLX_EXinst_N73068/GROM ;
  wire \DLX_EXinst_N73534/FROM ;
  wire \DLX_EXinst_N73534/GROM ;
  wire \DLX_EXinst_N74029/FROM ;
  wire \DLX_EXinst_N74029/GROM ;
  wire \DLX_IDinst_Mmux_IR_latched_Result<16>1_5/FROM ;
  wire \DLX_IDinst_Mmux_IR_latched_Result<16>1_5/GROM ;
  wire \DLX_IDinst_Mmux_IR_latched_Result<16>1_4/FROM ;
  wire \DLX_IDinst_Mmux_IR_latched_Result<16>1_4/GROM ;
  wire \DLX_EXinst_N74206/FROM ;
  wire \DLX_EXinst_N74206/GROM ;
  wire \DLX_EXinst_N73158/FROM ;
  wire \DLX_EXinst_N73158/GROM ;
  wire \DLX_EXinst_N73594/FROM ;
  wire \DLX_EXinst_N73594/GROM ;
  wire \DLX_IDinst_current_IR<16>/FROM ;
  wire \DLX_IDinst_current_IR<16>/GROM ;
  wire \N164579/FROM ;
  wire \N164579/GROM ;
  wire \DLX_EXinst_N73239/FROM ;
  wire \DLX_EXinst_N73239/GROM ;
  wire \DLX_EXinst_N73088/FROM ;
  wire \DLX_EXinst_N73088/GROM ;
  wire \DLX_EXinst_N73499/FROM ;
  wire \DLX_EXinst_N73499/GROM ;
  wire \DLX_EXinst_N73345/FROM ;
  wire \DLX_EXinst_N73345/GROM ;
  wire \DLX_EXinst_N73514/FROM ;
  wire \DLX_EXinst_N73514/GROM ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_133;
  wire \DLX_IDinst_RegFile_20_4/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_134;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_74;
  wire \DLX_IDinst_RegFile_20_4/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_20_4/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_597;
  wire \DLX_IDinst_RegFile_21_0/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_598;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_522;
  wire \DLX_IDinst_RegFile_21_0/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_21_0/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_145;
  wire \DLX_IDinst_RegFile_12_5/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_146;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_86;
  wire \DLX_IDinst_RegFile_12_5/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_12_5/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_609;
  wire \DLX_IDinst_RegFile_13_1/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_610;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_534;
  wire \DLX_IDinst_RegFile_13_1/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_13_1/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_149;
  wire \DLX_IDinst_RegFile_20_5/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_150;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_90;
  wire \DLX_IDinst_RegFile_20_5/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_20_5/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_613;
  wire \DLX_IDinst_RegFile_21_1/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_614;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_538;
  wire \DLX_IDinst_RegFile_21_1/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_21_1/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_161;
  wire \DLX_IDinst_RegFile_12_6/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_162;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_102;
  wire \DLX_IDinst_RegFile_12_6/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_12_6/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_625;
  wire \DLX_IDinst_RegFile_13_2/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_626;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_550;
  wire \DLX_IDinst_RegFile_13_2/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_13_2/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_165;
  wire \DLX_IDinst_RegFile_20_6/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_166;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_106;
  wire \DLX_IDinst_RegFile_20_6/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_20_6/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_629;
  wire \DLX_IDinst_RegFile_21_2/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_630;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_554;
  wire \DLX_IDinst_RegFile_21_2/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_21_2/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_177;
  wire \DLX_IDinst_RegFile_12_7/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_178;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_118;
  wire \DLX_IDinst_RegFile_12_7/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_12_7/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_641;
  wire \DLX_IDinst_RegFile_13_3/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_642;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_566;
  wire \DLX_IDinst_RegFile_13_3/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_13_3/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_181;
  wire \DLX_IDinst_RegFile_20_7/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_182;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_122;
  wire \DLX_IDinst_RegFile_20_7/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_20_7/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_645;
  wire \DLX_IDinst_RegFile_21_3/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_646;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_570;
  wire \DLX_IDinst_RegFile_21_3/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_21_3/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_193;
  wire \DLX_IDinst_RegFile_12_8/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_194;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_134;
  wire \DLX_IDinst_RegFile_12_8/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_12_8/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_657;
  wire \DLX_IDinst_RegFile_13_4/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_658;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_582;
  wire \DLX_IDinst_RegFile_13_4/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_13_4/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_197;
  wire \DLX_IDinst_RegFile_20_8/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_198;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_138;
  wire \DLX_IDinst_RegFile_20_8/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_20_8/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_661;
  wire \DLX_IDinst_RegFile_21_4/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_662;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_586;
  wire \DLX_IDinst_RegFile_21_4/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_21_4/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_73;
  wire \DLX_IDinst_RegFile_30_0/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_74;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_14;
  wire \DLX_IDinst_RegFile_30_0/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_30_0/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_209;
  wire \DLX_IDinst_RegFile_12_9/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_210;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_150;
  wire \DLX_IDinst_RegFile_12_9/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_12_9/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_673;
  wire \DLX_IDinst_RegFile_13_5/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_674;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_598;
  wire \DLX_IDinst_RegFile_13_5/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_13_5/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_213;
  wire \DLX_IDinst_RegFile_20_9/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_214;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_154;
  wire \DLX_IDinst_RegFile_20_9/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_20_9/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_677;
  wire \DLX_IDinst_RegFile_21_5/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_678;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_602;
  wire \DLX_IDinst_RegFile_21_5/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_21_5/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_89;
  wire \DLX_IDinst_RegFile_30_1/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_90;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_30;
  wire \DLX_IDinst_RegFile_30_1/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_30_1/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_689;
  wire \DLX_IDinst_RegFile_13_6/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_690;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_614;
  wire \DLX_IDinst_RegFile_13_6/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_13_6/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_693;
  wire \DLX_IDinst_RegFile_21_6/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_694;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_618;
  wire \DLX_IDinst_RegFile_21_6/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_21_6/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_105;
  wire \DLX_IDinst_RegFile_30_2/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_106;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_46;
  wire \DLX_IDinst_RegFile_30_2/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_30_2/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_705;
  wire \DLX_IDinst_RegFile_13_7/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_706;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_630;
  wire \DLX_IDinst_RegFile_13_7/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_13_7/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_709;
  wire \DLX_IDinst_RegFile_21_7/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_710;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_634;
  wire \DLX_IDinst_RegFile_21_7/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_21_7/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_121;
  wire \DLX_IDinst_RegFile_30_3/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_122;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_62;
  wire \DLX_IDinst_RegFile_30_3/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_30_3/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_721;
  wire \DLX_IDinst_RegFile_13_8/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_722;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_646;
  wire \DLX_IDinst_RegFile_13_8/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_13_8/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_725;
  wire \DLX_IDinst_RegFile_21_8/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_726;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_650;
  wire \DLX_IDinst_RegFile_21_8/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_21_8/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_137;
  wire \DLX_IDinst_RegFile_30_4/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_138;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_78;
  wire \DLX_IDinst_RegFile_30_4/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_30_4/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_601;
  wire \DLX_IDinst_RegFile_31_0/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_602;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_526;
  wire \DLX_IDinst_RegFile_31_0/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_31_0/CYINIT ;
  wire \N136748/FROM ;
  wire \N136748/GROM ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_737;
  wire \DLX_IDinst_RegFile_13_9/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_738;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_662;
  wire \DLX_IDinst_RegFile_13_9/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_13_9/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_741;
  wire \DLX_IDinst_RegFile_21_9/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_742;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_666;
  wire \DLX_IDinst_RegFile_21_9/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_21_9/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_153;
  wire \DLX_IDinst_RegFile_30_5/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_154;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_94;
  wire \DLX_IDinst_RegFile_30_5/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_30_5/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_617;
  wire \DLX_IDinst_RegFile_31_1/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_618;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_542;
  wire \DLX_IDinst_RegFile_31_1/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_31_1/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_169;
  wire \DLX_IDinst_RegFile_30_6/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_170;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_110;
  wire \DLX_IDinst_RegFile_30_6/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_30_6/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_633;
  wire \DLX_IDinst_RegFile_31_2/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_634;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_558;
  wire \DLX_IDinst_RegFile_31_2/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_31_2/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_185;
  wire \DLX_IDinst_RegFile_30_7/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_186;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_126;
  wire \DLX_IDinst_RegFile_30_7/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_30_7/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_649;
  wire \DLX_IDinst_RegFile_31_3/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_650;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_574;
  wire \DLX_IDinst_RegFile_31_3/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_31_3/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_67;
  wire \DLX_IDinst_RegFile_16_0/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_68;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_8;
  wire \DLX_IDinst_RegFile_16_0/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_16_0/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_71;
  wire \DLX_IDinst_RegFile_24_0/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_72;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_12;
  wire \DLX_IDinst_RegFile_24_0/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_24_0/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_201;
  wire \DLX_IDinst_RegFile_30_8/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_202;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_142;
  wire \DLX_IDinst_RegFile_30_8/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_30_8/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_665;
  wire \DLX_IDinst_RegFile_31_4/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_666;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_590;
  wire \DLX_IDinst_RegFile_31_4/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_31_4/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_83;
  wire \DLX_IDinst_RegFile_16_1/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_84;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_24;
  wire \DLX_IDinst_RegFile_16_1/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_16_1/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_87;
  wire \DLX_IDinst_RegFile_24_1/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_88;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_28;
  wire \DLX_IDinst_RegFile_24_1/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_24_1/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_217;
  wire \DLX_IDinst_RegFile_30_9/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_218;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_158;
  wire \DLX_IDinst_RegFile_30_9/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_30_9/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_681;
  wire \DLX_IDinst_RegFile_31_5/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_682;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_606;
  wire \DLX_IDinst_RegFile_31_5/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_31_5/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_627;
  wire \DLX_IDinst_RegFile_16_2/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_628;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_552;
  wire \DLX_IDinst_RegFile_16_2/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_16_2/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_103;
  wire \DLX_IDinst_RegFile_24_2/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_104;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_44;
  wire \DLX_IDinst_RegFile_24_2/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_24_2/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_697;
  wire \DLX_IDinst_RegFile_31_6/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_698;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_622;
  wire \DLX_IDinst_RegFile_31_6/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_31_6/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_115;
  wire \DLX_IDinst_RegFile_16_3/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_116;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_56;
  wire \DLX_IDinst_RegFile_16_3/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_16_3/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_119;
  wire \DLX_IDinst_RegFile_24_3/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_120;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_60;
  wire \DLX_IDinst_RegFile_24_3/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_24_3/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_713;
  wire \DLX_IDinst_RegFile_31_7/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_714;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_638;
  wire \DLX_IDinst_RegFile_31_7/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_31_7/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_131;
  wire \DLX_IDinst_RegFile_16_4/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_132;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_72;
  wire \DLX_IDinst_RegFile_16_4/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_16_4/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_595;
  wire \DLX_IDinst_RegFile_17_0/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_596;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_520;
  wire \DLX_IDinst_RegFile_17_0/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_17_0/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_135;
  wire \DLX_IDinst_RegFile_24_4/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_136;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_76;
  wire \DLX_IDinst_RegFile_24_4/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_24_4/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_599;
  wire \DLX_IDinst_RegFile_25_0/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_600;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_524;
  wire \DLX_IDinst_RegFile_25_0/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_25_0/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_729;
  wire \DLX_IDinst_RegFile_31_8/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_730;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_654;
  wire \DLX_IDinst_RegFile_31_8/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_31_8/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_147;
  wire \DLX_IDinst_RegFile_16_5/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_148;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_88;
  wire \DLX_IDinst_RegFile_16_5/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_16_5/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_611;
  wire \DLX_IDinst_RegFile_17_1/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_612;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_536;
  wire \DLX_IDinst_RegFile_17_1/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_17_1/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_151;
  wire \DLX_IDinst_RegFile_24_5/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_152;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_92;
  wire \DLX_IDinst_RegFile_24_5/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_24_5/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_615;
  wire \DLX_IDinst_RegFile_25_1/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_616;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_540;
  wire \DLX_IDinst_RegFile_25_1/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_25_1/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_745;
  wire \DLX_IDinst_RegFile_31_9/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_746;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_670;
  wire \DLX_IDinst_RegFile_31_9/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_31_9/CYINIT ;
  wire \CHOICE3139/GROM ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_163;
  wire \DLX_IDinst_RegFile_16_6/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_164;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_104;
  wire \DLX_IDinst_RegFile_16_6/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_16_6/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_167;
  wire \DLX_IDinst_RegFile_24_6/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_168;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_108;
  wire \DLX_IDinst_RegFile_24_6/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_24_6/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_707;
  wire \DLX_IDinst_RegFile_16_7/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_708;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_632;
  wire \DLX_IDinst_RegFile_16_7/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_16_7/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_643;
  wire \DLX_IDinst_RegFile_17_3/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_644;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_568;
  wire \DLX_IDinst_RegFile_17_3/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_17_3/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_183;
  wire \DLX_IDinst_RegFile_24_7/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_184;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_124;
  wire \DLX_IDinst_RegFile_24_7/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_24_7/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_647;
  wire \DLX_IDinst_RegFile_25_3/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_648;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_572;
  wire \DLX_IDinst_RegFile_25_3/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_25_3/CYINIT ;
  wire \CHOICE3455/GROM ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_195;
  wire \DLX_IDinst_RegFile_16_8/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_196;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_136;
  wire \DLX_IDinst_RegFile_16_8/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_16_8/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_659;
  wire \DLX_IDinst_RegFile_17_4/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_660;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_584;
  wire \DLX_IDinst_RegFile_17_4/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_17_4/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_199;
  wire \DLX_IDinst_RegFile_24_8/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_200;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_140;
  wire \DLX_IDinst_RegFile_24_8/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_24_8/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_663;
  wire \DLX_IDinst_RegFile_25_4/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_664;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_588;
  wire \DLX_IDinst_RegFile_25_4/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_25_4/CYINIT ;
  wire \CHOICE3251/FROM ;
  wire \CHOICE3251/GROM ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_211;
  wire \DLX_IDinst_RegFile_16_9/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_212;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_152;
  wire \DLX_IDinst_RegFile_16_9/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_16_9/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_675;
  wire \DLX_IDinst_RegFile_17_5/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_676;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_600;
  wire \DLX_IDinst_RegFile_17_5/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_17_5/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_215;
  wire \DLX_IDinst_RegFile_24_9/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_216;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_156;
  wire \DLX_IDinst_RegFile_24_9/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_24_9/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_679;
  wire \DLX_IDinst_RegFile_25_5/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_680;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_604;
  wire \DLX_IDinst_RegFile_25_5/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_25_5/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_691;
  wire \DLX_IDinst_RegFile_17_6/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_692;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_616;
  wire \DLX_IDinst_RegFile_17_6/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_17_6/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_695;
  wire \DLX_IDinst_RegFile_25_6/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_696;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_620;
  wire \DLX_IDinst_RegFile_25_6/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_25_6/CYINIT ;
  wire \vga_top_vga1_helpcounter<2>/GROM ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_711;
  wire \DLX_IDinst_RegFile_25_7/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_712;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_636;
  wire \DLX_IDinst_RegFile_25_7/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_25_7/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_727;
  wire \DLX_IDinst_RegFile_25_8/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_728;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_652;
  wire \DLX_IDinst_RegFile_25_8/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_25_8/CYINIT ;
  wire \DLX_IFinst_IR_previous<22>/FROM ;
  wire \DLX_IFinst_IR_previous<22>/GROM ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_739;
  wire \DLX_IDinst_RegFile_17_9/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_740;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_664;
  wire \DLX_IDinst_RegFile_17_9/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_17_9/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_743;
  wire \DLX_IDinst_RegFile_25_9/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_744;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_668;
  wire \DLX_IDinst_RegFile_25_9/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_25_9/CYINIT ;
  wire \DLX_IFinst_IR_curr_N3087/FROM ;
  wire \DLX_IFinst_IR_curr_N3087/GROM ;
  wire \DLX_IDinst_RegFile_6_9/FROM ;
  wire \DLX_IDinst_RegFile_6_9/GROM ;
  wire \N163432/FROM ;
  wire \N163432/GROM ;
  wire \CHOICE6002/FROM ;
  wire \CHOICE6002/GROM ;
  wire \DLX_EXinst__n0056/FROM ;
  wire \DLX_EXinst__n0056/GROM ;
  wire \DLX_IDinst_RegFile_2_14/FROM ;
  wire \DLX_IDinst_RegFile_2_14/GROM ;
  wire \DLX_EXinst__n0080/FROM ;
  wire \DLX_EXinst__n0080/GROM ;
  wire \DLX_EXinst__n0077/FROM ;
  wire \DLX_EXinst__n0077/GROM ;
  wire \DLX_EXinst__n0078/FROM ;
  wire \DLX_EXinst__n0078/GROM ;
  wire \DLX_IDinst_RegFile_0_21/FROM ;
  wire \DLX_IDinst_RegFile_0_21/GROM ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_221;
  wire \DLX_IDinst_RegFile_4_10/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_222;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_162;
  wire \DLX_IDinst_RegFile_4_10/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_4_10/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_237;
  wire \DLX_IDinst_RegFile_4_11/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_238;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_178;
  wire \DLX_IDinst_RegFile_4_11/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_4_11/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_253;
  wire \DLX_IDinst_RegFile_4_12/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_254;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_194;
  wire \DLX_IDinst_RegFile_4_12/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_4_12/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_381;
  wire \DLX_IDinst_RegFile_4_20/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_382;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_322;
  wire \DLX_IDinst_RegFile_4_20/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_4_20/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_269;
  wire \DLX_IDinst_RegFile_4_13/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_270;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_210;
  wire \DLX_IDinst_RegFile_4_13/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_4_13/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_397;
  wire \DLX_IDinst_RegFile_4_21/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_398;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_338;
  wire \DLX_IDinst_RegFile_4_21/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_4_21/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_285;
  wire \DLX_IDinst_RegFile_4_14/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_286;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_226;
  wire \DLX_IDinst_RegFile_4_14/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_4_14/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_413;
  wire \DLX_IDinst_RegFile_4_22/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_414;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_354;
  wire \DLX_IDinst_RegFile_4_22/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_4_22/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1069;
  wire \DLX_IDinst_RegFile_4_30/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1070;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_994;
  wire \DLX_IDinst_RegFile_4_30/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_4_30/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1085;
  wire \DLX_IDinst_RegFile_4_31/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1086;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_1010;
  wire \DLX_IDinst_RegFile_4_31/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_4_31/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_301;
  wire \DLX_IDinst_RegFile_4_15/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_302;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_242;
  wire \DLX_IDinst_RegFile_4_15/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_4_15/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_429;
  wire \DLX_IDinst_RegFile_4_23/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_430;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_370;
  wire \DLX_IDinst_RegFile_4_23/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_4_23/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_317;
  wire \DLX_IDinst_RegFile_4_16/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_318;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_258;
  wire \DLX_IDinst_RegFile_4_16/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_4_16/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_445;
  wire \DLX_IDinst_RegFile_4_24/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_446;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_386;
  wire \DLX_IDinst_RegFile_4_24/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_4_24/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_333;
  wire \DLX_IDinst_RegFile_4_17/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_334;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_274;
  wire \DLX_IDinst_RegFile_4_17/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_4_17/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_461;
  wire \DLX_IDinst_RegFile_4_25/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_462;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_402;
  wire \DLX_IDinst_RegFile_4_25/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_4_25/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_349;
  wire \DLX_IDinst_RegFile_4_18/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_350;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_290;
  wire \DLX_IDinst_RegFile_4_18/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_4_18/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_477;
  wire \DLX_IDinst_RegFile_4_26/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_478;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_418;
  wire \DLX_IDinst_RegFile_4_26/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_4_26/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_749;
  wire \DLX_IDinst_RegFile_5_10/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_750;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_674;
  wire \DLX_IDinst_RegFile_5_10/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_5_10/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_365;
  wire \DLX_IDinst_RegFile_4_19/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_366;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_306;
  wire \DLX_IDinst_RegFile_4_19/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_4_19/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_493;
  wire \DLX_IDinst_RegFile_4_27/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_494;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_434;
  wire \DLX_IDinst_RegFile_4_27/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_4_27/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_765;
  wire \DLX_IDinst_RegFile_5_11/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_766;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_690;
  wire \DLX_IDinst_RegFile_5_11/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_5_11/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1037;
  wire \DLX_IDinst_RegFile_4_28/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1038;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_962;
  wire \DLX_IDinst_RegFile_4_28/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_4_28/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_909;
  wire \DLX_IDinst_RegFile_5_20/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_910;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_834;
  wire \DLX_IDinst_RegFile_5_20/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_5_20/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_781;
  wire \DLX_IDinst_RegFile_5_12/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_782;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_706;
  wire \DLX_IDinst_RegFile_5_12/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_5_12/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1053;
  wire \DLX_IDinst_RegFile_4_29/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1054;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_978;
  wire \DLX_IDinst_RegFile_4_29/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_4_29/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_925;
  wire \DLX_IDinst_RegFile_5_21/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_926;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_850;
  wire \DLX_IDinst_RegFile_5_21/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_5_21/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_797;
  wire \DLX_IDinst_RegFile_5_13/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_798;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_722;
  wire \DLX_IDinst_RegFile_5_13/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_5_13/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_541;
  wire \DLX_IDinst_RegFile_5_30/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_542;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_482;
  wire \DLX_IDinst_RegFile_5_30/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_5_30/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_941;
  wire \DLX_IDinst_RegFile_5_22/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_942;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_866;
  wire \DLX_IDinst_RegFile_5_22/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_5_22/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_813;
  wire \DLX_IDinst_RegFile_5_14/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_814;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_738;
  wire \DLX_IDinst_RegFile_5_14/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_5_14/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_557;
  wire \DLX_IDinst_RegFile_5_31/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_558;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_498;
  wire \DLX_IDinst_RegFile_5_31/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_5_31/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_957;
  wire \DLX_IDinst_RegFile_5_23/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_958;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_882;
  wire \DLX_IDinst_RegFile_5_23/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_5_23/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_829;
  wire \DLX_IDinst_RegFile_5_15/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_830;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_754;
  wire \DLX_IDinst_RegFile_5_15/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_5_15/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_973;
  wire \DLX_IDinst_RegFile_5_24/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_974;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_898;
  wire \DLX_IDinst_RegFile_5_24/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_5_24/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_845;
  wire \DLX_IDinst_RegFile_5_16/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_846;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_770;
  wire \DLX_IDinst_RegFile_5_16/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_5_16/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_989;
  wire \DLX_IDinst_RegFile_5_25/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_990;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_914;
  wire \DLX_IDinst_RegFile_5_25/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_5_25/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_861;
  wire \DLX_IDinst_RegFile_5_17/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_862;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_786;
  wire \DLX_IDinst_RegFile_5_17/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_5_17/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1005;
  wire \DLX_IDinst_RegFile_5_26/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1006;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_930;
  wire \DLX_IDinst_RegFile_5_26/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_5_26/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_877;
  wire \DLX_IDinst_RegFile_5_18/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_878;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_802;
  wire \DLX_IDinst_RegFile_5_18/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_5_18/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1021;
  wire \DLX_IDinst_RegFile_5_27/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1022;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_946;
  wire \DLX_IDinst_RegFile_5_27/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_5_27/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_893;
  wire \DLX_IDinst_RegFile_5_19/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_894;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_818;
  wire \DLX_IDinst_RegFile_5_19/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_5_19/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_509;
  wire \DLX_IDinst_RegFile_5_28/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_510;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_450;
  wire \DLX_IDinst_RegFile_5_28/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_5_28/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_223;
  wire \DLX_IDinst_RegFile_8_10/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_224;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_164;
  wire \DLX_IDinst_RegFile_8_10/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_8_10/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_239;
  wire \DLX_IDinst_RegFile_8_11/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_240;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_180;
  wire \DLX_IDinst_RegFile_8_11/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_8_11/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_383;
  wire \DLX_IDinst_RegFile_8_20/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_384;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_324;
  wire \DLX_IDinst_RegFile_8_20/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_8_20/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_255;
  wire \DLX_IDinst_RegFile_8_12/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_256;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_196;
  wire \DLX_IDinst_RegFile_8_12/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_8_12/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_399;
  wire \DLX_IDinst_RegFile_8_21/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_400;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_340;
  wire \DLX_IDinst_RegFile_8_21/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_8_21/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_271;
  wire \DLX_IDinst_RegFile_8_13/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_272;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_212;
  wire \DLX_IDinst_RegFile_8_13/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_8_13/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1071;
  wire \DLX_IDinst_RegFile_8_30/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1072;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_996;
  wire \DLX_IDinst_RegFile_8_30/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_8_30/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_415;
  wire \DLX_IDinst_RegFile_8_22/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_416;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_356;
  wire \DLX_IDinst_RegFile_8_22/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_8_22/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_287;
  wire \DLX_IDinst_RegFile_8_14/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_288;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_228;
  wire \DLX_IDinst_RegFile_8_14/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_8_14/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_431;
  wire \DLX_IDinst_RegFile_8_23/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_432;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_372;
  wire \DLX_IDinst_RegFile_8_23/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_8_23/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_303;
  wire \DLX_IDinst_RegFile_8_15/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_304;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_244;
  wire \DLX_IDinst_RegFile_8_15/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_8_15/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1087;
  wire \DLX_IDinst_RegFile_8_31/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1088;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_1012;
  wire \DLX_IDinst_RegFile_8_31/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_8_31/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_447;
  wire \DLX_IDinst_RegFile_8_24/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_448;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_388;
  wire \DLX_IDinst_RegFile_8_24/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_8_24/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_319;
  wire \DLX_IDinst_RegFile_8_16/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_320;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_260;
  wire \DLX_IDinst_RegFile_8_16/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_8_16/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_463;
  wire \DLX_IDinst_RegFile_8_25/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_464;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_404;
  wire \DLX_IDinst_RegFile_8_25/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_8_25/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_335;
  wire \DLX_IDinst_RegFile_8_17/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_336;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_276;
  wire \DLX_IDinst_RegFile_8_17/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_8_17/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_479;
  wire \DLX_IDinst_RegFile_8_26/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_480;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_420;
  wire \DLX_IDinst_RegFile_8_26/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_8_26/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_351;
  wire \DLX_IDinst_RegFile_8_18/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_352;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_292;
  wire \DLX_IDinst_RegFile_8_18/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_8_18/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_751;
  wire \DLX_IDinst_RegFile_9_10/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_752;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_676;
  wire \DLX_IDinst_RegFile_9_10/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_9_10/CYINIT ;
  wire \N163827/FROM ;
  wire \N163827/GROM ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_495;
  wire \DLX_IDinst_RegFile_8_27/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_496;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_436;
  wire \DLX_IDinst_RegFile_8_27/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_8_27/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_367;
  wire \DLX_IDinst_RegFile_8_19/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_368;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_308;
  wire \DLX_IDinst_RegFile_8_19/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_8_19/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_767;
  wire \DLX_IDinst_RegFile_9_11/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_768;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_692;
  wire \DLX_IDinst_RegFile_9_11/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_9_11/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1039;
  wire \DLX_IDinst_RegFile_8_28/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1040;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_964;
  wire \DLX_IDinst_RegFile_8_28/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_8_28/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_911;
  wire \DLX_IDinst_RegFile_9_20/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_912;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_836;
  wire \DLX_IDinst_RegFile_9_20/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_9_20/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_783;
  wire \DLX_IDinst_RegFile_9_12/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_784;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_708;
  wire \DLX_IDinst_RegFile_9_12/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_9_12/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1055;
  wire \DLX_IDinst_RegFile_8_29/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1056;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_980;
  wire \DLX_IDinst_RegFile_8_29/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_8_29/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_927;
  wire \DLX_IDinst_RegFile_9_21/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_928;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_852;
  wire \DLX_IDinst_RegFile_9_21/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_9_21/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_799;
  wire \DLX_IDinst_RegFile_9_13/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_800;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_724;
  wire \DLX_IDinst_RegFile_9_13/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_9_13/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_543;
  wire \DLX_IDinst_RegFile_9_30/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_544;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_484;
  wire \DLX_IDinst_RegFile_9_30/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_9_30/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_943;
  wire \DLX_IDinst_RegFile_9_22/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_944;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_868;
  wire \DLX_IDinst_RegFile_9_22/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_9_22/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_959;
  wire \DLX_IDinst_RegFile_9_23/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_960;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_884;
  wire \DLX_IDinst_RegFile_9_23/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_9_23/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_831;
  wire \DLX_IDinst_RegFile_9_15/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_832;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_756;
  wire \DLX_IDinst_RegFile_9_15/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_9_15/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_559;
  wire \DLX_IDinst_RegFile_9_31/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_560;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_500;
  wire \DLX_IDinst_RegFile_9_31/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_9_31/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_975;
  wire \DLX_IDinst_RegFile_9_24/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_976;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_900;
  wire \DLX_IDinst_RegFile_9_24/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_9_24/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_847;
  wire \DLX_IDinst_RegFile_9_16/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_848;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_772;
  wire \DLX_IDinst_RegFile_9_16/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_9_16/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_991;
  wire \DLX_IDinst_RegFile_9_25/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_992;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_916;
  wire \DLX_IDinst_RegFile_9_25/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_9_25/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_863;
  wire \DLX_IDinst_RegFile_9_17/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_864;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_788;
  wire \DLX_IDinst_RegFile_9_17/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_9_17/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1007;
  wire \DLX_IDinst_RegFile_9_26/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1008;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_932;
  wire \DLX_IDinst_RegFile_9_26/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_9_26/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_879;
  wire \DLX_IDinst_RegFile_9_18/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_880;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_804;
  wire \DLX_IDinst_RegFile_9_18/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_9_18/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1023;
  wire \DLX_IDinst_RegFile_9_27/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1024;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_948;
  wire \DLX_IDinst_RegFile_9_27/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_9_27/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_895;
  wire \DLX_IDinst_RegFile_9_19/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_896;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_820;
  wire \DLX_IDinst_RegFile_9_19/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_9_19/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_511;
  wire \DLX_IDinst_RegFile_9_28/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_512;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_452;
  wire \DLX_IDinst_RegFile_9_28/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_9_28/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_527;
  wire \DLX_IDinst_RegFile_9_29/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_528;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_468;
  wire \DLX_IDinst_RegFile_9_29/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_9_29/CYINIT ;
  wire \N136625/FROM ;
  wire \N136625/GROM ;
  wire \DLX_MEMinst_opcode_of_WB<1>/GROM ;
  wire \DLX_IFinst_IR_previous<3>/FROM ;
  wire \DLX_IFinst_IR_previous<3>/GROM ;
  wire \DLX_IDinst_RegFile_3_28/FROM ;
  wire \DLX_IDinst_RegFile_3_28/GROM ;
  wire \DLX_IFinst_IR_previous<9>/FROM ;
  wire \DLX_IFinst_IR_previous<9>/GROM ;
  wire \N163210/FROM ;
  wire \N163210/GROM ;
  wire \DLX_IDinst_EPC<9>/FROM ;
  wire \DLX_IDinst_EPC<9>/GROM ;
  wire \DLX_IDinst_RegFile_0_10/FROM ;
  wire \DLX_IDinst_RegFile_0_10/GROM ;
  wire \DLX_IDinst_RegFile_2_1/FROM ;
  wire \DLX_IDinst_RegFile_2_1/GROM ;
  wire \DLX_IDinst_RegFile_0_20/FROM ;
  wire \DLX_IDinst_RegFile_0_20/GROM ;
  wire \N163708/FROM ;
  wire \N163708/GROM ;
  wire \DLX_IDinst_RegFile_30_31/FROM ;
  wire \DLX_IDinst_RegFile_30_31/GROM ;
  wire \N145644/FROM ;
  wire \N145644/GROM ;
  wire \N145073/FROM ;
  wire \N145073/GROM ;
  wire \DLX_IDinst_RegFile_2_2/FROM ;
  wire \DLX_IDinst_RegFile_2_2/GROM ;
  wire \N145258/FROM ;
  wire \N145258/GROM ;
  wire \N144481/FROM ;
  wire \N144481/GROM ;
  wire \DLX_IDinst_RegFile_2_3/FROM ;
  wire \DLX_IDinst_RegFile_2_3/GROM ;
  wire \N144646/FROM ;
  wire \N144646/GROM ;
  wire \CHOICE3449/FROM ;
  wire \CHOICE3449/GROM ;
  wire \DLX_IDinst_RegFile_2_4/FROM ;
  wire \DLX_IDinst_RegFile_2_4/GROM ;
  wire \N145443/FROM ;
  wire \N145443/GROM ;
  wire \DLX_IDinst_RegFile_31_13/FROM ;
  wire \DLX_IDinst_RegFile_31_13/GROM ;
  wire \DLX_IDinst__n0311/FROM ;
  wire \DLX_IDinst__n0311/GROM ;
  wire \CHOICE3321/FROM ;
  wire \CHOICE3321/GROM ;
  wire \DLX_IDinst_RegFile_31_22/FROM ;
  wire \DLX_IDinst_RegFile_31_22/GROM ;
  wire \DLX_IDinst_RegFile_15_31/FROM ;
  wire \DLX_IDinst_RegFile_15_31/GROM ;
  wire \DLX_IDinst_RegFile_31_16/FROM ;
  wire \DLX_IDinst_RegFile_31_16/GROM ;
  wire \DLX_IDinst_RegFile_15_18/FROM ;
  wire \DLX_IDinst_RegFile_15_18/GROM ;
  wire \DLX_IDinst_RegFile_15_19/FROM ;
  wire \DLX_IDinst_RegFile_15_19/GROM ;
  wire \DLX_IDinst_RegFile_19_0/FROM ;
  wire \DLX_IDinst_RegFile_19_0/GROM ;
  wire \DLX_IDinst__n0097/FROM ;
  wire \DLX_IDinst__n0097/GROM ;
  wire \DLX_IDinst__n0629<1>/FROM ;
  wire \DLX_IDinst__n0629<1>/GROM ;
  wire \DLX_IDinst__n0436/GROM ;
  wire \DLX_IFinst_IR_curr<13>/FROM ;
  wire \DLX_IFinst_IR_curr<13>/GROM ;
  wire \DLX_IDinst_RegFile_24_30/FROM ;
  wire \DLX_IDinst_RegFile_24_30/GROM ;
  wire \DLX_IFinst_IR_curr<30>/FROM ;
  wire \DLX_IFinst_IR_curr<30>/GROM ;
  wire \DLX_IDinst_RegFile_17_17/FROM ;
  wire \DLX_IDinst_RegFile_17_17/GROM ;
  wire \DLX_IFinst_IR_curr<22>/FROM ;
  wire \DLX_IFinst_IR_curr<22>/GROM ;
  wire \DLX_IFinst_IR_curr<14>/FROM ;
  wire \DLX_IFinst_IR_curr<14>/GROM ;
  wire \DLX_IFinst_IR_curr<23>/FROM ;
  wire \DLX_IFinst_IR_curr<23>/GROM ;
  wire \DLX_IDinst_RegFile_19_29/FROM ;
  wire \DLX_IDinst_RegFile_19_29/GROM ;
  wire \DLX_IDinst_RegFile_0_3/FROM ;
  wire \DLX_IDinst_RegFile_0_3/GROM ;
  wire \DLX_EXinst_ALU_result<5>/FROM ;
  wire \DLX_EXinst_ALU_result<5>/GROM ;
  wire \DLX_IDinst_RegFile_23_1/FROM ;
  wire \DLX_IDinst_RegFile_23_1/GROM ;
  wire \DLX_IDinst_RegFile_14_6/FROM ;
  wire \DLX_IDinst_RegFile_14_6/GROM ;
  wire \DLX_IDinst_RegFile_0_5/FROM ;
  wire \DLX_IDinst_RegFile_0_5/GROM ;
  wire \DLX_IFinst_IR_curr<17>/FROM ;
  wire \DLX_IFinst_IR_curr<17>/GROM ;
  wire \DLX_IFinst_IR_curr<26>/FROM ;
  wire \DLX_IFinst_IR_curr<26>/GROM ;
  wire \DLX_IFinst_IR_curr<18>/FROM ;
  wire \DLX_IFinst_IR_curr<18>/GROM ;
  wire \DLX_IDinst_RegFile_14_7/FROM ;
  wire \DLX_IDinst_RegFile_14_7/GROM ;
  wire \DLX_IDinst_RegFile_11_20/FROM ;
  wire \DLX_IDinst_RegFile_11_20/GROM ;
  wire \DLX_IDinst_RegFile_11_30/FROM ;
  wire \DLX_IDinst_RegFile_11_30/GROM ;
  wire \DLX_IDinst_RegFile_11_15/FROM ;
  wire \DLX_IDinst_RegFile_11_15/GROM ;
  wire \CHOICE3784/FROM ;
  wire \CHOICE3784/GROM ;
  wire \DLX_IDinst_RegFile_11_25/FROM ;
  wire \DLX_IDinst_RegFile_11_25/GROM ;
  wire \N163538/FROM ;
  wire \N163538/GROM ;
  wire \DLX_IDinst_RegFile_1_24/FROM ;
  wire \DLX_IDinst_RegFile_1_24/GROM ;
  wire \CHOICE3729/FROM ;
  wire \CHOICE3729/GROM ;
  wire \DLX_IDinst_RegFile_23_3/FROM ;
  wire \DLX_IDinst_RegFile_23_3/GROM ;
  wire \DLX_IDinst_RegFile_14_8/FROM ;
  wire \DLX_IDinst_RegFile_14_8/GROM ;
  wire \DLX_IDinst_RegFile_3_2/FROM ;
  wire \DLX_IDinst_RegFile_3_2/GROM ;
  wire \DLX_IDinst_RegFile_3_3/FROM ;
  wire \DLX_IDinst_RegFile_3_3/GROM ;
  wire \CHOICE3674/FROM ;
  wire \CHOICE3674/GROM ;
  wire \DLX_IDinst_RegFile_22_9/FROM ;
  wire \DLX_IDinst_RegFile_22_9/GROM ;
  wire \DLX_IDinst_RegFile_7_5/FROM ;
  wire \DLX_IDinst_RegFile_7_5/GROM ;
  wire \DLX_IDinst_RegFile_2_8/FROM ;
  wire \DLX_IDinst_RegFile_2_8/GROM ;
  wire \DLX_IDinst_RegFile_23_7/FROM ;
  wire \DLX_IDinst_RegFile_23_7/GROM ;
  wire \CHOICE4282/FROM ;
  wire \CHOICE4282/GROM ;
  wire \CHOICE4285/FROM ;
  wire \CHOICE4285/GROM ;
  wire \DLX_IDinst_RegFile_27_23/FROM ;
  wire \DLX_IDinst_RegFile_27_23/GROM ;
  wire \DLX_IDinst_RegFile_3_5/FROM ;
  wire \DLX_IDinst_RegFile_3_5/GROM ;
  wire \DLX_IFinst_IR_previous<11>/FROM ;
  wire \DLX_IFinst_IR_previous<11>/GROM ;
  wire \CHOICE5741/FROM ;
  wire \CHOICE5741/GROM ;
  wire \DLX_MEMinst_RF_data_in<24>/GROM ;
  wire \CHOICE5967/FROM ;
  wire \CHOICE5967/GROM ;
  wire \DLX_IDinst_RegFile_2_9/FROM ;
  wire \DLX_IDinst_RegFile_2_9/GROM ;
  wire \DLX_IFinst_IR_previous<23>/FROM ;
  wire \DLX_IFinst_IR_previous<23>/GROM ;
  wire \DLX_IDinst_RegFile_10_1/FROM ;
  wire \DLX_IDinst_RegFile_10_1/GROM ;
  wire \DLX_IDinst_RegFile_10_2/FROM ;
  wire \DLX_IDinst_RegFile_10_2/GROM ;
  wire \CHOICE5081/FROM ;
  wire \CHOICE5081/GROM ;
  wire \CHOICE5938/FROM ;
  wire \CHOICE5938/GROM ;
  wire \DLX_IDinst_RegFile_10_4/FROM ;
  wire \DLX_IDinst_RegFile_10_4/GROM ;
  wire \CHOICE6008/FROM ;
  wire \CHOICE6008/GROM ;
  wire \CHOICE5751/FROM ;
  wire \CHOICE5751/GROM ;
  wire \DLX_IDinst_RegFile_10_5/FROM ;
  wire \DLX_IDinst_RegFile_10_5/GROM ;
  wire \DLX_IDinst_RegFile_11_1/FROM ;
  wire \DLX_IDinst_RegFile_11_1/GROM ;
  wire \DLX_IFinst_IR_previous<28>/FROM ;
  wire \DLX_IFinst_IR_previous<28>/GROM ;
  wire \DLX_IFinst_IR_previous<29>/FROM ;
  wire \DLX_IFinst_IR_previous<29>/GROM ;
  wire \CHOICE5562/FROM ;
  wire \CHOICE5562/GROM ;
  wire \CHOICE4947/FROM ;
  wire \CHOICE4947/GROM ;
  wire \CHOICE5572/FROM ;
  wire \CHOICE5572/GROM ;
  wire \DLX_IDinst_RegFile_10_7/FROM ;
  wire \DLX_IDinst_RegFile_10_7/GROM ;
  wire \CHOICE5486/FROM ;
  wire \CHOICE5486/GROM ;
  wire \CHOICE5496/FROM ;
  wire \CHOICE5496/GROM ;
  wire \DLX_IDinst_RegFile_6_10/FROM ;
  wire \DLX_IDinst_RegFile_6_10/GROM ;
  wire \DLX_IDinst_RegFile_10_8/FROM ;
  wire \DLX_IDinst_RegFile_10_8/GROM ;
  wire \DLX_EXinst_ALU_result<4>/FROM ;
  wire \DLX_EXinst_ALU_result<4>/GROM ;
  wire \DLX_IDinst_RegFile_6_11/FROM ;
  wire \DLX_IDinst_RegFile_6_11/GROM ;
  wire \DLX_IFinst_PC<11>/FROM ;
  wire \DLX_IFinst_PC<11>/GROM ;
  wire \CHOICE3986/FROM ;
  wire \CHOICE3986/GROM ;
  wire \DLX_IDinst_RegFile_14_31/FROM ;
  wire \DLX_IDinst_RegFile_14_31/GROM ;
  wire \CHOICE3927/FROM ;
  wire \CHOICE3927/GROM ;
  wire \CHOICE3851/FROM ;
  wire \CHOICE3851/GROM ;
  wire \DLX_IDinst_RegFile_30_16/FROM ;
  wire \DLX_IDinst_RegFile_30_16/GROM ;
  wire \DLX_IDinst_RegFile_22_17/FROM ;
  wire \DLX_IDinst_RegFile_22_17/GROM ;
  wire \CHOICE3868/FROM ;
  wire \CHOICE3868/GROM ;
  wire \CHOICE5165/GROM ;
  wire \DLX_IDinst_RegFile_14_18/FROM ;
  wire \DLX_IDinst_RegFile_14_18/GROM ;
  wire \DLX_IDinst_RegFile_6_21/FROM ;
  wire \DLX_IDinst_RegFile_6_21/GROM ;
  wire \N163489/FROM ;
  wire \N163489/GROM ;
  wire \N164119/FROM ;
  wire \N164119/GROM ;
  wire \DLX_IDinst_RegFile_23_10/FROM ;
  wire \DLX_IDinst_RegFile_23_10/GROM ;
  wire \DLX_IDinst_RegFile_5_29/FROM ;
  wire \DLX_IDinst_RegFile_5_29/GROM ;
  wire \DLX_IDinst_RegFile_14_27/FROM ;
  wire \DLX_IDinst_RegFile_14_27/GROM ;
  wire \DLX_IDinst_RegFile_6_22/FROM ;
  wire \DLX_IDinst_RegFile_6_22/GROM ;
  wire \DLX_IDinst_RegFile_22_19/FROM ;
  wire \DLX_IDinst_RegFile_22_19/GROM ;
  wire \DLX_IDinst_RegFile_6_14/FROM ;
  wire \DLX_IDinst_RegFile_6_14/GROM ;
  wire \DLX_IDinst_RegFile_6_30/FROM ;
  wire \DLX_IDinst_RegFile_6_30/GROM ;
  wire \DLX_IDinst_RegFile_6_31/FROM ;
  wire \DLX_IDinst_RegFile_6_31/GROM ;
  wire \DLX_IDinst_RegFile_6_15/FROM ;
  wire \DLX_IDinst_RegFile_6_15/GROM ;
  wire \DM_read_data<1>/FROM ;
  wire \DM_read_data<1>/GROM ;
  wire \DM_read_data<2>/FROM ;
  wire \DM_read_data<2>/GROM ;
  wire \DLX_IDinst_RegFile_6_24/FROM ;
  wire \DLX_IDinst_RegFile_6_24/GROM ;
  wire \DLX_IDinst_RegFile_6_17/FROM ;
  wire \DLX_IDinst_RegFile_6_17/GROM ;
  wire \DLX_IDinst_RegFile_6_25/FROM ;
  wire \DLX_IDinst_RegFile_6_25/GROM ;
  wire \DLX_IDinst_RegFile_7_10/FROM ;
  wire \DLX_IDinst_RegFile_7_10/GROM ;
  wire \DLX_IDinst_RegFile_6_18/FROM ;
  wire \DLX_IDinst_RegFile_6_18/GROM ;
  wire \CHOICE1669/FROM ;
  wire \CHOICE1669/GROM ;
  wire \DLX_IDinst_RegFile_15_17/FROM ;
  wire \DLX_IDinst_RegFile_15_17/GROM ;
  wire \N163688/FROM ;
  wire \N163688/GROM ;
  wire \N132648/FROM ;
  wire \N132648/GROM ;
  wire \DLX_IFinst_stalled/CEMUXNOT ;
  wire \DLX_IFinst_stalled/FROM ;
  wire \DLX_IFinst_stalled/GROM ;
  wire \N127012/FROM ;
  wire \N127012/GROM ;
  wire \DLX_IDinst_RegFile_6_27/FROM ;
  wire \DLX_IDinst_RegFile_6_27/GROM ;
  wire \N163230/FROM ;
  wire \N163230/GROM ;
  wire \DLX_IDinst_RegFile_31_18/FROM ;
  wire \DLX_IDinst_RegFile_31_18/GROM ;
  wire \N163664/FROM ;
  wire \N163664/GROM ;
  wire \DLX_IDinst_RegFile_7_20/FROM ;
  wire \DLX_IDinst_RegFile_7_20/GROM ;
  wire \DLX_IDinst_RegFile_23_27/FROM ;
  wire \DLX_IDinst_RegFile_23_27/GROM ;
  wire \DLX_IDinst_RegFile_7_12/FROM ;
  wire \DLX_IDinst_RegFile_7_12/GROM ;
  wire \DLX_IDinst_RegFile_31_19/FROM ;
  wire \DLX_IDinst_RegFile_31_19/GROM ;
  wire \reset_IBUF_5/GROM ;
  wire \CHOICE2112/FROM ;
  wire \CHOICE2112/GROM ;
  wire \DLX_EXinst_Mshift__n0021_Sh<0>/FROM ;
  wire \DLX_EXinst_Mshift__n0021_Sh<0>/GROM ;
  wire \DLX_EXinst_Mshift__n0021_Sh<40>/FROM ;
  wire \DLX_EXinst_Mshift__n0021_Sh<40>/GROM ;
  wire \DLX_EXinst_Mshift__n0021_Sh<1>/FROM ;
  wire \DLX_EXinst_Mshift__n0021_Sh<1>/GROM ;
  wire \DLX_EXinst_Mshift__n0021_Sh<42>/FROM ;
  wire \DLX_EXinst_Mshift__n0021_Sh<42>/GROM ;
  wire \N163442/FROM ;
  wire \N163442/GROM ;
  wire \DLX_EXinst_Mshift__n0021_Sh<8>/FROM ;
  wire \DLX_EXinst_Mshift__n0021_Sh<8>/GROM ;
  wire \DLX_IDinst_RegFile_10_30/FROM ;
  wire \DLX_IDinst_RegFile_10_30/GROM ;
  wire \DLX_IDinst_EPC<10>/FROM ;
  wire \DLX_IDinst_EPC<10>/GROM ;
  wire \DLX_IDinst_EPC<11>/FROM ;
  wire \DLX_IDinst_EPC<11>/GROM ;
  wire \DLX_IDinst_EPC<20>/FROM ;
  wire \DLX_IDinst_EPC<20>/GROM ;
  wire \DLX_IDinst_EPC<12>/FROM ;
  wire \DLX_IDinst_EPC<12>/GROM ;
  wire \DLX_IDinst_EPC<21>/FROM ;
  wire \DLX_IDinst_EPC<21>/GROM ;
  wire \DLX_IDinst_EPC<13>/FROM ;
  wire \DLX_IDinst_EPC<13>/GROM ;
  wire \DLX_IDinst_EPC<22>/FROM ;
  wire \DLX_IDinst_EPC<22>/GROM ;
  wire \DLX_IDinst_EPC<14>/FROM ;
  wire \DLX_IDinst_EPC<14>/GROM ;
  wire \DLX_IDinst_EPC<31>/FROM ;
  wire \DLX_IDinst_EPC<31>/GROM ;
  wire \DLX_IDinst_EPC<16>/FROM ;
  wire \DLX_IDinst_EPC<16>/GROM ;
  wire \DLX_IDinst_EPC<25>/FROM ;
  wire \DLX_IDinst_EPC<25>/GROM ;
  wire \DLX_IDinst_EPC<18>/FROM ;
  wire \DLX_IDinst_EPC<18>/GROM ;
  wire \DLX_IDinst_EPC<19>/FROM ;
  wire \DLX_IDinst_EPC<19>/GROM ;
  wire \DLX_IDinst_EPC<28>/FROM ;
  wire \DLX_IDinst_EPC<28>/GROM ;
  wire \N163680/FROM ;
  wire \N163680/GROM ;
  wire \N163700/FROM ;
  wire \N163700/GROM ;
  wire \N163325/FROM ;
  wire \N163325/GROM ;
  wire \vga_top_vga1_N112904/FROM ;
  wire \vga_top_vga1_N112904/GROM ;
  wire \DLX_EXinst_Mshift__n0023_Sh<0>/FROM ;
  wire \DLX_EXinst_Mshift__n0023_Sh<0>/GROM ;
  wire \vga_top_vga1_N112910/FROM ;
  wire \vga_top_vga1_N112910/GROM ;
  wire \DLX_EXinst_Mshift__n0023_Sh<1>/FROM ;
  wire \DLX_EXinst_Mshift__n0023_Sh<1>/GROM ;
  wire \vga_top_vga1_N112921/FROM ;
  wire \vga_top_vga1_N112921/GROM ;
  wire \vga_top_vga1_N112946/FROM ;
  wire \vga_top_vga1_N112946/GROM ;
  wire \vga_top_vga1_N112941/GROM ;
  wire \N163510/FROM ;
  wire \N163510/GROM ;
  wire \DLX_EXinst_Mshift__n0023_Sh<7>/FROM ;
  wire \DLX_EXinst_Mshift__n0023_Sh<7>/GROM ;
  wire \DLX_EXinst_Mshift__n0023_Sh<8>/FROM ;
  wire \DLX_EXinst_Mshift__n0023_Sh<8>/GROM ;
  wire \DLX_EXinst_N73023/FROM ;
  wire \DLX_EXinst_N73023/GROM ;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_261/FROM ;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_261/GROM ;
  wire \N163639/GROM ;
  wire \DLX_IDinst_branch_address<0>/FROM ;
  wire N145826;
  wire \DLX_IDinst_branch_address<1>/FROM ;
  wire N139826;
  wire \DLX_IDinst_branch_address<2>/FROM ;
  wire N139889;
  wire \N163278/FROM ;
  wire \N163278/GROM ;
  wire \DLX_EXinst_Mshift__n0024_Sh<50>/FROM ;
  wire \DLX_EXinst_Mshift__n0024_Sh<50>/GROM ;
  wire \DLX_IDinst_branch_address<3>/FROM ;
  wire N139952;
  wire \DLX_IDinst_branch_address<4>/FROM ;
  wire N140015;
  wire \N163447/FROM ;
  wire \N163447/GROM ;
  wire \N163262/FROM ;
  wire \N163262/GROM ;
  wire \DLX_IDinst_EPC<0>/FROM ;
  wire N140078;
  wire \DLX_IDinst_branch_address<6>/FROM ;
  wire N145997;
  wire \DLX_IDinst_branch_address<7>/FROM ;
  wire N140126;
  wire \DLX_IDinst_branch_address<8>/FROM ;
  wire N140193;
  wire \DLX_IDinst_branch_address<9>/FROM ;
  wire N140256;
  wire \N163622/FROM ;
  wire \N163622/GROM ;
  wire \N163588/FROM ;
  wire \N163588/GROM ;
  wire \DLX_IDinst_counter<0>/FROM ;
  wire N144314;
  wire \N163456/FROM ;
  wire \N163456/GROM ;
  wire \N163477/FROM ;
  wire \N163477/GROM ;
  wire \N163465/FROM ;
  wire \N163465/GROM ;
  wire \N163452/FROM ;
  wire \N163452/GROM ;
  wire \N131077/FROM ;
  wire \N131077/GROM ;
  wire \DLX_IDinst_Cause_Reg<10>/FROM ;
  wire \DLX_IDinst_Cause_Reg<10>/GROM ;
  wire \DLX_IDinst_Cause_Reg<11>/FROM ;
  wire \DLX_IDinst_Cause_Reg<11>/GROM ;
  wire \DLX_IDinst_Cause_Reg<12>/FROM ;
  wire \DLX_IDinst_Cause_Reg<12>/GROM ;
  wire \DLX_IDinst_Cause_Reg<13>/FROM ;
  wire \DLX_IDinst_Cause_Reg<13>/GROM ;
  wire \DLX_IDinst_Cause_Reg<14>/FROM ;
  wire \DLX_IDinst_Cause_Reg<14>/GROM ;
  wire \DLX_IDinst_Cause_Reg<15>/FROM ;
  wire \DLX_IDinst_Cause_Reg<15>/GROM ;
  wire \DLX_IDinst_Cause_Reg<31>/FROM ;
  wire \DLX_IDinst_Cause_Reg<31>/GROM ;
  wire \DLX_EXinst_Mshift__n0019_Sh<23>/FROM ;
  wire \DLX_EXinst_Mshift__n0019_Sh<23>/GROM ;
  wire \vga_top_vga1_helpcounter<0>/BXMUXNOT ;
  wire \N163737/FROM ;
  wire \N163737/GROM ;
  wire \N163550/FROM ;
  wire \N163550/GROM ;
  wire \N163178/FROM ;
  wire \N163178/GROM ;
  wire \N163668/GROM ;
  wire \N163643/FROM ;
  wire \N163643/GROM ;
  wire \DLX_EXinst_N73013/FROM ;
  wire \DLX_EXinst_N73013/GROM ;
  wire \DLX_EXinst_N73424/FROM ;
  wire \DLX_EXinst_N73424/GROM ;
  wire \CHOICE1907/FROM ;
  wire \CHOICE1907/GROM ;
  wire \CHOICE1921/FROM ;
  wire \CHOICE1921/GROM ;
  wire \CHOICE1963/FROM ;
  wire \CHOICE1963/GROM ;
  wire \DLX_MEMinst_reg_dst_out<0>/FROM ;
  wire \DLX_MEMinst_reg_dst_out<0>/GROM ;
  wire \DLX_MEMinst_reg_dst_out<1>/FROM ;
  wire \DLX_MEMinst_reg_dst_out<1>/GROM ;
  wire \DLX_MEMinst_reg_dst_out<2>/FROM ;
  wire \DLX_MEMinst_reg_dst_out<2>/GROM ;
  wire \CHOICE3122/FROM ;
  wire \CHOICE3122/GROM ;
  wire \DLX_EXinst_N76388/FROM ;
  wire \DLX_EXinst_N76388/GROM ;
  wire \DLX_MEMinst_reg_dst_out<3>/FROM ;
  wire \DLX_MEMinst_reg_dst_out<3>/GROM ;
  wire \DLX_MEMinst_reg_dst_out<4>/LOGIC_ZERO ;
  wire DLX_IDinst_Mcompar__n0368_inst_lut4_42;
  wire \DLX_MEMinst_reg_dst_out<4>/CYMUXF ;
  wire \DLX_MEMinst_reg_dst_out<4>/CYINIT ;
  wire \CHOICE1870/FROM ;
  wire \CHOICE1870/GROM ;
  wire \CHOICE2053/FROM ;
  wire \CHOICE2053/GROM ;
  wire \N164172/FROM ;
  wire \N164172/GROM ;
  wire \CHOICE1280/FROM ;
  wire \CHOICE1280/GROM ;
  wire \N139189/FROM ;
  wire \N139189/GROM ;
  wire \N136960/FROM ;
  wire \N136960/GROM ;
  wire \CHOICE2945/FROM ;
  wire \CHOICE2945/GROM ;
  wire \DLX_EXinst_reg_out_B_EX<26>/GROM ;
  wire \CHOICE3615/FROM ;
  wire \CHOICE3615/GROM ;
  wire \N134683/FROM ;
  wire \N134683/GROM ;
  wire \DLX_EXinst_reg_out_B_EX<18>/GROM ;
  wire \N139297/FROM ;
  wire \N139297/GROM ;
  wire \CHOICE3081/FROM ;
  wire \CHOICE3081/GROM ;
  wire \CHOICE3091/FROM ;
  wire \CHOICE3091/GROM ;
  wire \CHOICE1295/FROM ;
  wire \CHOICE1295/GROM ;
  wire \CHOICE2020/FROM ;
  wire \CHOICE2020/GROM ;
  wire \DLX_EXinst_N73549/FROM ;
  wire \DLX_EXinst_N73549/GROM ;
  wire \DLX_IDinst_Mmux__COND_4_inst_lut4_54/FROM ;
  wire \DLX_IDinst_Mmux__COND_4_inst_lut4_54/GROM ;
  wire \DLX_IDinst_Mmux__COND_4_inst_lut4_53/FROM ;
  wire \DLX_IDinst_Mmux__COND_4_inst_lut4_53/GROM ;
  wire \CHOICE2025/FROM ;
  wire \CHOICE2025/GROM ;
  wire \N139405/FROM ;
  wire \N139405/GROM ;
  wire \DLX_IDinst_Mmux__COND_4_inst_lut4_49/FROM ;
  wire \DLX_IDinst_Mmux__COND_4_inst_lut4_49/GROM ;
  wire \DLX_IDinst_Mmux__COND_4_inst_lut4_48/FROM ;
  wire \DLX_IDinst_Mmux__COND_4_inst_lut4_48/GROM ;
  wire \DLX_EXinst_N73058/FROM ;
  wire \DLX_EXinst_N73058/GROM ;
  wire \N163506/FROM ;
  wire \N163506/GROM ;
  wire \N139100/FROM ;
  wire \N139100/GROM ;
  wire \DLX_IDinst_Mmux__COND_4_inst_lut4_47/FROM ;
  wire \DLX_IDinst_Mmux__COND_4_inst_lut4_47/GROM ;
  wire \DLX_IDinst_rt_addr<4>/GROM ;
  wire \CHOICE1888/FROM ;
  wire \CHOICE1888/GROM ;
  wire \CHOICE1939/FROM ;
  wire \CHOICE1939/GROM ;
  wire \DLX_EXinst_ALU_result<31>/FROM ;
  wire CHOICE5867;
  wire \N163246/FROM ;
  wire \N163246/GROM ;
  wire \N147200/FROM ;
  wire \N147200/GROM ;
  wire \DLX_IDinst__n0381/FROM ;
  wire \DLX_IDinst__n0381/GROM ;
  wire \CHOICE1348/FROM ;
  wire \CHOICE1348/GROM ;
  wire \vga_top_vga1_videoon/FROM ;
  wire \vga_top_vga1_videoon/GROM ;
  wire \vga_top_vga1_videoon/LOGIC_ONE ;
  wire \N163534/FROM ;
  wire \N163534/GROM ;
  wire \DLX_IDinst_Ker1084541_1/FROM ;
  wire \DLX_IDinst_Ker1084541_1/GROM ;
  wire \N163602/FROM ;
  wire \N163602/GROM ;
  wire \DM_read_data<9>/FROM ;
  wire \DM_read_data<9>/GROM ;
  wire \N163627/FROM ;
  wire \N163627/GROM ;
  wire \N163692/FROM ;
  wire \N163692/GROM ;
  wire \DLX_IDinst_EPC<1>/FROM ;
  wire \DLX_IDinst_EPC<1>/GROM ;
  wire \DLX_IDinst_EPC<7>/FROM ;
  wire \DLX_IDinst_EPC<7>/GROM ;
  wire \DLX_IDinst_EPC<8>/FROM ;
  wire \DLX_IDinst_EPC<8>/GROM ;
  wire \DLX_EXinst_ALU_result<1>/FROM ;
  wire \DLX_EXinst_ALU_result<1>/GROM ;
  wire \vga_top_vga1_N112931/FROM ;
  wire \vga_top_vga1_N112931/GROM ;
  wire \N163407/FROM ;
  wire \N163407/GROM ;
  wire \DLX_IDinst_rd_addr<0>/FROM ;
  wire \DLX_IDinst_rd_addr<1>/FROM ;
  wire \DLX_IDinst_Imm<5>/FROM ;
  wire DLX_IDinst__n0129;
  wire \DLX_IDinst_rd_addr<2>/FROM ;
  wire \DLX_EXinst_N76002/FROM ;
  wire \DLX_EXinst_N76002/GROM ;
  wire \DLX_EXinst_N73897/FROM ;
  wire \DLX_EXinst_N73897/GROM ;
  wire \DLX_EXinst_N73267/FROM ;
  wire \DLX_EXinst_N73267/GROM ;
  wire \DLX_EXinst_N72803/FROM ;
  wire \DLX_EXinst_N72803/GROM ;
  wire \DLX_EXinst_N73604/FROM ;
  wire \DLX_EXinst_N73604/GROM ;
  wire \DLX_EXinst_N73524/FROM ;
  wire \DLX_EXinst_N73524/GROM ;
  wire \DLX_EXinst_N74245/FROM ;
  wire \DLX_EXinst_N74245/GROM ;
  wire \DLX_EXinst_N73554/FROM ;
  wire \DLX_EXinst_N73554/GROM ;
  wire \DLX_EXinst_N73509/FROM ;
  wire \DLX_EXinst_N73509/GROM ;
  wire \DLX_EXinst_N72822/FROM ;
  wire \DLX_EXinst_N72822/GROM ;
  wire \DLX_EXinst_N72710/FROM ;
  wire \DLX_EXinst_N72710/GROM ;
  wire \DLX_EXinst_N73464/FROM ;
  wire \DLX_EXinst_N73464/GROM ;
  wire \DLX_EXinst_N73519/FROM ;
  wire \DLX_EXinst_N73519/GROM ;
  wire \DLX_EXinst_N72815/FROM ;
  wire \DLX_EXinst_N72815/GROM ;
  wire \DLX_EXinst_N73544/FROM ;
  wire \DLX_EXinst_N73544/GROM ;
  wire \DLX_EXinst_N73384/FROM ;
  wire \DLX_EXinst_N73384/GROM ;
  wire \DLX_EXinst_N72809/FROM ;
  wire \DLX_EXinst_N72809/GROM ;
  wire \DLX_EXinst_N73529/FROM ;
  wire \DLX_EXinst_N73529/GROM ;
  wire \DLX_EXinst_N73369/FROM ;
  wire \DLX_EXinst_N73369/GROM ;
  wire \DLX_EXinst_N73474/FROM ;
  wire \DLX_EXinst_N73474/GROM ;
  wire \DLX_EXinst_N73394/FROM ;
  wire \DLX_EXinst_N73394/GROM ;
  wire \DLX_EXinst_reg_out_B_EX<0>/FROM ;
  wire \DLX_EXinst_N73539/FROM ;
  wire \DLX_EXinst_N73539/GROM ;
  wire \DLX_EXinst_N76011/FROM ;
  wire \DLX_EXinst_N76011/GROM ;
  wire \DLX_EXinst_N73379/GROM ;
  wire \DLX_EXinst_N73564/FROM ;
  wire \DLX_EXinst_N73564/GROM ;
  wire \DLX_EXinst_N74196/FROM ;
  wire \DLX_EXinst_N74196/GROM ;
  wire \DLX_EXinst_N73579/FROM ;
  wire \DLX_EXinst_N73579/GROM ;
  wire \DLX_EXinst_N72853/FROM ;
  wire \DLX_EXinst_N72853/GROM ;
  wire \DLX_EXinst_N73389/FROM ;
  wire \DLX_EXinst_N73389/GROM ;
  wire \DLX_EXinst_N73469/FROM ;
  wire \DLX_EXinst_N73469/GROM ;
  wire \DLX_EXinst_N73494/FROM ;
  wire \DLX_EXinst_N73494/GROM ;
  wire \DLX_EXinst_N73574/FROM ;
  wire \DLX_EXinst_N73574/GROM ;
  wire \DLX_EXinst_N74686/FROM ;
  wire \DLX_EXinst_N74686/GROM ;
  wire \DLX_EXinst_N72943/FROM ;
  wire \DLX_EXinst_N72943/GROM ;
  wire \DLX_EXinst_N72863/FROM ;
  wire \DLX_EXinst_N72863/GROM ;
  wire \DLX_EXinst_N73399/FROM ;
  wire \DLX_EXinst_N73399/GROM ;
  wire \DLX_EXinst_word/FROM ;
  wire DLX_EXinst__n0011;
  wire \DLX_EXinst_N73479/FROM ;
  wire \DLX_EXinst_N73479/GROM ;
  wire \DLX_EXinst_N73559/FROM ;
  wire \DLX_EXinst_N73559/GROM ;
  wire DLX_EXinst__n0010;
  wire \DLX_EXinst_byte/GROM ;
  wire \DLX_EXinst_N73584/FROM ;
  wire \DLX_EXinst_N73584/GROM ;
  wire \DLX_EXinst_N72873/FROM ;
  wire \DLX_EXinst_N72873/GROM ;
  wire \DLX_EXinst_N73569/FROM ;
  wire \DLX_EXinst_N73569/GROM ;
  wire \DLX_EXinst_N73489/FROM ;
  wire \DLX_EXinst_N73489/GROM ;
  wire \DLX_EXinst_N74201/FROM ;
  wire \DLX_EXinst_N74201/GROM ;
  wire \DLX_EXinst_N76041/FROM ;
  wire \DLX_EXinst_N76041/GROM ;
  wire \DLX_EXinst_N72858/FROM ;
  wire \DLX_EXinst_N72858/GROM ;
  wire \DLX_EXinst_N75139/FROM ;
  wire \DLX_EXinst_N75139/GROM ;
  wire \DLX_EXinst_N72963/FROM ;
  wire \DLX_EXinst_N72963/GROM ;
  wire \DLX_EXinst_N72883/FROM ;
  wire \DLX_EXinst_N72883/GROM ;
  wire \DLX_EXinst_N72948/FROM ;
  wire \DLX_EXinst_N72948/GROM ;
  wire \DLX_EXinst_N72888/FROM ;
  wire \DLX_EXinst_N72888/GROM ;
  wire \DLX_EXinst_N72797/FROM ;
  wire \DLX_EXinst_N72797/GROM ;
  wire \DLX_EXinst_N73589/FROM ;
  wire \DLX_EXinst_N73589/GROM ;
  wire \DLX_EXinst_N76318/FROM ;
  wire \DLX_EXinst_N76318/GROM ;
  wire \DLX_EXinst_N72958/FROM ;
  wire \DLX_EXinst_N72958/GROM ;
  wire \DLX_EXinst_N72878/FROM ;
  wire \DLX_EXinst_N72878/GROM ;
  wire \DLX_EXinst_N72791/FROM ;
  wire \DLX_EXinst_N72791/GROM ;
  wire \DLX_EXinst_N72968/FROM ;
  wire \DLX_EXinst_N72968/GROM ;
  wire \CHOICE2103/GROM ;
  wire \DLX_EXinst_N74991/FROM ;
  wire \DLX_EXinst_N74991/GROM ;
  wire \DLX_EXinst_N76338/FROM ;
  wire \DLX_EXinst_N76338/GROM ;
  wire \DLX_EXinst_N72898/FROM ;
  wire \DLX_EXinst_N72898/GROM ;
  wire \DLX_EXinst_N73848/FROM ;
  wire \DLX_EXinst_N73848/GROM ;
  wire \DLX_EXinst_N76285/GROM ;
  wire \DLX_EXinst_N76431/FROM ;
  wire \DLX_EXinst_N76431/GROM ;
  wire \DLX_EXinst_ALU_result<9>/FROM ;
  wire \DLX_EXinst_ALU_result<9>/GROM ;
  wire \DLX_EXinst_N76463/FROM ;
  wire \DLX_EXinst_N76463/GROM ;
  wire \DLX_EXinst_N74701/FROM ;
  wire \DLX_EXinst_N74701/GROM ;
  wire \CHOICE2119/FROM ;
  wire \CHOICE2119/GROM ;
  wire \DLX_EXinst_N76457/FROM ;
  wire \DLX_EXinst_N76457/GROM ;
  wire \DLX_EXinst_N76473/FROM ;
  wire \DLX_EXinst_N76473/GROM ;
  wire \DLX_EXinst_N74681/GROM ;
  wire \DLX_EXinst_N74711/FROM ;
  wire \DLX_EXinst_N74711/GROM ;
  wire \N139656/GROM ;
  wire \DLX_EXinst_N74951/GROM ;
  wire \DLX_EXinst_N76496/FROM ;
  wire \DLX_EXinst_N76496/GROM ;
  wire \DLX_EXinst_N76490/FROM ;
  wire \DLX_EXinst_N76490/GROM ;
  wire \DLX_EXinst_N74971/FROM ;
  wire \DLX_EXinst_N74971/GROM ;
  wire \N164607/FROM ;
  wire \N164607/GROM ;
  wire \DLX_EXinst_N75993/FROM ;
  wire \DLX_EXinst_N75993/GROM ;
  wire \N134590/FROM ;
  wire \N134590/GROM ;
  wire \CHOICE3386/FROM ;
  wire \CHOICE3386/GROM ;
  wire \CHOICE3301/FROM ;
  wire \CHOICE3301/GROM ;
  wire \DLX_EXinst_Mcompar__n0069_inst_cy_261/FROM ;
  wire \DLX_EXinst_Mcompar__n0069_inst_cy_261/GROM ;
  wire \CHOICE1326/FROM ;
  wire \CHOICE1326/GROM ;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_229/FROM ;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_229/GROM ;
  wire \CHOICE1693/FROM ;
  wire \CHOICE1693/GROM ;
  wire \DLX_EXinst_ALU_result<2>/FROM ;
  wire \DLX_EXinst_ALU_result<2>/GROM ;
  wire \N132148/FROM ;
  wire \N132148/GROM ;
  wire \DLX_IDinst_mem_write/FROM ;
  wire DLX_IDinst__n0141;
  wire \N163222/GROM ;
  wire \DLX_IDinst_mem_to_reg/FROM ;
  wire DLX_IDinst__n0139;
  wire \N164089/FROM ;
  wire \N164089/GROM ;
  wire \DLX_EXinst_N74130/FROM ;
  wire \DLX_EXinst_N74130/GROM ;
  wire \DLX_EXinst_N73287/FROM ;
  wire \DLX_EXinst_N73287/GROM ;
  wire \DLX_EXinst_reg_out_B_EX<2>/FROM ;
  wire \N132193/FROM ;
  wire \N132193/GROM ;
  wire \DLX_EXinst_N74625/FROM ;
  wire \DLX_EXinst_N74625/GROM ;
  wire \DLX_IDinst_RegFile_10_11/FROM ;
  wire \DLX_IDinst_RegFile_10_11/GROM ;
  wire \DLX_IDinst_RegFile_10_12/FROM ;
  wire \DLX_IDinst_RegFile_10_12/GROM ;
  wire \DLX_IDinst_RegFile_10_13/FROM ;
  wire \DLX_IDinst_RegFile_10_13/GROM ;
  wire \DLX_IDinst_RegFile_10_14/FROM ;
  wire \DLX_IDinst_RegFile_10_14/GROM ;
  wire \DLX_IDinst_RegFile_10_15/FROM ;
  wire \DLX_IDinst_RegFile_10_15/GROM ;
  wire \DLX_IDinst_RegFile_0_8/FROM ;
  wire \DLX_IDinst_RegFile_0_8/GROM ;
  wire \N164094/FROM ;
  wire \N164094/GROM ;
  wire \DLX_IDinst_RegFile_0_9/FROM ;
  wire \DLX_IDinst_RegFile_0_9/GROM ;
  wire \DLX_IDinst_RegFile_10_10/FROM ;
  wire \DLX_IDinst_RegFile_10_10/GROM ;
  wire \N132252/FROM ;
  wire \N132252/GROM ;
  wire \DLX_EXinst_ALU_result<3>/FROM ;
  wire \DLX_EXinst_ALU_result<3>/GROM ;
  wire \N131191/FROM ;
  wire \N131191/GROM ;
  wire \N131255/FROM ;
  wire \N131255/GROM ;
  wire \N131315/FROM ;
  wire \N131315/GROM ;
  wire \N130105/FROM ;
  wire \N130105/GROM ;
  wire \N130157/FROM ;
  wire \N130157/GROM ;
  wire \DLX_EXinst_Mshift__n0021_Sh<2>/FROM ;
  wire \DLX_EXinst_Mshift__n0021_Sh<2>/GROM ;
  wire \DLX_EXinst_Mshift__n0021_Sh<7>/FROM ;
  wire \DLX_EXinst_Mshift__n0021_Sh<7>/GROM ;
  wire \DLX_EXinst_opcode_of_EX_reg<0>/FROM ;
  wire \DLX_EXinst_opcode_of_EX_reg<0>/GROM ;
  wire \DLX_EXinst_opcode_of_EX_reg<1>/FROM ;
  wire \DLX_EXinst_opcode_of_EX_reg<1>/GROM ;
  wire \DLX_EXinst_opcode_of_EX_reg<2>/FROM ;
  wire \DLX_EXinst_opcode_of_EX_reg<2>/GROM ;
  wire \DLX_EXinst_opcode_of_EX_reg<3>/FROM ;
  wire \DLX_EXinst_opcode_of_EX_reg<3>/GROM ;
  wire \DLX_EXinst_opcode_of_EX_reg<4>/FROM ;
  wire \DLX_EXinst_opcode_of_EX_reg<4>/GROM ;
  wire \DM_write/ENABLE ;
  wire \DM_write/TORGTS ;
  wire \DM_write/OUTMUX ;
  wire DLX_EXinst_mem_write_EX_1;
  wire \DM_write/OD ;
  wire \CLI/ENABLE ;
  wire \CLI/TORGTS ;
  wire \CLI/OUTMUX ;
  wire DLX_IDinst_CLI_1;
  wire \CLI/OD ;
  wire \INT/IBUF ;
  wire \NPC_eff<0>/ENABLE ;
  wire \NPC_eff<0>/TORGTS ;
  wire \NPC_eff<0>/OUTMUX ;
  wire DLX_IFinst_NPC_0_1;
  wire \NPC_eff<0>/OD ;
  wire \NPC_eff<1>/ENABLE ;
  wire \NPC_eff<1>/TORGTS ;
  wire \NPC_eff<1>/OUTMUX ;
  wire DLX_IFinst_NPC_1_1;
  wire \NPC_eff<1>/OD ;
  wire \NPC_eff<2>/ENABLE ;
  wire \NPC_eff<2>/TORGTS ;
  wire \NPC_eff<2>/OUTMUX ;
  wire DLX_IFinst_NPC_2_1;
  wire \NPC_eff<2>/OD ;
  wire \NPC_eff<3>/ENABLE ;
  wire \NPC_eff<3>/TORGTS ;
  wire \NPC_eff<3>/OUTMUX ;
  wire DLX_IFinst_NPC_3_1;
  wire \NPC_eff<3>/OD ;
  wire \NPC_eff<4>/ENABLE ;
  wire \NPC_eff<4>/TORGTS ;
  wire \NPC_eff<4>/OUTMUX ;
  wire DLX_IFinst_NPC_4_1;
  wire \NPC_eff<4>/OD ;
  wire \NPC_eff<5>/ENABLE ;
  wire \NPC_eff<5>/TORGTS ;
  wire \NPC_eff<5>/OUTMUX ;
  wire DLX_IFinst_NPC_5_1;
  wire \NPC_eff<5>/OD ;
  wire \NPC_eff<6>/ENABLE ;
  wire \NPC_eff<6>/TORGTS ;
  wire \NPC_eff<6>/OUTMUX ;
  wire DLX_IFinst_NPC_6_1;
  wire \NPC_eff<6>/OD ;
  wire \NPC_eff<7>/ENABLE ;
  wire \NPC_eff<7>/TORGTS ;
  wire \NPC_eff<7>/OUTMUX ;
  wire DLX_IFinst_NPC_7_1;
  wire \NPC_eff<7>/OD ;
  wire \NPC_eff<8>/ENABLE ;
  wire \NPC_eff<8>/TORGTS ;
  wire \NPC_eff<8>/OUTMUX ;
  wire DLX_IFinst_NPC_8_1;
  wire \NPC_eff<8>/OD ;
  wire \NPC_eff<9>/ENABLE ;
  wire \NPC_eff<9>/TORGTS ;
  wire \NPC_eff<9>/OUTMUX ;
  wire DLX_IFinst_NPC_9_1;
  wire \NPC_eff<9>/OD ;
  wire \mask<0>/ENABLE ;
  wire \mask<0>/TORGTS ;
  wire \mask<0>/OUTMUX ;
  wire \mask<3>/ENABLE ;
  wire \mask<3>/TORGTS ;
  wire \mask<3>/OUTMUX ;
  wire \NPC_eff<10>/ENABLE ;
  wire \NPC_eff<10>/TORGTS ;
  wire \NPC_eff<10>/OUTMUX ;
  wire DLX_IFinst_NPC_10_1;
  wire \NPC_eff<10>/OD ;
  wire \NPC_eff<11>/ENABLE ;
  wire \NPC_eff<11>/TORGTS ;
  wire \NPC_eff<11>/OUTMUX ;
  wire DLX_IFinst_NPC_11_1;
  wire \NPC_eff<11>/OD ;
  wire \NPC_eff<12>/ENABLE ;
  wire \NPC_eff<12>/TORGTS ;
  wire \NPC_eff<12>/OUTMUX ;
  wire DLX_IFinst_NPC_12_1;
  wire \NPC_eff<12>/OD ;
  wire \NPC_eff<13>/ENABLE ;
  wire \NPC_eff<13>/TORGTS ;
  wire \NPC_eff<13>/OUTMUX ;
  wire DLX_IFinst_NPC_13_1;
  wire \NPC_eff<13>/OD ;
  wire \NPC_eff<14>/ENABLE ;
  wire \NPC_eff<14>/TORGTS ;
  wire \NPC_eff<14>/OUTMUX ;
  wire DLX_IFinst_NPC_14_1;
  wire \NPC_eff<14>/OD ;
  wire \NPC_eff<15>/ENABLE ;
  wire \NPC_eff<15>/TORGTS ;
  wire \NPC_eff<15>/OUTMUX ;
  wire DLX_IFinst_NPC_15_1;
  wire \NPC_eff<15>/OD ;
  wire \DM_write_data<0>/ENABLE ;
  wire \DM_write_data<0>/TORGTS ;
  wire \DM_write_data<0>/OUTMUX ;
  wire DLX_EXinst_reg_out_B_EX_0_1;
  wire \DM_write_data<0>/OD ;
  wire \blue<0>/ENABLE ;
  wire \blue<0>/TORGTS ;
  wire \blue<0>/OUTMUX ;
  wire \blue<1>/ENABLE ;
  wire \blue<1>/TORGTS ;
  wire \blue<1>/OUTMUX ;
  wire \blue<2>/ENABLE ;
  wire \blue<2>/TORGTS ;
  wire \blue<2>/OUTMUX ;
  wire \mask<1>/ENABLE ;
  wire \mask<1>/TORGTS ;
  wire \mask<1>/OUTMUX ;
  wire \mask<2>/ENABLE ;
  wire \mask<2>/TORGTS ;
  wire \mask<2>/OUTMUX ;
  wire \hsync/ENABLE ;
  wire \hsync/TORGTS ;
  wire \hsync/OUTMUX ;
  wire vga_top_vga1_hsyncout;
  wire \hsync/LOGIC_ZERO ;
  wire \reset/IBUF ;
  wire \stall/ENABLE ;
  wire \stall/TORGTS ;
  wire \stall/OUTMUX ;
  wire DLX_IDinst_stall_1;
  wire \stall/OD ;
  wire \vsync/ENABLE ;
  wire \vsync/TORGTS ;
  wire \vsync/OUTMUX ;
  wire vga_top_vga1_vsyncout;
  wire \vsync/LOGIC_ZERO ;
  wire \FREEZE/IBUF ;
  wire \branch_sig/ENABLE ;
  wire \branch_sig/TORGTS ;
  wire \branch_sig/OUTMUX ;
  wire DLX_IDinst_branch_sig_1;
  wire \branch_sig/OD ;
  wire \red<0>/ENABLE ;
  wire \red<0>/TORGTS ;
  wire \red<0>/OUTMUX ;
  wire \red<1>/ENABLE ;
  wire \red<1>/TORGTS ;
  wire \red<1>/OUTMUX ;
  wire \green<0>/ENABLE ;
  wire \green<0>/TORGTS ;
  wire \green<0>/OUTMUX ;
  wire \green<1>/ENABLE ;
  wire \green<1>/TORGTS ;
  wire \green<1>/OUTMUX ;
  wire \green<2>/ENABLE ;
  wire \green<2>/TORGTS ;
  wire \green<2>/OUTMUX ;
  wire \DM_addr_eff<10>/ENABLE ;
  wire \DM_addr_eff<10>/TORGTS ;
  wire \DM_addr_eff<10>/OUTMUX ;
  wire \DM_addr_eff<11>/ENABLE ;
  wire \DM_addr_eff<11>/TORGTS ;
  wire \DM_addr_eff<11>/OUTMUX ;
  wire \DM_addr_eff<12>/ENABLE ;
  wire \DM_addr_eff<12>/TORGTS ;
  wire \DM_addr_eff<12>/OUTMUX ;
  wire \DM_addr_eff<13>/ENABLE ;
  wire \DM_addr_eff<13>/TORGTS ;
  wire \DM_addr_eff<13>/OUTMUX ;
  wire \DM_addr_eff<14>/ENABLE ;
  wire \DM_addr_eff<14>/TORGTS ;
  wire \DM_addr_eff<14>/OUTMUX ;
  wire \DM_addr_eff<0>/ENABLE ;
  wire \DM_addr_eff<0>/TORGTS ;
  wire \DM_addr_eff<0>/OUTMUX ;
  wire \DM_addr_eff<1>/ENABLE ;
  wire \DM_addr_eff<1>/TORGTS ;
  wire \DM_addr_eff<1>/OUTMUX ;
  wire \DM_addr_eff<2>/ENABLE ;
  wire \DM_addr_eff<2>/TORGTS ;
  wire \DM_addr_eff<2>/OUTMUX ;
  wire \DM_addr_eff<3>/ENABLE ;
  wire \DM_addr_eff<3>/TORGTS ;
  wire \DM_addr_eff<3>/OUTMUX ;
  wire \DM_addr_eff<4>/ENABLE ;
  wire \DM_addr_eff<4>/TORGTS ;
  wire \DM_addr_eff<4>/OUTMUX ;
  wire \DM_addr_eff<5>/ENABLE ;
  wire \DM_addr_eff<5>/TORGTS ;
  wire \DM_addr_eff<5>/OUTMUX ;
  wire \DM_addr_eff<6>/ENABLE ;
  wire \DM_addr_eff<6>/TORGTS ;
  wire \DM_addr_eff<6>/OUTMUX ;
  wire \DM_addr_eff<7>/ENABLE ;
  wire \DM_addr_eff<7>/TORGTS ;
  wire \DM_addr_eff<7>/OUTMUX ;
  wire \DM_addr_eff<8>/ENABLE ;
  wire \DM_addr_eff<8>/TORGTS ;
  wire \DM_addr_eff<8>/OUTMUX ;
  wire \DM_addr_eff<9>/ENABLE ;
  wire \DM_addr_eff<9>/TORGTS ;
  wire \DM_addr_eff<9>/OUTMUX ;
  wire \PIPEEMPTY/ENABLE ;
  wire \PIPEEMPTY/TORGTS ;
  wire \PIPEEMPTY/OUTMUX ;
  wire \DM_read/ENABLE ;
  wire \DM_read/TORGTS ;
  wire \DM_read/OUTMUX ;
  wire DLX_EXinst_mem_read_EX;
  wire \DM_read/OD ;
  wire \IR_MSB<0>/ENABLE ;
  wire \IR_MSB<0>/TORGTS ;
  wire \IR_MSB<0>/OUTMUX ;
  wire \IR_MSB<1>/ENABLE ;
  wire \IR_MSB<1>/TORGTS ;
  wire \IR_MSB<1>/OUTMUX ;
  wire \IR_MSB<2>/ENABLE ;
  wire \IR_MSB<2>/TORGTS ;
  wire \IR_MSB<2>/OUTMUX ;
  wire \IR_MSB<3>/ENABLE ;
  wire \IR_MSB<3>/TORGTS ;
  wire \IR_MSB<3>/OUTMUX ;
  wire \IR_MSB<4>/ENABLE ;
  wire \IR_MSB<4>/TORGTS ;
  wire \IR_MSB<4>/OUTMUX ;
  wire \IR_MSB<5>/ENABLE ;
  wire \IR_MSB<5>/TORGTS ;
  wire \IR_MSB<5>/OUTMUX ;
  wire \IR_MSB<6>/ENABLE ;
  wire \IR_MSB<6>/TORGTS ;
  wire \IR_MSB<6>/OUTMUX ;
  wire \IR_MSB<7>/ENABLE ;
  wire \IR_MSB<7>/TORGTS ;
  wire \IR_MSB<7>/OUTMUX ;
  wire \clkdivider/LOCKED ;
  wire \clkdivider/CLK2X180 ;
  wire \clkdivider/CLK2X ;
  wire \clkdivider/CLK270 ;
  wire \clkdivider/CLK180 ;
  wire \clkdivider/CLK90 ;
  wire \clkdivider/LOGIC_ZERO ;
  wire \vga0/DOB15 ;
  wire \vga0/DOB14 ;
  wire \vga0/DOB13 ;
  wire \vga0/DOB12 ;
  wire \vga0/DOB11 ;
  wire \vga0/DOB10 ;
  wire \vga0/DOB9 ;
  wire \vga0/DOB8 ;
  wire \vga0/DOB7 ;
  wire \vga0/DOB6 ;
  wire \vga0/DOB5 ;
  wire \vga0/DOB4 ;
  wire \vga0/DOB3 ;
  wire \vga0/DOB2 ;
  wire \vga0/DOB1 ;
  wire \vga0/DOA15 ;
  wire \vga0/DOA14 ;
  wire \vga0/DOA13 ;
  wire \vga0/DOA12 ;
  wire \vga0/DOA11 ;
  wire \vga0/DOA10 ;
  wire \vga0/DOA9 ;
  wire \vga0/DOA8 ;
  wire \vga0/DOA7 ;
  wire \vga0/DOA6 ;
  wire \vga0/DOA5 ;
  wire \vga0/DOA4 ;
  wire \vga0/DOA3 ;
  wire \vga0/DOA2 ;
  wire \vga0/DOA1 ;
  wire \vga0/DIB15 ;
  wire \vga0/DIB14 ;
  wire \vga0/DIB13 ;
  wire \vga0/DIB12 ;
  wire \vga0/DIB11 ;
  wire \vga0/DIB10 ;
  wire \vga0/DIB9 ;
  wire \vga0/DIB8 ;
  wire \vga0/DIB7 ;
  wire \vga0/DIB6 ;
  wire \vga0/DIB5 ;
  wire \vga0/DIB4 ;
  wire \vga0/DIB3 ;
  wire \vga0/DIB2 ;
  wire \vga0/DIB1 ;
  wire \vga0/DIB0 ;
  wire \vga0/DIA15 ;
  wire \vga0/DIA14 ;
  wire \vga0/DIA13 ;
  wire \vga0/DIA12 ;
  wire \vga0/DIA11 ;
  wire \vga0/DIA10 ;
  wire \vga0/DIA9 ;
  wire \vga0/DIA8 ;
  wire \vga0/DIA7 ;
  wire \vga0/DIA6 ;
  wire \vga0/DIA5 ;
  wire \vga0/DIA4 ;
  wire \vga0/DIA3 ;
  wire \vga0/DIA2 ;
  wire \vga0/DIA1 ;
  wire \vga0/LOGIC_ZERO ;
  wire \vga0/LOGIC_ONE ;
  wire \vga0/CLKA_INTNOT ;
  wire \vga1/DOB15 ;
  wire \vga1/DOB14 ;
  wire \vga1/DOB13 ;
  wire \vga1/DOB12 ;
  wire \vga1/DOB11 ;
  wire \vga1/DOB10 ;
  wire \vga1/DOB9 ;
  wire \vga1/DOB8 ;
  wire \vga1/DOB7 ;
  wire \vga1/DOB6 ;
  wire \vga1/DOB5 ;
  wire \vga1/DOB4 ;
  wire \vga1/DOB3 ;
  wire \vga1/DOB2 ;
  wire \vga1/DOB1 ;
  wire \vga1/DOA15 ;
  wire \vga1/DOA14 ;
  wire \vga1/DOA13 ;
  wire \vga1/DOA12 ;
  wire \vga1/DOA11 ;
  wire \vga1/DOA10 ;
  wire \vga1/DOA9 ;
  wire \vga1/DOA8 ;
  wire \vga1/DOA7 ;
  wire \vga1/DOA6 ;
  wire \vga1/DOA5 ;
  wire \vga1/DOA4 ;
  wire \vga1/DOA3 ;
  wire \vga1/DOA2 ;
  wire \vga1/DOA1 ;
  wire \vga1/DIB15 ;
  wire \vga1/DIB14 ;
  wire \vga1/DIB13 ;
  wire \vga1/DIB12 ;
  wire \vga1/DIB11 ;
  wire \vga1/DIB10 ;
  wire \vga1/DIB9 ;
  wire \vga1/DIB8 ;
  wire \vga1/DIB7 ;
  wire \vga1/DIB6 ;
  wire \vga1/DIB5 ;
  wire \vga1/DIB4 ;
  wire \vga1/DIB3 ;
  wire \vga1/DIB2 ;
  wire \vga1/DIB1 ;
  wire \vga1/DIB0 ;
  wire \vga1/DIA15 ;
  wire \vga1/DIA14 ;
  wire \vga1/DIA13 ;
  wire \vga1/DIA12 ;
  wire \vga1/DIA11 ;
  wire \vga1/DIA10 ;
  wire \vga1/DIA9 ;
  wire \vga1/DIA8 ;
  wire \vga1/DIA7 ;
  wire \vga1/DIA6 ;
  wire \vga1/DIA5 ;
  wire \vga1/DIA4 ;
  wire \vga1/DIA3 ;
  wire \vga1/DIA2 ;
  wire \vga1/DIA1 ;
  wire \vga1/LOGIC_ZERO ;
  wire \vga1/LOGIC_ONE ;
  wire \vga1/CLKA_INTNOT ;
  wire \vga2/DOB15 ;
  wire \vga2/DOB14 ;
  wire \vga2/DOB13 ;
  wire \vga2/DOB12 ;
  wire \vga2/DOB11 ;
  wire \vga2/DOB10 ;
  wire \vga2/DOB9 ;
  wire \vga2/DOB8 ;
  wire \vga2/DOB7 ;
  wire \vga2/DOB6 ;
  wire \vga2/DOB5 ;
  wire \vga2/DOB4 ;
  wire \vga2/DOB3 ;
  wire \vga2/DOB2 ;
  wire \vga2/DOB1 ;
  wire \vga2/DOA15 ;
  wire \vga2/DOA14 ;
  wire \vga2/DOA13 ;
  wire \vga2/DOA12 ;
  wire \vga2/DOA11 ;
  wire \vga2/DOA10 ;
  wire \vga2/DOA9 ;
  wire \vga2/DOA8 ;
  wire \vga2/DOA7 ;
  wire \vga2/DOA6 ;
  wire \vga2/DOA5 ;
  wire \vga2/DOA4 ;
  wire \vga2/DOA3 ;
  wire \vga2/DOA2 ;
  wire \vga2/DOA1 ;
  wire \vga2/DIB15 ;
  wire \vga2/DIB14 ;
  wire \vga2/DIB13 ;
  wire \vga2/DIB12 ;
  wire \vga2/DIB11 ;
  wire \vga2/DIB10 ;
  wire \vga2/DIB9 ;
  wire \vga2/DIB8 ;
  wire \vga2/DIB7 ;
  wire \vga2/DIB6 ;
  wire \vga2/DIB5 ;
  wire \vga2/DIB4 ;
  wire \vga2/DIB3 ;
  wire \vga2/DIB2 ;
  wire \vga2/DIB1 ;
  wire \vga2/DIB0 ;
  wire \vga2/DIA15 ;
  wire \vga2/DIA14 ;
  wire \vga2/DIA13 ;
  wire \vga2/DIA12 ;
  wire \vga2/DIA11 ;
  wire \vga2/DIA10 ;
  wire \vga2/DIA9 ;
  wire \vga2/DIA8 ;
  wire \vga2/DIA7 ;
  wire \vga2/DIA6 ;
  wire \vga2/DIA5 ;
  wire \vga2/DIA4 ;
  wire \vga2/DIA3 ;
  wire \vga2/DIA2 ;
  wire \vga2/DIA1 ;
  wire \vga2/LOGIC_ZERO ;
  wire \vga2/LOGIC_ONE ;
  wire \vga2/CLKA_INTNOT ;
  wire \vga3/DOB15 ;
  wire \vga3/DOB14 ;
  wire \vga3/DOB13 ;
  wire \vga3/DOB12 ;
  wire \vga3/DOB11 ;
  wire \vga3/DOB10 ;
  wire \vga3/DOB9 ;
  wire \vga3/DOB8 ;
  wire \vga3/DOB7 ;
  wire \vga3/DOB6 ;
  wire \vga3/DOB5 ;
  wire \vga3/DOB4 ;
  wire \vga3/DOB3 ;
  wire \vga3/DOB2 ;
  wire \vga3/DOB1 ;
  wire \vga3/DOA15 ;
  wire \vga3/DOA14 ;
  wire \vga3/DOA13 ;
  wire \vga3/DOA12 ;
  wire \vga3/DOA11 ;
  wire \vga3/DOA10 ;
  wire \vga3/DOA9 ;
  wire \vga3/DOA8 ;
  wire \vga3/DOA7 ;
  wire \vga3/DOA6 ;
  wire \vga3/DOA5 ;
  wire \vga3/DOA4 ;
  wire \vga3/DOA3 ;
  wire \vga3/DOA2 ;
  wire \vga3/DOA1 ;
  wire \vga3/DIB15 ;
  wire \vga3/DIB14 ;
  wire \vga3/DIB13 ;
  wire \vga3/DIB12 ;
  wire \vga3/DIB11 ;
  wire \vga3/DIB10 ;
  wire \vga3/DIB9 ;
  wire \vga3/DIB8 ;
  wire \vga3/DIB7 ;
  wire \vga3/DIB6 ;
  wire \vga3/DIB5 ;
  wire \vga3/DIB4 ;
  wire \vga3/DIB3 ;
  wire \vga3/DIB2 ;
  wire \vga3/DIB1 ;
  wire \vga3/DIB0 ;
  wire \vga3/DIA15 ;
  wire \vga3/DIA14 ;
  wire \vga3/DIA13 ;
  wire \vga3/DIA12 ;
  wire \vga3/DIA11 ;
  wire \vga3/DIA10 ;
  wire \vga3/DIA9 ;
  wire \vga3/DIA8 ;
  wire \vga3/DIA7 ;
  wire \vga3/DIA6 ;
  wire \vga3/DIA5 ;
  wire \vga3/DIA4 ;
  wire \vga3/DIA3 ;
  wire \vga3/DIA2 ;
  wire \vga3/DIA1 ;
  wire \vga3/LOGIC_ZERO ;
  wire \vga3/LOGIC_ONE ;
  wire \vga3/CLKA_INTNOT ;
  wire \vga4/DOB15 ;
  wire \vga4/DOB14 ;
  wire \vga4/DOB13 ;
  wire \vga4/DOB12 ;
  wire \vga4/DOB11 ;
  wire \vga4/DOB10 ;
  wire \vga4/DOB9 ;
  wire \vga4/DOB8 ;
  wire \vga4/DOB7 ;
  wire \vga4/DOB6 ;
  wire \vga4/DOB5 ;
  wire \vga4/DOB4 ;
  wire \vga4/DOB3 ;
  wire \vga4/DOB2 ;
  wire \vga4/DOB1 ;
  wire \vga4/DOA15 ;
  wire \vga4/DOA14 ;
  wire \vga4/DOA13 ;
  wire \vga4/DOA12 ;
  wire \vga4/DOA11 ;
  wire \vga4/DOA10 ;
  wire \vga4/DOA9 ;
  wire \vga4/DOA8 ;
  wire \vga4/DOA7 ;
  wire \vga4/DOA6 ;
  wire \vga4/DOA5 ;
  wire \vga4/DOA4 ;
  wire \vga4/DOA3 ;
  wire \vga4/DOA2 ;
  wire \vga4/DOA1 ;
  wire \vga4/DIB15 ;
  wire \vga4/DIB14 ;
  wire \vga4/DIB13 ;
  wire \vga4/DIB12 ;
  wire \vga4/DIB11 ;
  wire \vga4/DIB10 ;
  wire \vga4/DIB9 ;
  wire \vga4/DIB8 ;
  wire \vga4/DIB7 ;
  wire \vga4/DIB6 ;
  wire \vga4/DIB5 ;
  wire \vga4/DIB4 ;
  wire \vga4/DIB3 ;
  wire \vga4/DIB2 ;
  wire \vga4/DIB1 ;
  wire \vga4/DIB0 ;
  wire \vga4/DIA15 ;
  wire \vga4/DIA14 ;
  wire \vga4/DIA13 ;
  wire \vga4/DIA12 ;
  wire \vga4/DIA11 ;
  wire \vga4/DIA10 ;
  wire \vga4/DIA9 ;
  wire \vga4/DIA8 ;
  wire \vga4/DIA7 ;
  wire \vga4/DIA6 ;
  wire \vga4/DIA5 ;
  wire \vga4/DIA4 ;
  wire \vga4/DIA3 ;
  wire \vga4/DIA2 ;
  wire \vga4/DIA1 ;
  wire \vga4/LOGIC_ZERO ;
  wire \vga4/LOGIC_ONE ;
  wire \vga4/CLKA_INTNOT ;
  wire \block0/DOB15 ;
  wire \block0/DOB14 ;
  wire \block0/DOB13 ;
  wire \block0/DOB12 ;
  wire \block0/DOB11 ;
  wire \block0/DOB10 ;
  wire \block0/DOB9 ;
  wire \block0/DOB8 ;
  wire \block0/DOA15 ;
  wire \block0/DOA14 ;
  wire \block0/DOA13 ;
  wire \block0/DOA12 ;
  wire \block0/DOA11 ;
  wire \block0/DOA10 ;
  wire \block0/DOA9 ;
  wire \block0/DOA8 ;
  wire \block0/DIB15 ;
  wire \block0/DIB14 ;
  wire \block0/DIB13 ;
  wire \block0/DIB12 ;
  wire \block0/DIB11 ;
  wire \block0/DIB10 ;
  wire \block0/DIB9 ;
  wire \block0/DIB8 ;
  wire \block0/DIB7 ;
  wire \block0/DIB6 ;
  wire \block0/DIB5 ;
  wire \block0/DIB4 ;
  wire \block0/DIB3 ;
  wire \block0/DIB2 ;
  wire \block0/DIB1 ;
  wire \block0/DIB0 ;
  wire \block0/DIA15 ;
  wire \block0/DIA14 ;
  wire \block0/DIA13 ;
  wire \block0/DIA12 ;
  wire \block0/DIA11 ;
  wire \block0/DIA10 ;
  wire \block0/DIA9 ;
  wire \block0/DIA8 ;
  wire \block0/ADDRB2 ;
  wire \block0/ADDRB1 ;
  wire \block0/ADDRB0 ;
  wire \block0/ADDRA2 ;
  wire \block0/ADDRA1 ;
  wire \block0/ADDRA0 ;
  wire \block0/LOGIC_ZERO ;
  wire \block0/LOGIC_ONE ;
  wire \block0/CLKA_INTNOT ;
  wire \block1/DOB15 ;
  wire \block1/DOB14 ;
  wire \block1/DOB13 ;
  wire \block1/DOB12 ;
  wire \block1/DOB11 ;
  wire \block1/DOB10 ;
  wire \block1/DOB9 ;
  wire \block1/DOB8 ;
  wire \block1/DOA15 ;
  wire \block1/DOA14 ;
  wire \block1/DOA13 ;
  wire \block1/DOA12 ;
  wire \block1/DOA11 ;
  wire \block1/DOA10 ;
  wire \block1/DOA9 ;
  wire \block1/DOA8 ;
  wire \block1/DIB15 ;
  wire \block1/DIB14 ;
  wire \block1/DIB13 ;
  wire \block1/DIB12 ;
  wire \block1/DIB11 ;
  wire \block1/DIB10 ;
  wire \block1/DIB9 ;
  wire \block1/DIB8 ;
  wire \block1/DIB7 ;
  wire \block1/DIB6 ;
  wire \block1/DIB5 ;
  wire \block1/DIB4 ;
  wire \block1/DIB3 ;
  wire \block1/DIB2 ;
  wire \block1/DIB1 ;
  wire \block1/DIB0 ;
  wire \block1/DIA15 ;
  wire \block1/DIA14 ;
  wire \block1/DIA13 ;
  wire \block1/DIA12 ;
  wire \block1/DIA11 ;
  wire \block1/DIA10 ;
  wire \block1/DIA9 ;
  wire \block1/DIA8 ;
  wire \block1/ADDRB2 ;
  wire \block1/ADDRB1 ;
  wire \block1/ADDRB0 ;
  wire \block1/ADDRA2 ;
  wire \block1/ADDRA1 ;
  wire \block1/ADDRA0 ;
  wire \block1/LOGIC_ZERO ;
  wire \block1/LOGIC_ONE ;
  wire \block1/CLKA_INTNOT ;
  wire \block2/DOB15 ;
  wire \block2/DOB14 ;
  wire \block2/DOB13 ;
  wire \block2/DOB12 ;
  wire \block2/DOB11 ;
  wire \block2/DOB10 ;
  wire \block2/DOB9 ;
  wire \block2/DOB8 ;
  wire \block2/DOA15 ;
  wire \block2/DOA14 ;
  wire \block2/DOA13 ;
  wire \block2/DOA12 ;
  wire \block2/DOA11 ;
  wire \block2/DOA10 ;
  wire \block2/DOA9 ;
  wire \block2/DOA8 ;
  wire \block2/DIB15 ;
  wire \block2/DIB14 ;
  wire \block2/DIB13 ;
  wire \block2/DIB12 ;
  wire \block2/DIB11 ;
  wire \block2/DIB10 ;
  wire \block2/DIB9 ;
  wire \block2/DIB8 ;
  wire \block2/DIB7 ;
  wire \block2/DIB6 ;
  wire \block2/DIB5 ;
  wire \block2/DIB4 ;
  wire \block2/DIB3 ;
  wire \block2/DIB2 ;
  wire \block2/DIB1 ;
  wire \block2/DIB0 ;
  wire \block2/DIA15 ;
  wire \block2/DIA14 ;
  wire \block2/DIA13 ;
  wire \block2/DIA12 ;
  wire \block2/DIA11 ;
  wire \block2/DIA10 ;
  wire \block2/DIA9 ;
  wire \block2/DIA8 ;
  wire \block2/ADDRB2 ;
  wire \block2/ADDRB1 ;
  wire \block2/ADDRB0 ;
  wire \block2/ADDRA2 ;
  wire \block2/ADDRA1 ;
  wire \block2/ADDRA0 ;
  wire \block2/LOGIC_ZERO ;
  wire \block2/LOGIC_ONE ;
  wire \block2/CLKA_INTNOT ;
  wire \block3/DOB15 ;
  wire \block3/DOB14 ;
  wire \block3/DOB13 ;
  wire \block3/DOB12 ;
  wire \block3/DOB11 ;
  wire \block3/DOB10 ;
  wire \block3/DOB9 ;
  wire \block3/DOB8 ;
  wire \block3/DOA15 ;
  wire \block3/DOA14 ;
  wire \block3/DOA13 ;
  wire \block3/DOA12 ;
  wire \block3/DOA11 ;
  wire \block3/DOA10 ;
  wire \block3/DOA9 ;
  wire \block3/DOA8 ;
  wire \block3/DIB15 ;
  wire \block3/DIB14 ;
  wire \block3/DIB13 ;
  wire \block3/DIB12 ;
  wire \block3/DIB11 ;
  wire \block3/DIB10 ;
  wire \block3/DIB9 ;
  wire \block3/DIB8 ;
  wire \block3/DIB7 ;
  wire \block3/DIB6 ;
  wire \block3/DIB5 ;
  wire \block3/DIB4 ;
  wire \block3/DIB3 ;
  wire \block3/DIB2 ;
  wire \block3/DIB1 ;
  wire \block3/DIB0 ;
  wire \block3/DIA15 ;
  wire \block3/DIA14 ;
  wire \block3/DIA13 ;
  wire \block3/DIA12 ;
  wire \block3/DIA11 ;
  wire \block3/DIA10 ;
  wire \block3/DIA9 ;
  wire \block3/DIA8 ;
  wire \block3/ADDRB2 ;
  wire \block3/ADDRB1 ;
  wire \block3/ADDRB0 ;
  wire \block3/ADDRA2 ;
  wire \block3/ADDRA1 ;
  wire \block3/ADDRA0 ;
  wire \block3/LOGIC_ZERO ;
  wire \block3/LOGIC_ONE ;
  wire \block3/CLKA_INTNOT ;
  wire N165608;
  wire N165606;
  wire \DLX_EXinst_Mshift__n0019_Sh<24>/F5MUX ;
  wire N165528;
  wire N165526;
  wire \DLX_EXinst_Mshift__n0019_Sh<25>/F5MUX ;
  wire N165338;
  wire N165336;
  wire \DLX_EXinst_Mshift__n0019_Sh<26>/F5MUX ;
  wire N165588;
  wire N165586;
  wire \DLX_EXinst_Mshift__n0019_Sh<28>/F5MUX ;
  wire N165513;
  wire N165511;
  wire \DLX_EXinst_Mshift__n0021_Sh<43>/F5MUX ;
  wire N165943;
  wire N165941;
  wire \DLX_EXinst_Mshift__n0022_Sh<59>/F5MUX ;
  wire N165773;
  wire N165771;
  wire \DLX_EXinst_Mshift__n0023_Sh<40>/F5MUX ;
  wire N165373;
  wire N165371;
  wire \DLX_EXinst_Mshift__n0021_Sh<3>/F5MUX ;
  wire N165333;
  wire N165331;
  wire \DLX_EXinst_Mshift__n0021_Sh<4>/F5MUX ;
  wire N165638;
  wire N165636;
  wire \DLX_EXinst_Mshift__n0021_Sh<5>/F5MUX ;
  wire N165343;
  wire N165341;
  wire \DLX_EXinst_Mshift__n0021_Sh<6>/F5MUX ;
  wire N165368;
  wire N165366;
  wire \CHOICE4135/F5MUX ;
  wire N165363;
  wire N165361;
  wire \CHOICE4070/F5MUX ;
  wire N165498;
  wire N165496;
  wire \CHOICE4721/F5MUX ;
  wire N165533;
  wire N165531;
  wire \CHOICE4005/F5MUX ;
  wire N165848;
  wire N165846;
  wire \CHOICE4729/F5MUX ;
  wire N165523;
  wire N165521;
  wire \CHOICE5896/F5MUX ;
  wire N165633;
  wire N165631;
  wire \CHOICE4573/F5MUX ;
  wire N165518;
  wire N165516;
  wire \CHOICE5791/F5MUX ;
  wire N165593;
  wire N165591;
  wire \CHOICE5378/F5MUX ;
  wire N165418;
  wire N165416;
  wire \CHOICE5999/F5MUX ;
  wire N165453;
  wire N165451;
  wire \CHOICE5220/F5MUX ;
  wire N165413;
  wire N165411;
  wire \CHOICE5299/F5MUX ;
  wire N165423;
  wire N165421;
  wire \CHOICE4866/F5MUX ;
  wire N165493;
  wire N165491;
  wire \CHOICE4792/F5MUX ;
  wire N165573;
  wire N165571;
  wire \DLX_EXinst_Mshift__n0019_Sh<27>/F5MUX ;
  wire N165918;
  wire N165916;
  wire \CHOICE4800/F5MUX ;
  wire N165788;
  wire N165786;
  wire \CHOICE5191/F5MUX ;
  wire N165683;
  wire N165681;
  wire \CHOICE4558/F5MUX ;
  wire N165623;
  wire N165621;
  wire \DLX_EXinst_Mshift__n0020_Sh<25>/F5MUX ;
  wire N165448;
  wire N165446;
  wire \DLX_EXinst_Mshift__n0020_Sh<26>/F5MUX ;
  wire N165473;
  wire N165471;
  wire \DLX_EXinst_Mshift__n0020_Sh<28>/F5MUX ;
  wire N165618;
  wire N165616;
  wire \DLX_EXinst_Mshift__n0023_Sh<3>/F5MUX ;
  wire N165603;
  wire N165601;
  wire \DLX_EXinst_Mshift__n0023_Sh<4>/F5MUX ;
  wire N165578;
  wire N165576;
  wire \DLX_EXinst_Mshift__n0023_Sh<5>/F5MUX ;
  wire N165823;
  wire N165821;
  wire \N163716/F5MUX ;
  wire N165403;
  wire N165401;
  wire \N163242/F5MUX ;
  wire N165783;
  wire N165781;
  wire N165768;
  wire N165766;
  wire N165748;
  wire N165746;
  wire N165728;
  wire N165726;
  wire N165723;
  wire N165721;
  wire N165693;
  wire N165691;
  wire N165703;
  wire N165701;
  wire N165798;
  wire N165796;
  wire N165738;
  wire N165736;
  wire N165743;
  wire N165741;
  wire N165468;
  wire N165466;
  wire \CHOICE1987/F5MUX ;
  wire N165548;
  wire N165546;
  wire \DLX_IDinst_N107405/F5MUX ;
  wire N165893;
  wire N165891;
  wire \N163338/F5MUX ;
  wire N165708;
  wire N165706;
  wire \CHOICE4498/F5MUX ;
  wire N165353;
  wire N165351;
  wire \CHOICE4438/F5MUX ;
  wire N165348;
  wire N165346;
  wire \CHOICE3813/F5MUX ;
  wire N165733;
  wire N165731;
  wire \CHOICE3758/F5MUX ;
  wire N165563;
  wire N165561;
  wire \DLX_IDinst_RegFile_3_12/F5MUX ;
  wire N165443;
  wire N165441;
  wire \CHOICE4754/F5MUX ;
  wire N165698;
  wire N165696;
  wire \CHOICE3703/F5MUX ;
  wire N165393;
  wire N165391;
  wire \CHOICE4102/F5MUX ;
  wire N165818;
  wire N165816;
  wire \CHOICE5838/F5MUX ;
  wire N165463;
  wire N165461;
  wire \CHOICE4037/F5MUX ;
  wire N165713;
  wire N165711;
  wire \CHOICE5864/F5MUX ;
  wire N165668;
  wire N165666;
  wire \CHOICE4608/F5MUX ;
  wire N165758;
  wire N165756;
  wire \DLX_IDinst_RegFile_2_31/F5MUX ;
  wire N165828;
  wire N165826;
  wire \CHOICE5648/F5MUX ;
  wire N165538;
  wire N165536;
  wire \DLX_IFinst_IR_previous<21>/F5MUX ;
  wire N165568;
  wire N165566;
  wire \CHOICE5258/F5MUX ;
  wire N165598;
  wire N165596;
  wire \DLX_IDinst_RegFile_1_4/F5MUX ;
  wire N165863;
  wire N165861;
  wire \CHOICE4874/F5MUX ;
  wire N165583;
  wire N165581;
  wire \DLX_IDinst_RegFile_10_0/F5MUX ;
  wire N165483;
  wire N165481;
  wire \CHOICE4825/F5MUX ;
  wire N165878;
  wire N165876;
  wire \DLX_EXinst_ALU_result_5_1/F5MUX ;
  wire N165843;
  wire N165841;
  wire \DLX_EXinst_ALU_result_6_1/F5MUX ;
  wire N165803;
  wire N165801;
  wire \DLX_EXinst_ALU_result_7_1/F5MUX ;
  wire N165438;
  wire N165436;
  wire \CHOICE1765/F5MUX ;
  wire N165628;
  wire N165626;
  wire \DLX_IDinst_RegFile_30_10/F5MUX ;
  wire N165488;
  wire N165486;
  wire \N137952/F5MUX ;
  wire N165478;
  wire N165476;
  wire \DLX_IFinst_IR_previous<24>/F5MUX ;
  wire N165378;
  wire N165376;
  wire \N134488/F5MUX ;
  wire N165933;
  wire N165931;
  wire \DLX_IDinst_RegFile_2_20/F5MUX ;
  wire N165558;
  wire N165556;
  wire \N137859/F5MUX ;
  wire N165503;
  wire N165501;
  wire \DLX_IDinst_RegFile_26_0/F5MUX ;
  wire N165658;
  wire N165656;
  wire \N138037/F5MUX ;
  wire N165508;
  wire N165506;
  wire \DLX_IDinst_RegFile_17_7/F5MUX ;
  wire N165958;
  wire N165956;
  wire \N137774/F5MUX ;
  wire N165543;
  wire N165541;
  wire \DLX_IDinst_RegFile_10_3/F5MUX ;
  wire N165408;
  wire N165406;
  wire \CHOICE1727/F5MUX ;
  wire N165673;
  wire N165671;
  wire \DLX_IDinst_RegFile_2_28/F5MUX ;
  wire N165663;
  wire N165661;
  wire \N134128/F5MUX ;
  wire N165428;
  wire N165426;
  wire \DLX_IFinst_IR_previous<1>/F5MUX ;
  wire N165383;
  wire N165381;
  wire \N133552/F5MUX ;
  wire N165898;
  wire N165896;
  wire \DLX_IDinst_RegFile_14_21/F5MUX ;
  wire N165868;
  wire N165866;
  wire \CHOICE2965/F5MUX ;
  wire N165388;
  wire N165386;
  wire \DLX_IFinst_IR_previous<4>/F5MUX ;
  wire N165358;
  wire N165356;
  wire \N133984/F5MUX ;
  wire N165458;
  wire N165456;
  wire \DLX_IDinst_RegFile_14_10/F5MUX ;
  wire N165643;
  wire N165641;
  wire \N133048/F5MUX ;
  wire N165653;
  wire N165651;
  wire \DLX_IDinst_RegFile_11_0/F5MUX ;
  wire N165613;
  wire N165611;
  wire \N133120/F5MUX ;
  wire N165948;
  wire N165946;
  wire \DLX_IDinst_RegFile_14_22/F5MUX ;
  wire N165688;
  wire N165686;
  wire \DM_read_data<0>/F5MUX ;
  wire \vram_out_vga_eff/LOGIC_ONE ;
  wire \vram_out_vga<4>_rt ;
  wire \vram_out_vga_eff/F6MUX ;
  wire \Mmux__COND_2_inst_mux_f6_0.F51 ;
  wire N165648;
  wire N165646;
  wire N162847;
  wire Mmux__COND_2__net1;
  wire Mmux__COND_2__net0;
  wire \Mmux__COND_2__net2/F5MUX ;
  wire N165953;
  wire N165951;
  wire \DLX_MEMinst_opcode_of_WB<3>/F5MUX ;
  wire N165928;
  wire N165926;
  wire N165793;
  wire N165791;
  wire N165923;
  wire N165921;
  wire N165808;
  wire N165806;
  wire N165888;
  wire N165886;
  wire N165753;
  wire N165751;
  wire N165913;
  wire N165911;
  wire N165778;
  wire N165776;
  wire N165398;
  wire N165396;
  wire N165873;
  wire N165871;
  wire N165838;
  wire N165836;
  wire N165678;
  wire N165676;
  wire N165883;
  wire N165881;
  wire N165858;
  wire N165856;
  wire N165853;
  wire N165851;
  wire N165813;
  wire N165811;
  wire N165903;
  wire N165901;
  wire N165718;
  wire N165716;
  wire N165908;
  wire N165906;
  wire N165763;
  wire N165761;
  wire N165938;
  wire N165936;
  wire N165833;
  wire N165831;
  wire N165553;
  wire N165551;
  wire \DLX_EXinst_N75154/F5MUX ;
  wire N165433;
  wire N165431;
  wire \DLX_IDinst_RegFile_22_14/F5MUX ;
  wire vga_top_vga1_vcounter_Madd__n0000_inst_lut2_9;
  wire \vga_top_vga1_vcounter<0>/CYMUXG ;
  wire \vga_top_vga1_vcounter<0>/GROM ;
  wire vga_top_vga1_vcounter_Madd__n0000_inst_cy_9;
  wire \vga_top_vga1_vcounter<0>/LOGIC_ZERO ;
  wire \vga_top_vga1_vcounter<2>/FROM ;
  wire \vga_top_vga1_vcounter<2>/CYMUXG ;
  wire \vga_top_vga1_vcounter<2>/LOGIC_ZERO ;
  wire \vga_top_vga1_vcounter<2>/GROM ;
  wire vga_top_vga1_vcounter_Madd__n0000_inst_cy_11;
  wire \vga_top_vga1_vcounter<2>/CYINIT ;
  wire \vga_top_vga1_vcounter<4>/FROM ;
  wire \vga_top_vga1_vcounter<4>/CYMUXG ;
  wire \vga_top_vga1_vcounter<4>/LOGIC_ZERO ;
  wire \vga_top_vga1_vcounter<4>/GROM ;
  wire vga_top_vga1_vcounter_Madd__n0000_inst_cy_13;
  wire \vga_top_vga1_vcounter<4>/CYINIT ;
  wire \vga_top_vga1_vcounter<6>/FROM ;
  wire \vga_top_vga1_vcounter<6>/CYMUXG ;
  wire \vga_top_vga1_vcounter<6>/LOGIC_ZERO ;
  wire \vga_top_vga1_vcounter<6>/GROM ;
  wire vga_top_vga1_vcounter_Madd__n0000_inst_cy_15;
  wire \vga_top_vga1_vcounter<6>/CYINIT ;
  wire \vga_top_vga1_vcounter<8>/LOGIC_ZERO ;
  wire \vga_top_vga1_vcounter<8>/FROM ;
  wire \vga_top_vga1_vcounter<9>_rt ;
  wire vga_top_vga1_vcounter_Madd__n0000_inst_cy_17;
  wire \vga_top_vga1_vcounter<8>/CYINIT ;
  wire DLX_EXinst_Mcompar__n0059_inst_lut4_0;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_103/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0059_inst_lut4_1;
  wire DLX_EXinst_Mcompar__n0059_inst_cy_102;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_103/LOGIC_ZERO ;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_103/LOGIC_ONE ;
  wire DLX_EXinst_Mcompar__n0059_inst_lut4_2;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_105/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0059_inst_lut4_3;
  wire DLX_EXinst_Mcompar__n0059_inst_cy_104;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_105/LOGIC_ZERO ;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_105/CYINIT ;
  wire DLX_EXinst_Mcompar__n0059_inst_lut4_4;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_107/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0059_inst_lut4_5;
  wire DLX_EXinst_Mcompar__n0059_inst_cy_106;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_107/LOGIC_ZERO ;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_107/CYINIT ;
  wire DLX_EXinst_Mcompar__n0059_inst_lut4_6;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_109/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0059_inst_lut4_7;
  wire DLX_EXinst_Mcompar__n0059_inst_cy_108;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_109/LOGIC_ZERO ;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_109/CYINIT ;
  wire DLX_EXinst_Mcompar__n0059_inst_lut4_8;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_111/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0059_inst_lut4_9;
  wire DLX_EXinst_Mcompar__n0059_inst_cy_110;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_111/LOGIC_ZERO ;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_111/CYINIT ;
  wire DLX_EXinst_Mcompar__n0059_inst_lut4_10;
  wire \DLX_IDinst_RegFile_14_12/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0059_inst_lut4_11;
  wire DLX_EXinst_Mcompar__n0059_inst_cy_112;
  wire \DLX_IDinst_RegFile_14_12/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_14_12/CYINIT ;
  wire DLX_EXinst_Mcompar__n0059_inst_lut4_12;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_115/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0059_inst_lut4_13;
  wire DLX_EXinst_Mcompar__n0059_inst_cy_114;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_115/LOGIC_ZERO ;
  wire \DLX_EXinst_Mcompar__n0059_inst_cy_115/CYINIT ;
  wire DLX_EXinst_Mcompar__n0059_inst_lut4_14;
  wire \DLX_IDinst_RegFile_30_17/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0059_inst_lut4_15;
  wire DLX_EXinst_Mcompar__n0059_inst_cy_116;
  wire \DLX_IDinst_RegFile_30_17/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_30_17/CYINIT ;
  wire DLX_EXinst_Mcompar__n0067_inst_lut2_134;
  wire \DLX_EXinst_Mcompar__n0067_inst_cy_199/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0067_inst_lut2_135;
  wire DLX_EXinst_Mcompar__n0067_inst_cy_198;
  wire \DLX_EXinst_Mcompar__n0067_inst_cy_199/LOGIC_ZERO ;
  wire DLX_EXinst_Mcompar__n0067_inst_lut2_136;
  wire \DLX_IDinst_RegFile_11_3/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0067_inst_lut2_137;
  wire DLX_EXinst_Mcompar__n0067_inst_cy_200;
  wire \DLX_IDinst_RegFile_11_3/CYINIT ;
  wire DLX_EXinst_Mcompar__n0067_inst_lut2_138;
  wire \DLX_EXinst_Mcompar__n0067_inst_cy_203/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0067_inst_lut2_139;
  wire DLX_EXinst_Mcompar__n0067_inst_cy_202;
  wire \DLX_EXinst_Mcompar__n0067_inst_cy_203/CYINIT ;
  wire DLX_EXinst_Mcompar__n0067_inst_lut2_140;
  wire \DLX_IDinst_RegFile_14_17/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0067_inst_lut2_141;
  wire DLX_EXinst_Mcompar__n0067_inst_cy_204;
  wire \DLX_IDinst_RegFile_14_17/CYINIT ;
  wire DLX_EXinst_Mcompar__n0067_inst_lut2_142;
  wire \DLX_EXinst_Mcompar__n0067_inst_cy_207/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0067_inst_lut2_143;
  wire DLX_EXinst_Mcompar__n0067_inst_cy_206;
  wire \DLX_EXinst_Mcompar__n0067_inst_cy_207/CYINIT ;
  wire DLX_EXinst_Mcompar__n0067_inst_lut2_144;
  wire \DLX_IDinst_RegFile_30_20/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0067_inst_lut2_145;
  wire DLX_EXinst_Mcompar__n0067_inst_cy_208;
  wire \DLX_IDinst_RegFile_30_20/CYINIT ;
  wire DLX_EXinst_Mcompar__n0067_inst_lut2_146;
  wire \DLX_EXinst_Mcompar__n0067_inst_cy_211/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0067_inst_lut2_147;
  wire DLX_EXinst_Mcompar__n0067_inst_cy_210;
  wire \DLX_EXinst_Mcompar__n0067_inst_cy_211/CYINIT ;
  wire DLX_EXinst_Mcompar__n0067_inst_lut2_148;
  wire \DLX_IDinst_RegFile_11_27/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0067_inst_lut2_149;
  wire DLX_EXinst_Mcompar__n0067_inst_cy_212;
  wire \DLX_IDinst_RegFile_11_27/CYINIT ;
  wire DLX_EXinst_Mcompar__n0067_inst_lut2_150;
  wire \DLX_EXinst_Mcompar__n0067_inst_cy_215/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0067_inst_lut2_151;
  wire DLX_EXinst_Mcompar__n0067_inst_cy_214;
  wire \DLX_EXinst_Mcompar__n0067_inst_cy_215/CYINIT ;
  wire DLX_EXinst_Mcompar__n0067_inst_lut2_152;
  wire \DLX_IDinst_RegFile_18_3/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0067_inst_lut2_153;
  wire DLX_EXinst_Mcompar__n0067_inst_cy_216;
  wire \DLX_IDinst_RegFile_18_3/CYINIT ;
  wire DLX_EXinst_Mcompar__n0067_inst_lut2_154;
  wire \DLX_EXinst_Mcompar__n0067_inst_cy_219/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0067_inst_lut2_155;
  wire DLX_EXinst_Mcompar__n0067_inst_cy_218;
  wire \DLX_EXinst_Mcompar__n0067_inst_cy_219/CYINIT ;
  wire DLX_EXinst_Mcompar__n0067_inst_lut2_156;
  wire \DLX_IDinst_RegFile_22_26/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0067_inst_lut2_157;
  wire DLX_EXinst_Mcompar__n0067_inst_cy_220;
  wire \DLX_IDinst_RegFile_22_26/CYINIT ;
  wire DLX_EXinst_Mcompar__n0067_inst_lut2_158;
  wire \DLX_EXinst_Mcompar__n0067_inst_cy_223/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0067_inst_lut2_159;
  wire DLX_EXinst_Mcompar__n0067_inst_cy_222;
  wire \DLX_EXinst_Mcompar__n0067_inst_cy_223/CYINIT ;
  wire DLX_EXinst_Mcompar__n0067_inst_lut2_160;
  wire \DLX_IDinst_RegFile_30_13/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0067_inst_lut2_161;
  wire DLX_EXinst_Mcompar__n0067_inst_cy_224;
  wire \DLX_IDinst_RegFile_30_13/CYINIT ;
  wire DLX_EXinst_Mcompar__n0067_inst_lut2_162;
  wire \DLX_EXinst_Mcompar__n0067_inst_cy_227/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0067_inst_lut2_163;
  wire DLX_EXinst_Mcompar__n0067_inst_cy_226;
  wire \DLX_EXinst_Mcompar__n0067_inst_cy_227/CYINIT ;
  wire DLX_EXinst_Mcompar__n0067_inst_lut2_164;
  wire \DLX_EXinst_Mcompar__n0067_inst_cy_228/CYMUXF ;
  wire \DLX_EXinst_Mcompar__n0067_inst_cy_228/CYINIT ;
  wire vga_top_vga1_gridvcounter_Madd__n0000_inst_lut2_0;
  wire \vga_top_vga1_gridvcounter<0>/CYMUXG ;
  wire \vga_top_vga1_gridvcounter<0>/GROM ;
  wire vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_0;
  wire \vga_top_vga1_gridvcounter<0>/LOGIC_ZERO ;
  wire \vga_top_vga1_gridvcounter<2>/FROM ;
  wire \vga_top_vga1_gridvcounter<2>/CYMUXG ;
  wire \vga_top_vga1_gridvcounter<2>/LOGIC_ZERO ;
  wire \vga_top_vga1_gridvcounter<2>/GROM ;
  wire vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_2;
  wire \vga_top_vga1_gridvcounter<2>/CYINIT ;
  wire \vga_top_vga1_gridvcounter<4>/FROM ;
  wire \vga_top_vga1_gridvcounter<4>/CYMUXG ;
  wire \vga_top_vga1_gridvcounter<4>/LOGIC_ZERO ;
  wire \vga_top_vga1_gridvcounter<4>/GROM ;
  wire vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_4;
  wire \vga_top_vga1_gridvcounter<4>/CYINIT ;
  wire \vga_top_vga1_gridvcounter<6>/FROM ;
  wire \vga_top_vga1_gridvcounter<6>/CYMUXG ;
  wire \vga_top_vga1_gridvcounter<6>/LOGIC_ZERO ;
  wire \vga_top_vga1_gridvcounter<6>/GROM ;
  wire vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_6;
  wire \vga_top_vga1_gridvcounter<6>/CYINIT ;
  wire \vga_top_vga1_gridvcounter<8>_rt ;
  wire \vga_top_vga1_gridvcounter<8>/CYINIT ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_102;
  wire \DLX_IDinst_RegFile_30_27/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_103;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_166;
  wire \DLX_IDinst_RegFile_30_27/LOGIC_ZERO ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_104;
  wire \DLX_EXinst_Mcompar__n0091_inst_cy_169/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_105;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_168;
  wire \DLX_EXinst_Mcompar__n0091_inst_cy_169/CYINIT ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_106;
  wire \DLX_IDinst_RegFile_22_30/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_107;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_170;
  wire \DLX_IDinst_RegFile_22_30/CYINIT ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_108;
  wire \DLX_EXinst_Mcompar__n0091_inst_cy_173/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_109;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_172;
  wire \DLX_EXinst_Mcompar__n0091_inst_cy_173/CYINIT ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_110;
  wire \DLX_IDinst_RegFile_1_6/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_111;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_174;
  wire \DLX_IDinst_RegFile_1_6/CYINIT ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_112;
  wire \DLX_EXinst_Mcompar__n0091_inst_cy_177/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_113;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_176;
  wire \DLX_EXinst_Mcompar__n0091_inst_cy_177/CYINIT ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_114;
  wire \DLX_IDinst_RegFile_30_22/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_115;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_178;
  wire \DLX_IDinst_RegFile_30_22/CYINIT ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_116;
  wire \DLX_EXinst_Mcompar__n0091_inst_cy_181/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_117;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_180;
  wire \DLX_EXinst_Mcompar__n0091_inst_cy_181/CYINIT ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_118;
  wire \DLX_IDinst_RegFile_30_18/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_119;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_182;
  wire \DLX_IDinst_RegFile_30_18/CYINIT ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_120;
  wire \DLX_EXinst_Mcompar__n0091_inst_cy_185/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_121;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_184;
  wire \DLX_EXinst_Mcompar__n0091_inst_cy_185/CYINIT ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_122;
  wire \DLX_IDinst_RegFile_22_23/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_123;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_186;
  wire \DLX_IDinst_RegFile_22_23/CYINIT ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_124;
  wire \DLX_EXinst_Mcompar__n0091_inst_cy_189/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_125;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_188;
  wire \DLX_EXinst_Mcompar__n0091_inst_cy_189/CYINIT ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_126;
  wire \DLX_IDinst_RegFile_15_11/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_127;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_190;
  wire \DLX_IDinst_RegFile_15_11/CYINIT ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_128;
  wire \DLX_EXinst_Mcompar__n0091_inst_cy_193/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_129;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_192;
  wire \DLX_EXinst_Mcompar__n0091_inst_cy_193/CYINIT ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_130;
  wire \DLX_IDinst_RegFile_3_6/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_131;
  wire DLX_EXinst_Mcompar__n0091_inst_cy_194;
  wire \DLX_IDinst_RegFile_3_6/CYINIT ;
  wire DLX_EXinst_Mcompar__n0091_inst_lut2_132;
  wire \DLX_EXinst_mem_to_reg_EX/CYMUXF ;
  wire \DLX_EXinst_mem_to_reg_EX/CYINIT ;
  wire DLX_IDinst_Msub__n0157_inst_lut2_198;
  wire \DLX_IDinst_RegFile_23_21/XORF ;
  wire \DLX_IDinst_RegFile_23_21/CYMUXG ;
  wire \DLX_IDinst_RegFile_23_21/XORG ;
  wire DLX_IDinst_Msub__n0157_inst_lut2_199;
  wire DLX_IDinst_Msub__n0157_inst_cy_265;
  wire \DLX_IDinst_RegFile_23_21/CYINIT ;
  wire \DLX_IDinst_RegFile_23_21/LOGIC_ONE ;
  wire \DLX_IDinst__n0157<2>/FROM ;
  wire \DLX_IDinst__n0157<2>/XORF ;
  wire \DLX_IDinst__n0157<2>/CYMUXG ;
  wire \DLX_IDinst__n0157<2>/XORG ;
  wire DLX_IDinst_Msub__n0157_inst_lut2_201;
  wire DLX_IDinst_Msub__n0157_inst_cy_267;
  wire \DLX_IDinst__n0157<2>/CYINIT ;
  wire DLX_IDinst_Msub__n0157_inst_lut2_202;
  wire \DLX_IDinst__n0157<4>/XORF ;
  wire \DLX_IDinst__n0157<4>/CYMUXG ;
  wire \DLX_IDinst__n0157<4>/XORG ;
  wire DLX_IDinst_Msub__n0157_inst_lut2_203;
  wire DLX_IDinst_Msub__n0157_inst_cy_269;
  wire \DLX_IDinst__n0157<4>/CYINIT ;
  wire DLX_IDinst_Msub__n0157_inst_lut2_204;
  wire \DLX_IDinst_RegFile_6_20/XORF ;
  wire \DLX_IDinst_RegFile_6_20/CYMUXG ;
  wire \DLX_IDinst_RegFile_6_20/XORG ;
  wire DLX_IDinst_Msub__n0157_inst_lut2_205;
  wire DLX_IDinst_Msub__n0157_inst_cy_271;
  wire \DLX_IDinst_RegFile_6_20/CYINIT ;
  wire DLX_IDinst_Msub__n0157_inst_lut2_206;
  wire \DLX_IDinst__n0157<8>/XORF ;
  wire \DLX_IDinst__n0157<8>/CYMUXG ;
  wire \DLX_IDinst__n0157<8>/XORG ;
  wire DLX_IDinst_Msub__n0157_inst_lut2_207;
  wire DLX_IDinst_Msub__n0157_inst_cy_273;
  wire \DLX_IDinst__n0157<8>/CYINIT ;
  wire DLX_IDinst_Msub__n0157_inst_lut2_208;
  wire \DLX_IDinst_RegFile_15_20/XORF ;
  wire \DLX_IDinst_RegFile_15_20/CYMUXG ;
  wire \DLX_IDinst_RegFile_15_20/XORG ;
  wire DLX_IDinst_Msub__n0157_inst_lut2_209;
  wire DLX_IDinst_Msub__n0157_inst_cy_275;
  wire \DLX_IDinst_RegFile_15_20/CYINIT ;
  wire DLX_IDinst_Msub__n0157_inst_lut2_210;
  wire \DLX_IDinst__n0157<12>/XORF ;
  wire \DLX_IDinst__n0157<12>/CYMUXG ;
  wire \DLX_IDinst__n0157<12>/XORG ;
  wire DLX_IDinst_Msub__n0157_inst_lut2_211;
  wire DLX_IDinst_Msub__n0157_inst_cy_277;
  wire \DLX_IDinst__n0157<12>/CYINIT ;
  wire DLX_IDinst_Msub__n0157_inst_lut2_212;
  wire \DLX_IDinst_RegFile_14_16/XORF ;
  wire \DLX_IDinst_RegFile_14_16/CYMUXG ;
  wire \DLX_IDinst_RegFile_14_16/XORG ;
  wire DLX_IDinst_Msub__n0157_inst_lut2_213;
  wire DLX_IDinst_Msub__n0157_inst_cy_279;
  wire \DLX_IDinst_RegFile_14_16/CYINIT ;
  wire DLX_IDinst_Msub__n0157_inst_lut2_214;
  wire \DLX_IDinst__n0157<16>/XORF ;
  wire \DLX_IDinst__n0157<16>/CYMUXG ;
  wire \DLX_IDinst__n0157<16>/XORG ;
  wire DLX_IDinst_Msub__n0157_inst_lut2_215;
  wire DLX_IDinst_Msub__n0157_inst_cy_281;
  wire \DLX_IDinst__n0157<16>/CYINIT ;
  wire DLX_IDinst_Msub__n0157_inst_lut2_216;
  wire \DLX_IDinst_RegFile_23_12/XORF ;
  wire \DLX_IDinst_RegFile_23_12/CYMUXG ;
  wire \DLX_IDinst_RegFile_23_12/XORG ;
  wire DLX_IDinst_Msub__n0157_inst_lut2_217;
  wire DLX_IDinst_Msub__n0157_inst_cy_283;
  wire \DLX_IDinst_RegFile_23_12/CYINIT ;
  wire DLX_IDinst_Msub__n0157_inst_lut2_218;
  wire \DLX_IDinst__n0157<20>/XORF ;
  wire \DLX_IDinst__n0157<20>/CYMUXG ;
  wire \DLX_IDinst__n0157<20>/XORG ;
  wire DLX_IDinst_Msub__n0157_inst_lut2_219;
  wire DLX_IDinst_Msub__n0157_inst_cy_285;
  wire \DLX_IDinst__n0157<20>/CYINIT ;
  wire DLX_IDinst_Msub__n0157_inst_lut2_220;
  wire \DLX_IDinst_RegFile_6_12/XORF ;
  wire \DLX_IDinst_RegFile_6_12/CYMUXG ;
  wire \DLX_IDinst_RegFile_6_12/XORG ;
  wire DLX_IDinst_Msub__n0157_inst_lut2_221;
  wire DLX_IDinst_Msub__n0157_inst_cy_287;
  wire \DLX_IDinst_RegFile_6_12/CYINIT ;
  wire DLX_IDinst_Msub__n0157_inst_lut2_222;
  wire \DLX_IDinst__n0157<24>/XORF ;
  wire \DLX_IDinst__n0157<24>/CYMUXG ;
  wire \DLX_IDinst__n0157<24>/XORG ;
  wire DLX_IDinst_Msub__n0157_inst_lut2_223;
  wire DLX_IDinst_Msub__n0157_inst_cy_289;
  wire \DLX_IDinst__n0157<24>/CYINIT ;
  wire DLX_IDinst_Msub__n0157_inst_lut2_224;
  wire \DLX_IDinst_RegFile_1_7/XORF ;
  wire \DLX_IDinst_RegFile_1_7/CYMUXG ;
  wire \DLX_IDinst_RegFile_1_7/XORG ;
  wire DLX_IDinst_Msub__n0157_inst_lut2_225;
  wire DLX_IDinst_Msub__n0157_inst_cy_291;
  wire \DLX_IDinst_RegFile_1_7/CYINIT ;
  wire DLX_IDinst_Msub__n0157_inst_lut2_226;
  wire \DLX_IDinst__n0157<28>/XORF ;
  wire \DLX_IDinst__n0157<28>/CYMUXG ;
  wire \DLX_IDinst__n0157<28>/XORG ;
  wire DLX_IDinst_Msub__n0157_inst_lut2_227;
  wire DLX_IDinst_Msub__n0157_inst_cy_293;
  wire \DLX_IDinst__n0157<28>/CYINIT ;
  wire DLX_IDinst_Msub__n0157_inst_lut2_228;
  wire \DLX_IDinst_RegFile_10_9/XORF ;
  wire \DLX_IDinst_RegFile_10_9/XORG ;
  wire DLX_IDinst_Msub__n0157_inst_lut2_229;
  wire DLX_IDinst_Msub__n0157_inst_cy_295;
  wire \DLX_IDinst_RegFile_10_9/CYINIT ;
  wire vga_top_vga1_gridhcounter_Madd__n0000_inst_lut2_0;
  wire \vga_top_vga1_gridhcounter<0>/CYMUXG ;
  wire \vga_top_vga1_gridhcounter<0>/GROM ;
  wire vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_0;
  wire \vga_top_vga1_gridhcounter<0>/LOGIC_ZERO ;
  wire \vga_top_vga1_gridhcounter<2>/FROM ;
  wire \vga_top_vga1_gridhcounter<2>/CYMUXG ;
  wire \vga_top_vga1_gridhcounter<2>/LOGIC_ZERO ;
  wire \vga_top_vga1_gridhcounter<2>/GROM ;
  wire vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_2;
  wire \vga_top_vga1_gridhcounter<2>/CYINIT ;
  wire \vga_top_vga1_gridhcounter<4>/FROM ;
  wire \vga_top_vga1_gridhcounter<4>/CYMUXG ;
  wire \vga_top_vga1_gridhcounter<4>/LOGIC_ZERO ;
  wire \vga_top_vga1_gridhcounter<4>/GROM ;
  wire vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_4;
  wire \vga_top_vga1_gridhcounter<4>/CYINIT ;
  wire \vga_top_vga1_gridhcounter<6>/FROM ;
  wire \vga_top_vga1_gridhcounter<6>/CYMUXG ;
  wire \vga_top_vga1_gridhcounter<6>/LOGIC_ZERO ;
  wire \vga_top_vga1_gridhcounter<6>/GROM ;
  wire vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_6;
  wire \vga_top_vga1_gridhcounter<6>/CYINIT ;
  wire \vga_top_vga1_gridhcounter<8>_rt ;
  wire \vga_top_vga1_gridhcounter<8>/CYINIT ;
  wire vga_top_vga1_hcounter_Madd__n0000_inst_lut2_19;
  wire \vga_top_vga1_hcounter<0>/CYMUXG ;
  wire \vga_top_vga1_hcounter<0>/GROM ;
  wire vga_top_vga1_hcounter_Madd__n0000_inst_cy_19;
  wire \vga_top_vga1_hcounter<0>/LOGIC_ZERO ;
  wire \vga_top_vga1_hcounter<2>/FROM ;
  wire \vga_top_vga1_hcounter<2>/CYMUXG ;
  wire \vga_top_vga1_hcounter<2>/LOGIC_ZERO ;
  wire \vga_top_vga1_hcounter<2>/GROM ;
  wire vga_top_vga1_hcounter_Madd__n0000_inst_cy_21;
  wire \vga_top_vga1_hcounter<2>/CYINIT ;
  wire \vga_top_vga1_hcounter<4>/FROM ;
  wire \vga_top_vga1_hcounter<4>/CYMUXG ;
  wire \vga_top_vga1_hcounter<4>/LOGIC_ZERO ;
  wire \vga_top_vga1_hcounter<4>/GROM ;
  wire vga_top_vga1_hcounter_Madd__n0000_inst_cy_23;
  wire \vga_top_vga1_hcounter<4>/CYINIT ;
  wire \vga_top_vga1_hcounter<6>/FROM ;
  wire \vga_top_vga1_hcounter<6>/CYMUXG ;
  wire \vga_top_vga1_hcounter<6>/LOGIC_ZERO ;
  wire \vga_top_vga1_hcounter<6>/GROM ;
  wire vga_top_vga1_hcounter_Madd__n0000_inst_cy_25;
  wire \vga_top_vga1_hcounter<6>/CYINIT ;
  wire \vga_top_vga1_hcounter<8>/FROM ;
  wire \vga_top_vga1_hcounter<8>/CYMUXG ;
  wire \vga_top_vga1_hcounter<8>/LOGIC_ZERO ;
  wire \vga_top_vga1_hcounter<8>/GROM ;
  wire vga_top_vga1_hcounter_Madd__n0000_inst_cy_27;
  wire \vga_top_vga1_hcounter<8>/CYINIT ;
  wire \vga_top_vga1_hcounter<10>/FROM ;
  wire \vga_top_vga1_hcounter<10>/CYMUXG ;
  wire \vga_top_vga1_hcounter<10>/LOGIC_ZERO ;
  wire \vga_top_vga1_hcounter<10>/GROM ;
  wire vga_top_vga1_hcounter_Madd__n0000_inst_cy_29;
  wire \vga_top_vga1_hcounter<10>/CYINIT ;
  wire \vga_top_vga1_hcounter<12>/FROM ;
  wire \vga_top_vga1_hcounter<12>/CYMUXG ;
  wire \vga_top_vga1_hcounter<12>/LOGIC_ZERO ;
  wire \vga_top_vga1_hcounter<12>/GROM ;
  wire vga_top_vga1_hcounter_Madd__n0000_inst_cy_31;
  wire \vga_top_vga1_hcounter<12>/CYINIT ;
  wire \vga_top_vga1_hcounter<14>/LOGIC_ZERO ;
  wire \vga_top_vga1_hcounter<14>/FROM ;
  wire \vga_top_vga1_hcounter<15>_rt ;
  wire vga_top_vga1_hcounter_Madd__n0000_inst_cy_33;
  wire \vga_top_vga1_hcounter<14>/CYINIT ;
  wire vga_top_vga1_Mmult__n0043_inst_lut2_303;
  wire \vga_top_vga1_Mmult__n0043_inst_lut2_317/CYMUXG ;
  wire \vga_top_vga1_Mmult__n0043_inst_lut2_317/XORG ;
  wire vga_top_vga1_Mmult__n0043_inst_lut2_304;
  wire vga_top_vga1_Mmult__n0043_inst_cy_436;
  wire \vga_top_vga1_Mmult__n0043_inst_lut2_317/LOGIC_ZERO ;
  wire vga_top_vga1_Mmult__n0043_inst_lut2_305;
  wire \DLX_IDinst_RegFile_3_14/XORF ;
  wire \DLX_IDinst_RegFile_3_14/CYMUXG ;
  wire \DLX_IDinst_RegFile_3_14/XORG ;
  wire vga_top_vga1_Mmult__n0043_inst_lut2_306;
  wire vga_top_vga1_Mmult__n0043_inst_cy_438;
  wire \DLX_IDinst_RegFile_3_14/CYINIT ;
  wire vga_top_vga1_Mmult__n0043_inst_lut2_307;
  wire \vga_top_vga1_Mmult__n0043_inst_lut2_320/XORF ;
  wire \vga_top_vga1_Mmult__n0043_inst_lut2_320/CYMUXG ;
  wire \vga_top_vga1_Mmult__n0043_inst_lut2_320/XORG ;
  wire vga_top_vga1_Mmult__n0043_inst_lut2_308;
  wire vga_top_vga1_Mmult__n0043_inst_cy_440;
  wire \vga_top_vga1_Mmult__n0043_inst_lut2_320/CYINIT ;
  wire vga_top_vga1_Mmult__n0043_inst_lut2_309;
  wire \vga_top_vga1_Mmult__n0043_inst_lut2_322/XORF ;
  wire \vga_top_vga1_Mmult__n0043_inst_lut2_322/XORG ;
  wire \$SIG_0 ;
  wire vga_top_vga1_Mmult__n0043_inst_cy_442;
  wire \vga_top_vga1_Mmult__n0043_inst_lut2_322/CYINIT ;
  wire \$SIG_1 ;
  wire \vga_top_vga1_Mcompar__n0034_inst_cy_329/CYMUXG ;
  wire \$SIG_2 ;
  wire vga_top_vga1_Mcompar__n0034_inst_cy_328;
  wire \vga_top_vga1_Mcompar__n0034_inst_cy_329/LOGIC_ZERO ;
  wire \vga_top_vga1_Mcompar__n0034_inst_cy_329/LOGIC_ONE ;
  wire vga_top_vga1_Mcompar__n0034_inst_lut2_262;
  wire \DLX_IDinst_RegFile_6_13/CYMUXG ;
  wire vga_top_vga1_Mcompar__n0034_inst_lut2_263;
  wire vga_top_vga1_Mcompar__n0034_inst_cy_330;
  wire \DLX_IDinst_RegFile_6_13/LOGIC_ONE ;
  wire \DLX_IDinst_RegFile_6_13/CYINIT ;
  wire \$SIG_3 ;
  wire \vga_top_vga1_Mcompar__n0034_inst_cy_333/CYMUXG ;
  wire \$SIG_4 ;
  wire vga_top_vga1_Mcompar__n0034_inst_cy_332;
  wire \vga_top_vga1_Mcompar__n0034_inst_cy_333/LOGIC_ZERO ;
  wire \vga_top_vga1_Mcompar__n0034_inst_cy_333/CYINIT ;
  wire vga_top_vga1_Mcompar__n0034_inst_lut2_264;
  wire \vga_top_vga1_Mcompar__n0034_inst_cy_335/CYMUXG ;
  wire vga_top_vga1_Mcompar__n0034_inst_lut2_265;
  wire vga_top_vga1_Mcompar__n0034_inst_cy_334;
  wire \vga_top_vga1_Mcompar__n0034_inst_cy_335/LOGIC_ONE ;
  wire \vga_top_vga1_Mcompar__n0034_inst_cy_335/CYINIT ;
  wire vga_top_vga1_Mcompar__n0034_inst_lut2_266;
  wire \DLX_IDinst_RegFile_14_29/CYMUXG ;
  wire vga_top_vga1_Mcompar__n0034_inst_lut2_267;
  wire vga_top_vga1_Mcompar__n0034_inst_cy_336;
  wire \DLX_IDinst_RegFile_14_29/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_14_29/CYINIT ;
  wire vga_top_vga1_Mcompar__n0034_inst_lut4_1099;
  wire \vga_top_vga1__n0034/CYMUXG ;
  wire vga_top_vga1_Mcompar__n0034_inst_lut2_268;
  wire vga_top_vga1_Mcompar__n0034_inst_cy_338;
  wire \vga_top_vga1__n0034/LOGIC_ONE ;
  wire \vga_top_vga1__n0034/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_155;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_97/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_156;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_96;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_97/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_97/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_251;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_193/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_252;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_192;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_193/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_193/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_171;
  wire \DLX_EXinst_reg_write_EX/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_172;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_112;
  wire \DLX_EXinst_reg_write_EX/LOGIC_ZERO ;
  wire \DLX_EXinst_reg_write_EX/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_179;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_121/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_180;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_120;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_121/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_121/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_267;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_209/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_268;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_208;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_209/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_209/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_187;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_129/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_188;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_128;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_129/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_129/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_347;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_289/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_348;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_288;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_289/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_289/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_353;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_295/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_354;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_294;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_295/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_295/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_363;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_305/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_364;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_304;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_305/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_305/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_283;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_225/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_284;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_224;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_225/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_225/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_203;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_145/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_204;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_144;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_145/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_145/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_459;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_401/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_460;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_400;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_401/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_401/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_379;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_321/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_380;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_320;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_321/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_321/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_299;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_241/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_300;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_240;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_241/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_241/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_219;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_161/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_220;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_160;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_161/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_161/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_555;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_497/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_556;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_496;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_497/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_497/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_475;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_417/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_476;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_416;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_417/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_417/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_395;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_337/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_396;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_336;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_337/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_337/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_315;
  wire \DLX_EXinst_reg_out_B_EX<3>/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_316;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_256;
  wire \DLX_EXinst_reg_out_B_EX<3>/LOGIC_ZERO ;
  wire \DLX_EXinst_reg_out_B_EX<3>/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_235;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_177/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_236;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_176;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_177/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_177/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_491;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_433/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_492;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_432;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_433/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_433/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_411;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_353/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_412;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_352;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_353/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_353/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_331;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_273/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_332;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_272;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_273/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_273/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_507;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_449/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_508;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_448;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_449/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_449/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_427;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_369/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_428;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_368;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_369/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_369/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_439;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_381/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_440;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_380;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_381/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_381/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_523;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_465/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_524;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_464;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_465/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_465/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_525;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_467/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_526;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_466;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_467/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_467/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_443;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_385/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_444;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_384;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_385/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_385/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_539;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_481/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_540;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_480;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_481/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_481/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_59;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_1/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_60;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_0;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_1/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_1/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_75;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_17/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_76;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_16;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_17/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_17/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_91;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_33/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_92;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_32;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_33/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_33/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_99;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_41/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_100;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_40;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_41/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_41/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_107;
  wire \DLX_IDinst_Cause_Reg<6>/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_108;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_48;
  wire \DLX_IDinst_Cause_Reg<6>/LOGIC_ZERO ;
  wire \DLX_IDinst_Cause_Reg<6>/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_123;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_65/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_124;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_64;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_65/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_65/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_139;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_81/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_140;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_80;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_81/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_4_inst_cy_81/LOGIC_ONE ;
  wire DLX_EXinst_Mcompar__n0065_inst_lut2_102;
  wire \DLX_EXinst_Mcompar__n0065_inst_cy_167/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0065_inst_lut2_103;
  wire DLX_EXinst_Mcompar__n0065_inst_cy_166;
  wire \DLX_EXinst_Mcompar__n0065_inst_cy_167/LOGIC_ZERO ;
  wire DLX_EXinst_Mcompar__n0065_inst_lut2_104;
  wire \DLX_IDinst_RegFile_3_0/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0065_inst_lut2_105;
  wire DLX_EXinst_Mcompar__n0065_inst_cy_168;
  wire \DLX_IDinst_RegFile_3_0/CYINIT ;
  wire DLX_EXinst_Mcompar__n0065_inst_lut2_106;
  wire \DLX_EXinst_Mcompar__n0065_inst_cy_171/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0065_inst_lut2_107;
  wire DLX_EXinst_Mcompar__n0065_inst_cy_170;
  wire \DLX_EXinst_Mcompar__n0065_inst_cy_171/CYINIT ;
  wire DLX_EXinst_Mcompar__n0065_inst_lut2_108;
  wire \DLX_IDinst_RegFile_31_11/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0065_inst_lut2_109;
  wire DLX_EXinst_Mcompar__n0065_inst_cy_172;
  wire \DLX_IDinst_RegFile_31_11/CYINIT ;
  wire DLX_EXinst_Mcompar__n0065_inst_lut2_110;
  wire \DLX_EXinst_Mcompar__n0065_inst_cy_175/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0065_inst_lut2_111;
  wire DLX_EXinst_Mcompar__n0065_inst_cy_174;
  wire \DLX_EXinst_Mcompar__n0065_inst_cy_175/CYINIT ;
  wire DLX_EXinst_Mcompar__n0065_inst_lut2_112;
  wire \DLX_IDinst_RegFile_3_30/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0065_inst_lut2_113;
  wire DLX_EXinst_Mcompar__n0065_inst_cy_176;
  wire \DLX_IDinst_RegFile_3_30/CYINIT ;
  wire DLX_EXinst_Mcompar__n0065_inst_lut2_114;
  wire \DLX_EXinst_Mcompar__n0065_inst_cy_179/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0065_inst_lut2_115;
  wire DLX_EXinst_Mcompar__n0065_inst_cy_178;
  wire \DLX_EXinst_Mcompar__n0065_inst_cy_179/CYINIT ;
  wire DLX_EXinst_Mcompar__n0065_inst_lut2_116;
  wire \DLX_IDinst_RegFile_22_28/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0065_inst_lut2_117;
  wire DLX_EXinst_Mcompar__n0065_inst_cy_180;
  wire \DLX_IDinst_RegFile_22_28/CYINIT ;
  wire DLX_EXinst_Mcompar__n0065_inst_lut2_118;
  wire \DLX_EXinst_Mcompar__n0065_inst_cy_183/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0065_inst_lut2_119;
  wire DLX_EXinst_Mcompar__n0065_inst_cy_182;
  wire \DLX_EXinst_Mcompar__n0065_inst_cy_183/CYINIT ;
  wire DLX_EXinst_Mcompar__n0065_inst_lut2_120;
  wire \DLX_IDinst_RegFile_1_8/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0065_inst_lut2_121;
  wire DLX_EXinst_Mcompar__n0065_inst_cy_184;
  wire \DLX_IDinst_RegFile_1_8/CYINIT ;
  wire DLX_EXinst_Mcompar__n0065_inst_lut2_122;
  wire \DLX_EXinst_Mcompar__n0065_inst_cy_187/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0065_inst_lut2_123;
  wire DLX_EXinst_Mcompar__n0065_inst_cy_186;
  wire \DLX_EXinst_Mcompar__n0065_inst_cy_187/CYINIT ;
  wire DLX_EXinst_Mcompar__n0065_inst_lut2_124;
  wire \DLX_IDinst_RegFile_31_20/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0065_inst_lut2_125;
  wire DLX_EXinst_Mcompar__n0065_inst_cy_188;
  wire \DLX_IDinst_RegFile_31_20/CYINIT ;
  wire DLX_EXinst_Mcompar__n0065_inst_lut2_126;
  wire \DLX_EXinst_Mcompar__n0065_inst_cy_191/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0065_inst_lut2_127;
  wire DLX_EXinst_Mcompar__n0065_inst_cy_190;
  wire \DLX_EXinst_Mcompar__n0065_inst_cy_191/CYINIT ;
  wire DLX_EXinst_Mcompar__n0065_inst_lut2_128;
  wire \DLX_IDinst_RegFile_24_12/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0065_inst_lut2_129;
  wire DLX_EXinst_Mcompar__n0065_inst_cy_192;
  wire \DLX_IDinst_RegFile_24_12/CYINIT ;
  wire DLX_EXinst_Mcompar__n0065_inst_lut2_130;
  wire \DLX_EXinst_Mcompar__n0065_inst_cy_195/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0065_inst_lut2_131;
  wire DLX_EXinst_Mcompar__n0065_inst_cy_194;
  wire \DLX_EXinst_Mcompar__n0065_inst_cy_195/CYINIT ;
  wire DLX_EXinst_Mcompar__n0065_inst_lut2_132;
  wire \DLX_EXinst_Mcompar__n0065_inst_cy_196/CYMUXF ;
  wire \DLX_EXinst_Mcompar__n0065_inst_cy_196/CYINIT ;
  wire vga_top_vga1_Mcompar__n0029_inst_lut1_22;
  wire \DLX_IDinst_RegFile_15_13/CYMUXG ;
  wire vga_top_vga1_Mcompar__n0029_inst_lut1_23;
  wire vga_top_vga1_Mcompar__n0029_inst_cy_370;
  wire \DLX_IDinst_RegFile_15_13/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_15_13/LOGIC_ONE ;
  wire \$SIG_5 ;
  wire \vga_top_vga1_Mcompar__n0029_inst_cy_373/CYMUXG ;
  wire \$SIG_6 ;
  wire vga_top_vga1_Mcompar__n0029_inst_cy_372;
  wire \vga_top_vga1_Mcompar__n0029_inst_cy_373/LOGIC_ONE ;
  wire \vga_top_vga1_Mcompar__n0029_inst_cy_373/CYINIT ;
  wire vga_top_vga1_Mcompar__n0029_inst_lut4_1104;
  wire \vga_top_vga1_Mcompar__n0029_inst_cy_375/CYMUXG ;
  wire vga_top_vga1_Mcompar__n0029_inst_lut4_1105;
  wire vga_top_vga1_Mcompar__n0029_inst_cy_374;
  wire \vga_top_vga1_Mcompar__n0029_inst_cy_375/LOGIC_ZERO ;
  wire \vga_top_vga1_Mcompar__n0029_inst_cy_375/CYINIT ;
  wire vga_top_vga1_Mcompar__n0029_inst_lut4_1106;
  wire \DLX_IFinst_IR_curr<10>/CYMUXG ;
  wire vga_top_vga1_Mcompar__n0029_inst_lut2_275;
  wire vga_top_vga1_Mcompar__n0029_inst_cy_376;
  wire \DLX_IFinst_IR_curr<10>/LOGIC_ZERO ;
  wire \DLX_IFinst_IR_curr<10>/CYINIT ;
  wire vga_top_vga1_Mcompar__n0037_inst_lut2_341;
  wire \vga_top_vga1_Mcompar__n0037_inst_cy_472/CYMUXG ;
  wire vga_top_vga1_Mcompar__n0037_inst_lut2_342;
  wire vga_top_vga1_Mcompar__n0037_inst_cy_471;
  wire \vga_top_vga1_Mcompar__n0037_inst_cy_472/LOGIC_ZERO ;
  wire \vga_top_vga1_Mcompar__n0037_inst_cy_472/LOGIC_ONE ;
  wire vga_top_vga1_Mcompar__n0037_inst_lut4_1139;
  wire \DLX_IDinst_RegFile_30_29/CYMUXG ;
  wire vga_top_vga1_Mcompar__n0037_inst_lut4_1140;
  wire vga_top_vga1_Mcompar__n0037_inst_cy_473;
  wire \DLX_IDinst_RegFile_30_29/LOGIC_ONE ;
  wire \DLX_IDinst_RegFile_30_29/CYINIT ;
  wire vga_top_vga1_Mcompar__n0037_inst_lut4_1141;
  wire \vga_top_vga1__n0037/CYMUXG ;
  wire vga_top_vga1_Mcompar__n0037_inst_lut2_343;
  wire vga_top_vga1_Mcompar__n0037_inst_cy_475;
  wire \vga_top_vga1__n0037/LOGIC_ONE ;
  wire \vga_top_vga1__n0037/CYINIT ;
  wire DLX_IDinst_Mcompar__n0368_inst_lut4_40;
  wire \DLX_IDinst_Mcompar__n0368_inst_cy_263/CYMUXG ;
  wire DLX_IDinst_Mcompar__n0368_inst_lut4_41;
  wire DLX_IDinst_Mcompar__n0368_inst_cy_262;
  wire \DLX_IDinst_Mcompar__n0368_inst_cy_263/LOGIC_ZERO ;
  wire \DLX_IDinst_Mcompar__n0368_inst_cy_263/LOGIC_ONE ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_70;
  wire \DLX_EXinst_Mcompar__n0063_inst_cy_135/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_71;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_134;
  wire \DLX_EXinst_Mcompar__n0063_inst_cy_135/LOGIC_ZERO ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_72;
  wire \DLX_IDinst_RegFile_15_22/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_73;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_136;
  wire \DLX_IDinst_RegFile_15_22/CYINIT ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_74;
  wire \DLX_EXinst_Mcompar__n0063_inst_cy_139/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_75;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_138;
  wire \DLX_EXinst_Mcompar__n0063_inst_cy_139/CYINIT ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_76;
  wire \DLX_IFinst_IR_curr<11>/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_77;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_140;
  wire \DLX_IFinst_IR_curr<11>/CYINIT ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_78;
  wire \DLX_EXinst_Mcompar__n0063_inst_cy_143/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_79;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_142;
  wire \DLX_EXinst_Mcompar__n0063_inst_cy_143/CYINIT ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_80;
  wire \DLX_IDinst_RegFile_23_14/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_81;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_144;
  wire \DLX_IDinst_RegFile_23_14/CYINIT ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_82;
  wire \DLX_EXinst_Mcompar__n0063_inst_cy_147/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_83;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_146;
  wire \DLX_EXinst_Mcompar__n0063_inst_cy_147/CYINIT ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_84;
  wire \DLX_IDinst_RegFile_26_3/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_85;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_148;
  wire \DLX_IDinst_RegFile_26_3/CYINIT ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_86;
  wire \DLX_EXinst_Mcompar__n0063_inst_cy_151/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_87;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_150;
  wire \DLX_EXinst_Mcompar__n0063_inst_cy_151/CYINIT ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_88;
  wire \DLX_IDinst_RegFile_15_23/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_89;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_152;
  wire \DLX_IDinst_RegFile_15_23/CYINIT ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_90;
  wire \DLX_EXinst_Mcompar__n0063_inst_cy_155/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_91;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_154;
  wire \DLX_EXinst_Mcompar__n0063_inst_cy_155/CYINIT ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_92;
  wire \DLX_IFinst_IR_curr<20>/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_93;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_156;
  wire \DLX_IFinst_IR_curr<20>/CYINIT ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_94;
  wire \DLX_EXinst_Mcompar__n0063_inst_cy_159/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_95;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_158;
  wire \DLX_EXinst_Mcompar__n0063_inst_cy_159/CYINIT ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_96;
  wire \DLX_IDinst_RegFile_31_23/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_97;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_160;
  wire \DLX_IDinst_RegFile_31_23/CYINIT ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_98;
  wire \DLX_EXinst_Mcompar__n0063_inst_cy_163/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0063_inst_lut2_99;
  wire DLX_EXinst_Mcompar__n0063_inst_cy_162;
  wire \DLX_EXinst_Mcompar__n0063_inst_cy_163/CYINIT ;
  wire vga_top_vga1_Mcompar__n0030_inst_lut4_1101;
  wire \DLX_IDinst_RegFile_31_29/CYMUXG ;
  wire vga_top_vga1_Mcompar__n0030_inst_lut4_1102;
  wire vga_top_vga1_Mcompar__n0030_inst_cy_354;
  wire \DLX_IDinst_RegFile_31_29/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_31_29/LOGIC_ONE ;
  wire vga_top_vga1_Mcompar__n0030_inst_lut1_10;
  wire \vga_top_vga1_Mcompar__n0030_inst_cy_357/CYMUXG ;
  wire vga_top_vga1_Mcompar__n0030_inst_lut1_11;
  wire vga_top_vga1_Mcompar__n0030_inst_cy_356;
  wire \vga_top_vga1_Mcompar__n0030_inst_cy_357/LOGIC_ONE ;
  wire \vga_top_vga1_Mcompar__n0030_inst_cy_357/CYINIT ;
  wire \$SIG_7 ;
  wire \vga_top_vga1_Mcompar__n0030_inst_cy_359/CYMUXG ;
  wire \$SIG_8 ;
  wire vga_top_vga1_Mcompar__n0030_inst_cy_358;
  wire \vga_top_vga1_Mcompar__n0030_inst_cy_359/LOGIC_ZERO ;
  wire \vga_top_vga1_Mcompar__n0030_inst_cy_359/CYINIT ;
  wire vga_top_vga1_Mcompar__n0030_inst_lut1_14;
  wire \DLX_IDinst_RegFile_31_31/CYMUXG ;
  wire vga_top_vga1_Mcompar__n0030_inst_lut1_15;
  wire vga_top_vga1_Mcompar__n0030_inst_cy_360;
  wire \DLX_IDinst_RegFile_31_31/LOGIC_ONE ;
  wire \DLX_IDinst_RegFile_31_31/CYINIT ;
  wire \$SIG_9 ;
  wire \vga_top_vga1_Mcompar__n0030_inst_cy_363/CYMUXG ;
  wire \$SIG_10 ;
  wire vga_top_vga1_Mcompar__n0030_inst_cy_362;
  wire \vga_top_vga1_Mcompar__n0030_inst_cy_363/LOGIC_ZERO ;
  wire \vga_top_vga1_Mcompar__n0030_inst_cy_363/CYINIT ;
  wire vga_top_vga1_Mcompar__n0030_inst_lut1_18;
  wire \vga_top_vga1_Mcompar__n0030_inst_cy_365/CYMUXG ;
  wire vga_top_vga1_Mcompar__n0030_inst_lut1_19;
  wire vga_top_vga1_Mcompar__n0030_inst_cy_364;
  wire \vga_top_vga1_Mcompar__n0030_inst_cy_365/LOGIC_ONE ;
  wire \vga_top_vga1_Mcompar__n0030_inst_cy_365/CYINIT ;
  wire \$SIG_11 ;
  wire \vga_top_vga1_Mcompar__n0030_inst_cy_367/CYMUXG ;
  wire \$SIG_12 ;
  wire vga_top_vga1_Mcompar__n0030_inst_cy_366;
  wire \vga_top_vga1_Mcompar__n0030_inst_cy_367/LOGIC_ZERO ;
  wire \vga_top_vga1_Mcompar__n0030_inst_cy_367/CYINIT ;
  wire vga_top_vga1_Mcompar__n0030_inst_lut4_1103;
  wire \DLX_IFinst_IR_curr<12>/CYMUXG ;
  wire vga_top_vga1_Mcompar__n0030_inst_lut2_274;
  wire vga_top_vga1_Mcompar__n0030_inst_cy_368;
  wire \DLX_IFinst_IR_curr<12>/LOGIC_ONE ;
  wire \DLX_IFinst_IR_curr<12>/CYINIT ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_70;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_135/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_71;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_134;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_135/LOGIC_ZERO ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_72;
  wire \DLX_IDinst_RegFile_23_16/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_73;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_136;
  wire \DLX_IDinst_RegFile_23_16/CYINIT ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_74;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_139/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_75;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_138;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_139/CYINIT ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_76;
  wire \vga_top_vga1_clockcounter_FFd2/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_77;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_140;
  wire \vga_top_vga1_clockcounter_FFd2/CYINIT ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_78;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_143/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_79;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_142;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_143/CYINIT ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_80;
  wire \DLX_IDinst_RegFile_6_26/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_81;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_144;
  wire \DLX_IDinst_RegFile_6_26/CYINIT ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_82;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_147/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_83;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_146;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_147/CYINIT ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_84;
  wire \DLX_IFinst_IR_curr<21>/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_85;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_148;
  wire \DLX_IFinst_IR_curr<21>/CYINIT ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_86;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_151/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_87;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_150;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_151/CYINIT ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_88;
  wire \DLX_IDinst_RegFile_7_11/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_89;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_152;
  wire \DLX_IDinst_RegFile_7_11/CYINIT ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_90;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_155/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_91;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_154;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_155/CYINIT ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_92;
  wire \DLX_IDinst_RegFile_3_23/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_93;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_156;
  wire \DLX_IDinst_RegFile_3_23/CYINIT ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_94;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_159/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_95;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_158;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_159/CYINIT ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_96;
  wire \DLX_IDinst_RegFile_31_17/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_97;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_160;
  wire \DLX_IDinst_RegFile_31_17/CYINIT ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_98;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_163/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_99;
  wire DLX_EXinst_Mcompar__n0089_inst_cy_162;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_163/CYINIT ;
  wire DLX_EXinst_Mcompar__n0089_inst_lut2_100;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_164/CYMUXF ;
  wire \DLX_EXinst_Mcompar__n0089_inst_cy_164/CYINIT ;
  wire DLX_IDinst_Mcompar__n0104_inst_lut4_40;
  wire \DLX_IDinst_Mcompar__n0104_inst_cy_263/CYMUXG ;
  wire DLX_IDinst_Mcompar__n0104_inst_lut4_41;
  wire DLX_IDinst_Mcompar__n0104_inst_cy_262;
  wire \DLX_IDinst_Mcompar__n0104_inst_cy_263/LOGIC_ZERO ;
  wire \DLX_IDinst_Mcompar__n0104_inst_cy_263/LOGIC_ONE ;
  wire \DLX_IDinst__n0104/LOGIC_ZERO ;
  wire DLX_IDinst_Mcompar__n0104_inst_lut4_42;
  wire \DLX_IDinst__n0104/CYMUXF ;
  wire \DLX_IDinst__n0104/CYINIT ;
  wire DLX_EXinst_Mcompar__n0061_inst_lut4_16;
  wire \DLX_EXinst_Mcompar__n0061_inst_cy_119/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0061_inst_lut4_17;
  wire DLX_EXinst_Mcompar__n0061_inst_cy_118;
  wire \DLX_EXinst_Mcompar__n0061_inst_cy_119/LOGIC_ONE ;
  wire \DLX_EXinst_Mcompar__n0061_inst_cy_119/LOGIC_ZERO ;
  wire DLX_EXinst_Mcompar__n0061_inst_lut4_18;
  wire \DLX_EXinst_Mcompar__n0061_inst_cy_121/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0061_inst_lut4_19;
  wire DLX_EXinst_Mcompar__n0061_inst_cy_120;
  wire \DLX_EXinst_Mcompar__n0061_inst_cy_121/LOGIC_ONE ;
  wire \DLX_EXinst_Mcompar__n0061_inst_cy_121/CYINIT ;
  wire DLX_EXinst_Mcompar__n0061_inst_lut4_20;
  wire \DLX_EXinst_Mcompar__n0061_inst_cy_123/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0061_inst_lut4_21;
  wire DLX_EXinst_Mcompar__n0061_inst_cy_122;
  wire \DLX_EXinst_Mcompar__n0061_inst_cy_123/LOGIC_ONE ;
  wire \DLX_EXinst_Mcompar__n0061_inst_cy_123/CYINIT ;
  wire DLX_EXinst_Mcompar__n0061_inst_lut4_22;
  wire \DLX_MEMinst_opcode_of_WB<0>/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0061_inst_lut4_23;
  wire DLX_EXinst_Mcompar__n0061_inst_cy_124;
  wire \DLX_MEMinst_opcode_of_WB<0>/LOGIC_ONE ;
  wire \DLX_MEMinst_opcode_of_WB<0>/CYINIT ;
  wire DLX_EXinst_Mcompar__n0061_inst_lut4_24;
  wire \DLX_EXinst_Mcompar__n0061_inst_cy_127/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0061_inst_lut4_25;
  wire DLX_EXinst_Mcompar__n0061_inst_cy_126;
  wire \DLX_EXinst_Mcompar__n0061_inst_cy_127/LOGIC_ONE ;
  wire \DLX_EXinst_Mcompar__n0061_inst_cy_127/CYINIT ;
  wire DLX_EXinst_Mcompar__n0061_inst_lut4_26;
  wire \DLX_IDinst_RegFile_23_26/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0061_inst_lut4_27;
  wire DLX_EXinst_Mcompar__n0061_inst_cy_128;
  wire \DLX_IDinst_RegFile_23_26/LOGIC_ONE ;
  wire \DLX_IDinst_RegFile_23_26/CYINIT ;
  wire DLX_EXinst_Mcompar__n0061_inst_lut4_28;
  wire \DLX_EXinst_Mcompar__n0061_inst_cy_131/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0061_inst_lut4_29;
  wire DLX_EXinst_Mcompar__n0061_inst_cy_130;
  wire \DLX_EXinst_Mcompar__n0061_inst_cy_131/LOGIC_ONE ;
  wire \DLX_EXinst_Mcompar__n0061_inst_cy_131/CYINIT ;
  wire DLX_EXinst_Mcompar__n0061_inst_lut4_30;
  wire \DLX_IDinst_RegFile_16_13/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0061_inst_lut4_31;
  wire DLX_EXinst_Mcompar__n0061_inst_cy_132;
  wire \DLX_IDinst_RegFile_16_13/LOGIC_ONE ;
  wire \DLX_IDinst_RegFile_16_13/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_667;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_593/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_668;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_592;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_593/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_593/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_587;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_513/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_588;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_512;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_513/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_513/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_683;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_609/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_684;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_608;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_609/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_609/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_603;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_529/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_604;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_528;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_529/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_529/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_763;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_689/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_764;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_688;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_689/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_689/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_779;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_705/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_780;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_704;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_705/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_705/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_699;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_625/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_700;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_624;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_625/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_625/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_619;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_545/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_620;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_544;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_545/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_545/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_631;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_557/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_632;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_556;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_557/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_557/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_875;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_801/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_876;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_800;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_801/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_801/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_795;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_721/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_796;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_720;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_721/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_721/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_715;
  wire \DLX_EXinst_reg_out_B_EX<5>/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_716;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_640;
  wire \DLX_EXinst_reg_out_B_EX<5>/LOGIC_ZERO ;
  wire \DLX_EXinst_reg_out_B_EX<5>/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_723;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_649/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_724;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_648;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_649/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_649/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_635;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_561/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_636;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_560;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_561/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_561/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_971;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_897/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_972;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_896;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_897/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_897/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_891;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_817/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_892;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_816;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_817/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_817/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_811;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_737/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_812;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_736;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_737/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_737/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_815;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_741/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_816;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_740;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_741/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_741/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_731;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_657/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_732;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_656;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_657/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_657/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_651;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_577/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_652;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_576;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_577/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_577/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_987;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_913/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_988;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_912;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_913/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_913/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_999;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_925/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1000;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_924;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_925/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_925/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_907;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_833/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_908;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_832;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_833/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_833/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_827;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_753/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_828;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_752;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_753/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_753/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_747;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_673/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_748;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_672;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_673/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_673/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1003;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_929/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1004;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_928;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_929/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_929/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_923;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_849/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_924;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_848;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_849/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_849/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_843;
  wire \DLX_MEMinst_opcode_of_WB<4>/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_844;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_768;
  wire \DLX_MEMinst_opcode_of_WB<4>/LOGIC_ZERO ;
  wire \DLX_MEMinst_opcode_of_WB<4>/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_939;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_865/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_940;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_864;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_865/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_865/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_859;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_785/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_860;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_784;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_785/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_785/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1019;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_945/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1020;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_944;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_945/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_945/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_955;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_881/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_956;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_880;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_881/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_881/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1035;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_961/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1036;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_960;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_961/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_961/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1051;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_977/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1052;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_976;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_977/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_977/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1067;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_993/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1068;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_992;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_993/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_993/LOGIC_ONE ;
  wire DLX_EXinst_Maddsub__n0012_inst_lut3_2;
  wire \DLX_IDinst_RegFile_3_16/XORF ;
  wire \DLX_IDinst_RegFile_3_16/CYMUXG ;
  wire \DLX_IDinst_RegFile_3_16/XORG ;
  wire DLX_EXinst_Maddsub__n0012_inst_lut3_3;
  wire DLX_EXinst_Maddsub__n0012_inst_cy_70;
  wire \DLX_IDinst_RegFile_3_16/CYINIT ;
  wire DLX_EXinst_Maddsub__n0012_inst_lut3_4;
  wire \DLX_EXinst__n0012<2>/XORF ;
  wire \DLX_EXinst__n0012<2>/CYMUXG ;
  wire \DLX_EXinst__n0012<2>/XORG ;
  wire DLX_EXinst_Maddsub__n0012_inst_lut3_5;
  wire DLX_EXinst_Maddsub__n0012_inst_cy_72;
  wire \DLX_EXinst__n0012<2>/CYINIT ;
  wire DLX_EXinst_Maddsub__n0012_inst_lut3_6;
  wire \DLX_EXinst__n0012<4>/XORF ;
  wire \DLX_EXinst__n0012<4>/CYMUXG ;
  wire \DLX_EXinst__n0012<4>/XORG ;
  wire DLX_EXinst_Maddsub__n0012_inst_lut3_7;
  wire DLX_EXinst_Maddsub__n0012_inst_cy_74;
  wire \DLX_EXinst__n0012<4>/CYINIT ;
  wire DLX_EXinst_Maddsub__n0012_inst_lut3_8;
  wire \DLX_EXinst__n0012<6>/XORF ;
  wire \DLX_EXinst__n0012<6>/CYMUXG ;
  wire \DLX_EXinst__n0012<6>/XORG ;
  wire DLX_EXinst_Maddsub__n0012_inst_lut3_9;
  wire DLX_EXinst_Maddsub__n0012_inst_cy_76;
  wire \DLX_EXinst__n0012<6>/CYINIT ;
  wire DLX_EXinst_Maddsub__n0012_inst_lut3_10;
  wire \DLX_IDinst_RegFile_26_10/XORF ;
  wire \DLX_IDinst_RegFile_26_10/CYMUXG ;
  wire \DLX_IDinst_RegFile_26_10/XORG ;
  wire DLX_EXinst_Maddsub__n0012_inst_lut3_11;
  wire DLX_EXinst_Maddsub__n0012_inst_cy_78;
  wire \DLX_IDinst_RegFile_26_10/CYINIT ;
  wire DLX_EXinst_Maddsub__n0012_inst_lut3_12;
  wire \DLX_EXinst__n0012<10>/XORF ;
  wire \DLX_EXinst__n0012<10>/CYMUXG ;
  wire \DLX_EXinst__n0012<10>/XORG ;
  wire DLX_EXinst_Maddsub__n0012_inst_lut3_13;
  wire DLX_EXinst_Maddsub__n0012_inst_cy_80;
  wire \DLX_EXinst__n0012<10>/CYINIT ;
  wire DLX_EXinst_Maddsub__n0012_inst_lut3_14;
  wire \DLX_EXinst__n0012<12>/XORF ;
  wire \DLX_EXinst__n0012<12>/CYMUXG ;
  wire \DLX_EXinst__n0012<12>/XORG ;
  wire DLX_EXinst_Maddsub__n0012_inst_lut3_15;
  wire DLX_EXinst_Maddsub__n0012_inst_cy_82;
  wire \DLX_EXinst__n0012<12>/CYINIT ;
  wire DLX_EXinst_Maddsub__n0012_inst_lut3_16;
  wire \DLX_EXinst__n0012<14>/XORF ;
  wire \DLX_EXinst__n0012<14>/CYMUXG ;
  wire \DLX_EXinst__n0012<14>/XORG ;
  wire DLX_EXinst_Maddsub__n0012_inst_lut3_17;
  wire DLX_EXinst_Maddsub__n0012_inst_cy_84;
  wire \DLX_EXinst__n0012<14>/CYINIT ;
  wire DLX_EXinst_Maddsub__n0012_inst_lut3_18;
  wire \DLX_IDinst_RegFile_18_5/XORF ;
  wire \DLX_IDinst_RegFile_18_5/CYMUXG ;
  wire \DLX_IDinst_RegFile_18_5/XORG ;
  wire DLX_EXinst_Maddsub__n0012_inst_lut3_19;
  wire DLX_EXinst_Maddsub__n0012_inst_cy_86;
  wire \DLX_IDinst_RegFile_18_5/CYINIT ;
  wire DLX_EXinst_Maddsub__n0012_inst_lut3_20;
  wire \DLX_EXinst__n0012<18>/XORF ;
  wire \DLX_EXinst__n0012<18>/CYMUXG ;
  wire \DLX_EXinst__n0012<18>/XORG ;
  wire DLX_EXinst_Maddsub__n0012_inst_lut3_21;
  wire DLX_EXinst_Maddsub__n0012_inst_cy_88;
  wire \DLX_EXinst__n0012<18>/CYINIT ;
  wire DLX_EXinst_Maddsub__n0012_inst_lut3_22;
  wire \DLX_EXinst__n0012<20>/XORF ;
  wire \DLX_EXinst__n0012<20>/CYMUXG ;
  wire \DLX_EXinst__n0012<20>/XORG ;
  wire DLX_EXinst_Maddsub__n0012_inst_lut3_23;
  wire DLX_EXinst_Maddsub__n0012_inst_cy_90;
  wire \DLX_EXinst__n0012<20>/CYINIT ;
  wire DLX_EXinst_Maddsub__n0012_inst_lut3_24;
  wire \DLX_EXinst__n0012<22>/XORF ;
  wire \DLX_EXinst__n0012<22>/CYMUXG ;
  wire \DLX_EXinst__n0012<22>/XORG ;
  wire DLX_EXinst_Maddsub__n0012_inst_lut3_25;
  wire DLX_EXinst_Maddsub__n0012_inst_cy_92;
  wire \DLX_EXinst__n0012<22>/CYINIT ;
  wire DLX_EXinst_Maddsub__n0012_inst_lut3_26;
  wire \DLX_IDinst_EPC<29>/XORF ;
  wire \DLX_IDinst_EPC<29>/CYMUXG ;
  wire \DLX_IDinst_EPC<29>/XORG ;
  wire DLX_EXinst_Maddsub__n0012_inst_lut3_27;
  wire DLX_EXinst_Maddsub__n0012_inst_cy_94;
  wire \DLX_IDinst_EPC<29>/CYINIT ;
  wire DLX_EXinst_Maddsub__n0012_inst_lut3_28;
  wire \DLX_EXinst__n0012<26>/XORF ;
  wire \DLX_EXinst__n0012<26>/CYMUXG ;
  wire \DLX_EXinst__n0012<26>/XORG ;
  wire DLX_EXinst_Maddsub__n0012_inst_lut3_29;
  wire DLX_EXinst_Maddsub__n0012_inst_cy_96;
  wire \DLX_EXinst__n0012<26>/CYINIT ;
  wire DLX_EXinst_Maddsub__n0012_inst_lut3_30;
  wire \DLX_EXinst__n0012<28>/XORF ;
  wire \DLX_EXinst__n0012<28>/CYMUXG ;
  wire \DLX_EXinst__n0012<28>/XORG ;
  wire DLX_EXinst_Maddsub__n0012_inst_lut3_31;
  wire DLX_EXinst_Maddsub__n0012_inst_cy_98;
  wire \DLX_EXinst__n0012<28>/CYINIT ;
  wire DLX_EXinst_Maddsub__n0012_inst_lut3_32;
  wire \DLX_EXinst__n0012<30>/XORF ;
  wire \DLX_EXinst__n0012<30>/XORG ;
  wire DLX_EXinst_Maddsub__n0012_inst_lut3_33;
  wire DLX_EXinst_Maddsub__n0012_inst_cy_100;
  wire \DLX_EXinst__n0012<30>/CYINIT ;
  wire DLX_EXinst_Mcompar__n0087_inst_lut4_16;
  wire \DLX_EXinst_Mcompar__n0087_inst_cy_119/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0087_inst_lut4_17;
  wire DLX_EXinst_Mcompar__n0087_inst_cy_118;
  wire \DLX_EXinst_Mcompar__n0087_inst_cy_119/LOGIC_ONE ;
  wire \DLX_EXinst_Mcompar__n0087_inst_cy_119/LOGIC_ZERO ;
  wire DLX_EXinst_Mcompar__n0087_inst_lut4_18;
  wire \DLX_EXinst_Mcompar__n0087_inst_cy_121/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0087_inst_lut4_19;
  wire DLX_EXinst_Mcompar__n0087_inst_cy_120;
  wire \DLX_EXinst_Mcompar__n0087_inst_cy_121/LOGIC_ONE ;
  wire \DLX_EXinst_Mcompar__n0087_inst_cy_121/CYINIT ;
  wire DLX_EXinst_Mcompar__n0087_inst_lut4_20;
  wire \DLX_EXinst_Mcompar__n0087_inst_cy_123/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0087_inst_lut4_21;
  wire DLX_EXinst_Mcompar__n0087_inst_cy_122;
  wire \DLX_EXinst_Mcompar__n0087_inst_cy_123/LOGIC_ONE ;
  wire \DLX_EXinst_Mcompar__n0087_inst_cy_123/CYINIT ;
  wire DLX_EXinst_Mcompar__n0087_inst_lut4_22;
  wire \DLX_EXinst_Mcompar__n0087_inst_cy_125/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0087_inst_lut4_23;
  wire DLX_EXinst_Mcompar__n0087_inst_cy_124;
  wire \DLX_EXinst_Mcompar__n0087_inst_cy_125/LOGIC_ONE ;
  wire \DLX_EXinst_Mcompar__n0087_inst_cy_125/CYINIT ;
  wire DLX_EXinst_Mcompar__n0087_inst_lut4_24;
  wire \DLX_EXinst_Mcompar__n0087_inst_cy_127/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0087_inst_lut4_25;
  wire DLX_EXinst_Mcompar__n0087_inst_cy_126;
  wire \DLX_EXinst_Mcompar__n0087_inst_cy_127/LOGIC_ONE ;
  wire \DLX_EXinst_Mcompar__n0087_inst_cy_127/CYINIT ;
  wire DLX_EXinst_Mcompar__n0087_inst_lut4_26;
  wire \DLX_EXinst_Mcompar__n0087_inst_cy_129/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0087_inst_lut4_27;
  wire DLX_EXinst_Mcompar__n0087_inst_cy_128;
  wire \DLX_EXinst_Mcompar__n0087_inst_cy_129/LOGIC_ONE ;
  wire \DLX_EXinst_Mcompar__n0087_inst_cy_129/CYINIT ;
  wire DLX_EXinst_Mcompar__n0087_inst_lut4_28;
  wire \DLX_EXinst_Mcompar__n0087_inst_cy_131/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0087_inst_lut4_29;
  wire DLX_EXinst_Mcompar__n0087_inst_cy_130;
  wire \DLX_EXinst_Mcompar__n0087_inst_cy_131/LOGIC_ONE ;
  wire \DLX_EXinst_Mcompar__n0087_inst_cy_131/CYINIT ;
  wire DLX_EXinst_Mcompar__n0087_inst_lut4_30;
  wire \DLX_EXinst__n0087/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0087_inst_lut4_31;
  wire DLX_EXinst_Mcompar__n0087_inst_cy_132;
  wire \DLX_EXinst__n0087/LOGIC_ONE ;
  wire \DLX_EXinst__n0087/CYINIT ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_166;
  wire \DLX_IDinst_RegFile_2_25/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_167;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_230;
  wire \DLX_IDinst_RegFile_2_25/LOGIC_ZERO ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_168;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_233/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_169;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_232;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_233/CYINIT ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_170;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_235/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_171;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_234;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_235/CYINIT ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_172;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_237/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_173;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_236;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_237/CYINIT ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_174;
  wire \DLX_IFinst_IR_curr<15>/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_175;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_238;
  wire \DLX_IFinst_IR_curr<15>/CYINIT ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_176;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_241/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_177;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_240;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_241/CYINIT ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_178;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_243/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_179;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_242;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_243/CYINIT ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_180;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_245/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_181;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_244;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_245/CYINIT ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_182;
  wire \DLX_IFinst_IR_curr<4>/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_183;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_246;
  wire \DLX_IFinst_IR_curr<4>/CYINIT ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_184;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_249/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_185;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_248;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_249/CYINIT ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_186;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_251/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_187;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_250;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_251/CYINIT ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_188;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_253/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_189;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_252;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_253/CYINIT ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_190;
  wire \DLX_IFinst_IR_curr<31>/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_191;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_254;
  wire \DLX_IFinst_IR_curr<31>/CYINIT ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_192;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_257/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_193;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_256;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_257/CYINIT ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_194;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_259/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0095_inst_lut2_195;
  wire DLX_EXinst_Mcompar__n0095_inst_cy_258;
  wire \DLX_EXinst_Mcompar__n0095_inst_cy_259/CYINIT ;
  wire \DLX_IDinst_Madd__n0158_inst_lut2_230/FROM ;
  wire \DLX_IDinst_Madd__n0158_inst_lut2_230/CYMUXG ;
  wire \DLX_IDinst_Madd__n0158_inst_lut2_230/XORG ;
  wire DLX_IDinst_Madd__n0158_inst_lut2_231;
  wire DLX_IDinst_Madd__n0158_inst_cy_297;
  wire \DLX_IDinst_Madd__n0158_inst_lut2_230/LOGIC_ZERO ;
  wire DLX_IDinst_Madd__n0158_inst_lut2_232;
  wire \DLX_IDinst_RegFile_2_30/XORF ;
  wire \DLX_IDinst_RegFile_2_30/CYMUXG ;
  wire \DLX_IDinst_RegFile_2_30/XORG ;
  wire DLX_IDinst_Madd__n0158_inst_lut2_233;
  wire DLX_IDinst_Madd__n0158_inst_cy_299;
  wire \DLX_IDinst_RegFile_2_30/CYINIT ;
  wire DLX_IDinst_Madd__n0158_inst_lut2_234;
  wire \DLX_IDinst__n0158<4>/XORF ;
  wire \DLX_IDinst__n0158<4>/CYMUXG ;
  wire \DLX_IDinst__n0158<4>/XORG ;
  wire DLX_IDinst_Madd__n0158_inst_lut2_235;
  wire DLX_IDinst_Madd__n0158_inst_cy_301;
  wire \DLX_IDinst__n0158<4>/CYINIT ;
  wire DLX_IDinst_Madd__n0158_inst_lut2_236;
  wire \DLX_IDinst__n0158<6>/XORF ;
  wire \DLX_IDinst__n0158<6>/CYMUXG ;
  wire \DLX_IDinst__n0158<6>/XORG ;
  wire DLX_IDinst_Madd__n0158_inst_lut2_237;
  wire DLX_IDinst_Madd__n0158_inst_cy_303;
  wire \DLX_IDinst__n0158<6>/CYINIT ;
  wire DLX_IDinst_Madd__n0158_inst_lut2_238;
  wire \DLX_IDinst__n0158<8>/XORF ;
  wire \DLX_IDinst__n0158<8>/CYMUXG ;
  wire \DLX_IDinst__n0158<8>/XORG ;
  wire DLX_IDinst_Madd__n0158_inst_lut2_239;
  wire DLX_IDinst_Madd__n0158_inst_cy_305;
  wire \DLX_IDinst__n0158<8>/CYINIT ;
  wire DLX_IDinst_Madd__n0158_inst_lut2_240;
  wire \DLX_IFinst_IR_curr<24>/XORF ;
  wire \DLX_IFinst_IR_curr<24>/CYMUXG ;
  wire \DLX_IFinst_IR_curr<24>/XORG ;
  wire DLX_IDinst_Madd__n0158_inst_lut2_241;
  wire DLX_IDinst_Madd__n0158_inst_cy_307;
  wire \DLX_IFinst_IR_curr<24>/CYINIT ;
  wire DLX_IDinst_Madd__n0158_inst_lut2_242;
  wire \DLX_IDinst__n0158<12>/XORF ;
  wire \DLX_IDinst__n0158<12>/CYMUXG ;
  wire \DLX_IDinst__n0158<12>/XORG ;
  wire DLX_IDinst_Madd__n0158_inst_lut2_243;
  wire DLX_IDinst_Madd__n0158_inst_cy_309;
  wire \DLX_IDinst__n0158<12>/CYINIT ;
  wire DLX_IDinst_Madd__n0158_inst_lut2_244;
  wire \DLX_IDinst__n0158<14>/XORF ;
  wire \DLX_IDinst__n0158<14>/CYMUXG ;
  wire \DLX_IDinst__n0158<14>/XORG ;
  wire DLX_IDinst_Madd__n0158_inst_lut2_245;
  wire DLX_IDinst_Madd__n0158_inst_cy_311;
  wire \DLX_IDinst__n0158<14>/CYINIT ;
  wire DLX_IDinst_Madd__n0158_inst_lut2_246;
  wire \DLX_IDinst__n0158<16>/XORF ;
  wire \DLX_IDinst__n0158<16>/CYMUXG ;
  wire \DLX_IDinst__n0158<16>/XORG ;
  wire DLX_IDinst_Madd__n0158_inst_lut2_247;
  wire DLX_IDinst_Madd__n0158_inst_cy_313;
  wire \DLX_IDinst__n0158<16>/CYINIT ;
  wire DLX_IDinst_Madd__n0158_inst_lut2_248;
  wire \DLX_IDinst_RegFile_0_6/XORF ;
  wire \DLX_IDinst_RegFile_0_6/CYMUXG ;
  wire \DLX_IDinst_RegFile_0_6/XORG ;
  wire DLX_IDinst_Madd__n0158_inst_lut2_249;
  wire DLX_IDinst_Madd__n0158_inst_cy_315;
  wire \DLX_IDinst_RegFile_0_6/CYINIT ;
  wire DLX_IDinst_Madd__n0158_inst_lut2_250;
  wire \DLX_IDinst__n0158<20>/XORF ;
  wire \DLX_IDinst__n0158<20>/CYMUXG ;
  wire \DLX_IDinst__n0158<20>/XORG ;
  wire DLX_IDinst_Madd__n0158_inst_lut2_251;
  wire DLX_IDinst_Madd__n0158_inst_cy_317;
  wire \DLX_IDinst__n0158<20>/CYINIT ;
  wire DLX_IDinst_Madd__n0158_inst_lut2_252;
  wire \DLX_IDinst__n0158<22>/XORF ;
  wire \DLX_IDinst__n0158<22>/CYMUXG ;
  wire \DLX_IDinst__n0158<22>/XORG ;
  wire DLX_IDinst_Madd__n0158_inst_lut2_253;
  wire DLX_IDinst_Madd__n0158_inst_cy_319;
  wire \DLX_IDinst__n0158<22>/CYINIT ;
  wire DLX_IDinst_Madd__n0158_inst_lut2_254;
  wire \DLX_IDinst__n0158<24>/XORF ;
  wire \DLX_IDinst__n0158<24>/CYMUXG ;
  wire \DLX_IDinst__n0158<24>/XORG ;
  wire DLX_IDinst_Madd__n0158_inst_lut2_255;
  wire DLX_IDinst_Madd__n0158_inst_cy_321;
  wire \DLX_IDinst__n0158<24>/CYINIT ;
  wire DLX_IDinst_Madd__n0158_inst_lut2_256;
  wire \DLX_IFinst_IR_curr<16>/XORF ;
  wire \DLX_IFinst_IR_curr<16>/CYMUXG ;
  wire \DLX_IFinst_IR_curr<16>/XORG ;
  wire DLX_IDinst_Madd__n0158_inst_lut2_257;
  wire DLX_IDinst_Madd__n0158_inst_cy_323;
  wire \DLX_IFinst_IR_curr<16>/CYINIT ;
  wire DLX_IDinst_Madd__n0158_inst_lut2_258;
  wire \DLX_IDinst__n0158<28>/XORF ;
  wire \DLX_IDinst__n0158<28>/CYMUXG ;
  wire \DLX_IDinst__n0158<28>/XORG ;
  wire DLX_IDinst_Madd__n0158_inst_lut2_259;
  wire DLX_IDinst_Madd__n0158_inst_cy_325;
  wire \DLX_IDinst__n0158<28>/CYINIT ;
  wire DLX_IDinst_Madd__n0158_inst_lut2_260;
  wire \DLX_IDinst__n0158<30>/XORF ;
  wire \DLX_IDinst__n0158<30>/XORG ;
  wire DLX_IDinst_Madd__n0158_inst_lut2_261;
  wire DLX_IDinst_Madd__n0158_inst_cy_327;
  wire \DLX_IDinst__n0158<30>/CYINIT ;
  wire DLX_IDinst_Mcompar__n0102_inst_lut4_40;
  wire \DLX_IDinst_Mcompar__n0102_inst_cy_263/CYMUXG ;
  wire DLX_IDinst_Mcompar__n0102_inst_lut4_41;
  wire DLX_IDinst_Mcompar__n0102_inst_cy_262;
  wire \DLX_IDinst_Mcompar__n0102_inst_cy_263/LOGIC_ZERO ;
  wire \DLX_IDinst_Mcompar__n0102_inst_cy_263/LOGIC_ONE ;
  wire \DLX_IDinst__n0102/LOGIC_ZERO ;
  wire DLX_IDinst_Mcompar__n0102_inst_lut4_42;
  wire \DLX_IDinst__n0102/CYMUXF ;
  wire \DLX_IDinst__n0102/CYINIT ;
  wire vga_top_vga1_Mcompar__n0033_inst_lut1_4;
  wire \DLX_IDinst_RegFile_2_18/CYMUXG ;
  wire vga_top_vga1_Mcompar__n0033_inst_lut1_5;
  wire vga_top_vga1_Mcompar__n0033_inst_cy_340;
  wire \DLX_IDinst_RegFile_2_18/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_2_18/LOGIC_ONE ;
  wire vga_top_vga1_Mcompar__n0033_inst_lut2_269;
  wire \vga_top_vga1_Mcompar__n0033_inst_cy_343/CYMUXG ;
  wire vga_top_vga1_Mcompar__n0033_inst_lut2_270;
  wire vga_top_vga1_Mcompar__n0033_inst_cy_342;
  wire \vga_top_vga1_Mcompar__n0033_inst_cy_343/LOGIC_ONE ;
  wire \vga_top_vga1_Mcompar__n0033_inst_cy_343/CYINIT ;
  wire vga_top_vga1_Mcompar__n0033_inst_lut3_98;
  wire \vga_top_vga1_Mcompar__n0033_inst_cy_345/CYMUXG ;
  wire vga_top_vga1_Mcompar__n0033_inst_lut3_99;
  wire vga_top_vga1_Mcompar__n0033_inst_cy_344;
  wire \vga_top_vga1_Mcompar__n0033_inst_cy_345/LOGIC_ZERO ;
  wire \vga_top_vga1_Mcompar__n0033_inst_cy_345/CYINIT ;
  wire vga_top_vga1_Mcompar__n0033_inst_lut2_271;
  wire \vga_top_vga1_Mcompar__n0033_inst_cy_347/CYMUXG ;
  wire vga_top_vga1_Mcompar__n0033_inst_lut2_272;
  wire vga_top_vga1_Mcompar__n0033_inst_cy_346;
  wire \vga_top_vga1_Mcompar__n0033_inst_cy_347/LOGIC_ONE ;
  wire \vga_top_vga1_Mcompar__n0033_inst_cy_347/CYINIT ;
  wire vga_top_vga1_Mcompar__n0033_inst_lut1_6;
  wire \DLX_IFinst_IR_curr<25>/CYMUXG ;
  wire vga_top_vga1_Mcompar__n0033_inst_lut1_7;
  wire vga_top_vga1_Mcompar__n0033_inst_cy_348;
  wire \DLX_IFinst_IR_curr<25>/LOGIC_ZERO ;
  wire \DLX_IFinst_IR_curr<25>/CYINIT ;
  wire \$SIG_13 ;
  wire \vga_top_vga1_Mcompar__n0033_inst_cy_351/CYMUXG ;
  wire \$SIG_14 ;
  wire vga_top_vga1_Mcompar__n0033_inst_cy_350;
  wire \vga_top_vga1_Mcompar__n0033_inst_cy_351/LOGIC_ONE ;
  wire \vga_top_vga1_Mcompar__n0033_inst_cy_351/CYINIT ;
  wire vga_top_vga1_Mcompar__n0033_inst_lut4_1100;
  wire \vga_top_vga1__n0033/CYMUXG ;
  wire vga_top_vga1_Mcompar__n0033_inst_lut2_273;
  wire vga_top_vga1_Mcompar__n0033_inst_cy_352;
  wire \vga_top_vga1__n0033/LOGIC_ZERO ;
  wire \vga_top_vga1__n0033/CYINIT ;
  wire \vga_top_vga1_Madd_addressout_inst_lut2_331/FROM ;
  wire \vga_top_vga1_Madd_addressout_inst_lut2_331/CYMUXG ;
  wire \vga_top_vga1_Madd_addressout_inst_lut2_331/XORG ;
  wire vga_top_vga1_Madd_addressout_inst_lut2_332;
  wire vga_top_vga1_Madd_addressout_inst_cy_462;
  wire \vga_top_vga1_Madd_addressout_inst_lut2_331/LOGIC_ZERO ;
  wire vga_top_vga1_Madd_addressout_inst_lut2_333;
  wire \vga_address<7>/XORF ;
  wire \vga_address<7>/CYMUXG ;
  wire \vga_address<7>/XORG ;
  wire vga_top_vga1_Madd_addressout_inst_lut2_334;
  wire vga_top_vga1_Madd_addressout_inst_cy_464;
  wire \vga_address<7>/CYINIT ;
  wire \vga_address<9>/FROM ;
  wire \vga_address<9>/XORF ;
  wire \vga_address<9>/CYMUXG ;
  wire \vga_address<9>/LOGIC_ZERO ;
  wire \vga_address<9>/XORG ;
  wire \vga_address<9>/GROM ;
  wire vga_top_vga1_Madd_addressout_inst_cy_466;
  wire \vga_address<9>/CYINIT ;
  wire \vga_address<11>/FROM ;
  wire \vga_address<11>/XORF ;
  wire \vga_address<11>/CYMUXG ;
  wire \vga_address<11>/LOGIC_ZERO ;
  wire \vga_address<11>/XORG ;
  wire \vga_address<11>/GROM ;
  wire vga_top_vga1_Madd_addressout_inst_cy_468;
  wire \vga_address<11>/CYINIT ;
  wire \vga_address<13>/LOGIC_ZERO ;
  wire \vga_address<13>/FROM ;
  wire \vga_address<13>/XORF ;
  wire \vga_address<13>/XORG ;
  wire vga_top_vga1_Mmult__n0043_inst_lut2_323_rt;
  wire vga_top_vga1_Madd_addressout_inst_cy_470;
  wire \vga_address<13>/CYINIT ;
  wire DLX_IFinst_Madd__n0005_inst_lut2_40;
  wire \DLX_IFinst__n0015<3>/CYMUXG ;
  wire \DLX_IFinst__n0015<3>/XORG ;
  wire \DLX_IFinst__n0015<3>/GROM ;
  wire DLX_IFinst_Madd__n0005_inst_cy_40;
  wire \DLX_IFinst__n0015<3>/LOGIC_ZERO ;
  wire \DLX_IFinst__n0015<4>/FROM ;
  wire \DLX_IFinst__n0015<4>/XORF ;
  wire \DLX_IFinst__n0015<4>/CYMUXG ;
  wire \DLX_IFinst__n0015<4>/LOGIC_ZERO ;
  wire \DLX_IFinst__n0015<4>/XORG ;
  wire \DLX_IFinst__n0015<4>/GROM ;
  wire DLX_IFinst_Madd__n0005_inst_cy_42;
  wire \DLX_IFinst__n0015<4>/CYINIT ;
  wire \DLX_IFinst__n0015<6>/FROM ;
  wire \DLX_IFinst__n0015<6>/XORF ;
  wire \DLX_IFinst__n0015<6>/CYMUXG ;
  wire \DLX_IFinst__n0015<6>/LOGIC_ZERO ;
  wire \DLX_IFinst__n0015<6>/XORG ;
  wire \DLX_IFinst__n0015<6>/GROM ;
  wire DLX_IFinst_Madd__n0005_inst_cy_44;
  wire \DLX_IFinst__n0015<6>/CYINIT ;
  wire \DLX_IFinst__n0015<8>/FROM ;
  wire \DLX_IFinst__n0015<8>/XORF ;
  wire \DLX_IFinst__n0015<8>/CYMUXG ;
  wire \DLX_IFinst__n0015<8>/LOGIC_ZERO ;
  wire \DLX_IFinst__n0015<8>/XORG ;
  wire \DLX_IFinst__n0015<8>/GROM ;
  wire DLX_IFinst_Madd__n0005_inst_cy_46;
  wire \DLX_IFinst__n0015<8>/CYINIT ;
  wire \DLX_IFinst__n0015<10>/FROM ;
  wire \DLX_IFinst__n0015<10>/XORF ;
  wire \DLX_IFinst__n0015<10>/CYMUXG ;
  wire \DLX_IFinst__n0015<10>/LOGIC_ZERO ;
  wire \DLX_IFinst__n0015<10>/XORG ;
  wire \DLX_IFinst__n0015<10>/GROM ;
  wire DLX_IFinst_Madd__n0005_inst_cy_48;
  wire \DLX_IFinst__n0015<10>/CYINIT ;
  wire \DLX_IFinst__n0015<12>/FROM ;
  wire \DLX_IFinst__n0015<12>/XORF ;
  wire \DLX_IFinst__n0015<12>/CYMUXG ;
  wire \DLX_IFinst__n0015<12>/LOGIC_ZERO ;
  wire \DLX_IFinst__n0015<12>/XORG ;
  wire \DLX_IFinst__n0015<12>/GROM ;
  wire DLX_IFinst_Madd__n0005_inst_cy_50;
  wire \DLX_IFinst__n0015<12>/CYINIT ;
  wire \DLX_IFinst__n0015<14>/FROM ;
  wire \DLX_IFinst__n0015<14>/XORF ;
  wire \DLX_IFinst__n0015<14>/CYMUXG ;
  wire \DLX_IFinst__n0015<14>/LOGIC_ZERO ;
  wire \DLX_IFinst__n0015<14>/XORG ;
  wire \DLX_IFinst__n0015<14>/GROM ;
  wire DLX_IFinst_Madd__n0005_inst_cy_52;
  wire \DLX_IFinst__n0015<14>/CYINIT ;
  wire \DLX_IFinst__n0015<16>/FROM ;
  wire \DLX_IFinst__n0015<16>/XORF ;
  wire \DLX_IFinst__n0015<16>/CYMUXG ;
  wire \DLX_IFinst__n0015<16>/LOGIC_ZERO ;
  wire \DLX_IFinst__n0015<16>/XORG ;
  wire \DLX_IFinst__n0015<16>/GROM ;
  wire DLX_IFinst_Madd__n0005_inst_cy_54;
  wire \DLX_IFinst__n0015<16>/CYINIT ;
  wire \DLX_IFinst__n0015<18>/FROM ;
  wire \DLX_IFinst__n0015<18>/XORF ;
  wire \DLX_IFinst__n0015<18>/CYMUXG ;
  wire \DLX_IFinst__n0015<18>/LOGIC_ZERO ;
  wire \DLX_IFinst__n0015<18>/XORG ;
  wire \DLX_IFinst__n0015<18>/GROM ;
  wire DLX_IFinst_Madd__n0005_inst_cy_56;
  wire \DLX_IFinst__n0015<18>/CYINIT ;
  wire \DLX_IFinst__n0015<20>/FROM ;
  wire \DLX_IFinst__n0015<20>/XORF ;
  wire \DLX_IFinst__n0015<20>/CYMUXG ;
  wire \DLX_IFinst__n0015<20>/LOGIC_ZERO ;
  wire \DLX_IFinst__n0015<20>/XORG ;
  wire \DLX_IFinst__n0015<20>/GROM ;
  wire DLX_IFinst_Madd__n0005_inst_cy_58;
  wire \DLX_IFinst__n0015<20>/CYINIT ;
  wire \DLX_IFinst__n0015<22>/FROM ;
  wire \DLX_IFinst__n0015<22>/XORF ;
  wire \DLX_IFinst__n0015<22>/CYMUXG ;
  wire \DLX_IFinst__n0015<22>/LOGIC_ZERO ;
  wire \DLX_IFinst__n0015<22>/XORG ;
  wire \DLX_IFinst__n0015<22>/GROM ;
  wire DLX_IFinst_Madd__n0005_inst_cy_60;
  wire \DLX_IFinst__n0015<22>/CYINIT ;
  wire \DLX_IFinst__n0015<24>/FROM ;
  wire \DLX_IFinst__n0015<24>/XORF ;
  wire \DLX_IFinst__n0015<24>/CYMUXG ;
  wire \DLX_IFinst__n0015<24>/LOGIC_ZERO ;
  wire \DLX_IFinst__n0015<24>/XORG ;
  wire \DLX_IFinst__n0015<24>/GROM ;
  wire DLX_IFinst_Madd__n0005_inst_cy_62;
  wire \DLX_IFinst__n0015<24>/CYINIT ;
  wire \DLX_IFinst__n0015<26>/FROM ;
  wire \DLX_IFinst__n0015<26>/XORF ;
  wire \DLX_IFinst__n0015<26>/CYMUXG ;
  wire \DLX_IFinst__n0015<26>/LOGIC_ZERO ;
  wire \DLX_IFinst__n0015<26>/XORG ;
  wire \DLX_IFinst__n0015<26>/GROM ;
  wire DLX_IFinst_Madd__n0005_inst_cy_64;
  wire \DLX_IFinst__n0015<26>/CYINIT ;
  wire \DLX_IFinst__n0015<28>/FROM ;
  wire \DLX_IFinst__n0015<28>/XORF ;
  wire \DLX_IFinst__n0015<28>/CYMUXG ;
  wire \DLX_IFinst__n0015<28>/LOGIC_ZERO ;
  wire \DLX_IFinst__n0015<28>/XORG ;
  wire \DLX_IFinst__n0015<28>/GROM ;
  wire DLX_IFinst_Madd__n0005_inst_cy_66;
  wire \DLX_IFinst__n0015<28>/CYINIT ;
  wire \DLX_IFinst__n0015<30>/LOGIC_ZERO ;
  wire \DLX_IFinst__n0015<30>/FROM ;
  wire \DLX_IFinst__n0015<30>/XORF ;
  wire \DLX_IFinst__n0015<30>/XORG ;
  wire \DLX_IFinst_NPC<31>_rt ;
  wire DLX_IFinst_Madd__n0005_inst_cy_68;
  wire \DLX_IFinst__n0015<30>/CYINIT ;
  wire DLX_EXinst_Mcompar__n0085_inst_lut4_0;
  wire \DLX_EXinst_Mcompar__n0085_inst_cy_103/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0085_inst_lut4_1;
  wire DLX_EXinst_Mcompar__n0085_inst_cy_102;
  wire \DLX_EXinst_Mcompar__n0085_inst_cy_103/LOGIC_ZERO ;
  wire \DLX_EXinst_Mcompar__n0085_inst_cy_103/LOGIC_ONE ;
  wire DLX_EXinst_Mcompar__n0085_inst_lut4_2;
  wire \DLX_EXinst_Mcompar__n0085_inst_cy_105/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0085_inst_lut4_3;
  wire DLX_EXinst_Mcompar__n0085_inst_cy_104;
  wire \DLX_EXinst_Mcompar__n0085_inst_cy_105/LOGIC_ZERO ;
  wire \DLX_EXinst_Mcompar__n0085_inst_cy_105/CYINIT ;
  wire DLX_EXinst_Mcompar__n0085_inst_lut4_4;
  wire \DLX_EXinst_Mcompar__n0085_inst_cy_107/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0085_inst_lut4_5;
  wire DLX_EXinst_Mcompar__n0085_inst_cy_106;
  wire \DLX_EXinst_Mcompar__n0085_inst_cy_107/LOGIC_ZERO ;
  wire \DLX_EXinst_Mcompar__n0085_inst_cy_107/CYINIT ;
  wire DLX_EXinst_Mcompar__n0085_inst_lut4_6;
  wire \DLX_EXinst_Mcompar__n0085_inst_cy_109/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0085_inst_lut4_7;
  wire DLX_EXinst_Mcompar__n0085_inst_cy_108;
  wire \DLX_EXinst_Mcompar__n0085_inst_cy_109/LOGIC_ZERO ;
  wire \DLX_EXinst_Mcompar__n0085_inst_cy_109/CYINIT ;
  wire DLX_EXinst_Mcompar__n0085_inst_lut4_8;
  wire \DLX_EXinst_Mcompar__n0085_inst_cy_111/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0085_inst_lut4_9;
  wire DLX_EXinst_Mcompar__n0085_inst_cy_110;
  wire \DLX_EXinst_Mcompar__n0085_inst_cy_111/LOGIC_ZERO ;
  wire \DLX_EXinst_Mcompar__n0085_inst_cy_111/CYINIT ;
  wire DLX_EXinst_Mcompar__n0085_inst_lut4_10;
  wire \DLX_EXinst_Mcompar__n0085_inst_cy_113/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0085_inst_lut4_11;
  wire DLX_EXinst_Mcompar__n0085_inst_cy_112;
  wire \DLX_EXinst_Mcompar__n0085_inst_cy_113/LOGIC_ZERO ;
  wire \DLX_EXinst_Mcompar__n0085_inst_cy_113/CYINIT ;
  wire DLX_EXinst_Mcompar__n0085_inst_lut4_12;
  wire \DLX_EXinst_Mcompar__n0085_inst_cy_115/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0085_inst_lut4_13;
  wire DLX_EXinst_Mcompar__n0085_inst_cy_114;
  wire \DLX_EXinst_Mcompar__n0085_inst_cy_115/LOGIC_ZERO ;
  wire \DLX_EXinst_Mcompar__n0085_inst_cy_115/CYINIT ;
  wire DLX_EXinst_Mcompar__n0085_inst_lut4_14;
  wire \DLX_EXinst__n0085/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0085_inst_lut4_15;
  wire DLX_EXinst_Mcompar__n0085_inst_cy_116;
  wire \DLX_EXinst__n0085/LOGIC_ZERO ;
  wire \DLX_EXinst__n0085/CYINIT ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_134;
  wire \DLX_IDinst_RegFile_1_19/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_135;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_198;
  wire \DLX_IDinst_RegFile_1_19/LOGIC_ZERO ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_136;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_201/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_137;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_200;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_201/CYINIT ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_138;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_203/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_139;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_202;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_203/CYINIT ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_140;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_205/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_141;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_204;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_205/CYINIT ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_142;
  wire \DLX_IDinst_RegFile_23_2/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_143;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_206;
  wire \DLX_IDinst_RegFile_23_2/CYINIT ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_144;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_209/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_145;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_208;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_209/CYINIT ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_146;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_211/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_147;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_210;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_211/CYINIT ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_148;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_213/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_149;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_212;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_213/CYINIT ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_150;
  wire \DLX_IDinst_RegFile_3_18/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_151;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_214;
  wire \DLX_IDinst_RegFile_3_18/CYINIT ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_152;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_217/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_153;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_216;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_217/CYINIT ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_154;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_219/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_155;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_218;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_219/CYINIT ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_156;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_221/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_157;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_220;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_221/CYINIT ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_158;
  wire \DLX_IFinst_IR_curr<6>/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_159;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_222;
  wire \DLX_IFinst_IR_curr<6>/CYINIT ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_160;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_225/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_161;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_224;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_225/CYINIT ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_162;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_227/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_163;
  wire DLX_EXinst_Mcompar__n0093_inst_cy_226;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_227/CYINIT ;
  wire DLX_EXinst_Mcompar__n0093_inst_lut2_164;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_228/CYMUXF ;
  wire \DLX_EXinst_Mcompar__n0093_inst_cy_228/CYINIT ;
  wire DLX_EXinst_Mcompar__n0069_inst_lut2_166;
  wire \DLX_EXinst_Mcompar__n0069_inst_cy_231/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0069_inst_lut2_167;
  wire DLX_EXinst_Mcompar__n0069_inst_cy_230;
  wire \DLX_EXinst_Mcompar__n0069_inst_cy_231/LOGIC_ZERO ;
  wire DLX_EXinst_Mcompar__n0069_inst_lut2_168;
  wire \DLX_IDinst_RegFile_2_26/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0069_inst_lut2_169;
  wire DLX_EXinst_Mcompar__n0069_inst_cy_232;
  wire \DLX_IDinst_RegFile_2_26/CYINIT ;
  wire DLX_EXinst_Mcompar__n0069_inst_lut2_170;
  wire \DLX_EXinst_Mcompar__n0069_inst_cy_235/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0069_inst_lut2_171;
  wire DLX_EXinst_Mcompar__n0069_inst_cy_234;
  wire \DLX_EXinst_Mcompar__n0069_inst_cy_235/CYINIT ;
  wire DLX_EXinst_Mcompar__n0069_inst_lut2_172;
  wire \DLX_EXinst_Mcompar__n0069_inst_cy_237/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0069_inst_lut2_173;
  wire DLX_EXinst_Mcompar__n0069_inst_cy_236;
  wire \DLX_EXinst_Mcompar__n0069_inst_cy_237/CYINIT ;
  wire DLX_EXinst_Mcompar__n0069_inst_lut2_174;
  wire \DLX_EXinst_Mcompar__n0069_inst_cy_239/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0069_inst_lut2_175;
  wire DLX_EXinst_Mcompar__n0069_inst_cy_238;
  wire \DLX_EXinst_Mcompar__n0069_inst_cy_239/CYINIT ;
  wire DLX_EXinst_Mcompar__n0069_inst_lut2_176;
  wire \DLX_IFinst_IR_curr<27>/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0069_inst_lut2_177;
  wire DLX_EXinst_Mcompar__n0069_inst_cy_240;
  wire \DLX_IFinst_IR_curr<27>/CYINIT ;
  wire DLX_EXinst_Mcompar__n0069_inst_lut2_178;
  wire \DLX_EXinst_Mcompar__n0069_inst_cy_243/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0069_inst_lut2_179;
  wire DLX_EXinst_Mcompar__n0069_inst_cy_242;
  wire \DLX_EXinst_Mcompar__n0069_inst_cy_243/CYINIT ;
  wire DLX_EXinst_Mcompar__n0069_inst_lut2_180;
  wire \DLX_EXinst_Mcompar__n0069_inst_cy_245/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0069_inst_lut2_181;
  wire DLX_EXinst_Mcompar__n0069_inst_cy_244;
  wire \DLX_EXinst_Mcompar__n0069_inst_cy_245/CYINIT ;
  wire DLX_EXinst_Mcompar__n0069_inst_lut2_182;
  wire \DLX_EXinst_Mcompar__n0069_inst_cy_247/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0069_inst_lut2_183;
  wire DLX_EXinst_Mcompar__n0069_inst_cy_246;
  wire \DLX_EXinst_Mcompar__n0069_inst_cy_247/CYINIT ;
  wire DLX_EXinst_Mcompar__n0069_inst_lut2_184;
  wire \DLX_IDinst_RegFile_3_26/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0069_inst_lut2_185;
  wire DLX_EXinst_Mcompar__n0069_inst_cy_248;
  wire \DLX_IDinst_RegFile_3_26/CYINIT ;
  wire DLX_EXinst_Mcompar__n0069_inst_lut2_186;
  wire \DLX_EXinst_Mcompar__n0069_inst_cy_251/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0069_inst_lut2_187;
  wire DLX_EXinst_Mcompar__n0069_inst_cy_250;
  wire \DLX_EXinst_Mcompar__n0069_inst_cy_251/CYINIT ;
  wire DLX_EXinst_Mcompar__n0069_inst_lut2_188;
  wire \DLX_EXinst_Mcompar__n0069_inst_cy_253/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0069_inst_lut2_189;
  wire DLX_EXinst_Mcompar__n0069_inst_cy_252;
  wire \DLX_EXinst_Mcompar__n0069_inst_cy_253/CYINIT ;
  wire DLX_EXinst_Mcompar__n0069_inst_lut2_190;
  wire \DLX_EXinst_Mcompar__n0069_inst_cy_255/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0069_inst_lut2_191;
  wire DLX_EXinst_Mcompar__n0069_inst_cy_254;
  wire \DLX_EXinst_Mcompar__n0069_inst_cy_255/CYINIT ;
  wire DLX_EXinst_Mcompar__n0069_inst_lut2_192;
  wire \DLX_IFinst_IR_curr<19>/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0069_inst_lut2_193;
  wire DLX_EXinst_Mcompar__n0069_inst_cy_256;
  wire \DLX_IFinst_IR_curr<19>/CYINIT ;
  wire DLX_EXinst_Mcompar__n0069_inst_lut2_194;
  wire \DLX_EXinst_Mcompar__n0069_inst_cy_259/CYMUXG ;
  wire DLX_EXinst_Mcompar__n0069_inst_lut2_195;
  wire DLX_EXinst_Mcompar__n0069_inst_cy_258;
  wire \DLX_EXinst_Mcompar__n0069_inst_cy_259/CYINIT ;
  wire DLX_EXinst_Mcompar__n0069_inst_lut2_196;
  wire \DLX_EXinst_Mcompar__n0069_inst_cy_260/CYMUXF ;
  wire \DLX_EXinst_Mcompar__n0069_inst_cy_260/CYINIT ;
  wire DLX_IDinst_Mcompar__n0100_inst_lut4_40;
  wire \DLX_IDinst_Mcompar__n0100_inst_cy_263/CYMUXG ;
  wire DLX_IDinst_Mcompar__n0100_inst_lut4_41;
  wire DLX_IDinst_Mcompar__n0100_inst_cy_262;
  wire \DLX_IDinst_Mcompar__n0100_inst_cy_263/LOGIC_ZERO ;
  wire \DLX_IDinst_Mcompar__n0100_inst_cy_263/LOGIC_ONE ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1083;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_1009/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1084;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_1008;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_1009/LOGIC_ZERO ;
  wire \DLX_IDinst_Mmux__COND_5_inst_cy_1009/LOGIC_ONE ;
  wire DLX_IDinst_Mcompar__n0105_inst_lut4_40;
  wire \DLX_IDinst_Mcompar__n0105_inst_cy_263/CYMUXG ;
  wire DLX_IDinst_Mcompar__n0105_inst_lut4_41;
  wire DLX_IDinst_Mcompar__n0105_inst_cy_262;
  wire \DLX_IDinst_Mcompar__n0105_inst_cy_263/LOGIC_ZERO ;
  wire \DLX_IDinst_Mcompar__n0105_inst_cy_263/LOGIC_ONE ;
  wire \DLX_IDinst__n0105/LOGIC_ZERO ;
  wire DLX_IDinst_Mcompar__n0105_inst_lut4_42;
  wire \DLX_IDinst__n0105/CYMUXF ;
  wire \DLX_IDinst__n0105/CYINIT ;
  wire DLX_IDinst_Mcompar__n0367_inst_lut4_40;
  wire \DLX_IDinst_Mcompar__n0367_inst_cy_263/CYMUXG ;
  wire DLX_IDinst_Mcompar__n0367_inst_lut4_41;
  wire DLX_IDinst_Mcompar__n0367_inst_cy_262;
  wire \DLX_IDinst_Mcompar__n0367_inst_cy_263/LOGIC_ZERO ;
  wire \DLX_IDinst_Mcompar__n0367_inst_cy_263/LOGIC_ONE ;
  wire \DLX_IDinst__n0367/LOGIC_ZERO ;
  wire DLX_IDinst_Mcompar__n0367_inst_lut4_42;
  wire \DLX_IDinst__n0367/CYMUXF ;
  wire \DLX_IDinst__n0367/CYINIT ;
  wire \DLX_IDinst_RegFile_10_20/GROM ;
  wire \DLX_IDinst_RegFile_10_21/GROM ;
  wire \DLX_IDinst_RegFile_10_22/GROM ;
  wire \DLX_IDinst_RegFile_10_23/GROM ;
  wire \DLX_IDinst_RegFile_10_31/GROM ;
  wire \DLX_IDinst_RegFile_10_24/GROM ;
  wire \DLX_IDinst_RegFile_10_16/GROM ;
  wire \DLX_IDinst_RegFile_10_25/GROM ;
  wire \DLX_IDinst_RegFile_10_17/GROM ;
  wire \DLX_IDinst_RegFile_10_26/GROM ;
  wire \DLX_IDinst_RegFile_10_18/GROM ;
  wire \DLX_IDinst_RegFile_10_27/GROM ;
  wire \DLX_IDinst_RegFile_10_19/GROM ;
  wire \DLX_IDinst_RegFile_10_28/GROM ;
  wire \DLX_IDinst_RegFile_10_29/GROM ;
  wire DLX_IDinst__n0124;
  wire DLX_IDinst__n0125;
  wire \DLX_EXinst_ALU_result_10_1/GROM ;
  wire \DLX_EXinst_ALU_result_11_1/GROM ;
  wire \DLX_EXinst_ALU_result_12_1/GROM ;
  wire \DLX_EXinst_ALU_result_13_1/GROM ;
  wire \DLX_EXinst_ALU_result_14_1/GROM ;
  wire \DLX_IDinst_current_IR<0>/GROM ;
  wire \DLX_IDinst_current_IR<1>/GROM ;
  wire \DLX_IDinst_current_IR<2>/GROM ;
  wire \DLX_IDinst_current_IR<3>/GROM ;
  wire \DLX_IDinst_current_IR<4>/GROM ;
  wire \DLX_IDinst_current_IR<5>/GROM ;
  wire \DLX_IDinst_current_IR<6>/GROM ;
  wire \DLX_IDinst_current_IR<7>/GROM ;
  wire \DLX_IDinst_current_IR<8>/GROM ;
  wire \DLX_IDinst_current_IR<9>/GROM ;
  wire \DLX_EXinst_ALU_result<8>/GROM ;
  wire DLX_IDinst__n0155;
  wire DLX_IDinst__n0119;
  wire DLX_IDinst__n0126;
  wire DLX_IDinst__n0127;
  wire DLX_IDinst__n0128;
  wire \DLX_IDinst_Imm<1>/GROM ;
  wire \DLX_IDinst_Imm<2>/GROM ;
  wire \DLX_IDinst_Imm<3>/GROM ;
  wire DLX_IDinst__n0140;
  wire \DLX_IDinst_CLI/GROM ;
  wire \DLX_IDinst_current_IR<10>/GROM ;
  wire \DLX_IDinst_current_IR<11>/GROM ;
  wire \DLX_IDinst_current_IR<20>/FROM ;
  wire \DLX_IDinst_current_IR<20>/GROM ;
  wire \DLX_IDinst_current_IR<12>/GROM ;
  wire \DLX_IDinst_current_IR<13>/GROM ;
  wire \DLX_IDinst_current_IR<30>/FROM ;
  wire \DLX_IDinst_current_IR<30>/GROM ;
  wire \DLX_IDinst_current_IR<14>/GROM ;
  wire \DLX_IDinst_current_IR<22>/FROM ;
  wire \DLX_IDinst_current_IR<22>/GROM ;
  wire \DLX_IDinst_current_IR<23>/FROM ;
  wire \DLX_IDinst_current_IR<23>/GROM ;
  wire \DLX_IDinst_current_IR<31>/FROM ;
  wire \DLX_IDinst_current_IR<31>/GROM ;
  wire \DLX_IDinst_current_IR<15>/GROM ;
  wire \DLX_IDinst_current_IR<24>/FROM ;
  wire \DLX_IDinst_current_IR<24>/GROM ;
  wire \DLX_IDinst_current_IR<25>/FROM ;
  wire \DLX_IDinst_current_IR<25>/GROM ;
  wire \DLX_IDinst_current_IR<17>/FROM ;
  wire \DLX_IDinst_current_IR<17>/GROM ;
  wire \DLX_IDinst_current_IR<26>/FROM ;
  wire \DLX_IDinst_current_IR<26>/GROM ;
  wire \DLX_IDinst_current_IR<18>/FROM ;
  wire \DLX_IDinst_current_IR<18>/GROM ;
  wire \DLX_IDinst_current_IR<27>/FROM ;
  wire \DLX_IDinst_current_IR<27>/GROM ;
  wire \DLX_IDinst_current_IR<19>/FROM ;
  wire \DLX_IDinst_current_IR<19>/GROM ;
  wire \DLX_IDinst_current_IR<28>/FROM ;
  wire \DLX_IDinst_current_IR<28>/GROM ;
  wire \DLX_IDinst_current_IR<29>/FROM ;
  wire \DLX_IDinst_current_IR<29>/GROM ;
  wire DLX_IDinst__n0120;
  wire DLX_IDinst__n0123;
  wire DLX_IDinst__n0121;
  wire DLX_IDinst__n0122;
  wire \DLX_IDinst_reg_out_B<2>/GROM ;
  wire \DLX_IDinst_reg_out_B<3>/GROM ;
  wire N162904;
  wire N162907;
  wire N162910;
  wire N162934;
  wire N162913;
  wire N162937;
  wire N162916;
  wire N162940;
  wire N162871;
  wire N162919;
  wire N162943;
  wire N162922;
  wire N162946;
  wire N162925;
  wire N162949;
  wire N162928;
  wire N162952;
  wire N162931;
  wire N162955;
  wire N162958;
  wire N162961;
  wire N162874;
  wire N162877;
  wire N162880;
  wire N162883;
  wire N162886;
  wire N162889;
  wire N162892;
  wire N162895;
  wire N162898;
  wire N162901;
  wire \DLX_EXinst_reg_dst_out<0>/GROM ;
  wire \DLX_EXinst_reg_dst_out<1>/GROM ;
  wire \DLX_EXinst_reg_dst_out<2>/GROM ;
  wire \DLX_EXinst_reg_dst_out<3>/GROM ;
  wire \DLX_EXinst_reg_dst_out<4>/LOGIC_ZERO ;
  wire DLX_IDinst_Mcompar__n0100_inst_lut4_42;
  wire \DLX_EXinst_reg_dst_out<4>/CYMUXF ;
  wire \DLX_EXinst_reg_dst_out<4>/CYINIT ;
  wire \DLX_EXinst_reg_dst_out<4>/GROM ;
  wire \DLX_EXinst_reg_out_B_EX<6>/FROM ;
  wire \DLX_EXinst_reg_out_B_EX<6>/GROM ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_225;
  wire \DLX_IDinst_RegFile_12_10/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_226;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_166;
  wire \DLX_IDinst_RegFile_12_10/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_12_10/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_229;
  wire \DLX_IDinst_RegFile_20_10/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_230;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_170;
  wire \DLX_IDinst_RegFile_20_10/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_20_10/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_241;
  wire \DLX_IDinst_RegFile_12_11/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_242;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_182;
  wire \DLX_IDinst_RegFile_12_11/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_12_11/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_245;
  wire \DLX_IDinst_RegFile_20_11/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_246;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_186;
  wire \DLX_IDinst_RegFile_20_11/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_20_11/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_385;
  wire \DLX_IDinst_RegFile_12_20/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_386;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_326;
  wire \DLX_IDinst_RegFile_12_20/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_12_20/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_257;
  wire \DLX_IDinst_RegFile_12_12/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_258;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_198;
  wire \DLX_IDinst_RegFile_12_12/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_12_12/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_389;
  wire \DLX_IDinst_RegFile_20_20/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_390;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_330;
  wire \DLX_IDinst_RegFile_20_20/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_20_20/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_261;
  wire \DLX_IDinst_RegFile_20_12/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_262;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_202;
  wire \DLX_IDinst_RegFile_20_12/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_20_12/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_401;
  wire \DLX_IDinst_RegFile_12_21/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_402;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_342;
  wire \DLX_IDinst_RegFile_12_21/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_12_21/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_273;
  wire \DLX_IDinst_RegFile_12_13/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_274;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_214;
  wire \DLX_IDinst_RegFile_12_13/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_12_13/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_405;
  wire \DLX_IDinst_RegFile_20_21/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_406;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_346;
  wire \DLX_IDinst_RegFile_20_21/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_20_21/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_277;
  wire \DLX_IDinst_RegFile_20_13/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_278;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_218;
  wire \DLX_IDinst_RegFile_20_13/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_20_13/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1073;
  wire \DLX_IDinst_RegFile_12_30/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1074;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_998;
  wire \DLX_IDinst_RegFile_12_30/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_12_30/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_417;
  wire \DLX_IDinst_RegFile_12_22/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_418;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_358;
  wire \DLX_IDinst_RegFile_12_22/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_12_22/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_289;
  wire \DLX_IDinst_RegFile_12_14/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_290;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_230;
  wire \DLX_IDinst_RegFile_12_14/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_12_14/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1077;
  wire \DLX_IDinst_RegFile_20_30/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1078;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_1002;
  wire \DLX_IDinst_RegFile_20_30/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_20_30/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_421;
  wire \DLX_IDinst_RegFile_20_22/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_422;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_362;
  wire \DLX_IDinst_RegFile_20_22/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_20_22/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_293;
  wire \DLX_IDinst_RegFile_20_14/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_294;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_234;
  wire \DLX_IDinst_RegFile_20_14/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_20_14/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_433;
  wire \DLX_IDinst_RegFile_12_23/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_434;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_374;
  wire \DLX_IDinst_RegFile_12_23/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_12_23/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_305;
  wire \DLX_IDinst_RegFile_12_15/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_306;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_246;
  wire \DLX_IDinst_RegFile_12_15/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_12_15/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_437;
  wire \DLX_IDinst_RegFile_20_23/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_438;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_378;
  wire \DLX_IDinst_RegFile_20_23/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_20_23/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_309;
  wire \DLX_IDinst_RegFile_20_15/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_310;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_250;
  wire \DLX_IDinst_RegFile_20_15/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_20_15/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1089;
  wire \DLX_IDinst_RegFile_12_31/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1090;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_1014;
  wire \DLX_IDinst_RegFile_12_31/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_12_31/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1093;
  wire \DLX_IDinst_RegFile_20_31/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1094;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_1018;
  wire \DLX_IDinst_RegFile_20_31/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_20_31/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_449;
  wire \DLX_IDinst_RegFile_12_24/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_450;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_390;
  wire \DLX_IDinst_RegFile_12_24/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_12_24/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_321;
  wire \DLX_IDinst_RegFile_12_16/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_322;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_262;
  wire \DLX_IDinst_RegFile_12_16/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_12_16/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_453;
  wire \DLX_IDinst_RegFile_20_24/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_454;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_394;
  wire \DLX_IDinst_RegFile_20_24/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_20_24/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_325;
  wire \DLX_IDinst_RegFile_20_16/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_326;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_266;
  wire \DLX_IDinst_RegFile_20_16/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_20_16/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_465;
  wire \DLX_IDinst_RegFile_12_25/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_466;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_406;
  wire \DLX_IDinst_RegFile_12_25/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_12_25/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_337;
  wire \DLX_IDinst_RegFile_12_17/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_338;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_278;
  wire \DLX_IDinst_RegFile_12_17/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_12_17/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_469;
  wire \DLX_IDinst_RegFile_20_25/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_470;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_410;
  wire \DLX_IDinst_RegFile_20_25/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_20_25/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_341;
  wire \DLX_IDinst_RegFile_20_17/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_342;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_282;
  wire \DLX_IDinst_RegFile_20_17/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_20_17/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_481;
  wire \DLX_IDinst_RegFile_12_26/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_482;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_422;
  wire \DLX_IDinst_RegFile_12_26/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_12_26/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_881;
  wire \DLX_IDinst_RegFile_12_18/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_882;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_806;
  wire \DLX_IDinst_RegFile_12_18/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_12_18/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_753;
  wire \DLX_IDinst_RegFile_13_10/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_754;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_678;
  wire \DLX_IDinst_RegFile_13_10/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_13_10/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_485;
  wire \DLX_IDinst_RegFile_20_26/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_486;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_426;
  wire \DLX_IDinst_RegFile_20_26/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_20_26/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_357;
  wire \DLX_IDinst_RegFile_20_18/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_358;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_298;
  wire \DLX_IDinst_RegFile_20_18/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_20_18/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_757;
  wire \DLX_IDinst_RegFile_21_10/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_758;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_682;
  wire \DLX_IDinst_RegFile_21_10/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_21_10/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1025;
  wire \DLX_IDinst_RegFile_12_27/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1026;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_950;
  wire \DLX_IDinst_RegFile_12_27/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_12_27/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_369;
  wire \DLX_IDinst_RegFile_12_19/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_370;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_310;
  wire \DLX_IDinst_RegFile_12_19/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_12_19/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_769;
  wire \DLX_IDinst_RegFile_13_11/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_770;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_694;
  wire \DLX_IDinst_RegFile_13_11/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_13_11/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1029;
  wire \DLX_IDinst_RegFile_20_27/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1030;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_954;
  wire \DLX_IDinst_RegFile_20_27/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_20_27/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_373;
  wire \DLX_IDinst_RegFile_20_19/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_374;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_314;
  wire \DLX_IDinst_RegFile_20_19/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_20_19/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_773;
  wire \DLX_IDinst_RegFile_21_11/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_774;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_698;
  wire \DLX_IDinst_RegFile_21_11/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_21_11/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1041;
  wire \DLX_IDinst_RegFile_12_28/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1042;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_966;
  wire \DLX_IDinst_RegFile_12_28/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_12_28/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_913;
  wire \DLX_IDinst_RegFile_13_20/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_914;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_838;
  wire \DLX_IDinst_RegFile_13_20/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_13_20/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_785;
  wire \DLX_IDinst_RegFile_13_12/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_786;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_710;
  wire \DLX_IDinst_RegFile_13_12/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_13_12/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1045;
  wire \DLX_IDinst_RegFile_20_28/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1046;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_970;
  wire \DLX_IDinst_RegFile_20_28/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_20_28/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_917;
  wire \DLX_IDinst_RegFile_21_20/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_918;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_842;
  wire \DLX_IDinst_RegFile_21_20/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_21_20/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_789;
  wire \DLX_IDinst_RegFile_21_12/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_790;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_714;
  wire \DLX_IDinst_RegFile_21_12/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_21_12/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1057;
  wire \DLX_IDinst_RegFile_12_29/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1058;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_982;
  wire \DLX_IDinst_RegFile_12_29/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_12_29/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_929;
  wire \DLX_IDinst_RegFile_13_21/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_930;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_854;
  wire \DLX_IDinst_RegFile_13_21/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_13_21/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_801;
  wire \DLX_IDinst_RegFile_13_13/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_802;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_726;
  wire \DLX_IDinst_RegFile_13_13/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_13_13/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1061;
  wire \DLX_IDinst_RegFile_20_29/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1062;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_986;
  wire \DLX_IDinst_RegFile_20_29/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_20_29/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_933;
  wire \DLX_IDinst_RegFile_21_21/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_934;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_858;
  wire \DLX_IDinst_RegFile_21_21/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_21_21/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_805;
  wire \DLX_IDinst_RegFile_21_13/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_806;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_730;
  wire \DLX_IDinst_RegFile_21_13/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_21_13/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_545;
  wire \DLX_IDinst_RegFile_13_30/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_546;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_486;
  wire \DLX_IDinst_RegFile_13_30/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_13_30/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_945;
  wire \DLX_IDinst_RegFile_13_22/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_946;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_870;
  wire \DLX_IDinst_RegFile_13_22/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_13_22/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_817;
  wire \DLX_IDinst_RegFile_13_14/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_818;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_742;
  wire \DLX_IDinst_RegFile_13_14/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_13_14/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_549;
  wire \DLX_IDinst_RegFile_21_30/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_550;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_490;
  wire \DLX_IDinst_RegFile_21_30/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_21_30/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_949;
  wire \DLX_IDinst_RegFile_21_22/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_950;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_874;
  wire \DLX_IDinst_RegFile_21_22/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_21_22/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_821;
  wire \DLX_IDinst_RegFile_21_14/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_822;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_746;
  wire \DLX_IDinst_RegFile_21_14/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_21_14/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_961;
  wire \DLX_IDinst_RegFile_13_23/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_962;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_886;
  wire \DLX_IDinst_RegFile_13_23/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_13_23/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_833;
  wire \DLX_IDinst_RegFile_13_15/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_834;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_758;
  wire \DLX_IDinst_RegFile_13_15/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_13_15/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_965;
  wire \DLX_IDinst_RegFile_21_23/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_966;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_890;
  wire \DLX_IDinst_RegFile_21_23/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_21_23/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_837;
  wire \DLX_IDinst_RegFile_21_15/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_838;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_762;
  wire \DLX_IDinst_RegFile_21_15/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_21_15/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_561;
  wire \DLX_IDinst_RegFile_13_31/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_562;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_502;
  wire \DLX_IDinst_RegFile_13_31/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_13_31/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_565;
  wire \DLX_IDinst_RegFile_21_31/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_566;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_506;
  wire \DLX_IDinst_RegFile_21_31/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_21_31/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_977;
  wire \DLX_IDinst_RegFile_13_24/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_978;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_902;
  wire \DLX_IDinst_RegFile_13_24/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_13_24/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_849;
  wire \DLX_IDinst_RegFile_13_16/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_850;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_774;
  wire \DLX_IDinst_RegFile_13_16/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_13_16/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_981;
  wire \DLX_IDinst_RegFile_21_24/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_982;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_906;
  wire \DLX_IDinst_RegFile_21_24/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_21_24/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_853;
  wire \DLX_IDinst_RegFile_21_16/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_854;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_778;
  wire \DLX_IDinst_RegFile_21_16/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_21_16/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_993;
  wire \DLX_IDinst_RegFile_13_25/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_994;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_918;
  wire \DLX_IDinst_RegFile_13_25/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_13_25/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_865;
  wire \DLX_IDinst_RegFile_13_17/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_866;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_790;
  wire \DLX_IDinst_RegFile_13_17/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_13_17/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_997;
  wire \DLX_IDinst_RegFile_21_25/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_998;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_922;
  wire \DLX_IDinst_RegFile_21_25/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_21_25/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_869;
  wire \DLX_IDinst_RegFile_21_17/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_870;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_794;
  wire \DLX_IDinst_RegFile_21_17/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_21_17/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1009;
  wire \DLX_IDinst_RegFile_13_26/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1010;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_934;
  wire \DLX_IDinst_RegFile_13_26/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_13_26/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1013;
  wire \DLX_IDinst_RegFile_21_26/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_1014;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_938;
  wire \DLX_IDinst_RegFile_21_26/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_21_26/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_885;
  wire \DLX_IDinst_RegFile_21_18/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_886;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_810;
  wire \DLX_IDinst_RegFile_21_18/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_21_18/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_497;
  wire \DLX_IDinst_RegFile_13_27/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_498;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_438;
  wire \DLX_IDinst_RegFile_13_27/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_13_27/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_897;
  wire \DLX_IDinst_RegFile_13_19/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_898;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_822;
  wire \DLX_IDinst_RegFile_13_19/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_13_19/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_501;
  wire \DLX_IDinst_RegFile_21_27/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_502;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_442;
  wire \DLX_IDinst_RegFile_21_27/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_21_27/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_901;
  wire \DLX_IDinst_RegFile_21_19/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_902;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_826;
  wire \DLX_IDinst_RegFile_21_19/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_21_19/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_513;
  wire \DLX_IDinst_RegFile_13_28/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_514;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_454;
  wire \DLX_IDinst_RegFile_13_28/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_13_28/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_517;
  wire \DLX_IDinst_RegFile_21_28/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_518;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_458;
  wire \DLX_IDinst_RegFile_21_28/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_21_28/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_529;
  wire \DLX_IDinst_RegFile_13_29/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_530;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_470;
  wire \DLX_IDinst_RegFile_13_29/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_13_29/CYINIT ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_533;
  wire \DLX_IDinst_RegFile_21_29/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_4_inst_lut4_534;
  wire DLX_IDinst_Mmux__COND_4_inst_cy_474;
  wire \DLX_IDinst_RegFile_21_29/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_21_29/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_755;
  wire \DLX_IDinst_RegFile_16_10/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_756;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_680;
  wire \DLX_IDinst_RegFile_16_10/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_16_10/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_759;
  wire \DLX_IDinst_RegFile_24_10/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_760;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_684;
  wire \DLX_IDinst_RegFile_24_10/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_24_10/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_771;
  wire \DLX_IDinst_RegFile_16_11/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_772;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_696;
  wire \DLX_IDinst_RegFile_16_11/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_16_11/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_775;
  wire \DLX_IDinst_RegFile_24_11/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_776;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_700;
  wire \DLX_IDinst_RegFile_24_11/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_24_11/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_915;
  wire \DLX_IDinst_RegFile_16_20/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_916;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_840;
  wire \DLX_IDinst_RegFile_16_20/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_16_20/CYINIT ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_787;
  wire \DLX_IDinst_RegFile_16_12/CYMUXG ;
  wire DLX_IDinst_Mmux__COND_5_inst_lut4_788;
  wire DLX_IDinst_Mmux__COND_5_inst_cy_712;
  wire \DLX_IDinst_RegFile_16_12/LOGIC_ZERO ;
  wire \DLX_IDinst_RegFile_16_12/CYINIT ;
  wire \CHOICE3150/FROM ;
  wire \CHOICE3150/GROM ;
  wire \DLX_IDinst_Cause_Reg<0>/FFY/RST ;
  wire \DLX_IDinst_Cause_Reg<1>/FFY/RST ;
  wire \DLX_IDinst_Cause_Reg<3>/FFY/RST ;
  wire \DLX_IDinst_Cause_Reg<2>/FFY/RST ;
  wire \DLX_IDinst_Cause_Reg<4>/FFY/RST ;
  wire \DLX_IDinst_Cause_Reg<5>/FFY/RST ;
  wire \DLX_IDinst_Cause_Reg<7>/FFY/RST ;
  wire \DLX_IDinst_Cause_Reg<8>/FFY/RST ;
  wire \DLX_IDinst_Cause_Reg<9>/FFY/RST ;
  wire \DLX_IDinst_Cause_Reg<10>/FFY/RST ;
  wire \DLX_IDinst_Cause_Reg<12>/FFY/RST ;
  wire \DLX_IDinst_Cause_Reg<11>/FFY/RST ;
  wire \DLX_IDinst_Cause_Reg<13>/FFY/RST ;
  wire \DLX_IDinst_Cause_Reg<14>/FFY/RST ;
  wire \DLX_IDinst_Cause_Reg<15>/FFY/RST ;
  wire \DLX_IDinst_Cause_Reg<31>/FFY/RST ;
  wire \DLX_IDinst_Cause_Reg<6>/FFY/RST ;
  wire \clkbuf2/CE ;
  wire \clkbuf3/CE ;
  wire \PWR_GND_0/FROM ;
  wire \PWR_GND_0/GROM ;
  wire GND;
  wire VCC;
  wire \NLW_Mmux__COND_2_inst_mux_f6_0.F51_IA_UNCONNECTED ;
  wire [0 : 0] DM_write_data;
  wire [31 : 8] DLX_IDinst_WB_data_eff;
  wire [25 : 0] DLX_IDinst_jtarget;
  wire [31 : 0] DLX_IDinst__n0623;
  wire [31 : 0] DLX_IDinst__n0620;
  wire [5 : 5] DLX_IDinst_IR_function_field;
  wire [5 : 0] DLX_IDinst_IR_opcode_field;
  wire [31 : 0] DLX_IDinst_reg_out_B;
  wire [31 : 0] DLX_IFinst_IR_latched;
  wire [31 : 0] DLX_IFinst_IR_previous;
  wire [31 : 0] DLX_EXinst_reg_out_B_EX;
  wire [31 : 26] DLX_IDinst_IR_latched;
  wire [5 : 0] DLX_IDinst__n0143;
  wire [31 : 0] DLX_MEMinst_RF_data_in;
  wire [31 : 0] DLX_EXinst_ALU_result;
  wire [31 : 0] DLX_IFinst_NPC;
  wire [31 : 0] DLX_IFinst_PC;
  wire [31 : 0] DLX_IDinst_reg_out_A;
  wire [31 : 0] DLX_IDinst_EPC;
  wire [5 : 0] DLX_EXinst_opcode_of_EX_reg;
  wire [5 : 0] DLX_MEMinst_opcode_of_WB;
  wire [31 : 0] DLX_EXinst__n0013;
  wire [31 : 0] DLX_EXinst__n0012;
  wire [9 : 0] vga_top_vga1_vcounter;
  wire [15 : 0] vga_top_vga1_hcounter;
  wire [4 : 0] DLX_MEMinst_reg_dst_out;
  wire [1 : 1] DLX_IDinst__n0629;
  wire [31 : 0] DLX_IFinst_IR_curr;
  wire [31 : 0] DLX_IDinst_branch_address;
  wire [31 : 0] DLX_IFinst__n0001;
  wire [31 : 3] DLX_IFinst__n0015;
  wire [23 : 0] IR;
  wire [31 : 0] DLX_IDinst_current_IR;
  wire [1 : 0] DLX_IDinst_counter;
  wire [31 : 0] DLX_IDinst__n0157;
  wire [2 : 0] vga_top_vga1_helpcounter;
  wire [4 : 0] vram_out_cpu;
  wire [37 : 33] Mshift__n0000_Sh;
  wire [31 : 0] RAM_read_data;
  wire [31 : 0] DM_read_data;
  wire [4 : 0] DLX_EXinst_reg_dst_out;
  wire [4 : 0] DLX_IDinst_rt_addr;
  wire [4 : 0] DLX_IDinst__n0018;
  wire [4 : 0] DLX_IDinst_rd_addr;
  wire [5 : 5] DLX_IDinst__n0025;
  wire [47 : 40] DLX_IDinst__n0618;
  wire [14 : 6] vga_address;
  wire [8 : 0] vga_top_vga1_gridhcounter;
  wire [4 : 0] vram_out_vga;
  wire [8 : 0] vga_top_vga1_gridvcounter;
  wire [31 : 1] DLX_IDinst__n0158;
  wire [4 : 0] DLX_reg_dst_of_EX;
  wire [31 : 0] DLX_IDinst__n0147;
  wire [5 : 0] DLX_IDinst__n0142;
  wire [4 : 0] DLX_IDinst__n0136;
  wire [2 : 1] vga_top_vga1_helpcounter__n0000;
  wire [31 : 0] DLX_MEMinst__n0000;
  wire [31 : 8] DLX_EXinst__n0008;
  wire [4 : 0] DLX_IDinst__n0135;
  wire [31 : 0] DLX_IFinst__n0003;
  wire [9 : 1] vga_top_vga1_vcounter__n0000;
  wire [8 : 1] vga_top_vga1_gridvcounter__n0000;
  wire [8 : 1] vga_top_vga1_gridhcounter__n0000;
  wire [15 : 1] vga_top_vga1_hcounter__n0000;
  wire [1 : 1] DLX_IDinst__n0145;
  assign
    DM_write_data_0 = DM_write_data[0];
  initial $sdf_annotate("DLX_top_timesim.sdf");
  defparam DLX_IDinst_RegFile_25_28_0.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_25_28_0 (
    .I(DLX_IDinst_WB_data_eff[28]),
    .CE(DLX_IDinst__n0600),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_25_28)
  );
  X_ZERO \DLX_IDinst_RegFile_25_28/LOGIC_ZERO_1  (
    .O(\DLX_IDinst_RegFile_25_28/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_972_2 (
    .IA(\DLX_IDinst_RegFile_25_28/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_25_28/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1047),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_972)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10471.INIT = 16'hDDF5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10471 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_583),
    .ADR1(DLX_IDinst_RegFile_25_28),
    .ADR2(DLX_IDinst_RegFile_24_28),
    .ADR3(DLX_IDinst_jtarget[21]),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1047)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10481.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10481 (
    .ADR0(DLX_IDinst_RegFile_27_28),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_584),
    .ADR2(DLX_IDinst_RegFile_26_28),
    .ADR3(DLX_IDinst_jtarget[21]),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1048)
  );
  X_BUF \DLX_IDinst_RegFile_25_28/COUTUSED  (
    .I(\DLX_IDinst_RegFile_25_28/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_973)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_973_3 (
    .IA(\DLX_IDinst_RegFile_25_28/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_972),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1048),
    .O(\DLX_IDinst_RegFile_25_28/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_25_28/CYINIT_4  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_971),
    .O(\DLX_IDinst_RegFile_25_28/CYINIT )
  );
  defparam DLX_IDinst_RegFile_26_20_5.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_26_20_5 (
    .I(DLX_IDinst_WB_data_eff[20]),
    .CE(DLX_IDinst__n0602),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_26_20)
  );
  X_ZERO \DLX_IDinst_RegFile_26_20/LOGIC_ZERO_6  (
    .O(\DLX_IDinst_RegFile_26_20/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_332_7 (
    .IA(\DLX_IDinst_RegFile_26_20/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_26_20/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_391),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_332)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3911.INIT = 16'hAFCF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3911 (
    .ADR0(DLX_IDinst_RegFile_25_20),
    .ADR1(DLX_IDinst_RegFile_24_20),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_55),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_391)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3921.INIT = 16'hDDF5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3921 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_56),
    .ADR1(DLX_IDinst_RegFile_27_20),
    .ADR2(DLX_IDinst_RegFile_26_20),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_392)
  );
  X_BUF \DLX_IDinst_RegFile_26_20/COUTUSED  (
    .I(\DLX_IDinst_RegFile_26_20/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_333)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_333_8 (
    .IA(\DLX_IDinst_RegFile_26_20/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_332),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_392),
    .O(\DLX_IDinst_RegFile_26_20/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_26_20/CYINIT_9  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_331),
    .O(\DLX_IDinst_RegFile_26_20/CYINIT )
  );
  defparam DLX_IDinst_RegFile_26_12_10.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_26_12_10 (
    .I(DLX_IDinst_WB_data_eff[12]),
    .CE(DLX_IDinst__n0602),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_26_12)
  );
  X_ZERO \DLX_IDinst_RegFile_26_12/LOGIC_ZERO_11  (
    .O(\DLX_IDinst_RegFile_26_12/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_204_12 (
    .IA(\DLX_IDinst_RegFile_26_12/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_26_12/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_263),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_204)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2631.INIT = 16'hBFB3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2631 (
    .ADR0(DLX_IDinst_RegFile_25_12),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_55),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR3(DLX_IDinst_RegFile_24_12),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_263)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2641.INIT = 16'hDFD5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2641 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_56),
    .ADR1(DLX_IDinst_RegFile_27_12),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR3(DLX_IDinst_RegFile_26_12),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_264)
  );
  X_BUF \DLX_IDinst_RegFile_26_12/COUTUSED  (
    .I(\DLX_IDinst_RegFile_26_12/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_205)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_205_13 (
    .IA(\DLX_IDinst_RegFile_26_12/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_204),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_264),
    .O(\DLX_IDinst_RegFile_26_12/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_26_12/CYINIT_14  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_203),
    .O(\DLX_IDinst_RegFile_26_12/CYINIT )
  );
  defparam DLX_IDinst_RegFile_17_29_15.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_17_29_15 (
    .I(DLX_IDinst_WB_data_eff[29]),
    .CE(DLX_IDinst__n0584),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_17_29)
  );
  X_ZERO \DLX_IDinst_RegFile_17_29/LOGIC_ZERO_16  (
    .O(\DLX_IDinst_RegFile_17_29/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_984_17 (
    .IA(\DLX_IDinst_RegFile_17_29/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_17_29/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1059),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_984)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10591.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10591 (
    .ADR0(DLX_IDinst_RegFile_16_29),
    .ADR1(DLX_IDinst_RegFile_17_29),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_579),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1059)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10601.INIT = 16'hFD5D;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10601 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_580),
    .ADR1(DLX_IDinst_RegFile_18_29),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR3(DLX_IDinst_RegFile_19_29),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1060)
  );
  X_BUF \DLX_IDinst_RegFile_17_29/COUTUSED  (
    .I(\DLX_IDinst_RegFile_17_29/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_985)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_985_18 (
    .IA(\DLX_IDinst_RegFile_17_29/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_984),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1060),
    .O(\DLX_IDinst_RegFile_17_29/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_17_29/CYINIT_19  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_983),
    .O(\DLX_IDinst_RegFile_17_29/CYINIT )
  );
  defparam DLX_IDinst_RegFile_18_21_20.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_18_21_20 (
    .I(DLX_IDinst_WB_data_eff[21]),
    .CE(DLX_IDinst__n0586),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_18_21)
  );
  X_ZERO \DLX_IDinst_RegFile_18_21/LOGIC_ZERO_21  (
    .O(\DLX_IDinst_RegFile_18_21/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_344_22 (
    .IA(\DLX_IDinst_RegFile_18_21/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_18_21/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_403),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_344)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4031.INIT = 16'hDDF5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4031 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_51),
    .ADR1(DLX_IDinst_RegFile_17_21),
    .ADR2(DLX_IDinst_RegFile_16_21),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_403)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4041.INIT = 16'hCFAF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4041 (
    .ADR0(DLX_IDinst_RegFile_18_21),
    .ADR1(DLX_IDinst_RegFile_19_21),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_52),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_404)
  );
  X_BUF \DLX_IDinst_RegFile_18_21/COUTUSED  (
    .I(\DLX_IDinst_RegFile_18_21/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_345)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_345_23 (
    .IA(\DLX_IDinst_RegFile_18_21/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_344),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_404),
    .O(\DLX_IDinst_RegFile_18_21/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_18_21/CYINIT_24  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_343),
    .O(\DLX_IDinst_RegFile_18_21/CYINIT )
  );
  defparam DLX_IDinst_RegFile_18_13_25.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_18_13_25 (
    .I(DLX_IDinst_WB_data_eff[13]),
    .CE(DLX_IDinst__n0586),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_18_13)
  );
  X_ZERO \DLX_IDinst_RegFile_18_13/LOGIC_ZERO_26  (
    .O(\DLX_IDinst_RegFile_18_13/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_216_27 (
    .IA(\DLX_IDinst_RegFile_18_13/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_18_13/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_275),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_216)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2751.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2751 (
    .ADR0(DLX_IDinst_RegFile_16_13),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_51),
    .ADR2(DLX_IDinst_RegFile_17_13),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_275)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2761.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2761 (
    .ADR0(DLX_IDinst_RegFile_18_13),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_52),
    .ADR2(DLX_IDinst_RegFile_19_13),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_276)
  );
  X_BUF \DLX_IDinst_RegFile_18_13/COUTUSED  (
    .I(\DLX_IDinst_RegFile_18_13/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_217)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_217_28 (
    .IA(\DLX_IDinst_RegFile_18_13/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_216),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_276),
    .O(\DLX_IDinst_RegFile_18_13/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_18_13/CYINIT_29  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_215),
    .O(\DLX_IDinst_RegFile_18_13/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_25_29/LOGIC_ZERO_30  (
    .O(\DLX_IDinst_RegFile_25_29/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_988_31 (
    .IA(\DLX_IDinst_RegFile_25_29/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_25_29/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1063),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_988)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10631.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10631 (
    .ADR0(DLX_IDinst_RegFile_24_29),
    .ADR1(DLX_IDinst_RegFile_25_29),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_583),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1063)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10641.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10641 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR1(DLX_IDinst_RegFile_26_29),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_584),
    .ADR3(DLX_IDinst_RegFile_27_29),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1064)
  );
  X_BUF \DLX_IDinst_RegFile_25_29/COUTUSED  (
    .I(\DLX_IDinst_RegFile_25_29/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_989)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_989_32 (
    .IA(\DLX_IDinst_RegFile_25_29/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_988),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1064),
    .O(\DLX_IDinst_RegFile_25_29/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_25_29/CYINIT_33  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_987),
    .O(\DLX_IDinst_RegFile_25_29/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_26_21/LOGIC_ZERO_34  (
    .O(\DLX_IDinst_RegFile_26_21/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_348_35 (
    .IA(\DLX_IDinst_RegFile_26_21/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_26_21/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_407),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_348)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4071.INIT = 16'hF7B3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4071 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_55),
    .ADR2(DLX_IDinst_RegFile_25_21),
    .ADR3(DLX_IDinst_RegFile_24_21),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_407)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4081.INIT = 16'hDFD5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4081 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_56),
    .ADR1(DLX_IDinst_RegFile_27_21),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR3(DLX_IDinst_RegFile_26_21),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_408)
  );
  X_BUF \DLX_IDinst_RegFile_26_21/COUTUSED  (
    .I(\DLX_IDinst_RegFile_26_21/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_349)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_349_36 (
    .IA(\DLX_IDinst_RegFile_26_21/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_348),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_408),
    .O(\DLX_IDinst_RegFile_26_21/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_26_21/CYINIT_37  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_347),
    .O(\DLX_IDinst_RegFile_26_21/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_26_13/LOGIC_ZERO_38  (
    .O(\DLX_IDinst_RegFile_26_13/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_220_39 (
    .IA(\DLX_IDinst_RegFile_26_13/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_26_13/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_279),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_220)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2791.INIT = 16'hFB3B;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2791 (
    .ADR0(DLX_IDinst_RegFile_24_13),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_55),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR3(DLX_IDinst_RegFile_25_13),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_279)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2801.INIT = 16'hFB73;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2801 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_56),
    .ADR2(DLX_IDinst_RegFile_26_13),
    .ADR3(DLX_IDinst_RegFile_27_13),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_280)
  );
  X_BUF \DLX_IDinst_RegFile_26_13/COUTUSED  (
    .I(\DLX_IDinst_RegFile_26_13/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_221)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_221_40 (
    .IA(\DLX_IDinst_RegFile_26_13/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_220),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_280),
    .O(\DLX_IDinst_RegFile_26_13/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_26_13/CYINIT_41  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_219),
    .O(\DLX_IDinst_RegFile_26_13/CYINIT )
  );
  defparam vga_top_vga1__n000962.INIT = 16'hFFF0;
  X_LUT4 vga_top_vga1__n000962 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(vga_top_vga1__n0029),
    .ADR3(vga_top_vga1__n0030),
    .O(\CHOICE3470/GROM )
  );
  X_BUF \CHOICE3470/YUSED  (
    .I(\CHOICE3470/GROM ),
    .O(CHOICE3470)
  );
  X_ZERO \DLX_IDinst_RegFile_18_30/LOGIC_ZERO_42  (
    .O(\DLX_IDinst_RegFile_18_30/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_1000_43 (
    .IA(\DLX_IDinst_RegFile_18_30/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_18_30/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1075),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_1000)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10751.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10751 (
    .ADR0(DLX_IDinst_RegFile_16_30),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_579),
    .ADR2(DLX_IDinst_RegFile_17_30),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1075)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10761.INIT = 16'hACFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10761 (
    .ADR0(DLX_IDinst_RegFile_19_30),
    .ADR1(DLX_IDinst_RegFile_18_30),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_580),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1076)
  );
  X_BUF \DLX_IDinst_RegFile_18_30/COUTUSED  (
    .I(\DLX_IDinst_RegFile_18_30/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_1001)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_1001_44 (
    .IA(\DLX_IDinst_RegFile_18_30/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_1000),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1076),
    .O(\DLX_IDinst_RegFile_18_30/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_18_30/CYINIT_45  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_999),
    .O(\DLX_IDinst_RegFile_18_30/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_18_22/LOGIC_ZERO_46  (
    .O(\DLX_IDinst_RegFile_18_22/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_360_47 (
    .IA(\DLX_IDinst_RegFile_18_22/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_18_22/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_419),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_360)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4191.INIT = 16'hE4FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4191 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR1(DLX_IDinst_RegFile_16_22),
    .ADR2(DLX_IDinst_RegFile_17_22),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_51),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_419)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4201.INIT = 16'hD8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4201 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR1(DLX_IDinst_RegFile_19_22),
    .ADR2(DLX_IDinst_RegFile_18_22),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_52),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_420)
  );
  X_BUF \DLX_IDinst_RegFile_18_22/COUTUSED  (
    .I(\DLX_IDinst_RegFile_18_22/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_361)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_361_48 (
    .IA(\DLX_IDinst_RegFile_18_22/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_360),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_420),
    .O(\DLX_IDinst_RegFile_18_22/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_18_22/CYINIT_49  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_359),
    .O(\DLX_IDinst_RegFile_18_22/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_18_14/LOGIC_ZERO_50  (
    .O(\DLX_IDinst_RegFile_18_14/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_232_51 (
    .IA(\DLX_IDinst_RegFile_18_14/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_18_14/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_291),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_232)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2911.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2911 (
    .ADR0(DLX_IDinst_RegFile_16_14),
    .ADR1(DLX_IDinst_RegFile_17_14),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_51),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_291)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2921.INIT = 16'hFD5D;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2921 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_52),
    .ADR1(DLX_IDinst_RegFile_18_14),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR3(DLX_IDinst_RegFile_19_14),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_292)
  );
  X_BUF \DLX_IDinst_RegFile_18_14/COUTUSED  (
    .I(\DLX_IDinst_RegFile_18_14/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_233)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_233_52 (
    .IA(\DLX_IDinst_RegFile_18_14/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_232),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_292),
    .O(\DLX_IDinst_RegFile_18_14/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_18_14/CYINIT_53  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_231),
    .O(\DLX_IDinst_RegFile_18_14/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_26_30/LOGIC_ZERO_54  (
    .O(\DLX_IDinst_RegFile_26_30/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_1004_55 (
    .IA(\DLX_IDinst_RegFile_26_30/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_26_30/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1079),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_1004)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10791.INIT = 16'hFB3B;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10791 (
    .ADR0(DLX_IDinst_RegFile_24_30),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_583),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR3(DLX_IDinst_RegFile_25_30),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1079)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10801.INIT = 16'hBFB3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10801 (
    .ADR0(DLX_IDinst_RegFile_27_30),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_584),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR3(DLX_IDinst_RegFile_26_30),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1080)
  );
  X_BUF \DLX_IDinst_RegFile_26_30/COUTUSED  (
    .I(\DLX_IDinst_RegFile_26_30/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_1005)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_1005_56 (
    .IA(\DLX_IDinst_RegFile_26_30/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_1004),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1080),
    .O(\DLX_IDinst_RegFile_26_30/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_26_30/CYINIT_57  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_1003),
    .O(\DLX_IDinst_RegFile_26_30/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_26_22/LOGIC_ZERO_58  (
    .O(\DLX_IDinst_RegFile_26_22/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_364_59 (
    .IA(\DLX_IDinst_RegFile_26_22/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_26_22/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_423),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_364)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4231.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4231 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR1(DLX_IDinst_RegFile_24_22),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_55),
    .ADR3(DLX_IDinst_RegFile_25_22),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_423)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4241.INIT = 16'hF7B3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4241 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_56),
    .ADR2(DLX_IDinst_RegFile_27_22),
    .ADR3(DLX_IDinst_RegFile_26_22),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_424)
  );
  X_BUF \DLX_IDinst_RegFile_26_22/COUTUSED  (
    .I(\DLX_IDinst_RegFile_26_22/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_365)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_365_60 (
    .IA(\DLX_IDinst_RegFile_26_22/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_364),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_424),
    .O(\DLX_IDinst_RegFile_26_22/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_26_22/CYINIT_61  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_363),
    .O(\DLX_IDinst_RegFile_26_22/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_26_14/LOGIC_ZERO_62  (
    .O(\DLX_IDinst_RegFile_26_14/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_236_63 (
    .IA(\DLX_IDinst_RegFile_26_14/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_26_14/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_295),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_236)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2951.INIT = 16'hACFF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2951 (
    .ADR0(DLX_IDinst_RegFile_25_14),
    .ADR1(DLX_IDinst_RegFile_24_14),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_55),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_295)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2961.INIT = 16'hE2FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2961 (
    .ADR0(DLX_IDinst_RegFile_26_14),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR2(DLX_IDinst_RegFile_27_14),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_56),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_296)
  );
  X_BUF \DLX_IDinst_RegFile_26_14/COUTUSED  (
    .I(\DLX_IDinst_RegFile_26_14/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_237)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_237_64 (
    .IA(\DLX_IDinst_RegFile_26_14/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_236),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_296),
    .O(\DLX_IDinst_RegFile_26_14/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_26_14/CYINIT_65  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_235),
    .O(\DLX_IDinst_RegFile_26_14/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_18_23/LOGIC_ZERO_66  (
    .O(\DLX_IDinst_RegFile_18_23/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_376_67 (
    .IA(\DLX_IDinst_RegFile_18_23/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_18_23/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_435),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_376)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4351.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4351 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_51),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR2(DLX_IDinst_RegFile_16_23),
    .ADR3(DLX_IDinst_RegFile_17_23),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_435)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4361.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4361 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR1(DLX_IDinst_RegFile_18_23),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_52),
    .ADR3(DLX_IDinst_RegFile_19_23),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_436)
  );
  X_BUF \DLX_IDinst_RegFile_18_23/COUTUSED  (
    .I(\DLX_IDinst_RegFile_18_23/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_377)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_377_68 (
    .IA(\DLX_IDinst_RegFile_18_23/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_376),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_436),
    .O(\DLX_IDinst_RegFile_18_23/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_18_23/CYINIT_69  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_375),
    .O(\DLX_IDinst_RegFile_18_23/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_18_15/LOGIC_ZERO_70  (
    .O(\DLX_IDinst_RegFile_18_15/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_248_71 (
    .IA(\DLX_IDinst_RegFile_18_15/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_18_15/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_307),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_248)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3071.INIT = 16'hFD5D;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3071 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_51),
    .ADR1(DLX_IDinst_RegFile_16_15),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR3(DLX_IDinst_RegFile_17_15),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_307)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3081.INIT = 16'hDFD5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3081 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_52),
    .ADR1(DLX_IDinst_RegFile_19_15),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR3(DLX_IDinst_RegFile_18_15),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_308)
  );
  X_BUF \DLX_IDinst_RegFile_18_15/COUTUSED  (
    .I(\DLX_IDinst_RegFile_18_15/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_249)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_249_72 (
    .IA(\DLX_IDinst_RegFile_18_15/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_248),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_308),
    .O(\DLX_IDinst_RegFile_18_15/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_18_15/CYINIT_73  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_247),
    .O(\DLX_IDinst_RegFile_18_15/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_26_23/LOGIC_ZERO_74  (
    .O(\DLX_IDinst_RegFile_26_23/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_892_75 (
    .IA(\DLX_IDinst_RegFile_26_23/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_26_23/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_967),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_892)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9671.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9671 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR1(DLX_IDinst_RegFile_24_23),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_583),
    .ADR3(DLX_IDinst_RegFile_25_23),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_967)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9681.INIT = 16'hFD5D;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9681 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_584),
    .ADR1(DLX_IDinst_RegFile_26_23),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR3(DLX_IDinst_RegFile_27_23),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_968)
  );
  X_BUF \DLX_IDinst_RegFile_26_23/COUTUSED  (
    .I(\DLX_IDinst_RegFile_26_23/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_893)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_893_76 (
    .IA(\DLX_IDinst_RegFile_26_23/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_892),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_968),
    .O(\DLX_IDinst_RegFile_26_23/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_26_23/CYINIT_77  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_891),
    .O(\DLX_IDinst_RegFile_26_23/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_26_15/LOGIC_ZERO_78  (
    .O(\DLX_IDinst_RegFile_26_15/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_252_79 (
    .IA(\DLX_IDinst_RegFile_26_15/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_26_15/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_311),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_252)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3111.INIT = 16'hB8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3111 (
    .ADR0(DLX_IDinst_RegFile_25_15),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR2(DLX_IDinst_RegFile_24_15),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_55),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_311)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3121.INIT = 16'hB8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3121 (
    .ADR0(DLX_IDinst_RegFile_27_15),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR2(DLX_IDinst_RegFile_26_15),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_56),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_312)
  );
  X_BUF \DLX_IDinst_RegFile_26_15/COUTUSED  (
    .I(\DLX_IDinst_RegFile_26_15/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_253)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_253_80 (
    .IA(\DLX_IDinst_RegFile_26_15/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_252),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_312),
    .O(\DLX_IDinst_RegFile_26_15/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_26_15/CYINIT_81  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_251),
    .O(\DLX_IDinst_RegFile_26_15/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_18_31/LOGIC_ZERO_82  (
    .O(\DLX_IDinst_RegFile_18_31/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_1016_83 (
    .IA(\DLX_IDinst_RegFile_18_31/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_18_31/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1091),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_1016)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10911.INIT = 16'hAFCF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10911 (
    .ADR0(DLX_IDinst_RegFile_17_31),
    .ADR1(DLX_IDinst_RegFile_16_31),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_579),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1091)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10921.INIT = 16'hBFB3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10921 (
    .ADR0(DLX_IDinst_RegFile_19_31),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_580),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR3(DLX_IDinst_RegFile_18_31),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1092)
  );
  X_BUF \DLX_IDinst_RegFile_18_31/COUTUSED  (
    .I(\DLX_IDinst_RegFile_18_31/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_1017)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_1017_84 (
    .IA(\DLX_IDinst_RegFile_18_31/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_1016),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1092),
    .O(\DLX_IDinst_RegFile_18_31/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_18_31/CYINIT_85  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_1015),
    .O(\DLX_IDinst_RegFile_18_31/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_26_31/LOGIC_ZERO_86  (
    .O(\DLX_IDinst_RegFile_26_31/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_1020_87 (
    .IA(\DLX_IDinst_RegFile_26_31/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_26_31/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1095),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_1020)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10951.INIT = 16'hAFCF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10951 (
    .ADR0(DLX_IDinst_RegFile_25_31),
    .ADR1(DLX_IDinst_RegFile_24_31),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_583),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1095)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10961.INIT = 16'hDDF5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10961 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_584),
    .ADR1(DLX_IDinst_RegFile_27_31),
    .ADR2(DLX_IDinst_RegFile_26_31),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1096)
  );
  X_BUF \DLX_IDinst_RegFile_26_31/COUTUSED  (
    .I(\DLX_IDinst_RegFile_26_31/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_1021)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_1021_88 (
    .IA(\DLX_IDinst_RegFile_26_31/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_1020),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1096),
    .O(\DLX_IDinst_RegFile_26_31/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_26_31/CYINIT_89  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_1019),
    .O(\DLX_IDinst_RegFile_26_31/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_18_24/LOGIC_ZERO_90  (
    .O(\DLX_IDinst_RegFile_18_24/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_392_91 (
    .IA(\DLX_IDinst_RegFile_18_24/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_18_24/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_451),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_392)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4511.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4511 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_51),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR2(DLX_IDinst_RegFile_16_24),
    .ADR3(DLX_IDinst_RegFile_17_24),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_451)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4521.INIT = 16'hB8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4521 (
    .ADR0(DLX_IDinst_RegFile_19_24),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR2(DLX_IDinst_RegFile_18_24),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_52),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_452)
  );
  X_BUF \DLX_IDinst_RegFile_18_24/COUTUSED  (
    .I(\DLX_IDinst_RegFile_18_24/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_393)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_393_92 (
    .IA(\DLX_IDinst_RegFile_18_24/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_392),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_452),
    .O(\DLX_IDinst_RegFile_18_24/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_18_24/CYINIT_93  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_391),
    .O(\DLX_IDinst_RegFile_18_24/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_18_16/LOGIC_ZERO_94  (
    .O(\DLX_IDinst_RegFile_18_16/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_264_95 (
    .IA(\DLX_IDinst_RegFile_18_16/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_18_16/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_323),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_264)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3231.INIT = 16'hDF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3231 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR1(DLX_IDinst_RegFile_17_16),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_51),
    .ADR3(DLX_IDinst_RegFile_16_16),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_323)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3241.INIT = 16'hBFB3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3241 (
    .ADR0(DLX_IDinst_RegFile_19_16),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_52),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR3(DLX_IDinst_RegFile_18_16),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_324)
  );
  X_BUF \DLX_IDinst_RegFile_18_16/COUTUSED  (
    .I(\DLX_IDinst_RegFile_18_16/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_265)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_265_96 (
    .IA(\DLX_IDinst_RegFile_18_16/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_264),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_324),
    .O(\DLX_IDinst_RegFile_18_16/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_18_16/CYINIT_97  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_263),
    .O(\DLX_IDinst_RegFile_18_16/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_26_24/LOGIC_ZERO_98  (
    .O(\DLX_IDinst_RegFile_26_24/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_396_99 (
    .IA(\DLX_IDinst_RegFile_26_24/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_26_24/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_455),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_396)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4551.INIT = 16'hF7B3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4551 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_55),
    .ADR2(DLX_IDinst_RegFile_25_24),
    .ADR3(DLX_IDinst_RegFile_24_24),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_455)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4561.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4561 (
    .ADR0(DLX_IDinst_RegFile_27_24),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_56),
    .ADR2(DLX_IDinst_RegFile_26_24),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_456)
  );
  X_BUF \DLX_IDinst_RegFile_26_24/COUTUSED  (
    .I(\DLX_IDinst_RegFile_26_24/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_397)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_397_100 (
    .IA(\DLX_IDinst_RegFile_26_24/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_396),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_456),
    .O(\DLX_IDinst_RegFile_26_24/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_26_24/CYINIT_101  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_395),
    .O(\DLX_IDinst_RegFile_26_24/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_26_16/LOGIC_ZERO_102  (
    .O(\DLX_IDinst_RegFile_26_16/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_268_103 (
    .IA(\DLX_IDinst_RegFile_26_16/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_26_16/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_327),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_268)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3271.INIT = 16'hF7D5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3271 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_55),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR2(DLX_IDinst_RegFile_25_16),
    .ADR3(DLX_IDinst_RegFile_24_16),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_327)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3281.INIT = 16'hBFB3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3281 (
    .ADR0(DLX_IDinst_RegFile_27_16),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_56),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR3(DLX_IDinst_RegFile_26_16),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_328)
  );
  X_BUF \DLX_IDinst_RegFile_26_16/COUTUSED  (
    .I(\DLX_IDinst_RegFile_26_16/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_269)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_269_104 (
    .IA(\DLX_IDinst_RegFile_26_16/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_268),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_328),
    .O(\DLX_IDinst_RegFile_26_16/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_26_16/CYINIT_105  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_267),
    .O(\DLX_IDinst_RegFile_26_16/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_18_25/LOGIC_ZERO_106  (
    .O(\DLX_IDinst_RegFile_18_25/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_408_107 (
    .IA(\DLX_IDinst_RegFile_18_25/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_18_25/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_467),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_408)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4671.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4671 (
    .ADR0(DLX_IDinst_RegFile_16_25),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_51),
    .ADR2(DLX_IDinst_RegFile_17_25),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_467)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4681.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4681 (
    .ADR0(DLX_IDinst_RegFile_18_25),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_52),
    .ADR2(DLX_IDinst_RegFile_19_25),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_468)
  );
  X_BUF \DLX_IDinst_RegFile_18_25/COUTUSED  (
    .I(\DLX_IDinst_RegFile_18_25/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_409)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_409_108 (
    .IA(\DLX_IDinst_RegFile_18_25/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_408),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_468),
    .O(\DLX_IDinst_RegFile_18_25/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_18_25/CYINIT_109  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_407),
    .O(\DLX_IDinst_RegFile_18_25/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_18_17/LOGIC_ZERO_110  (
    .O(\DLX_IDinst_RegFile_18_17/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_280_111 (
    .IA(\DLX_IDinst_RegFile_18_17/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_18_17/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_339),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_280)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3391.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3391 (
    .ADR0(DLX_IDinst_RegFile_16_17),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_51),
    .ADR2(DLX_IDinst_RegFile_17_17),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_339)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3401.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3401 (
    .ADR0(DLX_IDinst_RegFile_18_17),
    .ADR1(DLX_IDinst_RegFile_19_17),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_52),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_340)
  );
  X_BUF \DLX_IDinst_RegFile_18_17/COUTUSED  (
    .I(\DLX_IDinst_RegFile_18_17/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_281)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_281_112 (
    .IA(\DLX_IDinst_RegFile_18_17/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_280),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_340),
    .O(\DLX_IDinst_RegFile_18_17/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_18_17/CYINIT_113  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_279),
    .O(\DLX_IDinst_RegFile_18_17/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_26_25/LOGIC_ZERO_114  (
    .O(\DLX_IDinst_RegFile_26_25/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_412_115 (
    .IA(\DLX_IDinst_RegFile_26_25/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_26_25/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_471),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_412)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4711.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4711 (
    .ADR0(DLX_IDinst_RegFile_24_25),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_55),
    .ADR2(DLX_IDinst_RegFile_25_25),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_471)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4721.INIT = 16'hDDF5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4721 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_56),
    .ADR1(DLX_IDinst_RegFile_27_25),
    .ADR2(DLX_IDinst_RegFile_26_25),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_472)
  );
  X_BUF \DLX_IDinst_RegFile_26_25/COUTUSED  (
    .I(\DLX_IDinst_RegFile_26_25/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_413)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_413_116 (
    .IA(\DLX_IDinst_RegFile_26_25/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_412),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_472),
    .O(\DLX_IDinst_RegFile_26_25/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_26_25/CYINIT_117  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_411),
    .O(\DLX_IDinst_RegFile_26_25/CYINIT )
  );
  defparam DLX_IDinst_RegFile_25_29_118.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_25_29_118 (
    .I(DLX_IDinst_WB_data_eff[29]),
    .CE(DLX_IDinst__n0600),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_25_29)
  );
  X_ZERO \DLX_IDinst_RegFile_26_17/LOGIC_ZERO_119  (
    .O(\DLX_IDinst_RegFile_26_17/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_284_120 (
    .IA(\DLX_IDinst_RegFile_26_17/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_26_17/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_343),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_284)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3431.INIT = 16'hF5DD;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3431 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_55),
    .ADR1(DLX_IDinst_RegFile_24_17),
    .ADR2(DLX_IDinst_RegFile_25_17),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_343)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3441.INIT = 16'hE2FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3441 (
    .ADR0(DLX_IDinst_RegFile_26_17),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR2(DLX_IDinst_RegFile_27_17),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_56),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_344)
  );
  X_BUF \DLX_IDinst_RegFile_26_17/COUTUSED  (
    .I(\DLX_IDinst_RegFile_26_17/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_285)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_285_121 (
    .IA(\DLX_IDinst_RegFile_26_17/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_284),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_344),
    .O(\DLX_IDinst_RegFile_26_17/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_26_17/CYINIT_122  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_283),
    .O(\DLX_IDinst_RegFile_26_17/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_18_26/LOGIC_ZERO_123  (
    .O(\DLX_IDinst_RegFile_18_26/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_424_124 (
    .IA(\DLX_IDinst_RegFile_18_26/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_18_26/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_483),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_424)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4831.INIT = 16'hE4FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4831 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR1(DLX_IDinst_RegFile_16_26),
    .ADR2(DLX_IDinst_RegFile_17_26),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_51),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_483)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4841.INIT = 16'hF7D5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4841 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_52),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR2(DLX_IDinst_RegFile_19_26),
    .ADR3(DLX_IDinst_RegFile_18_26),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_484)
  );
  X_BUF \DLX_IDinst_RegFile_18_26/COUTUSED  (
    .I(\DLX_IDinst_RegFile_18_26/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_425)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_425_125 (
    .IA(\DLX_IDinst_RegFile_18_26/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_424),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_484),
    .O(\DLX_IDinst_RegFile_18_26/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_18_26/CYINIT_126  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_423),
    .O(\DLX_IDinst_RegFile_18_26/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_18_18/LOGIC_ZERO_127  (
    .O(\DLX_IDinst_RegFile_18_18/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_296_128 (
    .IA(\DLX_IDinst_RegFile_18_18/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_18_18/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_355),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_296)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3551.INIT = 16'hDFD5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3551 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_51),
    .ADR1(DLX_IDinst_RegFile_17_18),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR3(DLX_IDinst_RegFile_16_18),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_355)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3561.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3561 (
    .ADR0(DLX_IDinst_RegFile_18_18),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_52),
    .ADR2(DLX_IDinst_RegFile_19_18),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_356)
  );
  X_BUF \DLX_IDinst_RegFile_18_18/COUTUSED  (
    .I(\DLX_IDinst_RegFile_18_18/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_297)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_297_129 (
    .IA(\DLX_IDinst_RegFile_18_18/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_296),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_356),
    .O(\DLX_IDinst_RegFile_18_18/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_18_18/CYINIT_130  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_295),
    .O(\DLX_IDinst_RegFile_18_18/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_19_10/LOGIC_ZERO_131  (
    .O(\DLX_IDinst_RegFile_19_10/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_168_132 (
    .IA(\DLX_IDinst_RegFile_19_10/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_19_10/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_227),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_168)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2271.INIT = 16'hDF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2271 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR1(DLX_IDinst_RegFile_17_10),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_51),
    .ADR3(DLX_IDinst_RegFile_16_10),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_227)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2281.INIT = 16'hD8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2281 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR1(DLX_IDinst_RegFile_19_10),
    .ADR2(DLX_IDinst_RegFile_18_10),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_52),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_228)
  );
  X_BUF \DLX_IDinst_RegFile_19_10/COUTUSED  (
    .I(\DLX_IDinst_RegFile_19_10/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_169)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_169_133 (
    .IA(\DLX_IDinst_RegFile_19_10/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_168),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_228),
    .O(\DLX_IDinst_RegFile_19_10/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_19_10/CYINIT_134  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_167),
    .O(\DLX_IDinst_RegFile_19_10/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_26_26/LOGIC_ZERO_135  (
    .O(\DLX_IDinst_RegFile_26_26/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_428_136 (
    .IA(\DLX_IDinst_RegFile_26_26/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_26_26/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_487),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_428)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4871.INIT = 16'hFD5D;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4871 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_55),
    .ADR1(DLX_IDinst_RegFile_24_26),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR3(DLX_IDinst_RegFile_25_26),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_487)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4881.INIT = 16'hACFF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4881 (
    .ADR0(DLX_IDinst_RegFile_27_26),
    .ADR1(DLX_IDinst_RegFile_26_26),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_56),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_488)
  );
  X_BUF \DLX_IDinst_RegFile_26_26/COUTUSED  (
    .I(\DLX_IDinst_RegFile_26_26/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_429)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_429_137 (
    .IA(\DLX_IDinst_RegFile_26_26/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_428),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_488),
    .O(\DLX_IDinst_RegFile_26_26/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_26_26/CYINIT_138  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_427),
    .O(\DLX_IDinst_RegFile_26_26/CYINIT )
  );
  defparam DLX_IDinst_RegFile_26_18_139.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_26_18_139 (
    .I(DLX_IDinst_WB_data_eff[18]),
    .CE(DLX_IDinst__n0602),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_26_18)
  );
  X_ZERO \DLX_IDinst_RegFile_26_18/LOGIC_ZERO_140  (
    .O(\DLX_IDinst_RegFile_26_18/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_300_141 (
    .IA(\DLX_IDinst_RegFile_26_18/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_26_18/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_359),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_300)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3591.INIT = 16'hF5DD;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3591 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_55),
    .ADR1(DLX_IDinst_RegFile_24_18),
    .ADR2(DLX_IDinst_RegFile_25_18),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_359)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3601.INIT = 16'hDDF5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3601 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_56),
    .ADR1(DLX_IDinst_RegFile_27_18),
    .ADR2(DLX_IDinst_RegFile_26_18),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_360)
  );
  X_BUF \DLX_IDinst_RegFile_26_18/COUTUSED  (
    .I(\DLX_IDinst_RegFile_26_18/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_301)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_301_142 (
    .IA(\DLX_IDinst_RegFile_26_18/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_300),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_360),
    .O(\DLX_IDinst_RegFile_26_18/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_26_18/CYINIT_143  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_299),
    .O(\DLX_IDinst_RegFile_26_18/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_27_10/LOGIC_ZERO_144  (
    .O(\DLX_IDinst_RegFile_27_10/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_172_145 (
    .IA(\DLX_IDinst_RegFile_27_10/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_27_10/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_231),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_172)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2311.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2311 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_55),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR2(DLX_IDinst_RegFile_24_10),
    .ADR3(DLX_IDinst_RegFile_25_10),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_231)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2321.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2321 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_56),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR2(DLX_IDinst_RegFile_26_10),
    .ADR3(DLX_IDinst_RegFile_27_10),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_232)
  );
  X_BUF \DLX_IDinst_RegFile_27_10/COUTUSED  (
    .I(\DLX_IDinst_RegFile_27_10/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_173)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_173_146 (
    .IA(\DLX_IDinst_RegFile_27_10/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_172),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_232),
    .O(\DLX_IDinst_RegFile_27_10/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_27_10/CYINIT_147  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_171),
    .O(\DLX_IDinst_RegFile_27_10/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_18_27/LOGIC_ZERO_148  (
    .O(\DLX_IDinst_RegFile_18_27/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_952_149 (
    .IA(\DLX_IDinst_RegFile_18_27/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_18_27/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1027),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_952)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10271.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10271 (
    .ADR0(DLX_IDinst_jtarget[21]),
    .ADR1(DLX_IDinst_RegFile_16_27),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_579),
    .ADR3(DLX_IDinst_RegFile_17_27),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1027)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10281.INIT = 16'hF7D5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10281 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_580),
    .ADR1(DLX_IDinst_jtarget[21]),
    .ADR2(DLX_IDinst_RegFile_19_27),
    .ADR3(DLX_IDinst_RegFile_18_27),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1028)
  );
  X_BUF \DLX_IDinst_RegFile_18_27/COUTUSED  (
    .I(\DLX_IDinst_RegFile_18_27/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_953)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_953_150 (
    .IA(\DLX_IDinst_RegFile_18_27/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_952),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1028),
    .O(\DLX_IDinst_RegFile_18_27/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_18_27/CYINIT_151  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_951),
    .O(\DLX_IDinst_RegFile_18_27/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_18_19/LOGIC_ZERO_152  (
    .O(\DLX_IDinst_RegFile_18_19/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_312_153 (
    .IA(\DLX_IDinst_RegFile_18_19/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_18_19/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_371),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_312)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3711.INIT = 16'hD8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3711 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR1(DLX_IDinst_RegFile_17_19),
    .ADR2(DLX_IDinst_RegFile_16_19),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_51),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_371)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3721.INIT = 16'hCFAF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3721 (
    .ADR0(DLX_IDinst_RegFile_18_19),
    .ADR1(DLX_IDinst_RegFile_19_19),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_52),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_372)
  );
  X_BUF \DLX_IDinst_RegFile_18_19/COUTUSED  (
    .I(\DLX_IDinst_RegFile_18_19/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_313)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_313_154 (
    .IA(\DLX_IDinst_RegFile_18_19/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_312),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_372),
    .O(\DLX_IDinst_RegFile_18_19/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_18_19/CYINIT_155  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_311),
    .O(\DLX_IDinst_RegFile_18_19/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_19_11/LOGIC_ZERO_156  (
    .O(\DLX_IDinst_RegFile_19_11/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_184_157 (
    .IA(\DLX_IDinst_RegFile_19_11/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_19_11/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_243),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_184)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2431.INIT = 16'hF7B3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2431 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_51),
    .ADR2(DLX_IDinst_RegFile_17_11),
    .ADR3(DLX_IDinst_RegFile_16_11),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_243)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2441.INIT = 16'hFB3B;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2441 (
    .ADR0(DLX_IDinst_RegFile_18_11),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_52),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR3(DLX_IDinst_RegFile_19_11),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_244)
  );
  X_BUF \DLX_IDinst_RegFile_19_11/COUTUSED  (
    .I(\DLX_IDinst_RegFile_19_11/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_185)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_185_158 (
    .IA(\DLX_IDinst_RegFile_19_11/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_184),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_244),
    .O(\DLX_IDinst_RegFile_19_11/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_19_11/CYINIT_159  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_183),
    .O(\DLX_IDinst_RegFile_19_11/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_26_27/LOGIC_ZERO_160  (
    .O(\DLX_IDinst_RegFile_26_27/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_956_161 (
    .IA(\DLX_IDinst_RegFile_26_27/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_26_27/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1031),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_956)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10311.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10311 (
    .ADR0(DLX_IDinst_jtarget[21]),
    .ADR1(DLX_IDinst_RegFile_24_27),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_583),
    .ADR3(DLX_IDinst_RegFile_25_27),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1031)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10321.INIT = 16'hE4FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10321 (
    .ADR0(DLX_IDinst_jtarget[21]),
    .ADR1(DLX_IDinst_RegFile_26_27),
    .ADR2(DLX_IDinst_RegFile_27_27),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_584),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1032)
  );
  X_BUF \DLX_IDinst_RegFile_26_27/COUTUSED  (
    .I(\DLX_IDinst_RegFile_26_27/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_957)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_957_162 (
    .IA(\DLX_IDinst_RegFile_26_27/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_956),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1032),
    .O(\DLX_IDinst_RegFile_26_27/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_26_27/CYINIT_163  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_955),
    .O(\DLX_IDinst_RegFile_26_27/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_26_19/LOGIC_ZERO_164  (
    .O(\DLX_IDinst_RegFile_26_19/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_316_165 (
    .IA(\DLX_IDinst_RegFile_26_19/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_26_19/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_375),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_316)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3751.INIT = 16'hFB3B;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3751 (
    .ADR0(DLX_IDinst_RegFile_24_19),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_55),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR3(DLX_IDinst_RegFile_25_19),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_375)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3761.INIT = 16'hB8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3761 (
    .ADR0(DLX_IDinst_RegFile_27_19),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR2(DLX_IDinst_RegFile_26_19),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_56),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_376)
  );
  X_BUF \DLX_IDinst_RegFile_26_19/COUTUSED  (
    .I(\DLX_IDinst_RegFile_26_19/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_317)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_317_166 (
    .IA(\DLX_IDinst_RegFile_26_19/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_316),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_376),
    .O(\DLX_IDinst_RegFile_26_19/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_26_19/CYINIT_167  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_315),
    .O(\DLX_IDinst_RegFile_26_19/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_27_11/LOGIC_ZERO_168  (
    .O(\DLX_IDinst_RegFile_27_11/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_188_169 (
    .IA(\DLX_IDinst_RegFile_27_11/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_27_11/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_247),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_188)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2471.INIT = 16'hBFB3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2471 (
    .ADR0(DLX_IDinst_RegFile_25_11),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_55),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR3(DLX_IDinst_RegFile_24_11),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_247)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2481.INIT = 16'hAFCF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2481 (
    .ADR0(DLX_IDinst_RegFile_27_11),
    .ADR1(DLX_IDinst_RegFile_26_11),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_56),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_248)
  );
  X_BUF \DLX_IDinst_RegFile_27_11/COUTUSED  (
    .I(\DLX_IDinst_RegFile_27_11/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_189)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_189_170 (
    .IA(\DLX_IDinst_RegFile_27_11/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_188),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_248),
    .O(\DLX_IDinst_RegFile_27_11/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_27_11/CYINIT_171  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_187),
    .O(\DLX_IDinst_RegFile_27_11/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_18_28/LOGIC_ZERO_172  (
    .O(\DLX_IDinst_RegFile_18_28/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_968_173 (
    .IA(\DLX_IDinst_RegFile_18_28/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_18_28/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1043),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_968)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10431.INIT = 16'hACFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10431 (
    .ADR0(DLX_IDinst_RegFile_17_28),
    .ADR1(DLX_IDinst_RegFile_16_28),
    .ADR2(DLX_IDinst_jtarget[21]),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_579),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1043)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10441.INIT = 16'hDF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10441 (
    .ADR0(DLX_IDinst_jtarget[21]),
    .ADR1(DLX_IDinst_RegFile_19_28),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_580),
    .ADR3(DLX_IDinst_RegFile_18_28),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1044)
  );
  X_BUF \DLX_IDinst_RegFile_18_28/COUTUSED  (
    .I(\DLX_IDinst_RegFile_18_28/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_969)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_969_174 (
    .IA(\DLX_IDinst_RegFile_18_28/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_968),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1044),
    .O(\DLX_IDinst_RegFile_18_28/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_18_28/CYINIT_175  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_967),
    .O(\DLX_IDinst_RegFile_18_28/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_19_20/LOGIC_ZERO_176  (
    .O(\DLX_IDinst_RegFile_19_20/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_328_177 (
    .IA(\DLX_IDinst_RegFile_19_20/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_19_20/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_387),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_328)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3871.INIT = 16'hCFAF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3871 (
    .ADR0(DLX_IDinst_RegFile_16_20),
    .ADR1(DLX_IDinst_RegFile_17_20),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_51),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_387)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3881.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3881 (
    .ADR0(DLX_IDinst_RegFile_18_20),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_52),
    .ADR2(DLX_IDinst_RegFile_19_20),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_388)
  );
  X_BUF \DLX_IDinst_RegFile_19_20/COUTUSED  (
    .I(\DLX_IDinst_RegFile_19_20/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_329)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_329_178 (
    .IA(\DLX_IDinst_RegFile_19_20/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_328),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_388),
    .O(\DLX_IDinst_RegFile_19_20/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_19_20/CYINIT_179  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_327),
    .O(\DLX_IDinst_RegFile_19_20/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_19_12/LOGIC_ZERO_180  (
    .O(\DLX_IDinst_RegFile_19_12/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_200_181 (
    .IA(\DLX_IDinst_RegFile_19_12/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_19_12/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_259),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_200)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2591.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2591 (
    .ADR0(DLX_IDinst_RegFile_16_12),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_51),
    .ADR2(DLX_IDinst_RegFile_17_12),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_259)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2601.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2601 (
    .ADR0(DLX_IDinst_RegFile_18_12),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_52),
    .ADR3(DLX_IDinst_RegFile_19_12),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_260)
  );
  X_BUF \DLX_IDinst_RegFile_19_12/COUTUSED  (
    .I(\DLX_IDinst_RegFile_19_12/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_201)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_201_182 (
    .IA(\DLX_IDinst_RegFile_19_12/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_200),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_260),
    .O(\DLX_IDinst_RegFile_19_12/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_19_12/CYINIT_183  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_199),
    .O(\DLX_IDinst_RegFile_19_12/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_26_28/LOGIC_ZERO_184  (
    .O(\DLX_IDinst_RegFile_26_28/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_460_185 (
    .IA(\DLX_IDinst_RegFile_26_28/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_26_28/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_519),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_460)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5191.INIT = 16'hF5DD;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5191 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_55),
    .ADR1(DLX_IDinst_RegFile_24_28),
    .ADR2(DLX_IDinst_RegFile_25_28),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_519)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5201.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5201 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR1(DLX_IDinst_RegFile_26_28),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_56),
    .ADR3(DLX_IDinst_RegFile_27_28),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_520)
  );
  X_BUF \DLX_IDinst_RegFile_26_28/COUTUSED  (
    .I(\DLX_IDinst_RegFile_26_28/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_461)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_461_186 (
    .IA(\DLX_IDinst_RegFile_26_28/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_460),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_520),
    .O(\DLX_IDinst_RegFile_26_28/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_26_28/CYINIT_187  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_459),
    .O(\DLX_IDinst_RegFile_26_28/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_27_20/LOGIC_ZERO_188  (
    .O(\DLX_IDinst_RegFile_27_20/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_844_189 (
    .IA(\DLX_IDinst_RegFile_27_20/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_27_20/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_919),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_844)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9191.INIT = 16'hAFCF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9191 (
    .ADR0(DLX_IDinst_RegFile_25_20),
    .ADR1(DLX_IDinst_RegFile_24_20),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_583),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_919)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9201.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9201 (
    .ADR0(DLX_IDinst_RegFile_27_20),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_584),
    .ADR2(DLX_IDinst_RegFile_26_20),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_920)
  );
  X_BUF \DLX_IDinst_RegFile_27_20/COUTUSED  (
    .I(\DLX_IDinst_RegFile_27_20/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_845)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_845_190 (
    .IA(\DLX_IDinst_RegFile_27_20/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_844),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_920),
    .O(\DLX_IDinst_RegFile_27_20/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_27_20/CYINIT_191  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_843),
    .O(\DLX_IDinst_RegFile_27_20/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_27_12/LOGIC_ZERO_192  (
    .O(\DLX_IDinst_RegFile_27_12/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_716_193 (
    .IA(\DLX_IDinst_RegFile_27_12/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_27_12/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_791),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_716)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7911.INIT = 16'hB8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7911 (
    .ADR0(DLX_IDinst_RegFile_25_12),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR2(DLX_IDinst_RegFile_24_12),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_583),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_791)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7921.INIT = 16'hBFB3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7921 (
    .ADR0(DLX_IDinst_RegFile_27_12),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_584),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR3(DLX_IDinst_RegFile_26_12),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_792)
  );
  X_BUF \DLX_IDinst_RegFile_27_12/COUTUSED  (
    .I(\DLX_IDinst_RegFile_27_12/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_717)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_717_194 (
    .IA(\DLX_IDinst_RegFile_27_12/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_716),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_792),
    .O(\DLX_IDinst_RegFile_27_12/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_27_12/CYINIT_195  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_715),
    .O(\DLX_IDinst_RegFile_27_12/CYINIT )
  );
  defparam DLX_IDinst_RegFile_26_21_196.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_26_21_196 (
    .I(DLX_IDinst_WB_data_eff[21]),
    .CE(DLX_IDinst__n0602),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_26_21)
  );
  X_ZERO \DLX_IDinst_RegFile_18_29/LOGIC_ZERO_197  (
    .O(\DLX_IDinst_RegFile_18_29/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_472_198 (
    .IA(\DLX_IDinst_RegFile_18_29/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_18_29/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_531),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_472)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5311.INIT = 16'hDFD5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5311 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_51),
    .ADR1(DLX_IDinst_RegFile_17_29),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR3(DLX_IDinst_RegFile_16_29),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_531)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5321.INIT = 16'hACFF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5321 (
    .ADR0(DLX_IDinst_RegFile_19_29),
    .ADR1(DLX_IDinst_RegFile_18_29),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_52),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_532)
  );
  X_BUF \DLX_IDinst_RegFile_18_29/COUTUSED  (
    .I(\DLX_IDinst_RegFile_18_29/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_473)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_473_199 (
    .IA(\DLX_IDinst_RegFile_18_29/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_472),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_532),
    .O(\DLX_IDinst_RegFile_18_29/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_18_29/CYINIT_200  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_471),
    .O(\DLX_IDinst_RegFile_18_29/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_19_21/LOGIC_ZERO_201  (
    .O(\DLX_IDinst_RegFile_19_21/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_856_202 (
    .IA(\DLX_IDinst_RegFile_19_21/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_19_21/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_931),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_856)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9311.INIT = 16'hFB3B;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9311 (
    .ADR0(DLX_IDinst_RegFile_16_21),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_579),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR3(DLX_IDinst_RegFile_17_21),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_931)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9321.INIT = 16'hFD5D;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9321 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_580),
    .ADR1(DLX_IDinst_RegFile_18_21),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR3(DLX_IDinst_RegFile_19_21),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_932)
  );
  X_BUF \DLX_IDinst_RegFile_19_21/COUTUSED  (
    .I(\DLX_IDinst_RegFile_19_21/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_857)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_857_203 (
    .IA(\DLX_IDinst_RegFile_19_21/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_856),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_932),
    .O(\DLX_IDinst_RegFile_19_21/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_19_21/CYINIT_204  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_855),
    .O(\DLX_IDinst_RegFile_19_21/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_19_13/LOGIC_ZERO_205  (
    .O(\DLX_IDinst_RegFile_19_13/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_728_206 (
    .IA(\DLX_IDinst_RegFile_19_13/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_19_13/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_803),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_728)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8031.INIT = 16'hF7B3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8031 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_579),
    .ADR2(DLX_IDinst_RegFile_17_13),
    .ADR3(DLX_IDinst_RegFile_16_13),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_803)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8041.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8041 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR1(DLX_IDinst_RegFile_18_13),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_580),
    .ADR3(DLX_IDinst_RegFile_19_13),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_804)
  );
  X_BUF \DLX_IDinst_RegFile_19_13/COUTUSED  (
    .I(\DLX_IDinst_RegFile_19_13/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_729)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_729_207 (
    .IA(\DLX_IDinst_RegFile_19_13/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_728),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_804),
    .O(\DLX_IDinst_RegFile_19_13/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_19_13/CYINIT_208  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_727),
    .O(\DLX_IDinst_RegFile_19_13/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_26_29/LOGIC_ZERO_209  (
    .O(\DLX_IDinst_RegFile_26_29/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_476_210 (
    .IA(\DLX_IDinst_RegFile_26_29/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_26_29/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_535),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_476)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5351.INIT = 16'hD8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5351 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR1(DLX_IDinst_RegFile_25_29),
    .ADR2(DLX_IDinst_RegFile_24_29),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_55),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_535)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5361.INIT = 16'hDFD5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5361 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_56),
    .ADR1(DLX_IDinst_RegFile_27_29),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR3(DLX_IDinst_RegFile_26_29),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_536)
  );
  X_BUF \DLX_IDinst_RegFile_26_29/COUTUSED  (
    .I(\DLX_IDinst_RegFile_26_29/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_477)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_477_211 (
    .IA(\DLX_IDinst_RegFile_26_29/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_476),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_536),
    .O(\DLX_IDinst_RegFile_26_29/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_26_29/CYINIT_212  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_475),
    .O(\DLX_IDinst_RegFile_26_29/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_27_21/LOGIC_ZERO_213  (
    .O(\DLX_IDinst_RegFile_27_21/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_860_214 (
    .IA(\DLX_IDinst_RegFile_27_21/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_27_21/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_935),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_860)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9351.INIT = 16'hD8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9351 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR1(DLX_IDinst_RegFile_25_21),
    .ADR2(DLX_IDinst_RegFile_24_21),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_583),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_935)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9361.INIT = 16'hB8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9361 (
    .ADR0(DLX_IDinst_RegFile_27_21),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR2(DLX_IDinst_RegFile_26_21),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_584),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_936)
  );
  X_BUF \DLX_IDinst_RegFile_27_21/COUTUSED  (
    .I(\DLX_IDinst_RegFile_27_21/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_861)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_861_215 (
    .IA(\DLX_IDinst_RegFile_27_21/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_860),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_936),
    .O(\DLX_IDinst_RegFile_27_21/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_27_21/CYINIT_216  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_859),
    .O(\DLX_IDinst_RegFile_27_21/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_27_13/LOGIC_ZERO_217  (
    .O(\DLX_IDinst_RegFile_27_13/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_732_218 (
    .IA(\DLX_IDinst_RegFile_27_13/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_27_13/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_807),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_732)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8071.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8071 (
    .ADR0(DLX_IDinst_RegFile_25_13),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_583),
    .ADR2(DLX_IDinst_RegFile_24_13),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_807)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8081.INIT = 16'hE2FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8081 (
    .ADR0(DLX_IDinst_RegFile_26_13),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR2(DLX_IDinst_RegFile_27_13),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_584),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_808)
  );
  X_BUF \DLX_IDinst_RegFile_27_13/COUTUSED  (
    .I(\DLX_IDinst_RegFile_27_13/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_733)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_733_219 (
    .IA(\DLX_IDinst_RegFile_27_13/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_732),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_808),
    .O(\DLX_IDinst_RegFile_27_13/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_27_13/CYINIT_220  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_731),
    .O(\DLX_IDinst_RegFile_27_13/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_19_30/LOGIC_ZERO_221  (
    .O(\DLX_IDinst_RegFile_19_30/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_488_222 (
    .IA(\DLX_IDinst_RegFile_19_30/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_19_30/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_547),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_488)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5471.INIT = 16'hAFCF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5471 (
    .ADR0(DLX_IDinst_RegFile_17_30),
    .ADR1(DLX_IDinst_RegFile_16_30),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_51),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_547)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5481.INIT = 16'hB8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5481 (
    .ADR0(DLX_IDinst_RegFile_19_30),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR2(DLX_IDinst_RegFile_18_30),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_52),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_548)
  );
  X_BUF \DLX_IDinst_RegFile_19_30/COUTUSED  (
    .I(\DLX_IDinst_RegFile_19_30/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_489)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_489_223 (
    .IA(\DLX_IDinst_RegFile_19_30/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_488),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_548),
    .O(\DLX_IDinst_RegFile_19_30/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_19_30/CYINIT_224  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_487),
    .O(\DLX_IDinst_RegFile_19_30/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_19_22/LOGIC_ZERO_225  (
    .O(\DLX_IDinst_RegFile_19_22/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_872_226 (
    .IA(\DLX_IDinst_RegFile_19_22/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_19_22/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_947),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_872)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9471.INIT = 16'hF7D5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9471 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_579),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR2(DLX_IDinst_RegFile_17_22),
    .ADR3(DLX_IDinst_RegFile_16_22),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_947)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9481.INIT = 16'hE4FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9481 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR1(DLX_IDinst_RegFile_18_22),
    .ADR2(DLX_IDinst_RegFile_19_22),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_580),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_948)
  );
  X_BUF \DLX_IDinst_RegFile_19_22/COUTUSED  (
    .I(\DLX_IDinst_RegFile_19_22/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_873)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_873_227 (
    .IA(\DLX_IDinst_RegFile_19_22/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_872),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_948),
    .O(\DLX_IDinst_RegFile_19_22/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_19_22/CYINIT_228  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_871),
    .O(\DLX_IDinst_RegFile_19_22/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_19_14/LOGIC_ZERO_229  (
    .O(\DLX_IDinst_RegFile_19_14/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_744_230 (
    .IA(\DLX_IDinst_RegFile_19_14/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_19_14/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_819),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_744)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8191.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8191 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_579),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR2(DLX_IDinst_RegFile_16_14),
    .ADR3(DLX_IDinst_RegFile_17_14),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_819)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8201.INIT = 16'hFB3B;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8201 (
    .ADR0(DLX_IDinst_RegFile_18_14),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_580),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR3(DLX_IDinst_RegFile_19_14),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_820)
  );
  X_BUF \DLX_IDinst_RegFile_19_14/COUTUSED  (
    .I(\DLX_IDinst_RegFile_19_14/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_745)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_745_231 (
    .IA(\DLX_IDinst_RegFile_19_14/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_744),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_820),
    .O(\DLX_IDinst_RegFile_19_14/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_19_14/CYINIT_232  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_743),
    .O(\DLX_IDinst_RegFile_19_14/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_27_30/LOGIC_ZERO_233  (
    .O(\DLX_IDinst_RegFile_27_30/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_492_234 (
    .IA(\DLX_IDinst_RegFile_27_30/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_27_30/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_551),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_492)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5511.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5511 (
    .ADR0(DLX_IDinst_RegFile_24_30),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_55),
    .ADR3(DLX_IDinst_RegFile_25_30),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_551)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5521.INIT = 16'hF7B3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5521 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_56),
    .ADR2(DLX_IDinst_RegFile_27_30),
    .ADR3(DLX_IDinst_RegFile_26_30),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_552)
  );
  X_BUF \DLX_IDinst_RegFile_27_30/COUTUSED  (
    .I(\DLX_IDinst_RegFile_27_30/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_493)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_493_235 (
    .IA(\DLX_IDinst_RegFile_27_30/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_492),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_552),
    .O(\DLX_IDinst_RegFile_27_30/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_27_30/CYINIT_236  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_491),
    .O(\DLX_IDinst_RegFile_27_30/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_27_22/LOGIC_ZERO_237  (
    .O(\DLX_IDinst_RegFile_27_22/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_876_238 (
    .IA(\DLX_IDinst_RegFile_27_22/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_27_22/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_951),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_876)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9511.INIT = 16'hF7B3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9511 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_583),
    .ADR2(DLX_IDinst_RegFile_25_22),
    .ADR3(DLX_IDinst_RegFile_24_22),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_951)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9521.INIT = 16'hE4FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9521 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR1(DLX_IDinst_RegFile_26_22),
    .ADR2(DLX_IDinst_RegFile_27_22),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_584),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_952)
  );
  X_BUF \DLX_IDinst_RegFile_27_22/COUTUSED  (
    .I(\DLX_IDinst_RegFile_27_22/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_877)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_877_239 (
    .IA(\DLX_IDinst_RegFile_27_22/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_876),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_952),
    .O(\DLX_IDinst_RegFile_27_22/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_27_22/CYINIT_240  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_875),
    .O(\DLX_IDinst_RegFile_27_22/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_27_14/LOGIC_ZERO_241  (
    .O(\DLX_IDinst_RegFile_27_14/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_748_242 (
    .IA(\DLX_IDinst_RegFile_27_14/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_27_14/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_823),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_748)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8231.INIT = 16'hE4FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8231 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR1(DLX_IDinst_RegFile_24_14),
    .ADR2(DLX_IDinst_RegFile_25_14),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_583),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_823)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8241.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8241 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_584),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR2(DLX_IDinst_RegFile_26_14),
    .ADR3(DLX_IDinst_RegFile_27_14),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_824)
  );
  X_BUF \DLX_IDinst_RegFile_27_14/COUTUSED  (
    .I(\DLX_IDinst_RegFile_27_14/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_749)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_749_243 (
    .IA(\DLX_IDinst_RegFile_27_14/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_748),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_824),
    .O(\DLX_IDinst_RegFile_27_14/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_27_14/CYINIT_244  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_747),
    .O(\DLX_IDinst_RegFile_27_14/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_19_23/LOGIC_ZERO_245  (
    .O(\DLX_IDinst_RegFile_19_23/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_888_246 (
    .IA(\DLX_IDinst_RegFile_19_23/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_19_23/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_963),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_888)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9631.INIT = 16'hAFCF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9631 (
    .ADR0(DLX_IDinst_RegFile_17_23),
    .ADR1(DLX_IDinst_RegFile_16_23),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_579),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_963)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9641.INIT = 16'hE2FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9641 (
    .ADR0(DLX_IDinst_RegFile_18_23),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR2(DLX_IDinst_RegFile_19_23),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_580),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_964)
  );
  X_BUF \DLX_IDinst_RegFile_19_23/COUTUSED  (
    .I(\DLX_IDinst_RegFile_19_23/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_889)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_889_247 (
    .IA(\DLX_IDinst_RegFile_19_23/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_888),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_964),
    .O(\DLX_IDinst_RegFile_19_23/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_19_23/CYINIT_248  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_887),
    .O(\DLX_IDinst_RegFile_19_23/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_19_15/LOGIC_ZERO_249  (
    .O(\DLX_IDinst_RegFile_19_15/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_760_250 (
    .IA(\DLX_IDinst_RegFile_19_15/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_19_15/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_835),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_760)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8351.INIT = 16'hF7B3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8351 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_579),
    .ADR2(DLX_IDinst_RegFile_17_15),
    .ADR3(DLX_IDinst_RegFile_16_15),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_835)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8361.INIT = 16'hDF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8361 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR1(DLX_IDinst_RegFile_19_15),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_580),
    .ADR3(DLX_IDinst_RegFile_18_15),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_836)
  );
  X_BUF \DLX_IDinst_RegFile_19_15/COUTUSED  (
    .I(\DLX_IDinst_RegFile_19_15/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_761)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_761_251 (
    .IA(\DLX_IDinst_RegFile_19_15/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_760),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_836),
    .O(\DLX_IDinst_RegFile_19_15/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_19_15/CYINIT_252  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_759),
    .O(\DLX_IDinst_RegFile_19_15/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_27_15/LOGIC_ZERO_253  (
    .O(\DLX_IDinst_RegFile_27_15/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_764_254 (
    .IA(\DLX_IDinst_RegFile_27_15/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_27_15/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_839),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_764)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8391.INIT = 16'hCFAF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8391 (
    .ADR0(DLX_IDinst_RegFile_24_15),
    .ADR1(DLX_IDinst_RegFile_25_15),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_583),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_839)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8401.INIT = 16'hDDF5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8401 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_584),
    .ADR1(DLX_IDinst_RegFile_27_15),
    .ADR2(DLX_IDinst_RegFile_26_15),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_840)
  );
  X_BUF \DLX_IDinst_RegFile_27_15/COUTUSED  (
    .I(\DLX_IDinst_RegFile_27_15/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_765)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_765_255 (
    .IA(\DLX_IDinst_RegFile_27_15/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_764),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_840),
    .O(\DLX_IDinst_RegFile_27_15/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_27_15/CYINIT_256  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_763),
    .O(\DLX_IDinst_RegFile_27_15/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_19_31/LOGIC_ZERO_257  (
    .O(\DLX_IDinst_RegFile_19_31/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_504_258 (
    .IA(\DLX_IDinst_RegFile_19_31/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_19_31/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_563),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_504)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5631.INIT = 16'hE2FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5631 (
    .ADR0(DLX_IDinst_RegFile_16_31),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR2(DLX_IDinst_RegFile_17_31),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_51),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_563)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5641.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5641 (
    .ADR0(DLX_IDinst_RegFile_18_31),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_52),
    .ADR3(DLX_IDinst_RegFile_19_31),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_564)
  );
  X_BUF \DLX_IDinst_RegFile_19_31/COUTUSED  (
    .I(\DLX_IDinst_RegFile_19_31/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_505)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_505_259 (
    .IA(\DLX_IDinst_RegFile_19_31/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_504),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_564),
    .O(\DLX_IDinst_RegFile_19_31/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_19_31/CYINIT_260  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_503),
    .O(\DLX_IDinst_RegFile_19_31/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_27_31/LOGIC_ZERO_261  (
    .O(\DLX_IDinst_RegFile_27_31/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_508_262 (
    .IA(\DLX_IDinst_RegFile_27_31/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_27_31/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_567),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_508)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5671.INIT = 16'hE4FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5671 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR1(DLX_IDinst_RegFile_24_31),
    .ADR2(DLX_IDinst_RegFile_25_31),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_55),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_567)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5681.INIT = 16'hBF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5681 (
    .ADR0(DLX_IDinst_RegFile_27_31),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_56),
    .ADR3(DLX_IDinst_RegFile_26_31),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_568)
  );
  X_BUF \DLX_IDinst_RegFile_27_31/COUTUSED  (
    .I(\DLX_IDinst_RegFile_27_31/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_509)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_509_263 (
    .IA(\DLX_IDinst_RegFile_27_31/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_508),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_568),
    .O(\DLX_IDinst_RegFile_27_31/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_27_31/CYINIT_264  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_507),
    .O(\DLX_IDinst_RegFile_27_31/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_19_24/LOGIC_ZERO_265  (
    .O(\DLX_IDinst_RegFile_19_24/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_904_266 (
    .IA(\DLX_IDinst_RegFile_19_24/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_19_24/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_979),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_904)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9791.INIT = 16'hDFD5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9791 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_579),
    .ADR1(DLX_IDinst_RegFile_17_24),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR3(DLX_IDinst_RegFile_16_24),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_979)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9801.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9801 (
    .ADR0(DLX_IDinst_RegFile_18_24),
    .ADR1(DLX_IDinst_RegFile_19_24),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_580),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_980)
  );
  X_BUF \DLX_IDinst_RegFile_19_24/COUTUSED  (
    .I(\DLX_IDinst_RegFile_19_24/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_905)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_905_267 (
    .IA(\DLX_IDinst_RegFile_19_24/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_904),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_980),
    .O(\DLX_IDinst_RegFile_19_24/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_19_24/CYINIT_268  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_903),
    .O(\DLX_IDinst_RegFile_19_24/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_19_16/LOGIC_ZERO_269  (
    .O(\DLX_IDinst_RegFile_19_16/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_776_270 (
    .IA(\DLX_IDinst_RegFile_19_16/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_19_16/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_851),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_776)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8511.INIT = 16'hE4FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8511 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR1(DLX_IDinst_RegFile_16_16),
    .ADR2(DLX_IDinst_RegFile_17_16),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_579),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_851)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8521.INIT = 16'hFD5D;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8521 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_580),
    .ADR1(DLX_IDinst_RegFile_18_16),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR3(DLX_IDinst_RegFile_19_16),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_852)
  );
  X_BUF \DLX_IDinst_RegFile_19_16/COUTUSED  (
    .I(\DLX_IDinst_RegFile_19_16/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_777)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_777_271 (
    .IA(\DLX_IDinst_RegFile_19_16/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_776),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_852),
    .O(\DLX_IDinst_RegFile_19_16/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_19_16/CYINIT_272  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_775),
    .O(\DLX_IDinst_RegFile_19_16/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_27_24/LOGIC_ZERO_273  (
    .O(\DLX_IDinst_RegFile_27_24/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_908_274 (
    .IA(\DLX_IDinst_RegFile_27_24/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_27_24/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_983),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_908)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9831.INIT = 16'hFD5D;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9831 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_583),
    .ADR1(DLX_IDinst_RegFile_24_24),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR3(DLX_IDinst_RegFile_25_24),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_983)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9841.INIT = 16'hCFAF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9841 (
    .ADR0(DLX_IDinst_RegFile_26_24),
    .ADR1(DLX_IDinst_RegFile_27_24),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_584),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_984)
  );
  X_BUF \DLX_IDinst_RegFile_27_24/COUTUSED  (
    .I(\DLX_IDinst_RegFile_27_24/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_909)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_909_275 (
    .IA(\DLX_IDinst_RegFile_27_24/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_908),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_984),
    .O(\DLX_IDinst_RegFile_27_24/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_27_24/CYINIT_276  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_907),
    .O(\DLX_IDinst_RegFile_27_24/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_27_16/LOGIC_ZERO_277  (
    .O(\DLX_IDinst_RegFile_27_16/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_780_278 (
    .IA(\DLX_IDinst_RegFile_27_16/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_27_16/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_855),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_780)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8551.INIT = 16'hF5DD;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8551 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_583),
    .ADR1(DLX_IDinst_RegFile_24_16),
    .ADR2(DLX_IDinst_RegFile_25_16),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_855)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8561.INIT = 16'hACFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8561 (
    .ADR0(DLX_IDinst_RegFile_27_16),
    .ADR1(DLX_IDinst_RegFile_26_16),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_584),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_856)
  );
  X_BUF \DLX_IDinst_RegFile_27_16/COUTUSED  (
    .I(\DLX_IDinst_RegFile_27_16/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_781)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_781_279 (
    .IA(\DLX_IDinst_RegFile_27_16/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_780),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_856),
    .O(\DLX_IDinst_RegFile_27_16/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_27_16/CYINIT_280  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_779),
    .O(\DLX_IDinst_RegFile_27_16/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_19_25/LOGIC_ZERO_281  (
    .O(\DLX_IDinst_RegFile_19_25/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_920_282 (
    .IA(\DLX_IDinst_RegFile_19_25/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_19_25/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_995),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_920)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9951.INIT = 16'hDF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9951 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR1(DLX_IDinst_RegFile_17_25),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_579),
    .ADR3(DLX_IDinst_RegFile_16_25),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_995)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9961.INIT = 16'hF5DD;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9961 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_580),
    .ADR1(DLX_IDinst_RegFile_18_25),
    .ADR2(DLX_IDinst_RegFile_19_25),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_996)
  );
  X_BUF \DLX_IDinst_RegFile_19_25/COUTUSED  (
    .I(\DLX_IDinst_RegFile_19_25/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_921)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_921_283 (
    .IA(\DLX_IDinst_RegFile_19_25/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_920),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_996),
    .O(\DLX_IDinst_RegFile_19_25/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_19_25/CYINIT_284  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_919),
    .O(\DLX_IDinst_RegFile_19_25/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_19_17/LOGIC_ZERO_285  (
    .O(\DLX_IDinst_RegFile_19_17/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_792_286 (
    .IA(\DLX_IDinst_RegFile_19_17/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_19_17/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_867),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_792)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8671.INIT = 16'hF7D5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8671 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_579),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR2(DLX_IDinst_RegFile_17_17),
    .ADR3(DLX_IDinst_RegFile_16_17),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_867)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8681.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8681 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR1(DLX_IDinst_RegFile_18_17),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_580),
    .ADR3(DLX_IDinst_RegFile_19_17),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_868)
  );
  X_BUF \DLX_IDinst_RegFile_19_17/COUTUSED  (
    .I(\DLX_IDinst_RegFile_19_17/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_793)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_793_287 (
    .IA(\DLX_IDinst_RegFile_19_17/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_792),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_868),
    .O(\DLX_IDinst_RegFile_19_17/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_19_17/CYINIT_288  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_791),
    .O(\DLX_IDinst_RegFile_19_17/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_27_17/LOGIC_ZERO_289  (
    .O(\DLX_IDinst_RegFile_27_17/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_796_290 (
    .IA(\DLX_IDinst_RegFile_27_17/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_27_17/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_871),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_796)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8711.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8711 (
    .ADR0(DLX_IDinst_RegFile_24_17),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_583),
    .ADR3(DLX_IDinst_RegFile_25_17),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_871)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8721.INIT = 16'hFB73;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8721 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_584),
    .ADR2(DLX_IDinst_RegFile_26_17),
    .ADR3(DLX_IDinst_RegFile_27_17),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_872)
  );
  X_BUF \DLX_IDinst_RegFile_27_17/COUTUSED  (
    .I(\DLX_IDinst_RegFile_27_17/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_797)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_797_291 (
    .IA(\DLX_IDinst_RegFile_27_17/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_796),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_872),
    .O(\DLX_IDinst_RegFile_27_17/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_27_17/CYINIT_292  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_795),
    .O(\DLX_IDinst_RegFile_27_17/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_19_26/LOGIC_ZERO_293  (
    .O(\DLX_IDinst_RegFile_19_26/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_936_294 (
    .IA(\DLX_IDinst_RegFile_19_26/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_19_26/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1011),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_936)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10111.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10111 (
    .ADR0(DLX_IDinst_RegFile_17_26),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_579),
    .ADR2(DLX_IDinst_RegFile_16_26),
    .ADR3(DLX_IDinst_jtarget[21]),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1011)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10121.INIT = 16'hF5DD;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10121 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_580),
    .ADR1(DLX_IDinst_RegFile_18_26),
    .ADR2(DLX_IDinst_RegFile_19_26),
    .ADR3(DLX_IDinst_jtarget[21]),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1012)
  );
  X_BUF \DLX_IDinst_RegFile_19_26/COUTUSED  (
    .I(\DLX_IDinst_RegFile_19_26/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_937)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_937_295 (
    .IA(\DLX_IDinst_RegFile_19_26/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_936),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1012),
    .O(\DLX_IDinst_RegFile_19_26/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_19_26/CYINIT_296  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_935),
    .O(\DLX_IDinst_RegFile_19_26/CYINIT )
  );
  defparam DLX_IDinst_RegFile_26_13_297.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_26_13_297 (
    .I(DLX_IDinst_WB_data_eff[13]),
    .CE(DLX_IDinst__n0602),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_26_13)
  );
  X_ZERO \DLX_IDinst_RegFile_19_18/LOGIC_ZERO_298  (
    .O(\DLX_IDinst_RegFile_19_18/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_808_299 (
    .IA(\DLX_IDinst_RegFile_19_18/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_19_18/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_883),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_808)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8831.INIT = 16'hDF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8831 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR1(DLX_IDinst_RegFile_17_18),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_579),
    .ADR3(DLX_IDinst_RegFile_16_18),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_883)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8841.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8841 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_580),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR2(DLX_IDinst_RegFile_18_18),
    .ADR3(DLX_IDinst_RegFile_19_18),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_884)
  );
  X_BUF \DLX_IDinst_RegFile_19_18/COUTUSED  (
    .I(\DLX_IDinst_RegFile_19_18/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_809)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_809_300 (
    .IA(\DLX_IDinst_RegFile_19_18/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_808),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_884),
    .O(\DLX_IDinst_RegFile_19_18/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_19_18/CYINIT_301  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_807),
    .O(\DLX_IDinst_RegFile_19_18/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_27_26/LOGIC_ZERO_302  (
    .O(\DLX_IDinst_RegFile_27_26/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_940_303 (
    .IA(\DLX_IDinst_RegFile_27_26/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_27_26/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1015),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_940)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10151.INIT = 16'hAFCF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10151 (
    .ADR0(DLX_IDinst_RegFile_25_26),
    .ADR1(DLX_IDinst_RegFile_24_26),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_583),
    .ADR3(DLX_IDinst_jtarget[21]),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1015)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10161.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10161 (
    .ADR0(DLX_IDinst_RegFile_26_26),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_584),
    .ADR2(DLX_IDinst_RegFile_27_26),
    .ADR3(DLX_IDinst_jtarget[21]),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1016)
  );
  X_BUF \DLX_IDinst_RegFile_27_26/COUTUSED  (
    .I(\DLX_IDinst_RegFile_27_26/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_941)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_941_304 (
    .IA(\DLX_IDinst_RegFile_27_26/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_940),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1016),
    .O(\DLX_IDinst_RegFile_27_26/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_27_26/CYINIT_305  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_939),
    .O(\DLX_IDinst_RegFile_27_26/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_27_18/LOGIC_ZERO_306  (
    .O(\DLX_IDinst_RegFile_27_18/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_812_307 (
    .IA(\DLX_IDinst_RegFile_27_18/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_27_18/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_887),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_812)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8871.INIT = 16'hDFD5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8871 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_583),
    .ADR1(DLX_IDinst_RegFile_25_18),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR3(DLX_IDinst_RegFile_24_18),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_887)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8881.INIT = 16'hDF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8881 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR1(DLX_IDinst_RegFile_27_18),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_584),
    .ADR3(DLX_IDinst_RegFile_26_18),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_888)
  );
  X_BUF \DLX_IDinst_RegFile_27_18/COUTUSED  (
    .I(\DLX_IDinst_RegFile_27_18/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_813)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_813_308 (
    .IA(\DLX_IDinst_RegFile_27_18/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_812),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_888),
    .O(\DLX_IDinst_RegFile_27_18/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_27_18/CYINIT_309  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_811),
    .O(\DLX_IDinst_RegFile_27_18/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_28_10/LOGIC_ZERO_310  (
    .O(\DLX_IDinst_RegFile_28_10/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_174_311 (
    .IA(\DLX_IDinst_RegFile_28_10/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_28_10/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_233),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_174)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2331.INIT = 16'hDDF5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2331 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_57),
    .ADR1(DLX_IDinst_RegFile_29_10),
    .ADR2(DLX_IDinst_RegFile_28_10),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_233)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2341.INIT = 16'hF5DD;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2341 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_58),
    .ADR1(DLX_IDinst_RegFile_30_10),
    .ADR2(DLX_IDinst_RegFile_31_10),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_234)
  );
  X_BUF \DLX_IDinst_RegFile_28_10/COUTUSED  (
    .I(\DLX_IDinst_RegFile_28_10/CYMUXG ),
    .O(DLX_IDinst__n0623[10])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_175 (
    .IA(\DLX_IDinst_RegFile_28_10/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_174),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_234),
    .O(\DLX_IDinst_RegFile_28_10/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_28_10/CYINIT_312  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_173),
    .O(\DLX_IDinst_RegFile_28_10/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_19_27/LOGIC_ZERO_313  (
    .O(\DLX_IDinst_RegFile_19_27/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_440_314 (
    .IA(\DLX_IDinst_RegFile_19_27/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_19_27/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_499),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_440)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4991.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4991 (
    .ADR0(DLX_IDinst_RegFile_16_27),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_51),
    .ADR3(DLX_IDinst_RegFile_17_27),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_499)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5001.INIT = 16'hACFF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5001 (
    .ADR0(DLX_IDinst_RegFile_19_27),
    .ADR1(DLX_IDinst_RegFile_18_27),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_52),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_500)
  );
  X_BUF \DLX_IDinst_RegFile_19_27/COUTUSED  (
    .I(\DLX_IDinst_RegFile_19_27/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_441)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_441_315 (
    .IA(\DLX_IDinst_RegFile_19_27/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_440),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_500),
    .O(\DLX_IDinst_RegFile_19_27/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_19_27/CYINIT_316  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_439),
    .O(\DLX_IDinst_RegFile_19_27/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_19_19/LOGIC_ZERO_317  (
    .O(\DLX_IDinst_RegFile_19_19/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_824_318 (
    .IA(\DLX_IDinst_RegFile_19_19/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_19_19/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_899),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_824)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8991.INIT = 16'hCFAF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8991 (
    .ADR0(DLX_IDinst_RegFile_16_19),
    .ADR1(DLX_IDinst_RegFile_17_19),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_579),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_899)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9001.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9001 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR1(DLX_IDinst_RegFile_18_19),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_580),
    .ADR3(DLX_IDinst_RegFile_19_19),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_900)
  );
  X_BUF \DLX_IDinst_RegFile_19_19/COUTUSED  (
    .I(\DLX_IDinst_RegFile_19_19/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_825)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_825_319 (
    .IA(\DLX_IDinst_RegFile_19_19/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_824),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_900),
    .O(\DLX_IDinst_RegFile_19_19/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_19_19/CYINIT_320  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_823),
    .O(\DLX_IDinst_RegFile_19_19/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_27_27/LOGIC_ZERO_321  (
    .O(\DLX_IDinst_RegFile_27_27/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_444_322 (
    .IA(\DLX_IDinst_RegFile_27_27/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_27_27/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_503),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_444)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5031.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5031 (
    .ADR0(DLX_IDinst_RegFile_24_27),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_55),
    .ADR3(DLX_IDinst_RegFile_25_27),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_503)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5041.INIT = 16'hCFAF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5041 (
    .ADR0(DLX_IDinst_RegFile_26_27),
    .ADR1(DLX_IDinst_RegFile_27_27),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_56),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_504)
  );
  X_BUF \DLX_IDinst_RegFile_27_27/COUTUSED  (
    .I(\DLX_IDinst_RegFile_27_27/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_445)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_445_323 (
    .IA(\DLX_IDinst_RegFile_27_27/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_444),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_504),
    .O(\DLX_IDinst_RegFile_27_27/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_27_27/CYINIT_324  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_443),
    .O(\DLX_IDinst_RegFile_27_27/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_27_19/LOGIC_ZERO_325  (
    .O(\DLX_IDinst_RegFile_27_19/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_828_326 (
    .IA(\DLX_IDinst_RegFile_27_19/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_27_19/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_903),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_828)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9031.INIT = 16'hB8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9031 (
    .ADR0(DLX_IDinst_RegFile_25_19),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR2(DLX_IDinst_RegFile_24_19),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_583),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_903)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9041.INIT = 16'hF7D5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9041 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_584),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR2(DLX_IDinst_RegFile_27_19),
    .ADR3(DLX_IDinst_RegFile_26_19),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_904)
  );
  X_BUF \DLX_IDinst_RegFile_27_19/COUTUSED  (
    .I(\DLX_IDinst_RegFile_27_19/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_829)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_829_327 (
    .IA(\DLX_IDinst_RegFile_27_19/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_828),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_904),
    .O(\DLX_IDinst_RegFile_27_19/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_27_19/CYINIT_328  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_827),
    .O(\DLX_IDinst_RegFile_27_19/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_28_11/LOGIC_ZERO_329  (
    .O(\DLX_IDinst_RegFile_28_11/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_190_330 (
    .IA(\DLX_IDinst_RegFile_28_11/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_28_11/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_249),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_190)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2491.INIT = 16'hCFAF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2491 (
    .ADR0(DLX_IDinst_RegFile_28_11),
    .ADR1(DLX_IDinst_RegFile_29_11),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_57),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_249)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2501.INIT = 16'hF5DD;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2501 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_58),
    .ADR1(DLX_IDinst_RegFile_30_11),
    .ADR2(DLX_IDinst_RegFile_31_11),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_250)
  );
  X_BUF \DLX_IDinst_RegFile_28_11/COUTUSED  (
    .I(\DLX_IDinst_RegFile_28_11/CYMUXG ),
    .O(DLX_IDinst__n0623[11])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_191 (
    .IA(\DLX_IDinst_RegFile_28_11/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_190),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_250),
    .O(\DLX_IDinst_RegFile_28_11/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_28_11/CYINIT_331  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_189),
    .O(\DLX_IDinst_RegFile_28_11/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_19_28/LOGIC_ZERO_332  (
    .O(\DLX_IDinst_RegFile_19_28/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_456_333 (
    .IA(\DLX_IDinst_RegFile_19_28/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_19_28/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_515),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_456)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5151.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5151 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR1(DLX_IDinst_RegFile_16_28),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_51),
    .ADR3(DLX_IDinst_RegFile_17_28),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_515)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5161.INIT = 16'hE2FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5161 (
    .ADR0(DLX_IDinst_RegFile_18_28),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR2(DLX_IDinst_RegFile_19_28),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_52),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_516)
  );
  X_BUF \DLX_IDinst_RegFile_19_28/COUTUSED  (
    .I(\DLX_IDinst_RegFile_19_28/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_457)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_457_334 (
    .IA(\DLX_IDinst_RegFile_19_28/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_456),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_516),
    .O(\DLX_IDinst_RegFile_19_28/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_19_28/CYINIT_335  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_455),
    .O(\DLX_IDinst_RegFile_19_28/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_28_20/LOGIC_ZERO_336  (
    .O(\DLX_IDinst_RegFile_28_20/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_334_337 (
    .IA(\DLX_IDinst_RegFile_28_20/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_28_20/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_393),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_334)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3931.INIT = 16'hD8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3931 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR1(DLX_IDinst_RegFile_29_20),
    .ADR2(DLX_IDinst_RegFile_28_20),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_57),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_393)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3941.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3941 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR1(DLX_IDinst_RegFile_30_20),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_58),
    .ADR3(DLX_IDinst_RegFile_31_20),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_394)
  );
  X_BUF \DLX_IDinst_RegFile_28_20/COUTUSED  (
    .I(\DLX_IDinst_RegFile_28_20/CYMUXG ),
    .O(DLX_IDinst__n0623[20])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_335 (
    .IA(\DLX_IDinst_RegFile_28_20/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_334),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_394),
    .O(\DLX_IDinst_RegFile_28_20/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_28_20/CYINIT_338  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_333),
    .O(\DLX_IDinst_RegFile_28_20/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_28_12/LOGIC_ZERO_339  (
    .O(\DLX_IDinst_RegFile_28_12/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_206_340 (
    .IA(\DLX_IDinst_RegFile_28_12/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_28_12/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_265),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_206)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2651.INIT = 16'hFD5D;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2651 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_57),
    .ADR1(DLX_IDinst_RegFile_28_12),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR3(DLX_IDinst_RegFile_29_12),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_265)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2661.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2661 (
    .ADR0(DLX_IDinst_RegFile_30_12),
    .ADR1(DLX_IDinst_RegFile_31_12),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_58),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_266)
  );
  X_BUF \DLX_IDinst_RegFile_28_12/COUTUSED  (
    .I(\DLX_IDinst_RegFile_28_12/CYMUXG ),
    .O(DLX_IDinst__n0623[12])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_207 (
    .IA(\DLX_IDinst_RegFile_28_12/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_206),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_266),
    .O(\DLX_IDinst_RegFile_28_12/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_28_12/CYINIT_341  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_205),
    .O(\DLX_IDinst_RegFile_28_12/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_28_21/LOGIC_ZERO_342  (
    .O(\DLX_IDinst_RegFile_28_21/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_350_343 (
    .IA(\DLX_IDinst_RegFile_28_21/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_28_21/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_409),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_350)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4091.INIT = 16'hCFAF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4091 (
    .ADR0(DLX_IDinst_RegFile_28_21),
    .ADR1(DLX_IDinst_RegFile_29_21),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_57),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_409)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4101.INIT = 16'hF7B3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4101 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_58),
    .ADR2(DLX_IDinst_RegFile_31_21),
    .ADR3(DLX_IDinst_RegFile_30_21),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_410)
  );
  X_BUF \DLX_IDinst_RegFile_28_21/COUTUSED  (
    .I(\DLX_IDinst_RegFile_28_21/CYMUXG ),
    .O(DLX_IDinst__n0623[21])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_351 (
    .IA(\DLX_IDinst_RegFile_28_21/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_350),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_410),
    .O(\DLX_IDinst_RegFile_28_21/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_28_21/CYINIT_344  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_349),
    .O(\DLX_IDinst_RegFile_28_21/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_28_13/LOGIC_ZERO_345  (
    .O(\DLX_IDinst_RegFile_28_13/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_222_346 (
    .IA(\DLX_IDinst_RegFile_28_13/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_28_13/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_281),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_222)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2811.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2811 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR1(DLX_IDinst_RegFile_28_13),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_57),
    .ADR3(DLX_IDinst_RegFile_29_13),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_281)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2821.INIT = 16'hACFF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2821 (
    .ADR0(DLX_IDinst_RegFile_31_13),
    .ADR1(DLX_IDinst_RegFile_30_13),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_58),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_282)
  );
  X_BUF \DLX_IDinst_RegFile_28_13/COUTUSED  (
    .I(\DLX_IDinst_RegFile_28_13/CYMUXG ),
    .O(DLX_IDinst__n0623[13])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_223 (
    .IA(\DLX_IDinst_RegFile_28_13/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_222),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_282),
    .O(\DLX_IDinst_RegFile_28_13/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_28_13/CYINIT_347  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_221),
    .O(\DLX_IDinst_RegFile_28_13/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_28_30/LOGIC_ZERO_348  (
    .O(\DLX_IDinst_RegFile_28_30/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_1006_349 (
    .IA(\DLX_IDinst_RegFile_28_30/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_28_30/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1081),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_1006)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10811.INIT = 16'hACFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10811 (
    .ADR0(DLX_IDinst_RegFile_29_30),
    .ADR1(DLX_IDinst_RegFile_28_30),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_585),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1081)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10821.INIT = 16'hBFB3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10821 (
    .ADR0(DLX_IDinst_RegFile_31_30),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_586),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR3(DLX_IDinst_RegFile_30_30),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1082)
  );
  X_BUF \DLX_IDinst_RegFile_28_30/COUTUSED  (
    .I(\DLX_IDinst_RegFile_28_30/CYMUXG ),
    .O(DLX_IDinst__n0620[30])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_1007 (
    .IA(\DLX_IDinst_RegFile_28_30/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_1006),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1082),
    .O(\DLX_IDinst_RegFile_28_30/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_28_30/CYINIT_350  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_1005),
    .O(\DLX_IDinst_RegFile_28_30/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_28_22/LOGIC_ZERO_351  (
    .O(\DLX_IDinst_RegFile_28_22/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_366_352 (
    .IA(\DLX_IDinst_RegFile_28_22/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_28_22/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_425),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_366)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4251.INIT = 16'hE4FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4251 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR1(DLX_IDinst_RegFile_28_22),
    .ADR2(DLX_IDinst_RegFile_29_22),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_57),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_425)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4261.INIT = 16'hD8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4261 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR1(DLX_IDinst_RegFile_31_22),
    .ADR2(DLX_IDinst_RegFile_30_22),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_58),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_426)
  );
  X_BUF \DLX_IDinst_RegFile_28_22/COUTUSED  (
    .I(\DLX_IDinst_RegFile_28_22/CYMUXG ),
    .O(DLX_IDinst__n0623[22])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_367 (
    .IA(\DLX_IDinst_RegFile_28_22/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_366),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_426),
    .O(\DLX_IDinst_RegFile_28_22/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_28_22/CYINIT_353  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_365),
    .O(\DLX_IDinst_RegFile_28_22/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_28_14/LOGIC_ZERO_354  (
    .O(\DLX_IDinst_RegFile_28_14/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_238_355 (
    .IA(\DLX_IDinst_RegFile_28_14/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_28_14/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_297),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_238)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2971.INIT = 16'hFB3B;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2971 (
    .ADR0(DLX_IDinst_RegFile_28_14),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_57),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR3(DLX_IDinst_RegFile_29_14),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_297)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2981.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2981 (
    .ADR0(DLX_IDinst_RegFile_30_14),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_58),
    .ADR3(DLX_IDinst_RegFile_31_14),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_298)
  );
  X_BUF \DLX_IDinst_RegFile_28_14/COUTUSED  (
    .I(\DLX_IDinst_RegFile_28_14/CYMUXG ),
    .O(DLX_IDinst__n0623[14])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_239 (
    .IA(\DLX_IDinst_RegFile_28_14/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_238),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_298),
    .O(\DLX_IDinst_RegFile_28_14/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_28_14/CYINIT_356  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_237),
    .O(\DLX_IDinst_RegFile_28_14/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_28_23/LOGIC_ZERO_357  (
    .O(\DLX_IDinst_RegFile_28_23/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_382_358 (
    .IA(\DLX_IDinst_RegFile_28_23/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_28_23/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_441),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_382)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4411.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4411 (
    .ADR0(DLX_IDinst_RegFile_29_23),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_57),
    .ADR2(DLX_IDinst_RegFile_28_23),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_441)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4421.INIT = 16'hF5DD;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4421 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_58),
    .ADR1(DLX_IDinst_RegFile_30_23),
    .ADR2(DLX_IDinst_RegFile_31_23),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_442)
  );
  X_BUF \DLX_IDinst_RegFile_28_23/COUTUSED  (
    .I(\DLX_IDinst_RegFile_28_23/CYMUXG ),
    .O(DLX_IDinst__n0623[23])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_383 (
    .IA(\DLX_IDinst_RegFile_28_23/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_382),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_442),
    .O(\DLX_IDinst_RegFile_28_23/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_28_23/CYINIT_359  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_381),
    .O(\DLX_IDinst_RegFile_28_23/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_28_15/LOGIC_ZERO_360  (
    .O(\DLX_IDinst_RegFile_28_15/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_254_361 (
    .IA(\DLX_IDinst_RegFile_28_15/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_28_15/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_313),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_254)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3131.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3131 (
    .ADR0(DLX_IDinst_RegFile_29_15),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_57),
    .ADR2(DLX_IDinst_RegFile_28_15),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_313)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3141.INIT = 16'hACFF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3141 (
    .ADR0(DLX_IDinst_RegFile_31_15),
    .ADR1(DLX_IDinst_RegFile_30_15),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_58),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_314)
  );
  X_BUF \DLX_IDinst_RegFile_28_15/COUTUSED  (
    .I(\DLX_IDinst_RegFile_28_15/CYMUXG ),
    .O(DLX_IDinst__n0623[15])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_255 (
    .IA(\DLX_IDinst_RegFile_28_15/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_254),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_314),
    .O(\DLX_IDinst_RegFile_28_15/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_28_15/CYINIT_362  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_253),
    .O(\DLX_IDinst_RegFile_28_15/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_28_31/LOGIC_ZERO_363  (
    .O(\DLX_IDinst_RegFile_28_31/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_1022_364 (
    .IA(\DLX_IDinst_RegFile_28_31/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_28_31/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1097),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_1022)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10971.INIT = 16'hACFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10971 (
    .ADR0(DLX_IDinst_RegFile_29_31),
    .ADR1(DLX_IDinst_RegFile_28_31),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_585),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1097)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10981.INIT = 16'hFB3B;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10981 (
    .ADR0(DLX_IDinst_RegFile_30_31),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_586),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR3(DLX_IDinst_RegFile_31_31),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1098)
  );
  X_BUF \DLX_IDinst_RegFile_28_31/COUTUSED  (
    .I(\DLX_IDinst_RegFile_28_31/CYMUXG ),
    .O(DLX_IDinst__n0620[31])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_1023 (
    .IA(\DLX_IDinst_RegFile_28_31/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_1022),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1098),
    .O(\DLX_IDinst_RegFile_28_31/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_28_31/CYINIT_365  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_1021),
    .O(\DLX_IDinst_RegFile_28_31/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_28_24/LOGIC_ZERO_366  (
    .O(\DLX_IDinst_RegFile_28_24/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_398_367 (
    .IA(\DLX_IDinst_RegFile_28_24/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_28_24/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_457),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_398)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4571.INIT = 16'hF7D5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4571 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_57),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR2(DLX_IDinst_RegFile_29_24),
    .ADR3(DLX_IDinst_RegFile_28_24),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_457)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4581.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4581 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR1(DLX_IDinst_RegFile_30_24),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_58),
    .ADR3(DLX_IDinst_RegFile_31_24),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_458)
  );
  X_BUF \DLX_IDinst_RegFile_28_24/COUTUSED  (
    .I(\DLX_IDinst_RegFile_28_24/CYMUXG ),
    .O(DLX_IDinst__n0623[24])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_399 (
    .IA(\DLX_IDinst_RegFile_28_24/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_398),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_458),
    .O(\DLX_IDinst_RegFile_28_24/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_28_24/CYINIT_368  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_397),
    .O(\DLX_IDinst_RegFile_28_24/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_28_16/LOGIC_ZERO_369  (
    .O(\DLX_IDinst_RegFile_28_16/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_270_370 (
    .IA(\DLX_IDinst_RegFile_28_16/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_28_16/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_329),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_270)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3291.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3291 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_57),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR2(DLX_IDinst_RegFile_28_16),
    .ADR3(DLX_IDinst_RegFile_29_16),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_329)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3301.INIT = 16'hBF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3301 (
    .ADR0(DLX_IDinst_RegFile_31_16),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_58),
    .ADR3(DLX_IDinst_RegFile_30_16),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_330)
  );
  X_BUF \DLX_IDinst_RegFile_28_16/COUTUSED  (
    .I(\DLX_IDinst_RegFile_28_16/CYMUXG ),
    .O(DLX_IDinst__n0623[16])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_271 (
    .IA(\DLX_IDinst_RegFile_28_16/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_270),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_330),
    .O(\DLX_IDinst_RegFile_28_16/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_28_16/CYINIT_371  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_269),
    .O(\DLX_IDinst_RegFile_28_16/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_28_25/LOGIC_ZERO_372  (
    .O(\DLX_IDinst_RegFile_28_25/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_414_373 (
    .IA(\DLX_IDinst_RegFile_28_25/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_28_25/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_473),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_414)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4731.INIT = 16'hCFAF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4731 (
    .ADR0(DLX_IDinst_RegFile_28_25),
    .ADR1(DLX_IDinst_RegFile_29_25),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_57),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_473)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4741.INIT = 16'hACFF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4741 (
    .ADR0(DLX_IDinst_RegFile_31_25),
    .ADR1(DLX_IDinst_RegFile_30_25),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_58),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_474)
  );
  X_BUF \DLX_IDinst_RegFile_28_25/COUTUSED  (
    .I(\DLX_IDinst_RegFile_28_25/CYMUXG ),
    .O(DLX_IDinst__n0623[25])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_415 (
    .IA(\DLX_IDinst_RegFile_28_25/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_414),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_474),
    .O(\DLX_IDinst_RegFile_28_25/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_28_25/CYINIT_374  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_413),
    .O(\DLX_IDinst_RegFile_28_25/CYINIT )
  );
  defparam DLX_IDinst_RegFile_18_22_375.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_18_22_375 (
    .I(DLX_IDinst_WB_data_eff[22]),
    .CE(DLX_IDinst__n0586),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_18_22)
  );
  X_ZERO \DLX_IDinst_RegFile_28_17/LOGIC_ZERO_376  (
    .O(\DLX_IDinst_RegFile_28_17/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_286_377 (
    .IA(\DLX_IDinst_RegFile_28_17/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_28_17/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_345),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_286)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3451.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3451 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_57),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR2(DLX_IDinst_RegFile_28_17),
    .ADR3(DLX_IDinst_RegFile_29_17),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_345)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3461.INIT = 16'hBF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3461 (
    .ADR0(DLX_IDinst_RegFile_31_17),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_58),
    .ADR3(DLX_IDinst_RegFile_30_17),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_346)
  );
  X_BUF \DLX_IDinst_RegFile_28_17/COUTUSED  (
    .I(\DLX_IDinst_RegFile_28_17/CYMUXG ),
    .O(DLX_IDinst__n0623[17])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_287 (
    .IA(\DLX_IDinst_RegFile_28_17/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_286),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_346),
    .O(\DLX_IDinst_RegFile_28_17/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_28_17/CYINIT_378  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_285),
    .O(\DLX_IDinst_RegFile_28_17/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_28_26/LOGIC_ZERO_379  (
    .O(\DLX_IDinst_RegFile_28_26/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_430_380 (
    .IA(\DLX_IDinst_RegFile_28_26/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_28_26/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_489),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_430)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4891.INIT = 16'hB8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4891 (
    .ADR0(DLX_IDinst_RegFile_29_26),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR2(DLX_IDinst_RegFile_28_26),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_57),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_489)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4901.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4901 (
    .ADR0(DLX_IDinst_RegFile_30_26),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_58),
    .ADR2(DLX_IDinst_RegFile_31_26),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_490)
  );
  X_BUF \DLX_IDinst_RegFile_28_26/COUTUSED  (
    .I(\DLX_IDinst_RegFile_28_26/CYMUXG ),
    .O(DLX_IDinst__n0623[26])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_431 (
    .IA(\DLX_IDinst_RegFile_28_26/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_430),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_490),
    .O(\DLX_IDinst_RegFile_28_26/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_28_26/CYINIT_381  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_429),
    .O(\DLX_IDinst_RegFile_28_26/CYINIT )
  );
  defparam DLX_IDinst_RegFile_18_30_382.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_18_30_382 (
    .I(DLX_IDinst_WB_data_eff[30]),
    .CE(DLX_IDinst__n0586),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_18_30)
  );
  X_ZERO \DLX_IDinst_RegFile_28_18/LOGIC_ZERO_383  (
    .O(\DLX_IDinst_RegFile_28_18/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_302_384 (
    .IA(\DLX_IDinst_RegFile_28_18/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_28_18/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_361),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_302)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3611.INIT = 16'hFB3B;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3611 (
    .ADR0(DLX_IDinst_RegFile_28_18),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_57),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR3(DLX_IDinst_RegFile_29_18),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_361)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3621.INIT = 16'hF5DD;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3621 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_58),
    .ADR1(DLX_IDinst_RegFile_30_18),
    .ADR2(DLX_IDinst_RegFile_31_18),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_362)
  );
  X_BUF \DLX_IDinst_RegFile_28_18/COUTUSED  (
    .I(\DLX_IDinst_RegFile_28_18/CYMUXG ),
    .O(DLX_IDinst__n0623[18])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_303 (
    .IA(\DLX_IDinst_RegFile_28_18/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_302),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_362),
    .O(\DLX_IDinst_RegFile_28_18/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_28_18/CYINIT_385  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_301),
    .O(\DLX_IDinst_RegFile_28_18/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_29_10/LOGIC_ZERO_386  (
    .O(\DLX_IDinst_RegFile_29_10/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_686_387 (
    .IA(\DLX_IDinst_RegFile_29_10/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_29_10/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_761),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_686)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7611.INIT = 16'hDDF5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7611 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_585),
    .ADR1(DLX_IDinst_RegFile_29_10),
    .ADR2(DLX_IDinst_RegFile_28_10),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_761)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7621.INIT = 16'hB8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7621 (
    .ADR0(DLX_IDinst_RegFile_31_10),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR2(DLX_IDinst_RegFile_30_10),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_586),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_762)
  );
  X_BUF \DLX_IDinst_RegFile_29_10/COUTUSED  (
    .I(\DLX_IDinst_RegFile_29_10/CYMUXG ),
    .O(DLX_IDinst__n0620[10])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_687 (
    .IA(\DLX_IDinst_RegFile_29_10/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_686),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_762),
    .O(\DLX_IDinst_RegFile_29_10/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_29_10/CYINIT_388  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_685),
    .O(\DLX_IDinst_RegFile_29_10/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_28_27/LOGIC_ZERO_389  (
    .O(\DLX_IDinst_RegFile_28_27/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_446_390 (
    .IA(\DLX_IDinst_RegFile_28_27/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_28_27/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_505),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_446)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5051.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5051 (
    .ADR0(DLX_IDinst_RegFile_29_27),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_57),
    .ADR2(DLX_IDinst_RegFile_28_27),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_505)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5061.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5061 (
    .ADR0(DLX_IDinst_RegFile_31_27),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_58),
    .ADR2(DLX_IDinst_RegFile_30_27),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_506)
  );
  X_BUF \DLX_IDinst_RegFile_28_27/COUTUSED  (
    .I(\DLX_IDinst_RegFile_28_27/CYMUXG ),
    .O(DLX_IDinst__n0623[27])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_447 (
    .IA(\DLX_IDinst_RegFile_28_27/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_446),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_506),
    .O(\DLX_IDinst_RegFile_28_27/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_28_27/CYINIT_391  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_445),
    .O(\DLX_IDinst_RegFile_28_27/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_28_19/LOGIC_ZERO_392  (
    .O(\DLX_IDinst_RegFile_28_19/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_318_393 (
    .IA(\DLX_IDinst_RegFile_28_19/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_28_19/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_377),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_318)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3771.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3771 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR1(DLX_IDinst_RegFile_28_19),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_57),
    .ADR3(DLX_IDinst_RegFile_29_19),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_377)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3781.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3781 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_58),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR2(DLX_IDinst_RegFile_30_19),
    .ADR3(DLX_IDinst_RegFile_31_19),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_378)
  );
  X_BUF \DLX_IDinst_RegFile_28_19/COUTUSED  (
    .I(\DLX_IDinst_RegFile_28_19/CYMUXG ),
    .O(DLX_IDinst__n0623[19])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_319 (
    .IA(\DLX_IDinst_RegFile_28_19/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_318),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_378),
    .O(\DLX_IDinst_RegFile_28_19/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_28_19/CYINIT_394  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_317),
    .O(\DLX_IDinst_RegFile_28_19/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_29_11/LOGIC_ZERO_395  (
    .O(\DLX_IDinst_RegFile_29_11/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_702_396 (
    .IA(\DLX_IDinst_RegFile_29_11/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_29_11/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_777),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_702)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7771.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7771 (
    .ADR0(DLX_IDinst_RegFile_28_11),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_585),
    .ADR2(DLX_IDinst_RegFile_29_11),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_777)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7781.INIT = 16'hE4FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7781 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR1(DLX_IDinst_RegFile_30_11),
    .ADR2(DLX_IDinst_RegFile_31_11),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_586),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_778)
  );
  X_BUF \DLX_IDinst_RegFile_29_11/COUTUSED  (
    .I(\DLX_IDinst_RegFile_29_11/CYMUXG ),
    .O(DLX_IDinst__n0620[11])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_703 (
    .IA(\DLX_IDinst_RegFile_29_11/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_702),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_778),
    .O(\DLX_IDinst_RegFile_29_11/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_29_11/CYINIT_397  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_701),
    .O(\DLX_IDinst_RegFile_29_11/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_28_28/LOGIC_ZERO_398  (
    .O(\DLX_IDinst_RegFile_28_28/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_974_399 (
    .IA(\DLX_IDinst_RegFile_28_28/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_28_28/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1049),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_974)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10491.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10491 (
    .ADR0(DLX_IDinst_RegFile_28_28),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_585),
    .ADR2(DLX_IDinst_RegFile_29_28),
    .ADR3(DLX_IDinst_jtarget[21]),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1049)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10501.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10501 (
    .ADR0(DLX_IDinst_RegFile_30_28),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_586),
    .ADR2(DLX_IDinst_RegFile_31_28),
    .ADR3(DLX_IDinst_jtarget[21]),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1050)
  );
  X_BUF \DLX_IDinst_RegFile_28_28/COUTUSED  (
    .I(\DLX_IDinst_RegFile_28_28/CYMUXG ),
    .O(DLX_IDinst__n0620[28])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_975 (
    .IA(\DLX_IDinst_RegFile_28_28/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_974),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1050),
    .O(\DLX_IDinst_RegFile_28_28/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_28_28/CYINIT_400  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_973),
    .O(\DLX_IDinst_RegFile_28_28/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_29_20/LOGIC_ZERO_401  (
    .O(\DLX_IDinst_RegFile_29_20/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_846_402 (
    .IA(\DLX_IDinst_RegFile_29_20/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_29_20/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_921),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_846)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9211.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9211 (
    .ADR0(DLX_IDinst_RegFile_28_20),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_585),
    .ADR2(DLX_IDinst_RegFile_29_20),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_921)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9221.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9221 (
    .ADR0(DLX_IDinst_RegFile_30_20),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_586),
    .ADR3(DLX_IDinst_RegFile_31_20),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_922)
  );
  X_BUF \DLX_IDinst_RegFile_29_20/COUTUSED  (
    .I(\DLX_IDinst_RegFile_29_20/CYMUXG ),
    .O(DLX_IDinst__n0620[20])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_847 (
    .IA(\DLX_IDinst_RegFile_29_20/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_846),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_922),
    .O(\DLX_IDinst_RegFile_29_20/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_29_20/CYINIT_403  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_845),
    .O(\DLX_IDinst_RegFile_29_20/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_29_12/LOGIC_ZERO_404  (
    .O(\DLX_IDinst_RegFile_29_12/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_718_405 (
    .IA(\DLX_IDinst_RegFile_29_12/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_29_12/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_793),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_718)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7931.INIT = 16'hF7D5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7931 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_585),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR2(DLX_IDinst_RegFile_29_12),
    .ADR3(DLX_IDinst_RegFile_28_12),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_793)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7941.INIT = 16'hD8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7941 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR1(DLX_IDinst_RegFile_31_12),
    .ADR2(DLX_IDinst_RegFile_30_12),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_586),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_794)
  );
  X_BUF \DLX_IDinst_RegFile_29_12/COUTUSED  (
    .I(\DLX_IDinst_RegFile_29_12/CYMUXG ),
    .O(DLX_IDinst__n0620[12])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_719 (
    .IA(\DLX_IDinst_RegFile_29_12/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_718),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_794),
    .O(\DLX_IDinst_RegFile_29_12/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_29_12/CYINIT_406  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_717),
    .O(\DLX_IDinst_RegFile_29_12/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_28_29/LOGIC_ZERO_407  (
    .O(\DLX_IDinst_RegFile_28_29/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_990_408 (
    .IA(\DLX_IDinst_RegFile_28_29/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_28_29/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1065),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_990)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10651.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10651 (
    .ADR0(DLX_IDinst_RegFile_28_29),
    .ADR1(DLX_IDinst_RegFile_29_29),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_585),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1065)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10661.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10661 (
    .ADR0(DLX_IDinst_RegFile_30_29),
    .ADR1(DLX_IDinst_RegFile_31_29),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_586),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1066)
  );
  X_BUF \DLX_IDinst_RegFile_28_29/COUTUSED  (
    .I(\DLX_IDinst_RegFile_28_29/CYMUXG ),
    .O(DLX_IDinst__n0620[29])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_991 (
    .IA(\DLX_IDinst_RegFile_28_29/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_990),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1066),
    .O(\DLX_IDinst_RegFile_28_29/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_28_29/CYINIT_409  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_989),
    .O(\DLX_IDinst_RegFile_28_29/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_29_21/LOGIC_ZERO_410  (
    .O(\DLX_IDinst_RegFile_29_21/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_862_411 (
    .IA(\DLX_IDinst_RegFile_29_21/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_29_21/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_937),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_862)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9371.INIT = 16'hD8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9371 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR1(DLX_IDinst_RegFile_29_21),
    .ADR2(DLX_IDinst_RegFile_28_21),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_585),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_937)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9381.INIT = 16'hB8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9381 (
    .ADR0(DLX_IDinst_RegFile_31_21),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR2(DLX_IDinst_RegFile_30_21),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_586),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_938)
  );
  X_BUF \DLX_IDinst_RegFile_29_21/COUTUSED  (
    .I(\DLX_IDinst_RegFile_29_21/CYMUXG ),
    .O(DLX_IDinst__n0620[21])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_863 (
    .IA(\DLX_IDinst_RegFile_29_21/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_862),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_938),
    .O(\DLX_IDinst_RegFile_29_21/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_29_21/CYINIT_412  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_861),
    .O(\DLX_IDinst_RegFile_29_21/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_29_13/LOGIC_ZERO_413  (
    .O(\DLX_IDinst_RegFile_29_13/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_734_414 (
    .IA(\DLX_IDinst_RegFile_29_13/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_29_13/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_809),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_734)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8091.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8091 (
    .ADR0(DLX_IDinst_RegFile_28_13),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_585),
    .ADR3(DLX_IDinst_RegFile_29_13),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_809)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8101.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8101 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_586),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR2(DLX_IDinst_RegFile_30_13),
    .ADR3(DLX_IDinst_RegFile_31_13),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_810)
  );
  X_BUF \DLX_IDinst_RegFile_29_13/COUTUSED  (
    .I(\DLX_IDinst_RegFile_29_13/CYMUXG ),
    .O(DLX_IDinst__n0620[13])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_735 (
    .IA(\DLX_IDinst_RegFile_29_13/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_734),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_810),
    .O(\DLX_IDinst_RegFile_29_13/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_29_13/CYINIT_415  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_733),
    .O(\DLX_IDinst_RegFile_29_13/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_29_30/LOGIC_ZERO_416  (
    .O(\DLX_IDinst_RegFile_29_30/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_494_417 (
    .IA(\DLX_IDinst_RegFile_29_30/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_29_30/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_553),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_494)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5531.INIT = 16'hCFAF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5531 (
    .ADR0(DLX_IDinst_RegFile_28_30),
    .ADR1(DLX_IDinst_RegFile_29_30),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_57),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_553)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5541.INIT = 16'hCFAF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5541 (
    .ADR0(DLX_IDinst_RegFile_30_30),
    .ADR1(DLX_IDinst_RegFile_31_30),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_58),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_554)
  );
  X_BUF \DLX_IDinst_RegFile_29_30/COUTUSED  (
    .I(\DLX_IDinst_RegFile_29_30/CYMUXG ),
    .O(DLX_IDinst__n0623[30])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_495 (
    .IA(\DLX_IDinst_RegFile_29_30/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_494),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_554),
    .O(\DLX_IDinst_RegFile_29_30/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_29_30/CYINIT_418  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_493),
    .O(\DLX_IDinst_RegFile_29_30/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_29_22/LOGIC_ZERO_419  (
    .O(\DLX_IDinst_RegFile_29_22/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_878_420 (
    .IA(\DLX_IDinst_RegFile_29_22/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_29_22/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_953),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_878)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9531.INIT = 16'hB8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9531 (
    .ADR0(DLX_IDinst_RegFile_29_22),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR2(DLX_IDinst_RegFile_28_22),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_585),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_953)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9541.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9541 (
    .ADR0(DLX_IDinst_RegFile_30_22),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_586),
    .ADR3(DLX_IDinst_RegFile_31_22),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_954)
  );
  X_BUF \DLX_IDinst_RegFile_29_22/COUTUSED  (
    .I(\DLX_IDinst_RegFile_29_22/CYMUXG ),
    .O(DLX_IDinst__n0620[22])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_879 (
    .IA(\DLX_IDinst_RegFile_29_22/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_878),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_954),
    .O(\DLX_IDinst_RegFile_29_22/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_29_22/CYINIT_421  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_877),
    .O(\DLX_IDinst_RegFile_29_22/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_29_14/LOGIC_ZERO_422  (
    .O(\DLX_IDinst_RegFile_29_14/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_750_423 (
    .IA(\DLX_IDinst_RegFile_29_14/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_29_14/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_825),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_750)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8251.INIT = 16'hF7D5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8251 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_585),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR2(DLX_IDinst_RegFile_29_14),
    .ADR3(DLX_IDinst_RegFile_28_14),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_825)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8261.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8261 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR1(DLX_IDinst_RegFile_30_14),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_586),
    .ADR3(DLX_IDinst_RegFile_31_14),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_826)
  );
  X_BUF \DLX_IDinst_RegFile_29_14/COUTUSED  (
    .I(\DLX_IDinst_RegFile_29_14/CYMUXG ),
    .O(DLX_IDinst__n0620[14])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_751 (
    .IA(\DLX_IDinst_RegFile_29_14/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_750),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_826),
    .O(\DLX_IDinst_RegFile_29_14/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_29_14/CYINIT_424  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_749),
    .O(\DLX_IDinst_RegFile_29_14/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_29_23/LOGIC_ZERO_425  (
    .O(\DLX_IDinst_RegFile_29_23/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_894_426 (
    .IA(\DLX_IDinst_RegFile_29_23/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_29_23/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_969),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_894)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9691.INIT = 16'hFB3B;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9691 (
    .ADR0(DLX_IDinst_RegFile_28_23),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_585),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR3(DLX_IDinst_RegFile_29_23),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_969)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9701.INIT = 16'hBF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9701 (
    .ADR0(DLX_IDinst_RegFile_31_23),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_586),
    .ADR3(DLX_IDinst_RegFile_30_23),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_970)
  );
  X_BUF \DLX_IDinst_RegFile_29_23/COUTUSED  (
    .I(\DLX_IDinst_RegFile_29_23/CYMUXG ),
    .O(DLX_IDinst__n0620[23])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_895 (
    .IA(\DLX_IDinst_RegFile_29_23/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_894),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_970),
    .O(\DLX_IDinst_RegFile_29_23/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_29_23/CYINIT_427  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_893),
    .O(\DLX_IDinst_RegFile_29_23/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_29_15/LOGIC_ZERO_428  (
    .O(\DLX_IDinst_RegFile_29_15/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_766_429 (
    .IA(\DLX_IDinst_RegFile_29_15/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_29_15/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_841),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_766)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8411.INIT = 16'hDDF5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8411 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_585),
    .ADR1(DLX_IDinst_RegFile_29_15),
    .ADR2(DLX_IDinst_RegFile_28_15),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_841)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8421.INIT = 16'hDDF5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8421 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_586),
    .ADR1(DLX_IDinst_RegFile_31_15),
    .ADR2(DLX_IDinst_RegFile_30_15),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_842)
  );
  X_BUF \DLX_IDinst_RegFile_29_15/COUTUSED  (
    .I(\DLX_IDinst_RegFile_29_15/CYMUXG ),
    .O(DLX_IDinst__n0620[15])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_767 (
    .IA(\DLX_IDinst_RegFile_29_15/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_766),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_842),
    .O(\DLX_IDinst_RegFile_29_15/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_29_15/CYINIT_430  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_765),
    .O(\DLX_IDinst_RegFile_29_15/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_29_31/LOGIC_ZERO_431  (
    .O(\DLX_IDinst_RegFile_29_31/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_510_432 (
    .IA(\DLX_IDinst_RegFile_29_31/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_29_31/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_569),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_510)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5691.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5691 (
    .ADR0(DLX_IDinst_RegFile_28_31),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_57),
    .ADR2(DLX_IDinst_RegFile_29_31),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_569)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5701.INIT = 16'hF5DD;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5701 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_58),
    .ADR1(DLX_IDinst_RegFile_30_31),
    .ADR2(DLX_IDinst_RegFile_31_31),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_570)
  );
  X_BUF \DLX_IDinst_RegFile_29_31/COUTUSED  (
    .I(\DLX_IDinst_RegFile_29_31/CYMUXG ),
    .O(DLX_IDinst__n0623[31])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_511 (
    .IA(\DLX_IDinst_RegFile_29_31/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_510),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_570),
    .O(\DLX_IDinst_RegFile_29_31/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_29_31/CYINIT_433  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_509),
    .O(\DLX_IDinst_RegFile_29_31/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_29_24/LOGIC_ZERO_434  (
    .O(\DLX_IDinst_RegFile_29_24/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_910_435 (
    .IA(\DLX_IDinst_RegFile_29_24/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_29_24/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_985),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_910)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9851.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9851 (
    .ADR0(DLX_IDinst_RegFile_29_24),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_585),
    .ADR2(DLX_IDinst_RegFile_28_24),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_985)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9861.INIT = 16'hB8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9861 (
    .ADR0(DLX_IDinst_RegFile_31_24),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR2(DLX_IDinst_RegFile_30_24),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_586),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_986)
  );
  X_BUF \DLX_IDinst_RegFile_29_24/COUTUSED  (
    .I(\DLX_IDinst_RegFile_29_24/CYMUXG ),
    .O(DLX_IDinst__n0620[24])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_911 (
    .IA(\DLX_IDinst_RegFile_29_24/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_910),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_986),
    .O(\DLX_IDinst_RegFile_29_24/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_29_24/CYINIT_436  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_909),
    .O(\DLX_IDinst_RegFile_29_24/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_29_16/LOGIC_ZERO_437  (
    .O(\DLX_IDinst_RegFile_29_16/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_782_438 (
    .IA(\DLX_IDinst_RegFile_29_16/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_29_16/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_857),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_782)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8571.INIT = 16'hAFCF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8571 (
    .ADR0(DLX_IDinst_RegFile_29_16),
    .ADR1(DLX_IDinst_RegFile_28_16),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_585),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_857)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8581.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8581 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR1(DLX_IDinst_RegFile_30_16),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_586),
    .ADR3(DLX_IDinst_RegFile_31_16),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_858)
  );
  X_BUF \DLX_IDinst_RegFile_29_16/COUTUSED  (
    .I(\DLX_IDinst_RegFile_29_16/CYMUXG ),
    .O(DLX_IDinst__n0620[16])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_783 (
    .IA(\DLX_IDinst_RegFile_29_16/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_782),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_858),
    .O(\DLX_IDinst_RegFile_29_16/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_29_16/CYINIT_439  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_781),
    .O(\DLX_IDinst_RegFile_29_16/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_29_25/LOGIC_ZERO_440  (
    .O(\DLX_IDinst_RegFile_29_25/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_926_441 (
    .IA(\DLX_IDinst_RegFile_29_25/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_29_25/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1001),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_926)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10011.INIT = 16'hDF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10011 (
    .ADR0(DLX_IDinst_jtarget[21]),
    .ADR1(DLX_IDinst_RegFile_29_25),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_585),
    .ADR3(DLX_IDinst_RegFile_28_25),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1001)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10021.INIT = 16'hBFB3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10021 (
    .ADR0(DLX_IDinst_RegFile_31_25),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_586),
    .ADR2(DLX_IDinst_jtarget[21]),
    .ADR3(DLX_IDinst_RegFile_30_25),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1002)
  );
  X_BUF \DLX_IDinst_RegFile_29_25/COUTUSED  (
    .I(\DLX_IDinst_RegFile_29_25/CYMUXG ),
    .O(DLX_IDinst__n0620[25])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_927 (
    .IA(\DLX_IDinst_RegFile_29_25/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_926),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1002),
    .O(\DLX_IDinst_RegFile_29_25/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_29_25/CYINIT_442  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_925),
    .O(\DLX_IDinst_RegFile_29_25/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_29_17/LOGIC_ZERO_443  (
    .O(\DLX_IDinst_RegFile_29_17/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_798_444 (
    .IA(\DLX_IDinst_RegFile_29_17/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_29_17/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_873),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_798)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8731.INIT = 16'hAFCF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8731 (
    .ADR0(DLX_IDinst_RegFile_29_17),
    .ADR1(DLX_IDinst_RegFile_28_17),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_585),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_873)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8741.INIT = 16'hFB3B;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8741 (
    .ADR0(DLX_IDinst_RegFile_30_17),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_586),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR3(DLX_IDinst_RegFile_31_17),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_874)
  );
  X_BUF \DLX_IDinst_RegFile_29_17/COUTUSED  (
    .I(\DLX_IDinst_RegFile_29_17/CYMUXG ),
    .O(DLX_IDinst__n0620[17])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_799 (
    .IA(\DLX_IDinst_RegFile_29_17/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_798),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_874),
    .O(\DLX_IDinst_RegFile_29_17/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_29_17/CYINIT_445  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_797),
    .O(\DLX_IDinst_RegFile_29_17/CYINIT )
  );
  defparam DLX_IDinst_RegFile_18_14_446.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_18_14_446 (
    .I(DLX_IDinst_WB_data_eff[14]),
    .CE(DLX_IDinst__n0586),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_18_14)
  );
  X_ZERO \DLX_IDinst_RegFile_29_26/LOGIC_ZERO_447  (
    .O(\DLX_IDinst_RegFile_29_26/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_942_448 (
    .IA(\DLX_IDinst_RegFile_29_26/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_29_26/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1017),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_942)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10171.INIT = 16'hBFB3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10171 (
    .ADR0(DLX_IDinst_RegFile_29_26),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_585),
    .ADR2(DLX_IDinst_jtarget[21]),
    .ADR3(DLX_IDinst_RegFile_28_26),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1017)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10181.INIT = 16'hDFD5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10181 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_586),
    .ADR1(DLX_IDinst_RegFile_31_26),
    .ADR2(DLX_IDinst_jtarget[21]),
    .ADR3(DLX_IDinst_RegFile_30_26),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1018)
  );
  X_BUF \DLX_IDinst_RegFile_29_26/COUTUSED  (
    .I(\DLX_IDinst_RegFile_29_26/CYMUXG ),
    .O(DLX_IDinst__n0620[26])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_943 (
    .IA(\DLX_IDinst_RegFile_29_26/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_942),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1018),
    .O(\DLX_IDinst_RegFile_29_26/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_29_26/CYINIT_449  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_941),
    .O(\DLX_IDinst_RegFile_29_26/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_29_18/LOGIC_ZERO_450  (
    .O(\DLX_IDinst_RegFile_29_18/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_814_451 (
    .IA(\DLX_IDinst_RegFile_29_18/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_29_18/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_889),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_814)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8891.INIT = 16'hBFB3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8891 (
    .ADR0(DLX_IDinst_RegFile_29_18),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_585),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR3(DLX_IDinst_RegFile_28_18),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_889)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8901.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8901 (
    .ADR0(DLX_IDinst_RegFile_30_18),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_586),
    .ADR3(DLX_IDinst_RegFile_31_18),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_890)
  );
  X_BUF \DLX_IDinst_RegFile_29_18/COUTUSED  (
    .I(\DLX_IDinst_RegFile_29_18/CYMUXG ),
    .O(DLX_IDinst__n0620[18])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_815 (
    .IA(\DLX_IDinst_RegFile_29_18/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_814),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_890),
    .O(\DLX_IDinst_RegFile_29_18/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_29_18/CYINIT_452  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_813),
    .O(\DLX_IDinst_RegFile_29_18/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_29_27/LOGIC_ZERO_453  (
    .O(\DLX_IDinst_RegFile_29_27/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_958_454 (
    .IA(\DLX_IDinst_RegFile_29_27/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_29_27/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1033),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_958)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10331.INIT = 16'hAFCF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10331 (
    .ADR0(DLX_IDinst_RegFile_29_27),
    .ADR1(DLX_IDinst_RegFile_28_27),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_585),
    .ADR3(DLX_IDinst_jtarget[21]),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1033)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10341.INIT = 16'hFB3B;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10341 (
    .ADR0(DLX_IDinst_RegFile_30_27),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_586),
    .ADR2(DLX_IDinst_jtarget[21]),
    .ADR3(DLX_IDinst_RegFile_31_27),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1034)
  );
  X_BUF \DLX_IDinst_RegFile_29_27/COUTUSED  (
    .I(\DLX_IDinst_RegFile_29_27/CYMUXG ),
    .O(DLX_IDinst__n0620[27])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_959 (
    .IA(\DLX_IDinst_RegFile_29_27/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_958),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1034),
    .O(\DLX_IDinst_RegFile_29_27/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_29_27/CYINIT_455  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_957),
    .O(\DLX_IDinst_RegFile_29_27/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_29_19/LOGIC_ZERO_456  (
    .O(\DLX_IDinst_RegFile_29_19/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_830_457 (
    .IA(\DLX_IDinst_RegFile_29_19/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_29_19/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_905),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_830)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9051.INIT = 16'hFD5D;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9051 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_585),
    .ADR1(DLX_IDinst_RegFile_28_19),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR3(DLX_IDinst_RegFile_29_19),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_905)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9061.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9061 (
    .ADR0(DLX_IDinst_RegFile_31_19),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_586),
    .ADR2(DLX_IDinst_RegFile_30_19),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_906)
  );
  X_BUF \DLX_IDinst_RegFile_29_19/COUTUSED  (
    .I(\DLX_IDinst_RegFile_29_19/CYMUXG ),
    .O(DLX_IDinst__n0620[19])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_831 (
    .IA(\DLX_IDinst_RegFile_29_19/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_830),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_906),
    .O(\DLX_IDinst_RegFile_29_19/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_29_19/CYINIT_458  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_829),
    .O(\DLX_IDinst_RegFile_29_19/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_29_28/LOGIC_ZERO_459  (
    .O(\DLX_IDinst_RegFile_29_28/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_462_460 (
    .IA(\DLX_IDinst_RegFile_29_28/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_29_28/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_521),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_462)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5211.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5211 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_57),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR2(DLX_IDinst_RegFile_28_28),
    .ADR3(DLX_IDinst_RegFile_29_28),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_521)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5221.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5221 (
    .ADR0(DLX_IDinst_RegFile_30_28),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_58),
    .ADR3(DLX_IDinst_RegFile_31_28),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_522)
  );
  X_BUF \DLX_IDinst_RegFile_29_28/COUTUSED  (
    .I(\DLX_IDinst_RegFile_29_28/CYMUXG ),
    .O(DLX_IDinst__n0623[28])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_463 (
    .IA(\DLX_IDinst_RegFile_29_28/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_462),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_522),
    .O(\DLX_IDinst_RegFile_29_28/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_29_28/CYINIT_461  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_461),
    .O(\DLX_IDinst_RegFile_29_28/CYINIT )
  );
  defparam DLX_EXinst__n01271.INIT = 16'h0010;
  X_LUT4 DLX_EXinst__n01271 (
    .ADR0(\DLX_IDinst_Imm[3] ),
    .ADR1(\DLX_IDinst_Imm[2] ),
    .ADR2(DLX_IDinst_IR_function_field[5]),
    .ADR3(\DLX_IDinst_Imm[4] ),
    .O(\DLX_EXinst__n0127/FROM )
  );
  defparam DLX_EXinst__n000521.INIT = 16'h0001;
  X_LUT4 DLX_EXinst__n000521 (
    .ADR0(\DLX_IDinst_Imm[1] ),
    .ADR1(\DLX_IDinst_Imm[3] ),
    .ADR2(\DLX_IDinst_Imm[2] ),
    .ADR3(\DLX_IDinst_Imm[4] ),
    .O(\DLX_EXinst__n0127/GROM )
  );
  X_BUF \DLX_EXinst__n0127/XUSED  (
    .I(\DLX_EXinst__n0127/FROM ),
    .O(DLX_EXinst__n0127)
  );
  X_BUF \DLX_EXinst__n0127/YUSED  (
    .I(\DLX_EXinst__n0127/GROM ),
    .O(CHOICE2089)
  );
  X_ZERO \DLX_IDinst_RegFile_29_29/LOGIC_ZERO_462  (
    .O(\DLX_IDinst_RegFile_29_29/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_478_463 (
    .IA(\DLX_IDinst_RegFile_29_29/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_29_29/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_537),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_478)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5371.INIT = 16'hF5DD;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5371 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_57),
    .ADR1(DLX_IDinst_RegFile_28_29),
    .ADR2(DLX_IDinst_RegFile_29_29),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_537)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5381.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5381 (
    .ADR0(DLX_IDinst_RegFile_30_29),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_58),
    .ADR3(DLX_IDinst_RegFile_31_29),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_538)
  );
  X_BUF \DLX_IDinst_RegFile_29_29/COUTUSED  (
    .I(\DLX_IDinst_RegFile_29_29/CYMUXG ),
    .O(DLX_IDinst__n0623[29])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_479 (
    .IA(\DLX_IDinst_RegFile_29_29/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_478),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_538),
    .O(\DLX_IDinst_RegFile_29_29/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_29_29/CYINIT_464  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_477),
    .O(\DLX_IDinst_RegFile_29_29/CYINIT )
  );
  defparam DLX_EXinst__n001410.INIT = 16'hFFFD;
  X_LUT4 DLX_EXinst__n001410 (
    .ADR0(DLX_IDinst_IR_function_field[5]),
    .ADR1(\DLX_IDinst_Imm[1] ),
    .ADR2(DLX_IDinst_IR_opcode_field[0]),
    .ADR3(\DLX_IDinst_Imm[4] ),
    .O(\CHOICE3008/FROM )
  );
  defparam DLX_EXinst__n001420.INIT = 16'h00FE;
  X_LUT4 DLX_EXinst__n001420 (
    .ADR0(CHOICE3008),
    .ADR1(\DLX_IDinst_Imm[3] ),
    .ADR2(\DLX_IDinst_Imm[2] ),
    .ADR3(DLX_IDinst_IR_opcode_field[3]),
    .O(\CHOICE3008/GROM )
  );
  X_BUF \CHOICE3008/XUSED  (
    .I(\CHOICE3008/FROM ),
    .O(CHOICE3008)
  );
  X_BUF \CHOICE3008/YUSED  (
    .I(\CHOICE3008/GROM ),
    .O(CHOICE3010)
  );
  defparam DLX_EXinst__n003212.INIT = 16'hFFFE;
  X_LUT4 DLX_EXinst__n003212 (
    .ADR0(DLX_IDinst_reg_out_B[26]),
    .ADR1(DLX_IDinst_reg_out_B[27]),
    .ADR2(DLX_IDinst_reg_out_B[24]),
    .ADR3(DLX_IDinst_reg_out_B[25]),
    .O(\CHOICE3575/FROM )
  );
  defparam DLX_EXinst__n003215.INIT = 16'hFFFE;
  X_LUT4 DLX_EXinst__n003215 (
    .ADR0(DLX_IDinst_reg_out_B[29]),
    .ADR1(DLX_IDinst_reg_out_B[28]),
    .ADR2(DLX_IDinst_reg_out_B[30]),
    .ADR3(CHOICE3575),
    .O(\CHOICE3575/GROM )
  );
  X_BUF \CHOICE3575/XUSED  (
    .I(\CHOICE3575/FROM ),
    .O(CHOICE3575)
  );
  X_BUF \CHOICE3575/YUSED  (
    .I(\CHOICE3575/GROM ),
    .O(CHOICE3576)
  );
  defparam DLX_EXinst_Ker76159116.INIT = 16'h0001;
  X_LUT4 DLX_EXinst_Ker76159116 (
    .ADR0(\DLX_IDinst_Imm[12] ),
    .ADR1(\DLX_IDinst_Imm[11] ),
    .ADR2(\DLX_IDinst_Imm[13] ),
    .ADR3(\DLX_IDinst_Imm[14] ),
    .O(\CHOICE3442/FROM )
  );
  defparam DLX_EXinst__n003150.INIT = 16'hFFFE;
  X_LUT4 DLX_EXinst__n003150 (
    .ADR0(\DLX_IDinst_Imm[15] ),
    .ADR1(\DLX_IDinst_Imm[14] ),
    .ADR2(\DLX_IDinst_Imm[12] ),
    .ADR3(\DLX_IDinst_Imm[13] ),
    .O(\CHOICE3442/GROM )
  );
  X_BUF \CHOICE3442/XUSED  (
    .I(\CHOICE3442/FROM ),
    .O(CHOICE3442)
  );
  X_BUF \CHOICE3442/YUSED  (
    .I(\CHOICE3442/GROM ),
    .O(CHOICE3272)
  );
  defparam DLX_EXinst_Ker76181120.INIT = 16'h0001;
  X_LUT4 DLX_EXinst_Ker76181120 (
    .ADR0(DLX_IDinst_reg_out_B[12]),
    .ADR1(DLX_IDinst_reg_out_B[11]),
    .ADR2(DLX_IDinst_reg_out_B[10]),
    .ADR3(DLX_IDinst_reg_out_B[13]),
    .O(\DLX_IFinst_IR_previous<26>/FROM )
  );
  defparam DLX_EXinst__n003250.INIT = 16'hFFFE;
  X_LUT4 DLX_EXinst__n003250 (
    .ADR0(DLX_IDinst_reg_out_B[15]),
    .ADR1(DLX_IDinst_reg_out_B[12]),
    .ADR2(DLX_IDinst_reg_out_B[13]),
    .ADR3(DLX_IDinst_reg_out_B[14]),
    .O(\DLX_IFinst_IR_previous<26>/GROM )
  );
  X_BUF \DLX_IFinst_IR_previous<26>/XUSED  (
    .I(\DLX_IFinst_IR_previous<26>/FROM ),
    .O(CHOICE3639)
  );
  X_BUF \DLX_IFinst_IR_previous<26>/YUSED  (
    .I(\DLX_IFinst_IR_previous<26>/GROM ),
    .O(CHOICE3587)
  );
  defparam DLX_IDinst_RegFile_1_28_465.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_1_28_465 (
    .I(DLX_IDinst_WB_data_eff[28]),
    .CE(DLX_IDinst__n0552),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_1_28)
  );
  defparam DLX_EXinst__n003155.INIT = 16'hFFFE;
  X_LUT4 DLX_EXinst__n003155 (
    .ADR0(\DLX_IDinst_Imm[8] ),
    .ADR1(\DLX_IDinst_Imm[9] ),
    .ADR2(\DLX_IDinst_Imm[10] ),
    .ADR3(\DLX_IDinst_Imm[11] ),
    .O(\DLX_IDinst_RegFile_1_28/FROM )
  );
  defparam DLX_EXinst__n003174_SW0.INIT = 16'hFFFA;
  X_LUT4 DLX_EXinst__n003174_SW0 (
    .ADR0(\DLX_IDinst_Imm[31] ),
    .ADR1(VCC),
    .ADR2(CHOICE3272),
    .ADR3(CHOICE3275),
    .O(\DLX_IDinst_RegFile_1_28/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_1_28/XUSED  (
    .I(\DLX_IDinst_RegFile_1_28/FROM ),
    .O(CHOICE3275)
  );
  X_BUF \DLX_IDinst_RegFile_1_28/YUSED  (
    .I(\DLX_IDinst_RegFile_1_28/GROM ),
    .O(N163162)
  );
  defparam DLX_EXinst_reg_out_B_EX_4.INIT = 1'b0;
  X_SFF DLX_EXinst_reg_out_B_EX_4 (
    .I(DLX_IDinst_reg_out_B[4]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_reg_out_B_EX[4])
  );
  defparam DLX_EXinst__n003174.INIT = 16'hFFFE;
  X_LUT4 DLX_EXinst__n003174 (
    .ADR0(\DLX_IDinst_Imm[7] ),
    .ADR1(\DLX_IDinst_Imm[5] ),
    .ADR2(N163162),
    .ADR3(\DLX_IDinst_Imm[6] ),
    .O(\DLX_EXinst_reg_out_B_EX<4>/FROM )
  );
  defparam DLX_EXinst_Ker764391.INIT = 16'h0040;
  X_LUT4 DLX_EXinst_Ker764391 (
    .ADR0(DLX_IDinst_IR_opcode_field[0]),
    .ADR1(DLX_EXinst_N76041),
    .ADR2(DLX_IDinst_IR_opcode_field[1]),
    .ADR3(N146478),
    .O(\DLX_EXinst_reg_out_B_EX<4>/GROM )
  );
  X_BUF \DLX_EXinst_reg_out_B_EX<4>/XUSED  (
    .I(\DLX_EXinst_reg_out_B_EX<4>/FROM ),
    .O(N146478)
  );
  X_BUF \DLX_EXinst_reg_out_B_EX<4>/YUSED  (
    .I(\DLX_EXinst_reg_out_B_EX<4>/GROM ),
    .O(DLX_EXinst_N76441)
  );
  defparam DLX_IDinst_RegFile_1_29_466.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_1_29_466 (
    .I(DLX_IDinst_WB_data_eff[29]),
    .CE(DLX_IDinst__n0552),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_1_29)
  );
  defparam DLX_EXinst_Ker7618196.INIT = 16'h0001;
  X_LUT4 DLX_EXinst_Ker7618196 (
    .ADR0(DLX_IDinst_reg_out_B[14]),
    .ADR1(DLX_IDinst_reg_out_B[15]),
    .ADR2(DLX_IDinst_reg_out_B[17]),
    .ADR3(DLX_IDinst_reg_out_B[16]),
    .O(\DLX_IDinst_RegFile_1_29/FROM )
  );
  defparam DLX_EXinst__n003238.INIT = 16'hFFFE;
  X_LUT4 DLX_EXinst__n003238 (
    .ADR0(DLX_IDinst_reg_out_B[18]),
    .ADR1(DLX_IDinst_reg_out_B[17]),
    .ADR2(DLX_IDinst_reg_out_B[19]),
    .ADR3(DLX_IDinst_reg_out_B[16]),
    .O(\DLX_IDinst_RegFile_1_29/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_1_29/XUSED  (
    .I(\DLX_IDinst_RegFile_1_29/FROM ),
    .O(CHOICE3631)
  );
  X_BUF \DLX_IDinst_RegFile_1_29/YUSED  (
    .I(\DLX_IDinst_RegFile_1_29/GROM ),
    .O(CHOICE3583)
  );
  defparam DLX_EXinst__n003255.INIT = 16'hFFFE;
  X_LUT4 DLX_EXinst__n003255 (
    .ADR0(DLX_IDinst_reg_out_B[9]),
    .ADR1(DLX_IDinst_reg_out_B[8]),
    .ADR2(DLX_IDinst_reg_out_B[10]),
    .ADR3(DLX_IDinst_reg_out_B[11]),
    .O(\CHOICE3590/FROM )
  );
  defparam DLX_EXinst__n003264_SW0.INIT = 16'hFFFE;
  X_LUT4 DLX_EXinst__n003264_SW0 (
    .ADR0(CHOICE3587),
    .ADR1(CHOICE3583),
    .ADR2(DLX_IDinst_reg_out_B[20]),
    .ADR3(CHOICE3590),
    .O(\CHOICE3590/GROM )
  );
  X_BUF \CHOICE3590/XUSED  (
    .I(\CHOICE3590/FROM ),
    .O(CHOICE3590)
  );
  X_BUF \CHOICE3590/YUSED  (
    .I(\CHOICE3590/GROM ),
    .O(N163386)
  );
  defparam DLX_EXinst__n003264.INIT = 16'hFFFE;
  X_LUT4 DLX_EXinst__n003264 (
    .ADR0(N163386),
    .ADR1(DLX_IDinst_reg_out_B[21]),
    .ADR2(DLX_IDinst_reg_out_B[23]),
    .ADR3(DLX_IDinst_reg_out_B[22]),
    .O(\CHOICE3592/FROM )
  );
  defparam DLX_EXinst_Ker764191.INIT = 16'h0010;
  X_LUT4 DLX_EXinst_Ker764191 (
    .ADR0(CHOICE3570),
    .ADR1(CHOICE3576),
    .ADR2(DLX_EXinst__n0081),
    .ADR3(CHOICE3592),
    .O(\CHOICE3592/GROM )
  );
  X_BUF \CHOICE3592/XUSED  (
    .I(\CHOICE3592/FROM ),
    .O(CHOICE3592)
  );
  X_BUF \CHOICE3592/YUSED  (
    .I(\CHOICE3592/GROM ),
    .O(DLX_EXinst_N76421)
  );
  defparam DLX_EXinst__n003275.INIT = 16'hFEFE;
  X_LUT4 DLX_EXinst__n003275 (
    .ADR0(CHOICE3592),
    .ADR1(CHOICE3576),
    .ADR2(CHOICE3570),
    .ADR3(VCC),
    .O(\DLX_IDinst_RegFile_22_20/FROM )
  );
  defparam \DLX_EXinst__n0007<19>298 .INIT = 16'hC0EA;
  X_LUT4 \DLX_EXinst__n0007<19>298  (
    .ADR0(N163696),
    .ADR1(N138371),
    .ADR2(N148609),
    .ADR3(N148323),
    .O(\DLX_IDinst_RegFile_22_20/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_22_20/XUSED  (
    .I(\DLX_IDinst_RegFile_22_20/FROM ),
    .O(N148323)
  );
  X_BUF \DLX_IDinst_RegFile_22_20/YUSED  (
    .I(\DLX_IDinst_RegFile_22_20/GROM ),
    .O(CHOICE5342)
  );
  defparam DLX_EXinst__n014045_SW0.INIT = 16'hFEFF;
  X_LUT4 DLX_EXinst__n014045_SW0 (
    .ADR0(\DLX_IDinst_Imm[3] ),
    .ADR1(\DLX_IDinst_Imm[1] ),
    .ADR2(\DLX_IDinst_Imm[2] ),
    .ADR3(\DLX_IDinst_Imm[0] ),
    .O(\N163298/FROM )
  );
  defparam DLX_EXinst__n014036.INIT = 16'hDFCF;
  X_LUT4 DLX_EXinst__n014036 (
    .ADR0(\DLX_IDinst_Imm[1] ),
    .ADR1(\DLX_IDinst_Imm[3] ),
    .ADR2(\DLX_IDinst_Imm[2] ),
    .ADR3(\DLX_IDinst_Imm[0] ),
    .O(\N163298/GROM )
  );
  X_BUF \N163298/XUSED  (
    .I(\N163298/FROM ),
    .O(N163298)
  );
  X_BUF \N163298/YUSED  (
    .I(\N163298/GROM ),
    .O(CHOICE1311)
  );
  defparam DLX_EXinst__n014045.INIT = 16'hF444;
  X_LUT4 DLX_EXinst__n014045 (
    .ADR0(DLX_IDinst_IR_function_field[5]),
    .ADR1(CHOICE1311),
    .ADR2(N163298),
    .ADR3(\DLX_IDinst_Imm[4] ),
    .O(\CHOICE1313/FROM )
  );
  defparam DLX_EXinst__n014058.INIT = 16'hFF88;
  X_LUT4 DLX_EXinst__n014058 (
    .ADR0(\DLX_IDinst_Imm[1] ),
    .ADR1(CHOICE1299),
    .ADR2(VCC),
    .ADR3(CHOICE1313),
    .O(\CHOICE1313/GROM )
  );
  X_BUF \CHOICE1313/XUSED  (
    .I(\CHOICE1313/FROM ),
    .O(CHOICE1313)
  );
  X_BUF \CHOICE1313/YUSED  (
    .I(\CHOICE1313/GROM ),
    .O(N134884)
  );
  defparam \DLX_IDinst__n0142<1>_SW0 .INIT = 16'h02FF;
  X_LUT4 \DLX_IDinst__n0142<1>_SW0  (
    .ADR0(DLX_IDinst_N108165),
    .ADR1(DLX_IDinst_IR_latched[26]),
    .ADR2(DLX_IDinst_IR_latched[30]),
    .ADR3(N139656),
    .O(\DLX_IDinst_IR_opcode_field<1>/FROM )
  );
  defparam \DLX_IDinst__n0142<1> .INIT = 16'h2030;
  X_LUT4 \DLX_IDinst__n0142<1>  (
    .ADR0(DLX_IDinst__n0453),
    .ADR1(DLX_IDinst_N108456),
    .ADR2(DLX_IDinst_IR_latched[27]),
    .ADR3(N132373),
    .O(DLX_IDinst__n0142[1])
  );
  X_BUF \DLX_IDinst_IR_opcode_field<1>/XUSED  (
    .I(\DLX_IDinst_IR_opcode_field<1>/FROM ),
    .O(N132373)
  );
  defparam DLX_IDinst_RegFile_26_30_467.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_26_30_467 (
    .I(DLX_IDinst_WB_data_eff[30]),
    .CE(DLX_IDinst__n0602),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_26_30)
  );
  defparam \DLX_IDinst_slot_num_FFd4-In59_SW0 .INIT = 16'hCCDC;
  X_LUT4 \DLX_IDinst_slot_num_FFd4-In59_SW0  (
    .ADR0(DLX_IDinst_intr_slot),
    .ADR1(DLX_IDinst_slot_num_FFd4),
    .ADR2(DLX_IDinst_slot_num_FFd1),
    .ADR3(DLX_IDinst_delay_slot),
    .O(\N163469/FROM )
  );
  defparam \DLX_IDinst_slot_num_FFd4-In59 .INIT = 16'h3332;
  X_LUT4 \DLX_IDinst_slot_num_FFd4-In59  (
    .ADR0(DLX_IDinst_slot_num_FFd3),
    .ADR1(DLX_EXinst__n0144),
    .ADR2(DLX_IDinst_slot_num_FFd2),
    .ADR3(N163469),
    .O(\N163469/GROM )
  );
  X_BUF \N163469/XUSED  (
    .I(\N163469/FROM ),
    .O(N163469)
  );
  X_BUF \N163469/YUSED  (
    .I(\N163469/GROM ),
    .O(CHOICE2993)
  );
  defparam \DLX_IDinst__n0142<3>_SW0 .INIT = 16'h4500;
  X_LUT4 \DLX_IDinst__n0142<3>_SW0  (
    .ADR0(DLX_IDinst__n0453),
    .ADR1(DLX_IDinst_N107405),
    .ADR2(N164150),
    .ADR3(DLX_IDinst_N107033),
    .O(\DLX_IDinst_IR_opcode_field<3>/FROM )
  );
  defparam \DLX_IDinst__n0142<3> .INIT = 16'h3020;
  X_LUT4 \DLX_IDinst__n0142<3>  (
    .ADR0(DLX_IDinst__n0453),
    .ADR1(DLX_IDinst_N108456),
    .ADR2(DLX_IDinst_IR_latched[29]),
    .ADR3(N127652),
    .O(DLX_IDinst__n0142[3])
  );
  X_BUF \DLX_IDinst_IR_opcode_field<3>/XUSED  (
    .I(\DLX_IDinst_IR_opcode_field<3>/FROM ),
    .O(N127652)
  );
  defparam \DLX_IDinst__n0142<4>_SW0 .INIT = 16'h1F0F;
  X_LUT4 \DLX_IDinst__n0142<4>_SW0  (
    .ADR0(DLX_IDinst_IR_latched[27]),
    .ADR1(DLX_IDinst_IR_latched[26]),
    .ADR2(N139656),
    .ADR3(DLX_IDinst_N108165),
    .O(\DLX_IDinst_IR_opcode_field<4>/FROM )
  );
  defparam \DLX_IDinst__n0142<4> .INIT = 16'h4050;
  X_LUT4 \DLX_IDinst__n0142<4>  (
    .ADR0(DLX_IDinst_Ker1084541_1),
    .ADR1(DLX_IDinst__n0453),
    .ADR2(DLX_IDinst_IR_latched[30]),
    .ADR3(N132324),
    .O(DLX_IDinst__n0142[4])
  );
  X_BUF \DLX_IDinst_IR_opcode_field<4>/XUSED  (
    .I(\DLX_IDinst_IR_opcode_field<4>/FROM ),
    .O(N132324)
  );
  defparam \DLX_IDinst__n0143<0>_SW0 .INIT = 16'h5400;
  X_LUT4 \DLX_IDinst__n0143<0>_SW0  (
    .ADR0(DLX_IDinst__n0453),
    .ADR1(CHOICE2119),
    .ADR2(DLX_IDinst_N107405),
    .ADR3(DLX_IDinst_N107033),
    .O(\DLX_IDinst_Imm<0>/FROM )
  );
  defparam \DLX_IDinst__n0143<0> .INIT = 16'h4440;
  X_LUT4 \DLX_IDinst__n0143<0>  (
    .ADR0(DLX_IDinst_Ker1084541_1),
    .ADR1(DLX_IDinst_jtarget[0]),
    .ADR2(DLX_IDinst__n0453),
    .ADR3(N127400),
    .O(\DLX_IDinst_Imm<0>/GROM )
  );
  X_BUF \DLX_IDinst_Imm<0>/XUSED  (
    .I(\DLX_IDinst_Imm<0>/FROM ),
    .O(N127400)
  );
  X_BUF \DLX_IDinst_Imm<0>/YUSED  (
    .I(\DLX_IDinst_Imm<0>/GROM ),
    .O(DLX_IDinst__n0143[0])
  );
  defparam \DLX_IDinst_slot_num_FFd4-In88_SW0 .INIT = 16'hFFCC;
  X_LUT4 \DLX_IDinst_slot_num_FFd4-In88_SW0  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_slot_num_FFd4),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_slot_num_FFd3),
    .O(\DLX_IDinst_RegFile_2_6/FROM )
  );
  defparam \DLX_IDinst_slot_num_FFd4-In88 .INIT = 16'hFCA0;
  X_LUT4 \DLX_IDinst_slot_num_FFd4-In88  (
    .ADR0(DLX_IDinst_slot_num_FFd2),
    .ADR1(DLX_IDinst_delay_slot),
    .ADR2(DLX_IDinst_intr_slot),
    .ADR3(N163132),
    .O(\DLX_IDinst_RegFile_2_6/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_2_6/XUSED  (
    .I(\DLX_IDinst_RegFile_2_6/FROM ),
    .O(N163132)
  );
  X_BUF \DLX_IDinst_RegFile_2_6/YUSED  (
    .I(\DLX_IDinst_RegFile_2_6/GROM ),
    .O(CHOICE3000)
  );
  defparam \mask<1>_SW122_SW0 .INIT = 16'hDD30;
  X_LUT4 \mask<1>_SW122_SW0  (
    .ADR0(DLX_EXinst_ALU_result[1]),
    .ADR1(DLX_EXinst_ALU_result[0]),
    .ADR2(DLX_EXinst_word),
    .ADR3(DLX_EXinst_byte),
    .O(\N164178/FROM )
  );
  defparam \mask<1>_SW122 .INIT = 16'h0001;
  X_LUT4 \mask<1>_SW122  (
    .ADR0(DLX_EXinst_ALU_result[14]),
    .ADR1(DLX_EXinst_ALU_result[13]),
    .ADR2(DLX_EXinst_ALU_result[12]),
    .ADR3(N164178),
    .O(\N164178/GROM )
  );
  X_BUF \N164178/XUSED  (
    .I(\N164178/FROM ),
    .O(N164178)
  );
  X_BUF \N164178/YUSED  (
    .I(\N164178/GROM ),
    .O(mask_1_OBUF)
  );
  defparam DLX_IFinst_PC_12.INIT = 1'b0;
  X_SFF DLX_IFinst_PC_12 (
    .I(DLX_IFinst_NPC[12]),
    .CE(DLX_IFinst_PC_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_PC[12])
  );
  defparam DLX_IFinst_PC_21.INIT = 1'b0;
  X_SFF DLX_IFinst_PC_21 (
    .I(DLX_IFinst_NPC[21]),
    .CE(DLX_IFinst_PC_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_IFinst_PC[21])
  );
  defparam DLX_IFinst_PC_13.INIT = 1'b0;
  X_SFF DLX_IFinst_PC_13 (
    .I(DLX_IFinst_NPC[13]),
    .CE(DLX_IFinst_PC_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_PC[13])
  );
  defparam DLX_IFinst_PC_22.INIT = 1'b0;
  X_SFF DLX_IFinst_PC_22 (
    .I(DLX_IFinst_NPC[22]),
    .CE(DLX_IFinst_PC_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_IFinst_PC[22])
  );
  defparam DLX_IFinst_PC_14.INIT = 1'b0;
  X_SFF DLX_IFinst_PC_14 (
    .I(DLX_IFinst_NPC[14]),
    .CE(DLX_IFinst_PC_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_PC[14])
  );
  defparam DLX_IFinst_PC_23.INIT = 1'b0;
  X_SFF DLX_IFinst_PC_23 (
    .I(DLX_IFinst_NPC[23]),
    .CE(DLX_IFinst_PC_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_IFinst_PC[23])
  );
  defparam DLX_IDinst_RegFile_26_14_468.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_26_14_468 (
    .I(DLX_IDinst_WB_data_eff[14]),
    .CE(DLX_IDinst__n0602),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_26_14)
  );
  defparam DLX_IFinst_PC_15.INIT = 1'b0;
  X_SFF DLX_IFinst_PC_15 (
    .I(DLX_IFinst_NPC[15]),
    .CE(DLX_IFinst_PC_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_IFinst_PC[15])
  );
  defparam DLX_IFinst_PC_31.INIT = 1'b0;
  X_SFF DLX_IFinst_PC_31 (
    .I(DLX_IFinst_NPC[31]),
    .CE(DLX_IFinst_PC_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_IFinst_PC[31])
  );
  defparam DLX_IFinst_PC_24.INIT = 1'b0;
  X_SFF DLX_IFinst_PC_24 (
    .I(DLX_IFinst_NPC[24]),
    .CE(DLX_IFinst_PC_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_IFinst_PC[24])
  );
  defparam DLX_IFinst_PC_16.INIT = 1'b0;
  X_SFF DLX_IFinst_PC_16 (
    .I(DLX_IFinst_NPC[16]),
    .CE(DLX_IFinst_PC_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_IFinst_PC[16])
  );
  defparam DLX_IFinst_PC_25.INIT = 1'b0;
  X_SFF DLX_IFinst_PC_25 (
    .I(DLX_IFinst_NPC[25]),
    .CE(DLX_IFinst_PC_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_IFinst_PC[25])
  );
  defparam DLX_IFinst_PC_17.INIT = 1'b0;
  X_SFF DLX_IFinst_PC_17 (
    .I(DLX_IFinst_NPC[17]),
    .CE(DLX_IFinst_PC_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_IFinst_PC[17])
  );
  defparam DLX_IFinst_PC_26.INIT = 1'b0;
  X_SFF DLX_IFinst_PC_26 (
    .I(DLX_IFinst_NPC[26]),
    .CE(DLX_IFinst_PC_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_IFinst_PC[26])
  );
  defparam DLX_IFinst_PC_18.INIT = 1'b0;
  X_SFF DLX_IFinst_PC_18 (
    .I(DLX_IFinst_NPC[18]),
    .CE(DLX_IFinst_PC_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_IFinst_PC[18])
  );
  defparam DLX_IFinst_PC_19.INIT = 1'b0;
  X_SFF DLX_IFinst_PC_19 (
    .I(DLX_IFinst_NPC[19]),
    .CE(DLX_IFinst_PC_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_IFinst_PC[19])
  );
  defparam DLX_IDinst_RegFile_26_22_469.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_26_22_469 (
    .I(DLX_IDinst_WB_data_eff[22]),
    .CE(DLX_IDinst__n0602),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_26_22)
  );
  defparam DLX_IFinst_PC_29.INIT = 1'b0;
  X_SFF DLX_IFinst_PC_29 (
    .I(DLX_IFinst_NPC[29]),
    .CE(DLX_IFinst_PC_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_IFinst_PC[29])
  );
  defparam \DLX_EXinst_Mshift__n0020_Sh<30>1 .INIT = 16'hAAB8;
  X_LUT4 \DLX_EXinst_Mshift__n0020_Sh<30>1  (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(DLX_IDinst_Imm_1_1),
    .ADR2(DLX_IDinst_reg_out_A[30]),
    .ADR3(DLX_IDinst_Imm_0_1),
    .O(\DLX_EXinst_Mshift__n0020_Sh<30>/FROM )
  );
  defparam DLX_EXinst_Ker7515726.INIT = 16'h3202;
  X_LUT4 DLX_EXinst_Ker7515726 (
    .ADR0(\DLX_EXinst_Mshift__n0020_Sh[26] ),
    .ADR1(\DLX_IDinst_Imm[5] ),
    .ADR2(DLX_IDinst_Imm_2_1),
    .ADR3(\DLX_EXinst_Mshift__n0020_Sh[30] ),
    .O(\DLX_EXinst_Mshift__n0020_Sh<30>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0020_Sh<30>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0020_Sh<30>/FROM ),
    .O(\DLX_EXinst_Mshift__n0020_Sh[30] )
  );
  X_BUF \DLX_EXinst_Mshift__n0020_Sh<30>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0020_Sh<30>/GROM ),
    .O(CHOICE1865)
  );
  defparam \DLX_EXinst_Mshift__n0020_Sh<61>1 .INIT = 16'h44CC;
  X_LUT4 \DLX_EXinst_Mshift__n0020_Sh<61>1  (
    .ADR0(DLX_IDinst_Imm_0_1),
    .ADR1(DLX_IDinst_reg_out_A[31]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_Imm_1_1),
    .O(\DLX_EXinst_Mshift__n0020_Sh<61>/FROM )
  );
  defparam DLX_EXinst_Ker7514713.INIT = 16'hC840;
  X_LUT4 DLX_EXinst_Ker7514713 (
    .ADR0(DLX_IDinst_Imm_2_1),
    .ADR1(\DLX_IDinst_Imm[5] ),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(\DLX_EXinst_Mshift__n0020_Sh[61] ),
    .O(\DLX_EXinst_Mshift__n0020_Sh<61>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0020_Sh<61>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0020_Sh<61>/FROM ),
    .O(\DLX_EXinst_Mshift__n0020_Sh[61] )
  );
  X_BUF \DLX_EXinst_Mshift__n0020_Sh<61>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0020_Sh<61>/GROM ),
    .O(CHOICE1915)
  );
  defparam \DLX_EXinst_Mshift__n0020_Sh<29>1 .INIT = 16'hBB88;
  X_LUT4 \DLX_EXinst_Mshift__n0020_Sh<29>1  (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(DLX_IDinst_Imm_1_1),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N72791),
    .O(\DLX_EXinst_Mshift__n0020_Sh<29>/FROM )
  );
  defparam DLX_EXinst_Ker7565714.INIT = 16'h0B08;
  X_LUT4 DLX_EXinst_Ker7565714 (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(DLX_EXinst_N72815),
    .ADR2(\DLX_IDinst_Imm[5] ),
    .ADR3(\DLX_EXinst_Mshift__n0020_Sh[29] ),
    .O(\DLX_EXinst_Mshift__n0020_Sh<29>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0020_Sh<29>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0020_Sh<29>/FROM ),
    .O(\DLX_EXinst_Mshift__n0020_Sh[29] )
  );
  X_BUF \DLX_EXinst_Mshift__n0020_Sh<29>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0020_Sh<29>/GROM ),
    .O(CHOICE2017)
  );
  defparam \DLX_EXinst__n0007<20>246 .INIT = 16'hF444;
  X_LUT4 \DLX_EXinst__n0007<20>246  (
    .ADR0(N148323),
    .ADR1(N163485),
    .ADR2(DLX_EXinst_N74966),
    .ADR3(N148609),
    .O(\CHOICE4693/FROM )
  );
  defparam \DLX_EXinst__n0007<20>269 .INIT = 16'hB3A0;
  X_LUT4 \DLX_EXinst__n0007<20>269  (
    .ADR0(N163481),
    .ADR1(DLX_IDinst_reg_out_B[4]),
    .ADR2(DLX_IDinst_reg_out_A[20]),
    .ADR3(CHOICE4693),
    .O(\CHOICE4693/GROM )
  );
  X_BUF \CHOICE4693/XUSED  (
    .I(\CHOICE4693/FROM ),
    .O(CHOICE4693)
  );
  X_BUF \CHOICE4693/YUSED  (
    .I(\CHOICE4693/GROM ),
    .O(CHOICE4696)
  );
  defparam \DLX_EXinst__n0007<12>183 .INIT = 16'hF020;
  X_LUT4 \DLX_EXinst__n0007<12>183  (
    .ADR0(DLX_EXinst__n0054),
    .ADR1(\DLX_IDinst_Imm[12] ),
    .ADR2(DLX_IDinst_reg_out_A[12]),
    .ADR3(DLX_EXinst__n0053),
    .O(\CHOICE3809/FROM )
  );
  defparam \DLX_EXinst__n0007<12>187 .INIT = 16'hFF0E;
  X_LUT4 \DLX_EXinst__n0007<12>187  (
    .ADR0(CHOICE3802),
    .ADR1(CHOICE3803),
    .ADR2(\DLX_IDinst_Imm[4] ),
    .ADR3(CHOICE3809),
    .O(\CHOICE3809/GROM )
  );
  X_BUF \CHOICE3809/XUSED  (
    .I(\CHOICE3809/FROM ),
    .O(CHOICE3809)
  );
  X_BUF \CHOICE3809/YUSED  (
    .I(\CHOICE3809/GROM ),
    .O(CHOICE3810)
  );
  defparam \DLX_EXinst__n0007<21>213 .INIT = 16'hEAC0;
  X_LUT4 \DLX_EXinst__n0007<21>213  (
    .ADR0(DLX_EXinst__n0012[21]),
    .ADR1(N134884),
    .ADR2(DLX_EXinst_ALU_result[21]),
    .ADR3(DLX_EXinst__n0127),
    .O(\CHOICE4172/FROM )
  );
  defparam \DLX_EXinst__n0007<20>193 .INIT = 16'hEAC0;
  X_LUT4 \DLX_EXinst__n0007<20>193  (
    .ADR0(DLX_EXinst__n0012[20]),
    .ADR1(DLX_EXinst_ALU_result[20]),
    .ADR2(N134884),
    .ADR3(DLX_EXinst__n0127),
    .O(\CHOICE4172/GROM )
  );
  X_BUF \CHOICE4172/XUSED  (
    .I(\CHOICE4172/FROM ),
    .O(CHOICE4172)
  );
  X_BUF \CHOICE4172/YUSED  (
    .I(\CHOICE4172/GROM ),
    .O(CHOICE4676)
  );
  defparam \DLX_EXinst__n0007<14>134 .INIT = 16'hCC00;
  X_LUT4 \DLX_EXinst__n0007<14>134  (
    .ADR0(VCC),
    .ADR1(\DLX_IDinst_Imm[4] ),
    .ADR2(VCC),
    .ADR3(N139405),
    .O(\CHOICE3685/FROM )
  );
  defparam \DLX_EXinst__n0007<13>134 .INIT = 16'hCC00;
  X_LUT4 \DLX_EXinst__n0007<13>134  (
    .ADR0(VCC),
    .ADR1(\DLX_IDinst_Imm[4] ),
    .ADR2(VCC),
    .ADR3(N139100),
    .O(\CHOICE3685/GROM )
  );
  X_BUF \CHOICE3685/XUSED  (
    .I(\CHOICE3685/FROM ),
    .O(CHOICE3685)
  );
  X_BUF \CHOICE3685/YUSED  (
    .I(\CHOICE3685/GROM ),
    .O(CHOICE3740)
  );
  defparam \DLX_EXinst__n0007<5>134 .INIT = 16'h4448;
  X_LUT4 \DLX_EXinst__n0007<5>134  (
    .ADR0(DLX_IDinst_IR_opcode_field[1]),
    .ADR1(DLX_EXinst_N76011),
    .ADR2(DLX_IDinst_IR_opcode_field[0]),
    .ADR3(DLX_IDinst_reg_out_A[5]),
    .O(\CHOICE3969/FROM )
  );
  defparam \DLX_EXinst__n0007<13>127 .INIT = 16'h4448;
  X_LUT4 \DLX_EXinst__n0007<13>127  (
    .ADR0(DLX_IDinst_IR_opcode_field[1]),
    .ADR1(DLX_EXinst_N76011),
    .ADR2(DLX_IDinst_IR_opcode_field[0]),
    .ADR3(DLX_IDinst_reg_out_A[13]),
    .O(\CHOICE3969/GROM )
  );
  X_BUF \CHOICE3969/XUSED  (
    .I(\CHOICE3969/FROM ),
    .O(CHOICE3969)
  );
  X_BUF \CHOICE3969/YUSED  (
    .I(\CHOICE3969/GROM ),
    .O(CHOICE3738)
  );
  defparam \DLX_EXinst__n0007<21>227 .INIT = 16'hFCEE;
  X_LUT4 \DLX_EXinst__n0007<21>227  (
    .ADR0(DLX_EXinst__n0079),
    .ADR1(DLX_EXinst_N74245),
    .ADR2(DLX_EXinst__n0077),
    .ADR3(DLX_IDinst_reg_out_B[21]),
    .O(\DLX_IDinst_RegFile_3_10/FROM )
  );
  defparam \DLX_EXinst__n0007<21>152 .INIT = 16'hC4C0;
  X_LUT4 \DLX_EXinst__n0007<21>152  (
    .ADR0(DLX_IDinst_reg_out_A[21]),
    .ADR1(DLX_IDinst_reg_out_B[21]),
    .ADR2(DLX_EXinst__n0078),
    .ADR3(DLX_EXinst__n0079),
    .O(\DLX_IDinst_RegFile_3_10/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_3_10/XUSED  (
    .I(\DLX_IDinst_RegFile_3_10/FROM ),
    .O(CHOICE4179)
  );
  X_BUF \DLX_IDinst_RegFile_3_10/YUSED  (
    .I(\DLX_IDinst_RegFile_3_10/GROM ),
    .O(CHOICE4157)
  );
  defparam \DLX_EXinst__n0007<7>162 .INIT = 16'hC808;
  X_LUT4 \DLX_EXinst__n0007<7>162  (
    .ADR0(N133984),
    .ADR1(DLX_EXinst_N73267),
    .ADR2(\DLX_IDinst_Imm[2] ),
    .ADR3(DLX_EXinst_N74941),
    .O(\CHOICE3859/FROM )
  );
  defparam \DLX_EXinst__n0007<13>156 .INIT = 16'hC0A0;
  X_LUT4 \DLX_EXinst__n0007<13>156  (
    .ADR0(DLX_EXinst_N74711),
    .ADR1(DLX_EXinst_N74981),
    .ADR2(DLX_EXinst_N73267),
    .ADR3(\DLX_IDinst_Imm[2] ),
    .O(\CHOICE3859/GROM )
  );
  X_BUF \CHOICE3859/XUSED  (
    .I(\CHOICE3859/FROM ),
    .O(CHOICE3859)
  );
  X_BUF \CHOICE3859/YUSED  (
    .I(\CHOICE3859/GROM ),
    .O(CHOICE3747)
  );
  defparam \DLX_EXinst__n0007<30>100 .INIT = 16'hFFF0;
  X_LUT4 \DLX_EXinst__n0007<30>100  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(CHOICE4721),
    .ADR3(CHOICE4729),
    .O(\CHOICE4730/GROM )
  );
  X_BUF \CHOICE4730/YUSED  (
    .I(\CHOICE4730/GROM ),
    .O(CHOICE4730)
  );
  defparam DLX_EXinst_Ker762661.INIT = 16'h00CC;
  X_LUT4 DLX_EXinst_Ker762661 (
    .ADR0(VCC),
    .ADR1(DLX_EXinst__n0080),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[4]),
    .O(\DLX_EXinst_N76268/FROM )
  );
  defparam \DLX_EXinst__n0007<21>237 .INIT = 16'h88F8;
  X_LUT4 \DLX_EXinst__n0007<21>237  (
    .ADR0(DLX_IDinst_reg_out_A[21]),
    .ADR1(CHOICE4179),
    .ADR2(N145073),
    .ADR3(DLX_IDinst_reg_out_B[4]),
    .O(\DLX_EXinst_N76268/GROM )
  );
  X_BUF \DLX_EXinst_N76268/XUSED  (
    .I(\DLX_EXinst_N76268/FROM ),
    .O(DLX_EXinst_N76268)
  );
  X_BUF \DLX_EXinst_N76268/YUSED  (
    .I(\DLX_EXinst_N76268/GROM ),
    .O(CHOICE4181)
  );
  defparam \DLX_EXinst__n0007<14>157 .INIT = 16'hC808;
  X_LUT4 \DLX_EXinst__n0007<14>157  (
    .ADR0(N130311),
    .ADR1(DLX_EXinst_N76318),
    .ADR2(\DLX_IDinst_Imm[3] ),
    .ADR3(DLX_EXinst_N72993),
    .O(\CHOICE3693/FROM )
  );
  defparam \DLX_EXinst__n0007<13>157 .INIT = 16'h8A80;
  X_LUT4 \DLX_EXinst__n0007<13>157  (
    .ADR0(DLX_EXinst_N76318),
    .ADR1(DLX_EXinst_N72988),
    .ADR2(\DLX_IDinst_Imm[3] ),
    .ADR3(N130363),
    .O(\CHOICE3693/GROM )
  );
  X_BUF \CHOICE3693/XUSED  (
    .I(\CHOICE3693/FROM ),
    .O(CHOICE3693)
  );
  X_BUF \CHOICE3693/YUSED  (
    .I(\CHOICE3693/GROM ),
    .O(CHOICE3748)
  );
  defparam \DLX_EXinst__n0007<13>183 .INIT = 16'h8C88;
  X_LUT4 \DLX_EXinst__n0007<13>183  (
    .ADR0(DLX_EXinst__n0053),
    .ADR1(DLX_IDinst_reg_out_A[13]),
    .ADR2(\DLX_IDinst_Imm[13] ),
    .ADR3(DLX_EXinst__n0054),
    .O(\CHOICE3754/FROM )
  );
  defparam \DLX_EXinst__n0007<13>187 .INIT = 16'hFF54;
  X_LUT4 \DLX_EXinst__n0007<13>187  (
    .ADR0(\DLX_IDinst_Imm[4] ),
    .ADR1(CHOICE3747),
    .ADR2(CHOICE3748),
    .ADR3(CHOICE3754),
    .O(\CHOICE3754/GROM )
  );
  X_BUF \CHOICE3754/XUSED  (
    .I(\CHOICE3754/FROM ),
    .O(CHOICE3754)
  );
  X_BUF \CHOICE3754/YUSED  (
    .I(\CHOICE3754/GROM ),
    .O(CHOICE3755)
  );
  defparam \DLX_EXinst__n0007<21>272 .INIT = 16'hAAA8;
  X_LUT4 \DLX_EXinst__n0007<21>272  (
    .ADR0(DLX_EXinst__n0036),
    .ADR1(CHOICE4157),
    .ADR2(N163639),
    .ADR3(CHOICE4172),
    .O(\DLX_EXinst_ALU_result<21>/FROM )
  );
  defparam \DLX_EXinst__n0007<21>284 .INIT = 16'hFF88;
  X_LUT4 \DLX_EXinst__n0007<21>284  (
    .ADR0(CHOICE929),
    .ADR1(DLX_IDinst_reg_out_A[31]),
    .ADR2(VCC),
    .ADR3(CHOICE4184),
    .O(CHOICE4185)
  );
  X_BUF \DLX_EXinst_ALU_result<21>/XUSED  (
    .I(\DLX_EXinst_ALU_result<21>/FROM ),
    .O(CHOICE4184)
  );
  defparam \DLX_EXinst__n0007<17>217 .INIT = 16'hEAC0;
  X_LUT4 \DLX_EXinst__n0007<17>217  (
    .ADR0(N134884),
    .ADR1(DLX_EXinst__n0012[17]),
    .ADR2(DLX_EXinst__n0127),
    .ADR3(DLX_EXinst_ALU_result[17]),
    .O(\CHOICE5400/FROM )
  );
  defparam \DLX_EXinst__n0007<22>213 .INIT = 16'hEAC0;
  X_LUT4 \DLX_EXinst__n0007<22>213  (
    .ADR0(N134884),
    .ADR1(DLX_EXinst__n0012[22]),
    .ADR2(DLX_EXinst__n0127),
    .ADR3(DLX_EXinst_ALU_result[22]),
    .O(\CHOICE5400/GROM )
  );
  X_BUF \CHOICE5400/XUSED  (
    .I(\CHOICE5400/FROM ),
    .O(CHOICE5400)
  );
  X_BUF \CHOICE5400/YUSED  (
    .I(\CHOICE5400/GROM ),
    .O(CHOICE4107)
  );
  defparam \DLX_EXinst__n0007<28>169 .INIT = 16'hECA0;
  X_LUT4 \DLX_EXinst__n0007<28>169  (
    .ADR0(DLX_EXinst__n0012[28]),
    .ADR1(DLX_IDinst_reg_out_A[31]),
    .ADR2(DLX_EXinst_N73959),
    .ADR3(CHOICE929),
    .O(\CHOICE4879/FROM )
  );
  defparam \DLX_EXinst__n0007<30>143 .INIT = 16'hEAC0;
  X_LUT4 \DLX_EXinst__n0007<30>143  (
    .ADR0(DLX_EXinst_N73959),
    .ADR1(CHOICE929),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(DLX_EXinst__n0012[30]),
    .O(\CHOICE4879/GROM )
  );
  X_BUF \CHOICE4879/XUSED  (
    .I(\CHOICE4879/FROM ),
    .O(CHOICE4879)
  );
  X_BUF \CHOICE4879/YUSED  (
    .I(\CHOICE4879/GROM ),
    .O(CHOICE4734)
  );
  defparam \DLX_EXinst__n0007<6>134 .INIT = 16'h4448;
  X_LUT4 \DLX_EXinst__n0007<6>134  (
    .ADR0(DLX_IDinst_IR_opcode_field[1]),
    .ADR1(DLX_EXinst_N76011),
    .ADR2(DLX_IDinst_IR_opcode_field[0]),
    .ADR3(DLX_IDinst_reg_out_A[6]),
    .O(\DLX_IDinst_RegFile_7_4/FROM )
  );
  defparam \DLX_EXinst__n0007<14>127 .INIT = 16'h5060;
  X_LUT4 \DLX_EXinst__n0007<14>127  (
    .ADR0(DLX_IDinst_IR_opcode_field[1]),
    .ADR1(DLX_IDinst_IR_opcode_field[0]),
    .ADR2(DLX_EXinst_N76011),
    .ADR3(DLX_IDinst_reg_out_A[14]),
    .O(\DLX_IDinst_RegFile_7_4/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_7_4/XUSED  (
    .I(\DLX_IDinst_RegFile_7_4/FROM ),
    .O(CHOICE3910)
  );
  X_BUF \DLX_IDinst_RegFile_7_4/YUSED  (
    .I(\DLX_IDinst_RegFile_7_4/GROM ),
    .O(CHOICE3683)
  );
  defparam \DLX_EXinst__n0007<22>227 .INIT = 16'hFFCA;
  X_LUT4 \DLX_EXinst__n0007<22>227  (
    .ADR0(DLX_EXinst__n0079),
    .ADR1(DLX_EXinst__n0077),
    .ADR2(DLX_IDinst_reg_out_B[22]),
    .ADR3(DLX_EXinst_N74245),
    .O(\CHOICE4114/FROM )
  );
  defparam \DLX_EXinst__n0007<22>152 .INIT = 16'hF020;
  X_LUT4 \DLX_EXinst__n0007<22>152  (
    .ADR0(DLX_EXinst__n0079),
    .ADR1(DLX_IDinst_reg_out_A[22]),
    .ADR2(DLX_IDinst_reg_out_B[22]),
    .ADR3(DLX_EXinst__n0078),
    .O(\CHOICE4114/GROM )
  );
  X_BUF \CHOICE4114/XUSED  (
    .I(\CHOICE4114/FROM ),
    .O(CHOICE4114)
  );
  X_BUF \CHOICE4114/YUSED  (
    .I(\CHOICE4114/GROM ),
    .O(CHOICE4092)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_260_470 (
    .IA(DLX_IDinst_reg_out_B[30]),
    .IB(\CHOICE4741/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_196),
    .O(\CHOICE4741/CYMUXF )
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1961.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1961 (
    .ADR0(DLX_IDinst_reg_out_B[30]),
    .ADR1(DLX_IDinst_reg_out_A[30]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_196)
  );
  defparam \DLX_EXinst__n0007<30>170 .INIT = 16'hF400;
  X_LUT4 \DLX_EXinst__n0007<30>170  (
    .ADR0(DLX_IDinst_reg_out_A[30]),
    .ADR1(DLX_EXinst__n0079),
    .ADR2(DLX_EXinst__n0078),
    .ADR3(DLX_IDinst_reg_out_B[30]),
    .O(\CHOICE4741/GROM )
  );
  X_BUF \CHOICE4741/XBUSED  (
    .I(\CHOICE4741/CYMUXF ),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_260)
  );
  X_BUF \CHOICE4741/YUSED  (
    .I(\CHOICE4741/GROM ),
    .O(CHOICE4741)
  );
  X_BUF \CHOICE4741/CYINIT_471  (
    .I(DLX_EXinst_Mcompar__n0095_inst_cy_259),
    .O(\CHOICE4741/CYINIT )
  );
  defparam \DLX_EXinst__n0007<26>246_SW0 .INIT = 16'hFAEE;
  X_LUT4 \DLX_EXinst__n0007<26>246_SW0  (
    .ADR0(DLX_EXinst_N74245),
    .ADR1(DLX_EXinst__n0079),
    .ADR2(DLX_EXinst__n0077),
    .ADR3(DLX_IDinst_reg_out_B[26]),
    .O(\N163672/FROM )
  );
  defparam \DLX_EXinst__n0007<30>242 .INIT = 16'hFCFA;
  X_LUT4 \DLX_EXinst__n0007<30>242  (
    .ADR0(DLX_EXinst__n0079),
    .ADR1(DLX_EXinst__n0077),
    .ADR2(DLX_EXinst_N74245),
    .ADR3(DLX_IDinst_reg_out_B[30]),
    .O(\N163672/GROM )
  );
  X_BUF \N163672/XUSED  (
    .I(\N163672/FROM ),
    .O(N163672)
  );
  X_BUF \N163672/YUSED  (
    .I(\N163672/GROM ),
    .O(CHOICE4760)
  );
  defparam \DLX_EXinst__n0007<30>251 .INIT = 16'hECA0;
  X_LUT4 \DLX_EXinst__n0007<30>251  (
    .ADR0(N134884),
    .ADR1(CHOICE4760),
    .ADR2(DLX_EXinst_ALU_result[30]),
    .ADR3(DLX_IDinst_reg_out_A[30]),
    .O(\DLX_IDinst_RegFile_1_9/FROM )
  );
  defparam \DLX_EXinst__n0007<30>257 .INIT = 16'hFFCC;
  X_LUT4 \DLX_EXinst__n0007<30>257  (
    .ADR0(VCC),
    .ADR1(CHOICE4754),
    .ADR2(VCC),
    .ADR3(CHOICE4762),
    .O(\DLX_IDinst_RegFile_1_9/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_1_9/XUSED  (
    .I(\DLX_IDinst_RegFile_1_9/FROM ),
    .O(CHOICE4762)
  );
  X_BUF \DLX_IDinst_RegFile_1_9/YUSED  (
    .I(\DLX_IDinst_RegFile_1_9/GROM ),
    .O(CHOICE4763)
  );
  defparam \DLX_EXinst__n0007<28>367 .INIT = 16'hECA0;
  X_LUT4 \DLX_EXinst__n0007<28>367  (
    .ADR0(DLX_EXinst_N74130),
    .ADR1(DLX_EXinst_N73794),
    .ADR2(DLX_IDinst_reg_out_A[27]),
    .ADR3(DLX_IDinst_reg_out_A[26]),
    .O(\CHOICE4918/FROM )
  );
  defparam \DLX_EXinst__n0007<30>315 .INIT = 16'hEAC0;
  X_LUT4 \DLX_EXinst__n0007<30>315  (
    .ADR0(DLX_IDinst_reg_out_A[29]),
    .ADR1(DLX_EXinst_N73794),
    .ADR2(DLX_IDinst_reg_out_A[28]),
    .ADR3(DLX_EXinst_N74130),
    .O(\CHOICE4918/GROM )
  );
  X_BUF \CHOICE4918/XUSED  (
    .I(\CHOICE4918/FROM ),
    .O(CHOICE4918)
  );
  X_BUF \CHOICE4918/YUSED  (
    .I(\CHOICE4918/GROM ),
    .O(CHOICE4770)
  );
  defparam \DLX_EXinst__n0007<22>237 .INIT = 16'hB3A0;
  X_LUT4 \DLX_EXinst__n0007<22>237  (
    .ADR0(CHOICE4114),
    .ADR1(DLX_IDinst_reg_out_B[4]),
    .ADR2(DLX_IDinst_reg_out_A[22]),
    .ADR3(N145644),
    .O(\CHOICE4116/FROM )
  );
  defparam \DLX_EXinst__n0007<22>272_SW0 .INIT = 16'hFF08;
  X_LUT4 \DLX_EXinst__n0007<22>272_SW0  (
    .ADR0(DLX_EXinst__n0080),
    .ADR1(CHOICE4102),
    .ADR2(N148323),
    .ADR3(CHOICE4116),
    .O(\CHOICE4116/GROM )
  );
  X_BUF \CHOICE4116/XUSED  (
    .I(\CHOICE4116/FROM ),
    .O(CHOICE4116)
  );
  X_BUF \CHOICE4116/YUSED  (
    .I(\CHOICE4116/GROM ),
    .O(N163321)
  );
  defparam \DLX_EXinst__n0007<30>318 .INIT = 16'hFFEA;
  X_LUT4 \DLX_EXinst__n0007<30>318  (
    .ADR0(CHOICE4766),
    .ADR1(DLX_EXinst__n0036),
    .ADR2(CHOICE4764),
    .ADR3(CHOICE4770),
    .O(\DLX_EXinst_ALU_result<30>/FROM )
  );
  defparam \DLX_EXinst__n0007<30>3321 .INIT = 16'hFF44;
  X_LUT4 \DLX_EXinst__n0007<30>3321  (
    .ADR0(DLX_EXinst__n0036),
    .ADR1(CHOICE4731),
    .ADR2(VCC),
    .ADR3(CHOICE4771),
    .O(N162838)
  );
  X_BUF \DLX_EXinst_ALU_result<30>/XUSED  (
    .I(\DLX_EXinst_ALU_result<30>/FROM ),
    .O(CHOICE4771)
  );
  defparam \DLX_EXinst__n0007<14>183 .INIT = 16'h8C88;
  X_LUT4 \DLX_EXinst__n0007<14>183  (
    .ADR0(DLX_EXinst__n0053),
    .ADR1(DLX_IDinst_reg_out_A[14]),
    .ADR2(\DLX_IDinst_Imm[14] ),
    .ADR3(DLX_EXinst__n0054),
    .O(\CHOICE3699/FROM )
  );
  defparam \DLX_EXinst__n0007<14>187 .INIT = 16'hFF0E;
  X_LUT4 \DLX_EXinst__n0007<14>187  (
    .ADR0(CHOICE3693),
    .ADR1(CHOICE3692),
    .ADR2(\DLX_IDinst_Imm[4] ),
    .ADR3(CHOICE3699),
    .O(\CHOICE3699/GROM )
  );
  X_BUF \CHOICE3699/XUSED  (
    .I(\CHOICE3699/FROM ),
    .O(CHOICE3699)
  );
  X_BUF \CHOICE3699/YUSED  (
    .I(\CHOICE3699/GROM ),
    .O(CHOICE3700)
  );
  defparam \DLX_EXinst__n0007<31>129 .INIT = 16'hC8C0;
  X_LUT4 \DLX_EXinst__n0007<31>129  (
    .ADR0(DLX_IDinst_reg_out_B[3]),
    .ADR1(DLX_IDinst_reg_out_B[2]),
    .ADR2(CHOICE1765),
    .ADR3(\DLX_EXinst_Mshift__n0023_Sh[19] ),
    .O(\CHOICE5797/FROM )
  );
  defparam \DLX_EXinst__n0007<31>120 .INIT = 16'h3022;
  X_LUT4 \DLX_EXinst__n0007<31>120  (
    .ADR0(CHOICE5791),
    .ADR1(DLX_IDinst_reg_out_B[2]),
    .ADR2(\DLX_EXinst_Mshift__n0023_Sh[23] ),
    .ADR3(DLX_IDinst_reg_out_B[3]),
    .O(\CHOICE5797/GROM )
  );
  X_BUF \CHOICE5797/XUSED  (
    .I(\CHOICE5797/FROM ),
    .O(CHOICE5797)
  );
  X_BUF \CHOICE5797/YUSED  (
    .I(\CHOICE5797/GROM ),
    .O(CHOICE5796)
  );
  defparam DLX_IDinst_RegFile_26_24_472.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_26_24_472 (
    .I(DLX_IDinst_WB_data_eff[24]),
    .CE(DLX_IDinst__n0602),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_26_24)
  );
  defparam \DLX_EXinst__n0007<22>272 .INIT = 16'hAAA8;
  X_LUT4 \DLX_EXinst__n0007<22>272  (
    .ADR0(DLX_EXinst__n0036),
    .ADR1(CHOICE4107),
    .ADR2(N163321),
    .ADR3(CHOICE4092),
    .O(\DLX_EXinst_ALU_result<22>/FROM )
  );
  defparam \DLX_EXinst__n0007<22>284 .INIT = 16'hFFA0;
  X_LUT4 \DLX_EXinst__n0007<22>284  (
    .ADR0(CHOICE929),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(CHOICE4119),
    .O(CHOICE4120)
  );
  X_BUF \DLX_EXinst_ALU_result<22>/XUSED  (
    .I(\DLX_EXinst_ALU_result<22>/FROM ),
    .O(CHOICE4119)
  );
  defparam \DLX_EXinst__n0007<3>172 .INIT = 16'hA0AC;
  X_LUT4 \DLX_EXinst__n0007<3>172  (
    .ADR0(\DLX_EXinst_Mshift__n0019_Sh[11] ),
    .ADR1(DLX_IDinst_reg_out_A[3]),
    .ADR2(DLX_IDinst_reg_out_B[3]),
    .ADR3(DLX_EXinst_N73239),
    .O(\CHOICE5474/FROM )
  );
  defparam \DLX_EXinst__n0007<30>185 .INIT = 16'hF404;
  X_LUT4 \DLX_EXinst__n0007<30>185  (
    .ADR0(DLX_EXinst_N73239),
    .ADR1(DLX_IDinst_reg_out_A[30]),
    .ADR2(DLX_IDinst_reg_out_B[3]),
    .ADR3(\DLX_EXinst_Mshift__n0023_Sh[22] ),
    .O(\CHOICE5474/GROM )
  );
  X_BUF \CHOICE5474/XUSED  (
    .I(\CHOICE5474/FROM ),
    .O(CHOICE5474)
  );
  X_BUF \CHOICE5474/YUSED  (
    .I(\CHOICE5474/GROM ),
    .O(CHOICE4748)
  );
  defparam DLX_IDinst_RegFile_26_16_473.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_26_16_473 (
    .I(DLX_IDinst_WB_data_eff[16]),
    .CE(DLX_IDinst__n0602),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_26_16)
  );
  defparam \DLX_EXinst__n0007<25>170 .INIT = 16'hEAC0;
  X_LUT4 \DLX_EXinst__n0007<25>170  (
    .ADR0(DLX_EXinst__n0127),
    .ADR1(DLX_EXinst_ALU_result[25]),
    .ADR2(N134884),
    .ADR3(DLX_EXinst__n0012[25]),
    .O(\CHOICE5096/FROM )
  );
  defparam \DLX_EXinst__n0007<23>213 .INIT = 16'hEAC0;
  X_LUT4 \DLX_EXinst__n0007<23>213  (
    .ADR0(DLX_EXinst__n0127),
    .ADR1(N134884),
    .ADR2(DLX_EXinst_ALU_result[23]),
    .ADR3(DLX_EXinst__n0012[23]),
    .O(\CHOICE5096/GROM )
  );
  X_BUF \CHOICE5096/XUSED  (
    .I(\CHOICE5096/FROM ),
    .O(CHOICE5096)
  );
  X_BUF \CHOICE5096/YUSED  (
    .I(\CHOICE5096/GROM ),
    .O(CHOICE4042)
  );
  defparam \DLX_EXinst__n0007<27>97_SW0 .INIT = 16'h3600;
  X_LUT4 \DLX_EXinst__n0007<27>97_SW0  (
    .ADR0(DLX_IDinst_IR_opcode_field[0]),
    .ADR1(DLX_IDinst_IR_opcode_field[1]),
    .ADR2(DLX_IDinst_reg_out_A[27]),
    .ADR3(DLX_EXinst_N76011),
    .O(\N163518/FROM )
  );
  defparam \DLX_EXinst__n0007<15>144 .INIT = 16'h4448;
  X_LUT4 \DLX_EXinst__n0007<15>144  (
    .ADR0(DLX_IDinst_IR_opcode_field[1]),
    .ADR1(DLX_EXinst_N76011),
    .ADR2(DLX_IDinst_reg_out_A[15]),
    .ADR3(DLX_IDinst_IR_opcode_field[0]),
    .O(\N163518/GROM )
  );
  X_BUF \N163518/XUSED  (
    .I(\N163518/FROM ),
    .O(N163518)
  );
  X_BUF \N163518/YUSED  (
    .I(\N163518/GROM ),
    .O(CHOICE4294)
  );
  defparam \DLX_EXinst__n0007<23>227 .INIT = 16'hFAEE;
  X_LUT4 \DLX_EXinst__n0007<23>227  (
    .ADR0(DLX_EXinst_N74245),
    .ADR1(DLX_EXinst__n0079),
    .ADR2(DLX_EXinst__n0077),
    .ADR3(DLX_IDinst_reg_out_B[23]),
    .O(\DLX_IDinst_RegFile_15_7/FROM )
  );
  defparam \DLX_EXinst__n0007<23>152 .INIT = 16'hF400;
  X_LUT4 \DLX_EXinst__n0007<23>152  (
    .ADR0(DLX_IDinst_reg_out_A[23]),
    .ADR1(DLX_EXinst__n0079),
    .ADR2(DLX_EXinst__n0078),
    .ADR3(DLX_IDinst_reg_out_B[23]),
    .O(\DLX_IDinst_RegFile_15_7/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_15_7/XUSED  (
    .I(\DLX_IDinst_RegFile_15_7/FROM ),
    .O(CHOICE4049)
  );
  X_BUF \DLX_IDinst_RegFile_15_7/YUSED  (
    .I(\DLX_IDinst_RegFile_15_7/GROM ),
    .O(CHOICE4027)
  );
  defparam DLX_EXinst_Ker73792_SW0.INIT = 16'h0800;
  X_LUT4 DLX_EXinst_Ker73792_SW0 (
    .ADR0(DLX_EXinst_N75964),
    .ADR1(DLX_EXinst_N76501),
    .ADR2(N148323),
    .ADR3(DLX_EXinst__n0080),
    .O(\N126777/FROM )
  );
  defparam DLX_EXinst_Ker73792.INIT = 16'hFF40;
  X_LUT4 DLX_EXinst_Ker73792 (
    .ADR0(\DLX_IDinst_Imm[0] ),
    .ADR1(DLX_EXinst_N76490),
    .ADR2(DLX_IDinst_Imm_1_1),
    .ADR3(N126777),
    .O(\N126777/GROM )
  );
  X_BUF \N126777/XUSED  (
    .I(\N126777/FROM ),
    .O(N126777)
  );
  X_BUF \N126777/YUSED  (
    .I(\N126777/GROM ),
    .O(DLX_EXinst_N73794)
  );
  defparam DLX_IDinst_RegFile_18_25_474.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_18_25_474 (
    .I(DLX_IDinst_WB_data_eff[25]),
    .CE(DLX_IDinst__n0586),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_18_25)
  );
  defparam \DLX_EXinst__n0007<3>29 .INIT = 16'h8C88;
  X_LUT4 \DLX_EXinst__n0007<3>29  (
    .ADR0(DLX_EXinst__n0053),
    .ADR1(DLX_IDinst_reg_out_A[3]),
    .ADR2(\DLX_IDinst_Imm[3] ),
    .ADR3(DLX_EXinst__n0054),
    .O(\CHOICE5441/FROM )
  );
  defparam \DLX_EXinst__n0007<15>209 .INIT = 16'hC4C0;
  X_LUT4 \DLX_EXinst__n0007<15>209  (
    .ADR0(\DLX_IDinst_Imm[15] ),
    .ADR1(DLX_IDinst_reg_out_A[15]),
    .ADR2(DLX_EXinst__n0053),
    .ADR3(DLX_EXinst__n0054),
    .O(\CHOICE5441/GROM )
  );
  X_BUF \CHOICE5441/XUSED  (
    .I(\CHOICE5441/FROM ),
    .O(CHOICE5441)
  );
  X_BUF \CHOICE5441/YUSED  (
    .I(\CHOICE5441/GROM ),
    .O(CHOICE4312)
  );
  defparam \DLX_EXinst__n0007<28>349 .INIT = 16'hA0A0;
  X_LUT4 \DLX_EXinst__n0007<28>349  (
    .ADR0(DLX_EXinst_N73287),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[25]),
    .ADR3(VCC),
    .O(\CHOICE4914/FROM )
  );
  defparam \DLX_EXinst__n0007<30>297 .INIT = 16'hC0C0;
  X_LUT4 \DLX_EXinst__n0007<30>297  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[27]),
    .ADR2(DLX_EXinst_N73287),
    .ADR3(VCC),
    .O(\CHOICE4914/GROM )
  );
  X_BUF \CHOICE4914/XUSED  (
    .I(\CHOICE4914/FROM ),
    .O(CHOICE4914)
  );
  X_BUF \CHOICE4914/YUSED  (
    .I(\CHOICE4914/GROM ),
    .O(CHOICE4766)
  );
  defparam \DLX_EXinst__n0007<31>162 .INIT = 16'hAFAC;
  X_LUT4 \DLX_EXinst__n0007<31>162  (
    .ADR0(\DLX_EXinst_Mshift__n0023_Sh[47] ),
    .ADR1(CHOICE5796),
    .ADR2(DLX_IDinst_reg_out_B[4]),
    .ADR3(CHOICE5797),
    .O(\CHOICE5801/FROM )
  );
  defparam \DLX_EXinst__n0007<31>208 .INIT = 16'h3222;
  X_LUT4 \DLX_EXinst__n0007<31>208  (
    .ADR0(CHOICE5805),
    .ADR1(N148323),
    .ADR2(DLX_EXinst__n0080),
    .ADR3(CHOICE5801),
    .O(\CHOICE5801/GROM )
  );
  X_BUF \CHOICE5801/XUSED  (
    .I(\CHOICE5801/FROM ),
    .O(CHOICE5801)
  );
  X_BUF \CHOICE5801/YUSED  (
    .I(\CHOICE5801/GROM ),
    .O(CHOICE5807)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_164_475 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(\CHOICE5829/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_100),
    .O(\CHOICE5829/CYMUXF )
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_1001.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_1001 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(DLX_IDinst_reg_out_A[30]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_100)
  );
  defparam \DLX_EXinst__n0007<31>306 .INIT = 16'hE400;
  X_LUT4 \DLX_EXinst__n0007<31>306  (
    .ADR0(\DLX_IDinst_Imm[1] ),
    .ADR1(DLX_IDinst_reg_out_A[30]),
    .ADR2(DLX_IDinst_reg_out_A[28]),
    .ADR3(\DLX_IDinst_Imm[0] ),
    .O(\CHOICE5829/GROM )
  );
  X_BUF \CHOICE5829/XBUSED  (
    .I(\CHOICE5829/CYMUXF ),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_164)
  );
  X_BUF \CHOICE5829/YUSED  (
    .I(\CHOICE5829/GROM ),
    .O(CHOICE5829)
  );
  X_BUF \CHOICE5829/CYINIT_476  (
    .I(DLX_EXinst_Mcompar__n0063_inst_cy_163),
    .O(\CHOICE5829/CYINIT )
  );
  defparam \DLX_EXinst__n0007<5>162 .INIT = 16'hC808;
  X_LUT4 \DLX_EXinst__n0007<5>162  (
    .ADR0(N134488),
    .ADR1(DLX_EXinst_N73267),
    .ADR2(\DLX_IDinst_Imm[2] ),
    .ADR3(DLX_EXinst_N74951),
    .O(\CHOICE3977/FROM )
  );
  defparam \DLX_EXinst__n0007<15>164 .INIT = 16'h8A80;
  X_LUT4 \DLX_EXinst__n0007<15>164  (
    .ADR0(DLX_EXinst_N73267),
    .ADR1(DLX_EXinst_N75352),
    .ADR2(\DLX_IDinst_Imm[2] ),
    .ADR3(DLX_EXinst_N75139),
    .O(\CHOICE3977/GROM )
  );
  X_BUF \CHOICE3977/XUSED  (
    .I(\CHOICE3977/FROM ),
    .O(CHOICE3977)
  );
  X_BUF \CHOICE3977/YUSED  (
    .I(\CHOICE3977/GROM ),
    .O(CHOICE4301)
  );
  defparam DLX_EXinst_Ker7377322.INIT = 16'hC0C0;
  X_LUT4 DLX_EXinst_Ker7377322 (
    .ADR0(VCC),
    .ADR1(CHOICE1661),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(VCC),
    .O(\N136886/FROM )
  );
  defparam \DLX_EXinst__n0007<15>245 .INIT = 16'hF0C0;
  X_LUT4 \DLX_EXinst__n0007<15>245  (
    .ADR0(VCC),
    .ADR1(CHOICE1661),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(CHOICE929),
    .O(\N136886/GROM )
  );
  X_BUF \N136886/XUSED  (
    .I(\N136886/FROM ),
    .O(N136886)
  );
  X_BUF \N136886/YUSED  (
    .I(\N136886/GROM ),
    .O(CHOICE4316)
  );
  defparam DLX_EXinst_Ker759811.INIT = 16'hC0C0;
  X_LUT4 DLX_EXinst_Ker759811 (
    .ADR0(VCC),
    .ADR1(N148609),
    .ADR2(DLX_IDinst_reg_out_B[4]),
    .ADR3(VCC),
    .O(\DLX_IDinst_RegFile_3_11/FROM )
  );
  defparam \DLX_EXinst__n0007<23>237 .INIT = 16'hCE0A;
  X_LUT4 \DLX_EXinst__n0007<23>237  (
    .ADR0(N145258),
    .ADR1(CHOICE4049),
    .ADR2(DLX_IDinst_reg_out_B[4]),
    .ADR3(DLX_IDinst_reg_out_A[23]),
    .O(\DLX_IDinst_RegFile_3_11/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_3_11/XUSED  (
    .I(\DLX_IDinst_RegFile_3_11/FROM ),
    .O(DLX_EXinst_N75983)
  );
  X_BUF \DLX_IDinst_RegFile_3_11/YUSED  (
    .I(\DLX_IDinst_RegFile_3_11/GROM ),
    .O(CHOICE4051)
  );
  defparam \DLX_EXinst__n0007<31>261_SW0_SW0 .INIT = 16'h4000;
  X_LUT4 \DLX_EXinst__n0007<31>261_SW0_SW0  (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(DLX_IDinst_reg_out_B[5]),
    .ADR2(\DLX_EXinst_Mshift__n0019_Sh[127] ),
    .ADR3(N148609),
    .O(\N164729/FROM )
  );
  defparam \DLX_EXinst__n0007<31>190 .INIT = 16'h0C00;
  X_LUT4 \DLX_EXinst__n0007<31>190  (
    .ADR0(VCC),
    .ADR1(\DLX_EXinst_Mshift__n0019_Sh[127] ),
    .ADR2(DLX_IDinst_reg_out_B[4]),
    .ADR3(DLX_EXinst__n0081),
    .O(\N164729/GROM )
  );
  X_BUF \N164729/XUSED  (
    .I(\N164729/FROM ),
    .O(N164729)
  );
  X_BUF \N164729/YUSED  (
    .I(\N164729/GROM ),
    .O(CHOICE5805)
  );
  defparam \DLX_EXinst__n0007<16>104 .INIT = 16'hAACC;
  X_LUT4 \DLX_EXinst__n0007<16>104  (
    .ADR0(DLX_EXinst__n0077),
    .ADR1(DLX_EXinst__n0079),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[16]),
    .O(\CHOICE4587/FROM )
  );
  defparam \DLX_EXinst__n0007<16>113 .INIT = 16'hFE00;
  X_LUT4 \DLX_EXinst__n0007<16>113  (
    .ADR0(CHOICE4587),
    .ADR1(DLX_EXinst__n0083),
    .ADR2(DLX_EXinst__n0078),
    .ADR3(DLX_IDinst_reg_out_A[16]),
    .O(\CHOICE4587/GROM )
  );
  X_BUF \CHOICE4587/XUSED  (
    .I(\CHOICE4587/FROM ),
    .O(CHOICE4587)
  );
  X_BUF \CHOICE4587/YUSED  (
    .I(\CHOICE4587/GROM ),
    .O(CHOICE4589)
  );
  defparam \DLX_EXinst__n0007<23>272 .INIT = 16'hCCC8;
  X_LUT4 \DLX_EXinst__n0007<23>272  (
    .ADR0(N163390),
    .ADR1(DLX_EXinst__n0036),
    .ADR2(CHOICE4042),
    .ADR3(CHOICE4027),
    .O(\DLX_EXinst_ALU_result<23>/FROM )
  );
  defparam \DLX_EXinst__n0007<23>284 .INIT = 16'hFFA0;
  X_LUT4 \DLX_EXinst__n0007<23>284  (
    .ADR0(CHOICE929),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(CHOICE4054),
    .O(CHOICE4055)
  );
  X_BUF \DLX_EXinst_ALU_result<23>/XUSED  (
    .I(\DLX_EXinst_ALU_result<23>/FROM ),
    .O(CHOICE4054)
  );
  defparam DLX_EXinst_Ker7436792.INIT = 16'h2E22;
  X_LUT4 DLX_EXinst_Ker7436792 (
    .ADR0(DLX_EXinst_N73093),
    .ADR1(DLX_IDinst_reg_out_B[2]),
    .ADR2(DLX_IDinst_reg_out_B[3]),
    .ADR3(\DLX_EXinst_Mshift__n0019_Sh[25] ),
    .O(\DLX_IDinst_RegFile_22_8/FROM )
  );
  defparam \DLX_EXinst__n0007<24>120 .INIT = 16'hCA00;
  X_LUT4 \DLX_EXinst__n0007<24>120  (
    .ADR0(\DLX_EXinst_Mshift__n0023_Sh[16] ),
    .ADR1(\DLX_EXinst_Mshift__n0023_Sh[12] ),
    .ADR2(DLX_IDinst_reg_out_B[2]),
    .ADR3(DLX_IDinst_reg_out_B[3]),
    .O(\DLX_IDinst_RegFile_22_8/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_22_8/XUSED  (
    .I(\DLX_IDinst_RegFile_22_8/FROM ),
    .O(CHOICE3043)
  );
  X_BUF \DLX_IDinst_RegFile_22_8/YUSED  (
    .I(\DLX_IDinst_RegFile_22_8/GROM ),
    .O(CHOICE5618)
  );
  defparam DLX_EXinst_Ker761221.INIT = 16'hC0C0;
  X_LUT4 DLX_EXinst_Ker761221 (
    .ADR0(VCC),
    .ADR1(N147520),
    .ADR2(\DLX_IDinst_Imm[5] ),
    .ADR3(VCC),
    .O(\DLX_EXinst_N76124/FROM )
  );
  defparam \DLX_EXinst__n0007<31>507 .INIT = 16'h7350;
  X_LUT4 \DLX_EXinst__n0007<31>507  (
    .ADR0(\DLX_IDinst_Imm[5] ),
    .ADR1(\DLX_IDinst_Imm[31] ),
    .ADR2(N147520),
    .ADR3(DLX_EXinst__n0054),
    .O(\DLX_EXinst_N76124/GROM )
  );
  X_BUF \DLX_EXinst_N76124/XUSED  (
    .I(\DLX_EXinst_N76124/FROM ),
    .O(DLX_EXinst_N76124)
  );
  X_BUF \DLX_EXinst_N76124/YUSED  (
    .I(\DLX_EXinst_N76124/GROM ),
    .O(CHOICE5861)
  );
  defparam \DLX_EXinst__n0007<16>140 .INIT = 16'hFFEC;
  X_LUT4 \DLX_EXinst__n0007<16>140  (
    .ADR0(CHOICE4574),
    .ADR1(CHOICE4579),
    .ADR2(DLX_EXinst_N76338),
    .ADR3(CHOICE4591),
    .O(\CHOICE4592/FROM )
  );
  defparam \DLX_EXinst__n0007<16>168 .INIT = 16'hEAC0;
  X_LUT4 \DLX_EXinst__n0007<16>168  (
    .ADR0(DLX_EXinst__n0036),
    .ADR1(DLX_EXinst_N73959),
    .ADR2(DLX_EXinst__n0012[16]),
    .ADR3(CHOICE4592),
    .O(\CHOICE4592/GROM )
  );
  X_BUF \CHOICE4592/XUSED  (
    .I(\CHOICE4592/FROM ),
    .O(CHOICE4592)
  );
  X_BUF \CHOICE4592/YUSED  (
    .I(\CHOICE4592/GROM ),
    .O(CHOICE4594)
  );
  defparam \DLX_EXinst__n0007<9>164 .INIT = 16'hA0C0;
  X_LUT4 \DLX_EXinst__n0007<9>164  (
    .ADR0(DLX_EXinst_N74711),
    .ADR1(DLX_EXinst_N74951),
    .ADR2(DLX_EXinst_N76473),
    .ADR3(\DLX_IDinst_Imm[2] ),
    .O(\CHOICE4545/FROM )
  );
  defparam \DLX_EXinst__n0007<16>301 .INIT = 16'hFFC0;
  X_LUT4 \DLX_EXinst__n0007<16>301  (
    .ADR0(VCC),
    .ADR1(\DLX_EXinst_Mshift__n0020_Sh[80] ),
    .ADR2(DLX_EXinst_N76473),
    .ADR3(CHOICE4624),
    .O(\CHOICE4545/GROM )
  );
  X_BUF \CHOICE4545/XUSED  (
    .I(\CHOICE4545/FROM ),
    .O(CHOICE4545)
  );
  X_BUF \CHOICE4545/YUSED  (
    .I(\CHOICE4545/GROM ),
    .O(CHOICE4625)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_5861.INIT = 16'h8000;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_5861 (
    .ADR0(DLX_IDinst_jtarget[22]),
    .ADR1(DLX_IDinst_jtarget[25]),
    .ADR2(DLX_IDinst_jtarget[23]),
    .ADR3(DLX_IDinst_jtarget[24]),
    .O(\DLX_IFinst_IR_previous<20>/FROM )
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_5801.INIT = 16'h0008;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_5801 (
    .ADR0(DLX_IDinst_jtarget[22]),
    .ADR1(DLX_IDinst_jtarget[25]),
    .ADR2(DLX_IDinst_jtarget[23]),
    .ADR3(DLX_IDinst_jtarget[24]),
    .O(\DLX_IFinst_IR_previous<20>/GROM )
  );
  X_BUF \DLX_IFinst_IR_previous<20>/XUSED  (
    .I(\DLX_IFinst_IR_previous<20>/FROM ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_586)
  );
  X_BUF \DLX_IFinst_IR_previous<20>/YUSED  (
    .I(\DLX_IFinst_IR_previous<20>/GROM ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_580)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_5851.INIT = 16'h2000;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_5851 (
    .ADR0(DLX_IDinst_jtarget[23]),
    .ADR1(DLX_IDinst_jtarget[22]),
    .ADR2(DLX_IDinst_jtarget[25]),
    .ADR3(DLX_IDinst_jtarget[24]),
    .O(\DLX_IDinst_RegFile_2_19/FROM )
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_5721.INIT = 16'h0010;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_5721 (
    .ADR0(DLX_IDinst_jtarget[25]),
    .ADR1(DLX_IDinst_jtarget[23]),
    .ADR2(DLX_IDinst_jtarget[22]),
    .ADR3(DLX_IDinst_jtarget[24]),
    .O(\DLX_IDinst_RegFile_2_19/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_2_19/XUSED  (
    .I(\DLX_IDinst_RegFile_2_19/FROM ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_585)
  );
  X_BUF \DLX_IDinst_RegFile_2_19/YUSED  (
    .I(\DLX_IDinst_RegFile_2_19/GROM ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_572)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_5841.INIT = 16'h0800;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_5841 (
    .ADR0(DLX_IDinst_jtarget[25]),
    .ADR1(DLX_IDinst_jtarget[24]),
    .ADR2(DLX_IDinst_jtarget[23]),
    .ADR3(DLX_IDinst_jtarget[22]),
    .O(\DLX_IDinst_Mmux__COND_5_inst_lut4_584/FROM )
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_5811.INIT = 16'h0040;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_5811 (
    .ADR0(DLX_IDinst_jtarget[22]),
    .ADR1(DLX_IDinst_jtarget[25]),
    .ADR2(DLX_IDinst_jtarget[23]),
    .ADR3(DLX_IDinst_jtarget[24]),
    .O(\DLX_IDinst_Mmux__COND_5_inst_lut4_584/GROM )
  );
  X_BUF \DLX_IDinst_Mmux__COND_5_inst_lut4_584/XUSED  (
    .I(\DLX_IDinst_Mmux__COND_5_inst_lut4_584/FROM ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_584)
  );
  X_BUF \DLX_IDinst_Mmux__COND_5_inst_lut4_584/YUSED  (
    .I(\DLX_IDinst_Mmux__COND_5_inst_lut4_584/GROM ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_581)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_5821.INIT = 16'h4000;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_5821 (
    .ADR0(DLX_IDinst_jtarget[24]),
    .ADR1(DLX_IDinst_jtarget[22]),
    .ADR2(DLX_IDinst_jtarget[23]),
    .ADR3(DLX_IDinst_jtarget[25]),
    .O(\DLX_IDinst_Mmux__COND_5_inst_lut4_582/FROM )
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_5731.INIT = 16'h0002;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_5731 (
    .ADR0(DLX_IDinst_jtarget[23]),
    .ADR1(DLX_IDinst_jtarget[24]),
    .ADR2(DLX_IDinst_jtarget[22]),
    .ADR3(DLX_IDinst_jtarget[25]),
    .O(\DLX_IDinst_Mmux__COND_5_inst_lut4_582/GROM )
  );
  X_BUF \DLX_IDinst_Mmux__COND_5_inst_lut4_582/XUSED  (
    .I(\DLX_IDinst_Mmux__COND_5_inst_lut4_582/FROM ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_582)
  );
  X_BUF \DLX_IDinst_Mmux__COND_5_inst_lut4_582/YUSED  (
    .I(\DLX_IDinst_Mmux__COND_5_inst_lut4_582/GROM ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_573)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_5781.INIT = 16'h0800;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_5781 (
    .ADR0(DLX_IDinst_jtarget[23]),
    .ADR1(DLX_IDinst_jtarget[24]),
    .ADR2(DLX_IDinst_jtarget[25]),
    .ADR3(DLX_IDinst_jtarget[22]),
    .O(\DLX_IDinst_Mmux__COND_5_inst_lut4_578/FROM )
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_5741.INIT = 16'h0020;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_5741 (
    .ADR0(DLX_IDinst_jtarget[23]),
    .ADR1(DLX_IDinst_jtarget[25]),
    .ADR2(DLX_IDinst_jtarget[22]),
    .ADR3(DLX_IDinst_jtarget[24]),
    .O(\DLX_IDinst_Mmux__COND_5_inst_lut4_578/GROM )
  );
  X_BUF \DLX_IDinst_Mmux__COND_5_inst_lut4_578/XUSED  (
    .I(\DLX_IDinst_Mmux__COND_5_inst_lut4_578/FROM ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_578)
  );
  X_BUF \DLX_IDinst_Mmux__COND_5_inst_lut4_578/YUSED  (
    .I(\DLX_IDinst_Mmux__COND_5_inst_lut4_578/GROM ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_574)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_5771.INIT = 16'h0400;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_5771 (
    .ADR0(DLX_IDinst_jtarget[25]),
    .ADR1(DLX_IDinst_jtarget[23]),
    .ADR2(DLX_IDinst_jtarget[22]),
    .ADR3(DLX_IDinst_jtarget[24]),
    .O(\DLX_IFinst_IR_previous<16>/FROM )
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_5751.INIT = 16'h0010;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_5751 (
    .ADR0(DLX_IDinst_jtarget[22]),
    .ADR1(DLX_IDinst_jtarget[25]),
    .ADR2(DLX_IDinst_jtarget[24]),
    .ADR3(DLX_IDinst_jtarget[23]),
    .O(\DLX_IFinst_IR_previous<16>/GROM )
  );
  X_BUF \DLX_IFinst_IR_previous<16>/XUSED  (
    .I(\DLX_IFinst_IR_previous<16>/FROM ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_577)
  );
  X_BUF \DLX_IFinst_IR_previous<16>/YUSED  (
    .I(\DLX_IFinst_IR_previous<16>/GROM ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_575)
  );
  defparam \DLX_IDinst__n0146<31>39 .INIT = 16'h4A40;
  X_LUT4 \DLX_IDinst__n0146<31>39  (
    .ADR0(DLX_IDinst_jtarget[22]),
    .ADR1(\DLX_IDinst_Cause_Reg[31] ),
    .ADR2(DLX_IDinst_jtarget[21]),
    .ADR3(DLX_IDinst_EPC[31]),
    .O(\DLX_IDinst_RegFile_2_27/FROM )
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_5761.INIT = 16'h0020;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_5761 (
    .ADR0(DLX_IDinst_jtarget[24]),
    .ADR1(DLX_IDinst_jtarget[25]),
    .ADR2(DLX_IDinst_jtarget[22]),
    .ADR3(DLX_IDinst_jtarget[23]),
    .O(\DLX_IDinst_RegFile_2_27/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_2_27/XUSED  (
    .I(\DLX_IDinst_RegFile_2_27/FROM ),
    .O(CHOICE3230)
  );
  X_BUF \DLX_IDinst_RegFile_2_27/YUSED  (
    .I(\DLX_IDinst_RegFile_2_27/GROM ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_576)
  );
  defparam DLX_IDinst_RegFile_18_11_477.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_18_11_477 (
    .I(DLX_IDinst_WB_data_eff[11]),
    .CE(DLX_IDinst__n0586),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_18_11)
  );
  defparam \DLX_EXinst_Mshift__n0020_Sh<88>1 .INIT = 16'hBB88;
  X_LUT4 \DLX_EXinst_Mshift__n0020_Sh<88>1  (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(DLX_IDinst_Imm_3_1),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N73379),
    .O(\DLX_IDinst_RegFile_18_11/FROM )
  );
  defparam \DLX_EXinst__n0007<8>228 .INIT = 16'hCAC0;
  X_LUT4 \DLX_EXinst__n0007<8>228  (
    .ADR0(\DLX_IDinst_Imm[4] ),
    .ADR1(DLX_EXinst_N76382),
    .ADR2(\DLX_IDinst_Imm[5] ),
    .ADR3(\DLX_EXinst_Mshift__n0020_Sh[88] ),
    .O(\DLX_IDinst_RegFile_18_11/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_18_11/XUSED  (
    .I(\DLX_IDinst_RegFile_18_11/FROM ),
    .O(\DLX_EXinst_Mshift__n0020_Sh[88] )
  );
  X_BUF \DLX_IDinst_RegFile_18_11/YUSED  (
    .I(\DLX_IDinst_RegFile_18_11/GROM ),
    .O(CHOICE5185)
  );
  defparam \DLX_IDinst_slot_num_FFd2-In46 .INIT = 16'h8A00;
  X_LUT4 \DLX_IDinst_slot_num_FFd2-In46  (
    .ADR0(N146700),
    .ADR1(DLX_IDinst_delay_slot),
    .ADR2(FREEZE_IBUF),
    .ADR3(DLX_IDinst_slot_num_FFd2),
    .O(\DLX_IDinst_slot_num_FFd2/FROM )
  );
  defparam \DLX_IDinst_slot_num_FFd2-In65 .INIT = 16'h5540;
  X_LUT4 \DLX_IDinst_slot_num_FFd2-In65  (
    .ADR0(DLX_IDinst_N108100),
    .ADR1(CHOICE2128),
    .ADR2(CHOICE2131),
    .ADR3(CHOICE2136),
    .O(\DLX_IDinst_slot_num_FFd2-In )
  );
  X_BUF \DLX_IDinst_slot_num_FFd2/XUSED  (
    .I(\DLX_IDinst_slot_num_FFd2/FROM ),
    .O(CHOICE2136)
  );
  defparam DLX_IDinst_RegFile_15_16_478.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_15_16_478 (
    .I(DLX_IDinst_WB_data_eff[16]),
    .CE(DLX_IDinst__n0580),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_15_16)
  );
  defparam \vga_top_vga1_blueout<2>1 .INIT = 16'h0300;
  X_LUT4 \vga_top_vga1_blueout<2>1  (
    .ADR0(VCC),
    .ADR1(vram_out_vga_eff),
    .ADR2(reset_IBUF_1),
    .ADR3(vga_top_vga1_videoon),
    .O(\DLX_IDinst_RegFile_15_16/FROM )
  );
  defparam \vga_top_vga1_greenout<0>1 .INIT = 16'h0300;
  X_LUT4 \vga_top_vga1_greenout<0>1  (
    .ADR0(VCC),
    .ADR1(reset_IBUF_1),
    .ADR2(vram_out_vga_eff),
    .ADR3(vga_top_vga1_videoon),
    .O(\DLX_IDinst_RegFile_15_16/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_15_16/XUSED  (
    .I(\DLX_IDinst_RegFile_15_16/FROM ),
    .O(blue_2_OBUF)
  );
  X_BUF \DLX_IDinst_RegFile_15_16/YUSED  (
    .I(\DLX_IDinst_RegFile_15_16/GROM ),
    .O(green_0_OBUF)
  );
  defparam DLX_IDinst_RegFile_26_5_479.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_26_5_479 (
    .I(DLX_MEMinst_RF_data_in[5]),
    .CE(DLX_IDinst__n0602),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_26_5)
  );
  defparam DLX_EXinst_Mcompar__n0067_inst_cy_229_480.INIT = 16'h8E8E;
  X_LUT4 DLX_EXinst_Mcompar__n0067_inst_cy_229_480 (
    .ADR0(DLX_EXinst_Mcompar__n0067_inst_cy_228),
    .ADR1(DLX_IDinst_Imm_31_1),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(VCC),
    .O(\DLX_IDinst_RegFile_26_5/FROM )
  );
  defparam \DLX_EXinst__n0007<0>429 .INIT = 16'h1032;
  X_LUT4 \DLX_EXinst__n0007<0>429  (
    .ADR0(DLX_IDinst_IR_opcode_field[2]),
    .ADR1(DLX_IDinst_IR_opcode_field[0]),
    .ADR2(DLX_EXinst__n0059),
    .ADR3(DLX_EXinst_Mcompar__n0067_inst_cy_229),
    .O(\DLX_IDinst_RegFile_26_5/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_26_5/XUSED  (
    .I(\DLX_IDinst_RegFile_26_5/FROM ),
    .O(DLX_EXinst_Mcompar__n0067_inst_cy_229)
  );
  X_BUF \DLX_IDinst_RegFile_26_5/YUSED  (
    .I(\DLX_IDinst_RegFile_26_5/GROM ),
    .O(CHOICE5958)
  );
  defparam \DLX_IDinst_slot_num_FFd3-In1 .INIT = 16'hC8C8;
  X_LUT4 \DLX_IDinst_slot_num_FFd3-In1  (
    .ADR0(DLX_IDinst_intr_slot),
    .ADR1(DLX_IDinst_slot_num_FFd1),
    .ADR2(DLX_IDinst_delay_slot),
    .ADR3(VCC),
    .O(\DLX_IDinst_slot_num_FFd3-In )
  );
  defparam \DLX_IDinst_slot_num_FFd4-In14 .INIT = 16'h0F02;
  X_LUT4 \DLX_IDinst_slot_num_FFd4-In14  (
    .ADR0(DLX_IDinst_slot_num_FFd1),
    .ADR1(DLX_IDinst_intr_slot),
    .ADR2(DLX_IDinst_delay_slot),
    .ADR3(DLX_IDinst_slot_num_FFd2),
    .O(\DLX_IDinst_slot_num_FFd3/GROM )
  );
  X_BUF \DLX_IDinst_slot_num_FFd3/YUSED  (
    .I(\DLX_IDinst_slot_num_FFd3/GROM ),
    .O(CHOICE2981)
  );
  defparam \DLX_IDinst_slot_num_FFd4-In30 .INIT = 16'hAAA8;
  X_LUT4 \DLX_IDinst_slot_num_FFd4-In30  (
    .ADR0(N164719),
    .ADR1(DLX_IDinst_slot_num_FFd4),
    .ADR2(DLX_IDinst_slot_num_FFd3),
    .ADR3(CHOICE2981),
    .O(\DLX_IDinst_slot_num_FFd4/FROM )
  );
  defparam \DLX_IDinst_slot_num_FFd4-In95 .INIT = 16'hFFFC;
  X_LUT4 \DLX_IDinst_slot_num_FFd4-In95  (
    .ADR0(VCC),
    .ADR1(CHOICE2993),
    .ADR2(CHOICE3000),
    .ADR3(CHOICE2984),
    .O(\DLX_IDinst_slot_num_FFd4-In )
  );
  X_BUF \DLX_IDinst_slot_num_FFd4/XUSED  (
    .I(\DLX_IDinst_slot_num_FFd4/FROM ),
    .O(CHOICE2984)
  );
  defparam \vga_top_vga1_blueout<0>1 .INIT = 16'h0404;
  X_LUT4 \vga_top_vga1_blueout<0>1  (
    .ADR0(reset_IBUF_1),
    .ADR1(vga_top_vga1_videoon),
    .ADR2(vram_out_vga_eff),
    .ADR3(VCC),
    .O(\DLX_IDinst_RegFile_2_21/FROM )
  );
  defparam \vga_top_vga1_greenout<2>1 .INIT = 16'h1100;
  X_LUT4 \vga_top_vga1_greenout<2>1  (
    .ADR0(vram_out_vga_eff),
    .ADR1(reset_IBUF_1),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_videoon),
    .O(\DLX_IDinst_RegFile_2_21/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_2_21/XUSED  (
    .I(\DLX_IDinst_RegFile_2_21/FROM ),
    .O(blue_0_OBUF)
  );
  X_BUF \DLX_IDinst_RegFile_2_21/YUSED  (
    .I(\DLX_IDinst_RegFile_2_21/GROM ),
    .O(green_2_OBUF)
  );
  X_ZERO \DLX_EXinst_noop/LOGIC_ZERO_481  (
    .O(\DLX_EXinst_noop/LOGIC_ZERO )
  );
  defparam DLX_IDinst_PIPEEMPTY1.INIT = 16'hC000;
  X_LUT4 DLX_IDinst_PIPEEMPTY1 (
    .ADR0(VCC),
    .ADR1(FREEZE_IBUF),
    .ADR2(DLX_EXinst_noop),
    .ADR3(DLX_MEMinst_noop),
    .O(\DLX_EXinst_noop/FROM )
  );
  defparam \DLX_IDinst_slot_num_FFd2-In25 .INIT = 16'h0033;
  X_LUT4 \DLX_IDinst_slot_num_FFd2-In25  (
    .ADR0(VCC),
    .ADR1(FREEZE_IBUF),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_delay_slot),
    .O(\DLX_EXinst_noop/GROM )
  );
  X_BUF \DLX_EXinst_noop/XUSED  (
    .I(\DLX_EXinst_noop/FROM ),
    .O(PIPEEMPTY_OBUF)
  );
  X_BUF \DLX_EXinst_noop/YUSED  (
    .I(\DLX_EXinst_noop/GROM ),
    .O(CHOICE2131)
  );
  defparam \DLX_EXinst_Mshift__n0021_Sh<10>1 .INIT = 16'hCACA;
  X_LUT4 \DLX_EXinst_Mshift__n0021_Sh<10>1  (
    .ADR0(DLX_EXinst_N73464),
    .ADR1(DLX_EXinst_N72938),
    .ADR2(DLX_IDinst_Imm_0_1),
    .ADR3(VCC),
    .O(\DLX_IDinst_RegFile_2_13/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0021_Sh<46>_SW0 .INIT = 16'hFC0C;
  X_LUT4 \DLX_EXinst_Mshift__n0021_Sh<46>_SW0  (
    .ADR0(VCC),
    .ADR1(\DLX_EXinst_Mshift__n0021_Sh[14] ),
    .ADR2(DLX_IDinst_Imm_2_1),
    .ADR3(\DLX_EXinst_Mshift__n0021_Sh[10] ),
    .O(\DLX_IDinst_RegFile_2_13/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_2_13/XUSED  (
    .I(\DLX_IDinst_RegFile_2_13/FROM ),
    .O(\DLX_EXinst_Mshift__n0021_Sh[10] )
  );
  X_BUF \DLX_IDinst_RegFile_2_13/YUSED  (
    .I(\DLX_IDinst_RegFile_2_13/GROM ),
    .O(N130311)
  );
  defparam \DLX_EXinst_Mshift__n0021_Sh<11>1 .INIT = 16'hBB88;
  X_LUT4 \DLX_EXinst_Mshift__n0021_Sh<11>1  (
    .ADR0(DLX_EXinst_N73464),
    .ADR1(DLX_IDinst_Imm_0_1),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N72943),
    .O(\DLX_IDinst_RegFile_1_1/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0021_Sh<47>_SW0 .INIT = 16'hFA0A;
  X_LUT4 \DLX_EXinst_Mshift__n0021_Sh<47>_SW0  (
    .ADR0(\DLX_EXinst_Mshift__n0021_Sh[15] ),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_Imm_2_1),
    .ADR3(\DLX_EXinst_Mshift__n0021_Sh[11] ),
    .O(\DLX_IDinst_RegFile_1_1/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_1_1/XUSED  (
    .I(\DLX_IDinst_RegFile_1_1/FROM ),
    .O(\DLX_EXinst_Mshift__n0021_Sh[11] )
  );
  X_BUF \DLX_IDinst_RegFile_1_1/YUSED  (
    .I(\DLX_IDinst_RegFile_1_1/GROM ),
    .O(N130415)
  );
  defparam DLX_IDinst_RegFile_11_21_482.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_11_21_482 (
    .I(DLX_IDinst_WB_data_eff[21]),
    .CE(DLX_IDinst__n0572),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_11_21)
  );
  defparam \DLX_EXinst_Mshift__n0021_Sh<24>1 .INIT = 16'hCCAA;
  X_LUT4 \DLX_EXinst_Mshift__n0021_Sh<24>1  (
    .ADR0(DLX_EXinst_N73499),
    .ADR1(DLX_EXinst_N72973),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_Imm_0_1),
    .O(\DLX_IDinst_RegFile_11_21/FROM )
  );
  defparam \DLX_EXinst__n0007<24>356 .INIT = 16'h2320;
  X_LUT4 \DLX_EXinst__n0007<24>356  (
    .ADR0(\DLX_EXinst_Mshift__n0021_Sh[20] ),
    .ADR1(\DLX_IDinst_Imm[3] ),
    .ADR2(\DLX_IDinst_Imm[2] ),
    .ADR3(\DLX_EXinst_Mshift__n0021_Sh[24] ),
    .O(\DLX_IDinst_RegFile_11_21/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_11_21/XUSED  (
    .I(\DLX_IDinst_RegFile_11_21/FROM ),
    .O(\DLX_EXinst_Mshift__n0021_Sh[24] )
  );
  X_BUF \DLX_IDinst_RegFile_11_21/YUSED  (
    .I(\DLX_IDinst_RegFile_11_21/GROM ),
    .O(CHOICE5667)
  );
  defparam DLX_IDinst_RegFile_2_22_483.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_2_22_483 (
    .I(DLX_IDinst_WB_data_eff[22]),
    .CE(DLX_IDinst__n0554),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_2_22)
  );
  defparam \DLX_EXinst_Mshift__n0021_Sh<16>1 .INIT = 16'hDD88;
  X_LUT4 \DLX_EXinst_Mshift__n0021_Sh<16>1  (
    .ADR0(DLX_IDinst_Imm_0_1),
    .ADR1(DLX_EXinst_N72953),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N73479),
    .O(\DLX_IDinst_RegFile_2_22/FROM )
  );
  defparam DLX_EXinst_Ker753751.INIT = 16'hFC30;
  X_LUT4 DLX_EXinst_Ker753751 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_Imm_2_1),
    .ADR2(\DLX_EXinst_Mshift__n0021_Sh[20] ),
    .ADR3(\DLX_EXinst_Mshift__n0021_Sh[16] ),
    .O(\DLX_IDinst_RegFile_2_22/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_2_22/XUSED  (
    .I(\DLX_IDinst_RegFile_2_22/FROM ),
    .O(\DLX_EXinst_Mshift__n0021_Sh[16] )
  );
  X_BUF \DLX_IDinst_RegFile_2_22/YUSED  (
    .I(\DLX_IDinst_RegFile_2_22/GROM ),
    .O(DLX_EXinst_N75377)
  );
  defparam \DLX_EXinst_Mshift__n0021_Sh<19>1 .INIT = 16'hAFA0;
  X_LUT4 \DLX_EXinst_Mshift__n0021_Sh<19>1  (
    .ADR0(DLX_EXinst_N73484),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_Imm_0_1),
    .ADR3(DLX_EXinst_N72963),
    .O(\DLX_IDinst_RegFile_15_5/FROM )
  );
  defparam DLX_EXinst_Ker7445937.INIT = 16'hFCCC;
  X_LUT4 DLX_EXinst_Ker7445937 (
    .ADR0(VCC),
    .ADR1(CHOICE1727),
    .ADR2(\DLX_IDinst_Imm[3] ),
    .ADR3(\DLX_EXinst_Mshift__n0021_Sh[19] ),
    .O(\DLX_IDinst_RegFile_15_5/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_15_5/XUSED  (
    .I(\DLX_IDinst_RegFile_15_5/FROM ),
    .O(\DLX_EXinst_Mshift__n0021_Sh[19] )
  );
  X_BUF \DLX_IDinst_RegFile_15_5/YUSED  (
    .I(\DLX_IDinst_RegFile_15_5/GROM ),
    .O(N137282)
  );
  defparam \DLX_EXinst_Mshift__n0022_Sh<12>1 .INIT = 16'hCCAA;
  X_LUT4 \DLX_EXinst_Mshift__n0022_Sh<12>1  (
    .ADR0(DLX_EXinst_N73519),
    .ADR1(DLX_EXinst_N73128),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_Imm_0_1),
    .O(\DLX_IFinst_IR_previous<13>/FROM )
  );
  defparam DLX_EXinst_Ker7467437.INIT = 16'hFCCC;
  X_LUT4 DLX_EXinst_Ker7467437 (
    .ADR0(VCC),
    .ADR1(CHOICE1791),
    .ADR2(DLX_IDinst_Imm_3_1),
    .ADR3(\DLX_EXinst_Mshift__n0022_Sh[12] ),
    .O(\DLX_IFinst_IR_previous<13>/GROM )
  );
  X_BUF \DLX_IFinst_IR_previous<13>/XUSED  (
    .I(\DLX_IFinst_IR_previous<13>/FROM ),
    .O(\DLX_EXinst_Mshift__n0022_Sh[12] )
  );
  X_BUF \DLX_IFinst_IR_previous<13>/YUSED  (
    .I(\DLX_IFinst_IR_previous<13>/GROM ),
    .O(N137680)
  );
  defparam \DLX_EXinst_Mshift__n0022_Sh<30>1 .INIT = 16'h0C0A;
  X_LUT4 \DLX_EXinst_Mshift__n0022_Sh<30>1  (
    .ADR0(DLX_IDinst_reg_out_A[30]),
    .ADR1(DLX_IDinst_reg_out_A[31]),
    .ADR2(DLX_IDinst_Imm_1_1),
    .ADR3(DLX_IDinst_Imm_0_1),
    .O(\DLX_EXinst_reg_out_B_EX<7>/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0022_Sh<58>1 .INIT = 16'h0E04;
  X_LUT4 \DLX_EXinst_Mshift__n0022_Sh<58>1  (
    .ADR0(DLX_IDinst_Imm_2_1),
    .ADR1(\DLX_EXinst_Mshift__n0020_Sh[26] ),
    .ADR2(DLX_IDinst_Imm_3_1),
    .ADR3(\DLX_EXinst_Mshift__n0022_Sh[30] ),
    .O(\DLX_EXinst_reg_out_B_EX<7>/GROM )
  );
  X_BUF \DLX_EXinst_reg_out_B_EX<7>/XUSED  (
    .I(\DLX_EXinst_reg_out_B_EX<7>/FROM ),
    .O(\DLX_EXinst_Mshift__n0022_Sh[30] )
  );
  X_BUF \DLX_EXinst_reg_out_B_EX<7>/YUSED  (
    .I(\DLX_EXinst_reg_out_B_EX<7>/GROM ),
    .O(\DLX_EXinst_Mshift__n0022_Sh[58] )
  );
  defparam DLX_IDinst_RegFile_2_23_484.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_2_23_484 (
    .I(DLX_IDinst_WB_data_eff[23]),
    .CE(DLX_IDinst__n0554),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_2_23)
  );
  defparam \DLX_EXinst_Mshift__n0022_Sh<22>1 .INIT = 16'hEE44;
  X_LUT4 \DLX_EXinst_Mshift__n0022_Sh<22>1  (
    .ADR0(DLX_IDinst_Imm_0_1),
    .ADR1(DLX_EXinst_N73544),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N73153),
    .O(\DLX_IDinst_RegFile_2_23/FROM )
  );
  defparam DLX_EXinst_Ker731611.INIT = 16'hBB88;
  X_LUT4 DLX_EXinst_Ker731611 (
    .ADR0(\DLX_EXinst_Mshift__n0022_Sh[30] ),
    .ADR1(\DLX_IDinst_Imm[3] ),
    .ADR2(VCC),
    .ADR3(\DLX_EXinst_Mshift__n0022_Sh[22] ),
    .O(\DLX_IDinst_RegFile_2_23/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_2_23/XUSED  (
    .I(\DLX_IDinst_RegFile_2_23/FROM ),
    .O(\DLX_EXinst_Mshift__n0022_Sh[22] )
  );
  X_BUF \DLX_IDinst_RegFile_2_23/YUSED  (
    .I(\DLX_IDinst_RegFile_2_23/GROM ),
    .O(DLX_EXinst_N73163)
  );
  defparam DLX_IDinst_RegFile_18_23_485.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_18_23_485 (
    .I(DLX_IDinst_WB_data_eff[23]),
    .CE(DLX_IDinst__n0586),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_18_23)
  );
  defparam \DLX_EXinst_Mshift__n0022_Sh<23>1 .INIT = 16'hDD88;
  X_LUT4 \DLX_EXinst_Mshift__n0022_Sh<23>1  (
    .ADR0(DLX_IDinst_Imm_0_1),
    .ADR1(DLX_EXinst_N73897),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N73153),
    .O(\DLX_IDinst_RegFile_2_15/FROM )
  );
  defparam DLX_EXinst_Ker731661.INIT = 16'h7340;
  X_LUT4 DLX_EXinst_Ker731661 (
    .ADR0(DLX_EXinst_N73211),
    .ADR1(\DLX_IDinst_Imm[3] ),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(\DLX_EXinst_Mshift__n0022_Sh[23] ),
    .O(\DLX_IDinst_RegFile_2_15/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_2_15/XUSED  (
    .I(\DLX_IDinst_RegFile_2_15/FROM ),
    .O(\DLX_EXinst_Mshift__n0022_Sh[23] )
  );
  X_BUF \DLX_IDinst_RegFile_2_15/YUSED  (
    .I(\DLX_IDinst_RegFile_2_15/GROM ),
    .O(DLX_EXinst_N73168)
  );
  defparam \DLX_EXinst_Mshift__n0022_Sh<16>1 .INIT = 16'hFA0A;
  X_LUT4 \DLX_EXinst_Mshift__n0022_Sh<16>1  (
    .ADR0(DLX_EXinst_N73529),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_Imm_0_1),
    .ADR3(DLX_EXinst_N73138),
    .O(\DLX_IDinst_RegFile_0_12/FROM )
  );
  defparam DLX_EXinst_Ker749441.INIT = 16'hFA50;
  X_LUT4 DLX_EXinst_Ker749441 (
    .ADR0(DLX_IDinst_Imm_3_1),
    .ADR1(VCC),
    .ADR2(\DLX_EXinst_Mshift__n0022_Sh[8] ),
    .ADR3(\DLX_EXinst_Mshift__n0022_Sh[16] ),
    .O(\DLX_IDinst_RegFile_0_12/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_0_12/XUSED  (
    .I(\DLX_IDinst_RegFile_0_12/FROM ),
    .O(\DLX_EXinst_Mshift__n0022_Sh[16] )
  );
  X_BUF \DLX_IDinst_RegFile_0_12/YUSED  (
    .I(\DLX_IDinst_RegFile_0_12/GROM ),
    .O(DLX_EXinst_N74946)
  );
  defparam DLX_IDinst_RegFile_23_30_486.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_23_30_486 (
    .I(DLX_IDinst_WB_data_eff[30]),
    .CE(DLX_IDinst__n0596),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_23_30)
  );
  defparam \DLX_EXinst_Mshift__n0022_Sh<17>1 .INIT = 16'hF0CC;
  X_LUT4 \DLX_EXinst_Mshift__n0022_Sh<17>1  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N73138),
    .ADR2(DLX_EXinst_N73534),
    .ADR3(DLX_IDinst_Imm_0_1),
    .O(\DLX_IDinst_RegFile_23_30/FROM )
  );
  defparam DLX_EXinst_Ker749791.INIT = 16'hBB88;
  X_LUT4 DLX_EXinst_Ker749791 (
    .ADR0(\DLX_EXinst_Mshift__n0020_Sh[25] ),
    .ADR1(DLX_IDinst_Imm_3_1),
    .ADR2(VCC),
    .ADR3(\DLX_EXinst_Mshift__n0022_Sh[17] ),
    .O(\DLX_IDinst_RegFile_23_30/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_23_30/XUSED  (
    .I(\DLX_IDinst_RegFile_23_30/FROM ),
    .O(\DLX_EXinst_Mshift__n0022_Sh[17] )
  );
  X_BUF \DLX_IDinst_RegFile_23_30/YUSED  (
    .I(\DLX_IDinst_RegFile_23_30/GROM ),
    .O(DLX_EXinst_N74981)
  );
  defparam DLX_IDinst_RegFile_2_24_487.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_2_24_487 (
    .I(DLX_IDinst_WB_data_eff[24]),
    .CE(DLX_IDinst__n0554),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_2_24)
  );
  defparam \DLX_EXinst_Mshift__n0022_Sh<50>1 .INIT = 16'hF5A0;
  X_LUT4 \DLX_EXinst_Mshift__n0022_Sh<50>1  (
    .ADR0(DLX_IDinst_Imm_2_1),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N73163),
    .ADR3(DLX_EXinst_N74986),
    .O(\DLX_IDinst_RegFile_2_24/FROM )
  );
  defparam \DLX_EXinst__n0007<18>109_SW0 .INIT = 16'hFAAA;
  X_LUT4 \DLX_EXinst__n0007<18>109_SW0  (
    .ADR0(CHOICE5220),
    .ADR1(VCC),
    .ADR2(DLX_EXinst__n0056),
    .ADR3(\DLX_EXinst_Mshift__n0022_Sh[50] ),
    .O(\DLX_IDinst_RegFile_2_24/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_2_24/XUSED  (
    .I(\DLX_IDinst_RegFile_2_24/FROM ),
    .O(\DLX_EXinst_Mshift__n0022_Sh[50] )
  );
  X_BUF \DLX_IDinst_RegFile_2_24/YUSED  (
    .I(\DLX_IDinst_RegFile_2_24/GROM ),
    .O(N163424)
  );
  defparam \DLX_EXinst_Mshift__n0022_Sh<18>1 .INIT = 16'hEE44;
  X_LUT4 \DLX_EXinst_Mshift__n0022_Sh<18>1  (
    .ADR0(DLX_IDinst_Imm_0_1),
    .ADR1(DLX_EXinst_N73534),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N73143),
    .O(\DLX_IDinst_RegFile_2_16/FROM )
  );
  defparam DLX_EXinst_Ker749841.INIT = 16'hCFC0;
  X_LUT4 DLX_EXinst_Ker749841 (
    .ADR0(VCC),
    .ADR1(\DLX_EXinst_Mshift__n0020_Sh[26] ),
    .ADR2(DLX_IDinst_Imm_3_1),
    .ADR3(\DLX_EXinst_Mshift__n0022_Sh[18] ),
    .O(\DLX_IDinst_RegFile_2_16/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_2_16/XUSED  (
    .I(\DLX_IDinst_RegFile_2_16/FROM ),
    .O(\DLX_EXinst_Mshift__n0022_Sh[18] )
  );
  X_BUF \DLX_IDinst_RegFile_2_16/YUSED  (
    .I(\DLX_IDinst_RegFile_2_16/GROM ),
    .O(DLX_EXinst_N74986)
  );
  defparam DLX_IDinst_RegFile_26_23_488.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_26_23_488 (
    .I(DLX_IDinst_WB_data_eff[23]),
    .CE(DLX_IDinst__n0602),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_26_23)
  );
  defparam \DLX_EXinst_Mshift__n0022_Sh<51>1 .INIT = 16'hFA0A;
  X_LUT4 \DLX_EXinst_Mshift__n0022_Sh<51>1  (
    .ADR0(DLX_EXinst_N75352),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_Imm_2_1),
    .ADR3(DLX_EXinst_N73168),
    .O(\DLX_IDinst_RegFile_16_15/FROM )
  );
  defparam \DLX_EXinst__n0007<19>109_SW0 .INIT = 16'hFCCC;
  X_LUT4 \DLX_EXinst__n0007<19>109_SW0  (
    .ADR0(VCC),
    .ADR1(CHOICE5299),
    .ADR2(DLX_EXinst__n0056),
    .ADR3(\DLX_EXinst_Mshift__n0022_Sh[51] ),
    .O(\DLX_IDinst_RegFile_16_15/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_16_15/XUSED  (
    .I(\DLX_IDinst_RegFile_16_15/FROM ),
    .O(\DLX_EXinst_Mshift__n0022_Sh[51] )
  );
  X_BUF \DLX_IDinst_RegFile_16_15/YUSED  (
    .I(\DLX_IDinst_RegFile_16_15/GROM ),
    .O(N163558)
  );
  defparam \DLX_EXinst_Mshift__n0022_Sh<57>1 .INIT = 16'h00E2;
  X_LUT4 \DLX_EXinst_Mshift__n0022_Sh<57>1  (
    .ADR0(\DLX_EXinst_Mshift__n0020_Sh[25] ),
    .ADR1(DLX_IDinst_Imm_2_1),
    .ADR2(\DLX_EXinst_Mshift__n0022_Sh[29] ),
    .ADR3(DLX_IDinst_Imm_3_1),
    .O(\DLX_IDinst_RegFile_2_17/FROM )
  );
  defparam \DLX_EXinst__n0007<25>75_SW0 .INIT = 16'hEEAA;
  X_LUT4 \DLX_EXinst__n0007<25>75_SW0  (
    .ADR0(CHOICE5076),
    .ADR1(DLX_EXinst__n0056),
    .ADR2(VCC),
    .ADR3(\DLX_EXinst_Mshift__n0022_Sh[57] ),
    .O(\DLX_IDinst_RegFile_2_17/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_2_17/XUSED  (
    .I(\DLX_IDinst_RegFile_2_17/FROM ),
    .O(\DLX_EXinst_Mshift__n0022_Sh[57] )
  );
  X_BUF \DLX_IDinst_RegFile_2_17/YUSED  (
    .I(\DLX_IDinst_RegFile_2_17/GROM ),
    .O(N163610)
  );
  defparam \DLX_EXinst_Mshift__n0022_Sh<49>1 .INIT = 16'hF3C0;
  X_LUT4 \DLX_EXinst_Mshift__n0022_Sh<49>1  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_Imm_2_1),
    .ADR2(DLX_EXinst_N73158),
    .ADR3(DLX_EXinst_N74981),
    .O(\DLX_IDinst_RegFile_22_6/FROM )
  );
  defparam \DLX_EXinst__n0007<17>109_SW0 .INIT = 16'hEECC;
  X_LUT4 \DLX_EXinst__n0007<17>109_SW0  (
    .ADR0(DLX_EXinst__n0056),
    .ADR1(CHOICE5378),
    .ADR2(VCC),
    .ADR3(\DLX_EXinst_Mshift__n0022_Sh[49] ),
    .O(\DLX_IDinst_RegFile_22_6/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_22_6/XUSED  (
    .I(\DLX_IDinst_RegFile_22_6/FROM ),
    .O(\DLX_EXinst_Mshift__n0022_Sh[49] )
  );
  X_BUF \DLX_IDinst_RegFile_22_6/YUSED  (
    .I(\DLX_IDinst_RegFile_22_6/GROM ),
    .O(N163635)
  );
  defparam DLX_IDinst__n01175.INIT = 16'hF080;
  X_LUT4 DLX_IDinst__n01175 (
    .ADR0(DLX_IDinst_N108465),
    .ADR1(DLX_IDinst_N108152),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(DLX_IDinst_N107405),
    .O(\DLX_IDinst_RegFile_1_23/FROM )
  );
  defparam DLX_IDinst_Ker10720631_SW0.INIT = 16'hF8F8;
  X_LUT4 DLX_IDinst_Ker10720631_SW0 (
    .ADR0(DLX_IDinst_N108465),
    .ADR1(DLX_IDinst_N108152),
    .ADR2(DLX_IDinst_N107405),
    .ADR3(VCC),
    .O(\DLX_IDinst_RegFile_1_23/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_1_23/XUSED  (
    .I(\DLX_IDinst_RegFile_1_23/FROM ),
    .O(CHOICE3348)
  );
  X_BUF \DLX_IDinst_RegFile_1_23/YUSED  (
    .I(\DLX_IDinst_RegFile_1_23/GROM ),
    .O(N163562)
  );
  defparam \DLX_EXinst_Mshift__n0020_Sh<127>1 .INIT = 16'h0100;
  X_LUT4 \DLX_EXinst_Mshift__n0020_Sh<127>1  (
    .ADR0(DLX_IDinst_Imm_1_1),
    .ADR1(DLX_EXinst_N72815),
    .ADR2(DLX_IDinst_Imm_0_1),
    .ADR3(DLX_IDinst_reg_out_A[31]),
    .O(\DLX_MEMinst_opcode_of_WB<5>/FROM )
  );
  defparam \DLX_EXinst__n0007<15>199 .INIT = 16'hA800;
  X_LUT4 \DLX_EXinst__n0007<15>199  (
    .ADR0(\DLX_IDinst_Imm[4] ),
    .ADR1(DLX_EXinst_N76441),
    .ADR2(DLX_EXinst_N76124),
    .ADR3(\DLX_EXinst_Mshift__n0020_Sh[127] ),
    .O(\DLX_MEMinst_opcode_of_WB<5>/GROM )
  );
  X_BUF \DLX_MEMinst_opcode_of_WB<5>/XUSED  (
    .I(\DLX_MEMinst_opcode_of_WB<5>/FROM ),
    .O(\DLX_EXinst_Mshift__n0020_Sh[127] )
  );
  X_BUF \DLX_MEMinst_opcode_of_WB<5>/YUSED  (
    .I(\DLX_MEMinst_opcode_of_WB<5>/GROM ),
    .O(CHOICE4308)
  );
  defparam DLX_IDinst_RegFile_11_24_489.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_11_24_489 (
    .I(DLX_IDinst_WB_data_eff[24]),
    .CE(DLX_IDinst__n0572),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_11_24)
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<24>1 .INIT = 16'hDD88;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<24>1  (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(DLX_EXinst_N72888),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N73594),
    .O(\DLX_IDinst_RegFile_11_24/FROM )
  );
  defparam \DLX_EXinst__n0007<24>119 .INIT = 16'h0D08;
  X_LUT4 \DLX_EXinst__n0007<24>119  (
    .ADR0(DLX_IDinst_reg_out_B[2]),
    .ADR1(\DLX_EXinst_Mshift__n0023_Sh[20] ),
    .ADR2(DLX_IDinst_reg_out_B[3]),
    .ADR3(\DLX_EXinst_Mshift__n0023_Sh[24] ),
    .O(\DLX_IDinst_RegFile_11_24/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_11_24/XUSED  (
    .I(\DLX_IDinst_RegFile_11_24/FROM ),
    .O(\DLX_EXinst_Mshift__n0023_Sh[24] )
  );
  X_BUF \DLX_IDinst_RegFile_11_24/YUSED  (
    .I(\DLX_IDinst_RegFile_11_24/GROM ),
    .O(CHOICE5617)
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<16>1 .INIT = 16'hAACC;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<16>1  (
    .ADR0(DLX_EXinst_N72868),
    .ADR1(DLX_EXinst_N73574),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[0]),
    .O(\DLX_IDinst_RegFile_6_6/FROM )
  );
  defparam DLX_EXinst_Ker750041.INIT = 16'hFC0C;
  X_LUT4 DLX_EXinst_Ker750041 (
    .ADR0(VCC),
    .ADR1(\DLX_EXinst_Mshift__n0023_Sh[20] ),
    .ADR2(DLX_IDinst_reg_out_B_2_1),
    .ADR3(\DLX_EXinst_Mshift__n0023_Sh[16] ),
    .O(\DLX_IDinst_RegFile_6_6/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_6_6/XUSED  (
    .I(\DLX_IDinst_RegFile_6_6/FROM ),
    .O(\DLX_EXinst_Mshift__n0023_Sh[16] )
  );
  X_BUF \DLX_IDinst_RegFile_6_6/YUSED  (
    .I(\DLX_IDinst_RegFile_6_6/GROM ),
    .O(DLX_EXinst_N75006)
  );
  defparam DLX_IFinst_PC_28.INIT = 1'b0;
  X_SFF DLX_IFinst_PC_28 (
    .I(DLX_IFinst_NPC[28]),
    .CE(DLX_IFinst_PC_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_IFinst_PC[28])
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<19>1 .INIT = 16'hB8B8;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<19>1  (
    .ADR0(DLX_EXinst_N73579),
    .ADR1(DLX_IDinst_reg_out_B[0]),
    .ADR2(DLX_EXinst_N72878),
    .ADR3(VCC),
    .O(\DLX_IFinst_PC<28>/FROM )
  );
  defparam DLX_EXinst_Ker7422637.INIT = 16'hFAAA;
  X_LUT4 DLX_EXinst_Ker7422637 (
    .ADR0(CHOICE1765),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[3]),
    .ADR3(\DLX_EXinst_Mshift__n0023_Sh[19] ),
    .O(\DLX_IFinst_PC<28>/GROM )
  );
  X_BUF \DLX_IFinst_PC<28>/XUSED  (
    .I(\DLX_IFinst_PC<28>/FROM ),
    .O(\DLX_EXinst_Mshift__n0023_Sh[19] )
  );
  X_BUF \DLX_IFinst_PC<28>/YUSED  (
    .I(\DLX_IFinst_PC<28>/GROM ),
    .O(N137518)
  );
  defparam DLX_EXinst_Ker764991.INIT = 16'h00F0;
  X_LUT4 DLX_EXinst_Ker764991 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[1]),
    .ADR3(DLX_IDinst_reg_out_B[0]),
    .O(\DLX_IDinst_RegFile_15_9/FROM )
  );
  defparam \DLX_EXinst__n0013<0>1 .INIT = 16'hFC0C;
  X_LUT4 \DLX_EXinst__n0013<0>1  (
    .ADR0(VCC),
    .ADR1(\DLX_IDinst_Imm[0] ),
    .ADR2(DLX_EXinst__n0036),
    .ADR3(DLX_IDinst_reg_out_B[0]),
    .O(\DLX_IDinst_RegFile_15_9/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_15_9/XUSED  (
    .I(\DLX_IDinst_RegFile_15_9/FROM ),
    .O(DLX_EXinst_N76501)
  );
  X_BUF \DLX_IDinst_RegFile_15_9/YUSED  (
    .I(\DLX_IDinst_RegFile_15_9/GROM ),
    .O(DLX_EXinst__n0013[0])
  );
  defparam DLX_IDinst_RegFile_1_26_490.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_1_26_490 (
    .I(DLX_IDinst_WB_data_eff[26]),
    .CE(DLX_IDinst__n0552),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_1_26)
  );
  defparam \DLX_IDinst__n0114<10>20 .INIT = 16'hE400;
  X_LUT4 \DLX_IDinst__n0114<10>20  (
    .ADR0(DLX_IDinst__n0175),
    .ADR1(DLX_IDinst__n0620[10]),
    .ADR2(DLX_MEMinst_RF_data_in[10]),
    .ADR3(DLX_IDinst_N107837),
    .O(\DLX_IDinst_RegFile_1_26/FROM )
  );
  defparam \DLX_IDinst_Mmux_regA_eff_Result<10>1 .INIT = 16'hAACC;
  X_LUT4 \DLX_IDinst_Mmux_regA_eff_Result<10>1  (
    .ADR0(DLX_MEMinst_RF_data_in[10]),
    .ADR1(DLX_IDinst__n0620[10]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst__n0175),
    .O(\DLX_IDinst_RegFile_1_26/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_1_26/XUSED  (
    .I(\DLX_IDinst_RegFile_1_26/FROM ),
    .O(CHOICE2235)
  );
  X_BUF \DLX_IDinst_RegFile_1_26/YUSED  (
    .I(\DLX_IDinst_RegFile_1_26/GROM ),
    .O(\DLX_IDinst_regA_eff[10] )
  );
  defparam \DLX_EXinst_Mshift__n0019_Sh<23>_SW0 .INIT = 16'hF5A0;
  X_LUT4 \DLX_EXinst_Mshift__n0019_Sh<23>_SW0  (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[26]),
    .ADR3(DLX_IDinst_reg_out_A[24]),
    .O(\DLX_IFinst_IR_previous<6>/FROM )
  );
  defparam \DLX_EXinst__n0013<1>1 .INIT = 16'hAFA0;
  X_LUT4 \DLX_EXinst__n0013<1>1  (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst__n0036),
    .ADR3(\DLX_IDinst_Imm[1] ),
    .O(\DLX_IFinst_IR_previous<6>/GROM )
  );
  X_BUF \DLX_IFinst_IR_previous<6>/XUSED  (
    .I(\DLX_IFinst_IR_previous<6>/FROM ),
    .O(N130927)
  );
  X_BUF \DLX_IFinst_IR_previous<6>/YUSED  (
    .I(\DLX_IFinst_IR_previous<6>/GROM ),
    .O(DLX_EXinst__n0013[1])
  );
  defparam DLX_IDinst_RegFile_26_2_491.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_26_2_491 (
    .I(DLX_MEMinst_RF_data_in[2]),
    .CE(DLX_IDinst__n0602),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_26_2)
  );
  defparam \DLX_IDinst__n0114<11>20 .INIT = 16'h88A0;
  X_LUT4 \DLX_IDinst__n0114<11>20  (
    .ADR0(DLX_IDinst_N107837),
    .ADR1(DLX_MEMinst_RF_data_in[11]),
    .ADR2(DLX_IDinst__n0620[11]),
    .ADR3(DLX_IDinst__n0175),
    .O(\DLX_IDinst_RegFile_26_2/FROM )
  );
  defparam \DLX_IDinst_Mmux_regA_eff_Result<11>1 .INIT = 16'hFA0A;
  X_LUT4 \DLX_IDinst_Mmux_regA_eff_Result<11>1  (
    .ADR0(DLX_IDinst__n0620[11]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst__n0175),
    .ADR3(DLX_MEMinst_RF_data_in[11]),
    .O(\DLX_IDinst_RegFile_26_2/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_26_2/XUSED  (
    .I(\DLX_IDinst_RegFile_26_2/FROM ),
    .O(CHOICE2246)
  );
  X_BUF \DLX_IDinst_RegFile_26_2/YUSED  (
    .I(\DLX_IDinst_RegFile_26_2/GROM ),
    .O(\DLX_IDinst_regA_eff[11] )
  );
  defparam DLX_IDinst_RegFile_22_13_492.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_22_13_492 (
    .I(DLX_IDinst_WB_data_eff[13]),
    .CE(DLX_IDinst__n0594),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_22_13)
  );
  defparam DLX_EXinst_Ker729061.INIT = 16'hD8D8;
  X_LUT4 DLX_EXinst_Ker729061 (
    .ADR0(DLX_IDinst_reg_out_B[2]),
    .ADR1(\DLX_EXinst_Mshift__n0023_Sh[2] ),
    .ADR2(\DLX_EXinst_Mshift__n0023_Sh[6] ),
    .ADR3(VCC),
    .O(\DLX_IDinst_RegFile_22_13/FROM )
  );
  defparam \DLX_EXinst__n0013<2>1 .INIT = 16'hAACC;
  X_LUT4 \DLX_EXinst__n0013<2>1  (
    .ADR0(DLX_IDinst_reg_out_B[2]),
    .ADR1(\DLX_IDinst_Imm[2] ),
    .ADR2(VCC),
    .ADR3(DLX_EXinst__n0036),
    .O(\DLX_IDinst_RegFile_22_13/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_22_13/XUSED  (
    .I(\DLX_IDinst_RegFile_22_13/FROM ),
    .O(DLX_EXinst_N72908)
  );
  X_BUF \DLX_IDinst_RegFile_22_13/YUSED  (
    .I(\DLX_IDinst_RegFile_22_13/GROM ),
    .O(DLX_EXinst__n0013[2])
  );
  defparam \DLX_IDinst__n0114<12>20 .INIT = 16'hA820;
  X_LUT4 \DLX_IDinst__n0114<12>20  (
    .ADR0(DLX_IDinst_N107837),
    .ADR1(DLX_IDinst__n0175),
    .ADR2(DLX_IDinst__n0620[12]),
    .ADR3(DLX_MEMinst_RF_data_in[12]),
    .O(\DLX_IDinst_RegFile_30_23/FROM )
  );
  defparam \DLX_IDinst_Mmux_regA_eff_Result<12>1 .INIT = 16'hFA50;
  X_LUT4 \DLX_IDinst_Mmux_regA_eff_Result<12>1  (
    .ADR0(DLX_IDinst__n0175),
    .ADR1(VCC),
    .ADR2(DLX_IDinst__n0620[12]),
    .ADR3(DLX_MEMinst_RF_data_in[12]),
    .O(\DLX_IDinst_RegFile_30_23/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_30_23/XUSED  (
    .I(\DLX_IDinst_RegFile_30_23/FROM ),
    .O(CHOICE2257)
  );
  X_BUF \DLX_IDinst_RegFile_30_23/YUSED  (
    .I(\DLX_IDinst_RegFile_30_23/GROM ),
    .O(\DLX_IDinst_regA_eff[12] )
  );
  defparam \DLX_IDinst_Mmux_regA_eff_Result<20>1 .INIT = 16'hCCF0;
  X_LUT4 \DLX_IDinst_Mmux_regA_eff_Result<20>1  (
    .ADR0(VCC),
    .ADR1(DLX_MEMinst_RF_data_in[20]),
    .ADR2(DLX_IDinst__n0620[20]),
    .ADR3(DLX_IDinst__n0175),
    .O(\DLX_IDinst_RegFile_3_13/FROM )
  );
  defparam DLX_IDinst__n0177169.INIT = 16'h0001;
  X_LUT4 DLX_IDinst__n0177169 (
    .ADR0(\DLX_IDinst_regA_eff[19] ),
    .ADR1(\DLX_IDinst_regA_eff[18] ),
    .ADR2(\DLX_IDinst_regA_eff[17] ),
    .ADR3(\DLX_IDinst_regA_eff[20] ),
    .O(\DLX_IDinst_RegFile_3_13/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_3_13/XUSED  (
    .I(\DLX_IDinst_RegFile_3_13/FROM ),
    .O(\DLX_IDinst_regA_eff[20] )
  );
  X_BUF \DLX_IDinst_RegFile_3_13/YUSED  (
    .I(\DLX_IDinst_RegFile_3_13/GROM ),
    .O(CHOICE4240)
  );
  defparam DLX_IDinst_RegFile_3_21_493.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_3_21_493 (
    .I(DLX_IDinst_WB_data_eff[21]),
    .CE(DLX_IDinst__n0556),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_3_21)
  );
  defparam \DLX_EXinst__n0007<24>45_SW0 .INIT = 16'hFFAA;
  X_LUT4 \DLX_EXinst__n0007<24>45_SW0  (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[3]),
    .O(\DLX_IDinst_RegFile_3_21/FROM )
  );
  defparam \DLX_EXinst__n0013<3>1 .INIT = 16'hCFC0;
  X_LUT4 \DLX_EXinst__n0013<3>1  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_B[3]),
    .ADR2(DLX_EXinst__n0036),
    .ADR3(\DLX_IDinst_Imm[3] ),
    .O(\DLX_IDinst_RegFile_3_21/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_3_21/XUSED  (
    .I(\DLX_IDinst_RegFile_3_21/FROM ),
    .O(N163790)
  );
  X_BUF \DLX_IDinst_RegFile_3_21/YUSED  (
    .I(\DLX_IDinst_RegFile_3_21/GROM ),
    .O(DLX_EXinst__n0013[3])
  );
  defparam DLX_IDinst_RegFile_18_15_494.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_18_15_494 (
    .I(DLX_IDinst_WB_data_eff[15]),
    .CE(DLX_IDinst__n0586),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_18_15)
  );
  defparam \DLX_IDinst__n0114<13>20 .INIT = 16'hD080;
  X_LUT4 \DLX_IDinst__n0114<13>20  (
    .ADR0(DLX_IDinst__n0175),
    .ADR1(DLX_MEMinst_RF_data_in[13]),
    .ADR2(DLX_IDinst_N107837),
    .ADR3(DLX_IDinst__n0620[13]),
    .O(\DLX_IDinst_RegFile_2_29/FROM )
  );
  defparam \DLX_IDinst_Mmux_regA_eff_Result<13>1 .INIT = 16'hF5A0;
  X_LUT4 \DLX_IDinst_Mmux_regA_eff_Result<13>1  (
    .ADR0(DLX_IDinst__n0175),
    .ADR1(VCC),
    .ADR2(DLX_MEMinst_RF_data_in[13]),
    .ADR3(DLX_IDinst__n0620[13]),
    .O(\DLX_IDinst_RegFile_2_29/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_2_29/XUSED  (
    .I(\DLX_IDinst_RegFile_2_29/FROM ),
    .O(CHOICE2268)
  );
  X_BUF \DLX_IDinst_RegFile_2_29/YUSED  (
    .I(\DLX_IDinst_RegFile_2_29/GROM ),
    .O(\DLX_IDinst_regA_eff[13] )
  );
  defparam \DLX_IDinst__n0114<21>20 .INIT = 16'h88A0;
  X_LUT4 \DLX_IDinst__n0114<21>20  (
    .ADR0(DLX_IDinst_N107837),
    .ADR1(DLX_MEMinst_RF_data_in[21]),
    .ADR2(DLX_IDinst__n0620[21]),
    .ADR3(DLX_IDinst__n0175),
    .O(\DLX_IDinst_RegFile_23_23/FROM )
  );
  defparam \DLX_IDinst_Mmux_regA_eff_Result<21>1 .INIT = 16'hD8D8;
  X_LUT4 \DLX_IDinst_Mmux_regA_eff_Result<21>1  (
    .ADR0(DLX_IDinst__n0175),
    .ADR1(DLX_MEMinst_RF_data_in[21]),
    .ADR2(DLX_IDinst__n0620[21]),
    .ADR3(VCC),
    .O(\DLX_IDinst_RegFile_23_23/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_23_23/XUSED  (
    .I(\DLX_IDinst_RegFile_23_23/FROM ),
    .O(CHOICE2368)
  );
  X_BUF \DLX_IDinst_RegFile_23_23/YUSED  (
    .I(\DLX_IDinst_RegFile_23_23/GROM ),
    .O(\DLX_IDinst_regA_eff[21] )
  );
  defparam DLX_EXinst_Ker759621.INIT = 16'h0010;
  X_LUT4 DLX_EXinst_Ker759621 (
    .ADR0(DLX_IDinst_reg_out_B_2_1),
    .ADR1(DLX_IDinst_reg_out_B_3_1),
    .ADR2(DLX_EXinst__n0036),
    .ADR3(DLX_IDinst_reg_out_B[4]),
    .O(\DLX_IDinst_RegFile_3_22/FROM )
  );
  defparam \DLX_EXinst__n0013<4>1 .INIT = 16'hBB88;
  X_LUT4 \DLX_EXinst__n0013<4>1  (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(DLX_EXinst__n0036),
    .ADR2(VCC),
    .ADR3(\DLX_IDinst_Imm[4] ),
    .O(\DLX_IDinst_RegFile_3_22/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_3_22/XUSED  (
    .I(\DLX_IDinst_RegFile_3_22/FROM ),
    .O(DLX_EXinst_N75964)
  );
  X_BUF \DLX_IDinst_RegFile_3_22/YUSED  (
    .I(\DLX_IDinst_RegFile_3_22/GROM ),
    .O(DLX_EXinst__n0013[4])
  );
  defparam \DLX_IDinst__n0114<14>20 .INIT = 16'hA088;
  X_LUT4 \DLX_IDinst__n0114<14>20  (
    .ADR0(DLX_IDinst_N107837),
    .ADR1(DLX_IDinst__n0620[14]),
    .ADR2(DLX_MEMinst_RF_data_in[14]),
    .ADR3(DLX_IDinst__n0175),
    .O(\DLX_IDinst_RegFile_23_17/FROM )
  );
  defparam \DLX_IDinst_Mmux_regA_eff_Result<14>1 .INIT = 16'hF0CC;
  X_LUT4 \DLX_IDinst_Mmux_regA_eff_Result<14>1  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst__n0620[14]),
    .ADR2(DLX_MEMinst_RF_data_in[14]),
    .ADR3(DLX_IDinst__n0175),
    .O(\DLX_IDinst_RegFile_23_17/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_23_17/XUSED  (
    .I(\DLX_IDinst_RegFile_23_17/FROM ),
    .O(CHOICE2279)
  );
  X_BUF \DLX_IDinst_RegFile_23_17/YUSED  (
    .I(\DLX_IDinst_RegFile_23_17/GROM ),
    .O(\DLX_IDinst_regA_eff[14] )
  );
  defparam \DLX_IDinst__n0114<22>20 .INIT = 16'h8A80;
  X_LUT4 \DLX_IDinst__n0114<22>20  (
    .ADR0(DLX_IDinst_N107837),
    .ADR1(DLX_MEMinst_RF_data_in[22]),
    .ADR2(DLX_IDinst__n0175),
    .ADR3(DLX_IDinst__n0620[22]),
    .O(\DLX_IDinst_RegFile_18_4/FROM )
  );
  defparam \DLX_IDinst_Mmux_regA_eff_Result<22>1 .INIT = 16'hFC0C;
  X_LUT4 \DLX_IDinst_Mmux_regA_eff_Result<22>1  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst__n0620[22]),
    .ADR2(DLX_IDinst__n0175),
    .ADR3(DLX_MEMinst_RF_data_in[22]),
    .O(\DLX_IDinst_RegFile_18_4/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_18_4/XUSED  (
    .I(\DLX_IDinst_RegFile_18_4/FROM ),
    .O(CHOICE2379)
  );
  X_BUF \DLX_IDinst_RegFile_18_4/YUSED  (
    .I(\DLX_IDinst_RegFile_18_4/GROM ),
    .O(\DLX_IDinst_regA_eff[22] )
  );
  defparam DLX_IDinst_RegFile_3_15_495.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_3_15_495 (
    .I(DLX_IDinst_WB_data_eff[15]),
    .CE(DLX_IDinst__n0556),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_3_15)
  );
  defparam \DLX_IDinst__n0114<30>20 .INIT = 16'hE200;
  X_LUT4 \DLX_IDinst__n0114<30>20  (
    .ADR0(DLX_IDinst__n0620[30]),
    .ADR1(DLX_IDinst__n0175),
    .ADR2(DLX_MEMinst_RF_data_in[30]),
    .ADR3(DLX_IDinst_N107837),
    .O(\DLX_IDinst_RegFile_3_15/FROM )
  );
  defparam \DLX_IDinst_Mmux_regA_eff_Result<30>1 .INIT = 16'hFC0C;
  X_LUT4 \DLX_IDinst_Mmux_regA_eff_Result<30>1  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst__n0620[30]),
    .ADR2(DLX_IDinst__n0175),
    .ADR3(DLX_MEMinst_RF_data_in[30]),
    .O(\DLX_IDinst_RegFile_3_15/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_3_15/XUSED  (
    .I(\DLX_IDinst_RegFile_3_15/FROM ),
    .O(CHOICE2390)
  );
  X_BUF \DLX_IDinst_RegFile_3_15/YUSED  (
    .I(\DLX_IDinst_RegFile_3_15/GROM ),
    .O(\DLX_IDinst_regA_eff[30] )
  );
  defparam DLX_EXinst_Ker760321.INIT = 16'hF000;
  X_LUT4 DLX_EXinst_Ker760321 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(N148609),
    .ADR3(DLX_IDinst_reg_out_B[5]),
    .O(\DLX_IDinst_RegFile_17_18/FROM )
  );
  defparam \DLX_EXinst__n0013<5>1 .INIT = 16'hFC30;
  X_LUT4 \DLX_EXinst__n0013<5>1  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst__n0036),
    .ADR2(\DLX_IDinst_Imm[5] ),
    .ADR3(DLX_IDinst_reg_out_B[5]),
    .O(\DLX_IDinst_RegFile_17_18/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_17_18/XUSED  (
    .I(\DLX_IDinst_RegFile_17_18/FROM ),
    .O(DLX_EXinst_N76034)
  );
  X_BUF \DLX_IDinst_RegFile_17_18/YUSED  (
    .I(\DLX_IDinst_RegFile_17_18/GROM ),
    .O(DLX_EXinst__n0013[5])
  );
  defparam \DLX_IDinst__n0114<15>20 .INIT = 16'hB080;
  X_LUT4 \DLX_IDinst__n0114<15>20  (
    .ADR0(DLX_MEMinst_RF_data_in[15]),
    .ADR1(DLX_IDinst__n0175),
    .ADR2(DLX_IDinst_N107837),
    .ADR3(DLX_IDinst__n0620[15]),
    .O(\DLX_IDinst_RegFile_3_31/FROM )
  );
  defparam \DLX_IDinst_Mmux_regA_eff_Result<15>1 .INIT = 16'hB8B8;
  X_LUT4 \DLX_IDinst_Mmux_regA_eff_Result<15>1  (
    .ADR0(DLX_MEMinst_RF_data_in[15]),
    .ADR1(DLX_IDinst__n0175),
    .ADR2(DLX_IDinst__n0620[15]),
    .ADR3(VCC),
    .O(\DLX_IDinst_RegFile_3_31/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_3_31/XUSED  (
    .I(\DLX_IDinst_RegFile_3_31/FROM ),
    .O(CHOICE2290)
  );
  X_BUF \DLX_IDinst_RegFile_3_31/YUSED  (
    .I(\DLX_IDinst_RegFile_3_31/GROM ),
    .O(\DLX_IDinst_regA_eff[15] )
  );
  defparam \DLX_IDinst__n0114<23>20 .INIT = 16'hC840;
  X_LUT4 \DLX_IDinst__n0114<23>20  (
    .ADR0(DLX_IDinst__n0175),
    .ADR1(DLX_IDinst_N107837),
    .ADR2(DLX_IDinst__n0620[23]),
    .ADR3(DLX_MEMinst_RF_data_in[23]),
    .O(\DLX_IDinst_RegFile_29_7/FROM )
  );
  defparam \DLX_IDinst_Mmux_regA_eff_Result<23>1 .INIT = 16'hBB88;
  X_LUT4 \DLX_IDinst_Mmux_regA_eff_Result<23>1  (
    .ADR0(DLX_MEMinst_RF_data_in[23]),
    .ADR1(DLX_IDinst__n0175),
    .ADR2(VCC),
    .ADR3(DLX_IDinst__n0620[23]),
    .O(\DLX_IDinst_RegFile_29_7/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_29_7/XUSED  (
    .I(\DLX_IDinst_RegFile_29_7/FROM ),
    .O(CHOICE2467)
  );
  X_BUF \DLX_IDinst_RegFile_29_7/YUSED  (
    .I(\DLX_IDinst_RegFile_29_7/GROM ),
    .O(\DLX_IDinst_regA_eff[23] )
  );
  defparam \DLX_EXinst__n0013<9>1 .INIT = 16'hE2E2;
  X_LUT4 \DLX_EXinst__n0013<9>1  (
    .ADR0(\DLX_IDinst_Imm[9] ),
    .ADR1(DLX_EXinst__n0036),
    .ADR2(DLX_IDinst_reg_out_B[9]),
    .ADR3(VCC),
    .O(\DLX_IDinst_RegFile_1_0/FROM )
  );
  defparam \DLX_EXinst__n0013<6>1 .INIT = 16'hFC30;
  X_LUT4 \DLX_EXinst__n0013<6>1  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst__n0036),
    .ADR2(\DLX_IDinst_Imm[6] ),
    .ADR3(DLX_IDinst_reg_out_B[6]),
    .O(\DLX_IDinst_RegFile_1_0/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_1_0/XUSED  (
    .I(\DLX_IDinst_RegFile_1_0/FROM ),
    .O(DLX_EXinst__n0013[9])
  );
  X_BUF \DLX_IDinst_RegFile_1_0/YUSED  (
    .I(\DLX_IDinst_RegFile_1_0/GROM ),
    .O(DLX_EXinst__n0013[6])
  );
  defparam DLX_IDinst_RegFile_3_24_496.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_3_24_496 (
    .I(DLX_IDinst_WB_data_eff[24]),
    .CE(DLX_IDinst__n0556),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_3_24)
  );
  defparam \DLX_IDinst_Mmux_regA_eff_Result<16>1 .INIT = 16'hAFA0;
  X_LUT4 \DLX_IDinst_Mmux_regA_eff_Result<16>1  (
    .ADR0(DLX_MEMinst_RF_data_in[16]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst__n0175),
    .ADR3(DLX_IDinst__n0620[16]),
    .O(\DLX_IDinst_RegFile_3_24/FROM )
  );
  defparam DLX_IDinst__n0177156.INIT = 16'h0001;
  X_LUT4 DLX_IDinst__n0177156 (
    .ADR0(\DLX_IDinst_regA_eff[14] ),
    .ADR1(\DLX_IDinst_regA_eff[13] ),
    .ADR2(\DLX_IDinst_regA_eff[15] ),
    .ADR3(\DLX_IDinst_regA_eff[16] ),
    .O(\DLX_IDinst_RegFile_3_24/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_3_24/XUSED  (
    .I(\DLX_IDinst_RegFile_3_24/FROM ),
    .O(\DLX_IDinst_regA_eff[16] )
  );
  X_BUF \DLX_IDinst_RegFile_3_24/YUSED  (
    .I(\DLX_IDinst_RegFile_3_24/GROM ),
    .O(CHOICE4233)
  );
  defparam \DLX_IDinst_Mmux_regA_eff_Result<24>1 .INIT = 16'hF0AA;
  X_LUT4 \DLX_IDinst_Mmux_regA_eff_Result<24>1  (
    .ADR0(DLX_IDinst__n0620[24]),
    .ADR1(VCC),
    .ADR2(DLX_MEMinst_RF_data_in[24]),
    .ADR3(DLX_IDinst__n0175),
    .O(\DLX_IDinst_RegFile_3_17/FROM )
  );
  defparam DLX_IDinst__n0177193.INIT = 16'h0001;
  X_LUT4 DLX_IDinst__n0177193 (
    .ADR0(\DLX_IDinst_regA_eff[23] ),
    .ADR1(\DLX_IDinst_regA_eff[21] ),
    .ADR2(\DLX_IDinst_regA_eff[22] ),
    .ADR3(\DLX_IDinst_regA_eff[24] ),
    .O(\DLX_IDinst_RegFile_3_17/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_3_17/XUSED  (
    .I(\DLX_IDinst_RegFile_3_17/FROM ),
    .O(\DLX_IDinst_regA_eff[24] )
  );
  X_BUF \DLX_IDinst_RegFile_3_17/YUSED  (
    .I(\DLX_IDinst_RegFile_3_17/GROM ),
    .O(CHOICE4248)
  );
  defparam \DLX_EXinst__n0013<13>1 .INIT = 16'hEE44;
  X_LUT4 \DLX_EXinst__n0013<13>1  (
    .ADR0(DLX_EXinst__n0036),
    .ADR1(\DLX_IDinst_Imm[13] ),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[13]),
    .O(\DLX_IDinst_RegFile_3_25/FROM )
  );
  defparam \DLX_EXinst__n0013<7>1 .INIT = 16'hAFA0;
  X_LUT4 \DLX_EXinst__n0013<7>1  (
    .ADR0(DLX_IDinst_reg_out_B[7]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst__n0036),
    .ADR3(\DLX_IDinst_Imm[7] ),
    .O(\DLX_IDinst_RegFile_3_25/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_3_25/XUSED  (
    .I(\DLX_IDinst_RegFile_3_25/FROM ),
    .O(DLX_EXinst__n0013[13])
  );
  X_BUF \DLX_IDinst_RegFile_3_25/YUSED  (
    .I(\DLX_IDinst_RegFile_3_25/GROM ),
    .O(DLX_EXinst__n0013[7])
  );
  defparam \DLX_IDinst__n0114<17>20 .INIT = 16'hE400;
  X_LUT4 \DLX_IDinst__n0114<17>20  (
    .ADR0(DLX_IDinst__n0175),
    .ADR1(DLX_IDinst__n0620[17]),
    .ADR2(DLX_MEMinst_RF_data_in[17]),
    .ADR3(DLX_IDinst_N107837),
    .O(\CHOICE2324/FROM )
  );
  defparam \DLX_IDinst_Mmux_regA_eff_Result<17>1 .INIT = 16'hEE44;
  X_LUT4 \DLX_IDinst_Mmux_regA_eff_Result<17>1  (
    .ADR0(DLX_IDinst__n0175),
    .ADR1(DLX_IDinst__n0620[17]),
    .ADR2(VCC),
    .ADR3(DLX_MEMinst_RF_data_in[17]),
    .O(\CHOICE2324/GROM )
  );
  X_BUF \CHOICE2324/XUSED  (
    .I(\CHOICE2324/FROM ),
    .O(CHOICE2324)
  );
  X_BUF \CHOICE2324/YUSED  (
    .I(\CHOICE2324/GROM ),
    .O(\DLX_IDinst_regA_eff[17] )
  );
  defparam \DLX_IDinst__n0114<25>20 .INIT = 16'h88C0;
  X_LUT4 \DLX_IDinst__n0114<25>20  (
    .ADR0(DLX_MEMinst_RF_data_in[25]),
    .ADR1(DLX_IDinst_N107837),
    .ADR2(DLX_IDinst__n0620[25]),
    .ADR3(DLX_IDinst__n0175),
    .O(\CHOICE2445/FROM )
  );
  defparam \DLX_IDinst_Mmux_regA_eff_Result<25>1 .INIT = 16'hFC30;
  X_LUT4 \DLX_IDinst_Mmux_regA_eff_Result<25>1  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst__n0175),
    .ADR2(DLX_IDinst__n0620[25]),
    .ADR3(DLX_MEMinst_RF_data_in[25]),
    .O(\CHOICE2445/GROM )
  );
  X_BUF \CHOICE2445/XUSED  (
    .I(\CHOICE2445/FROM ),
    .O(CHOICE2445)
  );
  X_BUF \CHOICE2445/YUSED  (
    .I(\CHOICE2445/GROM ),
    .O(\DLX_IDinst_regA_eff[25] )
  );
  defparam \DLX_EXinst__n0013<10>1 .INIT = 16'hAAF0;
  X_LUT4 \DLX_EXinst__n0013<10>1  (
    .ADR0(DLX_IDinst_reg_out_B[10]),
    .ADR1(VCC),
    .ADR2(\DLX_IDinst_Imm[10] ),
    .ADR3(DLX_EXinst__n0036),
    .O(\DLX_EXinst__n0013<10>/FROM )
  );
  defparam \DLX_EXinst__n0013<8>1 .INIT = 16'hB8B8;
  X_LUT4 \DLX_EXinst__n0013<8>1  (
    .ADR0(DLX_IDinst_reg_out_B[8]),
    .ADR1(DLX_EXinst__n0036),
    .ADR2(\DLX_IDinst_Imm[8] ),
    .ADR3(VCC),
    .O(\DLX_EXinst__n0013<10>/GROM )
  );
  X_BUF \DLX_EXinst__n0013<10>/XUSED  (
    .I(\DLX_EXinst__n0013<10>/FROM ),
    .O(DLX_EXinst__n0013[10])
  );
  X_BUF \DLX_EXinst__n0013<10>/YUSED  (
    .I(\DLX_EXinst__n0013<10>/GROM ),
    .O(DLX_EXinst__n0013[8])
  );
  defparam \DLX_EXinst__n0007<31>28 .INIT = 16'hEAC0;
  X_LUT4 \DLX_EXinst__n0007<31>28  (
    .ADR0(N134884),
    .ADR1(DLX_EXinst__n0127),
    .ADR2(DLX_EXinst__n0012[31]),
    .ADR3(DLX_EXinst_ALU_result[31]),
    .O(\CHOICE5771/FROM )
  );
  defparam \DLX_EXinst__n0007<0>4 .INIT = 16'hF888;
  X_LUT4 \DLX_EXinst__n0007<0>4  (
    .ADR0(DLX_EXinst__n0127),
    .ADR1(DLX_EXinst__n0012[0]),
    .ADR2(N134884),
    .ADR3(DLX_EXinst_ALU_result[0]),
    .O(\CHOICE5771/GROM )
  );
  X_BUF \CHOICE5771/XUSED  (
    .I(\CHOICE5771/FROM ),
    .O(CHOICE5771)
  );
  X_BUF \CHOICE5771/YUSED  (
    .I(\CHOICE5771/GROM ),
    .O(CHOICE5871)
  );
  defparam \DLX_IDinst__n0114<18>20 .INIT = 16'hC480;
  X_LUT4 \DLX_IDinst__n0114<18>20  (
    .ADR0(DLX_IDinst__n0175),
    .ADR1(DLX_IDinst_N107837),
    .ADR2(DLX_MEMinst_RF_data_in[18]),
    .ADR3(DLX_IDinst__n0620[18]),
    .O(\CHOICE2335/FROM )
  );
  defparam \DLX_IDinst_Mmux_regA_eff_Result<18>1 .INIT = 16'hF3C0;
  X_LUT4 \DLX_IDinst_Mmux_regA_eff_Result<18>1  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst__n0175),
    .ADR2(DLX_MEMinst_RF_data_in[18]),
    .ADR3(DLX_IDinst__n0620[18]),
    .O(\CHOICE2335/GROM )
  );
  X_BUF \CHOICE2335/XUSED  (
    .I(\CHOICE2335/FROM ),
    .O(CHOICE2335)
  );
  X_BUF \CHOICE2335/YUSED  (
    .I(\CHOICE2335/GROM ),
    .O(\DLX_IDinst_regA_eff[18] )
  );
  defparam \DLX_IDinst__n0114<26>20 .INIT = 16'hC0A0;
  X_LUT4 \DLX_IDinst__n0114<26>20  (
    .ADR0(DLX_IDinst__n0620[26]),
    .ADR1(DLX_MEMinst_RF_data_in[26]),
    .ADR2(DLX_IDinst_N107837),
    .ADR3(DLX_IDinst__n0175),
    .O(\CHOICE2434/FROM )
  );
  defparam \DLX_IDinst_Mmux_regA_eff_Result<26>1 .INIT = 16'hAACC;
  X_LUT4 \DLX_IDinst_Mmux_regA_eff_Result<26>1  (
    .ADR0(DLX_MEMinst_RF_data_in[26]),
    .ADR1(DLX_IDinst__n0620[26]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst__n0175),
    .O(\CHOICE2434/GROM )
  );
  X_BUF \CHOICE2434/XUSED  (
    .I(\CHOICE2434/FROM ),
    .O(CHOICE2434)
  );
  X_BUF \CHOICE2434/YUSED  (
    .I(\CHOICE2434/GROM ),
    .O(\DLX_IDinst_regA_eff[26] )
  );
  defparam \DLX_IDinst__n0114<19>20 .INIT = 16'hE200;
  X_LUT4 \DLX_IDinst__n0114<19>20  (
    .ADR0(DLX_IDinst__n0620[19]),
    .ADR1(DLX_IDinst__n0175),
    .ADR2(DLX_MEMinst_RF_data_in[19]),
    .ADR3(DLX_IDinst_N107837),
    .O(\CHOICE2346/FROM )
  );
  defparam \DLX_IDinst_Mmux_regA_eff_Result<19>1 .INIT = 16'hFC0C;
  X_LUT4 \DLX_IDinst_Mmux_regA_eff_Result<19>1  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst__n0620[19]),
    .ADR2(DLX_IDinst__n0175),
    .ADR3(DLX_MEMinst_RF_data_in[19]),
    .O(\CHOICE2346/GROM )
  );
  X_BUF \CHOICE2346/XUSED  (
    .I(\CHOICE2346/FROM ),
    .O(CHOICE2346)
  );
  X_BUF \CHOICE2346/YUSED  (
    .I(\CHOICE2346/GROM ),
    .O(\DLX_IDinst_regA_eff[19] )
  );
  defparam \DLX_EXinst__n0007<2>7 .INIT = 16'h0400;
  X_LUT4 \DLX_EXinst__n0007<2>7  (
    .ADR0(\DLX_IDinst_Imm[2] ),
    .ADR1(\DLX_EXinst_Mshift__n0021_Sh[2] ),
    .ADR2(\DLX_IDinst_Imm[3] ),
    .ADR3(DLX_EXinst_N76463),
    .O(\CHOICE5511/FROM )
  );
  defparam \DLX_EXinst__n0007<1>7 .INIT = 16'h1000;
  X_LUT4 \DLX_EXinst__n0007<1>7  (
    .ADR0(\DLX_IDinst_Imm[2] ),
    .ADR1(\DLX_IDinst_Imm[3] ),
    .ADR2(\DLX_EXinst_Mshift__n0021_Sh[1] ),
    .ADR3(DLX_EXinst_N76463),
    .O(\CHOICE5511/GROM )
  );
  X_BUF \CHOICE5511/XUSED  (
    .I(\CHOICE5511/FROM ),
    .O(CHOICE5511)
  );
  X_BUF \CHOICE5511/YUSED  (
    .I(\CHOICE5511/GROM ),
    .O(CHOICE5690)
  );
  defparam \DLX_IDinst_Mmux_regA_eff_Result<28>1 .INIT = 16'hF0CC;
  X_LUT4 \DLX_IDinst_Mmux_regA_eff_Result<28>1  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst__n0620[28]),
    .ADR2(DLX_MEMinst_RF_data_in[28]),
    .ADR3(DLX_IDinst__n0175),
    .O(\DLX_IDinst_regA_eff<28>/FROM )
  );
  defparam DLX_IDinst__n0177206.INIT = 16'h0001;
  X_LUT4 DLX_IDinst__n0177206 (
    .ADR0(\DLX_IDinst_regA_eff[27] ),
    .ADR1(\DLX_IDinst_regA_eff[26] ),
    .ADR2(\DLX_IDinst_regA_eff[25] ),
    .ADR3(\DLX_IDinst_regA_eff[28] ),
    .O(\DLX_IDinst_regA_eff<28>/GROM )
  );
  X_BUF \DLX_IDinst_regA_eff<28>/XUSED  (
    .I(\DLX_IDinst_regA_eff<28>/FROM ),
    .O(\DLX_IDinst_regA_eff[28] )
  );
  X_BUF \DLX_IDinst_regA_eff<28>/YUSED  (
    .I(\DLX_IDinst_regA_eff<28>/GROM ),
    .O(CHOICE4255)
  );
  defparam \DLX_IDinst__n0114<29>20 .INIT = 16'hB080;
  X_LUT4 \DLX_IDinst__n0114<29>20  (
    .ADR0(DLX_MEMinst_RF_data_in[29]),
    .ADR1(DLX_IDinst__n0175),
    .ADR2(DLX_IDinst_N107837),
    .ADR3(DLX_IDinst__n0620[29]),
    .O(\CHOICE2401/FROM )
  );
  defparam \DLX_IDinst_Mmux_regA_eff_Result<29>1 .INIT = 16'hAAF0;
  X_LUT4 \DLX_IDinst_Mmux_regA_eff_Result<29>1  (
    .ADR0(DLX_MEMinst_RF_data_in[29]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst__n0620[29]),
    .ADR3(DLX_IDinst__n0175),
    .O(\CHOICE2401/GROM )
  );
  X_BUF \CHOICE2401/XUSED  (
    .I(\CHOICE2401/FROM ),
    .O(CHOICE2401)
  );
  X_BUF \CHOICE2401/YUSED  (
    .I(\CHOICE2401/GROM ),
    .O(\DLX_IDinst_regA_eff[29] )
  );
  defparam \DLX_EXinst__n0007<3>7 .INIT = 16'h0200;
  X_LUT4 \DLX_EXinst__n0007<3>7  (
    .ADR0(DLX_EXinst_N76463),
    .ADR1(\DLX_IDinst_Imm[3] ),
    .ADR2(\DLX_IDinst_Imm[2] ),
    .ADR3(\DLX_EXinst_Mshift__n0021_Sh[3] ),
    .O(\CHOICE5435/FROM )
  );
  defparam \DLX_EXinst__n0007<3>16 .INIT = 16'h5450;
  X_LUT4 \DLX_EXinst__n0007<3>16  (
    .ADR0(N146478),
    .ADR1(\DLX_EXinst_Mshift__n0022_Sh[51] ),
    .ADR2(CHOICE5435),
    .ADR3(DLX_EXinst_N76285),
    .O(\CHOICE5435/GROM )
  );
  X_BUF \CHOICE5435/XUSED  (
    .I(\CHOICE5435/FROM ),
    .O(CHOICE5435)
  );
  X_BUF \CHOICE5435/YUSED  (
    .I(\CHOICE5435/GROM ),
    .O(CHOICE5437)
  );
  defparam vga_top_vga1__n0011_SW1.INIT = 16'hFDDD;
  X_LUT4 vga_top_vga1__n0011_SW1 (
    .ADR0(vga_top_vga1_N112941),
    .ADR1(vga_top_vga1_vcounter[5]),
    .ADR2(vga_top_vga1_vcounter[2]),
    .ADR3(vga_top_vga1_vcounter[3]),
    .O(\N164108/FROM )
  );
  defparam vga_top_vga1__n0011_497.INIT = 16'hF3F7;
  X_LUT4 vga_top_vga1__n0011_497 (
    .ADR0(vga_top_vga1_vcounter[4]),
    .ADR1(vga_top_vga1_vcounter[9]),
    .ADR2(vga_top_vga1_helpme),
    .ADR3(N164108),
    .O(\N164108/GROM )
  );
  X_BUF \N164108/XUSED  (
    .I(\N164108/FROM ),
    .O(N164108)
  );
  X_BUF \N164108/YUSED  (
    .I(\N164108/GROM ),
    .O(vga_top_vga1__n0011)
  );
  defparam vga_top_vga1__n0012_SW0.INIT = 16'h33FF;
  X_LUT4 vga_top_vga1__n0012_SW0 (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_N112904),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_N112946),
    .O(\N127166/FROM )
  );
  defparam vga_top_vga1__n0012_498.INIT = 16'hF0F1;
  X_LUT4 vga_top_vga1__n0012_498 (
    .ADR0(vga_top_vga1_hcounter[5]),
    .ADR1(vga_top_vga1_hcounter[9]),
    .ADR2(reset_IBUF_1),
    .ADR3(N127166),
    .O(\N127166/GROM )
  );
  X_BUF \N127166/XUSED  (
    .I(\N127166/FROM ),
    .O(N127166)
  );
  X_BUF \N127166/YUSED  (
    .I(\N127166/GROM ),
    .O(vga_top_vga1__n0012)
  );
  defparam \DLX_EXinst_Mshift__n0024_Sh<30>1 .INIT = 16'h0B08;
  X_LUT4 \DLX_EXinst_Mshift__n0024_Sh<30>1  (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(DLX_IDinst_reg_out_B[0]),
    .ADR2(DLX_IDinst_reg_out_B[1]),
    .ADR3(DLX_IDinst_reg_out_A[30]),
    .O(\DLX_EXinst_Mshift__n0024_Sh<30>/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0024_Sh<58>1 .INIT = 16'h3202;
  X_LUT4 \DLX_EXinst_Mshift__n0024_Sh<58>1  (
    .ADR0(\DLX_EXinst_Mshift__n0019_Sh[26] ),
    .ADR1(DLX_IDinst_reg_out_B_3_1),
    .ADR2(DLX_IDinst_reg_out_B_2_1),
    .ADR3(\DLX_EXinst_Mshift__n0024_Sh[30] ),
    .O(\DLX_EXinst_Mshift__n0024_Sh<30>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0024_Sh<30>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0024_Sh<30>/FROM ),
    .O(\DLX_EXinst_Mshift__n0024_Sh[30] )
  );
  X_BUF \DLX_EXinst_Mshift__n0024_Sh<30>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0024_Sh<30>/GROM ),
    .O(\DLX_EXinst_Mshift__n0024_Sh[58] )
  );
  defparam \DLX_EXinst_Mshift__n0024_Sh<31>1 .INIT = 16'h0300;
  X_LUT4 \DLX_EXinst_Mshift__n0024_Sh<31>1  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(DLX_IDinst_reg_out_B[0]),
    .ADR3(DLX_IDinst_reg_out_A[31]),
    .O(\DLX_EXinst_Mshift__n0024_Sh<31>/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0024_Sh<59>1 .INIT = 16'h0E04;
  X_LUT4 \DLX_EXinst_Mshift__n0024_Sh<59>1  (
    .ADR0(DLX_IDinst_reg_out_B_2_1),
    .ADR1(\DLX_EXinst_Mshift__n0019_Sh[27] ),
    .ADR2(DLX_IDinst_reg_out_B_3_1),
    .ADR3(\DLX_EXinst_Mshift__n0024_Sh[31] ),
    .O(\DLX_EXinst_Mshift__n0024_Sh<31>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0024_Sh<31>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0024_Sh<31>/FROM ),
    .O(\DLX_EXinst_Mshift__n0024_Sh[31] )
  );
  X_BUF \DLX_EXinst_Mshift__n0024_Sh<31>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0024_Sh<31>/GROM ),
    .O(\DLX_EXinst_Mshift__n0024_Sh[59] )
  );
  defparam \DLX_EXinst_Mshift__n0024_Sh<51>1 .INIT = 16'hBB88;
  X_LUT4 \DLX_EXinst_Mshift__n0024_Sh<51>1  (
    .ADR0(DLX_EXinst_N73103),
    .ADR1(DLX_IDinst_reg_out_B_2_1),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N74976),
    .O(\DLX_EXinst_Mshift__n0024_Sh<51>/FROM )
  );
  defparam \DLX_EXinst__n0007<19>298_SW0 .INIT = 16'hFAAA;
  X_LUT4 \DLX_EXinst__n0007<19>298_SW0  (
    .ADR0(CHOICE5337),
    .ADR1(VCC),
    .ADR2(DLX_EXinst__n0081),
    .ADR3(\DLX_EXinst_Mshift__n0024_Sh[51] ),
    .O(\DLX_EXinst_Mshift__n0024_Sh<51>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0024_Sh<51>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0024_Sh<51>/FROM ),
    .O(\DLX_EXinst_Mshift__n0024_Sh[51] )
  );
  X_BUF \DLX_EXinst_Mshift__n0024_Sh<51>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0024_Sh<51>/GROM ),
    .O(N163696)
  );
  defparam vga_top_vga1__n0006_SW0.INIT = 16'hFFCF;
  X_LUT4 vga_top_vga1__n0006_SW0 (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_hcounter[3]),
    .ADR2(vga_top_vga1_N112936),
    .ADR3(vga_top_vga1_hcounter[0]),
    .O(\N132499/FROM )
  );
  defparam vga_top_vga1__n0006_499.INIT = 16'hCCEC;
  X_LUT4 vga_top_vga1__n0006_499 (
    .ADR0(vga_top_vga1_hcounter[9]),
    .ADR1(vga_top_vga1_helpme),
    .ADR2(vga_top_vga1_hcounter[8]),
    .ADR3(N132499),
    .O(\N132499/GROM )
  );
  X_BUF \N132499/XUSED  (
    .I(\N132499/FROM ),
    .O(N132499)
  );
  X_BUF \N132499/YUSED  (
    .I(\N132499/GROM ),
    .O(vga_top_vga1__n0006)
  );
  defparam DLX_IDinst_RegFile_26_15_500.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_26_15_500 (
    .I(DLX_IDinst_WB_data_eff[15]),
    .CE(DLX_IDinst__n0602),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_26_15)
  );
  defparam vga_top_vga1__n0007_SW0.INIT = 16'hDFFF;
  X_LUT4 vga_top_vga1__n0007_SW0 (
    .ADR0(vga_top_vga1_vcounter[1]),
    .ADR1(vga_top_vga1_vcounter[0]),
    .ADR2(vga_top_vga1_vcounter[3]),
    .ADR3(vga_top_vga1_vcounter[2]),
    .O(\N136799/FROM )
  );
  defparam vga_top_vga1__n0007_501.INIT = 16'hAAEA;
  X_LUT4 vga_top_vga1__n0007_501 (
    .ADR0(vga_top_vga1_helpme),
    .ADR1(vga_top_vga1_vcounter[9]),
    .ADR2(vga_top_vga1_N112910),
    .ADR3(N136799),
    .O(\N136799/GROM )
  );
  X_BUF \N136799/XUSED  (
    .I(\N136799/FROM ),
    .O(N136799)
  );
  X_BUF \N136799/YUSED  (
    .I(\N136799/GROM ),
    .O(vga_top_vga1__n0007)
  );
  defparam DLX_EXinst_Ker7551347.INIT = 16'h0200;
  X_LUT4 DLX_EXinst_Ker7551347 (
    .ADR0(DLX_EXinst_N76421),
    .ADR1(DLX_IDinst_reg_out_B_3_1),
    .ADR2(DLX_IDinst_reg_out_B_2_1),
    .ADR3(\DLX_EXinst_Mshift__n0024_Sh[29] ),
    .O(\CHOICE2040/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0024_Sh<57>1 .INIT = 16'h3120;
  X_LUT4 \DLX_EXinst_Mshift__n0024_Sh<57>1  (
    .ADR0(DLX_IDinst_reg_out_B_2_1),
    .ADR1(DLX_IDinst_reg_out_B_3_1),
    .ADR2(\DLX_EXinst_Mshift__n0024_Sh[29] ),
    .ADR3(\DLX_EXinst_Mshift__n0019_Sh[25] ),
    .O(\CHOICE2040/GROM )
  );
  X_BUF \CHOICE2040/XUSED  (
    .I(\CHOICE2040/FROM ),
    .O(CHOICE2040)
  );
  X_BUF \CHOICE2040/YUSED  (
    .I(\CHOICE2040/GROM ),
    .O(\DLX_EXinst_Mshift__n0024_Sh[57] )
  );
  defparam DLX_IDinst_RegFile_18_31_502.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_18_31_502 (
    .I(DLX_IDinst_WB_data_eff[31]),
    .CE(DLX_IDinst__n0586),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_18_31)
  );
  defparam \DLX_EXinst_Mshift__n0024_Sh<49>1 .INIT = 16'hFC0C;
  X_LUT4 \DLX_EXinst_Mshift__n0024_Sh<49>1  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N74726),
    .ADR2(DLX_IDinst_reg_out_B_2_1),
    .ADR3(DLX_EXinst_N73093),
    .O(\DLX_IDinst_RegFile_3_20/FROM )
  );
  defparam \DLX_EXinst__n0007<17>298_SW0 .INIT = 16'hFAF0;
  X_LUT4 \DLX_EXinst__n0007<17>298_SW0  (
    .ADR0(DLX_EXinst__n0081),
    .ADR1(VCC),
    .ADR2(CHOICE5416),
    .ADR3(\DLX_EXinst_Mshift__n0024_Sh[49] ),
    .O(\DLX_IDinst_RegFile_3_20/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_3_20/XUSED  (
    .I(\DLX_IDinst_RegFile_3_20/FROM ),
    .O(\DLX_EXinst_Mshift__n0024_Sh[49] )
  );
  X_BUF \DLX_IDinst_RegFile_3_20/YUSED  (
    .I(\DLX_IDinst_RegFile_3_20/GROM ),
    .O(N163598)
  );
  defparam DLX_EXinst_Ker74439.INIT = 16'hB8B8;
  X_LUT4 DLX_EXinst_Ker74439 (
    .ADR0(\DLX_EXinst_Mshift__n0019_Sh[22] ),
    .ADR1(DLX_IDinst_reg_out_B_3_1),
    .ADR2(N130569),
    .ADR3(VCC),
    .O(\DLX_EXinst_N74441/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0024_Sh<50>_SW0 .INIT = 16'hFA50;
  X_LUT4 \DLX_EXinst_Mshift__n0024_Sh<50>_SW0  (
    .ADR0(DLX_IDinst_reg_out_B_3_1),
    .ADR1(VCC),
    .ADR2(\DLX_EXinst_Mshift__n0019_Sh[22] ),
    .ADR3(\DLX_EXinst_Mshift__n0024_Sh[30] ),
    .O(\DLX_EXinst_N74441/GROM )
  );
  X_BUF \DLX_EXinst_N74441/XUSED  (
    .I(\DLX_EXinst_N74441/FROM ),
    .O(DLX_EXinst_N74441)
  );
  X_BUF \DLX_EXinst_N74441/YUSED  (
    .I(\DLX_EXinst_N74441/GROM ),
    .O(N131027)
  );
  defparam \mask<0>_SW1 .INIT = 16'h30FA;
  X_LUT4 \mask<0>_SW1  (
    .ADR0(DLX_EXinst_word),
    .ADR1(DLX_EXinst_ALU_result[1]),
    .ADR2(DLX_EXinst_byte),
    .ADR3(DLX_EXinst_ALU_result[0]),
    .O(\N164125/FROM )
  );
  defparam \mask<0> .INIT = 16'h0001;
  X_LUT4 \mask<0>  (
    .ADR0(DLX_EXinst_ALU_result[14]),
    .ADR1(DLX_EXinst_ALU_result[13]),
    .ADR2(DLX_EXinst_ALU_result[12]),
    .ADR3(N164125),
    .O(\N164125/GROM )
  );
  X_BUF \N164125/XUSED  (
    .I(\N164125/FROM ),
    .O(N164125)
  );
  X_BUF \N164125/YUSED  (
    .I(\N164125/GROM ),
    .O(mask_0_OBUF)
  );
  defparam DLX_EXinst_Ker74623_SW0.INIT = 16'h8800;
  X_LUT4 DLX_EXinst_Ker74623_SW0 (
    .ADR0(DLX_EXinst_N73267),
    .ADR1(DLX_IDinst_Imm_1_1),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N76412),
    .O(\DLX_IDinst_RegFile_18_1/FROM )
  );
  defparam DLX_EXinst_Ker74134_SW0.INIT = 16'h2200;
  X_LUT4 DLX_EXinst_Ker74134_SW0 (
    .ADR0(DLX_EXinst_N73267),
    .ADR1(DLX_IDinst_Imm_1_1),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N76412),
    .O(\DLX_IDinst_RegFile_18_1/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_18_1/XUSED  (
    .I(\DLX_IDinst_RegFile_18_1/FROM ),
    .O(N132037)
  );
  X_BUF \DLX_IDinst_RegFile_18_1/YUSED  (
    .I(\DLX_IDinst_RegFile_18_1/GROM ),
    .O(N131955)
  );
  defparam \mask<3>_SW1 .INIT = 16'hF8C8;
  X_LUT4 \mask<3>_SW1  (
    .ADR0(DLX_EXinst_ALU_result[1]),
    .ADR1(DLX_EXinst_byte),
    .ADR2(DLX_EXinst_ALU_result[0]),
    .ADR3(DLX_EXinst_word),
    .O(\N164115/FROM )
  );
  defparam \mask<3> .INIT = 16'h0001;
  X_LUT4 \mask<3>  (
    .ADR0(DLX_EXinst_ALU_result[13]),
    .ADR1(DLX_EXinst_ALU_result[12]),
    .ADR2(DLX_EXinst_ALU_result[14]),
    .ADR3(N164115),
    .O(\N164115/GROM )
  );
  X_BUF \N164115/XUSED  (
    .I(\N164115/FROM ),
    .O(N164115)
  );
  X_BUF \N164115/YUSED  (
    .I(\N164115/GROM ),
    .O(mask_3_OBUF)
  );
  defparam DLX_IDinst_Ker10739796.INIT = 16'h0001;
  X_LUT4 DLX_IDinst_Ker10739796 (
    .ADR0(DLX_IDinst_IR_opcode_field[0]),
    .ADR1(DLX_IDinst_IR_opcode_field[4]),
    .ADR2(DLX_IDinst_IR_opcode_field[1]),
    .ADR3(DLX_IDinst_IR_opcode_field[2]),
    .O(\DLX_IFinst_IR_previous<19>/FROM )
  );
  defparam DLX_EXinst__n0036_SW0.INIT = 16'hFEFE;
  X_LUT4 DLX_EXinst__n0036_SW0 (
    .ADR0(DLX_IDinst_IR_opcode_field[3]),
    .ADR1(DLX_IDinst_IR_opcode_field[2]),
    .ADR2(DLX_IDinst_IR_opcode_field[4]),
    .ADR3(VCC),
    .O(\DLX_IFinst_IR_previous<19>/GROM )
  );
  X_BUF \DLX_IFinst_IR_previous<19>/XUSED  (
    .I(\DLX_IFinst_IR_previous<19>/FROM ),
    .O(CHOICE1346)
  );
  X_BUF \DLX_IFinst_IR_previous<19>/YUSED  (
    .I(\DLX_IFinst_IR_previous<19>/GROM ),
    .O(N132091)
  );
  defparam DLX_IDinst_Ker1085361.INIT = 16'h2000;
  X_LUT4 DLX_IDinst_Ker1085361 (
    .ADR0(DLX_MEMinst_reg_dst_out[0]),
    .ADR1(DLX_MEMinst_reg_dst_out[4]),
    .ADR2(DLX_MEMinst_reg_dst_out[2]),
    .ADR3(DLX_MEMinst_reg_write_MEM),
    .O(\DLX_MEMinst_reg_write_MEM/FROM )
  );
  defparam DLX_IDinst__n05801.INIT = 16'hC000;
  X_LUT4 DLX_IDinst__n05801 (
    .ADR0(VCC),
    .ADR1(DLX_MEMinst_reg_dst_out[1]),
    .ADR2(DLX_MEMinst_reg_dst_out[3]),
    .ADR3(DLX_IDinst_N108538),
    .O(\DLX_MEMinst_reg_write_MEM/GROM )
  );
  X_BUF \DLX_MEMinst_reg_write_MEM/XUSED  (
    .I(\DLX_MEMinst_reg_write_MEM/FROM ),
    .O(DLX_IDinst_N108538)
  );
  X_BUF \DLX_MEMinst_reg_write_MEM/YUSED  (
    .I(\DLX_MEMinst_reg_write_MEM/GROM ),
    .O(DLX_IDinst__n0580)
  );
  defparam DLX_IDinst_RegFile_14_23_503.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_14_23_503 (
    .I(DLX_IDinst_WB_data_eff[23]),
    .CE(DLX_IDinst__n0578),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_14_23)
  );
  defparam DLX_EXinst__n0109_SW0.INIT = 16'h0404;
  X_LUT4 DLX_EXinst__n0109_SW0 (
    .ADR0(DLX_IDinst_IR_opcode_field[5]),
    .ADR1(DLX_IDinst_IR_opcode_field[3]),
    .ADR2(DLX_IDinst_IR_opcode_field[2]),
    .ADR3(VCC),
    .O(\DLX_IDinst_RegFile_14_23/FROM )
  );
  defparam DLX_EXinst__n0109_504.INIT = 16'h5540;
  X_LUT4 DLX_EXinst__n0109_504 (
    .ADR0(DLX_IDinst_IR_opcode_field[4]),
    .ADR1(DLX_IDinst_IR_opcode_field[5]),
    .ADR2(DLX_EXinst_N73345),
    .ADR3(N126741),
    .O(\DLX_IDinst_RegFile_14_23/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_14_23/XUSED  (
    .I(\DLX_IDinst_RegFile_14_23/FROM ),
    .O(N126741)
  );
  X_BUF \DLX_IDinst_RegFile_14_23/YUSED  (
    .I(\DLX_IDinst_RegFile_14_23/GROM ),
    .O(DLX_EXinst__n0109)
  );
  defparam \DLX_EXinst__n0007<31>293 .INIT = 16'h0D08;
  X_LUT4 \DLX_EXinst__n0007<31>293  (
    .ADR0(\DLX_IDinst_Imm[1] ),
    .ADR1(DLX_IDinst_reg_out_A[29]),
    .ADR2(\DLX_IDinst_Imm[0] ),
    .ADR3(DLX_IDinst_reg_out_A[31]),
    .O(\CHOICE5824/FROM )
  );
  defparam DLX_EXinst_Ker73285_SW0.INIT = 16'h8800;
  X_LUT4 DLX_EXinst_Ker73285_SW0 (
    .ADR0(DLX_EXinst_N76490),
    .ADR1(\DLX_IDinst_Imm[0] ),
    .ADR2(VCC),
    .ADR3(\DLX_IDinst_Imm[1] ),
    .O(\CHOICE5824/GROM )
  );
  X_BUF \CHOICE5824/XUSED  (
    .I(\CHOICE5824/FROM ),
    .O(CHOICE5824)
  );
  X_BUF \CHOICE5824/YUSED  (
    .I(\CHOICE5824/GROM ),
    .O(N132064)
  );
  defparam DLX_IDinst__n011750.INIT = 16'hFFF8;
  X_LUT4 DLX_IDinst__n011750 (
    .ADR0(DLX_IDinst_N108496),
    .ADR1(CHOICE3352),
    .ADR2(DLX_IDinst__n0453),
    .ADR3(CHOICE3359),
    .O(\DLX_IDinst_branch_sig/FROM )
  );
  defparam DLX_IDinst__n011761.INIT = 16'hFFFC;
  X_LUT4 DLX_IDinst__n011761 (
    .ADR0(VCC),
    .ADR1(CHOICE3348),
    .ADR2(DLX_IDinst_N108456),
    .ADR3(CHOICE3361),
    .O(\DLX_IDinst_branch_sig/GROM )
  );
  X_BUF \DLX_IDinst_branch_sig/XUSED  (
    .I(\DLX_IDinst_branch_sig/FROM ),
    .O(CHOICE3361)
  );
  X_BUF \DLX_IDinst_branch_sig/YUSED  (
    .I(\DLX_IDinst_branch_sig/GROM ),
    .O(N146990)
  );
  defparam DLX_IDinst__n013851_SW0.INIT = 16'h0245;
  X_LUT4 DLX_IDinst__n013851_SW0 (
    .ADR0(DLX_IDinst_IR_latched[27]),
    .ADR1(DLX_IDinst_IR_latched[28]),
    .ADR2(DLX_IDinst_IR_latched[26]),
    .ADR3(DLX_IDinst_IR_latched[30]),
    .O(\N163128/FROM )
  );
  defparam DLX_IDinst__n011814.INIT = 16'hF3FF;
  X_LUT4 DLX_IDinst__n011814 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_IR_latched[26]),
    .ADR2(DLX_IDinst_IR_latched[28]),
    .ADR3(DLX_IDinst_IR_latched[29]),
    .O(\N163128/GROM )
  );
  X_BUF \N163128/XUSED  (
    .I(\N163128/FROM ),
    .O(N163128)
  );
  X_BUF \N163128/YUSED  (
    .I(\N163128/GROM ),
    .O(CHOICE2301)
  );
  defparam DLX_IDinst__n011823.INIT = 16'hF0E0;
  X_LUT4 DLX_IDinst__n011823 (
    .ADR0(DLX_IDinst_IR_latched[30]),
    .ADR1(DLX_IDinst_IR_latched[31]),
    .ADR2(N164702),
    .ADR3(CHOICE2301),
    .O(\DLX_IDinst_Imm<31>/FROM )
  );
  defparam DLX_IDinst__n011832.INIT = 16'h0C00;
  X_LUT4 DLX_IDinst__n011832 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_jtarget[15]),
    .ADR2(DLX_IDinst_N108456),
    .ADR3(CHOICE2303),
    .O(\DLX_IDinst_Imm<31>/GROM )
  );
  X_BUF \DLX_IDinst_Imm<31>/XUSED  (
    .I(\DLX_IDinst_Imm<31>/FROM ),
    .O(CHOICE2303)
  );
  X_BUF \DLX_IDinst_Imm<31>/YUSED  (
    .I(\DLX_IDinst_Imm<31>/GROM ),
    .O(N140698)
  );
  defparam DLX_IDinst_Ker1084541.INIT = 16'hA000;
  X_LUT4 DLX_IDinst_Ker1084541 (
    .ADR0(DLX_IDinst_N108165),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_IR_latched[27]),
    .ADR3(DLX_IDinst_IR_latched[26]),
    .O(\DLX_IDinst_RegFile_10_6/FROM )
  );
  defparam DLX_IDinst__n011736.INIT = 16'h1400;
  X_LUT4 DLX_IDinst__n011736 (
    .ADR0(DLX_IDinst_IR_latched[26]),
    .ADR1(DLX_IDinst_IR_latched[30]),
    .ADR2(DLX_IDinst_IR_latched[27]),
    .ADR3(DLX_IDinst_N108165),
    .O(\DLX_IDinst_RegFile_10_6/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_10_6/XUSED  (
    .I(\DLX_IDinst_RegFile_10_6/FROM ),
    .O(DLX_IDinst_N108456)
  );
  X_BUF \DLX_IDinst_RegFile_10_6/YUSED  (
    .I(\DLX_IDinst_RegFile_10_6/GROM ),
    .O(CHOICE3359)
  );
  defparam DLX_IDinst__n015149_SW0.INIT = 16'hFFCF;
  X_LUT4 DLX_IDinst__n015149_SW0 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_IR_latched[27]),
    .ADR2(DLX_IDinst_N108496),
    .ADR3(DLX_IDinst_IR_latched[30]),
    .O(\N163842/FROM )
  );
  defparam DLX_IDinst__n015135.INIT = 16'h008C;
  X_LUT4 DLX_IDinst__n015135 (
    .ADR0(DLX_IDinst_N108496),
    .ADR1(DLX_IDinst_IR_latched[27]),
    .ADR2(DLX_IDinst_IR_latched[30]),
    .ADR3(DLX_IDinst_IR_latched[28]),
    .O(\N163842/GROM )
  );
  X_BUF \N163842/XUSED  (
    .I(\N163842/FROM ),
    .O(N163842)
  );
  X_BUF \N163842/YUSED  (
    .I(\N163842/GROM ),
    .O(CHOICE3328)
  );
  defparam DLX_IDinst__n015149.INIT = 16'h4400;
  X_LUT4 DLX_IDinst__n015149 (
    .ADR0(N163842),
    .ADR1(DLX_IDinst_IR_latched[28]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst__n0462),
    .O(\DLX_IDinst_RegFile_11_2/FROM )
  );
  defparam DLX_IDinst__n015169.INIT = 16'h0504;
  X_LUT4 DLX_IDinst__n015169 (
    .ADR0(DLX_IDinst_IR_latched[29]),
    .ADR1(CHOICE3328),
    .ADR2(DLX_IDinst_IR_latched[31]),
    .ADR3(CHOICE3335),
    .O(\DLX_IDinst_RegFile_11_2/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_11_2/XUSED  (
    .I(\DLX_IDinst_RegFile_11_2/FROM ),
    .O(CHOICE3335)
  );
  X_BUF \DLX_IDinst_RegFile_11_2/YUSED  (
    .I(\DLX_IDinst_RegFile_11_2/GROM ),
    .O(CHOICE3337)
  );
  defparam DLX_IDinst__n013725.INIT = 16'h330A;
  X_LUT4 DLX_IDinst__n013725 (
    .ADR0(DLX_IDinst__n0434),
    .ADR1(DLX_IDinst__n0433),
    .ADR2(DLX_IDinst__n0436),
    .ADR3(DLX_IDinst__n0167),
    .O(\CHOICE3508/FROM )
  );
  defparam DLX_IDinst__n013796_SW0.INIT = 16'hA2A0;
  X_LUT4 DLX_IDinst__n013796_SW0 (
    .ADR0(DLX_IDinst__n0629[1]),
    .ADR1(DLX_IDinst__n0166),
    .ADR2(CHOICE3515),
    .ADR3(CHOICE3508),
    .O(\CHOICE3508/GROM )
  );
  X_BUF \CHOICE3508/XUSED  (
    .I(\CHOICE3508/FROM ),
    .O(CHOICE3508)
  );
  X_BUF \CHOICE3508/YUSED  (
    .I(\CHOICE3508/GROM ),
    .O(N163554)
  );
  defparam DLX_IDinst__n013851.INIT = 16'h07F7;
  X_LUT4 DLX_IDinst__n013851 (
    .ADR0(DLX_IDinst_N108443),
    .ADR1(N163128),
    .ADR2(DLX_IDinst__n0437),
    .ADR3(DLX_IDinst__n0439),
    .O(\CHOICE3547/FROM )
  );
  defparam DLX_IDinst__n013899.INIT = 16'hA8A0;
  X_LUT4 DLX_IDinst__n013899 (
    .ADR0(CHOICE3552),
    .ADR1(DLX_IDinst_N108152),
    .ADR2(DLX_IDinst_N107405),
    .ADR3(CHOICE3547),
    .O(\CHOICE3547/GROM )
  );
  X_BUF \CHOICE3547/XUSED  (
    .I(\CHOICE3547/FROM ),
    .O(CHOICE3547)
  );
  X_BUF \CHOICE3547/YUSED  (
    .I(\CHOICE3547/GROM ),
    .O(CHOICE3553)
  );
  defparam DLX_IDinst_Ker107103_SW0.INIT = 16'h8000;
  X_LUT4 DLX_IDinst_Ker107103_SW0 (
    .ADR0(DLX_IDinst_N108244),
    .ADR1(DLX_IDinst_IR_latched[26]),
    .ADR2(DLX_IDinst_IR_latched[31]),
    .ADR3(DLX_IDinst_N108264),
    .O(\N164734/FROM )
  );
  defparam DLX_IDinst_Ker10735446_SW0.INIT = 16'hC004;
  X_LUT4 DLX_IDinst_Ker10735446_SW0 (
    .ADR0(DLX_IDinst__n0453),
    .ADR1(DLX_IDinst_N108264),
    .ADR2(DLX_IDinst_IR_latched[26]),
    .ADR3(DLX_IDinst_IR_latched[31]),
    .O(\N164734/GROM )
  );
  X_BUF \N164734/XUSED  (
    .I(\N164734/FROM ),
    .O(N164734)
  );
  X_BUF \N164734/YUSED  (
    .I(\N164734/GROM ),
    .O(N163836)
  );
  defparam DLX_EXinst_Ker74345_SW0.INIT = 16'h0800;
  X_LUT4 DLX_EXinst_Ker74345_SW0 (
    .ADR0(DLX_IDinst_Imm_1_1),
    .ADR1(DLX_EXinst_N73267),
    .ADR2(\DLX_IDinst_Imm[0] ),
    .ADR3(DLX_EXinst_N76412),
    .O(\N136586/FROM )
  );
  defparam DLX_EXinst_Ker74345.INIT = 16'hFF80;
  X_LUT4 DLX_EXinst_Ker74345 (
    .ADR0(DLX_EXinst_N75964),
    .ADR1(DLX_EXinst_N72710),
    .ADR2(DLX_EXinst_N76501),
    .ADR3(N136586),
    .O(\N136586/GROM )
  );
  X_BUF \N136586/XUSED  (
    .I(\N136586/FROM ),
    .O(N136586)
  );
  X_BUF \N136586/YUSED  (
    .I(\N136586/GROM ),
    .O(DLX_EXinst_N74347)
  );
  defparam DLX_IDinst__n013789.INIT = 16'h2202;
  X_LUT4 DLX_IDinst__n013789 (
    .ADR0(DLX_IDinst_N107572),
    .ADR1(DLX_IDinst__n0453),
    .ADR2(DLX_IDinst__n0100),
    .ADR3(DLX_IDinst__n0382),
    .O(\CHOICE3524/FROM )
  );
  defparam DLX_IDinst__n013796.INIT = 16'hF1F0;
  X_LUT4 DLX_IDinst__n013796 (
    .ADR0(DLX_IDinst__n0434),
    .ADR1(DLX_IDinst__n0167),
    .ADR2(N163554),
    .ADR3(CHOICE3524),
    .O(\CHOICE3524/GROM )
  );
  X_BUF \CHOICE3524/XUSED  (
    .I(\CHOICE3524/FROM ),
    .O(CHOICE3524)
  );
  X_BUF \CHOICE3524/YUSED  (
    .I(\CHOICE3524/GROM ),
    .O(CHOICE3526)
  );
  defparam \DLX_IDinst__n0145<0>15 .INIT = 16'h8A80;
  X_LUT4 \DLX_IDinst__n0145<0>15  (
    .ADR0(DLX_IDinst_N108238),
    .ADR1(N138903),
    .ADR2(DLX_IDinst__n0166),
    .ADR3(N137212),
    .O(\DLX_IDinst_RegFile_1_5/FROM )
  );
  defparam DLX_IDinst__n014952.INIT = 16'hF080;
  X_LUT4 DLX_IDinst__n014952 (
    .ADR0(DLX_IDinst_N108238),
    .ADR1(N138903),
    .ADR2(DLX_IDinst__n0166),
    .ADR3(N135079),
    .O(\DLX_IDinst_RegFile_1_5/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_1_5/XUSED  (
    .I(\DLX_IDinst_RegFile_1_5/FROM ),
    .O(CHOICE2911)
  );
  X_BUF \DLX_IDinst_RegFile_1_5/YUSED  (
    .I(\DLX_IDinst_RegFile_1_5/GROM ),
    .O(CHOICE3490)
  );
  defparam DLX_IDinst__n0164_505.INIT = 16'h0444;
  X_LUT4 DLX_IDinst__n0164_505 (
    .ADR0(DLX_IDinst_IR_latched[29]),
    .ADR1(DLX_IDinst_N108476),
    .ADR2(N127043),
    .ADR3(DLX_IDinst_IR_latched[27]),
    .O(\DLX_IDinst__n0164/FROM )
  );
  defparam DLX_IDinst__n013896.INIT = 16'h7777;
  X_LUT4 DLX_IDinst__n013896 (
    .ADR0(DLX_IDinst__n0427),
    .ADR1(DLX_IDinst_N108476),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IDinst__n0164/GROM )
  );
  X_BUF \DLX_IDinst__n0164/XUSED  (
    .I(\DLX_IDinst__n0164/FROM ),
    .O(DLX_IDinst__n0164)
  );
  X_BUF \DLX_IDinst__n0164/YUSED  (
    .I(\DLX_IDinst__n0164/GROM ),
    .O(CHOICE3552)
  );
  defparam DLX_IDinst__n04621.INIT = 16'h4800;
  X_LUT4 DLX_IDinst__n04621 (
    .ADR0(DLX_IDinst_zflag),
    .ADR1(DLX_IDinst_N108221),
    .ADR2(DLX_IDinst_IR_latched[26]),
    .ADR3(DLX_IDinst_N108443),
    .O(\DLX_IDinst_RegFile_22_11/FROM )
  );
  defparam DLX_IDinst_Ker10822663_SW0.INIT = 16'h0020;
  X_LUT4 DLX_IDinst_Ker10822663_SW0 (
    .ADR0(DLX_IDinst_N108443),
    .ADR1(DLX_IDinst_zflag),
    .ADR2(DLX_IDinst_N108221),
    .ADR3(DLX_IDinst_IR_latched[26]),
    .O(\DLX_IDinst_RegFile_22_11/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_22_11/XUSED  (
    .I(\DLX_IDinst_RegFile_22_11/FROM ),
    .O(DLX_IDinst__n0462)
  );
  X_BUF \DLX_IDinst_RegFile_22_11/YUSED  (
    .I(\DLX_IDinst_RegFile_22_11/GROM ),
    .O(N163831)
  );
  defparam DLX_IDinst__n014984.INIT = 16'h2220;
  X_LUT4 DLX_IDinst__n014984 (
    .ADR0(DLX_IDinst_N107033),
    .ADR1(DLX_IDinst__n0453),
    .ADR2(CHOICE3490),
    .ADR3(CHOICE3487),
    .O(\DLX_IDinst_stall/FROM )
  );
  defparam DLX_IDinst__n0149116.INIT = 16'hCDCC;
  X_LUT4 DLX_IDinst__n0149116 (
    .ADR0(DLX_IDinst__n0637),
    .ADR1(CHOICE3495),
    .ADR2(DLX_IDinst_Ker1084541_1),
    .ADR3(CHOICE3493),
    .O(\DLX_IDinst_stall/GROM )
  );
  X_BUF \DLX_IDinst_stall/XUSED  (
    .I(\DLX_IDinst_stall/FROM ),
    .O(CHOICE3493)
  );
  X_BUF \DLX_IDinst_stall/YUSED  (
    .I(\DLX_IDinst_stall/GROM ),
    .O(N147786)
  );
  defparam DLX_EXinst_Ker76181161_SW0.INIT = 16'hBFFF;
  X_LUT4 DLX_EXinst_Ker76181161_SW0 (
    .ADR0(DLX_IDinst_reg_out_B[30]),
    .ADR1(CHOICE3631),
    .ADR2(CHOICE3647),
    .ADR3(CHOICE3624),
    .O(\N163733/FROM )
  );
  defparam DLX_EXinst_Ker76181161.INIT = 16'h0020;
  X_LUT4 DLX_EXinst_Ker76181161 (
    .ADR0(CHOICE3616),
    .ADR1(DLX_IDinst_reg_out_B[31]),
    .ADR2(CHOICE3600),
    .ADR3(N163733),
    .O(\N163733/GROM )
  );
  X_BUF \N163733/XUSED  (
    .I(\N163733/FROM ),
    .O(N163733)
  );
  X_BUF \N163733/YUSED  (
    .I(\N163733/GROM ),
    .O(N148609)
  );
  defparam \DLX_IDinst__n0146<0>48_SW0 .INIT = 16'hEE44;
  X_LUT4 \DLX_IDinst__n0146<0>48_SW0  (
    .ADR0(DLX_IDinst__n0175),
    .ADR1(DLX_IDinst__n0620[0]),
    .ADR2(VCC),
    .ADR3(DLX_MEMinst_RF_data_in[0]),
    .O(\N163574/FROM )
  );
  defparam DLX_IDinst__n017716.INIT = 16'h0001;
  X_LUT4 DLX_IDinst__n017716 (
    .ADR0(DLX_IDinst__n0175),
    .ADR1(DLX_IDinst__n0620[0]),
    .ADR2(DLX_IDinst__n0620[31]),
    .ADR3(DLX_IDinst__n0620[6]),
    .O(\N163574/GROM )
  );
  X_BUF \N163574/XUSED  (
    .I(\N163574/FROM ),
    .O(N163574)
  );
  X_BUF \N163574/YUSED  (
    .I(\N163574/GROM ),
    .O(CHOICE4196)
  );
  defparam \DLX_IDinst__n0146<6>48_SW0 .INIT = 16'hFA0A;
  X_LUT4 \DLX_IDinst__n0146<6>48_SW0  (
    .ADR0(DLX_IDinst__n0620[6]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst__n0175),
    .ADR3(DLX_MEMinst_RF_data_in[6]),
    .O(\DLX_IFinst_IR_curr<28>/FROM )
  );
  defparam DLX_IDinst__n017728.INIT = 16'h0100;
  X_LUT4 DLX_IDinst__n017728 (
    .ADR0(DLX_MEMinst_RF_data_in[0]),
    .ADR1(DLX_MEMinst_RF_data_in[31]),
    .ADR2(DLX_MEMinst_RF_data_in[6]),
    .ADR3(DLX_IDinst__n0175),
    .O(\DLX_IFinst_IR_curr<28>/GROM )
  );
  X_BUF \DLX_IFinst_IR_curr<28>/XUSED  (
    .I(\DLX_IFinst_IR_curr<28>/FROM ),
    .O(N163724)
  );
  X_BUF \DLX_IFinst_IR_curr<28>/YUSED  (
    .I(\DLX_IFinst_IR_curr<28>/GROM ),
    .O(CHOICE4202)
  );
  defparam DLX_IDinst__n042812.INIT = 16'h3130;
  X_LUT4 DLX_IDinst__n042812 (
    .ADR0(DLX_IDinst_IR_latched[26]),
    .ADR1(DLX_IDinst_IR_latched[29]),
    .ADR2(DLX_IDinst_IR_latched[27]),
    .ADR3(DLX_IDinst_IR_latched[28]),
    .O(\CHOICE1971/FROM )
  );
  defparam DLX_IDinst__n042891.INIT = 16'h3222;
  X_LUT4 DLX_IDinst__n042891 (
    .ADR0(CHOICE1987),
    .ADR1(DLX_IDinst_IR_latched[31]),
    .ADR2(DLX_IDinst_IR_latched[30]),
    .ADR3(CHOICE1971),
    .O(\CHOICE1971/GROM )
  );
  X_BUF \CHOICE1971/XUSED  (
    .I(\CHOICE1971/FROM ),
    .O(CHOICE1971)
  );
  X_BUF \CHOICE1971/YUSED  (
    .I(\CHOICE1971/GROM ),
    .O(CHOICE1989)
  );
  defparam DLX_IDinst__n017757.INIT = 16'h0407;
  X_LUT4 DLX_IDinst__n017757 (
    .ADR0(DLX_MEMinst_RF_data_in[2]),
    .ADR1(DLX_IDinst__n0175),
    .ADR2(\DLX_IDinst_regA_eff[3] ),
    .ADR3(DLX_IDinst__n0620[2]),
    .O(\CHOICE4208/FROM )
  );
  defparam DLX_IDinst__n017761.INIT = 16'h5400;
  X_LUT4 DLX_IDinst__n017761 (
    .ADR0(\DLX_IDinst_regA_eff[1] ),
    .ADR1(CHOICE4202),
    .ADR2(CHOICE4196),
    .ADR3(CHOICE4208),
    .O(\CHOICE4208/GROM )
  );
  X_BUF \CHOICE4208/XUSED  (
    .I(\CHOICE4208/FROM ),
    .O(CHOICE4208)
  );
  X_BUF \CHOICE4208/YUSED  (
    .I(\CHOICE4208/GROM ),
    .O(CHOICE4209)
  );
  defparam DLX_EXinst__n0083_SW0.INIT = 16'hFCFF;
  X_LUT4 DLX_EXinst__n0083_SW0 (
    .ADR0(VCC),
    .ADR1(\DLX_IDinst_Imm[3] ),
    .ADR2(\DLX_IDinst_Imm[2] ),
    .ADR3(DLX_IDinst_IR_function_field[5]),
    .O(\N131907/FROM )
  );
  defparam DLX_EXinst__n0083_506.INIT = 16'h0200;
  X_LUT4 DLX_EXinst__n0083_506 (
    .ADR0(\DLX_IDinst_Imm[0] ),
    .ADR1(\DLX_IDinst_Imm[1] ),
    .ADR2(N131907),
    .ADR3(\DLX_IDinst_Imm[4] ),
    .O(\N131907/GROM )
  );
  X_BUF \N131907/XUSED  (
    .I(\N131907/FROM ),
    .O(N131907)
  );
  X_BUF \N131907/YUSED  (
    .I(\N131907/GROM ),
    .O(DLX_EXinst__n0083)
  );
  defparam DLX_IDinst_Ker10739777.INIT = 16'h57FF;
  X_LUT4 DLX_IDinst_Ker10739777 (
    .ADR0(DLX_IDinst_IR_opcode_field[2]),
    .ADR1(DLX_IDinst_IR_opcode_field[1]),
    .ADR2(DLX_IDinst_IR_opcode_field[0]),
    .ADR3(DLX_IDinst_IR_opcode_field[4]),
    .O(\CHOICE1338/FROM )
  );
  defparam DLX_EXinst_Ker72763_SW1.INIT = 16'hFEFF;
  X_LUT4 DLX_EXinst_Ker72763_SW1 (
    .ADR0(DLX_IDinst_IR_opcode_field[4]),
    .ADR1(DLX_IDinst_IR_opcode_field[2]),
    .ADR2(DLX_IDinst_reg_dst),
    .ADR3(DLX_IDinst_IR_opcode_field[5]),
    .O(\CHOICE1338/GROM )
  );
  X_BUF \CHOICE1338/XUSED  (
    .I(\CHOICE1338/FROM ),
    .O(CHOICE1338)
  );
  X_BUF \CHOICE1338/YUSED  (
    .I(\CHOICE1338/GROM ),
    .O(N164077)
  );
  defparam \DLX_IDinst__n0146<30>491 .INIT = 16'h0080;
  X_LUT4 \DLX_IDinst__n0146<30>491  (
    .ADR0(DLX_IDinst_Ker1084541_1),
    .ADR1(DLX_IDinst__n0116),
    .ADR2(DLX_IFinst_NPC[30]),
    .ADR3(DLX_IDinst__n0387),
    .O(N162964)
  );
  defparam DLX_IDinst_Ker107103.INIT = 16'hBF00;
  X_LUT4 DLX_IDinst_Ker107103 (
    .ADR0(DLX_IDinst__n0387),
    .ADR1(DLX_IDinst__n0116),
    .ADR2(DLX_IDinst_Ker1084541_1),
    .ADR3(N164734),
    .O(\DLX_IDinst_reg_out_A<30>/GROM )
  );
  X_BUF \DLX_IDinst_reg_out_A<30>/YUSED  (
    .I(\DLX_IDinst_reg_out_A<30>/GROM ),
    .O(DLX_IDinst_N107105)
  );
  defparam DLX_IDinst_RegFile_26_31_507.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_26_31_507 (
    .I(DLX_IDinst_WB_data_eff[31]),
    .CE(DLX_IDinst__n0602),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_26_31)
  );
  defparam \DLX_IDinst__n0114<1>20 .INIT = 16'hA0C0;
  X_LUT4 \DLX_IDinst__n0114<1>20  (
    .ADR0(DLX_MEMinst_RF_data_in[1]),
    .ADR1(DLX_IDinst__n0620[1]),
    .ADR2(DLX_IDinst_N107837),
    .ADR3(DLX_IDinst__n0175),
    .O(\CHOICE2148/FROM )
  );
  defparam \DLX_IDinst_Mmux_regA_eff_Result<1>1 .INIT = 16'hACAC;
  X_LUT4 \DLX_IDinst_Mmux_regA_eff_Result<1>1  (
    .ADR0(DLX_MEMinst_RF_data_in[1]),
    .ADR1(DLX_IDinst__n0620[1]),
    .ADR2(DLX_IDinst__n0175),
    .ADR3(VCC),
    .O(\CHOICE2148/GROM )
  );
  X_BUF \CHOICE2148/XUSED  (
    .I(\CHOICE2148/FROM ),
    .O(CHOICE2148)
  );
  X_BUF \CHOICE2148/YUSED  (
    .I(\CHOICE2148/GROM ),
    .O(\DLX_IDinst_regA_eff[1] )
  );
  defparam \DLX_IDinst__n0114<2>20 .INIT = 16'hC808;
  X_LUT4 \DLX_IDinst__n0114<2>20  (
    .ADR0(DLX_IDinst__n0620[2]),
    .ADR1(DLX_IDinst_N107837),
    .ADR2(DLX_IDinst__n0175),
    .ADR3(DLX_MEMinst_RF_data_in[2]),
    .O(\DLX_IFinst_IR_curr<29>/FROM )
  );
  defparam \DLX_IDinst_Mmux_regA_eff_Result<2>1 .INIT = 16'hFC0C;
  X_LUT4 \DLX_IDinst_Mmux_regA_eff_Result<2>1  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst__n0620[2]),
    .ADR2(DLX_IDinst__n0175),
    .ADR3(DLX_MEMinst_RF_data_in[2]),
    .O(\DLX_IFinst_IR_curr<29>/GROM )
  );
  X_BUF \DLX_IFinst_IR_curr<29>/XUSED  (
    .I(\DLX_IFinst_IR_curr<29>/FROM ),
    .O(CHOICE2159)
  );
  X_BUF \DLX_IFinst_IR_curr<29>/YUSED  (
    .I(\DLX_IFinst_IR_curr<29>/GROM ),
    .O(\DLX_IDinst_regA_eff[2] )
  );
  defparam \DLX_IDinst__n0114<3>20 .INIT = 16'hAC00;
  X_LUT4 \DLX_IDinst__n0114<3>20  (
    .ADR0(DLX_MEMinst_RF_data_in[3]),
    .ADR1(DLX_IDinst__n0620[3]),
    .ADR2(DLX_IDinst__n0175),
    .ADR3(DLX_IDinst_N107837),
    .O(\CHOICE2170/FROM )
  );
  defparam \DLX_IDinst_Mmux_regA_eff_Result<3>1 .INIT = 16'hCFC0;
  X_LUT4 \DLX_IDinst_Mmux_regA_eff_Result<3>1  (
    .ADR0(VCC),
    .ADR1(DLX_MEMinst_RF_data_in[3]),
    .ADR2(DLX_IDinst__n0175),
    .ADR3(DLX_IDinst__n0620[3]),
    .O(\CHOICE2170/GROM )
  );
  X_BUF \CHOICE2170/XUSED  (
    .I(\CHOICE2170/FROM ),
    .O(CHOICE2170)
  );
  X_BUF \CHOICE2170/YUSED  (
    .I(\CHOICE2170/GROM ),
    .O(\DLX_IDinst_regA_eff[3] )
  );
  defparam DLX_IDinst_Ker107171.INIT = 16'hBABB;
  X_LUT4 DLX_IDinst_Ker107171 (
    .ADR0(N127094),
    .ADR1(DLX_IDinst_Ker1084541_1),
    .ADR2(DLX_IDinst__n0453),
    .ADR3(DLX_IDinst__n0098),
    .O(\DLX_IDinst_reg_out_B<0>/FROM )
  );
  defparam \DLX_IDinst__n0147<0>1 .INIT = 16'hD800;
  X_LUT4 \DLX_IDinst__n0147<0>1  (
    .ADR0(DLX_IDinst__n0176),
    .ADR1(DLX_MEMinst_RF_data_in[0]),
    .ADR2(DLX_IDinst__n0623[0]),
    .ADR3(DLX_IDinst_N107173),
    .O(DLX_IDinst__n0147[0])
  );
  X_BUF \DLX_IDinst_reg_out_B<0>/XUSED  (
    .I(\DLX_IDinst_reg_out_B<0>/FROM ),
    .O(DLX_IDinst_N107173)
  );
  defparam \DLX_IDinst__n0114<4>20 .INIT = 16'hA808;
  X_LUT4 \DLX_IDinst__n0114<4>20  (
    .ADR0(DLX_IDinst_N107837),
    .ADR1(DLX_IDinst__n0620[4]),
    .ADR2(DLX_IDinst__n0175),
    .ADR3(DLX_MEMinst_RF_data_in[4]),
    .O(\CHOICE2181/FROM )
  );
  defparam \DLX_IDinst_Mmux_regA_eff_Result<4>1 .INIT = 16'hACAC;
  X_LUT4 \DLX_IDinst_Mmux_regA_eff_Result<4>1  (
    .ADR0(DLX_MEMinst_RF_data_in[4]),
    .ADR1(DLX_IDinst__n0620[4]),
    .ADR2(DLX_IDinst__n0175),
    .ADR3(VCC),
    .O(\CHOICE2181/GROM )
  );
  X_BUF \CHOICE2181/XUSED  (
    .I(\CHOICE2181/FROM ),
    .O(CHOICE2181)
  );
  X_BUF \CHOICE2181/YUSED  (
    .I(\CHOICE2181/GROM ),
    .O(\DLX_IDinst_regA_eff[4] )
  );
  defparam \DLX_IDinst_slot_num_FFd1-In1 .INIT = 16'h2000;
  X_LUT4 \DLX_IDinst_slot_num_FFd1-In1  (
    .ADR0(DLX_IDinst_delay_slot),
    .ADR1(DLX_IDinst_N108100),
    .ADR2(DLX_IDinst_slot_num_FFd2),
    .ADR3(N147200),
    .O(\DLX_IDinst_slot_num_FFd1-In )
  );
  defparam DLX_IDinst_Ker108231.INIT = 16'h0005;
  X_LUT4 DLX_IDinst_Ker108231 (
    .ADR0(DLX_IDinst__n0376),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_N108100),
    .ADR3(N132648),
    .O(\DLX_IDinst_slot_num_FFd1/GROM )
  );
  X_BUF \DLX_IDinst_slot_num_FFd1/YUSED  (
    .I(\DLX_IDinst_slot_num_FFd1/GROM ),
    .O(DLX_IDinst_N108233)
  );
  defparam \DLX_IDinst__n0114<5>20 .INIT = 16'hC808;
  X_LUT4 \DLX_IDinst__n0114<5>20  (
    .ADR0(DLX_IDinst__n0620[5]),
    .ADR1(DLX_IDinst_N107837),
    .ADR2(DLX_IDinst__n0175),
    .ADR3(DLX_MEMinst_RF_data_in[5]),
    .O(\CHOICE2192/FROM )
  );
  defparam \DLX_IDinst_Mmux_regA_eff_Result<5>1 .INIT = 16'hEE44;
  X_LUT4 \DLX_IDinst_Mmux_regA_eff_Result<5>1  (
    .ADR0(DLX_IDinst__n0175),
    .ADR1(DLX_IDinst__n0620[5]),
    .ADR2(VCC),
    .ADR3(DLX_MEMinst_RF_data_in[5]),
    .O(\CHOICE2192/GROM )
  );
  X_BUF \CHOICE2192/XUSED  (
    .I(\CHOICE2192/FROM ),
    .O(CHOICE2192)
  );
  X_BUF \CHOICE2192/YUSED  (
    .I(\CHOICE2192/GROM ),
    .O(\DLX_IDinst_regA_eff[5] )
  );
  defparam \DLX_IDinst__n0146<31>48_SW0 .INIT = 16'hB8B8;
  X_LUT4 \DLX_IDinst__n0146<31>48_SW0  (
    .ADR0(DLX_MEMinst_RF_data_in[31]),
    .ADR1(DLX_IDinst__n0175),
    .ADR2(DLX_IDinst__n0620[31]),
    .ADR3(VCC),
    .O(\N163652/FROM )
  );
  defparam \DLX_IDinst_Mmux_regA_eff_Result<7>1 .INIT = 16'hBB88;
  X_LUT4 \DLX_IDinst_Mmux_regA_eff_Result<7>1  (
    .ADR0(DLX_MEMinst_RF_data_in[7]),
    .ADR1(DLX_IDinst__n0175),
    .ADR2(VCC),
    .ADR3(DLX_IDinst__n0620[7]),
    .O(\N163652/GROM )
  );
  X_BUF \N163652/XUSED  (
    .I(\N163652/FROM ),
    .O(N163652)
  );
  X_BUF \N163652/YUSED  (
    .I(\N163652/GROM ),
    .O(\DLX_IDinst_regA_eff[7] )
  );
  defparam \DLX_IDinst_Mmux_regA_eff_Result<8>1 .INIT = 16'hCCAA;
  X_LUT4 \DLX_IDinst_Mmux_regA_eff_Result<8>1  (
    .ADR0(DLX_IDinst__n0620[8]),
    .ADR1(DLX_MEMinst_RF_data_in[8]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst__n0175),
    .O(\DLX_IDinst_RegFile_3_19/FROM )
  );
  defparam DLX_IDinst__n0177103.INIT = 16'h0001;
  X_LUT4 DLX_IDinst__n0177103 (
    .ADR0(\DLX_IDinst_regA_eff[5] ),
    .ADR1(\DLX_IDinst_regA_eff[4] ),
    .ADR2(\DLX_IDinst_regA_eff[7] ),
    .ADR3(\DLX_IDinst_regA_eff[8] ),
    .O(\DLX_IDinst_RegFile_3_19/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_3_19/XUSED  (
    .I(\DLX_IDinst_RegFile_3_19/FROM ),
    .O(\DLX_IDinst_regA_eff[8] )
  );
  X_BUF \DLX_IDinst_RegFile_3_19/YUSED  (
    .I(\DLX_IDinst_RegFile_3_19/GROM ),
    .O(CHOICE4217)
  );
  defparam \DLX_IDinst__n0114<9>20 .INIT = 16'h88A0;
  X_LUT4 \DLX_IDinst__n0114<9>20  (
    .ADR0(DLX_IDinst_N107837),
    .ADR1(DLX_MEMinst_RF_data_in[9]),
    .ADR2(DLX_IDinst__n0620[9]),
    .ADR3(DLX_IDinst__n0175),
    .O(\CHOICE2224/FROM )
  );
  defparam \DLX_IDinst_Mmux_regA_eff_Result<9>1 .INIT = 16'hF5A0;
  X_LUT4 \DLX_IDinst_Mmux_regA_eff_Result<9>1  (
    .ADR0(DLX_IDinst__n0175),
    .ADR1(VCC),
    .ADR2(DLX_MEMinst_RF_data_in[9]),
    .ADR3(DLX_IDinst__n0620[9]),
    .O(\CHOICE2224/GROM )
  );
  X_BUF \CHOICE2224/XUSED  (
    .I(\CHOICE2224/FROM ),
    .O(CHOICE2224)
  );
  X_BUF \CHOICE2224/YUSED  (
    .I(\CHOICE2224/GROM ),
    .O(\DLX_IDinst_regA_eff[9] )
  );
  defparam DLX_IDinst_Ker107835.INIT = 16'hACA0;
  X_LUT4 DLX_IDinst_Ker107835 (
    .ADR0(DLX_IDinst_IR_latched[30]),
    .ADR1(N137086),
    .ADR2(DLX_IDinst_Ker1084541_1),
    .ADR3(DLX_IDinst_N108496),
    .O(\DLX_IDinst_N107837/FROM )
  );
  defparam \DLX_IDinst__n0114<6>32 .INIT = 16'hCA00;
  X_LUT4 \DLX_IDinst__n0114<6>32  (
    .ADR0(DLX_IDinst__n0620[6]),
    .ADR1(DLX_MEMinst_RF_data_in[6]),
    .ADR2(DLX_IDinst__n0175),
    .ADR3(DLX_IDinst_N107837),
    .O(\DLX_IDinst_N107837/GROM )
  );
  X_BUF \DLX_IDinst_N107837/XUSED  (
    .I(\DLX_IDinst_N107837/FROM ),
    .O(DLX_IDinst_N107837)
  );
  X_BUF \DLX_IDinst_N107837/YUSED  (
    .I(\DLX_IDinst_N107837/GROM ),
    .O(CHOICE3193)
  );
  defparam \DLX_EXinst__n0007<25>9 .INIT = 16'hCE00;
  X_LUT4 \DLX_EXinst__n0007<25>9  (
    .ADR0(DLX_EXinst__n0054),
    .ADR1(DLX_EXinst__n0053),
    .ADR2(\DLX_IDinst_Imm[31] ),
    .ADR3(DLX_IDinst_reg_out_A[25]),
    .O(\CHOICE5058/FROM )
  );
  defparam \DLX_EXinst__n0007<10>141 .INIT = 16'hC0E0;
  X_LUT4 \DLX_EXinst__n0007<10>141  (
    .ADR0(DLX_EXinst__n0054),
    .ADR1(DLX_EXinst__n0053),
    .ADR2(DLX_IDinst_reg_out_A[10]),
    .ADR3(\DLX_IDinst_Imm[10] ),
    .O(\CHOICE5058/GROM )
  );
  X_BUF \CHOICE5058/XUSED  (
    .I(\CHOICE5058/FROM ),
    .O(CHOICE5058)
  );
  X_BUF \CHOICE5058/YUSED  (
    .I(\CHOICE5058/GROM ),
    .O(CHOICE4479)
  );
  defparam \DLX_EXinst__n0007<9>126 .INIT = 16'hEAC0;
  X_LUT4 \DLX_EXinst__n0007<9>126  (
    .ADR0(\DLX_EXinst_Mshift__n0021_Sh[41] ),
    .ADR1(\DLX_EXinst_Mshift__n0022_Sh[57] ),
    .ADR2(DLX_EXinst_N76285),
    .ADR3(DLX_EXinst_N76463),
    .O(\DLX_IDinst_RegFile_2_5/FROM )
  );
  defparam \DLX_EXinst__n0007<10>126 .INIT = 16'hF888;
  X_LUT4 \DLX_EXinst__n0007<10>126  (
    .ADR0(\DLX_EXinst_Mshift__n0021_Sh[42] ),
    .ADR1(DLX_EXinst_N76463),
    .ADR2(DLX_EXinst_N76285),
    .ADR3(\DLX_EXinst_Mshift__n0022_Sh[58] ),
    .O(\DLX_IDinst_RegFile_2_5/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_2_5/XUSED  (
    .I(\DLX_IDinst_RegFile_2_5/FROM ),
    .O(CHOICE4534)
  );
  X_BUF \DLX_IDinst_RegFile_2_5/YUSED  (
    .I(\DLX_IDinst_RegFile_2_5/GROM ),
    .O(CHOICE4474)
  );
  defparam DLX_EXinst__n00541.INIT = 16'h0A00;
  X_LUT4 DLX_EXinst__n00541 (
    .ADR0(DLX_EXinst_N76011),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_IR_opcode_field[0]),
    .ADR3(DLX_IDinst_IR_opcode_field[1]),
    .O(\DLX_EXinst__n0054/FROM )
  );
  defparam \DLX_EXinst__n0007<10>175 .INIT = 16'h02A8;
  X_LUT4 \DLX_EXinst__n0007<10>175  (
    .ADR0(DLX_EXinst_N76011),
    .ADR1(DLX_IDinst_reg_out_A[10]),
    .ADR2(DLX_IDinst_IR_opcode_field[0]),
    .ADR3(DLX_IDinst_IR_opcode_field[1]),
    .O(\DLX_EXinst__n0054/GROM )
  );
  X_BUF \DLX_EXinst__n0054/XUSED  (
    .I(\DLX_EXinst__n0054/FROM ),
    .O(DLX_EXinst__n0054)
  );
  X_BUF \DLX_EXinst__n0054/YUSED  (
    .I(\DLX_EXinst__n0054/GROM ),
    .O(CHOICE4490)
  );
  defparam \DLX_EXinst__n0007<1>88 .INIT = 16'h8080;
  X_LUT4 \DLX_EXinst__n0007<1>88  (
    .ADR0(\DLX_IDinst_Imm[4] ),
    .ADR1(N138037),
    .ADR2(N147520),
    .ADR3(VCC),
    .O(\CHOICE5713/FROM )
  );
  defparam \DLX_EXinst__n0007<10>184 .INIT = 16'h8080;
  X_LUT4 \DLX_EXinst__n0007<10>184  (
    .ADR0(N138143),
    .ADR1(\DLX_IDinst_Imm[4] ),
    .ADR2(N147520),
    .ADR3(VCC),
    .O(\CHOICE5713/GROM )
  );
  X_BUF \CHOICE5713/XUSED  (
    .I(\CHOICE5713/FROM ),
    .O(CHOICE5713)
  );
  X_BUF \CHOICE5713/YUSED  (
    .I(\CHOICE5713/GROM ),
    .O(CHOICE4493)
  );
  defparam \DLX_EXinst__n0007<27>9 .INIT = 16'hAE00;
  X_LUT4 \DLX_EXinst__n0007<27>9  (
    .ADR0(DLX_EXinst__n0053),
    .ADR1(DLX_EXinst__n0054),
    .ADR2(\DLX_IDinst_Imm[31] ),
    .ADR3(DLX_IDinst_reg_out_A[27]),
    .O(\CHOICE4924/FROM )
  );
  defparam \DLX_EXinst__n0007<11>141 .INIT = 16'hA0E0;
  X_LUT4 \DLX_EXinst__n0007<11>141  (
    .ADR0(DLX_EXinst__n0053),
    .ADR1(DLX_EXinst__n0054),
    .ADR2(DLX_IDinst_reg_out_A[11]),
    .ADR3(\DLX_IDinst_Imm[11] ),
    .O(\CHOICE4924/GROM )
  );
  X_BUF \CHOICE4924/XUSED  (
    .I(\CHOICE4924/FROM ),
    .O(CHOICE4924)
  );
  X_BUF \CHOICE4924/YUSED  (
    .I(\CHOICE4924/GROM ),
    .O(CHOICE4419)
  );
  defparam DLX_EXinst__n00511.INIT = 16'h8080;
  X_LUT4 DLX_EXinst__n00511 (
    .ADR0(DLX_IDinst_IR_opcode_field[1]),
    .ADR1(DLX_EXinst_N76011),
    .ADR2(DLX_IDinst_IR_opcode_field[0]),
    .ADR3(VCC),
    .O(\DLX_IDinst_RegFile_27_25/FROM )
  );
  defparam \DLX_EXinst__n0007<11>175 .INIT = 16'h10E0;
  X_LUT4 \DLX_EXinst__n0007<11>175  (
    .ADR0(DLX_IDinst_IR_opcode_field[0]),
    .ADR1(DLX_IDinst_reg_out_A[11]),
    .ADR2(DLX_EXinst_N76011),
    .ADR3(DLX_IDinst_IR_opcode_field[1]),
    .O(\DLX_IDinst_RegFile_27_25/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_27_25/XUSED  (
    .I(\DLX_IDinst_RegFile_27_25/FROM ),
    .O(DLX_EXinst__n0051)
  );
  X_BUF \DLX_IDinst_RegFile_27_25/YUSED  (
    .I(\DLX_IDinst_RegFile_27_25/GROM ),
    .O(CHOICE4430)
  );
  defparam \DLX_EXinst__n0007<3>88 .INIT = 16'h8800;
  X_LUT4 \DLX_EXinst__n0007<3>88  (
    .ADR0(N138713),
    .ADR1(\DLX_IDinst_Imm[4] ),
    .ADR2(VCC),
    .ADR3(N147520),
    .O(\CHOICE5458/FROM )
  );
  defparam \DLX_EXinst__n0007<11>184 .INIT = 16'h8080;
  X_LUT4 \DLX_EXinst__n0007<11>184  (
    .ADR0(N137774),
    .ADR1(\DLX_IDinst_Imm[4] ),
    .ADR2(N147520),
    .ADR3(VCC),
    .O(\CHOICE5458/GROM )
  );
  X_BUF \CHOICE5458/XUSED  (
    .I(\CHOICE5458/FROM ),
    .O(CHOICE5458)
  );
  X_BUF \CHOICE5458/YUSED  (
    .I(\CHOICE5458/GROM ),
    .O(CHOICE4433)
  );
  defparam DLX_EXinst__n00521.INIT = 16'h000C;
  X_LUT4 DLX_EXinst__n00521 (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N76011),
    .ADR2(DLX_IDinst_IR_opcode_field[0]),
    .ADR3(DLX_IDinst_IR_opcode_field[1]),
    .O(\DLX_EXinst__n0052/FROM )
  );
  defparam \DLX_EXinst__n0007<20>107 .INIT = 16'h2228;
  X_LUT4 \DLX_EXinst__n0007<20>107  (
    .ADR0(DLX_EXinst_N76011),
    .ADR1(DLX_IDinst_IR_opcode_field[1]),
    .ADR2(DLX_IDinst_reg_out_A[20]),
    .ADR3(DLX_IDinst_IR_opcode_field[0]),
    .O(\DLX_EXinst__n0052/GROM )
  );
  X_BUF \DLX_EXinst__n0052/XUSED  (
    .I(\DLX_EXinst__n0052/FROM ),
    .O(DLX_EXinst__n0052)
  );
  X_BUF \DLX_EXinst__n0052/YUSED  (
    .I(\DLX_EXinst__n0052/GROM ),
    .O(CHOICE4659)
  );
  defparam \DLX_EXinst__n0007<20>116 .INIT = 16'hECA0;
  X_LUT4 \DLX_EXinst__n0007<20>116  (
    .ADR0(DLX_EXinst__n0109),
    .ADR1(CHOICE4659),
    .ADR2(DLX_EXinst__n0012[20]),
    .ADR3(\DLX_IDinst_Imm[31] ),
    .O(\CHOICE4661/FROM )
  );
  defparam \DLX_EXinst__n0007<20>137_SW0 .INIT = 16'hFFF0;
  X_LUT4 \DLX_EXinst__n0007<20>137_SW0  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(CHOICE4653),
    .ADR3(CHOICE4661),
    .O(\CHOICE4661/GROM )
  );
  X_BUF \CHOICE4661/XUSED  (
    .I(\CHOICE4661/FROM ),
    .O(CHOICE4661)
  );
  X_BUF \CHOICE4661/YUSED  (
    .I(\CHOICE4661/GROM ),
    .O(N163174)
  );
  defparam \DLX_EXinst__n0007<20>310 .INIT = 16'hF0E0;
  X_LUT4 \DLX_EXinst__n0007<20>310  (
    .ADR0(N163473),
    .ADR1(CHOICE4676),
    .ADR2(DLX_EXinst__n0036),
    .ADR3(CHOICE4669),
    .O(\DLX_IDinst_RegFile_3_1/FROM )
  );
  defparam \DLX_EXinst__n0007<20>321 .INIT = 16'hFFC0;
  X_LUT4 \DLX_EXinst__n0007<20>321  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[31]),
    .ADR2(CHOICE929),
    .ADR3(CHOICE4699),
    .O(\DLX_IDinst_RegFile_3_1/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_3_1/XUSED  (
    .I(\DLX_IDinst_RegFile_3_1/FROM ),
    .O(CHOICE4699)
  );
  X_BUF \DLX_IDinst_RegFile_3_1/YUSED  (
    .I(\DLX_IDinst_RegFile_3_1/GROM ),
    .O(CHOICE4700)
  );
  defparam DLX_IDinst_RegFile_18_16_508.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_18_16_508 (
    .I(DLX_IDinst_WB_data_eff[16]),
    .CE(DLX_IDinst__n0586),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_18_16)
  );
  defparam \DLX_EXinst__n0007<25>97_SW0 .INIT = 16'h5060;
  X_LUT4 \DLX_EXinst__n0007<25>97_SW0  (
    .ADR0(DLX_IDinst_IR_opcode_field[1]),
    .ADR1(DLX_IDinst_reg_out_A[25]),
    .ADR2(DLX_EXinst_N76011),
    .ADR3(DLX_IDinst_IR_opcode_field[0]),
    .O(\N163606/FROM )
  );
  defparam \DLX_EXinst__n0007<12>127 .INIT = 16'h10E0;
  X_LUT4 \DLX_EXinst__n0007<12>127  (
    .ADR0(DLX_IDinst_IR_opcode_field[0]),
    .ADR1(DLX_IDinst_reg_out_A[12]),
    .ADR2(DLX_EXinst_N76011),
    .ADR3(DLX_IDinst_IR_opcode_field[1]),
    .O(\N163606/GROM )
  );
  X_BUF \N163606/XUSED  (
    .I(\N163606/FROM ),
    .O(N163606)
  );
  X_BUF \N163606/YUSED  (
    .I(\N163606/GROM ),
    .O(CHOICE3793)
  );
  defparam \DLX_EXinst__n0007<20>224 .INIT = 16'hA820;
  X_LUT4 \DLX_EXinst__n0007<20>224  (
    .ADR0(DLX_EXinst__n0080),
    .ADR1(DLX_IDinst_reg_out_B[3]),
    .ADR2(DLX_EXinst_N75006),
    .ADR3(DLX_EXinst_N74051),
    .O(\CHOICE4688/FROM )
  );
  defparam \DLX_EXinst__n0007<20>246_SW0 .INIT = 16'hFFC0;
  X_LUT4 \DLX_EXinst__n0007<20>246_SW0  (
    .ADR0(VCC),
    .ADR1(\DLX_EXinst_Mshift__n0024_Sh[52] ),
    .ADR2(DLX_EXinst__n0081),
    .ADR3(CHOICE4688),
    .O(\CHOICE4688/GROM )
  );
  X_BUF \CHOICE4688/XUSED  (
    .I(\CHOICE4688/FROM ),
    .O(CHOICE4688)
  );
  X_BUF \CHOICE4688/YUSED  (
    .I(\CHOICE4688/GROM ),
    .O(N163485)
  );
  defparam \DLX_EXinst__n0007<20>137 .INIT = 16'hFFD8;
  X_LUT4 \DLX_EXinst__n0007<20>137  (
    .ADR0(\DLX_IDinst_Imm[4] ),
    .ADR1(CHOICE4634),
    .ADR2(CHOICE4647),
    .ADR3(N163174),
    .O(\DLX_EXinst_ALU_result<20>/FROM )
  );
  defparam \DLX_EXinst__n0007<20>3361 .INIT = 16'h0F00;
  X_LUT4 \DLX_EXinst__n0007<20>3361  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_EXinst__n0036),
    .ADR3(CHOICE4663),
    .O(N162820)
  );
  X_BUF \DLX_EXinst_ALU_result<20>/XUSED  (
    .I(\DLX_EXinst_ALU_result<20>/FROM ),
    .O(CHOICE4663)
  );
  defparam DLX_IDinst_RegFile_18_24_509.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_18_24_509 (
    .I(DLX_IDinst_WB_data_eff[24]),
    .CE(DLX_IDinst__n0586),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_18_24)
  );
  defparam \DLX_EXinst__n0007<14>156 .INIT = 16'hE400;
  X_LUT4 \DLX_EXinst__n0007<14>156  (
    .ADR0(\DLX_IDinst_Imm[2] ),
    .ADR1(DLX_EXinst_N74701),
    .ADR2(DLX_EXinst_N74986),
    .ADR3(DLX_EXinst_N73267),
    .O(\DLX_IDinst_RegFile_3_27/FROM )
  );
  defparam \DLX_EXinst__n0007<12>156 .INIT = 16'hC0A0;
  X_LUT4 \DLX_EXinst__n0007<12>156  (
    .ADR0(DLX_EXinst_N74706),
    .ADR1(DLX_EXinst_N74971),
    .ADR2(DLX_EXinst_N73267),
    .ADR3(\DLX_IDinst_Imm[2] ),
    .O(\DLX_IDinst_RegFile_3_27/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_3_27/XUSED  (
    .I(\DLX_IDinst_RegFile_3_27/FROM ),
    .O(CHOICE3692)
  );
  X_BUF \DLX_IDinst_RegFile_3_27/YUSED  (
    .I(\DLX_IDinst_RegFile_3_27/GROM ),
    .O(CHOICE3802)
  );
  defparam \DLX_EXinst__n0007<20>9 .INIT = 16'hCCEC;
  X_LUT4 \DLX_EXinst__n0007<20>9  (
    .ADR0(DLX_EXinst_N76318),
    .ADR1(DLX_EXinst__n0051),
    .ADR2(DLX_EXinst_N72983),
    .ADR3(\DLX_IDinst_Imm[3] ),
    .O(\CHOICE4634/FROM )
  );
  defparam \DLX_EXinst__n0007<12>157 .INIT = 16'hC808;
  X_LUT4 \DLX_EXinst__n0007<12>157  (
    .ADR0(DLX_EXinst_N74223),
    .ADR1(DLX_EXinst_N76318),
    .ADR2(\DLX_IDinst_Imm[3] ),
    .ADR3(DLX_EXinst_N72983),
    .O(\CHOICE4634/GROM )
  );
  X_BUF \CHOICE4634/XUSED  (
    .I(\CHOICE4634/FROM ),
    .O(CHOICE4634)
  );
  X_BUF \CHOICE4634/YUSED  (
    .I(\CHOICE4634/GROM ),
    .O(CHOICE3803)
  );
  defparam \DLX_EXinst__n0007<20>269_SW0 .INIT = 16'hFFE2;
  X_LUT4 \DLX_EXinst__n0007<20>269_SW0  (
    .ADR0(DLX_EXinst__n0079),
    .ADR1(DLX_IDinst_reg_out_B[20]),
    .ADR2(DLX_EXinst__n0077),
    .ADR3(DLX_EXinst_N74245),
    .O(\N163481/FROM )
  );
  defparam \DLX_EXinst__n0007<20>174 .INIT = 16'h8C88;
  X_LUT4 \DLX_EXinst__n0007<20>174  (
    .ADR0(DLX_EXinst__n0078),
    .ADR1(DLX_IDinst_reg_out_B[20]),
    .ADR2(DLX_IDinst_reg_out_A[20]),
    .ADR3(DLX_EXinst__n0079),
    .O(\N163481/GROM )
  );
  X_BUF \N163481/XUSED  (
    .I(\N163481/FROM ),
    .O(N163481)
  );
  X_BUF \N163481/YUSED  (
    .I(\N163481/GROM ),
    .O(CHOICE4669)
  );
  defparam \DLX_EXinst__n0007<31>464 .INIT = 16'h2000;
  X_LUT4 \DLX_EXinst__n0007<31>464  (
    .ADR0(N147520),
    .ADR1(\DLX_IDinst_Imm[4] ),
    .ADR2(\DLX_EXinst_Mshift__n0020_Sh[127] ),
    .ADR3(\DLX_IDinst_Imm[5] ),
    .O(\DLX_IDinst_RegFile_23_8/FROM )
  );
  defparam \DLX_EXinst__n0007<31>429 .INIT = 16'h00C0;
  X_LUT4 \DLX_EXinst__n0007<31>429  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst__n0056),
    .ADR2(\DLX_EXinst_Mshift__n0020_Sh[127] ),
    .ADR3(\DLX_IDinst_Imm[4] ),
    .O(\DLX_IDinst_RegFile_23_8/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_23_8/XUSED  (
    .I(\DLX_IDinst_RegFile_23_8/FROM ),
    .O(CHOICE5846)
  );
  X_BUF \DLX_IDinst_RegFile_23_8/YUSED  (
    .I(\DLX_IDinst_RegFile_23_8/GROM ),
    .O(CHOICE5841)
  );
  defparam \DLX_EXinst_Mshift__n0021_Sh<40>_SW0 .INIT = 16'h4747;
  X_LUT4 \DLX_EXinst_Mshift__n0021_Sh<40>_SW0  (
    .ADR0(\DLX_EXinst_Mshift__n0021_Sh[0] ),
    .ADR1(DLX_IDinst_Imm_3_1),
    .ADR2(\DLX_EXinst_Mshift__n0021_Sh[8] ),
    .ADR3(VCC),
    .O(\N131375/FROM )
  );
  defparam \DLX_EXinst__n0007<16>223 .INIT = 16'hFF08;
  X_LUT4 \DLX_EXinst__n0007<16>223  (
    .ADR0(\DLX_EXinst_Mshift__n0021_Sh[0] ),
    .ADR1(\DLX_IDinst_Imm[4] ),
    .ADR2(DLX_EXinst_N72815),
    .ADR3(CHOICE4608),
    .O(\N131375/GROM )
  );
  X_BUF \N131375/XUSED  (
    .I(\N131375/FROM ),
    .O(N131375)
  );
  X_BUF \N131375/YUSED  (
    .I(\N131375/GROM ),
    .O(CHOICE4609)
  );
  defparam \DLX_EXinst__n0007<16>312 .INIT = 16'hFEFA;
  X_LUT4 \DLX_EXinst__n0007<16>312  (
    .ADR0(CHOICE4614),
    .ADR1(CHOICE4609),
    .ADR2(CHOICE4625),
    .ADR3(DLX_EXinst_N76318),
    .O(\DLX_EXinst_ALU_result<16>/FROM )
  );
  defparam \DLX_EXinst__n0007<16>342 .INIT = 16'hDDCC;
  X_LUT4 \DLX_EXinst__n0007<16>342  (
    .ADR0(DLX_EXinst__n0036),
    .ADR1(CHOICE4316),
    .ADR2(VCC),
    .ADR3(CHOICE4626),
    .O(CHOICE4629)
  );
  X_BUF \DLX_EXinst_ALU_result<16>/XUSED  (
    .I(\DLX_EXinst_ALU_result<16>/FROM ),
    .O(CHOICE4626)
  );
  defparam \DLX_EXinst__n0007<24>144 .INIT = 16'hF5E4;
  X_LUT4 \DLX_EXinst__n0007<24>144  (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(CHOICE5617),
    .ADR2(\DLX_EXinst_Mshift__n0023_Sh[40] ),
    .ADR3(CHOICE5618),
    .O(\CHOICE5622/FROM )
  );
  defparam \DLX_EXinst__n0007<24>193 .INIT = 16'h3222;
  X_LUT4 \DLX_EXinst__n0007<24>193  (
    .ADR0(CHOICE5628),
    .ADR1(N148323),
    .ADR2(DLX_EXinst__n0080),
    .ADR3(CHOICE5622),
    .O(\CHOICE5622/GROM )
  );
  X_BUF \CHOICE5622/XUSED  (
    .I(\CHOICE5622/FROM ),
    .O(CHOICE5622)
  );
  X_BUF \CHOICE5622/YUSED  (
    .I(\CHOICE5622/GROM ),
    .O(CHOICE5630)
  );
  defparam \DLX_EXinst__n0007<21>70 .INIT = 16'hF888;
  X_LUT4 \DLX_EXinst__n0007<21>70  (
    .ADR0(DLX_EXinst__n0109),
    .ADR1(DLX_EXinst__n0012[21]),
    .ADR2(DLX_EXinst__n0051),
    .ADR3(\DLX_IDinst_Imm[5] ),
    .O(\DLX_IDinst_RegFile_7_3/FROM )
  );
  defparam \DLX_EXinst__n0007<31>483 .INIT = 16'hEAC0;
  X_LUT4 \DLX_EXinst__n0007<31>483  (
    .ADR0(DLX_EXinst__n0109),
    .ADR1(\DLX_IDinst_Imm[15] ),
    .ADR2(DLX_EXinst__n0051),
    .ADR3(DLX_EXinst__n0012[31]),
    .O(\DLX_IDinst_RegFile_7_3/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_7_3/XUSED  (
    .I(\DLX_IDinst_RegFile_7_3/FROM ),
    .O(CHOICE4140)
  );
  X_BUF \DLX_IDinst_RegFile_7_3/YUSED  (
    .I(\DLX_IDinst_RegFile_7_3/GROM ),
    .O(CHOICE5850)
  );
  defparam \DLX_EXinst__n0007<24>411 .INIT = 16'h0400;
  X_LUT4 \DLX_EXinst__n0007<24>411  (
    .ADR0(\DLX_IDinst_Imm[3] ),
    .ADR1(DLX_EXinst_N73379),
    .ADR2(\DLX_IDinst_Imm[4] ),
    .ADR3(DLX_EXinst__n0056),
    .O(\CHOICE5677/FROM )
  );
  defparam \DLX_EXinst__n0007<24>429 .INIT = 16'h3320;
  X_LUT4 \DLX_EXinst__n0007<24>429  (
    .ADR0(CHOICE5671),
    .ADR1(N146478),
    .ADR2(DLX_EXinst__n0055),
    .ADR3(CHOICE5677),
    .O(\CHOICE5677/GROM )
  );
  X_BUF \CHOICE5677/XUSED  (
    .I(\CHOICE5677/FROM ),
    .O(CHOICE5677)
  );
  X_BUF \CHOICE5677/YUSED  (
    .I(\CHOICE5677/GROM ),
    .O(CHOICE5679)
  );
  defparam \DLX_EXinst__n0007<28>13 .INIT = 16'h88C8;
  X_LUT4 \DLX_EXinst__n0007<28>13  (
    .ADR0(DLX_EXinst__n0053),
    .ADR1(DLX_IDinst_reg_out_A[28]),
    .ADR2(DLX_EXinst__n0054),
    .ADR3(\DLX_IDinst_Imm[31] ),
    .O(\CHOICE4850/FROM )
  );
  defparam \DLX_EXinst__n0007<16>258 .INIT = 16'hC0E0;
  X_LUT4 \DLX_EXinst__n0007<16>258  (
    .ADR0(DLX_EXinst__n0054),
    .ADR1(DLX_EXinst__n0053),
    .ADR2(DLX_IDinst_reg_out_A[16]),
    .ADR3(\DLX_IDinst_Imm[31] ),
    .O(\CHOICE4850/GROM )
  );
  X_BUF \CHOICE4850/XUSED  (
    .I(\CHOICE4850/FROM ),
    .O(CHOICE4850)
  );
  X_BUF \CHOICE4850/YUSED  (
    .I(\CHOICE4850/GROM ),
    .O(CHOICE4614)
  );
  defparam \DLX_EXinst__n0007<17>109 .INIT = 16'hF222;
  X_LUT4 \DLX_EXinst__n0007<17>109  (
    .ADR0(N163635),
    .ADR1(N146478),
    .ADR2(N147520),
    .ADR3(N138037),
    .O(\CHOICE5383/FROM )
  );
  defparam \DLX_EXinst__n0007<17>136 .INIT = 16'hD5C0;
  X_LUT4 \DLX_EXinst__n0007<17>136  (
    .ADR0(\DLX_IDinst_Imm[4] ),
    .ADR1(N163631),
    .ADR2(\DLX_IDinst_Imm[31] ),
    .ADR3(CHOICE5383),
    .O(\CHOICE5383/GROM )
  );
  X_BUF \CHOICE5383/XUSED  (
    .I(\CHOICE5383/FROM ),
    .O(CHOICE5383)
  );
  X_BUF \CHOICE5383/YUSED  (
    .I(\CHOICE5383/GROM ),
    .O(CHOICE5385)
  );
  defparam \DLX_EXinst__n0007<20>95 .INIT = 16'hC4C0;
  X_LUT4 \DLX_EXinst__n0007<20>95  (
    .ADR0(\DLX_IDinst_Imm[31] ),
    .ADR1(DLX_IDinst_reg_out_A[20]),
    .ADR2(DLX_EXinst__n0053),
    .ADR3(DLX_EXinst__n0054),
    .O(\DLX_IDinst_RegFile_22_16/FROM )
  );
  defparam \DLX_EXinst__n0007<24>269 .INIT = 16'hF400;
  X_LUT4 \DLX_EXinst__n0007<24>269  (
    .ADR0(\DLX_IDinst_Imm[31] ),
    .ADR1(DLX_EXinst__n0054),
    .ADR2(DLX_EXinst__n0053),
    .ADR3(DLX_IDinst_reg_out_A[24]),
    .O(\DLX_IDinst_RegFile_22_16/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_22_16/XUSED  (
    .I(\DLX_IDinst_RegFile_22_16/FROM ),
    .O(CHOICE4653)
  );
  X_BUF \DLX_IDinst_RegFile_22_16/YUSED  (
    .I(\DLX_IDinst_RegFile_22_16/GROM ),
    .O(CHOICE5639)
  );
  defparam \DLX_EXinst__n0007<8>163_SW0 .INIT = 16'h5410;
  X_LUT4 \DLX_EXinst__n0007<8>163_SW0  (
    .ADR0(\DLX_IDinst_Imm[3] ),
    .ADR1(\DLX_IDinst_Imm[2] ),
    .ADR2(\DLX_EXinst_Mshift__n0022_Sh[24] ),
    .ADR3(\DLX_EXinst_Mshift__n0020_Sh[28] ),
    .O(\N164155/FROM )
  );
  defparam \DLX_EXinst__n0007<24>357 .INIT = 16'hE400;
  X_LUT4 \DLX_EXinst__n0007<24>357  (
    .ADR0(\DLX_IDinst_Imm[2] ),
    .ADR1(\DLX_EXinst_Mshift__n0021_Sh[16] ),
    .ADR2(\DLX_EXinst_Mshift__n0021_Sh[12] ),
    .ADR3(\DLX_IDinst_Imm[3] ),
    .O(\N164155/GROM )
  );
  X_BUF \N164155/XUSED  (
    .I(\N164155/FROM ),
    .O(N164155)
  );
  X_BUF \N164155/YUSED  (
    .I(\N164155/GROM ),
    .O(CHOICE5668)
  );
  defparam \DLX_EXinst__n0007<24>454 .INIT = 16'hFEFA;
  X_LUT4 \DLX_EXinst__n0007<24>454  (
    .ADR0(CHOICE5679),
    .ADR1(DLX_EXinst__n0109),
    .ADR2(N163716),
    .ADR3(DLX_EXinst__n0012[24]),
    .O(\DLX_EXinst_ALU_result<24>/FROM )
  );
  defparam \DLX_EXinst__n0007<24>484 .INIT = 16'h0F0E;
  X_LUT4 \DLX_EXinst__n0007<24>484  (
    .ADR0(CHOICE5639),
    .ADR1(CHOICE5648),
    .ADR2(DLX_EXinst__n0036),
    .ADR3(CHOICE5681),
    .O(CHOICE5683)
  );
  X_BUF \DLX_EXinst_ALU_result<24>/XUSED  (
    .I(\DLX_EXinst_ALU_result<24>/FROM ),
    .O(CHOICE5681)
  );
  defparam \DLX_EXinst__n0007<25>246_SW0 .INIT = 16'hFFB8;
  X_LUT4 \DLX_EXinst__n0007<25>246_SW0  (
    .ADR0(DLX_EXinst__n0077),
    .ADR1(DLX_IDinst_reg_out_B[25]),
    .ADR2(DLX_EXinst__n0079),
    .ADR3(DLX_EXinst_N74245),
    .O(\N163522/FROM )
  );
  defparam \DLX_EXinst__n0007<25>158 .INIT = 16'h8A88;
  X_LUT4 \DLX_EXinst__n0007<25>158  (
    .ADR0(DLX_IDinst_reg_out_B[25]),
    .ADR1(DLX_EXinst__n0078),
    .ADR2(DLX_IDinst_reg_out_A[25]),
    .ADR3(DLX_EXinst__n0079),
    .O(\N163522/GROM )
  );
  X_BUF \N163522/XUSED  (
    .I(\N163522/FROM ),
    .O(N163522)
  );
  X_BUF \N163522/YUSED  (
    .I(\N163522/GROM ),
    .O(CHOICE5091)
  );
  defparam \DLX_EXinst__n0007<25>246 .INIT = 16'hF222;
  X_LUT4 \DLX_EXinst__n0007<25>246  (
    .ADR0(CHOICE5113),
    .ADR1(DLX_IDinst_reg_out_B[4]),
    .ADR2(N163522),
    .ADR3(DLX_IDinst_reg_out_A[25]),
    .O(\DLX_IDinst_RegFile_2_7/FROM )
  );
  defparam \DLX_EXinst__n0007<25>286_SW0 .INIT = 16'hFFC0;
  X_LUT4 \DLX_EXinst__n0007<25>286_SW0  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N75973),
    .ADR2(\DLX_EXinst_Mshift__n0023_Sh[41] ),
    .ADR3(CHOICE5116),
    .O(\DLX_IDinst_RegFile_2_7/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_2_7/XUSED  (
    .I(\DLX_IDinst_RegFile_2_7/FROM ),
    .O(CHOICE5116)
  );
  X_BUF \DLX_IDinst_RegFile_2_7/YUSED  (
    .I(\DLX_IDinst_RegFile_2_7/GROM ),
    .O(N163514)
  );
  defparam \DLX_EXinst__n0007<18>109 .INIT = 16'h88F8;
  X_LUT4 \DLX_EXinst__n0007<18>109  (
    .ADR0(N147520),
    .ADR1(N137608),
    .ADR2(N163424),
    .ADR3(N146478),
    .O(\CHOICE5225/FROM )
  );
  defparam \DLX_EXinst__n0007<18>136 .INIT = 16'hB3A0;
  X_LUT4 \DLX_EXinst__n0007<18>136  (
    .ADR0(N163420),
    .ADR1(\DLX_IDinst_Imm[4] ),
    .ADR2(\DLX_IDinst_Imm[31] ),
    .ADR3(CHOICE5225),
    .O(\CHOICE5225/GROM )
  );
  X_BUF \CHOICE5225/XUSED  (
    .I(\CHOICE5225/FROM ),
    .O(CHOICE5225)
  );
  X_BUF \CHOICE5225/YUSED  (
    .I(\CHOICE5225/GROM ),
    .O(CHOICE5227)
  );
  defparam \DLX_EXinst__n0007<25>286 .INIT = 16'hF0E0;
  X_LUT4 \DLX_EXinst__n0007<25>286  (
    .ADR0(CHOICE5096),
    .ADR1(CHOICE5091),
    .ADR2(DLX_EXinst__n0036),
    .ADR3(N163514),
    .O(\DLX_EXinst_ALU_result<25>/FROM )
  );
  defparam \DLX_EXinst__n0007<25>296 .INIT = 16'hFFA0;
  X_LUT4 \DLX_EXinst__n0007<25>296  (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(VCC),
    .ADR2(CHOICE929),
    .ADR3(CHOICE5119),
    .O(CHOICE5120)
  );
  X_BUF \DLX_EXinst_ALU_result<25>/XUSED  (
    .I(\DLX_EXinst_ALU_result<25>/FROM ),
    .O(CHOICE5119)
  );
  defparam \DLX_EXinst__n0007<17>326_SW0 .INIT = 16'hEFEC;
  X_LUT4 \DLX_EXinst__n0007<17>326_SW0  (
    .ADR0(DLX_EXinst__n0077),
    .ADR1(DLX_EXinst_N74245),
    .ADR2(DLX_IDinst_reg_out_B[17]),
    .ADR3(DLX_EXinst__n0079),
    .O(\N163593/FROM )
  );
  defparam \DLX_EXinst__n0007<17>199 .INIT = 16'hD0C0;
  X_LUT4 \DLX_EXinst__n0007<17>199  (
    .ADR0(DLX_IDinst_reg_out_A[17]),
    .ADR1(DLX_EXinst__n0078),
    .ADR2(DLX_IDinst_reg_out_B[17]),
    .ADR3(DLX_EXinst__n0079),
    .O(\N163593/GROM )
  );
  X_BUF \N163593/XUSED  (
    .I(\N163593/FROM ),
    .O(N163593)
  );
  X_BUF \N163593/YUSED  (
    .I(\N163593/GROM ),
    .O(CHOICE5393)
  );
  defparam \DLX_EXinst__n0007<17>367 .INIT = 16'hFE00;
  X_LUT4 \DLX_EXinst__n0007<17>367  (
    .ADR0(CHOICE5400),
    .ADR1(CHOICE5393),
    .ADR2(N163584),
    .ADR3(DLX_EXinst__n0036),
    .O(\DLX_EXinst_ALU_result<17>/FROM )
  );
  defparam \DLX_EXinst__n0007<17>378 .INIT = 16'hFFC0;
  X_LUT4 \DLX_EXinst__n0007<17>378  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[31]),
    .ADR2(CHOICE929),
    .ADR3(CHOICE5427),
    .O(CHOICE5428)
  );
  X_BUF \DLX_EXinst_ALU_result<17>/XUSED  (
    .I(\DLX_EXinst_ALU_result<17>/FROM ),
    .O(CHOICE5427)
  );
  defparam \DLX_EXinst__n0007<27>170 .INIT = 16'hEAC0;
  X_LUT4 \DLX_EXinst__n0007<27>170  (
    .ADR0(DLX_EXinst__n0012[27]),
    .ADR1(DLX_EXinst_ALU_result[27]),
    .ADR2(N134884),
    .ADR3(DLX_EXinst__n0127),
    .O(\CHOICE4962/FROM )
  );
  defparam \DLX_EXinst__n0007<18>217 .INIT = 16'hECA0;
  X_LUT4 \DLX_EXinst__n0007<18>217  (
    .ADR0(DLX_EXinst_ALU_result[18]),
    .ADR1(DLX_EXinst__n0012[18]),
    .ADR2(N134884),
    .ADR3(DLX_EXinst__n0127),
    .O(\CHOICE4962/GROM )
  );
  X_BUF \CHOICE4962/XUSED  (
    .I(\CHOICE4962/FROM ),
    .O(CHOICE4962)
  );
  X_BUF \CHOICE4962/YUSED  (
    .I(\CHOICE4962/GROM ),
    .O(CHOICE5242)
  );
  defparam \DLX_EXinst__n0007<17>298 .INIT = 16'h8F88;
  X_LUT4 \DLX_EXinst__n0007<17>298  (
    .ADR0(N137859),
    .ADR1(N148609),
    .ADR2(N148323),
    .ADR3(N163598),
    .O(\CHOICE5421/FROM )
  );
  defparam \DLX_EXinst__n0007<17>326 .INIT = 16'hD5C0;
  X_LUT4 \DLX_EXinst__n0007<17>326  (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(N163593),
    .ADR2(DLX_IDinst_reg_out_A[17]),
    .ADR3(CHOICE5421),
    .O(\CHOICE5421/GROM )
  );
  X_BUF \CHOICE5421/XUSED  (
    .I(\CHOICE5421/FROM ),
    .O(CHOICE5421)
  );
  X_BUF \CHOICE5421/YUSED  (
    .I(\CHOICE5421/GROM ),
    .O(CHOICE5424)
  );
  defparam \DLX_EXinst__n0007<19>217 .INIT = 16'hF888;
  X_LUT4 \DLX_EXinst__n0007<19>217  (
    .ADR0(N134884),
    .ADR1(DLX_EXinst_ALU_result[19]),
    .ADR2(DLX_EXinst__n0012[19]),
    .ADR3(DLX_EXinst__n0127),
    .O(\CHOICE5321/FROM )
  );
  defparam \DLX_EXinst__n0007<26>170 .INIT = 16'hEAC0;
  X_LUT4 \DLX_EXinst__n0007<26>170  (
    .ADR0(DLX_EXinst__n0012[26]),
    .ADR1(N134884),
    .ADR2(DLX_EXinst_ALU_result[26]),
    .ADR3(DLX_EXinst__n0127),
    .O(\CHOICE5321/GROM )
  );
  X_BUF \CHOICE5321/XUSED  (
    .I(\CHOICE5321/FROM ),
    .O(CHOICE5321)
  );
  X_BUF \CHOICE5321/YUSED  (
    .I(\CHOICE5321/GROM ),
    .O(CHOICE5029)
  );
  defparam \DLX_EXinst__n0007<31>9 .INIT = 16'h8C88;
  X_LUT4 \DLX_EXinst__n0007<31>9  (
    .ADR0(DLX_EXinst__n0078),
    .ADR1(DLX_IDinst_reg_out_B[31]),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(DLX_EXinst__n0079),
    .O(\DLX_IDinst_RegFile_3_4/FROM )
  );
  defparam \DLX_EXinst__n0007<26>158 .INIT = 16'hC0E0;
  X_LUT4 \DLX_EXinst__n0007<26>158  (
    .ADR0(DLX_EXinst__n0079),
    .ADR1(DLX_EXinst__n0078),
    .ADR2(DLX_IDinst_reg_out_B[26]),
    .ADR3(DLX_IDinst_reg_out_A[26]),
    .O(\DLX_IDinst_RegFile_3_4/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_3_4/XUSED  (
    .I(\DLX_IDinst_RegFile_3_4/FROM ),
    .O(CHOICE5764)
  );
  X_BUF \DLX_IDinst_RegFile_3_4/YUSED  (
    .I(\DLX_IDinst_RegFile_3_4/GROM ),
    .O(CHOICE5024)
  );
  defparam \DLX_EXinst__n0007<26>246 .INIT = 16'hAE0C;
  X_LUT4 \DLX_EXinst__n0007<26>246  (
    .ADR0(DLX_IDinst_reg_out_A[26]),
    .ADR1(CHOICE5046),
    .ADR2(DLX_IDinst_reg_out_B[4]),
    .ADR3(N163672),
    .O(\CHOICE5049/FROM )
  );
  defparam \DLX_EXinst__n0007<26>286_SW0 .INIT = 16'hFFA0;
  X_LUT4 \DLX_EXinst__n0007<26>286_SW0  (
    .ADR0(\DLX_EXinst_Mshift__n0023_Sh[42] ),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N75973),
    .ADR3(CHOICE5049),
    .O(\CHOICE5049/GROM )
  );
  X_BUF \CHOICE5049/XUSED  (
    .I(\CHOICE5049/FROM ),
    .O(CHOICE5049)
  );
  X_BUF \CHOICE5049/YUSED  (
    .I(\CHOICE5049/GROM ),
    .O(N163660)
  );
  defparam \DLX_EXinst__n0007<19>109 .INIT = 16'h8F88;
  X_LUT4 \DLX_EXinst__n0007<19>109  (
    .ADR0(N147520),
    .ADR1(N138713),
    .ADR2(N146478),
    .ADR3(N163558),
    .O(\CHOICE5304/FROM )
  );
  defparam \DLX_EXinst__n0007<19>121 .INIT = 16'h0F00;
  X_LUT4 \DLX_EXinst__n0007<19>121  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(\DLX_IDinst_Imm[4] ),
    .ADR3(CHOICE5304),
    .O(\CHOICE5304/GROM )
  );
  X_BUF \CHOICE5304/XUSED  (
    .I(\CHOICE5304/FROM ),
    .O(CHOICE5304)
  );
  X_BUF \CHOICE5304/YUSED  (
    .I(\CHOICE5304/GROM ),
    .O(CHOICE5305)
  );
  defparam \DLX_EXinst__n0007<26>286 .INIT = 16'hFE00;
  X_LUT4 \DLX_EXinst__n0007<26>286  (
    .ADR0(CHOICE5024),
    .ADR1(CHOICE5029),
    .ADR2(N163660),
    .ADR3(DLX_EXinst__n0036),
    .O(\DLX_EXinst_ALU_result<26>/FROM )
  );
  defparam \DLX_EXinst__n0007<26>296 .INIT = 16'hFFC0;
  X_LUT4 \DLX_EXinst__n0007<26>296  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[31]),
    .ADR2(CHOICE929),
    .ADR3(CHOICE5052),
    .O(CHOICE5053)
  );
  X_BUF \DLX_EXinst_ALU_result<26>/XUSED  (
    .I(\DLX_EXinst_ALU_result<26>/FROM ),
    .O(CHOICE5052)
  );
  defparam \DLX_EXinst__n0007<18>326_SW0 .INIT = 16'hEFEC;
  X_LUT4 \DLX_EXinst__n0007<18>326_SW0  (
    .ADR0(DLX_EXinst__n0077),
    .ADR1(DLX_EXinst_N74245),
    .ADR2(DLX_IDinst_reg_out_B[18]),
    .ADR3(DLX_EXinst__n0079),
    .O(\N163294/FROM )
  );
  defparam \DLX_EXinst__n0007<18>199 .INIT = 16'hBA00;
  X_LUT4 \DLX_EXinst__n0007<18>199  (
    .ADR0(DLX_EXinst__n0078),
    .ADR1(DLX_IDinst_reg_out_A[18]),
    .ADR2(DLX_EXinst__n0079),
    .ADR3(DLX_IDinst_reg_out_B[18]),
    .O(\N163294/GROM )
  );
  X_BUF \N163294/XUSED  (
    .I(\N163294/FROM ),
    .O(N163294)
  );
  X_BUF \N163294/YUSED  (
    .I(\N163294/GROM ),
    .O(CHOICE5235)
  );
  defparam \DLX_EXinst__n0007<18>367 .INIT = 16'hAAA8;
  X_LUT4 \DLX_EXinst__n0007<18>367  (
    .ADR0(DLX_EXinst__n0036),
    .ADR1(CHOICE5235),
    .ADR2(N163290),
    .ADR3(CHOICE5242),
    .O(\DLX_EXinst_ALU_result<18>/FROM )
  );
  defparam \DLX_EXinst__n0007<18>378 .INIT = 16'hFF88;
  X_LUT4 \DLX_EXinst__n0007<18>378  (
    .ADR0(CHOICE929),
    .ADR1(DLX_IDinst_reg_out_A[31]),
    .ADR2(VCC),
    .ADR3(CHOICE5269),
    .O(CHOICE5270)
  );
  X_BUF \DLX_EXinst_ALU_result<18>/XUSED  (
    .I(\DLX_EXinst_ALU_result<18>/FROM ),
    .O(CHOICE5269)
  );
  defparam \DLX_EXinst__n0007<18>298 .INIT = 16'hF222;
  X_LUT4 \DLX_EXinst__n0007<18>298  (
    .ADR0(N163302),
    .ADR1(N148323),
    .ADR2(N148609),
    .ADR3(N137372),
    .O(\CHOICE5263/FROM )
  );
  defparam \DLX_EXinst__n0007<18>326 .INIT = 16'hD5C0;
  X_LUT4 \DLX_EXinst__n0007<18>326  (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(DLX_IDinst_reg_out_A[18]),
    .ADR2(N163294),
    .ADR3(CHOICE5263),
    .O(\CHOICE5263/GROM )
  );
  X_BUF \CHOICE5263/XUSED  (
    .I(\CHOICE5263/FROM ),
    .O(CHOICE5263)
  );
  X_BUF \CHOICE5263/YUSED  (
    .I(\CHOICE5263/GROM ),
    .O(CHOICE5266)
  );
  defparam \DLX_EXinst__n0007<19>149 .INIT = 16'hFEFA;
  X_LUT4 \DLX_EXinst__n0007<19>149  (
    .ADR0(N163338),
    .ADR1(DLX_EXinst__n0109),
    .ADR2(CHOICE5305),
    .ADR3(DLX_EXinst__n0012[19]),
    .O(\CHOICE5307/FROM )
  );
  defparam \DLX_EXinst__n0007<19>179 .INIT = 16'h0F0E;
  X_LUT4 \DLX_EXinst__n0007<19>179  (
    .ADR0(CHOICE5275),
    .ADR1(CHOICE5278),
    .ADR2(DLX_EXinst__n0036),
    .ADR3(CHOICE5307),
    .O(\CHOICE5307/GROM )
  );
  X_BUF \CHOICE5307/XUSED  (
    .I(\CHOICE5307/FROM ),
    .O(CHOICE5307)
  );
  X_BUF \CHOICE5307/YUSED  (
    .I(\CHOICE5307/GROM ),
    .O(CHOICE5310)
  );
  defparam \DLX_EXinst__n0007<19>326 .INIT = 16'hA0EC;
  X_LUT4 \DLX_EXinst__n0007<19>326  (
    .ADR0(N163684),
    .ADR1(CHOICE5342),
    .ADR2(DLX_IDinst_reg_out_A[19]),
    .ADR3(DLX_IDinst_reg_out_B[4]),
    .O(\CHOICE5345/FROM )
  );
  defparam \DLX_EXinst__n0007<19>367_SW0 .INIT = 16'hFF40;
  X_LUT4 \DLX_EXinst__n0007<19>367_SW0  (
    .ADR0(DLX_EXinst_N72822),
    .ADR1(\DLX_EXinst_Mshift__n0023_Sh[3] ),
    .ADR2(DLX_EXinst_N75973),
    .ADR3(CHOICE5345),
    .O(\CHOICE5345/GROM )
  );
  X_BUF \CHOICE5345/XUSED  (
    .I(\CHOICE5345/FROM ),
    .O(CHOICE5345)
  );
  X_BUF \CHOICE5345/YUSED  (
    .I(\CHOICE5345/GROM ),
    .O(N163676)
  );
  defparam \DLX_EXinst__n0007<27>246_SW0 .INIT = 16'hFAEE;
  X_LUT4 \DLX_EXinst__n0007<27>246_SW0  (
    .ADR0(DLX_EXinst_N74245),
    .ADR1(DLX_EXinst__n0079),
    .ADR2(DLX_EXinst__n0077),
    .ADR3(DLX_IDinst_reg_out_B[27]),
    .O(\N163412/FROM )
  );
  defparam \DLX_EXinst__n0007<27>158 .INIT = 16'hAA08;
  X_LUT4 \DLX_EXinst__n0007<27>158  (
    .ADR0(DLX_IDinst_reg_out_B[27]),
    .ADR1(DLX_EXinst__n0079),
    .ADR2(DLX_IDinst_reg_out_A[27]),
    .ADR3(DLX_EXinst__n0078),
    .O(\N163412/GROM )
  );
  X_BUF \N163412/XUSED  (
    .I(\N163412/FROM ),
    .O(N163412)
  );
  X_BUF \N163412/YUSED  (
    .I(\N163412/GROM ),
    .O(CHOICE4957)
  );
  defparam \DLX_EXinst__n0007<27>246 .INIT = 16'hD5C0;
  X_LUT4 \DLX_EXinst__n0007<27>246  (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(DLX_IDinst_reg_out_A[27]),
    .ADR2(N163412),
    .ADR3(CHOICE4979),
    .O(\CHOICE4982/FROM )
  );
  defparam \DLX_EXinst__n0007<27>286_SW0 .INIT = 16'hFFA0;
  X_LUT4 \DLX_EXinst__n0007<27>286_SW0  (
    .ADR0(DLX_EXinst_N75973),
    .ADR1(VCC),
    .ADR2(\DLX_EXinst_Mshift__n0023_Sh[43] ),
    .ADR3(CHOICE4982),
    .O(\CHOICE4982/GROM )
  );
  X_BUF \CHOICE4982/XUSED  (
    .I(\CHOICE4982/FROM ),
    .O(CHOICE4982)
  );
  X_BUF \CHOICE4982/YUSED  (
    .I(\CHOICE4982/GROM ),
    .O(N163399)
  );
  defparam DLX_IDinst_RegFile_18_17_510.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_18_17_510 (
    .I(DLX_IDinst_WB_data_eff[17]),
    .CE(DLX_IDinst__n0586),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_18_17)
  );
  defparam \DLX_EXinst_Mshift__n0020_Sh<27>_SW0 .INIT = 16'hFC30;
  X_LUT4 \DLX_EXinst_Mshift__n0020_Sh<27>_SW0  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_Imm_0_1),
    .ADR2(DLX_IDinst_reg_out_A[27]),
    .ADR3(DLX_IDinst_reg_out_A[28]),
    .O(\N130467/FROM )
  );
  defparam \DLX_EXinst__n0007<28>221 .INIT = 16'hC0CA;
  X_LUT4 \DLX_EXinst__n0007<28>221  (
    .ADR0(DLX_IDinst_reg_out_A[28]),
    .ADR1(\DLX_EXinst_Mshift__n0023_Sh[24] ),
    .ADR2(DLX_IDinst_reg_out_B[2]),
    .ADR3(DLX_EXinst_N73239),
    .O(\N130467/GROM )
  );
  X_BUF \N130467/XUSED  (
    .I(\N130467/FROM ),
    .O(N130467)
  );
  X_BUF \N130467/YUSED  (
    .I(\N130467/GROM ),
    .O(CHOICE4896)
  );
  defparam \DLX_EXinst__n0007<28>302 .INIT = 16'hEAC0;
  X_LUT4 \DLX_EXinst__n0007<28>302  (
    .ADR0(DLX_IDinst_reg_out_A[28]),
    .ADR1(N134884),
    .ADR2(DLX_EXinst_ALU_result[28]),
    .ADR3(CHOICE4908),
    .O(\CHOICE4910/FROM )
  );
  defparam \DLX_EXinst__n0007<28>308 .INIT = 16'hFFF0;
  X_LUT4 \DLX_EXinst__n0007<28>308  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(CHOICE4902),
    .ADR3(CHOICE4910),
    .O(\CHOICE4910/GROM )
  );
  X_BUF \CHOICE4910/XUSED  (
    .I(\CHOICE4910/FROM ),
    .O(CHOICE4910)
  );
  X_BUF \CHOICE4910/YUSED  (
    .I(\CHOICE4910/GROM ),
    .O(CHOICE4911)
  );
  defparam \DLX_EXinst__n0007<27>286 .INIT = 16'hF0E0;
  X_LUT4 \DLX_EXinst__n0007<27>286  (
    .ADR0(CHOICE4962),
    .ADR1(CHOICE4957),
    .ADR2(DLX_EXinst__n0036),
    .ADR3(N163399),
    .O(\DLX_EXinst_ALU_result<27>/FROM )
  );
  defparam \DLX_EXinst__n0007<27>296 .INIT = 16'hFFA0;
  X_LUT4 \DLX_EXinst__n0007<27>296  (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(VCC),
    .ADR2(CHOICE929),
    .ADR3(CHOICE4985),
    .O(CHOICE4986)
  );
  X_BUF \DLX_EXinst_ALU_result<27>/XUSED  (
    .I(\DLX_EXinst_ALU_result<27>/FROM ),
    .O(CHOICE4985)
  );
  defparam \DLX_EXinst__n0007<19>367 .INIT = 16'hCCC8;
  X_LUT4 \DLX_EXinst__n0007<19>367  (
    .ADR0(CHOICE5321),
    .ADR1(DLX_EXinst__n0036),
    .ADR2(N163676),
    .ADR3(CHOICE5314),
    .O(\DLX_EXinst_ALU_result<19>/FROM )
  );
  defparam \DLX_EXinst__n0007<19>378 .INIT = 16'hFF88;
  X_LUT4 \DLX_EXinst__n0007<19>378  (
    .ADR0(CHOICE929),
    .ADR1(DLX_IDinst_reg_out_A[31]),
    .ADR2(VCC),
    .ADR3(CHOICE5348),
    .O(CHOICE5349)
  );
  X_BUF \DLX_EXinst_ALU_result<19>/XUSED  (
    .I(\DLX_EXinst_ALU_result<19>/FROM ),
    .O(CHOICE5348)
  );
  defparam \DLX_EXinst__n0007<19>326_SW0 .INIT = 16'hEFEA;
  X_LUT4 \DLX_EXinst__n0007<19>326_SW0  (
    .ADR0(DLX_EXinst_N74245),
    .ADR1(DLX_EXinst__n0077),
    .ADR2(DLX_IDinst_reg_out_B[19]),
    .ADR3(DLX_EXinst__n0079),
    .O(\N163684/FROM )
  );
  defparam \DLX_EXinst__n0007<19>199 .INIT = 16'hC0C8;
  X_LUT4 \DLX_EXinst__n0007<19>199  (
    .ADR0(DLX_EXinst__n0079),
    .ADR1(DLX_IDinst_reg_out_B[19]),
    .ADR2(DLX_EXinst__n0078),
    .ADR3(DLX_IDinst_reg_out_A[19]),
    .O(\N163684/GROM )
  );
  X_BUF \N163684/XUSED  (
    .I(\N163684/FROM ),
    .O(N163684)
  );
  X_BUF \N163684/YUSED  (
    .I(\N163684/GROM ),
    .O(CHOICE5314)
  );
  defparam \DLX_EXinst__n0007<29>100 .INIT = 16'hFCFC;
  X_LUT4 \DLX_EXinst__n0007<29>100  (
    .ADR0(VCC),
    .ADR1(CHOICE4800),
    .ADR2(CHOICE4792),
    .ADR3(VCC),
    .O(\CHOICE4801/GROM )
  );
  X_BUF \CHOICE4801/YUSED  (
    .I(\CHOICE4801/GROM ),
    .O(CHOICE4801)
  );
  defparam DLX_IDinst_RegFile_26_25_511.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_26_25_511 (
    .I(DLX_IDinst_WB_data_eff[25]),
    .CE(DLX_IDinst__n0602),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_26_25)
  );
  defparam \DLX_EXinst__n0007<28>370 .INIT = 16'hFEFA;
  X_LUT4 \DLX_EXinst__n0007<28>370  (
    .ADR0(CHOICE4914),
    .ADR1(CHOICE4912),
    .ADR2(CHOICE4918),
    .ADR3(DLX_EXinst__n0036),
    .O(\DLX_EXinst_ALU_result<28>/FROM )
  );
  defparam \DLX_EXinst__n0007<28>3841 .INIT = 16'hFF0C;
  X_LUT4 \DLX_EXinst__n0007<28>3841  (
    .ADR0(VCC),
    .ADR1(CHOICE4876),
    .ADR2(DLX_EXinst__n0036),
    .ADR3(CHOICE4919),
    .O(N162804)
  );
  X_BUF \DLX_EXinst_ALU_result<28>/XUSED  (
    .I(\DLX_EXinst_ALU_result<28>/FROM ),
    .O(CHOICE4919)
  );
  defparam \DLX_EXinst_Mshift__n0019_Sh<12>1 .INIT = 16'hCCAA;
  X_LUT4 \DLX_EXinst_Mshift__n0019_Sh<12>1  (
    .ADR0(DLX_EXinst_N73389),
    .ADR1(DLX_EXinst_N73043),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[0]),
    .O(\DLX_EXinst_Mshift__n0019_Sh<12>/FROM )
  );
  defparam DLX_EXinst_Ker7443439.INIT = 16'hCCFA;
  X_LUT4 DLX_EXinst_Ker7443439 (
    .ADR0(N163136),
    .ADR1(\DLX_EXinst_Mshift__n0019_Sh[12] ),
    .ADR2(CHOICE1749),
    .ADR3(DLX_IDinst_reg_out_B_3_1),
    .O(\DLX_EXinst_Mshift__n0019_Sh<12>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0019_Sh<12>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0019_Sh<12>/FROM ),
    .O(\DLX_EXinst_Mshift__n0019_Sh[12] )
  );
  X_BUF \DLX_EXinst_Mshift__n0019_Sh<12>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0019_Sh<12>/GROM ),
    .O(N137448)
  );
  defparam \DLX_EXinst__n0007<5>13 .INIT = 16'hEFEA;
  X_LUT4 \DLX_EXinst__n0007<5>13  (
    .ADR0(DLX_EXinst_N74245),
    .ADR1(DLX_EXinst__n0077),
    .ADR2(DLX_IDinst_reg_out_B[5]),
    .ADR3(DLX_EXinst__n0079),
    .O(\CHOICE3939/FROM )
  );
  defparam \DLX_EXinst__n0007<28>293 .INIT = 16'hFEAE;
  X_LUT4 \DLX_EXinst__n0007<28>293  (
    .ADR0(DLX_EXinst_N74245),
    .ADR1(DLX_EXinst__n0079),
    .ADR2(DLX_IDinst_reg_out_B[28]),
    .ADR3(DLX_EXinst__n0077),
    .O(\CHOICE3939/GROM )
  );
  X_BUF \CHOICE3939/XUSED  (
    .I(\CHOICE3939/FROM ),
    .O(CHOICE3939)
  );
  X_BUF \CHOICE3939/YUSED  (
    .I(\CHOICE3939/GROM ),
    .O(CHOICE4908)
  );
  defparam DLX_EXinst_Ker763801.INIT = 16'h00F0;
  X_LUT4 DLX_EXinst_Ker763801 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(DLX_IDinst_Imm_3_1),
    .O(\DLX_EXinst_N76382/FROM )
  );
  defparam \DLX_EXinst__n0007<29>143 .INIT = 16'hECA0;
  X_LUT4 \DLX_EXinst__n0007<29>143  (
    .ADR0(DLX_EXinst_N73959),
    .ADR1(CHOICE929),
    .ADR2(DLX_EXinst__n0012[29]),
    .ADR3(DLX_IDinst_reg_out_A[31]),
    .O(\DLX_EXinst_N76382/GROM )
  );
  X_BUF \DLX_EXinst_N76382/XUSED  (
    .I(\DLX_EXinst_N76382/FROM ),
    .O(DLX_EXinst_N76382)
  );
  X_BUF \DLX_EXinst_N76382/YUSED  (
    .I(\DLX_EXinst_N76382/GROM ),
    .O(CHOICE4805)
  );
  defparam \DLX_EXinst_Mshift__n0019_Sh<21>1 .INIT = 16'hF0AA;
  X_LUT4 \DLX_EXinst_Mshift__n0019_Sh<21>1  (
    .ADR0(DLX_EXinst_N73063),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N73414),
    .ADR3(DLX_IDinst_reg_out_B[0]),
    .O(\DLX_IDinst_RegFile_1_17/FROM )
  );
  defparam DLX_EXinst_Ker730911.INIT = 16'hF3C0;
  X_LUT4 DLX_EXinst_Ker730911 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_B[3]),
    .ADR2(\DLX_EXinst_Mshift__n0024_Sh[29] ),
    .ADR3(\DLX_EXinst_Mshift__n0019_Sh[21] ),
    .O(\DLX_IDinst_RegFile_1_17/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_1_17/XUSED  (
    .I(\DLX_IDinst_RegFile_1_17/FROM ),
    .O(\DLX_EXinst_Mshift__n0019_Sh[21] )
  );
  X_BUF \DLX_IDinst_RegFile_1_17/YUSED  (
    .I(\DLX_IDinst_RegFile_1_17/GROM ),
    .O(DLX_EXinst_N73093)
  );
  defparam \DLX_EXinst__n0007<13>13 .INIT = 16'hDC00;
  X_LUT4 \DLX_EXinst__n0007<13>13  (
    .ADR0(DLX_IDinst_reg_out_A[13]),
    .ADR1(DLX_EXinst__n0078),
    .ADR2(DLX_EXinst__n0079),
    .ADR3(DLX_IDinst_reg_out_B[13]),
    .O(\CHOICE3711/FROM )
  );
  defparam \DLX_EXinst__n0007<29>170 .INIT = 16'hAE00;
  X_LUT4 \DLX_EXinst__n0007<29>170  (
    .ADR0(DLX_EXinst__n0078),
    .ADR1(DLX_EXinst__n0079),
    .ADR2(DLX_IDinst_reg_out_A[29]),
    .ADR3(DLX_IDinst_reg_out_B[29]),
    .O(\CHOICE3711/GROM )
  );
  X_BUF \CHOICE3711/XUSED  (
    .I(\CHOICE3711/FROM ),
    .O(CHOICE3711)
  );
  X_BUF \CHOICE3711/YUSED  (
    .I(\CHOICE3711/GROM ),
    .O(CHOICE4812)
  );
  defparam \DLX_EXinst_Mshift__n0019_Sh<30>1 .INIT = 16'hAAAC;
  X_LUT4 \DLX_EXinst_Mshift__n0019_Sh<30>1  (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(DLX_IDinst_reg_out_A[30]),
    .ADR2(DLX_IDinst_reg_out_B[1]),
    .ADR3(DLX_IDinst_reg_out_B[0]),
    .O(\DLX_EXinst_Mshift__n0019_Sh<30>/FROM )
  );
  defparam DLX_EXinst_Ker7495426.INIT = 16'h0E04;
  X_LUT4 DLX_EXinst_Ker7495426 (
    .ADR0(DLX_IDinst_reg_out_B_2_1),
    .ADR1(\DLX_EXinst_Mshift__n0019_Sh[26] ),
    .ADR2(DLX_IDinst_reg_out_B[5]),
    .ADR3(\DLX_EXinst_Mshift__n0019_Sh[30] ),
    .O(\DLX_EXinst_Mshift__n0019_Sh<30>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0019_Sh<30>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0019_Sh<30>/FROM ),
    .O(\DLX_EXinst_Mshift__n0019_Sh[30] )
  );
  X_BUF \DLX_EXinst_Mshift__n0019_Sh<30>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0019_Sh<30>/GROM ),
    .O(CHOICE1883)
  );
  defparam \DLX_EXinst__n0007<29>251 .INIT = 16'hECA0;
  X_LUT4 \DLX_EXinst__n0007<29>251  (
    .ADR0(DLX_EXinst_ALU_result[29]),
    .ADR1(DLX_IDinst_reg_out_A[29]),
    .ADR2(N134884),
    .ADR3(CHOICE4831),
    .O(\CHOICE4833/FROM )
  );
  defparam \DLX_EXinst__n0007<29>257 .INIT = 16'hFFCC;
  X_LUT4 \DLX_EXinst__n0007<29>257  (
    .ADR0(VCC),
    .ADR1(CHOICE4825),
    .ADR2(VCC),
    .ADR3(CHOICE4833),
    .O(\CHOICE4833/GROM )
  );
  X_BUF \CHOICE4833/XUSED  (
    .I(\CHOICE4833/FROM ),
    .O(CHOICE4833)
  );
  X_BUF \CHOICE4833/YUSED  (
    .I(\CHOICE4833/GROM ),
    .O(CHOICE4834)
  );
  defparam \DLX_EXinst__n0007<29>318 .INIT = 16'hFEEE;
  X_LUT4 \DLX_EXinst__n0007<29>318  (
    .ADR0(CHOICE4841),
    .ADR1(CHOICE4837),
    .ADR2(DLX_EXinst__n0036),
    .ADR3(CHOICE4835),
    .O(\DLX_EXinst_ALU_result<29>/FROM )
  );
  defparam \DLX_EXinst__n0007<29>3321 .INIT = 16'hFF44;
  X_LUT4 \DLX_EXinst__n0007<29>3321  (
    .ADR0(DLX_EXinst__n0036),
    .ADR1(CHOICE4802),
    .ADR2(VCC),
    .ADR3(CHOICE4842),
    .O(N162835)
  );
  X_BUF \DLX_EXinst_ALU_result<29>/XUSED  (
    .I(\DLX_EXinst_ALU_result<29>/FROM ),
    .O(CHOICE4842)
  );
  defparam \DLX_EXinst__n0007<2>172 .INIT = 16'hF202;
  X_LUT4 \DLX_EXinst__n0007<2>172  (
    .ADR0(DLX_IDinst_reg_out_A[2]),
    .ADR1(DLX_EXinst_N73239),
    .ADR2(DLX_IDinst_reg_out_B[3]),
    .ADR3(\DLX_EXinst_Mshift__n0019_Sh[10] ),
    .O(\CHOICE5550/FROM )
  );
  defparam \DLX_EXinst__n0007<29>185 .INIT = 16'hDC10;
  X_LUT4 \DLX_EXinst__n0007<29>185  (
    .ADR0(DLX_EXinst_N73239),
    .ADR1(DLX_IDinst_reg_out_B[3]),
    .ADR2(DLX_IDinst_reg_out_A[29]),
    .ADR3(\DLX_EXinst_Mshift__n0023_Sh[21] ),
    .O(\CHOICE5550/GROM )
  );
  X_BUF \CHOICE5550/XUSED  (
    .I(\CHOICE5550/FROM ),
    .O(CHOICE5550)
  );
  X_BUF \CHOICE5550/YUSED  (
    .I(\CHOICE5550/GROM ),
    .O(CHOICE4819)
  );
  defparam \DLX_EXinst_Mshift__n0019_Sh<16>1 .INIT = 16'hBB88;
  X_LUT4 \DLX_EXinst_Mshift__n0019_Sh<16>1  (
    .ADR0(DLX_EXinst_N73053),
    .ADR1(DLX_IDinst_reg_out_B[0]),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N73399),
    .O(\DLX_EXinst_Mshift__n0019_Sh<16>/FROM )
  );
  defparam DLX_EXinst_Ker746891.INIT = 16'hFA0A;
  X_LUT4 DLX_EXinst_Ker746891 (
    .ADR0(\DLX_EXinst_Mshift__n0019_Sh[8] ),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B_3_1),
    .ADR3(\DLX_EXinst_Mshift__n0019_Sh[16] ),
    .O(\DLX_EXinst_Mshift__n0019_Sh<16>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0019_Sh<16>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0019_Sh<16>/FROM ),
    .O(\DLX_EXinst_Mshift__n0019_Sh[16] )
  );
  X_BUF \DLX_EXinst_Mshift__n0019_Sh<16>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0019_Sh<16>/GROM ),
    .O(DLX_EXinst_N74691)
  );
  defparam DLX_EXinst_Ker76159158_SW0.INIT = 16'hDDFF;
  X_LUT4 DLX_EXinst_Ker76159158_SW0 (
    .ADR0(DLX_EXinst_N76041),
    .ADR1(\DLX_IDinst_Imm[31] ),
    .ADR2(VCC),
    .ADR3(CHOICE3451),
    .O(\N163148/FROM )
  );
  defparam DLX_EXinst_Ker76159158.INIT = 16'h0020;
  X_LUT4 DLX_EXinst_Ker76159158 (
    .ADR0(DLX_IDinst_IR_opcode_field[1]),
    .ADR1(\DLX_IDinst_Imm[6] ),
    .ADR2(DLX_IDinst_IR_opcode_field[0]),
    .ADR3(N163148),
    .O(\N163148/GROM )
  );
  X_BUF \N163148/XUSED  (
    .I(\N163148/FROM ),
    .O(N163148)
  );
  X_BUF \N163148/YUSED  (
    .I(\N163148/GROM ),
    .O(N147520)
  );
  defparam \DLX_EXinst_Mshift__n0019_Sh<17>1 .INIT = 16'hCCF0;
  X_LUT4 \DLX_EXinst_Mshift__n0019_Sh<17>1  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N73404),
    .ADR2(DLX_EXinst_N73053),
    .ADR3(DLX_IDinst_reg_out_B[0]),
    .O(\DLX_IDinst_RegFile_27_29/FROM )
  );
  defparam DLX_EXinst_Ker747241.INIT = 16'hF3C0;
  X_LUT4 DLX_EXinst_Ker747241 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_B_3_1),
    .ADR2(\DLX_EXinst_Mshift__n0019_Sh[25] ),
    .ADR3(\DLX_EXinst_Mshift__n0019_Sh[17] ),
    .O(\DLX_IDinst_RegFile_27_29/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_27_29/XUSED  (
    .I(\DLX_IDinst_RegFile_27_29/FROM ),
    .O(\DLX_EXinst_Mshift__n0019_Sh[17] )
  );
  X_BUF \DLX_IDinst_RegFile_27_29/YUSED  (
    .I(\DLX_IDinst_RegFile_27_29/GROM ),
    .O(DLX_EXinst_N74726)
  );
  defparam \DLX_EXinst_Mshift__n0019_Sh<18>1 .INIT = 16'hD8D8;
  X_LUT4 \DLX_EXinst_Mshift__n0019_Sh<18>1  (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(DLX_EXinst_N73058),
    .ADR2(DLX_EXinst_N73404),
    .ADR3(VCC),
    .O(\DLX_EXinst_Mshift__n0019_Sh<18>/FROM )
  );
  defparam DLX_EXinst_Ker747291.INIT = 16'hAFA0;
  X_LUT4 DLX_EXinst_Ker747291 (
    .ADR0(\DLX_EXinst_Mshift__n0019_Sh[26] ),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B_3_1),
    .ADR3(\DLX_EXinst_Mshift__n0019_Sh[18] ),
    .O(\DLX_EXinst_Mshift__n0019_Sh<18>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0019_Sh<18>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0019_Sh<18>/FROM ),
    .O(\DLX_EXinst_Mshift__n0019_Sh[18] )
  );
  X_BUF \DLX_EXinst_Mshift__n0019_Sh<18>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0019_Sh<18>/GROM ),
    .O(DLX_EXinst_N74731)
  );
  defparam \DLX_EXinst_Mshift__n0019_Sh<19>1 .INIT = 16'hFA0A;
  X_LUT4 \DLX_EXinst_Mshift__n0019_Sh<19>1  (
    .ADR0(DLX_EXinst_N73058),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[0]),
    .ADR3(DLX_EXinst_N73409),
    .O(\DLX_EXinst_Mshift__n0019_Sh<19>/FROM )
  );
  defparam DLX_EXinst_Ker749741.INIT = 16'hBB88;
  X_LUT4 DLX_EXinst_Ker749741 (
    .ADR0(\DLX_EXinst_Mshift__n0019_Sh[27] ),
    .ADR1(DLX_IDinst_reg_out_B_3_1),
    .ADR2(VCC),
    .ADR3(\DLX_EXinst_Mshift__n0019_Sh[19] ),
    .O(\DLX_EXinst_Mshift__n0019_Sh<19>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0019_Sh<19>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0019_Sh<19>/FROM ),
    .O(\DLX_EXinst_Mshift__n0019_Sh[19] )
  );
  X_BUF \DLX_EXinst_Mshift__n0019_Sh<19>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0019_Sh<19>/GROM ),
    .O(DLX_EXinst_N74976)
  );
  defparam \DLX_EXinst_Mshift__n0019_Sh<61>1 .INIT = 16'h5F00;
  X_LUT4 \DLX_EXinst_Mshift__n0019_Sh<61>1  (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[1]),
    .ADR3(DLX_IDinst_reg_out_A[31]),
    .O(\DLX_EXinst_Mshift__n0019_Sh<61>/FROM )
  );
  defparam DLX_EXinst_Ker7495913.INIT = 16'hE020;
  X_LUT4 DLX_EXinst_Ker7495913 (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(DLX_IDinst_reg_out_B_2_1),
    .ADR2(DLX_IDinst_reg_out_B[5]),
    .ADR3(\DLX_EXinst_Mshift__n0019_Sh[61] ),
    .O(\DLX_EXinst_Mshift__n0019_Sh<61>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0019_Sh<61>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0019_Sh<61>/FROM ),
    .O(\DLX_EXinst_Mshift__n0019_Sh[61] )
  );
  X_BUF \DLX_EXinst_Mshift__n0019_Sh<61>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0019_Sh<61>/GROM ),
    .O(CHOICE1933)
  );
  defparam \DLX_EXinst_Mshift__n0019_Sh<29>1 .INIT = 16'hCFC0;
  X_LUT4 \DLX_EXinst_Mshift__n0019_Sh<29>1  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[31]),
    .ADR2(DLX_IDinst_reg_out_B[1]),
    .ADR3(DLX_EXinst_N72803),
    .O(\DLX_IDinst_EPC<6>/FROM )
  );
  defparam DLX_EXinst_Ker7551314.INIT = 16'h0D08;
  X_LUT4 DLX_EXinst_Ker7551314 (
    .ADR0(DLX_EXinst_N72822),
    .ADR1(DLX_IDinst_reg_out_A[31]),
    .ADR2(DLX_IDinst_reg_out_B[5]),
    .ADR3(\DLX_EXinst_Mshift__n0019_Sh[29] ),
    .O(\DLX_IDinst_EPC<6>/GROM )
  );
  X_BUF \DLX_IDinst_EPC<6>/XUSED  (
    .I(\DLX_IDinst_EPC<6>/FROM ),
    .O(\DLX_EXinst_Mshift__n0019_Sh[29] )
  );
  X_BUF \DLX_IDinst_EPC<6>/YUSED  (
    .I(\DLX_IDinst_EPC<6>/GROM ),
    .O(CHOICE2032)
  );
  defparam DLX_IFinst_IR_previous_10.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_10 (
    .I(DLX_IFinst_IR_latched[10]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[10])
  );
  defparam DLX_IFinst_IR_previous_12.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_12 (
    .I(DLX_IFinst_IR_latched[12]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[12])
  );
  defparam DLX_IFinst_IR_previous_14.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_14 (
    .I(DLX_IFinst_IR_latched[14]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[14])
  );
  defparam DLX_IFinst_IR_previous_15.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_15 (
    .I(DLX_IFinst_IR_latched[15]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[15])
  );
  defparam DLX_IFinst_IR_previous_31.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_31 (
    .I(DLX_IFinst_IR_latched[31]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[31])
  );
  defparam DLX_IFinst_IR_previous_25.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_25 (
    .I(DLX_IFinst_IR_latched[25]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[25])
  );
  defparam DLX_IFinst_IR_previous_17.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_17 (
    .I(DLX_IFinst_IR_latched[17]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[17])
  );
  defparam DLX_IFinst_IR_previous_18.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_18 (
    .I(DLX_IFinst_IR_latched[18]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[18])
  );
  defparam DLX_IFinst_IR_previous_27.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_27 (
    .I(DLX_IFinst_IR_latched[27]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[27])
  );
  defparam DLX_EXinst__n0036_512.INIT = 16'h0001;
  X_LUT4 DLX_EXinst__n0036_512 (
    .ADR0(DLX_IDinst_IR_opcode_field[0]),
    .ADR1(DLX_IDinst_IR_opcode_field[1]),
    .ADR2(N132091),
    .ADR3(DLX_IDinst_IR_opcode_field[5]),
    .O(\DLX_EXinst__n0036/FROM )
  );
  defparam DLX_EXinst_Ker764101.INIT = 16'h0001;
  X_LUT4 DLX_EXinst_Ker764101 (
    .ADR0(DLX_IDinst_Imm_2_1),
    .ADR1(DLX_IDinst_Imm_3_1),
    .ADR2(\DLX_IDinst_Imm[4] ),
    .ADR3(DLX_EXinst__n0036),
    .O(\DLX_EXinst__n0036/GROM )
  );
  X_BUF \DLX_EXinst__n0036/XUSED  (
    .I(\DLX_EXinst__n0036/FROM ),
    .O(DLX_EXinst__n0036)
  );
  X_BUF \DLX_EXinst__n0036/YUSED  (
    .I(\DLX_EXinst__n0036/GROM ),
    .O(DLX_EXinst_N76412)
  );
  defparam \DLX_EXinst_Mshift__n0019_Sh<88>1 .INIT = 16'hFA50;
  X_LUT4 \DLX_EXinst_Mshift__n0019_Sh<88>1  (
    .ADR0(DLX_IDinst_reg_out_B_3_1),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N73369),
    .ADR3(DLX_IDinst_reg_out_A[31]),
    .O(\DLX_EXinst_Mshift__n0019_Sh<88>/FROM )
  );
  defparam \DLX_EXinst__n0007<8>72 .INIT = 16'hE2C0;
  X_LUT4 \DLX_EXinst__n0007<8>72  (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(DLX_IDinst_reg_out_B[5]),
    .ADR2(DLX_EXinst_N76388),
    .ADR3(\DLX_EXinst_Mshift__n0019_Sh[88] ),
    .O(\DLX_EXinst_Mshift__n0019_Sh<88>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0019_Sh<88>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0019_Sh<88>/FROM ),
    .O(\DLX_EXinst_Mshift__n0019_Sh[88] )
  );
  X_BUF \DLX_EXinst_Mshift__n0019_Sh<88>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0019_Sh<88>/GROM ),
    .O(CHOICE5146)
  );
  defparam DLX_IDinst_RegFile_26_17_513.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_26_17_513 (
    .I(DLX_IDinst_WB_data_eff[17]),
    .CE(DLX_IDinst__n0602),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_26_17)
  );
  defparam \vga_top_vga1_redout<1>1 .INIT = 16'h0030;
  X_LUT4 \vga_top_vga1_redout<1>1  (
    .ADR0(VCC),
    .ADR1(vram_out_vga_eff),
    .ADR2(vga_top_vga1_videoon),
    .ADR3(reset_IBUF_1),
    .O(\red_1_OBUF/FROM )
  );
  defparam \vga_top_vga1_redout<0>1 .INIT = 16'h0500;
  X_LUT4 \vga_top_vga1_redout<0>1  (
    .ADR0(reset_IBUF_1),
    .ADR1(VCC),
    .ADR2(vram_out_vga_eff),
    .ADR3(vga_top_vga1_videoon),
    .O(\red_1_OBUF/GROM )
  );
  X_BUF \red_1_OBUF/XUSED  (
    .I(\red_1_OBUF/FROM ),
    .O(red_1_OBUF)
  );
  X_BUF \red_1_OBUF/YUSED  (
    .I(\red_1_OBUF/GROM ),
    .O(red_0_OBUF)
  );
  X_ZERO \DLX_IDinst_RegFile_4_0/LOGIC_ZERO_514  (
    .O(\DLX_IDinst_RegFile_4_0/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_2_515 (
    .IA(\DLX_IDinst_RegFile_4_0/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_4_0/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_61),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_2)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_611.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_611 (
    .ADR0(DLX_IDinst_RegFile_4_0),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_45),
    .ADR2(DLX_IDinst_RegFile_5_0),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_61)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_621.INIT = 16'hE2FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_621 (
    .ADR0(DLX_IDinst_RegFile_6_0),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR2(DLX_IDinst_RegFile_7_0),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_46),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_62)
  );
  X_BUF \DLX_IDinst_RegFile_4_0/COUTUSED  (
    .I(\DLX_IDinst_RegFile_4_0/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_3)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_3_516 (
    .IA(\DLX_IDinst_RegFile_4_0/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_2),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_62),
    .O(\DLX_IDinst_RegFile_4_0/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_4_0/CYINIT_517  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_1),
    .O(\DLX_IDinst_RegFile_4_0/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_4_1/LOGIC_ZERO_518  (
    .O(\DLX_IDinst_RegFile_4_1/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_18_519 (
    .IA(\DLX_IDinst_RegFile_4_1/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_4_1/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_77),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_18)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_771.INIT = 16'hB8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_771 (
    .ADR0(DLX_IDinst_RegFile_5_1),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR2(DLX_IDinst_RegFile_4_1),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_45),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_77)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_781.INIT = 16'hF7D5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_781 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_46),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR2(DLX_IDinst_RegFile_7_1),
    .ADR3(DLX_IDinst_RegFile_6_1),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_78)
  );
  X_BUF \DLX_IDinst_RegFile_4_1/COUTUSED  (
    .I(\DLX_IDinst_RegFile_4_1/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_19)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_19_520 (
    .IA(\DLX_IDinst_RegFile_4_1/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_18),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_78),
    .O(\DLX_IDinst_RegFile_4_1/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_4_1/CYINIT_521  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_17),
    .O(\DLX_IDinst_RegFile_4_1/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_4_2/LOGIC_ZERO_522  (
    .O(\DLX_IDinst_RegFile_4_2/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_34_523 (
    .IA(\DLX_IDinst_RegFile_4_2/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_4_2/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_93),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_34)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_931.INIT = 16'hE2FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_931 (
    .ADR0(DLX_IDinst_RegFile_4_2),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR2(DLX_IDinst_RegFile_5_2),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_45),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_93)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_941.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_941 (
    .ADR0(DLX_IDinst_RegFile_6_2),
    .ADR1(DLX_IDinst_RegFile_7_2),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_46),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_94)
  );
  X_BUF \DLX_IDinst_RegFile_4_2/COUTUSED  (
    .I(\DLX_IDinst_RegFile_4_2/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_35)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_35_524 (
    .IA(\DLX_IDinst_RegFile_4_2/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_34),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_94),
    .O(\DLX_IDinst_RegFile_4_2/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_4_2/CYINIT_525  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_33),
    .O(\DLX_IDinst_RegFile_4_2/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_4_3/LOGIC_ZERO_526  (
    .O(\DLX_IDinst_RegFile_4_3/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_50_527 (
    .IA(\DLX_IDinst_RegFile_4_3/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_4_3/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_109),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_50)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1091.INIT = 16'hFD5D;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1091 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_45),
    .ADR1(DLX_IDinst_RegFile_4_3),
    .ADR2(DLX_IDinst_jtarget[16]),
    .ADR3(DLX_IDinst_RegFile_5_3),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_109)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1101.INIT = 16'hDDF5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1101 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_46),
    .ADR1(DLX_IDinst_RegFile_7_3),
    .ADR2(DLX_IDinst_RegFile_6_3),
    .ADR3(DLX_IDinst_jtarget[16]),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_110)
  );
  X_BUF \DLX_IDinst_RegFile_4_3/COUTUSED  (
    .I(\DLX_IDinst_RegFile_4_3/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_51)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_51_528 (
    .IA(\DLX_IDinst_RegFile_4_3/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_50),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_110),
    .O(\DLX_IDinst_RegFile_4_3/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_4_3/CYINIT_529  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_49),
    .O(\DLX_IDinst_RegFile_4_3/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_4_4/LOGIC_ZERO_530  (
    .O(\DLX_IDinst_RegFile_4_4/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_66_531 (
    .IA(\DLX_IDinst_RegFile_4_4/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_4_4/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_125),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_66)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1251.INIT = 16'hDF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1251 (
    .ADR0(DLX_IDinst_jtarget[16]),
    .ADR1(DLX_IDinst_RegFile_5_4),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_45),
    .ADR3(DLX_IDinst_RegFile_4_4),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_125)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1261.INIT = 16'hFD5D;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1261 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_46),
    .ADR1(DLX_IDinst_RegFile_6_4),
    .ADR2(DLX_IDinst_jtarget[16]),
    .ADR3(DLX_IDinst_RegFile_7_4),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_126)
  );
  X_BUF \DLX_IDinst_RegFile_4_4/COUTUSED  (
    .I(\DLX_IDinst_RegFile_4_4/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_67)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_67_532 (
    .IA(\DLX_IDinst_RegFile_4_4/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_66),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_126),
    .O(\DLX_IDinst_RegFile_4_4/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_4_4/CYINIT_533  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_65),
    .O(\DLX_IDinst_RegFile_4_4/CYINIT )
  );
  defparam DLX_IDinst_Ker10825762_SW0.INIT = 16'hB1BB;
  X_LUT4 DLX_IDinst_Ker10825762_SW0 (
    .ADR0(DLX_IFinst_IR_latched[28]),
    .ADR1(DLX_IFinst_IR_latched[30]),
    .ADR2(DLX_IFinst_IR_latched[27]),
    .ADR3(CHOICE3293),
    .O(\DLX_IFinst_IR_previous<30>/FROM )
  );
  defparam DLX_IDinst_Ker10825762.INIT = 16'h00CD;
  X_LUT4 DLX_IDinst_Ker10825762 (
    .ADR0(DLX_IDinst__n0105),
    .ADR1(DLX_IDinst__n0381),
    .ADR2(DLX_IDinst__n0102),
    .ADR3(N163314),
    .O(\DLX_IFinst_IR_previous<30>/GROM )
  );
  X_BUF \DLX_IFinst_IR_previous<30>/XUSED  (
    .I(\DLX_IFinst_IR_previous<30>/FROM ),
    .O(N163314)
  );
  X_BUF \DLX_IFinst_IR_previous<30>/YUSED  (
    .I(\DLX_IFinst_IR_previous<30>/GROM ),
    .O(CHOICE3300)
  );
  defparam DLX_IDinst_RegFile_3_8_534.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_3_8_534 (
    .I(DLX_IDinst_WB_data_eff[8]),
    .CE(DLX_IDinst__n0556),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_3_8)
  );
  X_ZERO \DLX_IDinst_RegFile_5_0/LOGIC_ZERO_535  (
    .O(\DLX_IDinst_RegFile_5_0/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_514_536 (
    .IA(\DLX_IDinst_RegFile_5_0/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_5_0/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_589),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_514)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_5891.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_5891 (
    .ADR0(DLX_IDinst_RegFile_5_0),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_573),
    .ADR2(DLX_IDinst_RegFile_4_0),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_589)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_5901.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_5901 (
    .ADR0(DLX_IDinst_RegFile_7_0),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_574),
    .ADR2(DLX_IDinst_RegFile_6_0),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_590)
  );
  X_BUF \DLX_IDinst_RegFile_5_0/COUTUSED  (
    .I(\DLX_IDinst_RegFile_5_0/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_515)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_515_537 (
    .IA(\DLX_IDinst_RegFile_5_0/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_514),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_590),
    .O(\DLX_IDinst_RegFile_5_0/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_5_0/CYINIT_538  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_513),
    .O(\DLX_IDinst_RegFile_5_0/CYINIT )
  );
  defparam \DLX_IFinst__n0001<0>_SW0 .INIT = 16'h3535;
  X_LUT4 \DLX_IFinst__n0001<0>_SW0  (
    .ADR0(DLX_IFinst_NPC[0]),
    .ADR1(DLX_IFinst_PC[0]),
    .ADR2(DLX_IFinst__n0000),
    .ADR3(VCC),
    .O(\DLX_IFinst_NPC<0>/FROM )
  );
  defparam \DLX_IFinst__n0001<0> .INIT = 16'hA0AF;
  X_LUT4 \DLX_IFinst__n0001<0>  (
    .ADR0(DLX_IDinst_branch_address[0]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(N128287),
    .O(\DLX_IFinst_NPC<0>/GROM )
  );
  X_BUF \DLX_IFinst_NPC<0>/XUSED  (
    .I(\DLX_IFinst_NPC<0>/FROM ),
    .O(N128287)
  );
  X_BUF \DLX_IFinst_NPC<0>/YUSED  (
    .I(\DLX_IFinst_NPC<0>/GROM ),
    .O(DLX_IFinst__n0001[0])
  );
  X_ZERO \DLX_IDinst_RegFile_4_5/LOGIC_ZERO_539  (
    .O(\DLX_IDinst_RegFile_4_5/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_82_540 (
    .IA(\DLX_IDinst_RegFile_4_5/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_4_5/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_141),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_82)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1411.INIT = 16'hB8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1411 (
    .ADR0(DLX_IDinst_RegFile_5_5),
    .ADR1(DLX_IDinst_jtarget[16]),
    .ADR2(DLX_IDinst_RegFile_4_5),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_45),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_141)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1421.INIT = 16'hB8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1421 (
    .ADR0(DLX_IDinst_RegFile_7_5),
    .ADR1(DLX_IDinst_jtarget[16]),
    .ADR2(DLX_IDinst_RegFile_6_5),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_46),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_142)
  );
  X_BUF \DLX_IDinst_RegFile_4_5/COUTUSED  (
    .I(\DLX_IDinst_RegFile_4_5/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_83)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_83_541 (
    .IA(\DLX_IDinst_RegFile_4_5/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_82),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_142),
    .O(\DLX_IDinst_RegFile_4_5/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_4_5/CYINIT_542  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_81),
    .O(\DLX_IDinst_RegFile_4_5/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_5_1/LOGIC_ZERO_543  (
    .O(\DLX_IDinst_RegFile_5_1/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_530_544 (
    .IA(\DLX_IDinst_RegFile_5_1/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_5_1/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_605),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_530)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6051.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6051 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR1(DLX_IDinst_RegFile_4_1),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_573),
    .ADR3(DLX_IDinst_RegFile_5_1),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_605)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6061.INIT = 16'hE4FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6061 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR1(DLX_IDinst_RegFile_6_1),
    .ADR2(DLX_IDinst_RegFile_7_1),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_574),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_606)
  );
  X_BUF \DLX_IDinst_RegFile_5_1/COUTUSED  (
    .I(\DLX_IDinst_RegFile_5_1/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_531)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_531_545 (
    .IA(\DLX_IDinst_RegFile_5_1/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_530),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_606),
    .O(\DLX_IDinst_RegFile_5_1/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_5_1/CYINIT_546  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_529),
    .O(\DLX_IDinst_RegFile_5_1/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_4_6/LOGIC_ZERO_547  (
    .O(\DLX_IDinst_RegFile_4_6/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_98_548 (
    .IA(\DLX_IDinst_RegFile_4_6/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_4_6/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_157),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_98)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1571.INIT = 16'hBFB3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1571 (
    .ADR0(DLX_IDinst_RegFile_5_6),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_45),
    .ADR2(DLX_IDinst_jtarget[16]),
    .ADR3(DLX_IDinst_RegFile_4_6),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_157)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1581.INIT = 16'hACFF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1581 (
    .ADR0(DLX_IDinst_RegFile_7_6),
    .ADR1(DLX_IDinst_RegFile_6_6),
    .ADR2(DLX_IDinst_jtarget[16]),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_46),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_158)
  );
  X_BUF \DLX_IDinst_RegFile_4_6/COUTUSED  (
    .I(\DLX_IDinst_RegFile_4_6/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_99)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_99_549 (
    .IA(\DLX_IDinst_RegFile_4_6/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_98),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_158),
    .O(\DLX_IDinst_RegFile_4_6/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_4_6/CYINIT_550  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_97),
    .O(\DLX_IDinst_RegFile_4_6/CYINIT )
  );
  defparam DLX_IDinst_RegFile_18_18_551.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_18_18_551 (
    .I(DLX_IDinst_WB_data_eff[18]),
    .CE(DLX_IDinst__n0586),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_18_18)
  );
  X_ZERO \DLX_IDinst_RegFile_5_2/LOGIC_ZERO_552  (
    .O(\DLX_IDinst_RegFile_5_2/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_546_553 (
    .IA(\DLX_IDinst_RegFile_5_2/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_5_2/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_621),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_546)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6211.INIT = 16'hBF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6211 (
    .ADR0(DLX_IDinst_RegFile_5_2),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_573),
    .ADR3(DLX_IDinst_RegFile_4_2),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_621)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6221.INIT = 16'hBFB3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6221 (
    .ADR0(DLX_IDinst_RegFile_7_2),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_574),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR3(DLX_IDinst_RegFile_6_2),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_622)
  );
  X_BUF \DLX_IDinst_RegFile_5_2/COUTUSED  (
    .I(\DLX_IDinst_RegFile_5_2/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_547)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_547_554 (
    .IA(\DLX_IDinst_RegFile_5_2/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_546),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_622),
    .O(\DLX_IDinst_RegFile_5_2/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_5_2/CYINIT_555  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_545),
    .O(\DLX_IDinst_RegFile_5_2/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_4_7/LOGIC_ZERO_556  (
    .O(\DLX_IDinst_RegFile_4_7/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_114_557 (
    .IA(\DLX_IDinst_RegFile_4_7/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_4_7/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_173),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_114)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1731.INIT = 16'hAFCF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1731 (
    .ADR0(DLX_IDinst_RegFile_5_7),
    .ADR1(DLX_IDinst_RegFile_4_7),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_45),
    .ADR3(DLX_IDinst_jtarget[16]),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_173)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1741.INIT = 16'hDDF5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1741 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_46),
    .ADR1(DLX_IDinst_RegFile_7_7),
    .ADR2(DLX_IDinst_RegFile_6_7),
    .ADR3(DLX_IDinst_jtarget[16]),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_174)
  );
  X_BUF \DLX_IDinst_RegFile_4_7/COUTUSED  (
    .I(\DLX_IDinst_RegFile_4_7/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_115)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_115_558 (
    .IA(\DLX_IDinst_RegFile_4_7/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_114),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_174),
    .O(\DLX_IDinst_RegFile_4_7/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_4_7/CYINIT_559  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_113),
    .O(\DLX_IDinst_RegFile_4_7/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_5_3/LOGIC_ZERO_560  (
    .O(\DLX_IDinst_RegFile_5_3/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_562_561 (
    .IA(\DLX_IDinst_RegFile_5_3/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_5_3/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_637),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_562)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6371.INIT = 16'hDF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6371 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR1(DLX_IDinst_RegFile_5_3),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_573),
    .ADR3(DLX_IDinst_RegFile_4_3),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_637)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6381.INIT = 16'hFB73;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6381 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_574),
    .ADR2(DLX_IDinst_RegFile_6_3),
    .ADR3(DLX_IDinst_RegFile_7_3),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_638)
  );
  X_BUF \DLX_IDinst_RegFile_5_3/COUTUSED  (
    .I(\DLX_IDinst_RegFile_5_3/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_563)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_563_562 (
    .IA(\DLX_IDinst_RegFile_5_3/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_562),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_638),
    .O(\DLX_IDinst_RegFile_5_3/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_5_3/CYINIT_563  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_561),
    .O(\DLX_IDinst_RegFile_5_3/CYINIT )
  );
  defparam DLX_IDinst_RegFile_18_26_564.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_18_26_564 (
    .I(DLX_IDinst_WB_data_eff[26]),
    .CE(DLX_IDinst__n0586),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_18_26)
  );
  X_ZERO \DLX_IDinst_RegFile_4_8/LOGIC_ZERO_565  (
    .O(\DLX_IDinst_RegFile_4_8/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_130_566 (
    .IA(\DLX_IDinst_RegFile_4_8/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_4_8/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_189),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_130)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1891.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1891 (
    .ADR0(DLX_IDinst_RegFile_4_8),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_45),
    .ADR2(DLX_IDinst_RegFile_5_8),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_189)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1901.INIT = 16'hAFCF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1901 (
    .ADR0(DLX_IDinst_RegFile_7_8),
    .ADR1(DLX_IDinst_RegFile_6_8),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_46),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_190)
  );
  X_BUF \DLX_IDinst_RegFile_4_8/COUTUSED  (
    .I(\DLX_IDinst_RegFile_4_8/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_131)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_131_567 (
    .IA(\DLX_IDinst_RegFile_4_8/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_130),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_190),
    .O(\DLX_IDinst_RegFile_4_8/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_4_8/CYINIT_568  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_129),
    .O(\DLX_IDinst_RegFile_4_8/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_5_4/LOGIC_ZERO_569  (
    .O(\DLX_IDinst_RegFile_5_4/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_578_570 (
    .IA(\DLX_IDinst_RegFile_5_4/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_5_4/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_653),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_578)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6531.INIT = 16'hBF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6531 (
    .ADR0(DLX_IDinst_RegFile_5_4),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_573),
    .ADR3(DLX_IDinst_RegFile_4_4),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_653)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6541.INIT = 16'hDFD5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6541 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_574),
    .ADR1(DLX_IDinst_RegFile_7_4),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR3(DLX_IDinst_RegFile_6_4),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_654)
  );
  X_BUF \DLX_IDinst_RegFile_5_4/COUTUSED  (
    .I(\DLX_IDinst_RegFile_5_4/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_579)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_579_571 (
    .IA(\DLX_IDinst_RegFile_5_4/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_578),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_654),
    .O(\DLX_IDinst_RegFile_5_4/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_5_4/CYINIT_572  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_577),
    .O(\DLX_IDinst_RegFile_5_4/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_4_9/LOGIC_ZERO_573  (
    .O(\DLX_IDinst_RegFile_4_9/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_146_574 (
    .IA(\DLX_IDinst_RegFile_4_9/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_4_9/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_205),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_146)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2051.INIT = 16'hFD5D;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2051 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_45),
    .ADR1(DLX_IDinst_RegFile_4_9),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR3(DLX_IDinst_RegFile_5_9),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_205)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2061.INIT = 16'hCFAF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2061 (
    .ADR0(DLX_IDinst_RegFile_6_9),
    .ADR1(DLX_IDinst_RegFile_7_9),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_46),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_206)
  );
  X_BUF \DLX_IDinst_RegFile_4_9/COUTUSED  (
    .I(\DLX_IDinst_RegFile_4_9/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_147)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_147_575 (
    .IA(\DLX_IDinst_RegFile_4_9/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_146),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_206),
    .O(\DLX_IDinst_RegFile_4_9/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_4_9/CYINIT_576  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_145),
    .O(\DLX_IDinst_RegFile_4_9/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_5_5/LOGIC_ZERO_577  (
    .O(\DLX_IDinst_RegFile_5_5/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_594_578 (
    .IA(\DLX_IDinst_RegFile_5_5/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_5_5/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_669),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_594)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6691.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6691 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR1(DLX_IDinst_RegFile_4_5),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_573),
    .ADR3(DLX_IDinst_RegFile_5_5),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_669)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6701.INIT = 16'hACFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6701 (
    .ADR0(DLX_IDinst_RegFile_7_5),
    .ADR1(DLX_IDinst_RegFile_6_5),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_574),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_670)
  );
  X_BUF \DLX_IDinst_RegFile_5_5/COUTUSED  (
    .I(\DLX_IDinst_RegFile_5_5/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_595)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_595_579 (
    .IA(\DLX_IDinst_RegFile_5_5/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_594),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_670),
    .O(\DLX_IDinst_RegFile_5_5/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_5_5/CYINIT_580  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_593),
    .O(\DLX_IDinst_RegFile_5_5/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_5_6/LOGIC_ZERO_581  (
    .O(\DLX_IDinst_RegFile_5_6/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_610_582 (
    .IA(\DLX_IDinst_RegFile_5_6/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_5_6/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_685),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_610)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6851.INIT = 16'hBF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6851 (
    .ADR0(DLX_IDinst_RegFile_5_6),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_573),
    .ADR3(DLX_IDinst_RegFile_4_6),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_685)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6861.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6861 (
    .ADR0(DLX_IDinst_RegFile_6_6),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_574),
    .ADR3(DLX_IDinst_RegFile_7_6),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_686)
  );
  X_BUF \DLX_IDinst_RegFile_5_6/COUTUSED  (
    .I(\DLX_IDinst_RegFile_5_6/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_611)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_611_583 (
    .IA(\DLX_IDinst_RegFile_5_6/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_610),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_686),
    .O(\DLX_IDinst_RegFile_5_6/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_5_6/CYINIT_584  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_609),
    .O(\DLX_IDinst_RegFile_5_6/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_5_7/LOGIC_ZERO_585  (
    .O(\DLX_IDinst_RegFile_5_7/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_626_586 (
    .IA(\DLX_IDinst_RegFile_5_7/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_5_7/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_701),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_626)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7011.INIT = 16'hF5DD;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7011 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_573),
    .ADR1(DLX_IDinst_RegFile_4_7),
    .ADR2(DLX_IDinst_RegFile_5_7),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_701)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7021.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7021 (
    .ADR0(DLX_IDinst_RegFile_6_7),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_574),
    .ADR3(DLX_IDinst_RegFile_7_7),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_702)
  );
  X_BUF \DLX_IDinst_RegFile_5_7/COUTUSED  (
    .I(\DLX_IDinst_RegFile_5_7/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_627)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_627_587 (
    .IA(\DLX_IDinst_RegFile_5_7/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_626),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_702),
    .O(\DLX_IDinst_RegFile_5_7/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_5_7/CYINIT_588  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_625),
    .O(\DLX_IDinst_RegFile_5_7/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_5_8/LOGIC_ZERO_589  (
    .O(\DLX_IDinst_RegFile_5_8/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_642_590 (
    .IA(\DLX_IDinst_RegFile_5_8/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_5_8/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_717),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_642)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7171.INIT = 16'hFB73;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7171 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_573),
    .ADR2(DLX_IDinst_RegFile_4_8),
    .ADR3(DLX_IDinst_RegFile_5_8),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_717)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7181.INIT = 16'hF5DD;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7181 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_574),
    .ADR1(DLX_IDinst_RegFile_6_8),
    .ADR2(DLX_IDinst_RegFile_7_8),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_718)
  );
  X_BUF \DLX_IDinst_RegFile_5_8/COUTUSED  (
    .I(\DLX_IDinst_RegFile_5_8/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_643)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_643_591 (
    .IA(\DLX_IDinst_RegFile_5_8/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_642),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_718),
    .O(\DLX_IDinst_RegFile_5_8/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_5_8/CYINIT_592  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_641),
    .O(\DLX_IDinst_RegFile_5_8/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_5_9/LOGIC_ZERO_593  (
    .O(\DLX_IDinst_RegFile_5_9/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_658_594 (
    .IA(\DLX_IDinst_RegFile_5_9/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_5_9/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_733),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_658)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7331.INIT = 16'hE2FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7331 (
    .ADR0(DLX_IDinst_RegFile_4_9),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR2(DLX_IDinst_RegFile_5_9),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_573),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_733)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7341.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7341 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_574),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR2(DLX_IDinst_RegFile_6_9),
    .ADR3(DLX_IDinst_RegFile_7_9),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_734)
  );
  X_BUF \DLX_IDinst_RegFile_5_9/COUTUSED  (
    .I(\DLX_IDinst_RegFile_5_9/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_659)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_659_595 (
    .IA(\DLX_IDinst_RegFile_5_9/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_658),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_734),
    .O(\DLX_IDinst_RegFile_5_9/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_5_9/CYINIT_596  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_657),
    .O(\DLX_IDinst_RegFile_5_9/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_8_0/LOGIC_ZERO_597  (
    .O(\DLX_IDinst_RegFile_8_0/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_4_598 (
    .IA(\DLX_IDinst_RegFile_8_0/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_8_0/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_63),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_4)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_631.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_631 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_47),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR2(DLX_IDinst_RegFile_8_0),
    .ADR3(DLX_IDinst_RegFile_9_0),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_63)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_641.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_641 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR1(DLX_IDinst_RegFile_10_0),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_48),
    .ADR3(DLX_IDinst_RegFile_11_0),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_64)
  );
  X_BUF \DLX_IDinst_RegFile_8_0/COUTUSED  (
    .I(\DLX_IDinst_RegFile_8_0/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_5)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_5_599 (
    .IA(\DLX_IDinst_RegFile_8_0/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_4),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_64),
    .O(\DLX_IDinst_RegFile_8_0/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_8_0/CYINIT_600  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_3),
    .O(\DLX_IDinst_RegFile_8_0/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_8_1/LOGIC_ZERO_601  (
    .O(\DLX_IDinst_RegFile_8_1/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_20_602 (
    .IA(\DLX_IDinst_RegFile_8_1/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_8_1/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_79),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_20)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_791.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_791 (
    .ADR0(DLX_IDinst_RegFile_8_1),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_47),
    .ADR3(DLX_IDinst_RegFile_9_1),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_79)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_801.INIT = 16'hDDF5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_801 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_48),
    .ADR1(DLX_IDinst_RegFile_11_1),
    .ADR2(DLX_IDinst_RegFile_10_1),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_80)
  );
  X_BUF \DLX_IDinst_RegFile_8_1/COUTUSED  (
    .I(\DLX_IDinst_RegFile_8_1/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_21)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_21_603 (
    .IA(\DLX_IDinst_RegFile_8_1/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_20),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_80),
    .O(\DLX_IDinst_RegFile_8_1/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_8_1/CYINIT_604  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_19),
    .O(\DLX_IDinst_RegFile_8_1/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_8_2/LOGIC_ZERO_605  (
    .O(\DLX_IDinst_RegFile_8_2/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_36_606 (
    .IA(\DLX_IDinst_RegFile_8_2/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_8_2/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_95),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_36)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_951.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_951 (
    .ADR0(DLX_IDinst_RegFile_9_2),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_47),
    .ADR2(DLX_IDinst_RegFile_8_2),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_95)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_961.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_961 (
    .ADR0(DLX_IDinst_RegFile_11_2),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_48),
    .ADR2(DLX_IDinst_RegFile_10_2),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_96)
  );
  X_BUF \DLX_IDinst_RegFile_8_2/COUTUSED  (
    .I(\DLX_IDinst_RegFile_8_2/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_37)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_37_607 (
    .IA(\DLX_IDinst_RegFile_8_2/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_36),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_96),
    .O(\DLX_IDinst_RegFile_8_2/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_8_2/CYINIT_608  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_35),
    .O(\DLX_IDinst_RegFile_8_2/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_8_3/LOGIC_ZERO_609  (
    .O(\DLX_IDinst_RegFile_8_3/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_52_610 (
    .IA(\DLX_IDinst_RegFile_8_3/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_8_3/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_111),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_52)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1111.INIT = 16'hFB3B;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1111 (
    .ADR0(DLX_IDinst_RegFile_8_3),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_47),
    .ADR2(DLX_IDinst_jtarget[16]),
    .ADR3(DLX_IDinst_RegFile_9_3),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_111)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1121.INIT = 16'hF5DD;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1121 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_48),
    .ADR1(DLX_IDinst_RegFile_10_3),
    .ADR2(DLX_IDinst_RegFile_11_3),
    .ADR3(DLX_IDinst_jtarget[16]),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_112)
  );
  X_BUF \DLX_IDinst_RegFile_8_3/COUTUSED  (
    .I(\DLX_IDinst_RegFile_8_3/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_53)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_53_611 (
    .IA(\DLX_IDinst_RegFile_8_3/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_52),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_112),
    .O(\DLX_IDinst_RegFile_8_3/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_8_3/CYINIT_612  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_51),
    .O(\DLX_IDinst_RegFile_8_3/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_8_4/LOGIC_ZERO_613  (
    .O(\DLX_IDinst_RegFile_8_4/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_68_614 (
    .IA(\DLX_IDinst_RegFile_8_4/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_8_4/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_127),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_68)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1271.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1271 (
    .ADR0(DLX_IDinst_RegFile_8_4),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_47),
    .ADR2(DLX_IDinst_RegFile_9_4),
    .ADR3(DLX_IDinst_jtarget[16]),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_127)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1281.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1281 (
    .ADR0(DLX_IDinst_RegFile_10_4),
    .ADR1(DLX_IDinst_jtarget[16]),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_48),
    .ADR3(DLX_IDinst_RegFile_11_4),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_128)
  );
  X_BUF \DLX_IDinst_RegFile_8_4/COUTUSED  (
    .I(\DLX_IDinst_RegFile_8_4/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_69)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_69_615 (
    .IA(\DLX_IDinst_RegFile_8_4/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_68),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_128),
    .O(\DLX_IDinst_RegFile_8_4/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_8_4/CYINIT_616  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_67),
    .O(\DLX_IDinst_RegFile_8_4/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_9_0/LOGIC_ZERO_617  (
    .O(\DLX_IDinst_RegFile_9_0/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_516_618 (
    .IA(\DLX_IDinst_RegFile_9_0/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_9_0/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_591),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_516)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_5911.INIT = 16'hE4FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_5911 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR1(DLX_IDinst_RegFile_8_0),
    .ADR2(DLX_IDinst_RegFile_9_0),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_575),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_591)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_5921.INIT = 16'hBF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_5921 (
    .ADR0(DLX_IDinst_RegFile_11_0),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_576),
    .ADR3(DLX_IDinst_RegFile_10_0),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_592)
  );
  X_BUF \DLX_IDinst_RegFile_9_0/COUTUSED  (
    .I(\DLX_IDinst_RegFile_9_0/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_517)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_517_619 (
    .IA(\DLX_IDinst_RegFile_9_0/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_516),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_592),
    .O(\DLX_IDinst_RegFile_9_0/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_9_0/CYINIT_620  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_515),
    .O(\DLX_IDinst_RegFile_9_0/CYINIT )
  );
  defparam DLX_IDinst_RegFile_19_10_621.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_19_10_621 (
    .I(DLX_IDinst_WB_data_eff[10]),
    .CE(DLX_IDinst__n0588),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_19_10)
  );
  X_ZERO \DLX_IDinst_RegFile_8_5/LOGIC_ZERO_622  (
    .O(\DLX_IDinst_RegFile_8_5/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_84_623 (
    .IA(\DLX_IDinst_RegFile_8_5/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_8_5/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_143),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_84)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1431.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1431 (
    .ADR0(DLX_IDinst_RegFile_8_5),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_47),
    .ADR2(DLX_IDinst_RegFile_9_5),
    .ADR3(DLX_IDinst_jtarget[16]),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_143)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1441.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1441 (
    .ADR0(DLX_IDinst_RegFile_10_5),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_48),
    .ADR2(DLX_IDinst_RegFile_11_5),
    .ADR3(DLX_IDinst_jtarget[16]),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_144)
  );
  X_BUF \DLX_IDinst_RegFile_8_5/COUTUSED  (
    .I(\DLX_IDinst_RegFile_8_5/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_85)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_85_624 (
    .IA(\DLX_IDinst_RegFile_8_5/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_84),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_144),
    .O(\DLX_IDinst_RegFile_8_5/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_8_5/CYINIT_625  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_83),
    .O(\DLX_IDinst_RegFile_8_5/CYINIT )
  );
  defparam DLX_IDinst_RegFile_26_26_626.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_26_26_626 (
    .I(DLX_IDinst_WB_data_eff[26]),
    .CE(DLX_IDinst__n0602),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_26_26)
  );
  X_ZERO \DLX_IDinst_RegFile_9_1/LOGIC_ZERO_627  (
    .O(\DLX_IDinst_RegFile_9_1/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_532_628 (
    .IA(\DLX_IDinst_RegFile_9_1/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_9_1/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_607),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_532)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6071.INIT = 16'hDF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6071 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR1(DLX_IDinst_RegFile_9_1),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_575),
    .ADR3(DLX_IDinst_RegFile_8_1),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_607)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6081.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6081 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR1(DLX_IDinst_RegFile_10_1),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_576),
    .ADR3(DLX_IDinst_RegFile_11_1),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_608)
  );
  X_BUF \DLX_IDinst_RegFile_9_1/COUTUSED  (
    .I(\DLX_IDinst_RegFile_9_1/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_533)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_533_629 (
    .IA(\DLX_IDinst_RegFile_9_1/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_532),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_608),
    .O(\DLX_IDinst_RegFile_9_1/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_9_1/CYINIT_630  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_531),
    .O(\DLX_IDinst_RegFile_9_1/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_8_6/LOGIC_ZERO_631  (
    .O(\DLX_IDinst_RegFile_8_6/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_100_632 (
    .IA(\DLX_IDinst_RegFile_8_6/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_8_6/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_159),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_100)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1591.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1591 (
    .ADR0(DLX_IDinst_RegFile_8_6),
    .ADR1(DLX_IDinst_jtarget[16]),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_47),
    .ADR3(DLX_IDinst_RegFile_9_6),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_159)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1601.INIT = 16'hBF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1601 (
    .ADR0(DLX_IDinst_RegFile_11_6),
    .ADR1(DLX_IDinst_jtarget[16]),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_48),
    .ADR3(DLX_IDinst_RegFile_10_6),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_160)
  );
  X_BUF \DLX_IDinst_RegFile_8_6/COUTUSED  (
    .I(\DLX_IDinst_RegFile_8_6/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_101)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_101_633 (
    .IA(\DLX_IDinst_RegFile_8_6/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_100),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_160),
    .O(\DLX_IDinst_RegFile_8_6/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_8_6/CYINIT_634  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_99),
    .O(\DLX_IDinst_RegFile_8_6/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_9_2/LOGIC_ZERO_635  (
    .O(\DLX_IDinst_RegFile_9_2/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_548_636 (
    .IA(\DLX_IDinst_RegFile_9_2/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_9_2/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_623),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_548)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6231.INIT = 16'hDF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6231 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR1(DLX_IDinst_RegFile_9_2),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_575),
    .ADR3(DLX_IDinst_RegFile_8_2),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_623)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6241.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6241 (
    .ADR0(DLX_IDinst_RegFile_10_2),
    .ADR1(DLX_IDinst_RegFile_11_2),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_576),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_624)
  );
  X_BUF \DLX_IDinst_RegFile_9_2/COUTUSED  (
    .I(\DLX_IDinst_RegFile_9_2/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_549)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_549_637 (
    .IA(\DLX_IDinst_RegFile_9_2/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_548),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_624),
    .O(\DLX_IDinst_RegFile_9_2/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_9_2/CYINIT_638  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_547),
    .O(\DLX_IDinst_RegFile_9_2/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_8_7/LOGIC_ZERO_639  (
    .O(\DLX_IDinst_RegFile_8_7/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_116_640 (
    .IA(\DLX_IDinst_RegFile_8_7/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_8_7/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_175),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_116)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1751.INIT = 16'hE4FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1751 (
    .ADR0(DLX_IDinst_jtarget[16]),
    .ADR1(DLX_IDinst_RegFile_8_7),
    .ADR2(DLX_IDinst_RegFile_9_7),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_47),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_175)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1761.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1761 (
    .ADR0(DLX_IDinst_RegFile_10_7),
    .ADR1(DLX_IDinst_jtarget[16]),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_48),
    .ADR3(DLX_IDinst_RegFile_11_7),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_176)
  );
  X_BUF \DLX_IDinst_RegFile_8_7/COUTUSED  (
    .I(\DLX_IDinst_RegFile_8_7/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_117)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_117_641 (
    .IA(\DLX_IDinst_RegFile_8_7/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_116),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_176),
    .O(\DLX_IDinst_RegFile_8_7/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_8_7/CYINIT_642  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_115),
    .O(\DLX_IDinst_RegFile_8_7/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_9_3/LOGIC_ZERO_643  (
    .O(\DLX_IDinst_RegFile_9_3/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_564_644 (
    .IA(\DLX_IDinst_RegFile_9_3/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_9_3/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_639),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_564)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6391.INIT = 16'hDFD5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6391 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_575),
    .ADR1(DLX_IDinst_RegFile_9_3),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR3(DLX_IDinst_RegFile_8_3),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_639)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6401.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6401 (
    .ADR0(DLX_IDinst_RegFile_10_3),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_576),
    .ADR2(DLX_IDinst_RegFile_11_3),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_640)
  );
  X_BUF \DLX_IDinst_RegFile_9_3/COUTUSED  (
    .I(\DLX_IDinst_RegFile_9_3/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_565)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_565_645 (
    .IA(\DLX_IDinst_RegFile_9_3/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_564),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_640),
    .O(\DLX_IDinst_RegFile_9_3/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_9_3/CYINIT_646  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_563),
    .O(\DLX_IDinst_RegFile_9_3/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_8_8/LOGIC_ZERO_647  (
    .O(\DLX_IDinst_RegFile_8_8/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_132_648 (
    .IA(\DLX_IDinst_RegFile_8_8/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_8_8/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_191),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_132)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1911.INIT = 16'hE2FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1911 (
    .ADR0(DLX_IDinst_RegFile_8_8),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR2(DLX_IDinst_RegFile_9_8),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_47),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_191)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1921.INIT = 16'hDFD5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1921 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_48),
    .ADR1(DLX_IDinst_RegFile_11_8),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR3(DLX_IDinst_RegFile_10_8),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_192)
  );
  X_BUF \DLX_IDinst_RegFile_8_8/COUTUSED  (
    .I(\DLX_IDinst_RegFile_8_8/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_133)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_133_649 (
    .IA(\DLX_IDinst_RegFile_8_8/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_132),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_192),
    .O(\DLX_IDinst_RegFile_8_8/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_8_8/CYINIT_650  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_131),
    .O(\DLX_IDinst_RegFile_8_8/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_9_4/LOGIC_ZERO_651  (
    .O(\DLX_IDinst_RegFile_9_4/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_580_652 (
    .IA(\DLX_IDinst_RegFile_9_4/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_9_4/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_655),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_580)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6551.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6551 (
    .ADR0(DLX_IDinst_RegFile_8_4),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_575),
    .ADR3(DLX_IDinst_RegFile_9_4),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_655)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6561.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6561 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_576),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR2(DLX_IDinst_RegFile_10_4),
    .ADR3(DLX_IDinst_RegFile_11_4),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_656)
  );
  X_BUF \DLX_IDinst_RegFile_9_4/COUTUSED  (
    .I(\DLX_IDinst_RegFile_9_4/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_581)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_581_653 (
    .IA(\DLX_IDinst_RegFile_9_4/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_580),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_656),
    .O(\DLX_IDinst_RegFile_9_4/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_9_4/CYINIT_654  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_579),
    .O(\DLX_IDinst_RegFile_9_4/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_8_9/LOGIC_ZERO_655  (
    .O(\DLX_IDinst_RegFile_8_9/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_148_656 (
    .IA(\DLX_IDinst_RegFile_8_9/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_8_9/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_207),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_148)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2071.INIT = 16'hBFB3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2071 (
    .ADR0(DLX_IDinst_RegFile_9_9),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_47),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR3(DLX_IDinst_RegFile_8_9),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_207)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2081.INIT = 16'hACFF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2081 (
    .ADR0(DLX_IDinst_RegFile_11_9),
    .ADR1(DLX_IDinst_RegFile_10_9),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_48),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_208)
  );
  X_BUF \DLX_IDinst_RegFile_8_9/COUTUSED  (
    .I(\DLX_IDinst_RegFile_8_9/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_149)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_149_657 (
    .IA(\DLX_IDinst_RegFile_8_9/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_148),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_208),
    .O(\DLX_IDinst_RegFile_8_9/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_8_9/CYINIT_658  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_147),
    .O(\DLX_IDinst_RegFile_8_9/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_9_5/LOGIC_ZERO_659  (
    .O(\DLX_IDinst_RegFile_9_5/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_596_660 (
    .IA(\DLX_IDinst_RegFile_9_5/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_9_5/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_671),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_596)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6711.INIT = 16'hFB3B;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6711 (
    .ADR0(DLX_IDinst_RegFile_8_5),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_575),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR3(DLX_IDinst_RegFile_9_5),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_671)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6721.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6721 (
    .ADR0(DLX_IDinst_RegFile_10_5),
    .ADR1(DLX_IDinst_RegFile_11_5),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_576),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_672)
  );
  X_BUF \DLX_IDinst_RegFile_9_5/COUTUSED  (
    .I(\DLX_IDinst_RegFile_9_5/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_597)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_597_661 (
    .IA(\DLX_IDinst_RegFile_9_5/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_596),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_672),
    .O(\DLX_IDinst_RegFile_9_5/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_9_5/CYINIT_662  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_595),
    .O(\DLX_IDinst_RegFile_9_5/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_9_6/LOGIC_ZERO_663  (
    .O(\DLX_IDinst_RegFile_9_6/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_612_664 (
    .IA(\DLX_IDinst_RegFile_9_6/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_9_6/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_687),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_612)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6871.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6871 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_575),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR2(DLX_IDinst_RegFile_8_6),
    .ADR3(DLX_IDinst_RegFile_9_6),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_687)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6881.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6881 (
    .ADR0(DLX_IDinst_RegFile_10_6),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_576),
    .ADR3(DLX_IDinst_RegFile_11_6),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_688)
  );
  X_BUF \DLX_IDinst_RegFile_9_6/COUTUSED  (
    .I(\DLX_IDinst_RegFile_9_6/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_613)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_613_665 (
    .IA(\DLX_IDinst_RegFile_9_6/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_612),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_688),
    .O(\DLX_IDinst_RegFile_9_6/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_9_6/CYINIT_666  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_611),
    .O(\DLX_IDinst_RegFile_9_6/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_9_7/LOGIC_ZERO_667  (
    .O(\DLX_IDinst_RegFile_9_7/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_628_668 (
    .IA(\DLX_IDinst_RegFile_9_7/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_9_7/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_703),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_628)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7031.INIT = 16'hDFD5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7031 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_575),
    .ADR1(DLX_IDinst_RegFile_9_7),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR3(DLX_IDinst_RegFile_8_7),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_703)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7041.INIT = 16'hCFAF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7041 (
    .ADR0(DLX_IDinst_RegFile_10_7),
    .ADR1(DLX_IDinst_RegFile_11_7),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_576),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_704)
  );
  X_BUF \DLX_IDinst_RegFile_9_7/COUTUSED  (
    .I(\DLX_IDinst_RegFile_9_7/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_629)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_629_669 (
    .IA(\DLX_IDinst_RegFile_9_7/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_628),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_704),
    .O(\DLX_IDinst_RegFile_9_7/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_9_7/CYINIT_670  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_627),
    .O(\DLX_IDinst_RegFile_9_7/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_9_8/LOGIC_ZERO_671  (
    .O(\DLX_IDinst_RegFile_9_8/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_644_672 (
    .IA(\DLX_IDinst_RegFile_9_8/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_9_8/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_719),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_644)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7191.INIT = 16'hDF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7191 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR1(DLX_IDinst_RegFile_9_8),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_575),
    .ADR3(DLX_IDinst_RegFile_8_8),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_719)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7201.INIT = 16'hFB73;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7201 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_576),
    .ADR2(DLX_IDinst_RegFile_10_8),
    .ADR3(DLX_IDinst_RegFile_11_8),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_720)
  );
  X_BUF \DLX_IDinst_RegFile_9_8/COUTUSED  (
    .I(\DLX_IDinst_RegFile_9_8/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_645)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_645_673 (
    .IA(\DLX_IDinst_RegFile_9_8/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_644),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_720),
    .O(\DLX_IDinst_RegFile_9_8/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_9_8/CYINIT_674  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_643),
    .O(\DLX_IDinst_RegFile_9_8/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_9_9/LOGIC_ZERO_675  (
    .O(\DLX_IDinst_RegFile_9_9/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_660_676 (
    .IA(\DLX_IDinst_RegFile_9_9/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_9_9/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_735),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_660)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7351.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7351 (
    .ADR0(DLX_IDinst_RegFile_8_9),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_575),
    .ADR3(DLX_IDinst_RegFile_9_9),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_735)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7361.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7361 (
    .ADR0(DLX_IDinst_RegFile_11_9),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_576),
    .ADR2(DLX_IDinst_RegFile_10_9),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_736)
  );
  X_BUF \DLX_IDinst_RegFile_9_9/COUTUSED  (
    .I(\DLX_IDinst_RegFile_9_9/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_661)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_661_677 (
    .IA(\DLX_IDinst_RegFile_9_9/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_660),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_736),
    .O(\DLX_IDinst_RegFile_9_9/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_9_9/CYINIT_678  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_659),
    .O(\DLX_IDinst_RegFile_9_9/CYINIT )
  );
  defparam \DLX_IFinst__n0001<1>_SW0 .INIT = 16'h03F3;
  X_LUT4 \DLX_IFinst__n0001<1>_SW0  (
    .ADR0(VCC),
    .ADR1(DLX_IFinst_NPC[1]),
    .ADR2(DLX_IFinst__n0000),
    .ADR3(DLX_IFinst_PC[1]),
    .O(\DLX_IFinst_NPC<1>/FROM )
  );
  defparam \DLX_IFinst__n0001<1> .INIT = 16'hA0F5;
  X_LUT4 \DLX_IFinst__n0001<1>  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_branch_address[1]),
    .ADR3(N129899),
    .O(\DLX_IFinst_NPC<1>/GROM )
  );
  X_BUF \DLX_IFinst_NPC<1>/XUSED  (
    .I(\DLX_IFinst_NPC<1>/FROM ),
    .O(N129899)
  );
  X_BUF \DLX_IFinst_NPC<1>/YUSED  (
    .I(\DLX_IFinst_NPC<1>/GROM ),
    .O(DLX_IFinst__n0001[1])
  );
  defparam \DLX_IFinst__n0001<2>_SW0 .INIT = 16'h7272;
  X_LUT4 \DLX_IFinst__n0001<2>_SW0  (
    .ADR0(DLX_IFinst__n0000),
    .ADR1(DLX_IFinst_PC[2]),
    .ADR2(DLX_IFinst_NPC[2]),
    .ADR3(VCC),
    .O(\DLX_IFinst_NPC<2>/FROM )
  );
  defparam \DLX_IFinst__n0001<2> .INIT = 16'hA0F5;
  X_LUT4 \DLX_IFinst__n0001<2>  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_branch_address[2]),
    .ADR3(N129847),
    .O(\DLX_IFinst_NPC<2>/GROM )
  );
  X_BUF \DLX_IFinst_NPC<2>/XUSED  (
    .I(\DLX_IFinst_NPC<2>/FROM ),
    .O(N129847)
  );
  X_BUF \DLX_IFinst_NPC<2>/YUSED  (
    .I(\DLX_IFinst_NPC<2>/GROM ),
    .O(DLX_IFinst__n0001[2])
  );
  defparam \mask<2>_SW122_SW0 .INIT = 16'hD8AA;
  X_LUT4 \mask<2>_SW122_SW0  (
    .ADR0(DLX_EXinst_byte),
    .ADR1(DLX_EXinst_ALU_result[1]),
    .ADR2(DLX_EXinst_word),
    .ADR3(DLX_EXinst_ALU_result[0]),
    .O(\N164184/FROM )
  );
  defparam \mask<2>_SW122 .INIT = 16'h0001;
  X_LUT4 \mask<2>_SW122  (
    .ADR0(DLX_EXinst_ALU_result[12]),
    .ADR1(DLX_EXinst_ALU_result[14]),
    .ADR2(DLX_EXinst_ALU_result[13]),
    .ADR3(N164184),
    .O(\N164184/GROM )
  );
  X_BUF \N164184/XUSED  (
    .I(\N164184/FROM ),
    .O(N164184)
  );
  X_BUF \N164184/YUSED  (
    .I(\N164184/GROM ),
    .O(mask_2_OBUF)
  );
  defparam \DLX_IFinst__n0001<3>_SW0 .INIT = 16'h4477;
  X_LUT4 \DLX_IFinst__n0001<3>_SW0  (
    .ADR0(DLX_IFinst_PC[3]),
    .ADR1(DLX_IFinst__n0000),
    .ADR2(VCC),
    .ADR3(DLX_IFinst__n0015[3]),
    .O(\DLX_IFinst_NPC<3>/FROM )
  );
  defparam \DLX_IFinst__n0001<3> .INIT = 16'hA0F5;
  X_LUT4 \DLX_IFinst__n0001<3>  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_branch_address[3]),
    .ADR3(N129795),
    .O(\DLX_IFinst_NPC<3>/GROM )
  );
  X_BUF \DLX_IFinst_NPC<3>/XUSED  (
    .I(\DLX_IFinst_NPC<3>/FROM ),
    .O(N129795)
  );
  X_BUF \DLX_IFinst_NPC<3>/YUSED  (
    .I(\DLX_IFinst_NPC<3>/GROM ),
    .O(DLX_IFinst__n0001[3])
  );
  defparam \DLX_IFinst__n0001<4>_SW0 .INIT = 16'h2277;
  X_LUT4 \DLX_IFinst__n0001<4>_SW0  (
    .ADR0(DLX_IFinst__n0000),
    .ADR1(DLX_IFinst_PC[4]),
    .ADR2(VCC),
    .ADR3(DLX_IFinst__n0015[4]),
    .O(\DLX_IFinst_NPC<4>/FROM )
  );
  defparam \DLX_IFinst__n0001<4> .INIT = 16'h88BB;
  X_LUT4 \DLX_IFinst__n0001<4>  (
    .ADR0(DLX_IDinst_branch_address[4]),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(VCC),
    .ADR3(N129743),
    .O(\DLX_IFinst_NPC<4>/GROM )
  );
  X_BUF \DLX_IFinst_NPC<4>/XUSED  (
    .I(\DLX_IFinst_NPC<4>/FROM ),
    .O(N129743)
  );
  X_BUF \DLX_IFinst_NPC<4>/YUSED  (
    .I(\DLX_IFinst_NPC<4>/GROM ),
    .O(DLX_IFinst__n0001[4])
  );
  defparam \DLX_IFinst__n0001<5>_SW0 .INIT = 16'h4477;
  X_LUT4 \DLX_IFinst__n0001<5>_SW0  (
    .ADR0(DLX_IFinst_PC[5]),
    .ADR1(DLX_IFinst__n0000),
    .ADR2(VCC),
    .ADR3(DLX_IFinst__n0015[5]),
    .O(\DLX_IFinst_NPC<5>/FROM )
  );
  defparam \DLX_IFinst__n0001<5> .INIT = 16'hA0AF;
  X_LUT4 \DLX_IFinst__n0001<5>  (
    .ADR0(DLX_IDinst_branch_address[5]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(N129691),
    .O(\DLX_IFinst_NPC<5>/GROM )
  );
  X_BUF \DLX_IFinst_NPC<5>/XUSED  (
    .I(\DLX_IFinst_NPC<5>/FROM ),
    .O(N129691)
  );
  X_BUF \DLX_IFinst_NPC<5>/YUSED  (
    .I(\DLX_IFinst_NPC<5>/GROM ),
    .O(DLX_IFinst__n0001[5])
  );
  defparam \DLX_IFinst__n0001<6>_SW0 .INIT = 16'h2277;
  X_LUT4 \DLX_IFinst__n0001<6>_SW0  (
    .ADR0(DLX_IFinst__n0000),
    .ADR1(DLX_IFinst_PC[6]),
    .ADR2(VCC),
    .ADR3(DLX_IFinst__n0015[6]),
    .O(\DLX_IFinst_NPC<6>/FROM )
  );
  defparam \DLX_IFinst__n0001<6> .INIT = 16'hC0CF;
  X_LUT4 \DLX_IFinst__n0001<6>  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_branch_address[6]),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(N129639),
    .O(\DLX_IFinst_NPC<6>/GROM )
  );
  X_BUF \DLX_IFinst_NPC<6>/XUSED  (
    .I(\DLX_IFinst_NPC<6>/FROM ),
    .O(N129639)
  );
  X_BUF \DLX_IFinst_NPC<6>/YUSED  (
    .I(\DLX_IFinst_NPC<6>/GROM ),
    .O(DLX_IFinst__n0001[6])
  );
  defparam \DLX_IFinst__n0001<7>_SW0 .INIT = 16'h3355;
  X_LUT4 \DLX_IFinst__n0001<7>_SW0  (
    .ADR0(DLX_IFinst__n0015[7]),
    .ADR1(DLX_IFinst_PC[7]),
    .ADR2(VCC),
    .ADR3(DLX_IFinst__n0000),
    .O(\DLX_IFinst_NPC<7>/FROM )
  );
  defparam \DLX_IFinst__n0001<7> .INIT = 16'hC0CF;
  X_LUT4 \DLX_IFinst__n0001<7>  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_branch_address[7]),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(N129587),
    .O(\DLX_IFinst_NPC<7>/GROM )
  );
  X_BUF \DLX_IFinst_NPC<7>/XUSED  (
    .I(\DLX_IFinst_NPC<7>/FROM ),
    .O(N129587)
  );
  X_BUF \DLX_IFinst_NPC<7>/YUSED  (
    .I(\DLX_IFinst_NPC<7>/GROM ),
    .O(DLX_IFinst__n0001[7])
  );
  defparam \DLX_IFinst__n0001<8>_SW0 .INIT = 16'h550F;
  X_LUT4 \DLX_IFinst__n0001<8>_SW0  (
    .ADR0(DLX_IFinst_PC[8]),
    .ADR1(VCC),
    .ADR2(DLX_IFinst__n0015[8]),
    .ADR3(DLX_IFinst__n0000),
    .O(\DLX_IFinst_NPC<8>/FROM )
  );
  defparam \DLX_IFinst__n0001<8> .INIT = 16'hA0F5;
  X_LUT4 \DLX_IFinst__n0001<8>  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_branch_address[8]),
    .ADR3(N129535),
    .O(\DLX_IFinst_NPC<8>/GROM )
  );
  X_BUF \DLX_IFinst_NPC<8>/XUSED  (
    .I(\DLX_IFinst_NPC<8>/FROM ),
    .O(N129535)
  );
  X_BUF \DLX_IFinst_NPC<8>/YUSED  (
    .I(\DLX_IFinst_NPC<8>/GROM ),
    .O(DLX_IFinst__n0001[8])
  );
  defparam \DLX_IFinst__n0001<9>_SW0 .INIT = 16'h4477;
  X_LUT4 \DLX_IFinst__n0001<9>_SW0  (
    .ADR0(DLX_IFinst_PC[9]),
    .ADR1(DLX_IFinst__n0000),
    .ADR2(VCC),
    .ADR3(DLX_IFinst__n0015[9]),
    .O(\DLX_IFinst_NPC<9>/FROM )
  );
  defparam \DLX_IFinst__n0001<9> .INIT = 16'hC0CF;
  X_LUT4 \DLX_IFinst__n0001<9>  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_branch_address[9]),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(N129483),
    .O(\DLX_IFinst_NPC<9>/GROM )
  );
  X_BUF \DLX_IFinst_NPC<9>/XUSED  (
    .I(\DLX_IFinst_NPC<9>/FROM ),
    .O(N129483)
  );
  X_BUF \DLX_IFinst_NPC<9>/YUSED  (
    .I(\DLX_IFinst_NPC<9>/GROM ),
    .O(DLX_IFinst__n0001[9])
  );
  defparam \DLX_EXinst__n0013<14>1 .INIT = 16'hF0AA;
  X_LUT4 \DLX_EXinst__n0013<14>1  (
    .ADR0(\DLX_IDinst_Imm[14] ),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[14]),
    .ADR3(DLX_EXinst__n0036),
    .O(\DLX_IFinst_IR_curr<7>/FROM )
  );
  defparam \DLX_EXinst__n0013<11>1 .INIT = 16'hAFA0;
  X_LUT4 \DLX_EXinst__n0013<11>1  (
    .ADR0(DLX_IDinst_reg_out_B[11]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst__n0036),
    .ADR3(\DLX_IDinst_Imm[11] ),
    .O(\DLX_IFinst_IR_curr<7>/GROM )
  );
  X_BUF \DLX_IFinst_IR_curr<7>/XUSED  (
    .I(\DLX_IFinst_IR_curr<7>/FROM ),
    .O(DLX_EXinst__n0013[14])
  );
  X_BUF \DLX_IFinst_IR_curr<7>/YUSED  (
    .I(\DLX_IFinst_IR_curr<7>/GROM ),
    .O(DLX_EXinst__n0013[11])
  );
  defparam DLX_IDinst_RegFile_11_10_679.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_11_10_679 (
    .I(DLX_IDinst_WB_data_eff[10]),
    .CE(DLX_IDinst__n0572),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_11_10)
  );
  defparam \DLX_EXinst__n0013<21>1 .INIT = 16'hEAC0;
  X_LUT4 \DLX_EXinst__n0013<21>1  (
    .ADR0(\DLX_IDinst_Imm[31] ),
    .ADR1(DLX_IDinst_reg_out_B[21]),
    .ADR2(DLX_EXinst__n0036),
    .ADR3(N136960),
    .O(\DLX_IDinst_RegFile_11_10/FROM )
  );
  defparam \DLX_EXinst__n0013<20>1 .INIT = 16'hECA0;
  X_LUT4 \DLX_EXinst__n0013<20>1  (
    .ADR0(DLX_IDinst_reg_out_B[20]),
    .ADR1(\DLX_IDinst_Imm[31] ),
    .ADR2(DLX_EXinst__n0036),
    .ADR3(N136960),
    .O(\DLX_IDinst_RegFile_11_10/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_11_10/XUSED  (
    .I(\DLX_IDinst_RegFile_11_10/FROM ),
    .O(DLX_EXinst__n0013[21])
  );
  X_BUF \DLX_IDinst_RegFile_11_10/YUSED  (
    .I(\DLX_IDinst_RegFile_11_10/GROM ),
    .O(DLX_EXinst__n0013[20])
  );
  defparam \DLX_EXinst__n0013<15>1 .INIT = 16'hD8D8;
  X_LUT4 \DLX_EXinst__n0013<15>1  (
    .ADR0(DLX_EXinst__n0036),
    .ADR1(DLX_IDinst_reg_out_B[15]),
    .ADR2(\DLX_IDinst_Imm[15] ),
    .ADR3(VCC),
    .O(\DLX_IDinst_RegFile_11_14/FROM )
  );
  defparam \DLX_EXinst__n0013<12>1 .INIT = 16'hF5A0;
  X_LUT4 \DLX_EXinst__n0013<12>1  (
    .ADR0(DLX_EXinst__n0036),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[12]),
    .ADR3(\DLX_IDinst_Imm[12] ),
    .O(\DLX_IDinst_RegFile_11_14/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_11_14/XUSED  (
    .I(\DLX_IDinst_RegFile_11_14/FROM ),
    .O(DLX_EXinst__n0013[15])
  );
  X_BUF \DLX_IDinst_RegFile_11_14/YUSED  (
    .I(\DLX_IDinst_RegFile_11_14/GROM ),
    .O(DLX_EXinst__n0013[12])
  );
  defparam \DLX_EXinst__n0013<27>1 .INIT = 16'hECA0;
  X_LUT4 \DLX_EXinst__n0013<27>1  (
    .ADR0(N136960),
    .ADR1(DLX_IDinst_reg_out_B[27]),
    .ADR2(\DLX_IDinst_Imm[31] ),
    .ADR3(DLX_EXinst__n0036),
    .O(\DLX_IDinst_RegFile_11_26/FROM )
  );
  defparam \DLX_EXinst__n0013<30>1 .INIT = 16'hEAC0;
  X_LUT4 \DLX_EXinst__n0013<30>1  (
    .ADR0(DLX_IDinst_reg_out_B[30]),
    .ADR1(N136960),
    .ADR2(\DLX_IDinst_Imm[31] ),
    .ADR3(DLX_EXinst__n0036),
    .O(\DLX_IDinst_RegFile_11_26/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_11_26/XUSED  (
    .I(\DLX_IDinst_RegFile_11_26/FROM ),
    .O(DLX_EXinst__n0013[27])
  );
  X_BUF \DLX_IDinst_RegFile_11_26/YUSED  (
    .I(\DLX_IDinst_RegFile_11_26/GROM ),
    .O(DLX_EXinst__n0013[30])
  );
  defparam \DLX_EXinst__n0013<18>1 .INIT = 16'hECA0;
  X_LUT4 \DLX_EXinst__n0013<18>1  (
    .ADR0(DLX_EXinst__n0036),
    .ADR1(N136960),
    .ADR2(DLX_IDinst_reg_out_B[18]),
    .ADR3(\DLX_IDinst_Imm[31] ),
    .O(\DLX_IDinst_RegFile_11_28/FROM )
  );
  defparam \DLX_EXinst__n0013<22>1 .INIT = 16'hECA0;
  X_LUT4 \DLX_EXinst__n0013<22>1  (
    .ADR0(DLX_IDinst_reg_out_B[22]),
    .ADR1(N136960),
    .ADR2(DLX_EXinst__n0036),
    .ADR3(\DLX_IDinst_Imm[31] ),
    .O(\DLX_IDinst_RegFile_11_28/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_11_28/XUSED  (
    .I(\DLX_IDinst_RegFile_11_28/FROM ),
    .O(DLX_EXinst__n0013[18])
  );
  X_BUF \DLX_IDinst_RegFile_11_28/YUSED  (
    .I(\DLX_IDinst_RegFile_11_28/GROM ),
    .O(DLX_EXinst__n0013[22])
  );
  defparam \DLX_EXinst__n0013<29>1 .INIT = 16'hECA0;
  X_LUT4 \DLX_EXinst__n0013<29>1  (
    .ADR0(N136960),
    .ADR1(DLX_IDinst_reg_out_B[29]),
    .ADR2(\DLX_IDinst_Imm[31] ),
    .ADR3(DLX_EXinst__n0036),
    .O(\DLX_IDinst_RegFile_7_2/FROM )
  );
  defparam \DLX_EXinst__n0013<31>1 .INIT = 16'hEAC0;
  X_LUT4 \DLX_EXinst__n0013<31>1  (
    .ADR0(DLX_IDinst_reg_out_B[31]),
    .ADR1(N136960),
    .ADR2(\DLX_IDinst_Imm[31] ),
    .ADR3(DLX_EXinst__n0036),
    .O(\DLX_IDinst_RegFile_7_2/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_7_2/XUSED  (
    .I(\DLX_IDinst_RegFile_7_2/FROM ),
    .O(DLX_EXinst__n0013[29])
  );
  X_BUF \DLX_IDinst_RegFile_7_2/YUSED  (
    .I(\DLX_IDinst_RegFile_7_2/GROM ),
    .O(DLX_EXinst__n0013[31])
  );
  defparam \DLX_EXinst__n0013<17>1 .INIT = 16'hF888;
  X_LUT4 \DLX_EXinst__n0013<17>1  (
    .ADR0(DLX_EXinst__n0036),
    .ADR1(DLX_IDinst_reg_out_B[17]),
    .ADR2(\DLX_IDinst_Imm[31] ),
    .ADR3(N136960),
    .O(\DLX_IDinst_RegFile_2_0/FROM )
  );
  defparam \DLX_EXinst__n0013<23>1 .INIT = 16'hEAC0;
  X_LUT4 \DLX_EXinst__n0013<23>1  (
    .ADR0(\DLX_IDinst_Imm[31] ),
    .ADR1(DLX_IDinst_reg_out_B[23]),
    .ADR2(DLX_EXinst__n0036),
    .ADR3(N136960),
    .O(\DLX_IDinst_RegFile_2_0/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_2_0/XUSED  (
    .I(\DLX_IDinst_RegFile_2_0/FROM ),
    .O(DLX_EXinst__n0013[17])
  );
  X_BUF \DLX_IDinst_RegFile_2_0/YUSED  (
    .I(\DLX_IDinst_RegFile_2_0/GROM ),
    .O(DLX_EXinst__n0013[23])
  );
  defparam \DLX_EXinst__n0013<25>1 .INIT = 16'hEAC0;
  X_LUT4 \DLX_EXinst__n0013<25>1  (
    .ADR0(\DLX_IDinst_Imm[31] ),
    .ADR1(DLX_IDinst_reg_out_B[25]),
    .ADR2(DLX_EXinst__n0036),
    .ADR3(N136960),
    .O(\DLX_IDinst_EPC<2>/FROM )
  );
  defparam \DLX_EXinst__n0013<24>1 .INIT = 16'hF888;
  X_LUT4 \DLX_EXinst__n0013<24>1  (
    .ADR0(DLX_IDinst_reg_out_B[24]),
    .ADR1(DLX_EXinst__n0036),
    .ADR2(N136960),
    .ADR3(\DLX_IDinst_Imm[31] ),
    .O(\DLX_IDinst_EPC<2>/GROM )
  );
  X_BUF \DLX_IDinst_EPC<2>/XUSED  (
    .I(\DLX_IDinst_EPC<2>/FROM ),
    .O(DLX_EXinst__n0013[25])
  );
  X_BUF \DLX_IDinst_EPC<2>/YUSED  (
    .I(\DLX_IDinst_EPC<2>/GROM ),
    .O(DLX_EXinst__n0013[24])
  );
  defparam \DLX_EXinst__n0013<19>1 .INIT = 16'hECA0;
  X_LUT4 \DLX_EXinst__n0013<19>1  (
    .ADR0(DLX_IDinst_reg_out_B[19]),
    .ADR1(\DLX_IDinst_Imm[31] ),
    .ADR2(DLX_EXinst__n0036),
    .ADR3(N136960),
    .O(\DLX_IDinst_EPC<3>/FROM )
  );
  defparam \DLX_EXinst__n0013<26>1 .INIT = 16'hECA0;
  X_LUT4 \DLX_EXinst__n0013<26>1  (
    .ADR0(\DLX_IDinst_Imm[31] ),
    .ADR1(DLX_IDinst_reg_out_B[26]),
    .ADR2(N136960),
    .ADR3(DLX_EXinst__n0036),
    .O(\DLX_IDinst_EPC<3>/GROM )
  );
  X_BUF \DLX_IDinst_EPC<3>/XUSED  (
    .I(\DLX_IDinst_EPC<3>/FROM ),
    .O(DLX_EXinst__n0013[19])
  );
  X_BUF \DLX_IDinst_EPC<3>/YUSED  (
    .I(\DLX_IDinst_EPC<3>/GROM ),
    .O(DLX_EXinst__n0013[26])
  );
  defparam \DLX_EXinst__n0007<23>9 .INIT = 16'hAA20;
  X_LUT4 \DLX_EXinst__n0007<23>9  (
    .ADR0(DLX_IDinst_reg_out_A[23]),
    .ADR1(\DLX_IDinst_Imm[31] ),
    .ADR2(DLX_EXinst__n0054),
    .ADR3(DLX_EXinst__n0053),
    .O(\DLX_IDinst_EPC<4>/FROM )
  );
  defparam \DLX_EXinst__n0013<28>1 .INIT = 16'hEAC0;
  X_LUT4 \DLX_EXinst__n0013<28>1  (
    .ADR0(DLX_IDinst_reg_out_B[28]),
    .ADR1(N136960),
    .ADR2(\DLX_IDinst_Imm[31] ),
    .ADR3(DLX_EXinst__n0036),
    .O(\DLX_IDinst_EPC<4>/GROM )
  );
  X_BUF \DLX_IDinst_EPC<4>/XUSED  (
    .I(\DLX_IDinst_EPC<4>/FROM ),
    .O(CHOICE3995)
  );
  X_BUF \DLX_IDinst_EPC<4>/YUSED  (
    .I(\DLX_IDinst_EPC<4>/GROM ),
    .O(DLX_EXinst__n0013[28])
  );
  defparam \DLX_EXinst__n0007<18>9 .INIT = 16'hCE00;
  X_LUT4 \DLX_EXinst__n0007<18>9  (
    .ADR0(DLX_EXinst__n0054),
    .ADR1(DLX_EXinst__n0053),
    .ADR2(\DLX_IDinst_Imm[31] ),
    .ADR3(DLX_IDinst_reg_out_A[18]),
    .O(\DLX_IDinst_EPC<5>/FROM )
  );
  defparam \DLX_EXinst__n0007<21>9 .INIT = 16'hD0C0;
  X_LUT4 \DLX_EXinst__n0007<21>9  (
    .ADR0(\DLX_IDinst_Imm[31] ),
    .ADR1(DLX_EXinst__n0053),
    .ADR2(DLX_IDinst_reg_out_A[21]),
    .ADR3(DLX_EXinst__n0054),
    .O(\DLX_IDinst_EPC<5>/GROM )
  );
  X_BUF \DLX_IDinst_EPC<5>/XUSED  (
    .I(\DLX_IDinst_EPC<5>/FROM ),
    .O(CHOICE5196)
  );
  X_BUF \DLX_IDinst_EPC<5>/YUSED  (
    .I(\DLX_IDinst_EPC<5>/GROM ),
    .O(CHOICE4125)
  );
  defparam \DLX_EXinst__n0007<30>13 .INIT = 16'hBA00;
  X_LUT4 \DLX_EXinst__n0007<30>13  (
    .ADR0(DLX_EXinst__n0053),
    .ADR1(\DLX_IDinst_Imm[31] ),
    .ADR2(DLX_EXinst__n0054),
    .ADR3(DLX_IDinst_reg_out_A[30]),
    .O(\DLX_IFinst_PC<10>/FROM )
  );
  defparam \DLX_EXinst__n0007<22>9 .INIT = 16'hA0E0;
  X_LUT4 \DLX_EXinst__n0007<22>9  (
    .ADR0(DLX_EXinst__n0053),
    .ADR1(DLX_EXinst__n0054),
    .ADR2(DLX_IDinst_reg_out_A[22]),
    .ADR3(\DLX_IDinst_Imm[31] ),
    .O(\DLX_IFinst_PC<10>/GROM )
  );
  X_BUF \DLX_IFinst_PC<10>/XUSED  (
    .I(\DLX_IFinst_PC<10>/FROM ),
    .O(CHOICE4708)
  );
  X_BUF \DLX_IFinst_PC<10>/YUSED  (
    .I(\DLX_IFinst_PC<10>/GROM ),
    .O(CHOICE4060)
  );
  defparam DLX_IDinst_RegFile_11_4_680.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_11_4_680 (
    .I(DLX_MEMinst_RF_data_in[4]),
    .CE(DLX_IDinst__n0572),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_11_4)
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<2>_SW0 .INIT = 16'h5353;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<2>_SW0  (
    .ADR0(DLX_IDinst_reg_out_A[1]),
    .ADR1(DLX_IDinst_reg_out_A[2]),
    .ADR2(DLX_IDinst_reg_out_B[0]),
    .ADR3(VCC),
    .O(\DLX_IDinst_RegFile_11_4/FROM )
  );
  defparam \DLX_EXinst__n0007<0>23 .INIT = 16'h0B08;
  X_LUT4 \DLX_EXinst__n0007<0>23  (
    .ADR0(DLX_IDinst_reg_out_A[2]),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(DLX_IDinst_reg_out_B[0]),
    .ADR3(DLX_IDinst_reg_out_A[0]),
    .O(\DLX_IDinst_RegFile_11_4/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_11_4/XUSED  (
    .I(\DLX_IDinst_RegFile_11_4/FROM ),
    .O(N131631)
  );
  X_BUF \DLX_IDinst_RegFile_11_4/YUSED  (
    .I(\DLX_IDinst_RegFile_11_4/GROM ),
    .O(CHOICE5881)
  );
  defparam \DLX_EXinst__n0007<0>581_SW0 .INIT = 16'hFA50;
  X_LUT4 \DLX_EXinst__n0007<0>581_SW0  (
    .ADR0(\DLX_IDinst_Imm[1] ),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[1]),
    .ADR3(DLX_IDinst_reg_out_A[3]),
    .O(\DLX_IDinst_RegFile_6_23/FROM )
  );
  defparam \DLX_EXinst__n0007<0>36 .INIT = 16'hA808;
  X_LUT4 \DLX_EXinst__n0007<0>36  (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(DLX_IDinst_reg_out_A[1]),
    .ADR2(DLX_IDinst_reg_out_B[1]),
    .ADR3(DLX_IDinst_reg_out_A[3]),
    .O(\DLX_IDinst_RegFile_6_23/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_6_23/XUSED  (
    .I(\DLX_IDinst_RegFile_6_23/FROM ),
    .O(N164636)
  );
  X_BUF \DLX_IDinst_RegFile_6_23/YUSED  (
    .I(\DLX_IDinst_RegFile_6_23/GROM ),
    .O(CHOICE5886)
  );
  defparam \DLX_EXinst__n0007<16>79 .INIT = 16'hB0A0;
  X_LUT4 \DLX_EXinst__n0007<16>79  (
    .ADR0(DLX_EXinst__n0078),
    .ADR1(DLX_IDinst_reg_out_A[16]),
    .ADR2(DLX_IDinst_reg_out_B[16]),
    .ADR3(DLX_EXinst__n0079),
    .O(\DLX_IDinst_RegFile_6_16/FROM )
  );
  defparam \DLX_EXinst__n0007<24>9 .INIT = 16'hDC00;
  X_LUT4 \DLX_EXinst__n0007<24>9  (
    .ADR0(DLX_IDinst_reg_out_A[24]),
    .ADR1(DLX_EXinst__n0078),
    .ADR2(DLX_EXinst__n0079),
    .ADR3(DLX_IDinst_reg_out_B[24]),
    .O(\DLX_IDinst_RegFile_6_16/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_6_16/XUSED  (
    .I(\DLX_IDinst_RegFile_6_16/FROM ),
    .O(CHOICE4579)
  );
  X_BUF \DLX_IDinst_RegFile_6_16/YUSED  (
    .I(\DLX_IDinst_RegFile_6_16/GROM ),
    .O(CHOICE5585)
  );
  defparam \DLX_EXinst__n0007<7>241_SW0_SW0 .INIT = 16'hFF32;
  X_LUT4 \DLX_EXinst__n0007<7>241_SW0_SW0  (
    .ADR0(CHOICE3830),
    .ADR1(DLX_IDinst_reg_out_B[4]),
    .ADR2(CHOICE3827),
    .ADR3(CHOICE3841),
    .O(\N164583/FROM )
  );
  defparam \DLX_EXinst__n0007<7>241_SW0 .INIT = 16'hFFEC;
  X_LUT4 \DLX_EXinst__n0007<7>241_SW0  (
    .ADR0(CHOICE3821),
    .ADR1(CHOICE3838),
    .ADR2(DLX_IDinst_reg_out_A[7]),
    .ADR3(N164583),
    .O(\N164583/GROM )
  );
  X_BUF \N164583/XUSED  (
    .I(\N164583/FROM ),
    .O(N164583)
  );
  X_BUF \N164583/YUSED  (
    .I(\N164583/GROM ),
    .O(N163226)
  );
  defparam \DLX_EXinst__n0007<2>16 .INIT = 16'h3222;
  X_LUT4 \DLX_EXinst__n0007<2>16  (
    .ADR0(CHOICE5511),
    .ADR1(N146478),
    .ADR2(DLX_EXinst_N76285),
    .ADR3(\DLX_EXinst_Mshift__n0022_Sh[50] ),
    .O(\DLX_IDinst_RegFile_6_19/FROM )
  );
  defparam \DLX_EXinst__n0007<1>16 .INIT = 16'h3222;
  X_LUT4 \DLX_EXinst__n0007<1>16  (
    .ADR0(CHOICE5690),
    .ADR1(N146478),
    .ADR2(DLX_EXinst_N76285),
    .ADR3(\DLX_EXinst_Mshift__n0022_Sh[49] ),
    .O(\DLX_IDinst_RegFile_6_19/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_6_19/XUSED  (
    .I(\DLX_IDinst_RegFile_6_19/FROM ),
    .O(CHOICE5513)
  );
  X_BUF \DLX_IDinst_RegFile_6_19/YUSED  (
    .I(\DLX_IDinst_RegFile_6_19/GROM ),
    .O(CHOICE5692)
  );
  defparam \DLX_EXinst__n0007<29>13 .INIT = 16'hAA08;
  X_LUT4 \DLX_EXinst__n0007<29>13  (
    .ADR0(DLX_IDinst_reg_out_A[29]),
    .ADR1(DLX_EXinst__n0054),
    .ADR2(\DLX_IDinst_Imm[31] ),
    .ADR3(DLX_EXinst__n0053),
    .O(\CHOICE4779/FROM )
  );
  defparam \DLX_EXinst__n0007<17>9 .INIT = 16'hBA00;
  X_LUT4 \DLX_EXinst__n0007<17>9  (
    .ADR0(DLX_EXinst__n0053),
    .ADR1(\DLX_IDinst_Imm[31] ),
    .ADR2(DLX_EXinst__n0054),
    .ADR3(DLX_IDinst_reg_out_A[17]),
    .O(\CHOICE4779/GROM )
  );
  X_BUF \CHOICE4779/XUSED  (
    .I(\CHOICE4779/FROM ),
    .O(CHOICE4779)
  );
  X_BUF \CHOICE4779/YUSED  (
    .I(\CHOICE4779/GROM ),
    .O(CHOICE5354)
  );
  defparam DLX_EXinst_Ker74372113.INIT = 16'h00C0;
  X_LUT4 DLX_EXinst_Ker74372113 (
    .ADR0(VCC),
    .ADR1(\DLX_EXinst_Mshift__n0019_Sh[26] ),
    .ADR2(DLX_IDinst_reg_out_B_2_1),
    .ADR3(DLX_IDinst_reg_out_B[3]),
    .O(\CHOICE3133/FROM )
  );
  defparam \DLX_EXinst__n0007<0>68 .INIT = 16'hAFAC;
  X_LUT4 \DLX_EXinst__n0007<0>68  (
    .ADR0(\DLX_EXinst_Mshift__n0019_Sh[8] ),
    .ADR1(CHOICE5881),
    .ADR2(DLX_IDinst_reg_out_B[3]),
    .ADR3(CHOICE5886),
    .O(\CHOICE3133/GROM )
  );
  X_BUF \CHOICE3133/XUSED  (
    .I(\CHOICE3133/FROM ),
    .O(CHOICE3133)
  );
  X_BUF \CHOICE3133/YUSED  (
    .I(\CHOICE3133/GROM ),
    .O(CHOICE5890)
  );
  defparam \DLX_EXinst__n0007<26>9 .INIT = 16'hAA08;
  X_LUT4 \DLX_EXinst__n0007<26>9  (
    .ADR0(DLX_IDinst_reg_out_A[26]),
    .ADR1(DLX_EXinst__n0054),
    .ADR2(\DLX_IDinst_Imm[31] ),
    .ADR3(DLX_EXinst__n0053),
    .O(\CHOICE4991/FROM )
  );
  defparam \DLX_EXinst__n0007<26>139 .INIT = 16'h00FE;
  X_LUT4 \DLX_EXinst__n0007<26>139  (
    .ADR0(CHOICE4991),
    .ADR1(CHOICE5017),
    .ADR2(CHOICE4992),
    .ADR3(DLX_EXinst__n0036),
    .O(\CHOICE4991/GROM )
  );
  X_BUF \CHOICE4991/XUSED  (
    .I(\CHOICE4991/FROM ),
    .O(CHOICE4991)
  );
  X_BUF \CHOICE4991/YUSED  (
    .I(\CHOICE4991/GROM ),
    .O(CHOICE5020)
  );
  defparam \DLX_EXinst__n0007<9>141 .INIT = 16'hB0A0;
  X_LUT4 \DLX_EXinst__n0007<9>141  (
    .ADR0(DLX_EXinst__n0053),
    .ADR1(\DLX_IDinst_Imm[9] ),
    .ADR2(DLX_IDinst_reg_out_A[9]),
    .ADR3(DLX_EXinst__n0054),
    .O(\CHOICE4539/FROM )
  );
  defparam \DLX_EXinst__n0007<1>29 .INIT = 16'hDC00;
  X_LUT4 \DLX_EXinst__n0007<1>29  (
    .ADR0(\DLX_IDinst_Imm[1] ),
    .ADR1(DLX_EXinst__n0053),
    .ADR2(DLX_EXinst__n0054),
    .ADR3(DLX_IDinst_reg_out_A[1]),
    .O(\CHOICE4539/GROM )
  );
  X_BUF \CHOICE4539/XUSED  (
    .I(\CHOICE4539/FROM ),
    .O(CHOICE4539)
  );
  X_BUF \CHOICE4539/YUSED  (
    .I(\CHOICE4539/GROM ),
    .O(CHOICE5696)
  );
  defparam \DLX_EXinst__n0007<3>48 .INIT = 16'hAE04;
  X_LUT4 \DLX_EXinst__n0007<3>48  (
    .ADR0(\DLX_IDinst_Imm[3] ),
    .ADR1(DLX_IDinst_reg_out_A[3]),
    .ADR2(DLX_EXinst_N73211),
    .ADR3(\DLX_EXinst_Mshift__n0022_Sh[11] ),
    .O(\CHOICE5447/FROM )
  );
  defparam \DLX_EXinst__n0007<1>48 .INIT = 16'hC5C0;
  X_LUT4 \DLX_EXinst__n0007<1>48  (
    .ADR0(DLX_EXinst_N73211),
    .ADR1(\DLX_EXinst_Mshift__n0022_Sh[9] ),
    .ADR2(\DLX_IDinst_Imm[3] ),
    .ADR3(DLX_IDinst_reg_out_A[1]),
    .O(\CHOICE5447/GROM )
  );
  X_BUF \CHOICE5447/XUSED  (
    .I(\CHOICE5447/FROM ),
    .O(CHOICE5447)
  );
  X_BUF \CHOICE5447/YUSED  (
    .I(\CHOICE5447/GROM ),
    .O(CHOICE5702)
  );
  defparam \DLX_EXinst__n0007<8>181 .INIT = 16'hF040;
  X_LUT4 \DLX_EXinst__n0007<8>181  (
    .ADR0(\DLX_IDinst_Imm[8] ),
    .ADR1(DLX_EXinst__n0054),
    .ADR2(DLX_IDinst_reg_out_A[8]),
    .ADR3(DLX_EXinst__n0053),
    .O(\CHOICE5170/FROM )
  );
  defparam \DLX_EXinst__n0007<19>9 .INIT = 16'hCE00;
  X_LUT4 \DLX_EXinst__n0007<19>9  (
    .ADR0(DLX_EXinst__n0054),
    .ADR1(DLX_EXinst__n0053),
    .ADR2(\DLX_IDinst_Imm[31] ),
    .ADR3(DLX_IDinst_reg_out_A[19]),
    .O(\CHOICE5170/GROM )
  );
  X_BUF \CHOICE5170/XUSED  (
    .I(\CHOICE5170/FROM ),
    .O(CHOICE5170)
  );
  X_BUF \CHOICE5170/YUSED  (
    .I(\CHOICE5170/GROM ),
    .O(CHOICE5275)
  );
  defparam \DLX_EXinst_Mshift__n0021_Sh<2>_SW0 .INIT = 16'h505F;
  X_LUT4 \DLX_EXinst_Mshift__n0021_Sh<2>_SW0  (
    .ADR0(DLX_IDinst_reg_out_A[1]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_Imm_0_1),
    .ADR3(DLX_IDinst_reg_out_A[2]),
    .O(\N131693/FROM )
  );
  defparam \DLX_EXinst__n0007<2>29 .INIT = 16'hF040;
  X_LUT4 \DLX_EXinst__n0007<2>29  (
    .ADR0(\DLX_IDinst_Imm[2] ),
    .ADR1(DLX_EXinst__n0054),
    .ADR2(DLX_IDinst_reg_out_A[2]),
    .ADR3(DLX_EXinst__n0053),
    .O(\N131693/GROM )
  );
  X_BUF \N131693/XUSED  (
    .I(\N131693/FROM ),
    .O(N131693)
  );
  X_BUF \N131693/YUSED  (
    .I(\N131693/GROM ),
    .O(CHOICE5517)
  );
  defparam \DLX_EXinst__n0007<3>79 .INIT = 16'h4448;
  X_LUT4 \DLX_EXinst__n0007<3>79  (
    .ADR0(DLX_IDinst_IR_opcode_field[1]),
    .ADR1(DLX_EXinst_N76011),
    .ADR2(DLX_IDinst_reg_out_A[3]),
    .ADR3(DLX_IDinst_IR_opcode_field[0]),
    .O(\CHOICE5455/FROM )
  );
  defparam \DLX_EXinst__n0007<1>79 .INIT = 16'h2228;
  X_LUT4 \DLX_EXinst__n0007<1>79  (
    .ADR0(DLX_EXinst_N76011),
    .ADR1(DLX_IDinst_IR_opcode_field[1]),
    .ADR2(DLX_IDinst_reg_out_A[1]),
    .ADR3(DLX_IDinst_IR_opcode_field[0]),
    .O(\CHOICE5455/GROM )
  );
  X_BUF \CHOICE5455/XUSED  (
    .I(\CHOICE5455/FROM ),
    .O(CHOICE5455)
  );
  X_BUF \CHOICE5455/YUSED  (
    .I(\CHOICE5455/GROM ),
    .O(CHOICE5710)
  );
  defparam DLX_IDinst_RegFile_27_10_681.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_27_10_681 (
    .I(DLX_IDinst_WB_data_eff[10]),
    .CE(DLX_IDinst__n0604),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_27_10)
  );
  defparam \DLX_EXinst__n0007<30>29 .INIT = 16'hF044;
  X_LUT4 \DLX_EXinst__n0007<30>29  (
    .ADR0(DLX_EXinst_N73211),
    .ADR1(DLX_IDinst_reg_out_A[30]),
    .ADR2(\DLX_EXinst_Mshift__n0021_Sh[22] ),
    .ADR3(\DLX_IDinst_Imm[3] ),
    .O(\CHOICE4716/FROM )
  );
  defparam \DLX_EXinst__n0007<2>48 .INIT = 16'hF202;
  X_LUT4 \DLX_EXinst__n0007<2>48  (
    .ADR0(DLX_IDinst_reg_out_A[2]),
    .ADR1(DLX_EXinst_N73211),
    .ADR2(\DLX_IDinst_Imm[3] ),
    .ADR3(\DLX_EXinst_Mshift__n0022_Sh[10] ),
    .O(\CHOICE4716/GROM )
  );
  X_BUF \CHOICE4716/XUSED  (
    .I(\CHOICE4716/FROM ),
    .O(CHOICE4716)
  );
  X_BUF \CHOICE4716/YUSED  (
    .I(\CHOICE4716/GROM ),
    .O(CHOICE5523)
  );
  defparam \DLX_EXinst__n0007<1>98 .INIT = 16'hFEEE;
  X_LUT4 \DLX_EXinst__n0007<1>98  (
    .ADR0(N163668),
    .ADR1(CHOICE5713),
    .ADR2(CHOICE5710),
    .ADR3(\DLX_IDinst_Imm[1] ),
    .O(\CHOICE5715/FROM )
  );
  defparam \DLX_EXinst__n0007<1>127 .INIT = 16'h3332;
  X_LUT4 \DLX_EXinst__n0007<1>127  (
    .ADR0(CHOICE5692),
    .ADR1(DLX_EXinst__n0036),
    .ADR2(CHOICE5696),
    .ADR3(CHOICE5715),
    .O(\CHOICE5715/GROM )
  );
  X_BUF \CHOICE5715/XUSED  (
    .I(\CHOICE5715/FROM ),
    .O(CHOICE5715)
  );
  X_BUF \CHOICE5715/YUSED  (
    .I(\CHOICE5715/GROM ),
    .O(CHOICE5717)
  );
  defparam \DLX_EXinst__n0007<21>92_SW0 .INIT = 16'h5600;
  X_LUT4 \DLX_EXinst__n0007<21>92_SW0  (
    .ADR0(DLX_IDinst_IR_opcode_field[1]),
    .ADR1(DLX_IDinst_IR_opcode_field[0]),
    .ADR2(DLX_IDinst_reg_out_A[21]),
    .ADR3(DLX_EXinst_N76011),
    .O(\N163704/FROM )
  );
  defparam \DLX_EXinst__n0007<2>79 .INIT = 16'h3600;
  X_LUT4 \DLX_EXinst__n0007<2>79  (
    .ADR0(DLX_IDinst_IR_opcode_field[0]),
    .ADR1(DLX_IDinst_IR_opcode_field[1]),
    .ADR2(DLX_IDinst_reg_out_A[2]),
    .ADR3(DLX_EXinst_N76011),
    .O(\N163704/GROM )
  );
  X_BUF \N163704/XUSED  (
    .I(\N163704/FROM ),
    .O(N163704)
  );
  X_BUF \N163704/YUSED  (
    .I(\N163704/GROM ),
    .O(CHOICE5531)
  );
  defparam \DLX_EXinst__n0007<31>45_SW0 .INIT = 16'hFCFE;
  X_LUT4 \DLX_EXinst__n0007<31>45_SW0  (
    .ADR0(N148609),
    .ADR1(DLX_EXinst__n0083),
    .ADR2(DLX_EXinst__n0078),
    .ADR3(DLX_IDinst_reg_out_B[5]),
    .O(\N163931/FROM )
  );
  defparam \DLX_EXinst__n0007<4>15 .INIT = 16'hF8F8;
  X_LUT4 \DLX_EXinst__n0007<4>15  (
    .ADR0(N148609),
    .ADR1(DLX_EXinst_N74966),
    .ADR2(DLX_EXinst__n0078),
    .ADR3(VCC),
    .O(\N163931/GROM )
  );
  X_BUF \N163931/XUSED  (
    .I(\N163931/FROM ),
    .O(N163931)
  );
  X_BUF \N163931/YUSED  (
    .I(\N163931/GROM ),
    .O(CHOICE4328)
  );
  defparam \DLX_EXinst__n0007<4>24 .INIT = 16'hFBF8;
  X_LUT4 \DLX_EXinst__n0007<4>24  (
    .ADR0(DLX_EXinst__n0077),
    .ADR1(DLX_IDinst_reg_out_A[4]),
    .ADR2(CHOICE4329),
    .ADR3(DLX_EXinst__n0079),
    .O(\CHOICE4330/FROM )
  );
  defparam \DLX_EXinst__n0007<4>41 .INIT = 16'hF888;
  X_LUT4 \DLX_EXinst__n0007<4>41  (
    .ADR0(N134884),
    .ADR1(DLX_EXinst_ALU_result[4]),
    .ADR2(DLX_IDinst_reg_out_B[4]),
    .ADR3(CHOICE4330),
    .O(\CHOICE4330/GROM )
  );
  X_BUF \CHOICE4330/XUSED  (
    .I(\CHOICE4330/FROM ),
    .O(CHOICE4330)
  );
  X_BUF \CHOICE4330/YUSED  (
    .I(\CHOICE4330/GROM ),
    .O(CHOICE4332)
  );
  defparam DLX_IDinst_RegFile_18_27_682.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_18_27_682 (
    .I(DLX_IDinst_WB_data_eff[27]),
    .CE(DLX_IDinst__n0586),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_18_27)
  );
  defparam \DLX_EXinst__n0007<8>229 .INIT = 16'hC0C0;
  X_LUT4 \DLX_EXinst__n0007<8>229  (
    .ADR0(VCC),
    .ADR1(CHOICE5185),
    .ADR2(N147520),
    .ADR3(VCC),
    .O(\CHOICE5186/FROM )
  );
  defparam \DLX_EXinst__n0007<2>88 .INIT = 16'h8080;
  X_LUT4 \DLX_EXinst__n0007<2>88  (
    .ADR0(\DLX_IDinst_Imm[4] ),
    .ADR1(N137608),
    .ADR2(N147520),
    .ADR3(VCC),
    .O(\CHOICE5186/GROM )
  );
  X_BUF \CHOICE5186/XUSED  (
    .I(\CHOICE5186/FROM ),
    .O(CHOICE5186)
  );
  X_BUF \CHOICE5186/YUSED  (
    .I(\CHOICE5186/GROM ),
    .O(CHOICE5534)
  );
  defparam DLX_EXinst_Ker7551863.INIT = 16'h0040;
  X_LUT4 DLX_EXinst_Ker7551863 (
    .ADR0(DLX_IDinst_reg_out_B_2_1),
    .ADR1(DLX_EXinst_N76421),
    .ADR2(\DLX_EXinst_Mshift__n0024_Sh[30] ),
    .ADR3(DLX_IDinst_reg_out_B_3_1),
    .O(\CHOICE2058/FROM )
  );
  defparam \DLX_EXinst__n0007<4>17 .INIT = 16'hFCF0;
  X_LUT4 \DLX_EXinst__n0007<4>17  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N76421),
    .ADR2(CHOICE4328),
    .ADR3(\DLX_EXinst_Mshift__n0024_Sh[52] ),
    .O(\CHOICE2058/GROM )
  );
  X_BUF \CHOICE2058/XUSED  (
    .I(\CHOICE2058/FROM ),
    .O(CHOICE2058)
  );
  X_BUF \CHOICE2058/YUSED  (
    .I(\CHOICE2058/GROM ),
    .O(CHOICE4329)
  );
  defparam \DLX_EXinst__n0007<2>98 .INIT = 16'hFFF8;
  X_LUT4 \DLX_EXinst__n0007<2>98  (
    .ADR0(CHOICE5531),
    .ADR1(\DLX_IDinst_Imm[2] ),
    .ADR2(CHOICE5534),
    .ADR3(CHOICE5526),
    .O(\CHOICE5536/FROM )
  );
  defparam \DLX_EXinst__n0007<2>127 .INIT = 16'h5554;
  X_LUT4 \DLX_EXinst__n0007<2>127  (
    .ADR0(DLX_EXinst__n0036),
    .ADR1(CHOICE5513),
    .ADR2(CHOICE5517),
    .ADR3(CHOICE5536),
    .O(\CHOICE5536/GROM )
  );
  X_BUF \CHOICE5536/XUSED  (
    .I(\CHOICE5536/FROM ),
    .O(CHOICE5536)
  );
  X_BUF \CHOICE5536/YUSED  (
    .I(\CHOICE5536/GROM ),
    .O(CHOICE5538)
  );
  defparam \DLX_EXinst__n0007<13>33 .INIT = 16'hCA00;
  X_LUT4 \DLX_EXinst__n0007<13>33  (
    .ADR0(DLX_EXinst_N74451),
    .ADR1(DLX_EXinst_N74726),
    .ADR2(DLX_IDinst_reg_out_B[2]),
    .ADR3(DLX_EXinst_N72710),
    .O(\CHOICE3718/FROM )
  );
  defparam \DLX_EXinst__n0007<5>32 .INIT = 16'hC480;
  X_LUT4 \DLX_EXinst__n0007<5>32  (
    .ADR0(DLX_IDinst_reg_out_B[2]),
    .ADR1(DLX_EXinst_N72710),
    .ADR2(DLX_EXinst_N74696),
    .ADR3(N133480),
    .O(\CHOICE3718/GROM )
  );
  X_BUF \CHOICE3718/XUSED  (
    .I(\CHOICE3718/FROM ),
    .O(CHOICE3718)
  );
  X_BUF \CHOICE3718/YUSED  (
    .I(\CHOICE3718/GROM ),
    .O(CHOICE3945)
  );
  defparam \DLX_EXinst__n0007<3>98 .INIT = 16'hFFEC;
  X_LUT4 \DLX_EXinst__n0007<3>98  (
    .ADR0(CHOICE5455),
    .ADR1(CHOICE5458),
    .ADR2(\DLX_IDinst_Imm[3] ),
    .ADR3(N163542),
    .O(\CHOICE5460/FROM )
  );
  defparam \DLX_EXinst__n0007<3>127 .INIT = 16'h3332;
  X_LUT4 \DLX_EXinst__n0007<3>127  (
    .ADR0(CHOICE5441),
    .ADR1(DLX_EXinst__n0036),
    .ADR2(CHOICE5437),
    .ADR3(CHOICE5460),
    .O(\CHOICE5460/GROM )
  );
  X_BUF \CHOICE5460/XUSED  (
    .I(\CHOICE5460/FROM ),
    .O(CHOICE5460)
  );
  X_BUF \CHOICE5460/YUSED  (
    .I(\CHOICE5460/GROM ),
    .O(CHOICE5462)
  );
  defparam \DLX_EXinst__n0007<9>51 .INIT = 16'hEFEA;
  X_LUT4 \DLX_EXinst__n0007<9>51  (
    .ADR0(DLX_EXinst_N74245),
    .ADR1(DLX_EXinst__n0077),
    .ADR2(DLX_IDinst_reg_out_B[9]),
    .ADR3(DLX_EXinst__n0079),
    .O(\CHOICE4519/FROM )
  );
  defparam \DLX_EXinst__n0007<6>13 .INIT = 16'hFDEC;
  X_LUT4 \DLX_EXinst__n0007<6>13  (
    .ADR0(DLX_IDinst_reg_out_B[6]),
    .ADR1(DLX_EXinst_N74245),
    .ADR2(DLX_EXinst__n0077),
    .ADR3(DLX_EXinst__n0079),
    .O(\CHOICE4519/GROM )
  );
  X_BUF \CHOICE4519/XUSED  (
    .I(\CHOICE4519/FROM ),
    .O(CHOICE4519)
  );
  X_BUF \CHOICE4519/YUSED  (
    .I(\CHOICE4519/GROM ),
    .O(CHOICE3880)
  );
  defparam \DLX_EXinst__n0007<6>38 .INIT = 16'h0008;
  X_LUT4 \DLX_EXinst__n0007<6>38  (
    .ADR0(DLX_EXinst_N72908),
    .ADR1(DLX_EXinst__n0080),
    .ADR2(N148323),
    .ADR3(DLX_IDinst_reg_out_B[3]),
    .O(\CHOICE3889/FROM )
  );
  defparam \DLX_EXinst__n0007<5>38 .INIT = 16'h0020;
  X_LUT4 \DLX_EXinst__n0007<5>38  (
    .ADR0(DLX_EXinst_N72903),
    .ADR1(DLX_IDinst_reg_out_B[3]),
    .ADR2(DLX_EXinst__n0080),
    .ADR3(N148323),
    .O(\CHOICE3889/GROM )
  );
  X_BUF \CHOICE3889/XUSED  (
    .I(\CHOICE3889/FROM ),
    .O(CHOICE3889)
  );
  X_BUF \CHOICE3889/YUSED  (
    .I(\CHOICE3889/GROM ),
    .O(CHOICE3948)
  );
  defparam \DLX_EXinst__n0007<15>38 .INIT = 16'hA0C0;
  X_LUT4 \DLX_EXinst__n0007<15>38  (
    .ADR0(DLX_EXinst_N74976),
    .ADR1(DLX_EXinst_N74686),
    .ADR2(DLX_EXinst_N72710),
    .ADR3(DLX_IDinst_reg_out_B[2]),
    .O(\CHOICE4273/FROM )
  );
  defparam \DLX_EXinst__n0007<6>32 .INIT = 16'h8A80;
  X_LUT4 \DLX_EXinst__n0007<6>32  (
    .ADR0(DLX_EXinst_N72710),
    .ADR1(DLX_EXinst_N74681),
    .ADR2(DLX_IDinst_reg_out_B[2]),
    .ADR3(N133408),
    .O(\CHOICE4273/GROM )
  );
  X_BUF \CHOICE4273/XUSED  (
    .I(\CHOICE4273/FROM ),
    .O(CHOICE4273)
  );
  X_BUF \CHOICE4273/YUSED  (
    .I(\CHOICE4273/GROM ),
    .O(CHOICE3886)
  );
  defparam \DLX_EXinst__n0007<8>12 .INIT = 16'hCC40;
  X_LUT4 \DLX_EXinst__n0007<8>12  (
    .ADR0(DLX_IDinst_reg_out_A[8]),
    .ADR1(DLX_IDinst_reg_out_B[8]),
    .ADR2(DLX_EXinst__n0079),
    .ADR3(DLX_EXinst__n0078),
    .O(\CHOICE5127/FROM )
  );
  defparam \DLX_EXinst__n0007<5>82 .INIT = 16'hCC40;
  X_LUT4 \DLX_EXinst__n0007<5>82  (
    .ADR0(DLX_IDinst_reg_out_A[5]),
    .ADR1(DLX_IDinst_reg_out_B[5]),
    .ADR2(DLX_EXinst__n0079),
    .ADR3(DLX_EXinst__n0078),
    .O(\CHOICE5127/GROM )
  );
  X_BUF \CHOICE5127/XUSED  (
    .I(\CHOICE5127/FROM ),
    .O(CHOICE5127)
  );
  X_BUF \CHOICE5127/YUSED  (
    .I(\CHOICE5127/GROM ),
    .O(CHOICE3956)
  );
  defparam \DLX_EXinst__n0007<8>47 .INIT = 16'hFBEA;
  X_LUT4 \DLX_EXinst__n0007<8>47  (
    .ADR0(DLX_EXinst_N74245),
    .ADR1(DLX_IDinst_reg_out_B[8]),
    .ADR2(DLX_EXinst__n0077),
    .ADR3(DLX_EXinst__n0079),
    .O(\CHOICE5139/FROM )
  );
  defparam \DLX_EXinst__n0007<7>13 .INIT = 16'hFCEE;
  X_LUT4 \DLX_EXinst__n0007<7>13  (
    .ADR0(DLX_EXinst__n0079),
    .ADR1(DLX_EXinst_N74245),
    .ADR2(DLX_EXinst__n0077),
    .ADR3(DLX_IDinst_reg_out_B[7]),
    .O(\CHOICE5139/GROM )
  );
  X_BUF \CHOICE5139/XUSED  (
    .I(\CHOICE5139/FROM ),
    .O(CHOICE5139)
  );
  X_BUF \CHOICE5139/YUSED  (
    .I(\CHOICE5139/GROM ),
    .O(CHOICE3821)
  );
  defparam \DLX_EXinst__n0007<12>33 .INIT = 16'hC088;
  X_LUT4 \DLX_EXinst__n0007<12>33  (
    .ADR0(DLX_EXinst_N74446),
    .ADR1(DLX_EXinst_N72710),
    .ADR2(DLX_EXinst_N74721),
    .ADR3(DLX_IDinst_reg_out_B[2]),
    .O(\CHOICE3773/FROM )
  );
  defparam \DLX_EXinst__n0007<7>32 .INIT = 16'hC808;
  X_LUT4 \DLX_EXinst__n0007<7>32  (
    .ADR0(N133552),
    .ADR1(DLX_EXinst_N72710),
    .ADR2(DLX_IDinst_reg_out_B[2]),
    .ADR3(DLX_EXinst_N74991),
    .O(\CHOICE3773/GROM )
  );
  X_BUF \CHOICE3773/XUSED  (
    .I(\CHOICE3773/FROM ),
    .O(CHOICE3773)
  );
  X_BUF \CHOICE3773/YUSED  (
    .I(\CHOICE3773/GROM ),
    .O(CHOICE3827)
  );
  defparam \DLX_EXinst__n0007<1>165 .INIT = 16'hB0A0;
  X_LUT4 \DLX_EXinst__n0007<1>165  (
    .ADR0(DLX_EXinst__n0078),
    .ADR1(DLX_IDinst_reg_out_A[1]),
    .ADR2(DLX_IDinst_reg_out_B[1]),
    .ADR3(DLX_EXinst__n0079),
    .O(\CHOICE5724/FROM )
  );
  defparam \DLX_EXinst__n0007<6>82 .INIT = 16'hCC08;
  X_LUT4 \DLX_EXinst__n0007<6>82  (
    .ADR0(DLX_EXinst__n0079),
    .ADR1(DLX_IDinst_reg_out_B[6]),
    .ADR2(DLX_IDinst_reg_out_A[6]),
    .ADR3(DLX_EXinst__n0078),
    .O(\CHOICE5724/GROM )
  );
  X_BUF \CHOICE5724/XUSED  (
    .I(\CHOICE5724/FROM ),
    .O(CHOICE5724)
  );
  X_BUF \CHOICE5724/YUSED  (
    .I(\CHOICE5724/GROM ),
    .O(CHOICE3897)
  );
  defparam DLX_EXinst_Ker764771.INIT = 16'h4400;
  X_LUT4 DLX_EXinst_Ker764771 (
    .ADR0(N148323),
    .ADR1(DLX_EXinst_N75964),
    .ADR2(VCC),
    .ADR3(DLX_EXinst__n0080),
    .O(\DLX_EXinst_N76479/FROM )
  );
  defparam \DLX_EXinst__n0007<7>38 .INIT = 16'h0200;
  X_LUT4 \DLX_EXinst__n0007<7>38  (
    .ADR0(DLX_EXinst_N72913),
    .ADR1(N148323),
    .ADR2(DLX_IDinst_reg_out_B[3]),
    .ADR3(DLX_EXinst__n0080),
    .O(\DLX_EXinst_N76479/GROM )
  );
  X_BUF \DLX_EXinst_N76479/XUSED  (
    .I(\DLX_EXinst_N76479/FROM ),
    .O(DLX_EXinst_N76479)
  );
  X_BUF \DLX_EXinst_N76479/YUSED  (
    .I(\DLX_EXinst_N76479/GROM ),
    .O(CHOICE3830)
  );
  defparam \DLX_EXinst__n0007<1>189 .INIT = 16'hD800;
  X_LUT4 \DLX_EXinst__n0007<1>189  (
    .ADR0(DLX_IDinst_reg_out_B[2]),
    .ADR1(N133480),
    .ADR2(CHOICE5729),
    .ADR3(DLX_EXinst_N76457),
    .O(\CHOICE5732/FROM )
  );
  defparam \DLX_EXinst__n0007<8>25 .INIT = 16'hA088;
  X_LUT4 \DLX_EXinst__n0007<8>25  (
    .ADR0(DLX_EXinst_N76457),
    .ADR1(DLX_EXinst_N74691),
    .ADR2(DLX_EXinst_N74446),
    .ADR3(DLX_IDinst_reg_out_B[2]),
    .O(\CHOICE5732/GROM )
  );
  X_BUF \CHOICE5732/XUSED  (
    .I(\CHOICE5732/FROM ),
    .O(CHOICE5732)
  );
  X_BUF \CHOICE5732/YUSED  (
    .I(\CHOICE5732/GROM ),
    .O(CHOICE5132)
  );
  defparam \DLX_EXinst__n0007<14>13 .INIT = 16'hF020;
  X_LUT4 \DLX_EXinst__n0007<14>13  (
    .ADR0(DLX_EXinst__n0079),
    .ADR1(DLX_IDinst_reg_out_A[14]),
    .ADR2(DLX_IDinst_reg_out_B[14]),
    .ADR3(DLX_EXinst__n0078),
    .O(\CHOICE3656/FROM )
  );
  defparam \DLX_EXinst__n0007<7>82 .INIT = 16'hF400;
  X_LUT4 \DLX_EXinst__n0007<7>82  (
    .ADR0(DLX_IDinst_reg_out_A[7]),
    .ADR1(DLX_EXinst__n0079),
    .ADR2(DLX_EXinst__n0078),
    .ADR3(DLX_IDinst_reg_out_B[7]),
    .O(\CHOICE3656/GROM )
  );
  X_BUF \CHOICE3656/XUSED  (
    .I(\CHOICE3656/FROM ),
    .O(CHOICE3656)
  );
  X_BUF \CHOICE3656/YUSED  (
    .I(\CHOICE3656/GROM ),
    .O(CHOICE3838)
  );
  defparam \DLX_EXinst__n0007<15>10 .INIT = 16'hCC40;
  X_LUT4 \DLX_EXinst__n0007<15>10  (
    .ADR0(DLX_IDinst_reg_out_A[15]),
    .ADR1(DLX_IDinst_reg_out_B[15]),
    .ADR2(DLX_EXinst__n0079),
    .ADR3(DLX_EXinst__n0078),
    .O(\CHOICE4263/FROM )
  );
  defparam \DLX_EXinst__n0007<9>12 .INIT = 16'hC0E0;
  X_LUT4 \DLX_EXinst__n0007<9>12  (
    .ADR0(DLX_EXinst__n0079),
    .ADR1(DLX_EXinst__n0078),
    .ADR2(DLX_IDinst_reg_out_B[9]),
    .ADR3(DLX_IDinst_reg_out_A[9]),
    .O(\CHOICE4263/GROM )
  );
  X_BUF \CHOICE4263/XUSED  (
    .I(\CHOICE4263/FROM ),
    .O(CHOICE4263)
  );
  X_BUF \CHOICE4263/YUSED  (
    .I(\CHOICE4263/GROM ),
    .O(CHOICE4505)
  );
  defparam \DLX_EXinst__n0007<3>189 .INIT = 16'hB080;
  X_LUT4 \DLX_EXinst__n0007<3>189  (
    .ADR0(N133552),
    .ADR1(DLX_IDinst_reg_out_B[2]),
    .ADR2(DLX_EXinst_N76457),
    .ADR3(CHOICE5474),
    .O(\CHOICE5477/FROM )
  );
  defparam \DLX_EXinst__n0007<9>25 .INIT = 16'hC480;
  X_LUT4 \DLX_EXinst__n0007<9>25  (
    .ADR0(DLX_IDinst_reg_out_B[2]),
    .ADR1(DLX_EXinst_N76457),
    .ADR2(DLX_EXinst_N74451),
    .ADR3(DLX_EXinst_N74696),
    .O(\CHOICE5477/GROM )
  );
  X_BUF \CHOICE5477/XUSED  (
    .I(\CHOICE5477/FROM ),
    .O(CHOICE5477)
  );
  X_BUF \CHOICE5477/YUSED  (
    .I(\CHOICE5477/GROM ),
    .O(CHOICE4510)
  );
  X_ZERO \vga_top_vga1_helpme/LOGIC_ZERO_683  (
    .O(\vga_top_vga1_helpme/LOGIC_ZERO )
  );
  defparam vga_top_vga1__n00101.INIT = 16'hFFFC;
  X_LUT4 vga_top_vga1__n00101 (
    .ADR0(VCC),
    .ADR1(vga_top_vga1__n0033),
    .ADR2(vga_top_vga1_helpme),
    .ADR3(vga_top_vga1__n0034),
    .O(\vga_top_vga1_helpme/GROM )
  );
  X_BUF \vga_top_vga1_helpme/YUSED  (
    .I(\vga_top_vga1_helpme/GROM ),
    .O(vga_top_vga1__n0010)
  );
  defparam \DLX_EXinst__n0007<10>81_SW0 .INIT = 16'hF888;
  X_LUT4 \DLX_EXinst__n0007<10>81_SW0  (
    .ADR0(DLX_EXinst_N75983),
    .ADR1(N138249),
    .ADR2(CHOICE4459),
    .ADR3(DLX_IDinst_reg_out_A[10]),
    .O(\N163728/FROM )
  );
  defparam \DLX_EXinst__n0007<10>81 .INIT = 16'hFFEA;
  X_LUT4 \DLX_EXinst__n0007<10>81  (
    .ADR0(CHOICE4465),
    .ADR1(N134884),
    .ADR2(DLX_EXinst_ALU_result[10]),
    .ADR3(N163728),
    .O(\N163728/GROM )
  );
  X_BUF \N163728/XUSED  (
    .I(\N163728/FROM ),
    .O(N163728)
  );
  X_BUF \N163728/YUSED  (
    .I(\N163728/GROM ),
    .O(CHOICE4467)
  );
  defparam \DLX_EXinst__n0007<10>65_SW0 .INIT = 16'h0777;
  X_LUT4 \DLX_EXinst__n0007<10>65_SW0  (
    .ADR0(DLX_EXinst_N76268),
    .ADR1(\DLX_EXinst_Mshift__n0023_Sh[42] ),
    .ADR2(DLX_EXinst_N76431),
    .ADR3(\DLX_EXinst_Mshift__n0024_Sh[58] ),
    .O(\N164228/FROM )
  );
  defparam \DLX_EXinst__n0007<10>65 .INIT = 16'h0001;
  X_LUT4 \DLX_EXinst__n0007<10>65  (
    .ADR0(CHOICE3592),
    .ADR1(CHOICE3576),
    .ADR2(CHOICE3570),
    .ADR3(N164228),
    .O(\N164228/GROM )
  );
  X_BUF \N164228/XUSED  (
    .I(\N164228/FROM ),
    .O(N164228)
  );
  X_BUF \N164228/YUSED  (
    .I(\N164228/GROM ),
    .O(CHOICE4465)
  );
  defparam \DLX_EXinst__n0007<11>65_SW0 .INIT = 16'h0777;
  X_LUT4 \DLX_EXinst__n0007<11>65_SW0  (
    .ADR0(DLX_EXinst_N76268),
    .ADR1(\DLX_EXinst_Mshift__n0023_Sh[43] ),
    .ADR2(DLX_EXinst_N76431),
    .ADR3(\DLX_EXinst_Mshift__n0024_Sh[59] ),
    .O(\N163979/FROM )
  );
  defparam \DLX_EXinst__n0007<11>65 .INIT = 16'h0001;
  X_LUT4 \DLX_EXinst__n0007<11>65  (
    .ADR0(CHOICE3576),
    .ADR1(CHOICE3570),
    .ADR2(CHOICE3592),
    .ADR3(N163979),
    .O(\N163979/GROM )
  );
  X_BUF \N163979/XUSED  (
    .I(\N163979/FROM ),
    .O(N163979)
  );
  X_BUF \N163979/YUSED  (
    .I(\N163979/GROM ),
    .O(CHOICE4405)
  );
  defparam \DLX_EXinst__n0007<11>81_SW0 .INIT = 16'hF888;
  X_LUT4 \DLX_EXinst__n0007<11>81_SW0  (
    .ADR0(CHOICE4399),
    .ADR1(DLX_IDinst_reg_out_A[11]),
    .ADR2(N137952),
    .ADR3(DLX_EXinst_N75983),
    .O(\N163286/FROM )
  );
  defparam \DLX_EXinst__n0007<11>81 .INIT = 16'hFFEC;
  X_LUT4 \DLX_EXinst__n0007<11>81  (
    .ADR0(DLX_EXinst_ALU_result[11]),
    .ADR1(CHOICE4405),
    .ADR2(N134884),
    .ADR3(N163286),
    .O(\N163286/GROM )
  );
  X_BUF \N163286/XUSED  (
    .I(\N163286/FROM ),
    .O(N163286)
  );
  X_BUF \N163286/YUSED  (
    .I(\N163286/GROM ),
    .O(CHOICE4407)
  );
  defparam reset_IBUF_14_684.INIT = 16'hAAAA;
  X_LUT4 reset_IBUF_14_684 (
    .ADR0(reset_IBUF),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\reset_IBUF_14/FROM )
  );
  defparam reset_IBUF_10_685.INIT = 16'hAAAA;
  X_LUT4 reset_IBUF_10_685 (
    .ADR0(reset_IBUF),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\reset_IBUF_14/GROM )
  );
  X_BUF \reset_IBUF_14/XUSED  (
    .I(\reset_IBUF_14/FROM ),
    .O(reset_IBUF_14)
  );
  X_BUF \reset_IBUF_14/YUSED  (
    .I(\reset_IBUF_14/GROM ),
    .O(reset_IBUF_10)
  );
  defparam reset_IBUF_13_686.INIT = 16'hAAAA;
  X_LUT4 reset_IBUF_13_686 (
    .ADR0(reset_IBUF),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\reset_IBUF_13/FROM )
  );
  defparam reset_IBUF_11_687.INIT = 16'hAAAA;
  X_LUT4 reset_IBUF_11_687 (
    .ADR0(reset_IBUF),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\reset_IBUF_13/GROM )
  );
  X_BUF \reset_IBUF_13/XUSED  (
    .I(\reset_IBUF_13/FROM ),
    .O(reset_IBUF_13)
  );
  X_BUF \reset_IBUF_13/YUSED  (
    .I(\reset_IBUF_13/GROM ),
    .O(reset_IBUF_11)
  );
  defparam reset_IBUF_9_688.INIT = 16'hAAAA;
  X_LUT4 reset_IBUF_9_688 (
    .ADR0(reset_IBUF),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\reset_IBUF_9/FROM )
  );
  defparam reset_IBUF_12_689.INIT = 16'hAAAA;
  X_LUT4 reset_IBUF_12_689 (
    .ADR0(reset_IBUF),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\reset_IBUF_9/GROM )
  );
  X_BUF \reset_IBUF_9/XUSED  (
    .I(\reset_IBUF_9/FROM ),
    .O(reset_IBUF_9)
  );
  X_BUF \reset_IBUF_9/YUSED  (
    .I(\reset_IBUF_9/GROM ),
    .O(reset_IBUF_12)
  );
  defparam \DLX_IDinst__n0146<0>39 .INIT = 16'h5088;
  X_LUT4 \DLX_IDinst__n0146<0>39  (
    .ADR0(DLX_IDinst_jtarget[22]),
    .ADR1(DLX_IDinst_EPC[0]),
    .ADR2(\DLX_IDinst_Cause_Reg[0] ),
    .ADR3(DLX_IDinst_jtarget[21]),
    .O(\DLX_IDinst_Cause_Reg<0>/GROM )
  );
  X_BUF \DLX_IDinst_Cause_Reg<0>/YUSED  (
    .I(\DLX_IDinst_Cause_Reg<0>/GROM ),
    .O(CHOICE3249)
  );
  defparam \DLX_IDinst__n0146<1>36_SW0 .INIT = 16'hCF77;
  X_LUT4 \DLX_IDinst__n0146<1>36_SW0  (
    .ADR0(DLX_IDinst_EPC[1]),
    .ADR1(DLX_IDinst_jtarget[22]),
    .ADR2(\DLX_IDinst_Cause_Reg[1] ),
    .ADR3(DLX_IDinst_jtarget[21]),
    .O(\DLX_IDinst_Cause_Reg<1>/FROM )
  );
  defparam \DLX_IDinst__n0146<1>36 .INIT = 16'h8F88;
  X_LUT4 \DLX_IDinst__n0146<1>36  (
    .ADR0(\DLX_IDinst_regA_eff[1] ),
    .ADR1(N134590),
    .ADR2(N163614),
    .ADR3(DLX_IDinst_N107105),
    .O(\DLX_IDinst_Cause_Reg<1>/GROM )
  );
  X_BUF \DLX_IDinst_Cause_Reg<1>/XUSED  (
    .I(\DLX_IDinst_Cause_Reg<1>/FROM ),
    .O(N163614)
  );
  X_BUF \DLX_IDinst_Cause_Reg<1>/YUSED  (
    .I(\DLX_IDinst_Cause_Reg<1>/GROM ),
    .O(CHOICE2903)
  );
  defparam \DLX_IDinst__n0146<2>36_SW0 .INIT = 16'hA7F7;
  X_LUT4 \DLX_IDinst__n0146<2>36_SW0  (
    .ADR0(DLX_IDinst_jtarget[22]),
    .ADR1(DLX_IDinst_EPC[2]),
    .ADR2(DLX_IDinst_jtarget[21]),
    .ADR3(\DLX_IDinst_Cause_Reg[2] ),
    .O(\DLX_IDinst_Cause_Reg<2>/FROM )
  );
  defparam \DLX_IDinst__n0146<2>36 .INIT = 16'hC0EA;
  X_LUT4 \DLX_IDinst__n0146<2>36  (
    .ADR0(DLX_IDinst_N107105),
    .ADR1(N134590),
    .ADR2(\DLX_IDinst_regA_eff[2] ),
    .ADR3(N163720),
    .O(\DLX_IDinst_Cause_Reg<2>/GROM )
  );
  X_BUF \DLX_IDinst_Cause_Reg<2>/XUSED  (
    .I(\DLX_IDinst_Cause_Reg<2>/FROM ),
    .O(N163720)
  );
  X_BUF \DLX_IDinst_Cause_Reg<2>/YUSED  (
    .I(\DLX_IDinst_Cause_Reg<2>/GROM ),
    .O(CHOICE2888)
  );
  defparam \DLX_IDinst__n0146<3>36_SW0 .INIT = 16'hD3DF;
  X_LUT4 \DLX_IDinst__n0146<3>36_SW0  (
    .ADR0(\DLX_IDinst_Cause_Reg[3] ),
    .ADR1(DLX_IDinst_jtarget[22]),
    .ADR2(DLX_IDinst_jtarget[21]),
    .ADR3(DLX_IDinst_EPC[3]),
    .O(\DLX_IDinst_Cause_Reg<3>/FROM )
  );
  defparam \DLX_IDinst__n0146<3>36 .INIT = 16'hC0EA;
  X_LUT4 \DLX_IDinst__n0146<3>36  (
    .ADR0(DLX_IDinst_N107105),
    .ADR1(N134590),
    .ADR2(\DLX_IDinst_regA_eff[3] ),
    .ADR3(N163437),
    .O(\DLX_IDinst_Cause_Reg<3>/GROM )
  );
  X_BUF \DLX_IDinst_Cause_Reg<3>/XUSED  (
    .I(\DLX_IDinst_Cause_Reg<3>/FROM ),
    .O(N163437)
  );
  X_BUF \DLX_IDinst_Cause_Reg<3>/YUSED  (
    .I(\DLX_IDinst_Cause_Reg<3>/GROM ),
    .O(CHOICE2483)
  );
  defparam \DLX_IDinst__n0146<4>36_SW0 .INIT = 16'h9DBF;
  X_LUT4 \DLX_IDinst__n0146<4>36_SW0  (
    .ADR0(DLX_IDinst_jtarget[21]),
    .ADR1(DLX_IDinst_jtarget[22]),
    .ADR2(DLX_IDinst_EPC[4]),
    .ADR3(\DLX_IDinst_Cause_Reg[4] ),
    .O(\DLX_IDinst_Cause_Reg<4>/FROM )
  );
  defparam \DLX_IDinst__n0146<4>36 .INIT = 16'hA0EC;
  X_LUT4 \DLX_IDinst__n0146<4>36  (
    .ADR0(N134590),
    .ADR1(DLX_IDinst_N107105),
    .ADR2(\DLX_IDinst_regA_eff[4] ),
    .ADR3(N163334),
    .O(\DLX_IDinst_Cause_Reg<4>/GROM )
  );
  X_BUF \DLX_IDinst_Cause_Reg<4>/XUSED  (
    .I(\DLX_IDinst_Cause_Reg<4>/FROM ),
    .O(N163334)
  );
  X_BUF \DLX_IDinst_Cause_Reg<4>/YUSED  (
    .I(\DLX_IDinst_Cause_Reg<4>/GROM ),
    .O(CHOICE2498)
  );
  defparam \DLX_IDinst__n0146<5>36_SW0 .INIT = 16'hC7F7;
  X_LUT4 \DLX_IDinst__n0146<5>36_SW0  (
    .ADR0(\DLX_IDinst_Cause_Reg[5] ),
    .ADR1(DLX_IDinst_jtarget[21]),
    .ADR2(DLX_IDinst_jtarget[22]),
    .ADR3(DLX_IDinst_EPC[5]),
    .O(\DLX_IDinst_Cause_Reg<5>/FROM )
  );
  defparam \DLX_IDinst__n0146<5>36 .INIT = 16'h88F8;
  X_LUT4 \DLX_IDinst__n0146<5>36  (
    .ADR0(\DLX_IDinst_regA_eff[5] ),
    .ADR1(N134590),
    .ADR2(DLX_IDinst_N107105),
    .ADR3(N163365),
    .O(\DLX_IDinst_Cause_Reg<5>/GROM )
  );
  X_BUF \DLX_IDinst_Cause_Reg<5>/XUSED  (
    .I(\DLX_IDinst_Cause_Reg<5>/FROM ),
    .O(N163365)
  );
  X_BUF \DLX_IDinst_Cause_Reg<5>/YUSED  (
    .I(\DLX_IDinst_Cause_Reg<5>/GROM ),
    .O(CHOICE2513)
  );
  defparam DLX_IDinst_RegFile_18_19_690.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_18_19_690 (
    .I(DLX_IDinst_WB_data_eff[19]),
    .CE(DLX_IDinst__n0586),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_18_19)
  );
  defparam \DLX_IDinst__n0146<7>36_SW0 .INIT = 16'hB5BF;
  X_LUT4 \DLX_IDinst__n0146<7>36_SW0  (
    .ADR0(DLX_IDinst_jtarget[22]),
    .ADR1(\DLX_IDinst_Cause_Reg[7] ),
    .ADR2(DLX_IDinst_jtarget[21]),
    .ADR3(DLX_IDinst_EPC[7]),
    .O(\DLX_IDinst_Cause_Reg<7>/FROM )
  );
  defparam \DLX_IDinst__n0146<7>36 .INIT = 16'h88F8;
  X_LUT4 \DLX_IDinst__n0146<7>36  (
    .ADR0(N134590),
    .ADR1(\DLX_IDinst_regA_eff[7] ),
    .ADR2(DLX_IDinst_N107105),
    .ADR3(N163712),
    .O(\DLX_IDinst_Cause_Reg<7>/GROM )
  );
  X_BUF \DLX_IDinst_Cause_Reg<7>/XUSED  (
    .I(\DLX_IDinst_Cause_Reg<7>/FROM ),
    .O(N163712)
  );
  X_BUF \DLX_IDinst_Cause_Reg<7>/YUSED  (
    .I(\DLX_IDinst_Cause_Reg<7>/GROM ),
    .O(CHOICE2528)
  );
  defparam \DLX_IDinst__n0146<8>36_SW0 .INIT = 16'hA7F7;
  X_LUT4 \DLX_IDinst__n0146<8>36_SW0  (
    .ADR0(DLX_IDinst_jtarget[21]),
    .ADR1(\DLX_IDinst_Cause_Reg[8] ),
    .ADR2(DLX_IDinst_jtarget[22]),
    .ADR3(DLX_IDinst_EPC[8]),
    .O(\DLX_IDinst_Cause_Reg<8>/FROM )
  );
  defparam \DLX_IDinst__n0146<8>36 .INIT = 16'h88F8;
  X_LUT4 \DLX_IDinst__n0146<8>36  (
    .ADR0(N134590),
    .ADR1(\DLX_IDinst_regA_eff[8] ),
    .ADR2(DLX_IDinst_N107105),
    .ADR3(N163403),
    .O(\DLX_IDinst_Cause_Reg<8>/GROM )
  );
  X_BUF \DLX_IDinst_Cause_Reg<8>/XUSED  (
    .I(\DLX_IDinst_Cause_Reg<8>/FROM ),
    .O(N163403)
  );
  X_BUF \DLX_IDinst_Cause_Reg<8>/YUSED  (
    .I(\DLX_IDinst_Cause_Reg<8>/GROM ),
    .O(CHOICE2543)
  );
  defparam \DLX_IDinst__n0146<9>36_SW0 .INIT = 16'hAF77;
  X_LUT4 \DLX_IDinst__n0146<9>36_SW0  (
    .ADR0(DLX_IDinst_jtarget[22]),
    .ADR1(DLX_IDinst_EPC[9]),
    .ADR2(\DLX_IDinst_Cause_Reg[9] ),
    .ADR3(DLX_IDinst_jtarget[21]),
    .O(\DLX_IDinst_Cause_Reg<9>/FROM )
  );
  defparam \DLX_IDinst__n0146<9>36 .INIT = 16'h88F8;
  X_LUT4 \DLX_IDinst__n0146<9>36  (
    .ADR0(N134590),
    .ADR1(\DLX_IDinst_regA_eff[9] ),
    .ADR2(DLX_IDinst_N107105),
    .ADR3(N163570),
    .O(\DLX_IDinst_Cause_Reg<9>/GROM )
  );
  X_BUF \DLX_IDinst_Cause_Reg<9>/XUSED  (
    .I(\DLX_IDinst_Cause_Reg<9>/FROM ),
    .O(N163570)
  );
  X_BUF \DLX_IDinst_Cause_Reg<9>/YUSED  (
    .I(\DLX_IDinst_Cause_Reg<9>/GROM ),
    .O(CHOICE2558)
  );
  defparam \DLX_EXinst__n0007<8>217 .INIT = 16'h4448;
  X_LUT4 \DLX_EXinst__n0007<8>217  (
    .ADR0(DLX_IDinst_IR_opcode_field[1]),
    .ADR1(DLX_EXinst_N76011),
    .ADR2(DLX_IDinst_reg_out_A[8]),
    .ADR3(DLX_IDinst_IR_opcode_field[0]),
    .O(\CHOICE5181/FROM )
  );
  defparam \DLX_EXinst__n0007<22>92_SW0 .INIT = 16'h4448;
  X_LUT4 \DLX_EXinst__n0007<22>92_SW0  (
    .ADR0(DLX_IDinst_IR_opcode_field[1]),
    .ADR1(DLX_EXinst_N76011),
    .ADR2(DLX_IDinst_reg_out_A[22]),
    .ADR3(DLX_IDinst_IR_opcode_field[0]),
    .O(\CHOICE5181/GROM )
  );
  X_BUF \CHOICE5181/XUSED  (
    .I(\CHOICE5181/FROM ),
    .O(CHOICE5181)
  );
  X_BUF \CHOICE5181/YUSED  (
    .I(\CHOICE5181/GROM ),
    .O(N163282)
  );
  defparam DLX_IDinst__n0428117.INIT = 16'h0C04;
  X_LUT4 DLX_IDinst__n0428117 (
    .ADR0(DLX_IDinst_IR_latched[27]),
    .ADR1(DLX_IDinst_N108476),
    .ADR2(DLX_IDinst_IR_latched[28]),
    .ADR3(DLX_IDinst_IR_latched[26]),
    .O(\CHOICE1994/FROM )
  );
  defparam DLX_IDinst__n0151115.INIT = 16'h2000;
  X_LUT4 DLX_IDinst__n0151115 (
    .ADR0(DLX_IDinst_IR_latched[26]),
    .ADR1(DLX_IDinst_IR_latched[28]),
    .ADR2(DLX_IDinst_N108443),
    .ADR3(DLX_IDinst_IR_latched[27]),
    .O(\CHOICE1994/GROM )
  );
  X_BUF \CHOICE1994/XUSED  (
    .I(\CHOICE1994/FROM ),
    .O(CHOICE1994)
  );
  X_BUF \CHOICE1994/YUSED  (
    .I(\CHOICE1994/GROM ),
    .O(CHOICE3343)
  );
  defparam DLX_IDinst__n0151119.INIT = 16'hFF0E;
  X_LUT4 DLX_IDinst__n0151119 (
    .ADR0(CHOICE3337),
    .ADR1(CHOICE3323),
    .ADR2(DLX_IDinst__n0453),
    .ADR3(CHOICE3343),
    .O(\DLX_IDinst_delay_slot/FROM )
  );
  defparam DLX_IDinst__n0151130.INIT = 16'h5500;
  X_LUT4 DLX_IDinst__n0151130 (
    .ADR0(DLX_IDinst__n0387),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(CHOICE3344),
    .O(N146881)
  );
  X_BUF \DLX_IDinst_delay_slot/XUSED  (
    .I(\DLX_IDinst_delay_slot/FROM ),
    .O(CHOICE3344)
  );
  defparam \DLX_EXinst__n0007<18>136_SW0 .INIT = 16'h04C8;
  X_LUT4 \DLX_EXinst__n0007<18>136_SW0  (
    .ADR0(DLX_IDinst_reg_out_A[18]),
    .ADR1(DLX_EXinst_N76011),
    .ADR2(DLX_IDinst_IR_opcode_field[0]),
    .ADR3(DLX_IDinst_IR_opcode_field[1]),
    .O(\N163420/FROM )
  );
  defparam \DLX_EXinst__n0007<23>92_SW0 .INIT = 16'h2228;
  X_LUT4 \DLX_EXinst__n0007<23>92_SW0  (
    .ADR0(DLX_EXinst_N76011),
    .ADR1(DLX_IDinst_IR_opcode_field[1]),
    .ADR2(DLX_IDinst_reg_out_A[23]),
    .ADR3(DLX_IDinst_IR_opcode_field[0]),
    .O(\N163420/GROM )
  );
  X_BUF \N163420/XUSED  (
    .I(\N163420/FROM ),
    .O(N163420)
  );
  X_BUF \N163420/YUSED  (
    .I(\N163420/GROM ),
    .O(N163460)
  );
  defparam DLX_IDinst__n0137116.INIT = 16'hC4CC;
  X_LUT4 DLX_IDinst__n0137116 (
    .ADR0(DLX_IDinst_N108503),
    .ADR1(CHOICE3526),
    .ADR2(DLX_IDinst_IR_latched[30]),
    .ADR3(DLX_IDinst_IR_latched[27]),
    .O(\DLX_IDinst_reg_dst/FROM )
  );
  defparam DLX_IDinst__n0137152.INIT = 16'hFFFA;
  X_LUT4 DLX_IDinst__n0137152 (
    .ADR0(DLX_IDinst_N108456),
    .ADR1(VCC),
    .ADR2(N163190),
    .ADR3(CHOICE3527),
    .O(N147993)
  );
  X_BUF \DLX_IDinst_reg_dst/XUSED  (
    .I(\DLX_IDinst_reg_dst/FROM ),
    .O(CHOICE3527)
  );
  defparam DLX_IDinst__n0138131.INIT = 16'hECA0;
  X_LUT4 DLX_IDinst__n0138131 (
    .ADR0(DLX_IDinst_N107405),
    .ADR1(DLX_IDinst_N107572),
    .ADR2(DLX_IDinst__n0629[1]),
    .ADR3(DLX_IDinst_N108152),
    .O(\CHOICE3558/FROM )
  );
  defparam DLX_IDinst__n0138169_SW0.INIT = 16'hFFA0;
  X_LUT4 DLX_IDinst__n0138169_SW0 (
    .ADR0(CHOICE3553),
    .ADR1(VCC),
    .ADR2(DLX_IDinst__n0163),
    .ADR3(CHOICE3558),
    .O(\CHOICE3558/GROM )
  );
  X_BUF \CHOICE3558/XUSED  (
    .I(\CHOICE3558/FROM ),
    .O(CHOICE3558)
  );
  X_BUF \CHOICE3558/YUSED  (
    .I(\CHOICE3558/GROM ),
    .O(N163120)
  );
  defparam DLX_IDinst__n0138160.INIT = 16'h0400;
  X_LUT4 DLX_IDinst__n0138160 (
    .ADR0(DLX_IDinst__n0453),
    .ADR1(DLX_IDinst_IR_latched[30]),
    .ADR2(DLX_IDinst_IR_latched[27]),
    .ADR3(DLX_IDinst_N108503),
    .O(\DLX_IDinst_reg_write/FROM )
  );
  defparam DLX_IDinst__n0138169.INIT = 16'hFFEA;
  X_LUT4 DLX_IDinst__n0138169 (
    .ADR0(DLX_IDinst_N108456),
    .ADR1(DLX_IDinst_N107223),
    .ADR2(N163120),
    .ADR3(CHOICE3565),
    .O(N148197)
  );
  X_BUF \DLX_IDinst_reg_write/XUSED  (
    .I(\DLX_IDinst_reg_write/FROM ),
    .O(CHOICE3565)
  );
  defparam DLX_IFinst_IR_curr_1.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_1 (
    .I(IR[1]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[1])
  );
  defparam DLX_IFinst_IR_curr_2.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_2 (
    .I(IR[2]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[2])
  );
  defparam DLX_IDinst_RegFile_26_27_691.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_26_27_691 (
    .I(DLX_IDinst_WB_data_eff[27]),
    .CE(DLX_IDinst__n0602),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_26_27)
  );
  defparam DLX_IFinst_IR_curr_3.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_3 (
    .I(IR[3]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[3])
  );
  defparam DLX_IFinst_IR_curr_5.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_5 (
    .I(IR[5]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[5])
  );
  defparam DLX_IFinst_IR_curr_8.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_8 (
    .I(IR[8]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[8])
  );
  defparam DLX_IFinst_IR_curr_9.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_9 (
    .I(IR[9]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[9])
  );
  defparam DLX_IDinst__n0177116.INIT = 16'h0001;
  X_LUT4 DLX_IDinst__n0177116 (
    .ADR0(\DLX_IDinst_regA_eff[10] ),
    .ADR1(\DLX_IDinst_regA_eff[9] ),
    .ADR2(\DLX_IDinst_regA_eff[11] ),
    .ADR3(\DLX_IDinst_regA_eff[12] ),
    .O(\CHOICE4224/FROM )
  );
  defparam DLX_IDinst__n0177117.INIT = 16'hCC00;
  X_LUT4 DLX_IDinst__n0177117 (
    .ADR0(VCC),
    .ADR1(CHOICE4217),
    .ADR2(VCC),
    .ADR3(CHOICE4224),
    .O(\CHOICE4224/GROM )
  );
  X_BUF \CHOICE4224/XUSED  (
    .I(\CHOICE4224/FROM ),
    .O(CHOICE4224)
  );
  X_BUF \CHOICE4224/YUSED  (
    .I(\CHOICE4224/GROM ),
    .O(CHOICE4225)
  );
  defparam DLX_IDinst__n0177207.INIT = 16'hF000;
  X_LUT4 DLX_IDinst__n0177207 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(CHOICE4255),
    .ADR3(CHOICE4248),
    .O(\CHOICE4256/FROM )
  );
  defparam DLX_IDinst__n0177234_SW0.INIT = 16'hDFFF;
  X_LUT4 DLX_IDinst__n0177234_SW0 (
    .ADR0(CHOICE4240),
    .ADR1(\DLX_IDinst_regA_eff[30] ),
    .ADR2(CHOICE4233),
    .ADR3(CHOICE4256),
    .O(\CHOICE4256/GROM )
  );
  X_BUF \CHOICE4256/XUSED  (
    .I(\CHOICE4256/FROM ),
    .O(CHOICE4256)
  );
  X_BUF \CHOICE4256/YUSED  (
    .I(\CHOICE4256/GROM ),
    .O(N163546)
  );
  defparam DLX_IDinst__n0177234.INIT = 16'h1000;
  X_LUT4 DLX_IDinst__n0177234 (
    .ADR0(\DLX_IDinst_regA_eff[29] ),
    .ADR1(N163546),
    .ADR2(CHOICE4209),
    .ADR3(CHOICE4225),
    .O(\DLX_IDinst_zflag/FROM )
  );
  defparam DLX_IDinst_Ker10825731.INIT = 16'h0330;
  X_LUT4 DLX_IDinst_Ker10825731 (
    .ADR0(VCC),
    .ADR1(DLX_IFinst_IR_latched[30]),
    .ADR2(DLX_IFinst_IR_latched[26]),
    .ADR3(DLX_IDinst_zflag),
    .O(\DLX_IDinst_zflag/GROM )
  );
  X_BUF \DLX_IDinst_zflag/XUSED  (
    .I(\DLX_IDinst_zflag/FROM ),
    .O(DLX_IDinst_zflag)
  );
  X_BUF \DLX_IDinst_zflag/YUSED  (
    .I(\DLX_IDinst_zflag/GROM ),
    .O(CHOICE3293)
  );
  defparam DLX_IDinst__n0428118.INIT = 16'hEEEE;
  X_LUT4 DLX_IDinst__n0428118 (
    .ADR0(CHOICE1989),
    .ADR1(CHOICE1994),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\N138903/FROM )
  );
  defparam DLX_IDinst__n013747.INIT = 16'h040C;
  X_LUT4 DLX_IDinst__n013747 (
    .ADR0(DLX_IDinst_N108238),
    .ADR1(DLX_IDinst__n0166),
    .ADR2(N135079),
    .ADR3(N138903),
    .O(\N138903/GROM )
  );
  X_BUF \N138903/XUSED  (
    .I(\N138903/FROM ),
    .O(N138903)
  );
  X_BUF \N138903/YUSED  (
    .I(\N138903/GROM ),
    .O(CHOICE3515)
  );
  defparam DLX_IDinst_Ker1072211.INIT = 16'h090F;
  X_LUT4 DLX_IDinst_Ker1072211 (
    .ADR0(DLX_IDinst_IR_latched[27]),
    .ADR1(DLX_IDinst_IR_latched[30]),
    .ADR2(DLX_IDinst__n0453),
    .ADR3(DLX_IDinst_N108503),
    .O(\DLX_IDinst_N107223/FROM )
  );
  defparam DLX_IDinst__n0140_SW0.INIT = 16'h80FF;
  X_LUT4 DLX_IDinst__n0140_SW0 (
    .ADR0(DLX_IDinst_IR_latched[27]),
    .ADR1(DLX_IDinst_IR_latched[26]),
    .ADR2(DLX_IDinst_N108165),
    .ADR3(DLX_IDinst_N107223),
    .O(\DLX_IDinst_N107223/GROM )
  );
  X_BUF \DLX_IDinst_N107223/XUSED  (
    .I(\DLX_IDinst_N107223/FROM ),
    .O(DLX_IDinst_N107223)
  );
  X_BUF \DLX_IDinst_N107223/YUSED  (
    .I(\DLX_IDinst_N107223/GROM ),
    .O(N127137)
  );
  defparam DLX_IDinst_RegFile_19_11_692.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_19_11_692 (
    .I(DLX_IDinst_WB_data_eff[11]),
    .CE(DLX_IDinst__n0588),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_19_11)
  );
  defparam \DLX_EXinst__n0007<0>390_SW0 .INIT = 16'hFEFA;
  X_LUT4 \DLX_EXinst__n0007<0>390_SW0  (
    .ADR0(CHOICE5908),
    .ADR1(CHOICE5901),
    .ADR2(N164591),
    .ADR3(DLX_IDinst_reg_out_A[0]),
    .O(\N163416/FROM )
  );
  defparam \DLX_EXinst__n0007<0>390 .INIT = 16'hAAA8;
  X_LUT4 \DLX_EXinst__n0007<0>390  (
    .ADR0(DLX_EXinst__n0036),
    .ADR1(CHOICE5896),
    .ADR2(CHOICE5871),
    .ADR3(N163416),
    .O(\N163416/GROM )
  );
  X_BUF \N163416/XUSED  (
    .I(\N163416/FROM ),
    .O(N163416)
  );
  X_BUF \N163416/YUSED  (
    .I(\N163416/GROM ),
    .O(CHOICE5945)
  );
  defparam \DLX_IFinst__n0001<10>_SW0 .INIT = 16'h0F55;
  X_LUT4 \DLX_IFinst__n0001<10>_SW0  (
    .ADR0(DLX_IFinst__n0015[10]),
    .ADR1(VCC),
    .ADR2(DLX_IFinst_PC[10]),
    .ADR3(DLX_IFinst__n0000),
    .O(\DLX_IFinst_NPC<10>/FROM )
  );
  defparam \DLX_IFinst__n0001<10> .INIT = 16'h88BB;
  X_LUT4 \DLX_IFinst__n0001<10>  (
    .ADR0(DLX_IDinst_branch_address[10]),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(VCC),
    .ADR3(N129431),
    .O(\DLX_IFinst_NPC<10>/GROM )
  );
  X_BUF \DLX_IFinst_NPC<10>/XUSED  (
    .I(\DLX_IFinst_NPC<10>/FROM ),
    .O(N129431)
  );
  X_BUF \DLX_IFinst_NPC<10>/YUSED  (
    .I(\DLX_IFinst_NPC<10>/GROM ),
    .O(DLX_IFinst__n0001[10])
  );
  defparam DLX_IDinst_Ker1083031.INIT = 16'hAA80;
  X_LUT4 DLX_IDinst_Ker1083031 (
    .ADR0(DLX_IDinst_N107033),
    .ADR1(DLX_IDinst_N108465),
    .ADR2(DLX_IDinst_N108152),
    .ADR3(DLX_IDinst_N107405),
    .O(\DLX_IDinst_N108305/FROM )
  );
  defparam \DLX_IDinst__n0114<26>6 .INIT = 16'hEAC0;
  X_LUT4 \DLX_IDinst__n0114<26>6  (
    .ADR0(DLX_IDinst_branch_address[26]),
    .ADR1(DLX_IDinst_EPC[26]),
    .ADR2(DLX_IDinst__n0098),
    .ADR3(DLX_IDinst_N108305),
    .O(\DLX_IDinst_N108305/GROM )
  );
  X_BUF \DLX_IDinst_N108305/XUSED  (
    .I(\DLX_IDinst_N108305/FROM ),
    .O(DLX_IDinst_N108305)
  );
  X_BUF \DLX_IDinst_N108305/YUSED  (
    .I(\DLX_IDinst_N108305/GROM ),
    .O(CHOICE2430)
  );
  defparam \DLX_EXinst__n0007<0>471_SW1 .INIT = 16'h7F57;
  X_LUT4 \DLX_EXinst__n0007<0>471_SW1  (
    .ADR0(DLX_IDinst_IR_opcode_field[1]),
    .ADR1(DLX_EXinst_Mcompar__n0065_inst_cy_196),
    .ADR2(\DLX_IDinst_Imm[31] ),
    .ADR3(DLX_IDinst_reg_out_A[31]),
    .O(\N164614/FROM )
  );
  defparam \DLX_EXinst__n0007<0>471_SW0 .INIT = 16'h2FBF;
  X_LUT4 \DLX_EXinst__n0007<0>471_SW0  (
    .ADR0(\DLX_IDinst_Imm[31] ),
    .ADR1(DLX_EXinst_Mcompar__n0063_inst_cy_164),
    .ADR2(DLX_IDinst_IR_opcode_field[1]),
    .ADR3(DLX_IDinst_reg_out_A[31]),
    .O(\N164614/GROM )
  );
  X_BUF \N164614/XUSED  (
    .I(\N164614/FROM ),
    .O(N164614)
  );
  X_BUF \N164614/YUSED  (
    .I(\N164614/GROM ),
    .O(N164612)
  );
  defparam DLX_IDinst_Ker1082421.INIT = 16'h0011;
  X_LUT4 DLX_IDinst_Ker1082421 (
    .ADR0(DLX_IDinst_jtarget[24]),
    .ADR1(DLX_IDinst_jtarget[23]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_jtarget[25]),
    .O(\DLX_IDinst_N108244/FROM )
  );
  defparam DLX_IDinst__n03821.INIT = 16'h1100;
  X_LUT4 DLX_IDinst__n03821 (
    .ADR0(DLX_IDinst_jtarget[22]),
    .ADR1(DLX_IDinst_jtarget[21]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_N108244),
    .O(\DLX_IDinst_N108244/GROM )
  );
  X_BUF \DLX_IDinst_N108244/XUSED  (
    .I(\DLX_IDinst_N108244/FROM ),
    .O(DLX_IDinst_N108244)
  );
  X_BUF \DLX_IDinst_N108244/YUSED  (
    .I(\DLX_IDinst_N108244/GROM ),
    .O(DLX_IDinst__n0382)
  );
  defparam DLX_IDinst_Ker1074501.INIT = 16'hFAFA;
  X_LUT4 DLX_IDinst_Ker1074501 (
    .ADR0(DLX_IDinst_slot_num_FFd1),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_slot_num_FFd3),
    .ADR3(VCC),
    .O(\DLX_IDinst_N107452/FROM )
  );
  defparam DLX_IDinst__n03761.INIT = 16'hF0D0;
  X_LUT4 DLX_IDinst__n03761 (
    .ADR0(DLX_IDinst_slot_num_FFd2),
    .ADR1(DLX_IDinst_slot_num_FFd4),
    .ADR2(DLX_IDinst_delay_slot),
    .ADR3(DLX_IDinst_N107452),
    .O(\DLX_IDinst_N107452/GROM )
  );
  X_BUF \DLX_IDinst_N107452/XUSED  (
    .I(\DLX_IDinst_N107452/FROM ),
    .O(DLX_IDinst_N107452)
  );
  X_BUF \DLX_IDinst_N107452/YUSED  (
    .I(\DLX_IDinst_N107452/GROM ),
    .O(DLX_IDinst__n0376)
  );
  defparam DLX_IDinst_Ker1082191.INIT = 16'h0300;
  X_LUT4 DLX_IDinst_Ker1082191 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_IR_latched[27]),
    .ADR2(DLX_IDinst_IR_latched[30]),
    .ADR3(DLX_IDinst_IR_latched[28]),
    .O(\DLX_IDinst_N108221/FROM )
  );
  defparam DLX_IDinst__n01061.INIT = 16'h0100;
  X_LUT4 DLX_IDinst__n01061 (
    .ADR0(DLX_IDinst_IR_latched[29]),
    .ADR1(DLX_IDinst_IR_latched[26]),
    .ADR2(DLX_IDinst_IR_latched[31]),
    .ADR3(DLX_IDinst_N108221),
    .O(\DLX_IDinst_N108221/GROM )
  );
  X_BUF \DLX_IDinst_N108221/XUSED  (
    .I(\DLX_IDinst_N108221/FROM ),
    .O(DLX_IDinst_N108221)
  );
  X_BUF \DLX_IDinst_N108221/YUSED  (
    .I(\DLX_IDinst_N108221/GROM ),
    .O(DLX_IDinst__n0106)
  );
  defparam DLX_IDinst_Ker1081631.INIT = 16'h04C4;
  X_LUT4 DLX_IDinst_Ker1081631 (
    .ADR0(DLX_IDinst_current_IR[28]),
    .ADR1(DLX_IDinst_N108443),
    .ADR2(DLX_EXinst__n0144),
    .ADR3(DLX_IFinst_IR_latched[28]),
    .O(\DLX_IDinst_N108165/FROM )
  );
  defparam DLX_IDinst_N1070331.INIT = 16'hF9FF;
  X_LUT4 DLX_IDinst_N1070331 (
    .ADR0(DLX_IDinst_IR_latched[30]),
    .ADR1(DLX_IDinst_IR_latched[27]),
    .ADR2(DLX_IDinst_IR_latched[26]),
    .ADR3(DLX_IDinst_N108165),
    .O(\DLX_IDinst_N108165/GROM )
  );
  X_BUF \DLX_IDinst_N108165/XUSED  (
    .I(\DLX_IDinst_N108165/FROM ),
    .O(DLX_IDinst_N108165)
  );
  X_BUF \DLX_IDinst_N108165/YUSED  (
    .I(\DLX_IDinst_N108165/GROM ),
    .O(DLX_IDinst_N107033)
  );
  defparam DLX_IDinst_Ker1082361.INIT = 16'h0022;
  X_LUT4 DLX_IDinst_Ker1082361 (
    .ADR0(DLX_IDinst_IR_opcode_field[3]),
    .ADR1(DLX_IDinst_IR_opcode_field[1]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_IR_opcode_field[5]),
    .O(\DLX_IDinst_N108238/FROM )
  );
  defparam DLX_IDinst__n04331.INIT = 16'hFCCC;
  X_LUT4 DLX_IDinst__n04331 (
    .ADR0(VCC),
    .ADR1(N135079),
    .ADR2(N137212),
    .ADR3(DLX_IDinst_N108238),
    .O(\DLX_IDinst_N108238/GROM )
  );
  X_BUF \DLX_IDinst_N108238/XUSED  (
    .I(\DLX_IDinst_N108238/FROM ),
    .O(DLX_IDinst_N108238)
  );
  X_BUF \DLX_IDinst_N108238/YUSED  (
    .I(\DLX_IDinst_N108238/GROM ),
    .O(DLX_IDinst__n0433)
  );
  defparam DLX_IDinst_Ker108257139_SW0.INIT = 16'h3122;
  X_LUT4 DLX_IDinst_Ker108257139_SW0 (
    .ADR0(DLX_IFinst_IR_latched[30]),
    .ADR1(DLX_IFinst_IR_latched[28]),
    .ADR2(DLX_IFinst_IR_latched[26]),
    .ADR3(DLX_IFinst_IR_latched[27]),
    .O(\N163258/GROM )
  );
  X_BUF \N163258/YUSED  (
    .I(\N163258/GROM ),
    .O(N163258)
  );
  defparam DLX_IDinst_Ker1076211.INIT = 16'hAAFF;
  X_LUT4 DLX_IDinst_Ker1076211 (
    .ADR0(DLX_IDinst_CLI),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(INT_IBUF),
    .O(\DLX_IDinst_N107623/FROM )
  );
  defparam \DLX_IDinst_slot_num_FFd2-In17 .INIT = 16'h88FA;
  X_LUT4 \DLX_IDinst_slot_num_FFd2-In17  (
    .ADR0(N163222),
    .ADR1(N146700),
    .ADR2(DLX_IDinst_slot_num_FFd2),
    .ADR3(DLX_IDinst_N107623),
    .O(\DLX_IDinst_N107623/GROM )
  );
  X_BUF \DLX_IDinst_N107623/XUSED  (
    .I(\DLX_IDinst_N107623/FROM ),
    .O(DLX_IDinst_N107623)
  );
  X_BUF \DLX_IDinst_N107623/YUSED  (
    .I(\DLX_IDinst_N107623/GROM ),
    .O(CHOICE2128)
  );
  defparam DLX_IDinst_Ker1085011.INIT = 16'h2222;
  X_LUT4 DLX_IDinst_Ker1085011 (
    .ADR0(DLX_IDinst_N108165),
    .ADR1(DLX_IDinst_IR_latched[26]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IDinst_N108503/FROM )
  );
  defparam DLX_IDinst_Ker10757410.INIT = 16'hDCCC;
  X_LUT4 DLX_IDinst_Ker10757410 (
    .ADR0(DLX_IDinst__n0453),
    .ADR1(DLX_IDinst_Ker1084541_1),
    .ADR2(DLX_IDinst_IR_latched[27]),
    .ADR3(DLX_IDinst_N108503),
    .O(\DLX_IDinst_N108503/GROM )
  );
  X_BUF \DLX_IDinst_N108503/XUSED  (
    .I(\DLX_IDinst_N108503/FROM ),
    .O(DLX_IDinst_N108503)
  );
  X_BUF \DLX_IDinst_N108503/YUSED  (
    .I(\DLX_IDinst_N108503/GROM ),
    .O(CHOICE1689)
  );
  defparam DLX_IDinst_Ker1082621.INIT = 16'h0010;
  X_LUT4 DLX_IDinst_Ker1082621 (
    .ADR0(DLX_IDinst_IR_latched[29]),
    .ADR1(DLX_IDinst_IR_latched[28]),
    .ADR2(DLX_IDinst_IR_latched[30]),
    .ADR3(DLX_IDinst_IR_latched[27]),
    .O(\DLX_IDinst_N108264/FROM )
  );
  defparam DLX_IDinst_Ker10735446_SW1.INIT = 16'h8800;
  X_LUT4 DLX_IDinst_Ker10735446_SW1 (
    .ADR0(DLX_IDinst_IR_latched[26]),
    .ADR1(DLX_IDinst_IR_latched[31]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_N108264),
    .O(\DLX_IDinst_N108264/GROM )
  );
  X_BUF \DLX_IDinst_N108264/XUSED  (
    .I(\DLX_IDinst_N108264/FROM ),
    .O(DLX_IDinst_N108264)
  );
  X_BUF \DLX_IDinst_N108264/YUSED  (
    .I(\DLX_IDinst_N108264/GROM ),
    .O(N163838)
  );
  defparam DLX_IDinst_Ker1082471.INIT = 16'h004C;
  X_LUT4 DLX_IDinst_Ker1082471 (
    .ADR0(DLX_IDinst_delay_slot),
    .ADR1(FREEZE_IBUF),
    .ADR2(DLX_IDinst_N107452),
    .ADR3(DLX_IDinst_intr_slot),
    .O(\DLX_IDinst_N108249/FROM )
  );
  defparam DLX_IDinst__n0149112.INIT = 16'hF000;
  X_LUT4 DLX_IDinst__n0149112 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IDinst__n0387),
    .ADR3(DLX_IDinst_N108249),
    .O(\DLX_IDinst_N108249/GROM )
  );
  X_BUF \DLX_IDinst_N108249/XUSED  (
    .I(\DLX_IDinst_N108249/FROM ),
    .O(DLX_IDinst_N108249)
  );
  X_BUF \DLX_IDinst_N108249/YUSED  (
    .I(\DLX_IDinst_N108249/GROM ),
    .O(CHOICE3495)
  );
  defparam DLX_IDinst_Ker1080981.INIT = 16'hFFFA;
  X_LUT4 DLX_IDinst_Ker1080981 (
    .ADR0(DLX_IDinst_counter[0]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_intr_slot),
    .ADR3(DLX_IDinst_counter[1]),
    .O(\DLX_IDinst_N108100/FROM )
  );
  defparam DLX_IDinst__n03911.INIT = 16'h0002;
  X_LUT4 DLX_IDinst__n03911 (
    .ADR0(DLX_IDinst_stall),
    .ADR1(DLX_IDinst_delay_slot),
    .ADR2(FREEZE_IBUF),
    .ADR3(DLX_IDinst_N108100),
    .O(\DLX_IDinst_N108100/GROM )
  );
  X_BUF \DLX_IDinst_N108100/XUSED  (
    .I(\DLX_IDinst_N108100/FROM ),
    .O(DLX_IDinst_N108100)
  );
  X_BUF \DLX_IDinst_N108100/YUSED  (
    .I(\DLX_IDinst_N108100/GROM ),
    .O(DLX_IDinst__n0391)
  );
  defparam DLX_IDinst_Ker1085151.INIT = 16'h0100;
  X_LUT4 DLX_IDinst_Ker1085151 (
    .ADR0(DLX_MEMinst_reg_dst_out[0]),
    .ADR1(DLX_MEMinst_reg_dst_out[2]),
    .ADR2(DLX_MEMinst_reg_dst_out[4]),
    .ADR3(DLX_MEMinst_reg_write_MEM),
    .O(\DLX_IDinst_N108517/FROM )
  );
  defparam DLX_IDinst__n05541.INIT = 16'h3000;
  X_LUT4 DLX_IDinst__n05541 (
    .ADR0(VCC),
    .ADR1(DLX_MEMinst_reg_dst_out[3]),
    .ADR2(DLX_MEMinst_reg_dst_out[1]),
    .ADR3(DLX_IDinst_N108517),
    .O(\DLX_IDinst_N108517/GROM )
  );
  X_BUF \DLX_IDinst_N108517/XUSED  (
    .I(\DLX_IDinst_N108517/FROM ),
    .O(DLX_IDinst_N108517)
  );
  X_BUF \DLX_IDinst_N108517/YUSED  (
    .I(\DLX_IDinst_N108517/GROM ),
    .O(DLX_IDinst__n0554)
  );
  defparam \DLX_IFinst__n0001<11>_SW0 .INIT = 16'h2727;
  X_LUT4 \DLX_IFinst__n0001<11>_SW0  (
    .ADR0(DLX_IFinst__n0000),
    .ADR1(DLX_IFinst_PC[11]),
    .ADR2(DLX_IFinst__n0015[11]),
    .ADR3(VCC),
    .O(\DLX_IFinst_NPC<11>/FROM )
  );
  defparam \DLX_IFinst__n0001<11> .INIT = 16'hA0AF;
  X_LUT4 \DLX_IFinst__n0001<11>  (
    .ADR0(DLX_IDinst_branch_address[11]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(N129379),
    .O(\DLX_IFinst_NPC<11>/GROM )
  );
  X_BUF \DLX_IFinst_NPC<11>/XUSED  (
    .I(\DLX_IFinst_NPC<11>/FROM ),
    .O(N129379)
  );
  X_BUF \DLX_IFinst_NPC<11>/YUSED  (
    .I(\DLX_IFinst_NPC<11>/GROM ),
    .O(DLX_IFinst__n0001[11])
  );
  defparam DLX_IDinst_Ker1085501.INIT = 16'h0008;
  X_LUT4 DLX_IDinst_Ker1085501 (
    .ADR0(DLX_MEMinst_reg_dst_out[4]),
    .ADR1(DLX_MEMinst_reg_write_MEM),
    .ADR2(DLX_MEMinst_reg_dst_out[0]),
    .ADR3(DLX_MEMinst_reg_dst_out[2]),
    .O(\DLX_IDinst_N108552/FROM )
  );
  defparam DLX_IDinst__n06021.INIT = 16'h8800;
  X_LUT4 DLX_IDinst__n06021 (
    .ADR0(DLX_MEMinst_reg_dst_out[3]),
    .ADR1(DLX_MEMinst_reg_dst_out[1]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_N108552),
    .O(\DLX_IDinst_N108552/GROM )
  );
  X_BUF \DLX_IDinst_N108552/XUSED  (
    .I(\DLX_IDinst_N108552/FROM ),
    .O(DLX_IDinst_N108552)
  );
  X_BUF \DLX_IDinst_N108552/YUSED  (
    .I(\DLX_IDinst_N108552/GROM ),
    .O(DLX_IDinst__n0602)
  );
  defparam \DLX_EXinst__n0007<1>241_SW0 .INIT = 16'h4555;
  X_LUT4 \DLX_EXinst__n0007<1>241_SW0  (
    .ADR0(CHOICE5747),
    .ADR1(DLX_EXinst_N72822),
    .ADR2(DLX_EXinst_N76268),
    .ADR3(\DLX_EXinst_Mshift__n0023_Sh[1] ),
    .O(\N164200/FROM )
  );
  defparam \DLX_EXinst__n0007<1>241 .INIT = 16'h0001;
  X_LUT4 \DLX_EXinst__n0007<1>241  (
    .ADR0(CHOICE3570),
    .ADR1(CHOICE3592),
    .ADR2(CHOICE3576),
    .ADR3(N164200),
    .O(\N164200/GROM )
  );
  X_BUF \N164200/XUSED  (
    .I(\N164200/FROM ),
    .O(N164200)
  );
  X_BUF \N164200/YUSED  (
    .I(\N164200/GROM ),
    .O(CHOICE5749)
  );
  defparam DLX_IDinst_Ker1073978.INIT = 16'h2222;
  X_LUT4 DLX_IDinst_Ker1073978 (
    .ADR0(DLX_IDinst_IR_opcode_field[4]),
    .ADR1(DLX_IDinst_IR_opcode_field[5]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\CHOICE1319/FROM )
  );
  defparam DLX_IDinst_Ker10739712.INIT = 16'hC400;
  X_LUT4 DLX_IDinst_Ker10739712 (
    .ADR0(DLX_IDinst_IR_opcode_field[0]),
    .ADR1(DLX_IDinst_IR_opcode_field[2]),
    .ADR2(DLX_IDinst_IR_opcode_field[1]),
    .ADR3(CHOICE1319),
    .O(\CHOICE1319/GROM )
  );
  X_BUF \CHOICE1319/XUSED  (
    .I(\CHOICE1319/FROM ),
    .O(CHOICE1319)
  );
  X_BUF \CHOICE1319/YUSED  (
    .I(\CHOICE1319/GROM ),
    .O(CHOICE1320)
  );
  defparam DLX_IDinst_Ker1085721.INIT = 16'h0800;
  X_LUT4 DLX_IDinst_Ker1085721 (
    .ADR0(DLX_IDinst_N108496),
    .ADR1(DLX_IDinst_N108443),
    .ADR2(DLX_IDinst_Ker1084541_1),
    .ADR3(DLX_IDinst_N107033),
    .O(\DLX_IDinst_N108574/FROM )
  );
  defparam DLX_IDinst_Ker1078681.INIT = 16'hECA0;
  X_LUT4 DLX_IDinst_Ker1078681 (
    .ADR0(DLX_IDinst_Ker1084541_1),
    .ADR1(DLX_IDinst__n0311),
    .ADR2(DLX_IDinst_IR_latched[30]),
    .ADR3(DLX_IDinst_N108574),
    .O(\DLX_IDinst_N108574/GROM )
  );
  X_BUF \DLX_IDinst_N108574/XUSED  (
    .I(\DLX_IDinst_N108574/FROM ),
    .O(DLX_IDinst_N108574)
  );
  X_BUF \DLX_IDinst_N108574/YUSED  (
    .I(\DLX_IDinst_N108574/GROM ),
    .O(DLX_IDinst_N107870)
  );
  defparam DLX_IDinst_Ker1085571.INIT = 16'h0020;
  X_LUT4 DLX_IDinst_Ker1085571 (
    .ADR0(DLX_MEMinst_reg_dst_out[2]),
    .ADR1(DLX_MEMinst_reg_dst_out[4]),
    .ADR2(DLX_MEMinst_reg_write_MEM),
    .ADR3(DLX_MEMinst_reg_dst_out[0]),
    .O(\DLX_IDinst_N108559/FROM )
  );
  defparam DLX_IDinst__n05781.INIT = 16'hC000;
  X_LUT4 DLX_IDinst__n05781 (
    .ADR0(VCC),
    .ADR1(DLX_MEMinst_reg_dst_out[3]),
    .ADR2(DLX_MEMinst_reg_dst_out[1]),
    .ADR3(DLX_IDinst_N108559),
    .O(\DLX_IDinst_N108559/GROM )
  );
  X_BUF \DLX_IDinst_N108559/XUSED  (
    .I(\DLX_IDinst_N108559/FROM ),
    .O(DLX_IDinst_N108559)
  );
  X_BUF \DLX_IDinst_N108559/YUSED  (
    .I(\DLX_IDinst_N108559/GROM ),
    .O(DLX_IDinst__n0578)
  );
  defparam \DLX_IFinst__n0001<20>_SW0 .INIT = 16'h0F55;
  X_LUT4 \DLX_IFinst__n0001<20>_SW0  (
    .ADR0(DLX_IFinst__n0015[20]),
    .ADR1(VCC),
    .ADR2(DLX_IFinst_PC[20]),
    .ADR3(DLX_IFinst__n0000),
    .O(\DLX_IFinst_NPC<20>/FROM )
  );
  defparam \DLX_IFinst__n0001<20> .INIT = 16'hC0F3;
  X_LUT4 \DLX_IFinst__n0001<20>  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(DLX_IDinst_branch_address[20]),
    .ADR3(N128911),
    .O(DLX_IFinst__n0001[20])
  );
  X_BUF \DLX_IFinst_NPC<20>/XUSED  (
    .I(\DLX_IFinst_NPC<20>/FROM ),
    .O(N128911)
  );
  defparam \DLX_IFinst__n0001<12>_SW0 .INIT = 16'h2277;
  X_LUT4 \DLX_IFinst__n0001<12>_SW0  (
    .ADR0(DLX_IFinst__n0000),
    .ADR1(DLX_IFinst_PC[12]),
    .ADR2(VCC),
    .ADR3(DLX_IFinst__n0015[12]),
    .O(\DLX_IFinst_NPC<12>/FROM )
  );
  defparam \DLX_IFinst__n0001<12> .INIT = 16'hC0CF;
  X_LUT4 \DLX_IFinst__n0001<12>  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_branch_address[12]),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(N129327),
    .O(\DLX_IFinst_NPC<12>/GROM )
  );
  X_BUF \DLX_IFinst_NPC<12>/XUSED  (
    .I(\DLX_IFinst_NPC<12>/FROM ),
    .O(N129327)
  );
  X_BUF \DLX_IFinst_NPC<12>/YUSED  (
    .I(\DLX_IFinst_NPC<12>/GROM ),
    .O(DLX_IFinst__n0001[12])
  );
  defparam \DLX_EXinst__n0007<0>299_SW1 .INIT = 16'h73F7;
  X_LUT4 \DLX_EXinst__n0007<0>299_SW1  (
    .ADR0(DLX_EXinst_Mcompar__n0091_inst_cy_196),
    .ADR1(\DLX_IDinst_Imm[1] ),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(DLX_IDinst_reg_out_B[31]),
    .O(\N164620/FROM )
  );
  defparam \DLX_EXinst__n0007<0>299_SW0 .INIT = 16'h4DFF;
  X_LUT4 \DLX_EXinst__n0007<0>299_SW0  (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(DLX_IDinst_reg_out_B[31]),
    .ADR2(DLX_EXinst_Mcompar__n0089_inst_cy_164),
    .ADR3(\DLX_IDinst_Imm[1] ),
    .O(\N164620/GROM )
  );
  X_BUF \N164620/XUSED  (
    .I(\N164620/FROM ),
    .O(N164620)
  );
  X_BUF \N164620/YUSED  (
    .I(\N164620/GROM ),
    .O(N164618)
  );
  defparam \DLX_IFinst__n0001<21>_SW0 .INIT = 16'h0A5F;
  X_LUT4 \DLX_IFinst__n0001<21>_SW0  (
    .ADR0(DLX_IFinst__n0000),
    .ADR1(VCC),
    .ADR2(DLX_IFinst_PC[21]),
    .ADR3(DLX_IFinst__n0015[21]),
    .O(\DLX_IFinst_NPC<21>/FROM )
  );
  defparam \DLX_IFinst__n0001<21> .INIT = 16'hC0CF;
  X_LUT4 \DLX_IFinst__n0001<21>  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_branch_address[21]),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(N128859),
    .O(DLX_IFinst__n0001[21])
  );
  X_BUF \DLX_IFinst_NPC<21>/XUSED  (
    .I(\DLX_IFinst_NPC<21>/FROM ),
    .O(N128859)
  );
  defparam \DLX_IFinst__n0001<13>_SW0 .INIT = 16'h4747;
  X_LUT4 \DLX_IFinst__n0001<13>_SW0  (
    .ADR0(DLX_IFinst_PC[13]),
    .ADR1(DLX_IFinst__n0000),
    .ADR2(DLX_IFinst__n0015[13]),
    .ADR3(VCC),
    .O(\DLX_IFinst_NPC<13>/FROM )
  );
  defparam \DLX_IFinst__n0001<13> .INIT = 16'h88DD;
  X_LUT4 \DLX_IFinst__n0001<13>  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(DLX_IDinst_branch_address[13]),
    .ADR2(VCC),
    .ADR3(N129275),
    .O(\DLX_IFinst_NPC<13>/GROM )
  );
  X_BUF \DLX_IFinst_NPC<13>/XUSED  (
    .I(\DLX_IFinst_NPC<13>/FROM ),
    .O(N129275)
  );
  X_BUF \DLX_IFinst_NPC<13>/YUSED  (
    .I(\DLX_IFinst_NPC<13>/GROM ),
    .O(DLX_IFinst__n0001[13])
  );
  defparam \DLX_IDinst__n0114<10>25 .INIT = 16'hF0F4;
  X_LUT4 \DLX_IDinst__n0114<10>25  (
    .ADR0(DLX_IDinst__n0453),
    .ADR1(CHOICE2231),
    .ADR2(CHOICE2235),
    .ADR3(DLX_IDinst_N108456),
    .O(\DLX_IDinst_branch_address<10>/FROM )
  );
  defparam \DLX_IDinst__n0114<10>31 .INIT = 16'hFFA0;
  X_LUT4 \DLX_IDinst__n0114<10>31  (
    .ADR0(DLX_IDinst__n0157[10]),
    .ADR1(VCC),
    .ADR2(N137082),
    .ADR3(CHOICE2236),
    .O(N140319)
  );
  X_BUF \DLX_IDinst_branch_address<10>/XUSED  (
    .I(\DLX_IDinst_branch_address<10>/FROM ),
    .O(CHOICE2236)
  );
  defparam DLX_IDinst_RegFile_26_19_693.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_26_19_693 (
    .I(DLX_IDinst_WB_data_eff[19]),
    .CE(DLX_IDinst__n0602),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_26_19)
  );
  defparam \DLX_IDinst__n0114<11>25 .INIT = 16'hFF04;
  X_LUT4 \DLX_IDinst__n0114<11>25  (
    .ADR0(DLX_IDinst__n0453),
    .ADR1(CHOICE2242),
    .ADR2(DLX_IDinst_N108456),
    .ADR3(CHOICE2246),
    .O(\DLX_IDinst_branch_address<11>/FROM )
  );
  defparam \DLX_IDinst__n0114<11>31 .INIT = 16'hFFC0;
  X_LUT4 \DLX_IDinst__n0114<11>31  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst__n0157[11]),
    .ADR2(N137082),
    .ADR3(CHOICE2247),
    .O(N140382)
  );
  X_BUF \DLX_IDinst_branch_address<11>/XUSED  (
    .I(\DLX_IDinst_branch_address<11>/FROM ),
    .O(CHOICE2247)
  );
  defparam \DLX_IDinst__n0114<27>20 .INIT = 16'hC0A0;
  X_LUT4 \DLX_IDinst__n0114<27>20  (
    .ADR0(DLX_IDinst__n0620[27]),
    .ADR1(DLX_MEMinst_RF_data_in[27]),
    .ADR2(DLX_IDinst_N107837),
    .ADR3(DLX_IDinst__n0175),
    .O(\DLX_IDinst_RegFile_2_12/FROM )
  );
  defparam \DLX_IDinst__n0114<20>20 .INIT = 16'h88C0;
  X_LUT4 \DLX_IDinst__n0114<20>20  (
    .ADR0(DLX_MEMinst_RF_data_in[20]),
    .ADR1(DLX_IDinst_N107837),
    .ADR2(DLX_IDinst__n0620[20]),
    .ADR3(DLX_IDinst__n0175),
    .O(\DLX_IDinst_RegFile_2_12/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_2_12/XUSED  (
    .I(\DLX_IDinst_RegFile_2_12/FROM ),
    .O(CHOICE2423)
  );
  X_BUF \DLX_IDinst_RegFile_2_12/YUSED  (
    .I(\DLX_IDinst_RegFile_2_12/GROM ),
    .O(CHOICE2357)
  );
  defparam \DLX_IDinst__n0114<20>25 .INIT = 16'hFF04;
  X_LUT4 \DLX_IDinst__n0114<20>25  (
    .ADR0(DLX_IDinst_N108456),
    .ADR1(CHOICE2353),
    .ADR2(DLX_IDinst__n0453),
    .ADR3(CHOICE2357),
    .O(\DLX_IDinst_branch_address<20>/FROM )
  );
  defparam \DLX_IDinst__n0114<20>31 .INIT = 16'hFFC0;
  X_LUT4 \DLX_IDinst__n0114<20>31  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst__n0157[20]),
    .ADR2(N137082),
    .ADR3(CHOICE2358),
    .O(N141013)
  );
  X_BUF \DLX_IDinst_branch_address<20>/XUSED  (
    .I(\DLX_IDinst_branch_address<20>/FROM ),
    .O(CHOICE2358)
  );
  defparam \DLX_IDinst__n0114<12>25 .INIT = 16'hF1F0;
  X_LUT4 \DLX_IDinst__n0114<12>25  (
    .ADR0(DLX_IDinst_N108456),
    .ADR1(DLX_IDinst__n0453),
    .ADR2(CHOICE2257),
    .ADR3(CHOICE2253),
    .O(\DLX_IDinst_branch_address<12>/FROM )
  );
  defparam \DLX_IDinst__n0114<12>31 .INIT = 16'hFF88;
  X_LUT4 \DLX_IDinst__n0114<12>31  (
    .ADR0(N137082),
    .ADR1(DLX_IDinst__n0157[12]),
    .ADR2(VCC),
    .ADR3(CHOICE2258),
    .O(N140445)
  );
  X_BUF \DLX_IDinst_branch_address<12>/XUSED  (
    .I(\DLX_IDinst_branch_address<12>/FROM ),
    .O(CHOICE2258)
  );
  defparam \DLX_IDinst__n0114<13>25 .INIT = 16'hFF04;
  X_LUT4 \DLX_IDinst__n0114<13>25  (
    .ADR0(DLX_IDinst__n0453),
    .ADR1(CHOICE2264),
    .ADR2(DLX_IDinst_N108456),
    .ADR3(CHOICE2268),
    .O(\DLX_IDinst_branch_address<13>/FROM )
  );
  defparam \DLX_IDinst__n0114<13>31 .INIT = 16'hFF88;
  X_LUT4 \DLX_IDinst__n0114<13>31  (
    .ADR0(DLX_IDinst__n0157[13]),
    .ADR1(N137082),
    .ADR2(VCC),
    .ADR3(CHOICE2269),
    .O(N140508)
  );
  X_BUF \DLX_IDinst_branch_address<13>/XUSED  (
    .I(\DLX_IDinst_branch_address<13>/FROM ),
    .O(CHOICE2269)
  );
  defparam DLX_IDinst_RegFile_27_11_694.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_27_11_694 (
    .I(DLX_IDinst_WB_data_eff[11]),
    .CE(DLX_IDinst__n0604),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_27_11)
  );
  defparam \DLX_IDinst__n0114<21>25 .INIT = 16'hAABA;
  X_LUT4 \DLX_IDinst__n0114<21>25  (
    .ADR0(CHOICE2368),
    .ADR1(DLX_IDinst__n0453),
    .ADR2(CHOICE2364),
    .ADR3(DLX_IDinst_N108456),
    .O(\DLX_IDinst_branch_address<21>/FROM )
  );
  defparam \DLX_IDinst__n0114<21>31 .INIT = 16'hFF88;
  X_LUT4 \DLX_IDinst__n0114<21>31  (
    .ADR0(DLX_IDinst__n0157[21]),
    .ADR1(N137082),
    .ADR2(VCC),
    .ADR3(CHOICE2369),
    .O(N141076)
  );
  X_BUF \DLX_IDinst_branch_address<21>/XUSED  (
    .I(\DLX_IDinst_branch_address<21>/FROM ),
    .O(CHOICE2369)
  );
  defparam \DLX_IFinst__n0001<30>_SW0 .INIT = 16'h05AF;
  X_LUT4 \DLX_IFinst__n0001<30>_SW0  (
    .ADR0(DLX_IFinst__n0000),
    .ADR1(VCC),
    .ADR2(DLX_IFinst__n0015[30]),
    .ADR3(DLX_IFinst_PC[30]),
    .O(\DLX_IFinst_NPC<30>/FROM )
  );
  defparam \DLX_IFinst__n0001<30> .INIT = 16'hC0CF;
  X_LUT4 \DLX_IFinst__n0001<30>  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_branch_address[30]),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(N128391),
    .O(DLX_IFinst__n0001[30])
  );
  X_BUF \DLX_IFinst_NPC<30>/XUSED  (
    .I(\DLX_IFinst_NPC<30>/FROM ),
    .O(N128391)
  );
  defparam \DLX_IFinst__n0001<14>_SW0 .INIT = 16'h4477;
  X_LUT4 \DLX_IFinst__n0001<14>_SW0  (
    .ADR0(DLX_IFinst_PC[14]),
    .ADR1(DLX_IFinst__n0000),
    .ADR2(VCC),
    .ADR3(DLX_IFinst__n0015[14]),
    .O(\DLX_IFinst_NPC<14>/FROM )
  );
  defparam \DLX_IFinst__n0001<14> .INIT = 16'h88BB;
  X_LUT4 \DLX_IFinst__n0001<14>  (
    .ADR0(DLX_IDinst_branch_address[14]),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(VCC),
    .ADR3(N129223),
    .O(\DLX_IFinst_NPC<14>/GROM )
  );
  X_BUF \DLX_IFinst_NPC<14>/XUSED  (
    .I(\DLX_IFinst_NPC<14>/FROM ),
    .O(N129223)
  );
  X_BUF \DLX_IFinst_NPC<14>/YUSED  (
    .I(\DLX_IFinst_NPC<14>/GROM ),
    .O(DLX_IFinst__n0001[14])
  );
  defparam \DLX_IFinst__n0001<22>_SW0 .INIT = 16'h3535;
  X_LUT4 \DLX_IFinst__n0001<22>_SW0  (
    .ADR0(DLX_IFinst__n0015[22]),
    .ADR1(DLX_IFinst_PC[22]),
    .ADR2(DLX_IFinst__n0000),
    .ADR3(VCC),
    .O(\DLX_IFinst_NPC<22>/FROM )
  );
  defparam \DLX_IFinst__n0001<22> .INIT = 16'h88BB;
  X_LUT4 \DLX_IFinst__n0001<22>  (
    .ADR0(DLX_IDinst_branch_address[22]),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(VCC),
    .ADR3(N128807),
    .O(DLX_IFinst__n0001[22])
  );
  X_BUF \DLX_IFinst_NPC<22>/XUSED  (
    .I(\DLX_IFinst_NPC<22>/FROM ),
    .O(N128807)
  );
  defparam \DLX_IDinst__n0114<22>25 .INIT = 16'hF0F2;
  X_LUT4 \DLX_IDinst__n0114<22>25  (
    .ADR0(CHOICE2375),
    .ADR1(DLX_IDinst_N108456),
    .ADR2(CHOICE2379),
    .ADR3(DLX_IDinst__n0453),
    .O(\DLX_IDinst_branch_address<22>/FROM )
  );
  defparam \DLX_IDinst__n0114<22>31 .INIT = 16'hFFC0;
  X_LUT4 \DLX_IDinst__n0114<22>31  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst__n0157[22]),
    .ADR2(N137082),
    .ADR3(CHOICE2380),
    .O(N141139)
  );
  X_BUF \DLX_IDinst_branch_address<22>/XUSED  (
    .I(\DLX_IDinst_branch_address<22>/FROM ),
    .O(CHOICE2380)
  );
  defparam \DLX_IDinst__n0114<14>25 .INIT = 16'hCCCE;
  X_LUT4 \DLX_IDinst__n0114<14>25  (
    .ADR0(CHOICE2275),
    .ADR1(CHOICE2279),
    .ADR2(DLX_IDinst__n0453),
    .ADR3(DLX_IDinst_N108456),
    .O(\DLX_IDinst_branch_address<14>/FROM )
  );
  defparam \DLX_IDinst__n0114<14>31 .INIT = 16'hFFC0;
  X_LUT4 \DLX_IDinst__n0114<14>31  (
    .ADR0(VCC),
    .ADR1(N137082),
    .ADR2(DLX_IDinst__n0157[14]),
    .ADR3(CHOICE2280),
    .O(N140571)
  );
  X_BUF \DLX_IDinst_branch_address<14>/XUSED  (
    .I(\DLX_IDinst_branch_address<14>/FROM ),
    .O(CHOICE2280)
  );
  defparam \DLX_IDinst__n0114<30>25 .INIT = 16'hCCDC;
  X_LUT4 \DLX_IDinst__n0114<30>25  (
    .ADR0(DLX_IDinst_N108456),
    .ADR1(CHOICE2390),
    .ADR2(CHOICE2386),
    .ADR3(DLX_IDinst__n0453),
    .O(\DLX_IDinst_branch_address<30>/FROM )
  );
  defparam \DLX_IDinst__n0114<30>31 .INIT = 16'hFF88;
  X_LUT4 \DLX_IDinst__n0114<30>31  (
    .ADR0(DLX_IDinst__n0157[30]),
    .ADR1(N137082),
    .ADR2(VCC),
    .ADR3(CHOICE2391),
    .O(N141202)
  );
  X_BUF \DLX_IDinst_branch_address<30>/XUSED  (
    .I(\DLX_IDinst_branch_address<30>/FROM ),
    .O(CHOICE2391)
  );
  defparam \DLX_IDinst__n0114<15>25 .INIT = 16'hCCCE;
  X_LUT4 \DLX_IDinst__n0114<15>25  (
    .ADR0(CHOICE2286),
    .ADR1(CHOICE2290),
    .ADR2(DLX_IDinst__n0453),
    .ADR3(DLX_IDinst_N108456),
    .O(\DLX_IDinst_branch_address<15>/FROM )
  );
  defparam \DLX_IDinst__n0114<15>31 .INIT = 16'hFFA0;
  X_LUT4 \DLX_IDinst__n0114<15>31  (
    .ADR0(DLX_IDinst__n0157[15]),
    .ADR1(VCC),
    .ADR2(N137082),
    .ADR3(CHOICE2291),
    .O(N140634)
  );
  X_BUF \DLX_IDinst_branch_address<15>/XUSED  (
    .I(\DLX_IDinst_branch_address<15>/FROM ),
    .O(CHOICE2291)
  );
  defparam \DLX_IDinst__n0114<23>25 .INIT = 16'hF1F0;
  X_LUT4 \DLX_IDinst__n0114<23>25  (
    .ADR0(DLX_IDinst_N108456),
    .ADR1(DLX_IDinst__n0453),
    .ADR2(CHOICE2467),
    .ADR3(CHOICE2463),
    .O(\DLX_IDinst_branch_address<23>/FROM )
  );
  defparam \DLX_IDinst__n0114<23>31 .INIT = 16'hFFA0;
  X_LUT4 \DLX_IDinst__n0114<23>31  (
    .ADR0(DLX_IDinst__n0157[23]),
    .ADR1(VCC),
    .ADR2(N137082),
    .ADR3(CHOICE2468),
    .O(N141643)
  );
  X_BUF \DLX_IDinst_branch_address<23>/XUSED  (
    .I(\DLX_IDinst_branch_address<23>/FROM ),
    .O(CHOICE2468)
  );
  defparam \DLX_IDinst__n0114<0>32 .INIT = 16'hC0A0;
  X_LUT4 \DLX_IDinst__n0114<0>32  (
    .ADR0(DLX_IDinst__n0620[0]),
    .ADR1(DLX_MEMinst_RF_data_in[0]),
    .ADR2(DLX_IDinst_N107837),
    .ADR3(DLX_IDinst__n0175),
    .O(\CHOICE3164/FROM )
  );
  defparam \DLX_IDinst__n0114<16>20 .INIT = 16'h8A80;
  X_LUT4 \DLX_IDinst__n0114<16>20  (
    .ADR0(DLX_IDinst_N107837),
    .ADR1(DLX_MEMinst_RF_data_in[16]),
    .ADR2(DLX_IDinst__n0175),
    .ADR3(DLX_IDinst__n0620[16]),
    .O(\CHOICE3164/GROM )
  );
  X_BUF \CHOICE3164/XUSED  (
    .I(\CHOICE3164/FROM ),
    .O(CHOICE3164)
  );
  X_BUF \CHOICE3164/YUSED  (
    .I(\CHOICE3164/GROM ),
    .O(CHOICE2313)
  );
  defparam \DLX_IDinst__n0114<31>28 .INIT = 16'hA280;
  X_LUT4 \DLX_IDinst__n0114<31>28  (
    .ADR0(DLX_IDinst_N107870),
    .ADR1(DLX_IDinst__n0175),
    .ADR2(DLX_MEMinst_RF_data_in[31]),
    .ADR3(DLX_IDinst__n0620[31]),
    .O(\DLX_IDinst_branch_address<31>/FROM )
  );
  defparam \DLX_IDinst__n0114<31>43 .INIT = 16'hFFEC;
  X_LUT4 \DLX_IDinst__n0114<31>43  (
    .ADR0(DLX_IDinst_N107609),
    .ADR1(CHOICE3173),
    .ADR2(DLX_IDinst__n0157[31]),
    .ADR3(CHOICE3178),
    .O(N145908)
  );
  X_BUF \DLX_IDinst_branch_address<31>/XUSED  (
    .I(\DLX_IDinst_branch_address<31>/FROM ),
    .O(CHOICE3178)
  );
  defparam \DLX_IDinst__n0114<8>20 .INIT = 16'hE200;
  X_LUT4 \DLX_IDinst__n0114<8>20  (
    .ADR0(DLX_IDinst__n0620[8]),
    .ADR1(DLX_IDinst__n0175),
    .ADR2(DLX_MEMinst_RF_data_in[8]),
    .ADR3(DLX_IDinst_N107837),
    .O(\CHOICE2213/FROM )
  );
  defparam \DLX_IDinst__n0114<24>20 .INIT = 16'hE200;
  X_LUT4 \DLX_IDinst__n0114<24>20  (
    .ADR0(DLX_IDinst__n0620[24]),
    .ADR1(DLX_IDinst__n0175),
    .ADR2(DLX_MEMinst_RF_data_in[24]),
    .ADR3(DLX_IDinst_N107837),
    .O(\CHOICE2213/GROM )
  );
  X_BUF \CHOICE2213/XUSED  (
    .I(\CHOICE2213/FROM ),
    .O(CHOICE2213)
  );
  X_BUF \CHOICE2213/YUSED  (
    .I(\CHOICE2213/GROM ),
    .O(CHOICE2456)
  );
  defparam DLX_EXinst_Ker7514760.INIT = 16'h00C0;
  X_LUT4 DLX_EXinst_Ker7514760 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_Imm_3_1),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(\DLX_IDinst_Imm[5] ),
    .O(\DLX_IDinst_RegFile_3_29/FROM )
  );
  defparam \DLX_EXinst__n0007<0>728_SW0 .INIT = 16'h8080;
  X_LUT4 \DLX_EXinst__n0007<0>728_SW0  (
    .ADR0(\DLX_IDinst_Imm[5] ),
    .ADR1(N147520),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(VCC),
    .O(\DLX_IDinst_RegFile_3_29/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_3_29/XUSED  (
    .I(\DLX_IDinst_RegFile_3_29/FROM ),
    .O(CHOICE1926)
  );
  X_BUF \DLX_IDinst_RegFile_3_29/YUSED  (
    .I(\DLX_IDinst_RegFile_3_29/GROM ),
    .O(N163953)
  );
  defparam \DLX_EXinst__n0007<0>760_SW0 .INIT = 16'hFF80;
  X_LUT4 \DLX_EXinst__n0007<0>760_SW0  (
    .ADR0(DLX_IDinst_IR_opcode_field[4]),
    .ADR1(DLX_EXinst_N76312),
    .ADR2(CHOICE5968),
    .ADR3(CHOICE6013),
    .O(\DLX_EXinst_ALU_result<0>/FROM )
  );
  defparam \DLX_EXinst__n0007<0>760 .INIT = 16'h0F0E;
  X_LUT4 \DLX_EXinst__n0007<0>760  (
    .ADR0(CHOICE6009),
    .ADR1(CHOICE5978),
    .ADR2(DLX_EXinst__n0036),
    .ADR3(N163238),
    .O(\DLX_EXinst_ALU_result<0>/GROM )
  );
  X_BUF \DLX_EXinst_ALU_result<0>/XUSED  (
    .I(\DLX_EXinst_ALU_result<0>/FROM ),
    .O(N163238)
  );
  X_BUF \DLX_EXinst_ALU_result<0>/YUSED  (
    .I(\DLX_EXinst_ALU_result<0>/GROM ),
    .O(CHOICE6016)
  );
  defparam DLX_IDinst_branch_address_16.INIT = 1'b0;
  X_SFF DLX_IDinst_branch_address_16 (
    .I(N140761),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_branch_address[16])
  );
  defparam \DLX_IDinst__n0114<16>25 .INIT = 16'hCCCE;
  X_LUT4 \DLX_IDinst__n0114<16>25  (
    .ADR0(CHOICE2309),
    .ADR1(CHOICE2313),
    .ADR2(DLX_IDinst__n0453),
    .ADR3(DLX_IDinst_N108456),
    .O(\DLX_IDinst_branch_address<16>/FROM )
  );
  defparam \DLX_IDinst__n0114<16>31 .INIT = 16'hFFA0;
  X_LUT4 \DLX_IDinst__n0114<16>31  (
    .ADR0(DLX_IDinst__n0157[16]),
    .ADR1(VCC),
    .ADR2(N137082),
    .ADR3(CHOICE2314),
    .O(N140761)
  );
  X_BUF \DLX_IDinst_branch_address<16>/XUSED  (
    .I(\DLX_IDinst_branch_address<16>/FROM ),
    .O(CHOICE2314)
  );
  defparam \DLX_IDinst__n0114<24>25 .INIT = 16'hCCCE;
  X_LUT4 \DLX_IDinst__n0114<24>25  (
    .ADR0(CHOICE2452),
    .ADR1(CHOICE2456),
    .ADR2(DLX_IDinst_N108456),
    .ADR3(DLX_IDinst__n0453),
    .O(\DLX_IDinst_branch_address<24>/FROM )
  );
  defparam \DLX_IDinst__n0114<24>31 .INIT = 16'hFCF0;
  X_LUT4 \DLX_IDinst__n0114<24>31  (
    .ADR0(VCC),
    .ADR1(N137082),
    .ADR2(CHOICE2457),
    .ADR3(DLX_IDinst__n0157[24]),
    .O(N141580)
  );
  X_BUF \DLX_IDinst_branch_address<24>/XUSED  (
    .I(\DLX_IDinst_branch_address<24>/FROM ),
    .O(CHOICE2457)
  );
  defparam \DLX_IDinst__n0114<25>25 .INIT = 16'hABAA;
  X_LUT4 \DLX_IDinst__n0114<25>25  (
    .ADR0(CHOICE2445),
    .ADR1(DLX_IDinst_N108456),
    .ADR2(DLX_IDinst__n0453),
    .ADR3(CHOICE2441),
    .O(\DLX_IDinst_branch_address<25>/FROM )
  );
  defparam \DLX_IDinst__n0114<25>31 .INIT = 16'hFF88;
  X_LUT4 \DLX_IDinst__n0114<25>31  (
    .ADR0(DLX_IDinst__n0157[25]),
    .ADR1(N137082),
    .ADR2(VCC),
    .ADR3(CHOICE2446),
    .O(N141517)
  );
  X_BUF \DLX_IDinst_branch_address<25>/XUSED  (
    .I(\DLX_IDinst_branch_address<25>/FROM ),
    .O(CHOICE2446)
  );
  defparam \DLX_IDinst__n0114<17>25 .INIT = 16'hFF10;
  X_LUT4 \DLX_IDinst__n0114<17>25  (
    .ADR0(DLX_IDinst_N108456),
    .ADR1(DLX_IDinst__n0453),
    .ADR2(CHOICE2320),
    .ADR3(CHOICE2324),
    .O(\DLX_IDinst_branch_address<17>/FROM )
  );
  defparam \DLX_IDinst__n0114<17>31 .INIT = 16'hFFA0;
  X_LUT4 \DLX_IDinst__n0114<17>31  (
    .ADR0(DLX_IDinst__n0157[17]),
    .ADR1(VCC),
    .ADR2(N137082),
    .ADR3(CHOICE2325),
    .O(N140824)
  );
  X_BUF \DLX_IDinst_branch_address<17>/XUSED  (
    .I(\DLX_IDinst_branch_address<17>/FROM ),
    .O(CHOICE2325)
  );
  defparam \DLX_IFinst__n0001<31>_SW0 .INIT = 16'h3355;
  X_LUT4 \DLX_IFinst__n0001<31>_SW0  (
    .ADR0(DLX_IFinst__n0015[31]),
    .ADR1(DLX_IFinst_PC[31]),
    .ADR2(VCC),
    .ADR3(DLX_IFinst__n0000),
    .O(\DLX_IFinst_NPC<31>/FROM )
  );
  defparam \DLX_IFinst__n0001<31> .INIT = 16'h88DD;
  X_LUT4 \DLX_IFinst__n0001<31>  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(DLX_IDinst_branch_address[31]),
    .ADR2(VCC),
    .ADR3(N128339),
    .O(DLX_IFinst__n0001[31])
  );
  X_BUF \DLX_IFinst_NPC<31>/XUSED  (
    .I(\DLX_IFinst_NPC<31>/FROM ),
    .O(N128339)
  );
  defparam \DLX_IFinst__n0001<15>_SW0 .INIT = 16'h03F3;
  X_LUT4 \DLX_IFinst__n0001<15>_SW0  (
    .ADR0(VCC),
    .ADR1(DLX_IFinst__n0015[15]),
    .ADR2(DLX_IFinst__n0000),
    .ADR3(DLX_IFinst_PC[15]),
    .O(\DLX_IFinst_NPC<15>/FROM )
  );
  defparam \DLX_IFinst__n0001<15> .INIT = 16'hC0F3;
  X_LUT4 \DLX_IFinst__n0001<15>  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(DLX_IDinst_branch_address[15]),
    .ADR3(N129171),
    .O(\DLX_IFinst_NPC<15>/GROM )
  );
  X_BUF \DLX_IFinst_NPC<15>/XUSED  (
    .I(\DLX_IFinst_NPC<15>/FROM ),
    .O(N129171)
  );
  X_BUF \DLX_IFinst_NPC<15>/YUSED  (
    .I(\DLX_IFinst_NPC<15>/GROM ),
    .O(DLX_IFinst__n0001[15])
  );
  defparam \DLX_IFinst__n0001<23>_SW0 .INIT = 16'h303F;
  X_LUT4 \DLX_IFinst__n0001<23>_SW0  (
    .ADR0(VCC),
    .ADR1(DLX_IFinst_PC[23]),
    .ADR2(DLX_IFinst__n0000),
    .ADR3(DLX_IFinst__n0015[23]),
    .O(\DLX_IFinst_NPC<23>/FROM )
  );
  defparam \DLX_IFinst__n0001<23> .INIT = 16'hC0CF;
  X_LUT4 \DLX_IFinst__n0001<23>  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_branch_address[23]),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(N128703),
    .O(DLX_IFinst__n0001[23])
  );
  X_BUF \DLX_IFinst_NPC<23>/XUSED  (
    .I(\DLX_IFinst_NPC<23>/FROM ),
    .O(N128703)
  );
  defparam \DLX_IDinst__n0114<26>25 .INIT = 16'hF0F4;
  X_LUT4 \DLX_IDinst__n0114<26>25  (
    .ADR0(DLX_IDinst_N108456),
    .ADR1(CHOICE2430),
    .ADR2(CHOICE2434),
    .ADR3(DLX_IDinst__n0453),
    .O(\DLX_IDinst_branch_address<26>/FROM )
  );
  defparam \DLX_IDinst__n0114<26>31 .INIT = 16'hFFA0;
  X_LUT4 \DLX_IDinst__n0114<26>31  (
    .ADR0(DLX_IDinst__n0157[26]),
    .ADR1(VCC),
    .ADR2(N137082),
    .ADR3(CHOICE2435),
    .O(N141454)
  );
  X_BUF \DLX_IDinst_branch_address<26>/XUSED  (
    .I(\DLX_IDinst_branch_address<26>/FROM ),
    .O(CHOICE2435)
  );
  defparam \DLX_IDinst__n0114<18>25 .INIT = 16'hAAAE;
  X_LUT4 \DLX_IDinst__n0114<18>25  (
    .ADR0(CHOICE2335),
    .ADR1(CHOICE2331),
    .ADR2(DLX_IDinst__n0453),
    .ADR3(DLX_IDinst_N108456),
    .O(\DLX_IDinst_branch_address<18>/FROM )
  );
  defparam \DLX_IDinst__n0114<18>31 .INIT = 16'hFF88;
  X_LUT4 \DLX_IDinst__n0114<18>31  (
    .ADR0(DLX_IDinst__n0157[18]),
    .ADR1(N137082),
    .ADR2(VCC),
    .ADR3(CHOICE2336),
    .O(N140887)
  );
  X_BUF \DLX_IDinst_branch_address<18>/XUSED  (
    .I(\DLX_IDinst_branch_address<18>/FROM ),
    .O(CHOICE2336)
  );
  defparam \DLX_IDinst__n0114<19>25 .INIT = 16'hABAA;
  X_LUT4 \DLX_IDinst__n0114<19>25  (
    .ADR0(CHOICE2346),
    .ADR1(DLX_IDinst__n0453),
    .ADR2(DLX_IDinst_N108456),
    .ADR3(CHOICE2342),
    .O(\DLX_IDinst_branch_address<19>/FROM )
  );
  defparam \DLX_IDinst__n0114<19>31 .INIT = 16'hFF88;
  X_LUT4 \DLX_IDinst__n0114<19>31  (
    .ADR0(N137082),
    .ADR1(DLX_IDinst__n0157[19]),
    .ADR2(VCC),
    .ADR3(CHOICE2347),
    .O(N140950)
  );
  X_BUF \DLX_IDinst_branch_address<19>/XUSED  (
    .I(\DLX_IDinst_branch_address<19>/FROM ),
    .O(CHOICE2347)
  );
  defparam \DLX_IDinst__n0114<27>25 .INIT = 16'hCCDC;
  X_LUT4 \DLX_IDinst__n0114<27>25  (
    .ADR0(DLX_IDinst_N108456),
    .ADR1(CHOICE2423),
    .ADR2(CHOICE2419),
    .ADR3(DLX_IDinst__n0453),
    .O(\DLX_IDinst_branch_address<27>/FROM )
  );
  defparam \DLX_IDinst__n0114<27>31 .INIT = 16'hFF88;
  X_LUT4 \DLX_IDinst__n0114<27>31  (
    .ADR0(DLX_IDinst__n0157[27]),
    .ADR1(N137082),
    .ADR2(VCC),
    .ADR3(CHOICE2424),
    .O(N141391)
  );
  X_BUF \DLX_IDinst_branch_address<27>/XUSED  (
    .I(\DLX_IDinst_branch_address<27>/FROM ),
    .O(CHOICE2424)
  );
  defparam \DLX_IDinst__n0147<28>1 .INIT = 16'hA280;
  X_LUT4 \DLX_IDinst__n0147<28>1  (
    .ADR0(DLX_IDinst_N107173),
    .ADR1(DLX_IDinst__n0176),
    .ADR2(DLX_MEMinst_RF_data_in[28]),
    .ADR3(DLX_IDinst__n0623[28]),
    .O(DLX_IDinst__n0147[28])
  );
  defparam \DLX_IDinst__n0114<28>20 .INIT = 16'hC480;
  X_LUT4 \DLX_IDinst__n0114<28>20  (
    .ADR0(DLX_IDinst__n0175),
    .ADR1(DLX_IDinst_N107837),
    .ADR2(DLX_MEMinst_RF_data_in[28]),
    .ADR3(DLX_IDinst__n0620[28]),
    .O(\DLX_IDinst_reg_out_B<28>/GROM )
  );
  X_BUF \DLX_IDinst_reg_out_B<28>/YUSED  (
    .I(\DLX_IDinst_reg_out_B<28>/GROM ),
    .O(CHOICE2412)
  );
  defparam \DLX_IDinst__n0114<28>25 .INIT = 16'hFF04;
  X_LUT4 \DLX_IDinst__n0114<28>25  (
    .ADR0(DLX_IDinst__n0453),
    .ADR1(CHOICE2408),
    .ADR2(DLX_IDinst_N108456),
    .ADR3(CHOICE2412),
    .O(\DLX_IDinst_branch_address<28>/FROM )
  );
  defparam \DLX_IDinst__n0114<28>31 .INIT = 16'hFFC0;
  X_LUT4 \DLX_IDinst__n0114<28>31  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst__n0157[28]),
    .ADR2(N137082),
    .ADR3(CHOICE2413),
    .O(N141328)
  );
  X_BUF \DLX_IDinst_branch_address<28>/XUSED  (
    .I(\DLX_IDinst_branch_address<28>/FROM ),
    .O(CHOICE2413)
  );
  defparam \DLX_IDinst__n0114<29>25 .INIT = 16'hFF02;
  X_LUT4 \DLX_IDinst__n0114<29>25  (
    .ADR0(CHOICE2397),
    .ADR1(DLX_IDinst_N108456),
    .ADR2(DLX_IDinst__n0453),
    .ADR3(CHOICE2401),
    .O(\DLX_IDinst_branch_address<29>/FROM )
  );
  defparam \DLX_IDinst__n0114<29>31 .INIT = 16'hFFA0;
  X_LUT4 \DLX_IDinst__n0114<29>31  (
    .ADR0(N137082),
    .ADR1(VCC),
    .ADR2(DLX_IDinst__n0157[29]),
    .ADR3(CHOICE2402),
    .O(N141265)
  );
  X_BUF \DLX_IDinst_branch_address<29>/XUSED  (
    .I(\DLX_IDinst_branch_address<29>/FROM ),
    .O(CHOICE2402)
  );
  defparam DLX_IDinst_RegFile_18_28_695.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_18_28_695 (
    .I(DLX_IDinst_WB_data_eff[28]),
    .CE(DLX_IDinst__n0586),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_18_28)
  );
  defparam \DLX_IFinst__n0001<24>_SW0 .INIT = 16'h05F5;
  X_LUT4 \DLX_IFinst__n0001<24>_SW0  (
    .ADR0(DLX_IFinst__n0015[24]),
    .ADR1(VCC),
    .ADR2(DLX_IFinst__n0000),
    .ADR3(DLX_IFinst_PC[24]),
    .O(\DLX_IFinst_NPC<24>/FROM )
  );
  defparam \DLX_IFinst__n0001<24> .INIT = 16'hA0AF;
  X_LUT4 \DLX_IFinst__n0001<24>  (
    .ADR0(DLX_IDinst_branch_address[24]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(N128755),
    .O(DLX_IFinst__n0001[24])
  );
  X_BUF \DLX_IFinst_NPC<24>/XUSED  (
    .I(\DLX_IFinst_NPC<24>/FROM ),
    .O(N128755)
  );
  defparam \DLX_IFinst__n0001<16>_SW0 .INIT = 16'h05AF;
  X_LUT4 \DLX_IFinst__n0001<16>_SW0  (
    .ADR0(DLX_IFinst__n0000),
    .ADR1(VCC),
    .ADR2(DLX_IFinst__n0015[16]),
    .ADR3(DLX_IFinst_PC[16]),
    .O(\DLX_IFinst_NPC<16>/FROM )
  );
  defparam \DLX_IFinst__n0001<16> .INIT = 16'h88DD;
  X_LUT4 \DLX_IFinst__n0001<16>  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(DLX_IDinst_branch_address[16]),
    .ADR2(VCC),
    .ADR3(N129119),
    .O(DLX_IFinst__n0001[16])
  );
  X_BUF \DLX_IFinst_NPC<16>/XUSED  (
    .I(\DLX_IFinst_NPC<16>/FROM ),
    .O(N129119)
  );
  defparam \DLX_EXinst__n0007<26>75_SW0 .INIT = 16'hEAEA;
  X_LUT4 \DLX_EXinst__n0007<26>75_SW0  (
    .ADR0(CHOICE5009),
    .ADR1(\DLX_EXinst_Mshift__n0022_Sh[58] ),
    .ADR2(DLX_EXinst__n0056),
    .ADR3(VCC),
    .O(\DLX_IDinst_RegFile_0_7/FROM )
  );
  defparam \DLX_EXinst__n0007<26>75 .INIT = 16'hD5C0;
  X_LUT4 \DLX_EXinst__n0007<26>75  (
    .ADR0(N146478),
    .ADR1(N138143),
    .ADR2(N147520),
    .ADR3(N163250),
    .O(\DLX_IDinst_RegFile_0_7/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_0_7/XUSED  (
    .I(\DLX_IDinst_RegFile_0_7/FROM ),
    .O(N163250)
  );
  X_BUF \DLX_IDinst_RegFile_0_7/YUSED  (
    .I(\DLX_IDinst_RegFile_0_7/GROM ),
    .O(CHOICE5014)
  );
  defparam \DLX_IFinst__n0001<25>_SW0 .INIT = 16'h330F;
  X_LUT4 \DLX_IFinst__n0001<25>_SW0  (
    .ADR0(VCC),
    .ADR1(DLX_IFinst_PC[25]),
    .ADR2(DLX_IFinst__n0015[25]),
    .ADR3(DLX_IFinst__n0000),
    .O(\DLX_IFinst_NPC<25>/FROM )
  );
  defparam \DLX_IFinst__n0001<25> .INIT = 16'h88DD;
  X_LUT4 \DLX_IFinst__n0001<25>  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(DLX_IDinst_branch_address[25]),
    .ADR2(VCC),
    .ADR3(N128651),
    .O(DLX_IFinst__n0001[25])
  );
  X_BUF \DLX_IFinst_NPC<25>/XUSED  (
    .I(\DLX_IFinst_NPC<25>/FROM ),
    .O(N128651)
  );
  defparam \DLX_IFinst__n0001<17>_SW0 .INIT = 16'h2727;
  X_LUT4 \DLX_IFinst__n0001<17>_SW0  (
    .ADR0(DLX_IFinst__n0000),
    .ADR1(DLX_IFinst_PC[17]),
    .ADR2(DLX_IFinst__n0015[17]),
    .ADR3(VCC),
    .O(\DLX_IFinst_NPC<17>/FROM )
  );
  defparam \DLX_IFinst__n0001<17> .INIT = 16'hA0F5;
  X_LUT4 \DLX_IFinst__n0001<17>  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_branch_address[17]),
    .ADR3(N129067),
    .O(DLX_IFinst__n0001[17])
  );
  X_BUF \DLX_IFinst_NPC<17>/XUSED  (
    .I(\DLX_IFinst_NPC<17>/FROM ),
    .O(N129067)
  );
  defparam \DLX_IFinst__n0001<26>_SW0 .INIT = 16'h3355;
  X_LUT4 \DLX_IFinst__n0001<26>_SW0  (
    .ADR0(DLX_IFinst__n0015[26]),
    .ADR1(DLX_IFinst_PC[26]),
    .ADR2(VCC),
    .ADR3(DLX_IFinst__n0000),
    .O(\DLX_IFinst_NPC<26>/FROM )
  );
  defparam \DLX_IFinst__n0001<26> .INIT = 16'hA0F5;
  X_LUT4 \DLX_IFinst__n0001<26>  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_branch_address[26]),
    .ADR3(N128599),
    .O(DLX_IFinst__n0001[26])
  );
  X_BUF \DLX_IFinst_NPC<26>/XUSED  (
    .I(\DLX_IFinst_NPC<26>/FROM ),
    .O(N128599)
  );
  defparam \DLX_IFinst__n0001<18>_SW0 .INIT = 16'h550F;
  X_LUT4 \DLX_IFinst__n0001<18>_SW0  (
    .ADR0(DLX_IFinst_PC[18]),
    .ADR1(VCC),
    .ADR2(DLX_IFinst__n0015[18]),
    .ADR3(DLX_IFinst__n0000),
    .O(\DLX_IFinst_NPC<18>/FROM )
  );
  defparam \DLX_IFinst__n0001<18> .INIT = 16'hA0AF;
  X_LUT4 \DLX_IFinst__n0001<18>  (
    .ADR0(DLX_IDinst_branch_address[18]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(N129015),
    .O(DLX_IFinst__n0001[18])
  );
  X_BUF \DLX_IFinst_NPC<18>/XUSED  (
    .I(\DLX_IFinst_NPC<18>/FROM ),
    .O(N129015)
  );
  defparam DLX_EXinst_Ker735971.INIT = 16'hF0CC;
  X_LUT4 DLX_EXinst_Ker735971 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[6]),
    .ADR2(DLX_IDinst_reg_out_A[4]),
    .ADR3(DLX_IDinst_reg_out_B[1]),
    .O(\DLX_EXinst_N73599/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0021_Sh<7>_SW0 .INIT = 16'hAFA0;
  X_LUT4 \DLX_EXinst_Mshift__n0021_Sh<7>_SW0  (
    .ADR0(DLX_IDinst_reg_out_A[4]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_Imm_1_1),
    .ADR3(DLX_IDinst_reg_out_A[6]),
    .O(\DLX_EXinst_N73599/GROM )
  );
  X_BUF \DLX_EXinst_N73599/XUSED  (
    .I(\DLX_EXinst_N73599/FROM ),
    .O(DLX_EXinst_N73599)
  );
  X_BUF \DLX_EXinst_N73599/YUSED  (
    .I(\DLX_EXinst_N73599/GROM ),
    .O(N130725)
  );
  defparam \DLX_IFinst__n0001<27>_SW0 .INIT = 16'h5353;
  X_LUT4 \DLX_IFinst__n0001<27>_SW0  (
    .ADR0(DLX_IFinst_PC[27]),
    .ADR1(DLX_IFinst__n0015[27]),
    .ADR2(DLX_IFinst__n0000),
    .ADR3(VCC),
    .O(\DLX_IFinst_NPC<27>/FROM )
  );
  defparam \DLX_IFinst__n0001<27> .INIT = 16'hC0CF;
  X_LUT4 \DLX_IFinst__n0001<27>  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_branch_address[27]),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(N128547),
    .O(DLX_IFinst__n0001[27])
  );
  X_BUF \DLX_IFinst_NPC<27>/XUSED  (
    .I(\DLX_IFinst_NPC<27>/FROM ),
    .O(N128547)
  );
  defparam \DLX_IFinst__n0001<19>_SW0 .INIT = 16'h11DD;
  X_LUT4 \DLX_IFinst__n0001<19>_SW0  (
    .ADR0(DLX_IFinst__n0015[19]),
    .ADR1(DLX_IFinst__n0000),
    .ADR2(VCC),
    .ADR3(DLX_IFinst_PC[19]),
    .O(\DLX_IFinst_NPC<19>/FROM )
  );
  defparam \DLX_IFinst__n0001<19> .INIT = 16'hA0F5;
  X_LUT4 \DLX_IFinst__n0001<19>  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_branch_address[19]),
    .ADR3(N128963),
    .O(DLX_IFinst__n0001[19])
  );
  X_BUF \DLX_IFinst_NPC<19>/XUSED  (
    .I(\DLX_IFinst_NPC<19>/FROM ),
    .O(N128963)
  );
  defparam \DLX_EXinst__n0007<2>241_SW0 .INIT = 16'h0F07;
  X_LUT4 \DLX_EXinst__n0007<2>241_SW0  (
    .ADR0(\DLX_EXinst_Mshift__n0023_Sh[2] ),
    .ADR1(DLX_EXinst_N76268),
    .ADR2(CHOICE5568),
    .ADR3(DLX_EXinst_N72822),
    .O(\DLX_MEMinst_opcode_of_WB<2>/FROM )
  );
  defparam \DLX_EXinst__n0007<2>241 .INIT = 16'h0001;
  X_LUT4 \DLX_EXinst__n0007<2>241  (
    .ADR0(CHOICE3576),
    .ADR1(CHOICE3570),
    .ADR2(CHOICE3592),
    .ADR3(N164082),
    .O(\DLX_MEMinst_opcode_of_WB<2>/GROM )
  );
  X_BUF \DLX_MEMinst_opcode_of_WB<2>/XUSED  (
    .I(\DLX_MEMinst_opcode_of_WB<2>/FROM ),
    .O(N164082)
  );
  X_BUF \DLX_MEMinst_opcode_of_WB<2>/YUSED  (
    .I(\DLX_MEMinst_opcode_of_WB<2>/GROM ),
    .O(CHOICE5570)
  );
  defparam DLX_IFinst_NPC_28.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_28 (
    .I(DLX_IFinst__n0001[28]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC[28])
  );
  defparam \DLX_IFinst__n0001<28>_SW0 .INIT = 16'h05F5;
  X_LUT4 \DLX_IFinst__n0001<28>_SW0  (
    .ADR0(DLX_IFinst__n0015[28]),
    .ADR1(VCC),
    .ADR2(DLX_IFinst__n0000),
    .ADR3(DLX_IFinst_PC[28]),
    .O(\DLX_IFinst_NPC<28>/FROM )
  );
  defparam \DLX_IFinst__n0001<28> .INIT = 16'hC0CF;
  X_LUT4 \DLX_IFinst__n0001<28>  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_branch_address[28]),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(N128495),
    .O(DLX_IFinst__n0001[28])
  );
  X_BUF \DLX_IFinst_NPC<28>/XUSED  (
    .I(\DLX_IFinst_NPC<28>/FROM ),
    .O(N128495)
  );
  defparam \DLX_IFinst__n0001<29>_SW0 .INIT = 16'h0A5F;
  X_LUT4 \DLX_IFinst__n0001<29>_SW0  (
    .ADR0(DLX_IFinst__n0000),
    .ADR1(VCC),
    .ADR2(DLX_IFinst_PC[29]),
    .ADR3(DLX_IFinst__n0015[29]),
    .O(\DLX_IFinst_NPC<29>/FROM )
  );
  defparam \DLX_IFinst__n0001<29> .INIT = 16'h88DD;
  X_LUT4 \DLX_IFinst__n0001<29>  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(DLX_IDinst_branch_address[29]),
    .ADR2(VCC),
    .ADR3(N128443),
    .O(DLX_IFinst__n0001[29])
  );
  X_BUF \DLX_IFinst_NPC<29>/XUSED  (
    .I(\DLX_IFinst_NPC<29>/FROM ),
    .O(N128443)
  );
  defparam \DLX_EXinst__n0007<5>241_SW0_SW0 .INIT = 16'hAAFE;
  X_LUT4 \DLX_EXinst__n0007<5>241_SW0_SW0  (
    .ADR0(CHOICE3959),
    .ADR1(CHOICE3948),
    .ADR2(CHOICE3945),
    .ADR3(DLX_IDinst_reg_out_B[4]),
    .O(\N164596/FROM )
  );
  defparam \DLX_EXinst__n0007<5>241_SW0 .INIT = 16'hFFEC;
  X_LUT4 \DLX_EXinst__n0007<5>241_SW0  (
    .ADR0(CHOICE3939),
    .ADR1(CHOICE3956),
    .ADR2(DLX_IDinst_reg_out_A[5]),
    .ADR3(N164596),
    .O(\N164596/GROM )
  );
  X_BUF \N164596/XUSED  (
    .I(\N164596/FROM ),
    .O(N164596)
  );
  X_BUF \N164596/YUSED  (
    .I(\N164596/GROM ),
    .O(N163182)
  );
  defparam \DLX_EXinst_Mshift__n0019_Sh<127>1 .INIT = 16'h0002;
  X_LUT4 \DLX_EXinst_Mshift__n0019_Sh<127>1  (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(DLX_IDinst_reg_out_B_2_1),
    .ADR2(DLX_IDinst_reg_out_B_3_1),
    .ADR3(DLX_EXinst_N73239),
    .O(\DLX_EXinst_Mshift__n0019_Sh<127>/FROM )
  );
  defparam \DLX_EXinst__n0007<15>16 .INIT = 16'hC800;
  X_LUT4 \DLX_EXinst__n0007<15>16  (
    .ADR0(DLX_EXinst_N76034),
    .ADR1(DLX_IDinst_reg_out_B[4]),
    .ADR2(DLX_EXinst_N76421),
    .ADR3(\DLX_EXinst_Mshift__n0019_Sh[127] ),
    .O(\DLX_EXinst_Mshift__n0019_Sh<127>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0019_Sh<127>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0019_Sh<127>/FROM ),
    .O(\DLX_EXinst_Mshift__n0019_Sh[127] )
  );
  X_BUF \DLX_EXinst_Mshift__n0019_Sh<127>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0019_Sh<127>/GROM ),
    .O(CHOICE4266)
  );
  defparam \DLX_EXinst__n0007<3>241_SW0 .INIT = 16'h0D0F;
  X_LUT4 \DLX_EXinst__n0007<3>241_SW0  (
    .ADR0(DLX_EXinst_N76268),
    .ADR1(DLX_EXinst_N72822),
    .ADR2(CHOICE5492),
    .ADR3(\DLX_EXinst_Mshift__n0023_Sh[3] ),
    .O(\N164138/FROM )
  );
  defparam \DLX_EXinst__n0007<3>241 .INIT = 16'h0001;
  X_LUT4 \DLX_EXinst__n0007<3>241  (
    .ADR0(CHOICE3576),
    .ADR1(CHOICE3592),
    .ADR2(CHOICE3570),
    .ADR3(N164138),
    .O(\N164138/GROM )
  );
  X_BUF \N164138/XUSED  (
    .I(\N164138/FROM ),
    .O(N164138)
  );
  X_BUF \N164138/YUSED  (
    .I(\N164138/GROM ),
    .O(CHOICE5494)
  );
  X_ZERO \DLX_IDinst_RegFile_12_0/LOGIC_ZERO_696  (
    .O(\DLX_IDinst_RegFile_12_0/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_6_697 (
    .IA(\DLX_IDinst_RegFile_12_0/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_12_0/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_65),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_6)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_651.INIT = 16'hF7B3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_651 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_49),
    .ADR2(DLX_IDinst_RegFile_13_0),
    .ADR3(DLX_IDinst_RegFile_12_0),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_65)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_661.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_661 (
    .ADR0(DLX_IDinst_RegFile_14_0),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_50),
    .ADR3(DLX_IDinst_RegFile_15_0),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_66)
  );
  X_BUF \DLX_IDinst_RegFile_12_0/COUTUSED  (
    .I(\DLX_IDinst_RegFile_12_0/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_7)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_7_698 (
    .IA(\DLX_IDinst_RegFile_12_0/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_6),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_66),
    .O(\DLX_IDinst_RegFile_12_0/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_12_0/CYINIT_699  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_5),
    .O(\DLX_IDinst_RegFile_12_0/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_20_0/LOGIC_ZERO_700  (
    .O(\DLX_IDinst_RegFile_20_0/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_10_701 (
    .IA(\DLX_IDinst_RegFile_20_0/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_20_0/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_69),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_10)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_691.INIT = 16'hF7D5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_691 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_53),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR2(DLX_IDinst_RegFile_21_0),
    .ADR3(DLX_IDinst_RegFile_20_0),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_69)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_701.INIT = 16'hF7D5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_701 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_54),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR2(DLX_IDinst_RegFile_23_0),
    .ADR3(DLX_IDinst_RegFile_22_0),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_70)
  );
  X_BUF \DLX_IDinst_RegFile_20_0/COUTUSED  (
    .I(\DLX_IDinst_RegFile_20_0/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_11)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_11_702 (
    .IA(\DLX_IDinst_RegFile_20_0/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_10),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_70),
    .O(\DLX_IDinst_RegFile_20_0/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_20_0/CYINIT_703  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_9),
    .O(\DLX_IDinst_RegFile_20_0/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_12_1/LOGIC_ZERO_704  (
    .O(\DLX_IDinst_RegFile_12_1/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_22_705 (
    .IA(\DLX_IDinst_RegFile_12_1/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_12_1/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_81),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_22)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_811.INIT = 16'hF5DD;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_811 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_49),
    .ADR1(DLX_IDinst_RegFile_12_1),
    .ADR2(DLX_IDinst_RegFile_13_1),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_81)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_821.INIT = 16'hCFAF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_821 (
    .ADR0(DLX_IDinst_RegFile_14_1),
    .ADR1(DLX_IDinst_RegFile_15_1),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_50),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_82)
  );
  X_BUF \DLX_IDinst_RegFile_12_1/COUTUSED  (
    .I(\DLX_IDinst_RegFile_12_1/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_23)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_23_706 (
    .IA(\DLX_IDinst_RegFile_12_1/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_22),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_82),
    .O(\DLX_IDinst_RegFile_12_1/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_12_1/CYINIT_707  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_21),
    .O(\DLX_IDinst_RegFile_12_1/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_20_1/LOGIC_ZERO_708  (
    .O(\DLX_IDinst_RegFile_20_1/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_26_709 (
    .IA(\DLX_IDinst_RegFile_20_1/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_20_1/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_85),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_26)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_851.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_851 (
    .ADR0(DLX_IDinst_RegFile_20_1),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_53),
    .ADR3(DLX_IDinst_RegFile_21_1),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_85)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_861.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_861 (
    .ADR0(DLX_IDinst_RegFile_23_1),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_54),
    .ADR2(DLX_IDinst_RegFile_22_1),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_86)
  );
  X_BUF \DLX_IDinst_RegFile_20_1/COUTUSED  (
    .I(\DLX_IDinst_RegFile_20_1/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_27)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_27_710 (
    .IA(\DLX_IDinst_RegFile_20_1/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_26),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_86),
    .O(\DLX_IDinst_RegFile_20_1/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_20_1/CYINIT_711  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_25),
    .O(\DLX_IDinst_RegFile_20_1/CYINIT )
  );
  defparam DLX_IDinst_RegFile_19_12_712.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_19_12_712 (
    .I(DLX_IDinst_WB_data_eff[12]),
    .CE(DLX_IDinst__n0588),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_19_12)
  );
  X_ZERO \DLX_IDinst_RegFile_12_2/LOGIC_ZERO_713  (
    .O(\DLX_IDinst_RegFile_12_2/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_38_714 (
    .IA(\DLX_IDinst_RegFile_12_2/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_12_2/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_97),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_38)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_971.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_971 (
    .ADR0(DLX_IDinst_RegFile_12_2),
    .ADR1(DLX_IDinst_RegFile_13_2),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_49),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_97)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_981.INIT = 16'hAFCF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_981 (
    .ADR0(DLX_IDinst_RegFile_15_2),
    .ADR1(DLX_IDinst_RegFile_14_2),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_50),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_98)
  );
  X_BUF \DLX_IDinst_RegFile_12_2/COUTUSED  (
    .I(\DLX_IDinst_RegFile_12_2/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_39)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_39_715 (
    .IA(\DLX_IDinst_RegFile_12_2/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_38),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_98),
    .O(\DLX_IDinst_RegFile_12_2/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_12_2/CYINIT_716  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_37),
    .O(\DLX_IDinst_RegFile_12_2/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_20_2/LOGIC_ZERO_717  (
    .O(\DLX_IDinst_RegFile_20_2/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_42_718 (
    .IA(\DLX_IDinst_RegFile_20_2/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_20_2/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_101),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_42)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1011.INIT = 16'hF7D5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1011 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_53),
    .ADR1(DLX_IDinst_jtarget[16]),
    .ADR2(DLX_IDinst_RegFile_21_2),
    .ADR3(DLX_IDinst_RegFile_20_2),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_101)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1021.INIT = 16'hDFD5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1021 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_54),
    .ADR1(DLX_IDinst_RegFile_23_2),
    .ADR2(DLX_IDinst_jtarget[16]),
    .ADR3(DLX_IDinst_RegFile_22_2),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_102)
  );
  X_BUF \DLX_IDinst_RegFile_20_2/COUTUSED  (
    .I(\DLX_IDinst_RegFile_20_2/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_43)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_43_719 (
    .IA(\DLX_IDinst_RegFile_20_2/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_42),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_102),
    .O(\DLX_IDinst_RegFile_20_2/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_20_2/CYINIT_720  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_41),
    .O(\DLX_IDinst_RegFile_20_2/CYINIT )
  );
  defparam DLX_IDinst_RegFile_19_20_721.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_19_20_721 (
    .I(DLX_IDinst_WB_data_eff[20]),
    .CE(DLX_IDinst__n0588),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_19_20)
  );
  X_ZERO \DLX_IDinst_RegFile_12_3/LOGIC_ZERO_722  (
    .O(\DLX_IDinst_RegFile_12_3/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_54_723 (
    .IA(\DLX_IDinst_RegFile_12_3/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_12_3/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_113),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_54)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1131.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1131 (
    .ADR0(DLX_IDinst_jtarget[16]),
    .ADR1(DLX_IDinst_RegFile_12_3),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_49),
    .ADR3(DLX_IDinst_RegFile_13_3),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_113)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1141.INIT = 16'hBFB3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1141 (
    .ADR0(DLX_IDinst_RegFile_15_3),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_50),
    .ADR2(DLX_IDinst_jtarget[16]),
    .ADR3(DLX_IDinst_RegFile_14_3),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_114)
  );
  X_BUF \DLX_IDinst_RegFile_12_3/COUTUSED  (
    .I(\DLX_IDinst_RegFile_12_3/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_55)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_55_724 (
    .IA(\DLX_IDinst_RegFile_12_3/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_54),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_114),
    .O(\DLX_IDinst_RegFile_12_3/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_12_3/CYINIT_725  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_53),
    .O(\DLX_IDinst_RegFile_12_3/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_20_3/LOGIC_ZERO_726  (
    .O(\DLX_IDinst_RegFile_20_3/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_58_727 (
    .IA(\DLX_IDinst_RegFile_20_3/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_20_3/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_117),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_58)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1171.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1171 (
    .ADR0(DLX_IDinst_RegFile_21_3),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_53),
    .ADR2(DLX_IDinst_RegFile_20_3),
    .ADR3(DLX_IDinst_jtarget[16]),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_117)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1181.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1181 (
    .ADR0(DLX_IDinst_jtarget[16]),
    .ADR1(DLX_IDinst_RegFile_22_3),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_54),
    .ADR3(DLX_IDinst_RegFile_23_3),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_118)
  );
  X_BUF \DLX_IDinst_RegFile_20_3/COUTUSED  (
    .I(\DLX_IDinst_RegFile_20_3/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_59)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_59_728 (
    .IA(\DLX_IDinst_RegFile_20_3/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_58),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_118),
    .O(\DLX_IDinst_RegFile_20_3/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_20_3/CYINIT_729  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_57),
    .O(\DLX_IDinst_RegFile_20_3/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_12_4/LOGIC_ZERO_730  (
    .O(\DLX_IDinst_RegFile_12_4/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_70_731 (
    .IA(\DLX_IDinst_RegFile_12_4/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_12_4/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_129),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_70)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1291.INIT = 16'hDFD5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1291 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_49),
    .ADR1(DLX_IDinst_RegFile_13_4),
    .ADR2(DLX_IDinst_jtarget[16]),
    .ADR3(DLX_IDinst_RegFile_12_4),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_129)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1301.INIT = 16'hFB3B;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1301 (
    .ADR0(DLX_IDinst_RegFile_14_4),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_50),
    .ADR2(DLX_IDinst_jtarget[16]),
    .ADR3(DLX_IDinst_RegFile_15_4),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_130)
  );
  X_BUF \DLX_IDinst_RegFile_12_4/COUTUSED  (
    .I(\DLX_IDinst_RegFile_12_4/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_71)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_71_732 (
    .IA(\DLX_IDinst_RegFile_12_4/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_70),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_130),
    .O(\DLX_IDinst_RegFile_12_4/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_12_4/CYINIT_733  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_69),
    .O(\DLX_IDinst_RegFile_12_4/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_13_0/LOGIC_ZERO_734  (
    .O(\DLX_IDinst_RegFile_13_0/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_518_735 (
    .IA(\DLX_IDinst_RegFile_13_0/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_13_0/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_593),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_518)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_5931.INIT = 16'hFB3B;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_5931 (
    .ADR0(DLX_IDinst_RegFile_12_0),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_577),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR3(DLX_IDinst_RegFile_13_0),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_593)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_5941.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_5941 (
    .ADR0(DLX_IDinst_RegFile_14_0),
    .ADR1(DLX_IDinst_RegFile_15_0),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_578),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_594)
  );
  X_BUF \DLX_IDinst_RegFile_13_0/COUTUSED  (
    .I(\DLX_IDinst_RegFile_13_0/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_519)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_519_736 (
    .IA(\DLX_IDinst_RegFile_13_0/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_518),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_594),
    .O(\DLX_IDinst_RegFile_13_0/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_13_0/CYINIT_737  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_517),
    .O(\DLX_IDinst_RegFile_13_0/CYINIT )
  );
  defparam \DLX_IDinst__n0018<3>1 .INIT = 16'hA888;
  X_LUT4 \DLX_IDinst__n0018<3>1  (
    .ADR0(DLX_IDinst_jtarget[14]),
    .ADR1(DLX_IDinst__n0453),
    .ADR2(DLX_IDinst_N107033),
    .ADR3(N139656),
    .O(\DLX_IDinst_rd_addr<3>/FROM )
  );
  defparam \DLX_IDinst__n0136<3>1 .INIT = 16'hFF80;
  X_LUT4 \DLX_IDinst__n0136<3>1  (
    .ADR0(DLX_IDinst_IR_latched[26]),
    .ADR1(DLX_IDinst_N108165),
    .ADR2(DLX_IDinst_IR_latched[27]),
    .ADR3(DLX_IDinst__n0018[3]),
    .O(DLX_IDinst__n0136[3])
  );
  X_BUF \DLX_IDinst_rd_addr<3>/XUSED  (
    .I(\DLX_IDinst_rd_addr<3>/FROM ),
    .O(DLX_IDinst__n0018[3])
  );
  defparam \DLX_IDinst__n0018<4>1 .INIT = 16'hA888;
  X_LUT4 \DLX_IDinst__n0018<4>1  (
    .ADR0(DLX_IDinst_jtarget[15]),
    .ADR1(DLX_IDinst__n0453),
    .ADR2(DLX_IDinst_N107033),
    .ADR3(N139656),
    .O(\DLX_IDinst_rd_addr<4>/FROM )
  );
  defparam \DLX_IDinst__n0136<4>1 .INIT = 16'hFF80;
  X_LUT4 \DLX_IDinst__n0136<4>1  (
    .ADR0(DLX_IDinst_N108165),
    .ADR1(DLX_IDinst_IR_latched[27]),
    .ADR2(DLX_IDinst_IR_latched[26]),
    .ADR3(DLX_IDinst__n0018[4]),
    .O(DLX_IDinst__n0136[4])
  );
  X_BUF \DLX_IDinst_rd_addr<4>/XUSED  (
    .I(\DLX_IDinst_rd_addr<4>/FROM ),
    .O(DLX_IDinst__n0018[4])
  );
  defparam \DLX_EXinst__n0007<27>223_SW0 .INIT = 16'hFAAA;
  X_LUT4 \DLX_EXinst__n0007<27>223_SW0  (
    .ADR0(CHOICE4974),
    .ADR1(VCC),
    .ADR2(\DLX_EXinst_Mshift__n0024_Sh[59] ),
    .ADR3(DLX_EXinst__n0081),
    .O(\N163428/FROM )
  );
  defparam \DLX_EXinst__n0007<27>223 .INIT = 16'hD5C0;
  X_LUT4 \DLX_EXinst__n0007<27>223  (
    .ADR0(N148323),
    .ADR1(N148609),
    .ADR2(N137952),
    .ADR3(N163428),
    .O(\N163428/GROM )
  );
  X_BUF \N163428/XUSED  (
    .I(\N163428/FROM ),
    .O(N163428)
  );
  X_BUF \N163428/YUSED  (
    .I(\N163428/GROM ),
    .O(CHOICE4979)
  );
  defparam \DLX_EXinst__n0007<9>65_SW0 .INIT = 16'h0777;
  X_LUT4 \DLX_EXinst__n0007<9>65_SW0  (
    .ADR0(DLX_EXinst_N76431),
    .ADR1(\DLX_EXinst_Mshift__n0024_Sh[57] ),
    .ADR2(DLX_EXinst_N76268),
    .ADR3(\DLX_EXinst_Mshift__n0023_Sh[41] ),
    .O(\N164207/FROM )
  );
  defparam \DLX_EXinst__n0007<9>65 .INIT = 16'h0001;
  X_LUT4 \DLX_EXinst__n0007<9>65  (
    .ADR0(CHOICE3576),
    .ADR1(N164207),
    .ADR2(CHOICE3592),
    .ADR3(CHOICE3570),
    .O(\N164207/GROM )
  );
  X_BUF \N164207/XUSED  (
    .I(\N164207/FROM ),
    .O(N164207)
  );
  X_BUF \N164207/YUSED  (
    .I(\N164207/GROM ),
    .O(CHOICE4525)
  );
  defparam \DLX_EXinst__n0007<9>81_SW0 .INIT = 16'hECA0;
  X_LUT4 \DLX_EXinst__n0007<9>81_SW0  (
    .ADR0(DLX_IDinst_reg_out_A[9]),
    .ADR1(DLX_EXinst_N75983),
    .ADR2(CHOICE4519),
    .ADR3(N138591),
    .O(\N163656/FROM )
  );
  defparam \DLX_EXinst__n0007<9>81 .INIT = 16'hFFEA;
  X_LUT4 \DLX_EXinst__n0007<9>81  (
    .ADR0(CHOICE4525),
    .ADR1(DLX_EXinst_ALU_result[9]),
    .ADR2(N134884),
    .ADR3(N163656),
    .O(\N163656/GROM )
  );
  X_BUF \N163656/XUSED  (
    .I(\N163656/FROM ),
    .O(N163656)
  );
  X_BUF \N163656/YUSED  (
    .I(\N163656/GROM ),
    .O(CHOICE4527)
  );
  defparam \DLX_EXinst__n0007<27>139_SW0 .INIT = 16'hFEFE;
  X_LUT4 \DLX_EXinst__n0007<27>139_SW0  (
    .ADR0(CHOICE4949),
    .ADR1(CHOICE4929),
    .ADR2(CHOICE4924),
    .ADR3(VCC),
    .O(\N163501/FROM )
  );
  defparam \DLX_EXinst__n0007<27>139 .INIT = 16'h3320;
  X_LUT4 \DLX_EXinst__n0007<27>139  (
    .ADR0(DLX_EXinst_N75993),
    .ADR1(DLX_EXinst__n0036),
    .ADR2(\DLX_EXinst_Mshift__n0021_Sh[43] ),
    .ADR3(N163501),
    .O(\N163501/GROM )
  );
  X_BUF \N163501/XUSED  (
    .I(\N163501/FROM ),
    .O(N163501)
  );
  X_BUF \N163501/YUSED  (
    .I(\N163501/GROM ),
    .O(CHOICE4953)
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<21>1_5_738 .INIT = 16'hCCCA;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<21>1_5_738  (
    .ADR0(DLX_IFinst_IR_latched[21]),
    .ADR1(DLX_IDinst_current_IR[21]),
    .ADR2(DLX_IDinst_counter[0]),
    .ADR3(DLX_IDinst_counter[1]),
    .O(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5/FROM )
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<21>1_1_739 .INIT = 16'hFE04;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<21>1_1_739  (
    .ADR0(DLX_IDinst_counter[1]),
    .ADR1(DLX_IFinst_IR_latched[21]),
    .ADR2(DLX_IDinst_counter[0]),
    .ADR3(DLX_IDinst_current_IR[21]),
    .O(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5/GROM )
  );
  X_BUF \DLX_IDinst_Mmux_IR_latched_Result<21>1_5/XUSED  (
    .I(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5/FROM ),
    .O(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 )
  );
  X_BUF \DLX_IDinst_Mmux_IR_latched_Result<21>1_5/YUSED  (
    .I(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5/GROM ),
    .O(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 )
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<21>1_4_740 .INIT = 16'hCCD8;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<21>1_4_740  (
    .ADR0(DLX_IDinst_counter[0]),
    .ADR1(DLX_IDinst_current_IR[21]),
    .ADR2(DLX_IFinst_IR_latched[21]),
    .ADR3(DLX_IDinst_counter[1]),
    .O(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4/FROM )
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<21>1_2_741 .INIT = 16'hFE10;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<21>1_2_741  (
    .ADR0(DLX_IDinst_counter[0]),
    .ADR1(DLX_IDinst_counter[1]),
    .ADR2(DLX_IFinst_IR_latched[21]),
    .ADR3(DLX_IDinst_current_IR[21]),
    .O(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4/GROM )
  );
  X_BUF \DLX_IDinst_Mmux_IR_latched_Result<21>1_4/XUSED  (
    .I(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4/FROM ),
    .O(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 )
  );
  X_BUF \DLX_IDinst_Mmux_IR_latched_Result<21>1_4/YUSED  (
    .I(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4/GROM ),
    .O(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 )
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<21>1 .INIT = 16'hF0E2;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<21>1  (
    .ADR0(DLX_IFinst_IR_latched[21]),
    .ADR1(DLX_IDinst_counter[0]),
    .ADR2(DLX_IDinst_current_IR[21]),
    .ADR3(DLX_IDinst_counter[1]),
    .O(\DLX_IDinst_current_IR<21>/FROM )
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<21>1_3_742 .INIT = 16'hCCD8;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<21>1_3_742  (
    .ADR0(DLX_IDinst_counter[0]),
    .ADR1(DLX_IDinst_current_IR[21]),
    .ADR2(DLX_IFinst_IR_latched[21]),
    .ADR3(DLX_IDinst_counter[1]),
    .O(\DLX_IDinst_current_IR<21>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<21>/XUSED  (
    .I(\DLX_IDinst_current_IR<21>/FROM ),
    .O(DLX_IDinst_jtarget[21])
  );
  X_BUF \DLX_IDinst_current_IR<21>/YUSED  (
    .I(\DLX_IDinst_current_IR<21>/GROM ),
    .O(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 )
  );
  defparam DLX_EXinst_Ker729361.INIT = 16'hAAF0;
  X_LUT4 DLX_EXinst_Ker729361 (
    .ADR0(DLX_IDinst_reg_out_A[7]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[9]),
    .ADR3(\DLX_IDinst_Imm[1] ),
    .O(\DLX_EXinst_N72938/FROM )
  );
  defparam DLX_EXinst_Ker731111.INIT = 16'hAAF0;
  X_LUT4 DLX_EXinst_Ker731111 (
    .ADR0(DLX_IDinst_reg_out_A[9]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[7]),
    .ADR3(\DLX_IDinst_Imm[1] ),
    .O(\DLX_EXinst_N72938/GROM )
  );
  X_BUF \DLX_EXinst_N72938/XUSED  (
    .I(\DLX_EXinst_N72938/FROM ),
    .O(DLX_EXinst_N72938)
  );
  X_BUF \DLX_EXinst_N72938/YUSED  (
    .I(\DLX_EXinst_N72938/GROM ),
    .O(DLX_EXinst_N73113)
  );
  defparam DLX_EXinst_Ker730311.INIT = 16'hB8B8;
  X_LUT4 DLX_EXinst_Ker730311 (
    .ADR0(DLX_IDinst_reg_out_A[11]),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(DLX_IDinst_reg_out_A[9]),
    .ADR3(VCC),
    .O(\DLX_EXinst_N73033/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0019_Sh<8>1 .INIT = 16'hEE44;
  X_LUT4 \DLX_EXinst_Mshift__n0019_Sh<8>1  (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(DLX_EXinst_N73429),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N73033),
    .O(\DLX_EXinst_N73033/GROM )
  );
  X_BUF \DLX_EXinst_N73033/XUSED  (
    .I(\DLX_EXinst_N73033/FROM ),
    .O(DLX_EXinst_N73033)
  );
  X_BUF \DLX_EXinst_N73033/YUSED  (
    .I(\DLX_EXinst_N73033/GROM ),
    .O(\DLX_EXinst_Mshift__n0019_Sh[8] )
  );
  defparam DLX_EXinst_Ker731211.INIT = 16'hCCF0;
  X_LUT4 DLX_EXinst_Ker731211 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[13]),
    .ADR2(DLX_IDinst_reg_out_A[11]),
    .ADR3(\DLX_IDinst_Imm[1] ),
    .O(\DLX_EXinst_N73123/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0022_Sh<10>1 .INIT = 16'hFA0A;
  X_LUT4 \DLX_EXinst_Mshift__n0022_Sh<10>1  (
    .ADR0(DLX_EXinst_N73514),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_Imm_0_1),
    .ADR3(DLX_EXinst_N73123),
    .O(\DLX_EXinst_N73123/GROM )
  );
  X_BUF \DLX_EXinst_N73123/XUSED  (
    .I(\DLX_EXinst_N73123/FROM ),
    .O(DLX_EXinst_N73123)
  );
  X_BUF \DLX_EXinst_N73123/YUSED  (
    .I(\DLX_EXinst_N73123/GROM ),
    .O(\DLX_EXinst_Mshift__n0022_Sh[10] )
  );
  defparam DLX_EXinst_Ker728661.INIT = 16'hCACA;
  X_LUT4 DLX_EXinst_Ker728661 (
    .ADR0(DLX_IDinst_reg_out_A[15]),
    .ADR1(DLX_IDinst_reg_out_A[13]),
    .ADR2(DLX_IDinst_reg_out_B[1]),
    .ADR3(VCC),
    .O(\DLX_EXinst_N72868/FROM )
  );
  defparam DLX_EXinst_Ker730411.INIT = 16'hF5A0;
  X_LUT4 DLX_EXinst_Ker730411 (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[15]),
    .ADR3(DLX_IDinst_reg_out_A[13]),
    .O(\DLX_EXinst_N72868/GROM )
  );
  X_BUF \DLX_EXinst_N72868/XUSED  (
    .I(\DLX_EXinst_N72868/FROM ),
    .O(DLX_EXinst_N72868)
  );
  X_BUF \DLX_EXinst_N72868/YUSED  (
    .I(\DLX_EXinst_N72868/GROM ),
    .O(DLX_EXinst_N73043)
  );
  defparam DLX_EXinst_Ker740011.INIT = 16'hACAC;
  X_LUT4 DLX_EXinst_Ker740011 (
    .ADR0(\DLX_EXinst_Mshift__n0021_Sh[11] ),
    .ADR1(\DLX_EXinst_Mshift__n0021_Sh[19] ),
    .ADR2(\DLX_IDinst_Imm[3] ),
    .ADR3(VCC),
    .O(\DLX_EXinst_N74003/GROM )
  );
  X_BUF \DLX_EXinst_N74003/YUSED  (
    .I(\DLX_EXinst_N74003/GROM ),
    .O(DLX_EXinst_N74003)
  );
  defparam DLX_EXinst_Ker729311.INIT = 16'hFC30;
  X_LUT4 DLX_EXinst_Ker729311 (
    .ADR0(VCC),
    .ADR1(\DLX_IDinst_Imm[1] ),
    .ADR2(DLX_IDinst_reg_out_A[7]),
    .ADR3(DLX_IDinst_reg_out_A[5]),
    .O(\DLX_EXinst_N72933/FROM )
  );
  defparam DLX_EXinst_Ker731061.INIT = 16'hACAC;
  X_LUT4 DLX_EXinst_Ker731061 (
    .ADR0(DLX_IDinst_reg_out_A[7]),
    .ADR1(DLX_IDinst_reg_out_A[5]),
    .ADR2(\DLX_IDinst_Imm[1] ),
    .ADR3(VCC),
    .O(\DLX_EXinst_N72933/GROM )
  );
  X_BUF \DLX_EXinst_N72933/XUSED  (
    .I(\DLX_EXinst_N72933/FROM ),
    .O(DLX_EXinst_N72933)
  );
  X_BUF \DLX_EXinst_N72933/YUSED  (
    .I(\DLX_EXinst_N72933/GROM ),
    .O(DLX_EXinst_N73108)
  );
  defparam DLX_EXinst_Ker728461.INIT = 16'hE2E2;
  X_LUT4 DLX_EXinst_Ker728461 (
    .ADR0(DLX_IDinst_reg_out_A[7]),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(DLX_IDinst_reg_out_A[5]),
    .ADR3(VCC),
    .O(\DLX_EXinst_N72848/FROM )
  );
  defparam DLX_EXinst_Ker730261.INIT = 16'hE2E2;
  X_LUT4 DLX_EXinst_Ker730261 (
    .ADR0(DLX_IDinst_reg_out_A[7]),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(DLX_IDinst_reg_out_A[9]),
    .ADR3(VCC),
    .O(\DLX_EXinst_N72848/GROM )
  );
  X_BUF \DLX_EXinst_N72848/XUSED  (
    .I(\DLX_EXinst_N72848/FROM ),
    .O(DLX_EXinst_N72848)
  );
  X_BUF \DLX_EXinst_N72848/YUSED  (
    .I(\DLX_EXinst_N72848/GROM ),
    .O(DLX_EXinst_N73028)
  );
  defparam DLX_EXinst_Ker731311.INIT = 16'hDD88;
  X_LUT4 DLX_EXinst_Ker731311 (
    .ADR0(\DLX_IDinst_Imm[1] ),
    .ADR1(DLX_IDinst_reg_out_A[17]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[15]),
    .O(\DLX_EXinst_N73133/FROM )
  );
  defparam DLX_EXinst_Ker74699_SW0.INIT = 16'hFA50;
  X_LUT4 DLX_EXinst_Ker74699_SW0 (
    .ADR0(\DLX_IDinst_Imm[0] ),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N73524),
    .ADR3(DLX_EXinst_N73133),
    .O(\DLX_EXinst_N73133/GROM )
  );
  X_BUF \DLX_EXinst_N73133/XUSED  (
    .I(\DLX_EXinst_N73133/FROM ),
    .O(DLX_EXinst_N73133)
  );
  X_BUF \DLX_EXinst_N73133/YUSED  (
    .I(\DLX_EXinst_N73133/GROM ),
    .O(N130825)
  );
  defparam DLX_EXinst_Ker731361.INIT = 16'hCCAA;
  X_LUT4 DLX_EXinst_Ker731361 (
    .ADR0(DLX_IDinst_reg_out_A[17]),
    .ADR1(DLX_IDinst_reg_out_A[19]),
    .ADR2(VCC),
    .ADR3(\DLX_IDinst_Imm[1] ),
    .O(\DLX_EXinst_N73138/FROM )
  );
  defparam DLX_EXinst_Ker730511.INIT = 16'hEE44;
  X_LUT4 DLX_EXinst_Ker730511 (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(DLX_IDinst_reg_out_A[17]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[19]),
    .O(\DLX_EXinst_N73138/GROM )
  );
  X_BUF \DLX_EXinst_N73138/XUSED  (
    .I(\DLX_EXinst_N73138/FROM ),
    .O(DLX_EXinst_N73138)
  );
  X_BUF \DLX_EXinst_N73138/YUSED  (
    .I(\DLX_EXinst_N73138/GROM ),
    .O(DLX_EXinst_N73053)
  );
  defparam DLX_EXinst_Ker731161.INIT = 16'hCFC0;
  X_LUT4 DLX_EXinst_Ker731161 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[11]),
    .ADR2(\DLX_IDinst_Imm[1] ),
    .ADR3(DLX_IDinst_reg_out_A[9]),
    .O(\DLX_EXinst_N73118/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0022_Sh<8>1 .INIT = 16'hEE22;
  X_LUT4 \DLX_EXinst_Mshift__n0022_Sh<8>1  (
    .ADR0(DLX_EXinst_N73554),
    .ADR1(DLX_IDinst_Imm_0_1),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N73118),
    .O(\DLX_EXinst_N73118/GROM )
  );
  X_BUF \DLX_EXinst_N73118/XUSED  (
    .I(\DLX_EXinst_N73118/FROM ),
    .O(DLX_EXinst_N73118)
  );
  X_BUF \DLX_EXinst_N73118/YUSED  (
    .I(\DLX_EXinst_N73118/GROM ),
    .O(\DLX_EXinst_Mshift__n0022_Sh[8] )
  );
  defparam DLX_EXinst_Ker730361.INIT = 16'hE2E2;
  X_LUT4 DLX_EXinst_Ker730361 (
    .ADR0(DLX_IDinst_reg_out_A[11]),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(DLX_IDinst_reg_out_A[13]),
    .ADR3(VCC),
    .O(\DLX_EXinst_N73038/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0019_Sh<10>1 .INIT = 16'hFA0A;
  X_LUT4 \DLX_EXinst_Mshift__n0019_Sh<10>1  (
    .ADR0(DLX_EXinst_N73384),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[0]),
    .ADR3(DLX_EXinst_N73038),
    .O(\DLX_EXinst_N73038/GROM )
  );
  X_BUF \DLX_EXinst_N73038/XUSED  (
    .I(\DLX_EXinst_N73038/FROM ),
    .O(DLX_EXinst_N73038)
  );
  X_BUF \DLX_EXinst_N73038/YUSED  (
    .I(\DLX_EXinst_N73038/GROM ),
    .O(\DLX_EXinst_Mshift__n0019_Sh[10] )
  );
  defparam DLX_EXinst_Ker729711.INIT = 16'hFA50;
  X_LUT4 DLX_EXinst_Ker729711 (
    .ADR0(\DLX_IDinst_Imm[1] ),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[23]),
    .ADR3(DLX_IDinst_reg_out_A[21]),
    .O(\DLX_EXinst_N72973/FROM )
  );
  defparam DLX_EXinst_Ker731411.INIT = 16'hDD88;
  X_LUT4 DLX_EXinst_Ker731411 (
    .ADR0(\DLX_IDinst_Imm[1] ),
    .ADR1(DLX_IDinst_reg_out_A[21]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[19]),
    .O(\DLX_EXinst_N72973/GROM )
  );
  X_BUF \DLX_EXinst_N72973/XUSED  (
    .I(\DLX_EXinst_N72973/FROM ),
    .O(DLX_EXinst_N72973)
  );
  X_BUF \DLX_EXinst_N72973/YUSED  (
    .I(\DLX_EXinst_N72973/GROM ),
    .O(DLX_EXinst_N73143)
  );
  defparam DLX_IDinst_RegFile_19_28_743.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_19_28_743 (
    .I(DLX_IDinst_WB_data_eff[28]),
    .CE(DLX_IDinst__n0588),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_19_28)
  );
  defparam DLX_EXinst_Ker730611.INIT = 16'hFC30;
  X_LUT4 DLX_EXinst_Ker730611 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(DLX_IDinst_reg_out_A[21]),
    .ADR3(DLX_IDinst_reg_out_A[23]),
    .O(\DLX_EXinst_N73063/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0019_Sh<20>1 .INIT = 16'hEE22;
  X_LUT4 \DLX_EXinst_Mshift__n0019_Sh<20>1  (
    .ADR0(DLX_EXinst_N73409),
    .ADR1(DLX_IDinst_reg_out_B[0]),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N73063),
    .O(\DLX_EXinst_N73063/GROM )
  );
  X_BUF \DLX_EXinst_N73063/XUSED  (
    .I(\DLX_EXinst_N73063/FROM ),
    .O(DLX_EXinst_N73063)
  );
  X_BUF \DLX_EXinst_N73063/YUSED  (
    .I(\DLX_EXinst_N73063/GROM ),
    .O(\DLX_EXinst_Mshift__n0019_Sh[20] )
  );
  defparam DLX_EXinst_Ker729511.INIT = 16'hAFA0;
  X_LUT4 DLX_EXinst_Ker729511 (
    .ADR0(DLX_IDinst_reg_out_A[13]),
    .ADR1(VCC),
    .ADR2(\DLX_IDinst_Imm[1] ),
    .ADR3(DLX_IDinst_reg_out_A[15]),
    .O(\DLX_EXinst_N72953/FROM )
  );
  defparam DLX_EXinst_Ker731261.INIT = 16'hFA0A;
  X_LUT4 DLX_EXinst_Ker731261 (
    .ADR0(DLX_IDinst_reg_out_A[13]),
    .ADR1(VCC),
    .ADR2(\DLX_IDinst_Imm[1] ),
    .ADR3(DLX_IDinst_reg_out_A[15]),
    .O(\DLX_EXinst_N72953/GROM )
  );
  X_BUF \DLX_EXinst_N72953/XUSED  (
    .I(\DLX_EXinst_N72953/FROM ),
    .O(DLX_EXinst_N72953)
  );
  X_BUF \DLX_EXinst_N72953/YUSED  (
    .I(\DLX_EXinst_N72953/GROM ),
    .O(DLX_EXinst_N73128)
  );
  defparam DLX_EXinst_Ker730461.INIT = 16'hFC0C;
  X_LUT4 DLX_EXinst_Ker730461 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[15]),
    .ADR2(DLX_IDinst_reg_out_B[1]),
    .ADR3(DLX_IDinst_reg_out_A[17]),
    .O(\DLX_EXinst_N73048/FROM )
  );
  defparam DLX_EXinst_Ker74439_SW0.INIT = 16'hFC0C;
  X_LUT4 DLX_EXinst_Ker74439_SW0 (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N73394),
    .ADR2(DLX_IDinst_reg_out_B[0]),
    .ADR3(DLX_EXinst_N73048),
    .O(\DLX_EXinst_N73048/GROM )
  );
  X_BUF \DLX_EXinst_N73048/XUSED  (
    .I(\DLX_EXinst_N73048/FROM ),
    .O(DLX_EXinst_N73048)
  );
  X_BUF \DLX_EXinst_N73048/YUSED  (
    .I(\DLX_EXinst_N73048/GROM ),
    .O(N130569)
  );
  defparam DLX_EXinst_Ker740221.INIT = 16'hAAF0;
  X_LUT4 DLX_EXinst_Ker740221 (
    .ADR0(\DLX_EXinst_Mshift__n0023_Sh[13] ),
    .ADR1(VCC),
    .ADR2(\DLX_EXinst_Mshift__n0023_Sh[21] ),
    .ADR3(DLX_IDinst_reg_out_B[3]),
    .O(\DLX_EXinst_N74024/FROM )
  );
  defparam \DLX_EXinst__n0007<25>201 .INIT = 16'hA808;
  X_LUT4 \DLX_EXinst__n0007<25>201  (
    .ADR0(DLX_EXinst__n0080),
    .ADR1(N133048),
    .ADR2(DLX_IDinst_reg_out_B[2]),
    .ADR3(DLX_EXinst_N74024),
    .O(\DLX_EXinst_N74024/GROM )
  );
  X_BUF \DLX_EXinst_N74024/XUSED  (
    .I(\DLX_EXinst_N74024/FROM ),
    .O(DLX_EXinst_N74024)
  );
  X_BUF \DLX_EXinst_N74024/YUSED  (
    .I(\DLX_EXinst_N74024/GROM ),
    .O(CHOICE5108)
  );
  defparam DLX_EXinst_Ker729761.INIT = 16'hFA50;
  X_LUT4 DLX_EXinst_Ker729761 (
    .ADR0(\DLX_IDinst_Imm[1] ),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[25]),
    .ADR3(DLX_IDinst_reg_out_A[23]),
    .O(\DLX_EXinst_N72978/FROM )
  );
  defparam DLX_EXinst_Ker731511.INIT = 16'hFA50;
  X_LUT4 DLX_EXinst_Ker731511 (
    .ADR0(\DLX_IDinst_Imm[1] ),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[23]),
    .ADR3(DLX_IDinst_reg_out_A[25]),
    .O(\DLX_EXinst_N72978/GROM )
  );
  X_BUF \DLX_EXinst_N72978/XUSED  (
    .I(\DLX_EXinst_N72978/FROM ),
    .O(DLX_EXinst_N72978)
  );
  X_BUF \DLX_EXinst_N72978/YUSED  (
    .I(\DLX_EXinst_N72978/GROM ),
    .O(DLX_EXinst_N73153)
  );
  defparam DLX_EXinst_Ker740321.INIT = 16'hFA50;
  X_LUT4 DLX_EXinst_Ker740321 (
    .ADR0(DLX_IDinst_reg_out_B[3]),
    .ADR1(VCC),
    .ADR2(\DLX_EXinst_Mshift__n0023_Sh[23] ),
    .ADR3(\DLX_EXinst_Mshift__n0023_Sh[15] ),
    .O(\DLX_EXinst_N74034/FROM )
  );
  defparam \DLX_EXinst__n0007<27>201 .INIT = 16'hA820;
  X_LUT4 \DLX_EXinst__n0007<27>201  (
    .ADR0(DLX_EXinst__n0080),
    .ADR1(DLX_IDinst_reg_out_B[2]),
    .ADR2(N137518),
    .ADR3(DLX_EXinst_N74034),
    .O(\DLX_EXinst_N74034/GROM )
  );
  X_BUF \DLX_EXinst_N74034/XUSED  (
    .I(\DLX_EXinst_N74034/FROM ),
    .O(DLX_EXinst_N74034)
  );
  X_BUF \DLX_EXinst_N74034/YUSED  (
    .I(\DLX_EXinst_N74034/GROM ),
    .O(CHOICE4974)
  );
  defparam DLX_EXinst_Ker732091.INIT = 16'hFFCC;
  X_LUT4 DLX_EXinst_Ker732091 (
    .ADR0(VCC),
    .ADR1(\DLX_IDinst_Imm[0] ),
    .ADR2(VCC),
    .ADR3(\DLX_IDinst_Imm[1] ),
    .O(\DLX_EXinst_N73211/FROM )
  );
  defparam DLX_EXinst_Ker7534028.INIT = 16'h78F8;
  X_LUT4 DLX_EXinst_Ker7534028 (
    .ADR0(DLX_IDinst_Imm_2_1),
    .ADR1(DLX_IDinst_Imm_3_1),
    .ADR2(\DLX_IDinst_Imm[5] ),
    .ADR3(DLX_EXinst_N73211),
    .O(\DLX_EXinst_N73211/GROM )
  );
  X_BUF \DLX_EXinst_N73211/XUSED  (
    .I(\DLX_EXinst_N73211/FROM ),
    .O(DLX_EXinst_N73211)
  );
  X_BUF \DLX_EXinst_N73211/YUSED  (
    .I(\DLX_EXinst_N73211/GROM ),
    .O(CHOICE1955)
  );
  defparam DLX_EXinst_Ker74449.INIT = 16'hCFC0;
  X_LUT4 DLX_EXinst_Ker74449 (
    .ADR0(VCC),
    .ADR1(\DLX_EXinst_Mshift__n0019_Sh[21] ),
    .ADR2(DLX_IDinst_reg_out_B_3_1),
    .ADR3(N130519),
    .O(\DLX_EXinst_N74451/FROM )
  );
  defparam DLX_EXinst_Ker730811.INIT = 16'hB8B8;
  X_LUT4 DLX_EXinst_Ker730811 (
    .ADR0(\DLX_EXinst_Mshift__n0019_Sh[29] ),
    .ADR1(DLX_IDinst_reg_out_B[3]),
    .ADR2(\DLX_EXinst_Mshift__n0019_Sh[21] ),
    .ADR3(VCC),
    .O(\DLX_EXinst_N74451/GROM )
  );
  X_BUF \DLX_EXinst_N74451/XUSED  (
    .I(\DLX_EXinst_N74451/FROM ),
    .O(DLX_EXinst_N74451)
  );
  X_BUF \DLX_EXinst_N74451/YUSED  (
    .I(\DLX_EXinst_N74451/GROM ),
    .O(DLX_EXinst_N73083)
  );
  defparam DLX_EXinst_Ker731461.INIT = 16'hAAF0;
  X_LUT4 DLX_EXinst_Ker731461 (
    .ADR0(DLX_IDinst_reg_out_A[23]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[21]),
    .ADR3(\DLX_IDinst_Imm[1] ),
    .O(\DLX_EXinst_N73148/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0022_Sh<20>1 .INIT = 16'hFC0C;
  X_LUT4 \DLX_EXinst_Mshift__n0022_Sh<20>1  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N73539),
    .ADR2(DLX_IDinst_Imm_0_1),
    .ADR3(DLX_EXinst_N73148),
    .O(\DLX_EXinst_N73148/GROM )
  );
  X_BUF \DLX_EXinst_N73148/XUSED  (
    .I(\DLX_EXinst_N73148/FROM ),
    .O(DLX_EXinst_N73148)
  );
  X_BUF \DLX_EXinst_N73148/YUSED  (
    .I(\DLX_EXinst_N73148/GROM ),
    .O(\DLX_EXinst_Mshift__n0022_Sh[20] )
  );
  defparam DLX_EXinst_Ker730661.INIT = 16'hEE44;
  X_LUT4 DLX_EXinst_Ker730661 (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(DLX_IDinst_reg_out_A[23]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[25]),
    .O(\DLX_EXinst_N73068/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0019_Sh<22>1 .INIT = 16'hEE44;
  X_LUT4 \DLX_EXinst_Mshift__n0019_Sh<22>1  (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(DLX_EXinst_N73414),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N73068),
    .O(\DLX_EXinst_N73068/GROM )
  );
  X_BUF \DLX_EXinst_N73068/XUSED  (
    .I(\DLX_EXinst_N73068/FROM ),
    .O(DLX_EXinst_N73068)
  );
  X_BUF \DLX_EXinst_N73068/YUSED  (
    .I(\DLX_EXinst_N73068/GROM ),
    .O(\DLX_EXinst_Mshift__n0019_Sh[22] )
  );
  defparam DLX_EXinst_Ker735321.INIT = 16'hE2E2;
  X_LUT4 DLX_EXinst_Ker735321 (
    .ADR0(DLX_IDinst_reg_out_A[18]),
    .ADR1(DLX_IDinst_Imm_1_1),
    .ADR2(DLX_IDinst_reg_out_A[20]),
    .ADR3(VCC),
    .O(\DLX_EXinst_N73534/FROM )
  );
  defparam DLX_EXinst_Ker734021.INIT = 16'hE2E2;
  X_LUT4 DLX_EXinst_Ker734021 (
    .ADR0(DLX_IDinst_reg_out_A[18]),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(DLX_IDinst_reg_out_A[20]),
    .ADR3(VCC),
    .O(\DLX_EXinst_N73534/GROM )
  );
  X_BUF \DLX_EXinst_N73534/XUSED  (
    .I(\DLX_EXinst_N73534/FROM ),
    .O(DLX_EXinst_N73534)
  );
  X_BUF \DLX_EXinst_N73534/YUSED  (
    .I(\DLX_EXinst_N73534/GROM ),
    .O(DLX_EXinst_N73404)
  );
  defparam DLX_EXinst_Ker740271.INIT = 16'hE4E4;
  X_LUT4 DLX_EXinst_Ker740271 (
    .ADR0(DLX_IDinst_reg_out_B[3]),
    .ADR1(\DLX_EXinst_Mshift__n0023_Sh[22] ),
    .ADR2(\DLX_EXinst_Mshift__n0023_Sh[14] ),
    .ADR3(VCC),
    .O(\DLX_EXinst_N74029/FROM )
  );
  defparam \DLX_EXinst__n0007<26>201 .INIT = 16'hE040;
  X_LUT4 \DLX_EXinst__n0007<26>201  (
    .ADR0(DLX_IDinst_reg_out_B[2]),
    .ADR1(N133120),
    .ADR2(DLX_EXinst__n0080),
    .ADR3(DLX_EXinst_N74029),
    .O(\DLX_EXinst_N74029/GROM )
  );
  X_BUF \DLX_EXinst_N74029/XUSED  (
    .I(\DLX_EXinst_N74029/FROM ),
    .O(DLX_EXinst_N74029)
  );
  X_BUF \DLX_EXinst_N74029/YUSED  (
    .I(\DLX_EXinst_N74029/GROM ),
    .O(CHOICE5041)
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<16>1_5_744 .INIT = 16'hAAAC;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<16>1_5_744  (
    .ADR0(DLX_IDinst_current_IR[16]),
    .ADR1(DLX_IFinst_IR_latched[16]),
    .ADR2(DLX_IDinst_counter[0]),
    .ADR3(DLX_IDinst_counter[1]),
    .O(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5/FROM )
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<16>1_1_745 .INIT = 16'hFE02;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<16>1_1_745  (
    .ADR0(DLX_IFinst_IR_latched[16]),
    .ADR1(DLX_IDinst_counter[1]),
    .ADR2(DLX_IDinst_counter[0]),
    .ADR3(DLX_IDinst_current_IR[16]),
    .O(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5/GROM )
  );
  X_BUF \DLX_IDinst_Mmux_IR_latched_Result<16>1_5/XUSED  (
    .I(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5/FROM ),
    .O(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 )
  );
  X_BUF \DLX_IDinst_Mmux_IR_latched_Result<16>1_5/YUSED  (
    .I(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5/GROM ),
    .O(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 )
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<16>1_4_746 .INIT = 16'hCDC8;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<16>1_4_746  (
    .ADR0(DLX_IDinst_counter[0]),
    .ADR1(DLX_IDinst_current_IR[16]),
    .ADR2(DLX_IDinst_counter[1]),
    .ADR3(DLX_IFinst_IR_latched[16]),
    .O(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4/FROM )
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<16>1_2_747 .INIT = 16'hCDC8;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<16>1_2_747  (
    .ADR0(DLX_IDinst_counter[0]),
    .ADR1(DLX_IDinst_current_IR[16]),
    .ADR2(DLX_IDinst_counter[1]),
    .ADR3(DLX_IFinst_IR_latched[16]),
    .O(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4/GROM )
  );
  X_BUF \DLX_IDinst_Mmux_IR_latched_Result<16>1_4/XUSED  (
    .I(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4/FROM ),
    .O(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 )
  );
  X_BUF \DLX_IDinst_Mmux_IR_latched_Result<16>1_4/YUSED  (
    .I(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4/GROM ),
    .O(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 )
  );
  defparam DLX_IDinst_RegFile_28_20_748.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_28_20_748 (
    .I(DLX_IDinst_WB_data_eff[20]),
    .CE(DLX_IDinst__n0606),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_28_20)
  );
  defparam DLX_EXinst_Ker742041.INIT = 16'hCACA;
  X_LUT4 DLX_EXinst_Ker742041 (
    .ADR0(\DLX_EXinst_Mshift__n0021_Sh[23] ),
    .ADR1(\DLX_EXinst_Mshift__n0021_Sh[15] ),
    .ADR2(\DLX_IDinst_Imm[3] ),
    .ADR3(VCC),
    .O(\DLX_EXinst_N74206/FROM )
  );
  defparam \DLX_EXinst__n0007<27>53 .INIT = 16'hC808;
  X_LUT4 \DLX_EXinst__n0007<27>53  (
    .ADR0(N137282),
    .ADR1(DLX_EXinst__n0055),
    .ADR2(\DLX_IDinst_Imm[2] ),
    .ADR3(DLX_EXinst_N74206),
    .O(\DLX_EXinst_N74206/GROM )
  );
  X_BUF \DLX_EXinst_N74206/XUSED  (
    .I(\DLX_EXinst_N74206/FROM ),
    .O(DLX_EXinst_N74206)
  );
  X_BUF \DLX_EXinst_N74206/YUSED  (
    .I(\DLX_EXinst_N74206/GROM ),
    .O(CHOICE4942)
  );
  defparam DLX_EXinst_Ker731561.INIT = 16'hFA0A;
  X_LUT4 DLX_EXinst_Ker731561 (
    .ADR0(\DLX_EXinst_Mshift__n0022_Sh[21] ),
    .ADR1(VCC),
    .ADR2(\DLX_IDinst_Imm[3] ),
    .ADR3(\DLX_EXinst_Mshift__n0022_Sh[29] ),
    .O(\DLX_EXinst_N73158/FROM )
  );
  defparam DLX_EXinst_Ker7464799.INIT = 16'h7340;
  X_LUT4 DLX_EXinst_Ker7464799 (
    .ADR0(DLX_IDinst_Imm_3_1),
    .ADR1(DLX_IDinst_Imm_2_1),
    .ADR2(\DLX_EXinst_Mshift__n0020_Sh[25] ),
    .ADR3(DLX_EXinst_N73158),
    .O(\DLX_EXinst_N73158/GROM )
  );
  X_BUF \DLX_EXinst_N73158/XUSED  (
    .I(\DLX_EXinst_N73158/FROM ),
    .O(DLX_EXinst_N73158)
  );
  X_BUF \DLX_EXinst_N73158/YUSED  (
    .I(\DLX_EXinst_N73158/GROM ),
    .O(CHOICE2972)
  );
  defparam DLX_EXinst_Ker735921.INIT = 16'hF3C0;
  X_LUT4 DLX_EXinst_Ker735921 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(DLX_IDinst_reg_out_A[22]),
    .ADR3(DLX_IDinst_reg_out_A[24]),
    .O(\DLX_EXinst_N73594/FROM )
  );
  defparam DLX_EXinst_Ker734121.INIT = 16'hE2E2;
  X_LUT4 DLX_EXinst_Ker734121 (
    .ADR0(DLX_IDinst_reg_out_A[22]),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(DLX_IDinst_reg_out_A[24]),
    .ADR3(VCC),
    .O(\DLX_EXinst_N73594/GROM )
  );
  X_BUF \DLX_EXinst_N73594/XUSED  (
    .I(\DLX_EXinst_N73594/FROM ),
    .O(DLX_EXinst_N73594)
  );
  X_BUF \DLX_EXinst_N73594/YUSED  (
    .I(\DLX_EXinst_N73594/GROM ),
    .O(DLX_EXinst_N73414)
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<16>1 .INIT = 16'hCDC8;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<16>1  (
    .ADR0(DLX_IDinst_counter[1]),
    .ADR1(DLX_IDinst_current_IR[16]),
    .ADR2(DLX_IDinst_counter[0]),
    .ADR3(DLX_IFinst_IR_latched[16]),
    .O(\DLX_IDinst_current_IR<16>/FROM )
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<16>1_3_749 .INIT = 16'hCCCA;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<16>1_3_749  (
    .ADR0(DLX_IFinst_IR_latched[16]),
    .ADR1(DLX_IDinst_current_IR[16]),
    .ADR2(DLX_IDinst_counter[1]),
    .ADR3(DLX_IDinst_counter[0]),
    .O(\DLX_IDinst_current_IR<16>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<16>/XUSED  (
    .I(\DLX_IDinst_current_IR<16>/FROM ),
    .O(DLX_IDinst_jtarget[16])
  );
  X_BUF \DLX_IDinst_current_IR<16>/YUSED  (
    .I(\DLX_IDinst_current_IR<16>/GROM ),
    .O(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 )
  );
  defparam \DLX_EXinst__n0007<28>142_SW0 .INIT = 16'h0E0A;
  X_LUT4 \DLX_EXinst__n0007<28>142_SW0  (
    .ADR0(CHOICE1295),
    .ADR1(N147520),
    .ADR2(\DLX_IDinst_Imm[4] ),
    .ADR3(CHOICE1291),
    .O(\N164579/FROM )
  );
  defparam \DLX_EXinst__n0007<28>142 .INIT = 16'hFFFE;
  X_LUT4 \DLX_EXinst__n0007<28>142  (
    .ADR0(CHOICE4850),
    .ADR1(CHOICE4866),
    .ADR2(CHOICE4874),
    .ADR3(N164579),
    .O(\N164579/GROM )
  );
  X_BUF \N164579/XUSED  (
    .I(\N164579/FROM ),
    .O(N164579)
  );
  X_BUF \N164579/YUSED  (
    .I(\N164579/GROM ),
    .O(CHOICE4876)
  );
  defparam DLX_EXinst_Ker732371.INIT = 16'hEEEE;
  X_LUT4 DLX_EXinst_Ker732371 (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(DLX_IDinst_reg_out_B[0]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_EXinst_N73239/FROM )
  );
  defparam DLX_EXinst_Ker7516228.INIT = 16'h78F8;
  X_LUT4 DLX_EXinst_Ker7516228 (
    .ADR0(DLX_IDinst_reg_out_B_2_1),
    .ADR1(DLX_IDinst_reg_out_B_3_1),
    .ADR2(DLX_IDinst_reg_out_B[5]),
    .ADR3(DLX_EXinst_N73239),
    .O(\DLX_EXinst_N73239/GROM )
  );
  X_BUF \DLX_EXinst_N73239/XUSED  (
    .I(\DLX_EXinst_N73239/FROM ),
    .O(DLX_EXinst_N73239)
  );
  X_BUF \DLX_EXinst_N73239/YUSED  (
    .I(\DLX_EXinst_N73239/GROM ),
    .O(CHOICE1899)
  );
  defparam DLX_EXinst_Ker730861.INIT = 16'hEE44;
  X_LUT4 DLX_EXinst_Ker730861 (
    .ADR0(DLX_IDinst_reg_out_B[3]),
    .ADR1(\DLX_EXinst_Mshift__n0019_Sh[22] ),
    .ADR2(VCC),
    .ADR3(\DLX_EXinst_Mshift__n0019_Sh[30] ),
    .O(\DLX_EXinst_N73088/FROM )
  );
  defparam DLX_EXinst_Ker7437254.INIT = 16'h5D08;
  X_LUT4 DLX_EXinst_Ker7437254 (
    .ADR0(DLX_IDinst_reg_out_B_2_1),
    .ADR1(\DLX_EXinst_Mshift__n0019_Sh[26] ),
    .ADR2(DLX_IDinst_reg_out_B[3]),
    .ADR3(DLX_EXinst_N73088),
    .O(\DLX_EXinst_N73088/GROM )
  );
  X_BUF \DLX_EXinst_N73088/XUSED  (
    .I(\DLX_EXinst_N73088/FROM ),
    .O(DLX_EXinst_N73088)
  );
  X_BUF \DLX_EXinst_N73088/YUSED  (
    .I(\DLX_EXinst_N73088/GROM ),
    .O(CHOICE3121)
  );
  defparam DLX_EXinst_Ker734971.INIT = 16'hFC30;
  X_LUT4 DLX_EXinst_Ker734971 (
    .ADR0(VCC),
    .ADR1(\DLX_IDinst_Imm[1] ),
    .ADR2(DLX_IDinst_reg_out_A[24]),
    .ADR3(DLX_IDinst_reg_out_A[22]),
    .O(\DLX_EXinst_N73499/FROM )
  );
  defparam DLX_EXinst_Ker734071.INIT = 16'hDD88;
  X_LUT4 DLX_EXinst_Ker734071 (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(DLX_IDinst_reg_out_A[22]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[20]),
    .O(\DLX_EXinst_N73499/GROM )
  );
  X_BUF \DLX_EXinst_N73499/XUSED  (
    .I(\DLX_EXinst_N73499/FROM ),
    .O(DLX_EXinst_N73499)
  );
  X_BUF \DLX_EXinst_N73499/YUSED  (
    .I(\DLX_EXinst_N73499/GROM ),
    .O(DLX_EXinst_N73409)
  );
  defparam DLX_EXinst_Ker733431.INIT = 16'h03BB;
  X_LUT4 DLX_EXinst_Ker733431 (
    .ADR0(DLX_IDinst_IR_opcode_field[0]),
    .ADR1(DLX_IDinst_IR_opcode_field[1]),
    .ADR2(DLX_IDinst_IR_opcode_field[3]),
    .ADR3(DLX_IDinst_IR_opcode_field[2]),
    .O(\DLX_EXinst_N73345/FROM )
  );
  defparam DLX_EXinst_Ker7621813.INIT = 16'hF000;
  X_LUT4 DLX_EXinst_Ker7621813 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_IR_opcode_field[5]),
    .ADR3(DLX_EXinst_N73345),
    .O(\DLX_EXinst_N73345/GROM )
  );
  X_BUF \DLX_EXinst_N73345/XUSED  (
    .I(\DLX_EXinst_N73345/FROM ),
    .O(DLX_EXinst_N73345)
  );
  X_BUF \DLX_EXinst_N73345/YUSED  (
    .I(\DLX_EXinst_N73345/GROM ),
    .O(CHOICE1670)
  );
  defparam DLX_IDinst_RegFile_27_28_750.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_27_28_750 (
    .I(DLX_IDinst_WB_data_eff[28]),
    .CE(DLX_IDinst__n0604),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_27_28)
  );
  defparam DLX_EXinst_Ker735121.INIT = 16'hD8D8;
  X_LUT4 DLX_EXinst_Ker735121 (
    .ADR0(DLX_IDinst_Imm_1_1),
    .ADR1(DLX_IDinst_reg_out_A[12]),
    .ADR2(DLX_IDinst_reg_out_A[10]),
    .ADR3(VCC),
    .O(\DLX_EXinst_N73514/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0022_Sh<9>1 .INIT = 16'hFC30;
  X_LUT4 \DLX_EXinst_Mshift__n0022_Sh<9>1  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_Imm_0_1),
    .ADR2(DLX_EXinst_N73118),
    .ADR3(DLX_EXinst_N73514),
    .O(\DLX_EXinst_N73514/GROM )
  );
  X_BUF \DLX_EXinst_N73514/XUSED  (
    .I(\DLX_EXinst_N73514/FROM ),
    .O(DLX_EXinst_N73514)
  );
  X_BUF \DLX_EXinst_N73514/YUSED  (
    .I(\DLX_EXinst_N73514/GROM ),
    .O(\DLX_EXinst_Mshift__n0022_Sh[9] )
  );
  X_ZERO \DLX_IDinst_RegFile_20_4/LOGIC_ZERO_751  (
    .O(\DLX_IDinst_RegFile_20_4/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_74_752 (
    .IA(\DLX_IDinst_RegFile_20_4/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_20_4/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_133),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_74)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1331.INIT = 16'hDF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1331 (
    .ADR0(DLX_IDinst_jtarget[16]),
    .ADR1(DLX_IDinst_RegFile_21_4),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_53),
    .ADR3(DLX_IDinst_RegFile_20_4),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_133)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1341.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1341 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_54),
    .ADR1(DLX_IDinst_jtarget[16]),
    .ADR2(DLX_IDinst_RegFile_22_4),
    .ADR3(DLX_IDinst_RegFile_23_4),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_134)
  );
  X_BUF \DLX_IDinst_RegFile_20_4/COUTUSED  (
    .I(\DLX_IDinst_RegFile_20_4/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_75)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_75_753 (
    .IA(\DLX_IDinst_RegFile_20_4/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_74),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_134),
    .O(\DLX_IDinst_RegFile_20_4/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_20_4/CYINIT_754  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_73),
    .O(\DLX_IDinst_RegFile_20_4/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_21_0/LOGIC_ZERO_755  (
    .O(\DLX_IDinst_RegFile_21_0/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_522_756 (
    .IA(\DLX_IDinst_RegFile_21_0/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_21_0/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_597),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_522)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_5971.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_5971 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_581),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR2(DLX_IDinst_RegFile_20_0),
    .ADR3(DLX_IDinst_RegFile_21_0),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_597)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_5981.INIT = 16'hFD5D;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_5981 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_582),
    .ADR1(DLX_IDinst_RegFile_22_0),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR3(DLX_IDinst_RegFile_23_0),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_598)
  );
  X_BUF \DLX_IDinst_RegFile_21_0/COUTUSED  (
    .I(\DLX_IDinst_RegFile_21_0/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_523)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_523_757 (
    .IA(\DLX_IDinst_RegFile_21_0/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_522),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_598),
    .O(\DLX_IDinst_RegFile_21_0/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_21_0/CYINIT_758  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_521),
    .O(\DLX_IDinst_RegFile_21_0/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_12_5/LOGIC_ZERO_759  (
    .O(\DLX_IDinst_RegFile_12_5/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_86_760 (
    .IA(\DLX_IDinst_RegFile_12_5/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_12_5/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_145),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_86)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1451.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1451 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_49),
    .ADR1(DLX_IDinst_jtarget[16]),
    .ADR2(DLX_IDinst_RegFile_12_5),
    .ADR3(DLX_IDinst_RegFile_13_5),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_145)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1461.INIT = 16'hE2FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1461 (
    .ADR0(DLX_IDinst_RegFile_14_5),
    .ADR1(DLX_IDinst_jtarget[16]),
    .ADR2(DLX_IDinst_RegFile_15_5),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_50),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_146)
  );
  X_BUF \DLX_IDinst_RegFile_12_5/COUTUSED  (
    .I(\DLX_IDinst_RegFile_12_5/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_87)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_87_761 (
    .IA(\DLX_IDinst_RegFile_12_5/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_86),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_146),
    .O(\DLX_IDinst_RegFile_12_5/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_12_5/CYINIT_762  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_85),
    .O(\DLX_IDinst_RegFile_12_5/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_13_1/LOGIC_ZERO_763  (
    .O(\DLX_IDinst_RegFile_13_1/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_534_764 (
    .IA(\DLX_IDinst_RegFile_13_1/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_13_1/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_609),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_534)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6091.INIT = 16'hE4FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6091 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR1(DLX_IDinst_RegFile_12_1),
    .ADR2(DLX_IDinst_RegFile_13_1),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_577),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_609)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6101.INIT = 16'hE4FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6101 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR1(DLX_IDinst_RegFile_14_1),
    .ADR2(DLX_IDinst_RegFile_15_1),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_578),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_610)
  );
  X_BUF \DLX_IDinst_RegFile_13_1/COUTUSED  (
    .I(\DLX_IDinst_RegFile_13_1/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_535)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_535_765 (
    .IA(\DLX_IDinst_RegFile_13_1/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_534),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_610),
    .O(\DLX_IDinst_RegFile_13_1/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_13_1/CYINIT_766  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_533),
    .O(\DLX_IDinst_RegFile_13_1/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_20_5/LOGIC_ZERO_767  (
    .O(\DLX_IDinst_RegFile_20_5/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_90_768 (
    .IA(\DLX_IDinst_RegFile_20_5/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_20_5/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_149),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_90)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1491.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1491 (
    .ADR0(DLX_IDinst_RegFile_20_5),
    .ADR1(DLX_IDinst_RegFile_21_5),
    .ADR2(DLX_IDinst_jtarget[16]),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_53),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_149)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1501.INIT = 16'hFD5D;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1501 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_54),
    .ADR1(DLX_IDinst_RegFile_22_5),
    .ADR2(DLX_IDinst_jtarget[16]),
    .ADR3(DLX_IDinst_RegFile_23_5),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_150)
  );
  X_BUF \DLX_IDinst_RegFile_20_5/COUTUSED  (
    .I(\DLX_IDinst_RegFile_20_5/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_91)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_91_769 (
    .IA(\DLX_IDinst_RegFile_20_5/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_90),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_150),
    .O(\DLX_IDinst_RegFile_20_5/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_20_5/CYINIT_770  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_89),
    .O(\DLX_IDinst_RegFile_20_5/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_21_1/LOGIC_ZERO_771  (
    .O(\DLX_IDinst_RegFile_21_1/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_538_772 (
    .IA(\DLX_IDinst_RegFile_21_1/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_21_1/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_613),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_538)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6131.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6131 (
    .ADR0(DLX_IDinst_RegFile_20_1),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_581),
    .ADR2(DLX_IDinst_RegFile_21_1),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_613)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6141.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6141 (
    .ADR0(DLX_IDinst_RegFile_22_1),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_582),
    .ADR3(DLX_IDinst_RegFile_23_1),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_614)
  );
  X_BUF \DLX_IDinst_RegFile_21_1/COUTUSED  (
    .I(\DLX_IDinst_RegFile_21_1/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_539)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_539_773 (
    .IA(\DLX_IDinst_RegFile_21_1/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_538),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_614),
    .O(\DLX_IDinst_RegFile_21_1/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_21_1/CYINIT_774  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_537),
    .O(\DLX_IDinst_RegFile_21_1/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_12_6/LOGIC_ZERO_775  (
    .O(\DLX_IDinst_RegFile_12_6/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_102_776 (
    .IA(\DLX_IDinst_RegFile_12_6/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_12_6/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_161),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_102)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1611.INIT = 16'hDF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1611 (
    .ADR0(DLX_IDinst_jtarget[16]),
    .ADR1(DLX_IDinst_RegFile_13_6),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_49),
    .ADR3(DLX_IDinst_RegFile_12_6),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_161)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1621.INIT = 16'hACFF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1621 (
    .ADR0(DLX_IDinst_RegFile_15_6),
    .ADR1(DLX_IDinst_RegFile_14_6),
    .ADR2(DLX_IDinst_jtarget[16]),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_50),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_162)
  );
  X_BUF \DLX_IDinst_RegFile_12_6/COUTUSED  (
    .I(\DLX_IDinst_RegFile_12_6/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_103)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_103_777 (
    .IA(\DLX_IDinst_RegFile_12_6/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_102),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_162),
    .O(\DLX_IDinst_RegFile_12_6/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_12_6/CYINIT_778  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_101),
    .O(\DLX_IDinst_RegFile_12_6/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_13_2/LOGIC_ZERO_779  (
    .O(\DLX_IDinst_RegFile_13_2/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_550_780 (
    .IA(\DLX_IDinst_RegFile_13_2/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_13_2/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_625),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_550)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6251.INIT = 16'hF7B3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6251 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_577),
    .ADR2(DLX_IDinst_RegFile_13_2),
    .ADR3(DLX_IDinst_RegFile_12_2),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_625)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6261.INIT = 16'hB8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6261 (
    .ADR0(DLX_IDinst_RegFile_15_2),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR2(DLX_IDinst_RegFile_14_2),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_578),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_626)
  );
  X_BUF \DLX_IDinst_RegFile_13_2/COUTUSED  (
    .I(\DLX_IDinst_RegFile_13_2/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_551)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_551_781 (
    .IA(\DLX_IDinst_RegFile_13_2/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_550),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_626),
    .O(\DLX_IDinst_RegFile_13_2/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_13_2/CYINIT_782  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_549),
    .O(\DLX_IDinst_RegFile_13_2/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_20_6/LOGIC_ZERO_783  (
    .O(\DLX_IDinst_RegFile_20_6/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_106_784 (
    .IA(\DLX_IDinst_RegFile_20_6/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_20_6/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_165),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_106)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1651.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1651 (
    .ADR0(DLX_IDinst_RegFile_21_6),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_53),
    .ADR2(DLX_IDinst_RegFile_20_6),
    .ADR3(DLX_IDinst_jtarget[16]),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_165)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1661.INIT = 16'hF5DD;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1661 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_54),
    .ADR1(DLX_IDinst_RegFile_22_6),
    .ADR2(DLX_IDinst_RegFile_23_6),
    .ADR3(DLX_IDinst_jtarget[16]),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_166)
  );
  X_BUF \DLX_IDinst_RegFile_20_6/COUTUSED  (
    .I(\DLX_IDinst_RegFile_20_6/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_107)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_107_785 (
    .IA(\DLX_IDinst_RegFile_20_6/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_106),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_166),
    .O(\DLX_IDinst_RegFile_20_6/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_20_6/CYINIT_786  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_105),
    .O(\DLX_IDinst_RegFile_20_6/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_21_2/LOGIC_ZERO_787  (
    .O(\DLX_IDinst_RegFile_21_2/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_554_788 (
    .IA(\DLX_IDinst_RegFile_21_2/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_21_2/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_629),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_554)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6291.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6291 (
    .ADR0(DLX_IDinst_RegFile_20_2),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_581),
    .ADR2(DLX_IDinst_RegFile_21_2),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_629)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6301.INIT = 16'hF5DD;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6301 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_582),
    .ADR1(DLX_IDinst_RegFile_22_2),
    .ADR2(DLX_IDinst_RegFile_23_2),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_630)
  );
  X_BUF \DLX_IDinst_RegFile_21_2/COUTUSED  (
    .I(\DLX_IDinst_RegFile_21_2/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_555)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_555_789 (
    .IA(\DLX_IDinst_RegFile_21_2/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_554),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_630),
    .O(\DLX_IDinst_RegFile_21_2/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_21_2/CYINIT_790  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_553),
    .O(\DLX_IDinst_RegFile_21_2/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_12_7/LOGIC_ZERO_791  (
    .O(\DLX_IDinst_RegFile_12_7/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_118_792 (
    .IA(\DLX_IDinst_RegFile_12_7/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_12_7/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_177),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_118)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1771.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1771 (
    .ADR0(DLX_IDinst_RegFile_12_7),
    .ADR1(DLX_IDinst_RegFile_13_7),
    .ADR2(DLX_IDinst_jtarget[16]),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_49),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_177)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1781.INIT = 16'hBFB3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1781 (
    .ADR0(DLX_IDinst_RegFile_15_7),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_50),
    .ADR2(DLX_IDinst_jtarget[16]),
    .ADR3(DLX_IDinst_RegFile_14_7),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_178)
  );
  X_BUF \DLX_IDinst_RegFile_12_7/COUTUSED  (
    .I(\DLX_IDinst_RegFile_12_7/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_119)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_119_793 (
    .IA(\DLX_IDinst_RegFile_12_7/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_118),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_178),
    .O(\DLX_IDinst_RegFile_12_7/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_12_7/CYINIT_794  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_117),
    .O(\DLX_IDinst_RegFile_12_7/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_13_3/LOGIC_ZERO_795  (
    .O(\DLX_IDinst_RegFile_13_3/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_566_796 (
    .IA(\DLX_IDinst_RegFile_13_3/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_13_3/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_641),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_566)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6411.INIT = 16'hDF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6411 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR1(DLX_IDinst_RegFile_13_3),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_577),
    .ADR3(DLX_IDinst_RegFile_12_3),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_641)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6421.INIT = 16'hAFCF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6421 (
    .ADR0(DLX_IDinst_RegFile_15_3),
    .ADR1(DLX_IDinst_RegFile_14_3),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_578),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_642)
  );
  X_BUF \DLX_IDinst_RegFile_13_3/COUTUSED  (
    .I(\DLX_IDinst_RegFile_13_3/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_567)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_567_797 (
    .IA(\DLX_IDinst_RegFile_13_3/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_566),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_642),
    .O(\DLX_IDinst_RegFile_13_3/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_13_3/CYINIT_798  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_565),
    .O(\DLX_IDinst_RegFile_13_3/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_20_7/LOGIC_ZERO_799  (
    .O(\DLX_IDinst_RegFile_20_7/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_122_800 (
    .IA(\DLX_IDinst_RegFile_20_7/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_20_7/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_181),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_122)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1811.INIT = 16'hFB3B;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1811 (
    .ADR0(DLX_IDinst_RegFile_20_7),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_53),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR3(DLX_IDinst_RegFile_21_7),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_181)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1821.INIT = 16'hF7D5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1821 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_54),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR2(DLX_IDinst_RegFile_23_7),
    .ADR3(DLX_IDinst_RegFile_22_7),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_182)
  );
  X_BUF \DLX_IDinst_RegFile_20_7/COUTUSED  (
    .I(\DLX_IDinst_RegFile_20_7/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_123)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_123_801 (
    .IA(\DLX_IDinst_RegFile_20_7/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_122),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_182),
    .O(\DLX_IDinst_RegFile_20_7/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_20_7/CYINIT_802  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_121),
    .O(\DLX_IDinst_RegFile_20_7/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_21_3/LOGIC_ZERO_803  (
    .O(\DLX_IDinst_RegFile_21_3/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_570_804 (
    .IA(\DLX_IDinst_RegFile_21_3/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_21_3/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_645),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_570)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6451.INIT = 16'hF7B3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6451 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_581),
    .ADR2(DLX_IDinst_RegFile_21_3),
    .ADR3(DLX_IDinst_RegFile_20_3),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_645)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6461.INIT = 16'hDF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6461 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR1(DLX_IDinst_RegFile_23_3),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_582),
    .ADR3(DLX_IDinst_RegFile_22_3),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_646)
  );
  X_BUF \DLX_IDinst_RegFile_21_3/COUTUSED  (
    .I(\DLX_IDinst_RegFile_21_3/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_571)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_571_805 (
    .IA(\DLX_IDinst_RegFile_21_3/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_570),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_646),
    .O(\DLX_IDinst_RegFile_21_3/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_21_3/CYINIT_806  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_569),
    .O(\DLX_IDinst_RegFile_21_3/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_12_8/LOGIC_ZERO_807  (
    .O(\DLX_IDinst_RegFile_12_8/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_134_808 (
    .IA(\DLX_IDinst_RegFile_12_8/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_12_8/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_193),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_134)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1931.INIT = 16'hE4FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1931 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR1(DLX_IDinst_RegFile_12_8),
    .ADR2(DLX_IDinst_RegFile_13_8),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_49),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_193)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1941.INIT = 16'hCFAF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1941 (
    .ADR0(DLX_IDinst_RegFile_14_8),
    .ADR1(DLX_IDinst_RegFile_15_8),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_50),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_194)
  );
  X_BUF \DLX_IDinst_RegFile_12_8/COUTUSED  (
    .I(\DLX_IDinst_RegFile_12_8/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_135)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_135_809 (
    .IA(\DLX_IDinst_RegFile_12_8/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_134),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_194),
    .O(\DLX_IDinst_RegFile_12_8/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_12_8/CYINIT_810  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_133),
    .O(\DLX_IDinst_RegFile_12_8/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_13_4/LOGIC_ZERO_811  (
    .O(\DLX_IDinst_RegFile_13_4/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_582_812 (
    .IA(\DLX_IDinst_RegFile_13_4/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_13_4/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_657),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_582)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6571.INIT = 16'hF7D5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6571 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_577),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR2(DLX_IDinst_RegFile_13_4),
    .ADR3(DLX_IDinst_RegFile_12_4),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_657)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6581.INIT = 16'hB8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6581 (
    .ADR0(DLX_IDinst_RegFile_15_4),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR2(DLX_IDinst_RegFile_14_4),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_578),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_658)
  );
  X_BUF \DLX_IDinst_RegFile_13_4/COUTUSED  (
    .I(\DLX_IDinst_RegFile_13_4/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_583)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_583_813 (
    .IA(\DLX_IDinst_RegFile_13_4/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_582),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_658),
    .O(\DLX_IDinst_RegFile_13_4/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_13_4/CYINIT_814  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_581),
    .O(\DLX_IDinst_RegFile_13_4/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_20_8/LOGIC_ZERO_815  (
    .O(\DLX_IDinst_RegFile_20_8/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_138_816 (
    .IA(\DLX_IDinst_RegFile_20_8/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_20_8/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_197),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_138)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1971.INIT = 16'hE2FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1971 (
    .ADR0(DLX_IDinst_RegFile_20_8),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR2(DLX_IDinst_RegFile_21_8),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_53),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_197)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1981.INIT = 16'hB8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1981 (
    .ADR0(DLX_IDinst_RegFile_23_8),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR2(DLX_IDinst_RegFile_22_8),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_54),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_198)
  );
  X_BUF \DLX_IDinst_RegFile_20_8/COUTUSED  (
    .I(\DLX_IDinst_RegFile_20_8/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_139)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_139_817 (
    .IA(\DLX_IDinst_RegFile_20_8/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_138),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_198),
    .O(\DLX_IDinst_RegFile_20_8/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_20_8/CYINIT_818  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_137),
    .O(\DLX_IDinst_RegFile_20_8/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_21_4/LOGIC_ZERO_819  (
    .O(\DLX_IDinst_RegFile_21_4/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_586_820 (
    .IA(\DLX_IDinst_RegFile_21_4/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_21_4/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_661),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_586)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6611.INIT = 16'hB8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6611 (
    .ADR0(DLX_IDinst_RegFile_21_4),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR2(DLX_IDinst_RegFile_20_4),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_581),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_661)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6621.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6621 (
    .ADR0(DLX_IDinst_RegFile_22_4),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_582),
    .ADR3(DLX_IDinst_RegFile_23_4),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_662)
  );
  X_BUF \DLX_IDinst_RegFile_21_4/COUTUSED  (
    .I(\DLX_IDinst_RegFile_21_4/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_587)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_587_821 (
    .IA(\DLX_IDinst_RegFile_21_4/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_586),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_662),
    .O(\DLX_IDinst_RegFile_21_4/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_21_4/CYINIT_822  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_585),
    .O(\DLX_IDinst_RegFile_21_4/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_30_0/LOGIC_ZERO_823  (
    .O(\DLX_IDinst_RegFile_30_0/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_14_824 (
    .IA(\DLX_IDinst_RegFile_30_0/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_30_0/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_73),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_14)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_731.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_731 (
    .ADR0(DLX_IDinst_RegFile_29_0),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_57),
    .ADR2(DLX_IDinst_RegFile_28_0),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_73)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_741.INIT = 16'hB8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_741 (
    .ADR0(DLX_IDinst_RegFile_31_0),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR2(DLX_IDinst_RegFile_30_0),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_58),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_74)
  );
  X_BUF \DLX_IDinst_RegFile_30_0/COUTUSED  (
    .I(\DLX_IDinst_RegFile_30_0/CYMUXG ),
    .O(DLX_IDinst__n0623[0])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_15 (
    .IA(\DLX_IDinst_RegFile_30_0/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_14),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_74),
    .O(\DLX_IDinst_RegFile_30_0/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_30_0/CYINIT_825  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_13),
    .O(\DLX_IDinst_RegFile_30_0/CYINIT )
  );
  defparam DLX_IDinst_RegFile_26_28_826.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_26_28_826 (
    .I(DLX_IDinst_WB_data_eff[28]),
    .CE(DLX_IDinst__n0602),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_26_28)
  );
  X_ZERO \DLX_IDinst_RegFile_12_9/LOGIC_ZERO_827  (
    .O(\DLX_IDinst_RegFile_12_9/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_150_828 (
    .IA(\DLX_IDinst_RegFile_12_9/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_12_9/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_209),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_150)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2091.INIT = 16'hAFCF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2091 (
    .ADR0(DLX_IDinst_RegFile_13_9),
    .ADR1(DLX_IDinst_RegFile_12_9),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_49),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_209)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2101.INIT = 16'hACFF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2101 (
    .ADR0(DLX_IDinst_RegFile_15_9),
    .ADR1(DLX_IDinst_RegFile_14_9),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_50),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_210)
  );
  X_BUF \DLX_IDinst_RegFile_12_9/COUTUSED  (
    .I(\DLX_IDinst_RegFile_12_9/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_151)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_151_829 (
    .IA(\DLX_IDinst_RegFile_12_9/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_150),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_210),
    .O(\DLX_IDinst_RegFile_12_9/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_12_9/CYINIT_830  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_149),
    .O(\DLX_IDinst_RegFile_12_9/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_13_5/LOGIC_ZERO_831  (
    .O(\DLX_IDinst_RegFile_13_5/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_598_832 (
    .IA(\DLX_IDinst_RegFile_13_5/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_13_5/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_673),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_598)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6731.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6731 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_577),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR2(DLX_IDinst_RegFile_12_5),
    .ADR3(DLX_IDinst_RegFile_13_5),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_673)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6741.INIT = 16'hE2FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6741 (
    .ADR0(DLX_IDinst_RegFile_14_5),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR2(DLX_IDinst_RegFile_15_5),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_578),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_674)
  );
  X_BUF \DLX_IDinst_RegFile_13_5/COUTUSED  (
    .I(\DLX_IDinst_RegFile_13_5/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_599)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_599_833 (
    .IA(\DLX_IDinst_RegFile_13_5/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_598),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_674),
    .O(\DLX_IDinst_RegFile_13_5/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_13_5/CYINIT_834  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_597),
    .O(\DLX_IDinst_RegFile_13_5/CYINIT )
  );
  defparam DLX_IDinst_RegFile_27_12_835.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_27_12_835 (
    .I(DLX_IDinst_WB_data_eff[12]),
    .CE(DLX_IDinst__n0604),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_27_12)
  );
  X_ZERO \DLX_IDinst_RegFile_20_9/LOGIC_ZERO_836  (
    .O(\DLX_IDinst_RegFile_20_9/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_154_837 (
    .IA(\DLX_IDinst_RegFile_20_9/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_20_9/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_213),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_154)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2131.INIT = 16'hF5DD;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2131 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_53),
    .ADR1(DLX_IDinst_RegFile_20_9),
    .ADR2(DLX_IDinst_RegFile_21_9),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_213)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2141.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2141 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_54),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR2(DLX_IDinst_RegFile_22_9),
    .ADR3(DLX_IDinst_RegFile_23_9),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_214)
  );
  X_BUF \DLX_IDinst_RegFile_20_9/COUTUSED  (
    .I(\DLX_IDinst_RegFile_20_9/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_155)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_155_838 (
    .IA(\DLX_IDinst_RegFile_20_9/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_154),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_214),
    .O(\DLX_IDinst_RegFile_20_9/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_20_9/CYINIT_839  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_153),
    .O(\DLX_IDinst_RegFile_20_9/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_21_5/LOGIC_ZERO_840  (
    .O(\DLX_IDinst_RegFile_21_5/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_602_841 (
    .IA(\DLX_IDinst_RegFile_21_5/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_21_5/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_677),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_602)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6771.INIT = 16'hF7B3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6771 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_581),
    .ADR2(DLX_IDinst_RegFile_21_5),
    .ADR3(DLX_IDinst_RegFile_20_5),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_677)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6781.INIT = 16'hB8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6781 (
    .ADR0(DLX_IDinst_RegFile_23_5),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR2(DLX_IDinst_RegFile_22_5),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_582),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_678)
  );
  X_BUF \DLX_IDinst_RegFile_21_5/COUTUSED  (
    .I(\DLX_IDinst_RegFile_21_5/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_603)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_603_842 (
    .IA(\DLX_IDinst_RegFile_21_5/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_602),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_678),
    .O(\DLX_IDinst_RegFile_21_5/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_21_5/CYINIT_843  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_601),
    .O(\DLX_IDinst_RegFile_21_5/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_30_1/LOGIC_ZERO_844  (
    .O(\DLX_IDinst_RegFile_30_1/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_30_845 (
    .IA(\DLX_IDinst_RegFile_30_1/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_30_1/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_89),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_30)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_891.INIT = 16'hBFB3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_891 (
    .ADR0(DLX_IDinst_RegFile_29_1),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_57),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR3(DLX_IDinst_RegFile_28_1),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_89)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_901.INIT = 16'hFB3B;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_901 (
    .ADR0(DLX_IDinst_RegFile_30_1),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_58),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR3(DLX_IDinst_RegFile_31_1),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_90)
  );
  X_BUF \DLX_IDinst_RegFile_30_1/COUTUSED  (
    .I(\DLX_IDinst_RegFile_30_1/CYMUXG ),
    .O(DLX_IDinst__n0623[1])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_31 (
    .IA(\DLX_IDinst_RegFile_30_1/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_30),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_90),
    .O(\DLX_IDinst_RegFile_30_1/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_30_1/CYINIT_846  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_29),
    .O(\DLX_IDinst_RegFile_30_1/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_13_6/LOGIC_ZERO_847  (
    .O(\DLX_IDinst_RegFile_13_6/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_614_848 (
    .IA(\DLX_IDinst_RegFile_13_6/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_13_6/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_689),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_614)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6891.INIT = 16'hDFD5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6891 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_577),
    .ADR1(DLX_IDinst_RegFile_13_6),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR3(DLX_IDinst_RegFile_12_6),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_689)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6901.INIT = 16'hFB3B;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6901 (
    .ADR0(DLX_IDinst_RegFile_14_6),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_578),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR3(DLX_IDinst_RegFile_15_6),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_690)
  );
  X_BUF \DLX_IDinst_RegFile_13_6/COUTUSED  (
    .I(\DLX_IDinst_RegFile_13_6/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_615)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_615_849 (
    .IA(\DLX_IDinst_RegFile_13_6/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_614),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_690),
    .O(\DLX_IDinst_RegFile_13_6/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_13_6/CYINIT_850  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_613),
    .O(\DLX_IDinst_RegFile_13_6/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_21_6/LOGIC_ZERO_851  (
    .O(\DLX_IDinst_RegFile_21_6/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_618_852 (
    .IA(\DLX_IDinst_RegFile_21_6/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_21_6/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_693),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_618)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6931.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6931 (
    .ADR0(DLX_IDinst_RegFile_20_6),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_581),
    .ADR2(DLX_IDinst_RegFile_21_6),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_693)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6941.INIT = 16'hCFAF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6941 (
    .ADR0(DLX_IDinst_RegFile_22_6),
    .ADR1(DLX_IDinst_RegFile_23_6),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_582),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_694)
  );
  X_BUF \DLX_IDinst_RegFile_21_6/COUTUSED  (
    .I(\DLX_IDinst_RegFile_21_6/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_619)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_619_853 (
    .IA(\DLX_IDinst_RegFile_21_6/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_618),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_694),
    .O(\DLX_IDinst_RegFile_21_6/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_21_6/CYINIT_854  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_617),
    .O(\DLX_IDinst_RegFile_21_6/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_30_2/LOGIC_ZERO_855  (
    .O(\DLX_IDinst_RegFile_30_2/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_46_856 (
    .IA(\DLX_IDinst_RegFile_30_2/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_30_2/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_105),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_46)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1051.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1051 (
    .ADR0(DLX_IDinst_RegFile_29_2),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_57),
    .ADR2(DLX_IDinst_RegFile_28_2),
    .ADR3(DLX_IDinst_jtarget[16]),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_105)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1061.INIT = 16'hE2FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1061 (
    .ADR0(DLX_IDinst_RegFile_30_2),
    .ADR1(DLX_IDinst_jtarget[16]),
    .ADR2(DLX_IDinst_RegFile_31_2),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_58),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_106)
  );
  X_BUF \DLX_IDinst_RegFile_30_2/COUTUSED  (
    .I(\DLX_IDinst_RegFile_30_2/CYMUXG ),
    .O(DLX_IDinst__n0623[2])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_47 (
    .IA(\DLX_IDinst_RegFile_30_2/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_46),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_106),
    .O(\DLX_IDinst_RegFile_30_2/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_30_2/CYINIT_857  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_45),
    .O(\DLX_IDinst_RegFile_30_2/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_13_7/LOGIC_ZERO_858  (
    .O(\DLX_IDinst_RegFile_13_7/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_630_859 (
    .IA(\DLX_IDinst_RegFile_13_7/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_13_7/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_705),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_630)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7051.INIT = 16'hF7D5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7051 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_577),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR2(DLX_IDinst_RegFile_13_7),
    .ADR3(DLX_IDinst_RegFile_12_7),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_705)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7061.INIT = 16'hE4FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7061 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR1(DLX_IDinst_RegFile_14_7),
    .ADR2(DLX_IDinst_RegFile_15_7),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_578),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_706)
  );
  X_BUF \DLX_IDinst_RegFile_13_7/COUTUSED  (
    .I(\DLX_IDinst_RegFile_13_7/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_631)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_631_860 (
    .IA(\DLX_IDinst_RegFile_13_7/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_630),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_706),
    .O(\DLX_IDinst_RegFile_13_7/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_13_7/CYINIT_861  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_629),
    .O(\DLX_IDinst_RegFile_13_7/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_21_7/LOGIC_ZERO_862  (
    .O(\DLX_IDinst_RegFile_21_7/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_634_863 (
    .IA(\DLX_IDinst_RegFile_21_7/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_21_7/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_709),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_634)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7091.INIT = 16'hBFB3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7091 (
    .ADR0(DLX_IDinst_RegFile_21_7),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_581),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR3(DLX_IDinst_RegFile_20_7),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_709)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7101.INIT = 16'hFD5D;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7101 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_582),
    .ADR1(DLX_IDinst_RegFile_22_7),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR3(DLX_IDinst_RegFile_23_7),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_710)
  );
  X_BUF \DLX_IDinst_RegFile_21_7/COUTUSED  (
    .I(\DLX_IDinst_RegFile_21_7/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_635)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_635_864 (
    .IA(\DLX_IDinst_RegFile_21_7/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_634),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_710),
    .O(\DLX_IDinst_RegFile_21_7/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_21_7/CYINIT_865  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_633),
    .O(\DLX_IDinst_RegFile_21_7/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_30_3/LOGIC_ZERO_866  (
    .O(\DLX_IDinst_RegFile_30_3/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_62_867 (
    .IA(\DLX_IDinst_RegFile_30_3/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_30_3/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_121),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_62)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1211.INIT = 16'hACFF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1211 (
    .ADR0(DLX_IDinst_RegFile_29_3),
    .ADR1(DLX_IDinst_RegFile_28_3),
    .ADR2(DLX_IDinst_jtarget[16]),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_57),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_121)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1221.INIT = 16'hAFCF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1221 (
    .ADR0(DLX_IDinst_RegFile_31_3),
    .ADR1(DLX_IDinst_RegFile_30_3),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_58),
    .ADR3(DLX_IDinst_jtarget[16]),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_122)
  );
  X_BUF \DLX_IDinst_RegFile_30_3/COUTUSED  (
    .I(\DLX_IDinst_RegFile_30_3/CYMUXG ),
    .O(DLX_IDinst__n0623[3])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_63 (
    .IA(\DLX_IDinst_RegFile_30_3/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_62),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_122),
    .O(\DLX_IDinst_RegFile_30_3/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_30_3/CYINIT_868  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_61),
    .O(\DLX_IDinst_RegFile_30_3/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_13_8/LOGIC_ZERO_869  (
    .O(\DLX_IDinst_RegFile_13_8/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_646_870 (
    .IA(\DLX_IDinst_RegFile_13_8/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_13_8/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_721),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_646)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7211.INIT = 16'hB8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7211 (
    .ADR0(DLX_IDinst_RegFile_13_8),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR2(DLX_IDinst_RegFile_12_8),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_577),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_721)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7221.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7221 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR1(DLX_IDinst_RegFile_14_8),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_578),
    .ADR3(DLX_IDinst_RegFile_15_8),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_722)
  );
  X_BUF \DLX_IDinst_RegFile_13_8/COUTUSED  (
    .I(\DLX_IDinst_RegFile_13_8/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_647)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_647_871 (
    .IA(\DLX_IDinst_RegFile_13_8/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_646),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_722),
    .O(\DLX_IDinst_RegFile_13_8/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_13_8/CYINIT_872  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_645),
    .O(\DLX_IDinst_RegFile_13_8/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_21_8/LOGIC_ZERO_873  (
    .O(\DLX_IDinst_RegFile_21_8/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_650_874 (
    .IA(\DLX_IDinst_RegFile_21_8/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_21_8/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_725),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_650)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7251.INIT = 16'hD8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7251 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR1(DLX_IDinst_RegFile_21_8),
    .ADR2(DLX_IDinst_RegFile_20_8),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_581),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_725)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7261.INIT = 16'hBF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7261 (
    .ADR0(DLX_IDinst_RegFile_23_8),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_582),
    .ADR3(DLX_IDinst_RegFile_22_8),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_726)
  );
  X_BUF \DLX_IDinst_RegFile_21_8/COUTUSED  (
    .I(\DLX_IDinst_RegFile_21_8/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_651)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_651_875 (
    .IA(\DLX_IDinst_RegFile_21_8/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_650),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_726),
    .O(\DLX_IDinst_RegFile_21_8/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_21_8/CYINIT_876  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_649),
    .O(\DLX_IDinst_RegFile_21_8/CYINIT )
  );
  defparam DLX_IDinst_RegFile_27_20_877.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_27_20_877 (
    .I(DLX_IDinst_WB_data_eff[20]),
    .CE(DLX_IDinst__n0604),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_27_20)
  );
  X_ZERO \DLX_IDinst_RegFile_30_4/LOGIC_ZERO_878  (
    .O(\DLX_IDinst_RegFile_30_4/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_78_879 (
    .IA(\DLX_IDinst_RegFile_30_4/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_30_4/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_137),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_78)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1371.INIT = 16'hF7B3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1371 (
    .ADR0(DLX_IDinst_jtarget[16]),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_57),
    .ADR2(DLX_IDinst_RegFile_29_4),
    .ADR3(DLX_IDinst_RegFile_28_4),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_137)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1381.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1381 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_58),
    .ADR1(DLX_IDinst_jtarget[16]),
    .ADR2(DLX_IDinst_RegFile_30_4),
    .ADR3(DLX_IDinst_RegFile_31_4),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_138)
  );
  X_BUF \DLX_IDinst_RegFile_30_4/COUTUSED  (
    .I(\DLX_IDinst_RegFile_30_4/CYMUXG ),
    .O(DLX_IDinst__n0623[4])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_79 (
    .IA(\DLX_IDinst_RegFile_30_4/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_78),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_138),
    .O(\DLX_IDinst_RegFile_30_4/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_30_4/CYINIT_880  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_77),
    .O(\DLX_IDinst_RegFile_30_4/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_31_0/LOGIC_ZERO_881  (
    .O(\DLX_IDinst_RegFile_31_0/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_526_882 (
    .IA(\DLX_IDinst_RegFile_31_0/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_31_0/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_601),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_526)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6011.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6011 (
    .ADR0(DLX_IDinst_RegFile_28_0),
    .ADR1(DLX_IDinst_RegFile_29_0),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_585),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_601)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6021.INIT = 16'hBFB3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6021 (
    .ADR0(DLX_IDinst_RegFile_31_0),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_586),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR3(DLX_IDinst_RegFile_30_0),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_602)
  );
  X_BUF \DLX_IDinst_RegFile_31_0/COUTUSED  (
    .I(\DLX_IDinst_RegFile_31_0/CYMUXG ),
    .O(DLX_IDinst__n0620[0])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_527 (
    .IA(\DLX_IDinst_RegFile_31_0/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_526),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_602),
    .O(\DLX_IDinst_RegFile_31_0/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_31_0/CYINIT_883  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_525),
    .O(\DLX_IDinst_RegFile_31_0/CYINIT )
  );
  defparam vga_top_vga1_Ker112929_SW0.INIT = 16'hFFBF;
  X_LUT4 vga_top_vga1_Ker112929_SW0 (
    .ADR0(vga_top_vga1_hcounter[8]),
    .ADR1(vga_top_vga1_hcounter[3]),
    .ADR2(vga_top_vga1_hcounter[0]),
    .ADR3(vga_top_vga1_hcounter[9]),
    .O(\N136748/FROM )
  );
  defparam vga_top_vga1__n00131.INIT = 16'h8080;
  X_LUT4 vga_top_vga1__n00131 (
    .ADR0(vga_top_vga1_hcounter[0]),
    .ADR1(vga_top_vga1__n0037),
    .ADR2(vga_top_vga1_hcounter[1]),
    .ADR3(VCC),
    .O(\N136748/GROM )
  );
  X_BUF \N136748/XUSED  (
    .I(\N136748/FROM ),
    .O(N136748)
  );
  X_BUF \N136748/YUSED  (
    .I(\N136748/GROM ),
    .O(vga_top_vga1__n0013)
  );
  X_ZERO \DLX_IDinst_RegFile_13_9/LOGIC_ZERO_884  (
    .O(\DLX_IDinst_RegFile_13_9/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_662_885 (
    .IA(\DLX_IDinst_RegFile_13_9/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_13_9/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_737),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_662)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7371.INIT = 16'hE2FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7371 (
    .ADR0(DLX_IDinst_RegFile_12_9),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR2(DLX_IDinst_RegFile_13_9),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_577),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_737)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7381.INIT = 16'hF7D5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7381 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_578),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR2(DLX_IDinst_RegFile_15_9),
    .ADR3(DLX_IDinst_RegFile_14_9),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_738)
  );
  X_BUF \DLX_IDinst_RegFile_13_9/COUTUSED  (
    .I(\DLX_IDinst_RegFile_13_9/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_663)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_663_886 (
    .IA(\DLX_IDinst_RegFile_13_9/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_662),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_738),
    .O(\DLX_IDinst_RegFile_13_9/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_13_9/CYINIT_887  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_661),
    .O(\DLX_IDinst_RegFile_13_9/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_21_9/LOGIC_ZERO_888  (
    .O(\DLX_IDinst_RegFile_21_9/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_666_889 (
    .IA(\DLX_IDinst_RegFile_21_9/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_21_9/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_741),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_666)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7411.INIT = 16'hE2FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7411 (
    .ADR0(DLX_IDinst_RegFile_20_9),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR2(DLX_IDinst_RegFile_21_9),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_581),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_741)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7421.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7421 (
    .ADR0(DLX_IDinst_RegFile_22_9),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_582),
    .ADR2(DLX_IDinst_RegFile_23_9),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_742)
  );
  X_BUF \DLX_IDinst_RegFile_21_9/COUTUSED  (
    .I(\DLX_IDinst_RegFile_21_9/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_667)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_667_890 (
    .IA(\DLX_IDinst_RegFile_21_9/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_666),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_742),
    .O(\DLX_IDinst_RegFile_21_9/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_21_9/CYINIT_891  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_665),
    .O(\DLX_IDinst_RegFile_21_9/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_30_5/LOGIC_ZERO_892  (
    .O(\DLX_IDinst_RegFile_30_5/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_94_893 (
    .IA(\DLX_IDinst_RegFile_30_5/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_30_5/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_153),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_94)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1531.INIT = 16'hBF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1531 (
    .ADR0(DLX_IDinst_RegFile_29_5),
    .ADR1(DLX_IDinst_jtarget[16]),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_57),
    .ADR3(DLX_IDinst_RegFile_28_5),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_153)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1541.INIT = 16'hB8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1541 (
    .ADR0(DLX_IDinst_RegFile_31_5),
    .ADR1(DLX_IDinst_jtarget[16]),
    .ADR2(DLX_IDinst_RegFile_30_5),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_58),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_154)
  );
  X_BUF \DLX_IDinst_RegFile_30_5/COUTUSED  (
    .I(\DLX_IDinst_RegFile_30_5/CYMUXG ),
    .O(DLX_IDinst__n0623[5])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_95 (
    .IA(\DLX_IDinst_RegFile_30_5/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_94),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_154),
    .O(\DLX_IDinst_RegFile_30_5/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_30_5/CYINIT_894  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_93),
    .O(\DLX_IDinst_RegFile_30_5/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_31_1/LOGIC_ZERO_895  (
    .O(\DLX_IDinst_RegFile_31_1/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_542_896 (
    .IA(\DLX_IDinst_RegFile_31_1/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_31_1/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_617),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_542)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6171.INIT = 16'hF7D5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6171 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_585),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR2(DLX_IDinst_RegFile_29_1),
    .ADR3(DLX_IDinst_RegFile_28_1),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_617)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6181.INIT = 16'hF5DD;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6181 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_586),
    .ADR1(DLX_IDinst_RegFile_30_1),
    .ADR2(DLX_IDinst_RegFile_31_1),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_618)
  );
  X_BUF \DLX_IDinst_RegFile_31_1/COUTUSED  (
    .I(\DLX_IDinst_RegFile_31_1/CYMUXG ),
    .O(DLX_IDinst__n0620[1])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_543 (
    .IA(\DLX_IDinst_RegFile_31_1/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_542),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_618),
    .O(\DLX_IDinst_RegFile_31_1/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_31_1/CYINIT_897  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_541),
    .O(\DLX_IDinst_RegFile_31_1/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_30_6/LOGIC_ZERO_898  (
    .O(\DLX_IDinst_RegFile_30_6/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_110_899 (
    .IA(\DLX_IDinst_RegFile_30_6/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_30_6/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_169),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_110)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1691.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1691 (
    .ADR0(DLX_IDinst_RegFile_28_6),
    .ADR1(DLX_IDinst_jtarget[16]),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_57),
    .ADR3(DLX_IDinst_RegFile_29_6),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_169)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1701.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1701 (
    .ADR0(DLX_IDinst_jtarget[16]),
    .ADR1(DLX_IDinst_RegFile_30_6),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_58),
    .ADR3(DLX_IDinst_RegFile_31_6),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_170)
  );
  X_BUF \DLX_IDinst_RegFile_30_6/COUTUSED  (
    .I(\DLX_IDinst_RegFile_30_6/CYMUXG ),
    .O(DLX_IDinst__n0623[6])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_111 (
    .IA(\DLX_IDinst_RegFile_30_6/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_110),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_170),
    .O(\DLX_IDinst_RegFile_30_6/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_30_6/CYINIT_900  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_109),
    .O(\DLX_IDinst_RegFile_30_6/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_31_2/LOGIC_ZERO_901  (
    .O(\DLX_IDinst_RegFile_31_2/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_558_902 (
    .IA(\DLX_IDinst_RegFile_31_2/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_31_2/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_633),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_558)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6331.INIT = 16'hFB3B;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6331 (
    .ADR0(DLX_IDinst_RegFile_28_2),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_585),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR3(DLX_IDinst_RegFile_29_2),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_633)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6341.INIT = 16'hDF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6341 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR1(DLX_IDinst_RegFile_31_2),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_586),
    .ADR3(DLX_IDinst_RegFile_30_2),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_634)
  );
  X_BUF \DLX_IDinst_RegFile_31_2/COUTUSED  (
    .I(\DLX_IDinst_RegFile_31_2/CYMUXG ),
    .O(DLX_IDinst__n0620[2])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_559 (
    .IA(\DLX_IDinst_RegFile_31_2/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_558),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_634),
    .O(\DLX_IDinst_RegFile_31_2/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_31_2/CYINIT_903  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_557),
    .O(\DLX_IDinst_RegFile_31_2/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_30_7/LOGIC_ZERO_904  (
    .O(\DLX_IDinst_RegFile_30_7/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_126_905 (
    .IA(\DLX_IDinst_RegFile_30_7/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_30_7/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_185),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_126)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1851.INIT = 16'hB8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1851 (
    .ADR0(DLX_IDinst_RegFile_29_7),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR2(DLX_IDinst_RegFile_28_7),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_57),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_185)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1861.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1861 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_58),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR2(DLX_IDinst_RegFile_30_7),
    .ADR3(DLX_IDinst_RegFile_31_7),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_186)
  );
  X_BUF \DLX_IDinst_RegFile_30_7/COUTUSED  (
    .I(\DLX_IDinst_RegFile_30_7/CYMUXG ),
    .O(DLX_IDinst__n0623[7])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_127 (
    .IA(\DLX_IDinst_RegFile_30_7/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_126),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_186),
    .O(\DLX_IDinst_RegFile_30_7/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_30_7/CYINIT_906  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_125),
    .O(\DLX_IDinst_RegFile_30_7/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_31_3/LOGIC_ZERO_907  (
    .O(\DLX_IDinst_RegFile_31_3/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_574_908 (
    .IA(\DLX_IDinst_RegFile_31_3/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_31_3/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_649),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_574)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6491.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6491 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_585),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR2(DLX_IDinst_RegFile_28_3),
    .ADR3(DLX_IDinst_RegFile_29_3),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_649)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6501.INIT = 16'hF5DD;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6501 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_586),
    .ADR1(DLX_IDinst_RegFile_30_3),
    .ADR2(DLX_IDinst_RegFile_31_3),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_650)
  );
  X_BUF \DLX_IDinst_RegFile_31_3/COUTUSED  (
    .I(\DLX_IDinst_RegFile_31_3/CYMUXG ),
    .O(DLX_IDinst__n0620[3])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_575 (
    .IA(\DLX_IDinst_RegFile_31_3/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_574),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_650),
    .O(\DLX_IDinst_RegFile_31_3/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_31_3/CYINIT_909  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_573),
    .O(\DLX_IDinst_RegFile_31_3/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_16_0/LOGIC_ZERO_910  (
    .O(\DLX_IDinst_RegFile_16_0/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_8_911 (
    .IA(\DLX_IDinst_RegFile_16_0/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_16_0/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_67),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_8)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_671.INIT = 16'hFB73;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_671 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_51),
    .ADR2(DLX_IDinst_RegFile_16_0),
    .ADR3(DLX_IDinst_RegFile_17_0),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_67)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_681.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_681 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR1(DLX_IDinst_RegFile_18_0),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_52),
    .ADR3(DLX_IDinst_RegFile_19_0),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_68)
  );
  X_BUF \DLX_IDinst_RegFile_16_0/COUTUSED  (
    .I(\DLX_IDinst_RegFile_16_0/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_9)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_9_912 (
    .IA(\DLX_IDinst_RegFile_16_0/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_8),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_68),
    .O(\DLX_IDinst_RegFile_16_0/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_16_0/CYINIT_913  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_7),
    .O(\DLX_IDinst_RegFile_16_0/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_24_0/LOGIC_ZERO_914  (
    .O(\DLX_IDinst_RegFile_24_0/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_12_915 (
    .IA(\DLX_IDinst_RegFile_24_0/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_24_0/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_71),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_12)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_711.INIT = 16'hE4FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_711 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR1(DLX_IDinst_RegFile_24_0),
    .ADR2(DLX_IDinst_RegFile_25_0),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_55),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_71)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_721.INIT = 16'hD8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_721 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR1(DLX_IDinst_RegFile_27_0),
    .ADR2(DLX_IDinst_RegFile_26_0),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_56),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_72)
  );
  X_BUF \DLX_IDinst_RegFile_24_0/COUTUSED  (
    .I(\DLX_IDinst_RegFile_24_0/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_13)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_13_916 (
    .IA(\DLX_IDinst_RegFile_24_0/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_12),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_72),
    .O(\DLX_IDinst_RegFile_24_0/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_24_0/CYINIT_917  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_11),
    .O(\DLX_IDinst_RegFile_24_0/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_30_8/LOGIC_ZERO_918  (
    .O(\DLX_IDinst_RegFile_30_8/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_142_919 (
    .IA(\DLX_IDinst_RegFile_30_8/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_30_8/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_201),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_142)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2011.INIT = 16'hDFD5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2011 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_57),
    .ADR1(DLX_IDinst_RegFile_29_8),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR3(DLX_IDinst_RegFile_28_8),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_201)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2021.INIT = 16'hE2FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2021 (
    .ADR0(DLX_IDinst_RegFile_30_8),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR2(DLX_IDinst_RegFile_31_8),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_58),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_202)
  );
  X_BUF \DLX_IDinst_RegFile_30_8/COUTUSED  (
    .I(\DLX_IDinst_RegFile_30_8/CYMUXG ),
    .O(DLX_IDinst__n0623[8])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_143 (
    .IA(\DLX_IDinst_RegFile_30_8/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_142),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_202),
    .O(\DLX_IDinst_RegFile_30_8/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_30_8/CYINIT_920  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_141),
    .O(\DLX_IDinst_RegFile_30_8/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_31_4/LOGIC_ZERO_921  (
    .O(\DLX_IDinst_RegFile_31_4/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_590_922 (
    .IA(\DLX_IDinst_RegFile_31_4/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_31_4/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_665),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_590)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6651.INIT = 16'hD8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6651 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR1(DLX_IDinst_RegFile_29_4),
    .ADR2(DLX_IDinst_RegFile_28_4),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_585),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_665)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6661.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6661 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_586),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR2(DLX_IDinst_RegFile_30_4),
    .ADR3(DLX_IDinst_RegFile_31_4),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_666)
  );
  X_BUF \DLX_IDinst_RegFile_31_4/COUTUSED  (
    .I(\DLX_IDinst_RegFile_31_4/CYMUXG ),
    .O(DLX_IDinst__n0620[4])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_591 (
    .IA(\DLX_IDinst_RegFile_31_4/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_590),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_666),
    .O(\DLX_IDinst_RegFile_31_4/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_31_4/CYINIT_923  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_589),
    .O(\DLX_IDinst_RegFile_31_4/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_16_1/LOGIC_ZERO_924  (
    .O(\DLX_IDinst_RegFile_16_1/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_24_925 (
    .IA(\DLX_IDinst_RegFile_16_1/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_16_1/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_83),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_24)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_831.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_831 (
    .ADR0(DLX_IDinst_RegFile_17_1),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_51),
    .ADR2(DLX_IDinst_RegFile_16_1),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_83)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_841.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_841 (
    .ADR0(DLX_IDinst_RegFile_18_1),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_52),
    .ADR2(DLX_IDinst_RegFile_19_1),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_84)
  );
  X_BUF \DLX_IDinst_RegFile_16_1/COUTUSED  (
    .I(\DLX_IDinst_RegFile_16_1/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_25)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_25_926 (
    .IA(\DLX_IDinst_RegFile_16_1/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_24),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_84),
    .O(\DLX_IDinst_RegFile_16_1/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_16_1/CYINIT_927  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_23),
    .O(\DLX_IDinst_RegFile_16_1/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_24_1/LOGIC_ZERO_928  (
    .O(\DLX_IDinst_RegFile_24_1/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_28_929 (
    .IA(\DLX_IDinst_RegFile_24_1/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_24_1/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_87),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_28)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_871.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_871 (
    .ADR0(DLX_IDinst_RegFile_24_1),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_55),
    .ADR3(DLX_IDinst_RegFile_25_1),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_87)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_881.INIT = 16'hACFF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_881 (
    .ADR0(DLX_IDinst_RegFile_27_1),
    .ADR1(DLX_IDinst_RegFile_26_1),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_56),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_88)
  );
  X_BUF \DLX_IDinst_RegFile_24_1/COUTUSED  (
    .I(\DLX_IDinst_RegFile_24_1/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_29)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_29_930 (
    .IA(\DLX_IDinst_RegFile_24_1/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_28),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_88),
    .O(\DLX_IDinst_RegFile_24_1/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_24_1/CYINIT_931  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_27),
    .O(\DLX_IDinst_RegFile_24_1/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_30_9/LOGIC_ZERO_932  (
    .O(\DLX_IDinst_RegFile_30_9/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_158_933 (
    .IA(\DLX_IDinst_RegFile_30_9/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_30_9/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_217),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_158)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2171.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2171 (
    .ADR0(DLX_IDinst_RegFile_28_9),
    .ADR1(DLX_IDinst_RegFile_29_9),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_57),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_217)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2181.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2181 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_58),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR2(DLX_IDinst_RegFile_30_9),
    .ADR3(DLX_IDinst_RegFile_31_9),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_218)
  );
  X_BUF \DLX_IDinst_RegFile_30_9/COUTUSED  (
    .I(\DLX_IDinst_RegFile_30_9/CYMUXG ),
    .O(DLX_IDinst__n0623[9])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_159 (
    .IA(\DLX_IDinst_RegFile_30_9/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_158),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_218),
    .O(\DLX_IDinst_RegFile_30_9/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_30_9/CYINIT_934  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_157),
    .O(\DLX_IDinst_RegFile_30_9/CYINIT )
  );
  defparam DLX_IDinst_RegFile_18_29_935.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_18_29_935 (
    .I(DLX_IDinst_WB_data_eff[29]),
    .CE(DLX_IDinst__n0586),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_18_29)
  );
  X_ZERO \DLX_IDinst_RegFile_31_5/LOGIC_ZERO_936  (
    .O(\DLX_IDinst_RegFile_31_5/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_606_937 (
    .IA(\DLX_IDinst_RegFile_31_5/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_31_5/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_681),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_606)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6811.INIT = 16'hFD5D;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6811 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_585),
    .ADR1(DLX_IDinst_RegFile_28_5),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR3(DLX_IDinst_RegFile_29_5),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_681)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6821.INIT = 16'hFD5D;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6821 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_586),
    .ADR1(DLX_IDinst_RegFile_30_5),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR3(DLX_IDinst_RegFile_31_5),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_682)
  );
  X_BUF \DLX_IDinst_RegFile_31_5/COUTUSED  (
    .I(\DLX_IDinst_RegFile_31_5/CYMUXG ),
    .O(DLX_IDinst__n0620[5])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_607 (
    .IA(\DLX_IDinst_RegFile_31_5/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_606),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_682),
    .O(\DLX_IDinst_RegFile_31_5/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_31_5/CYINIT_938  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_605),
    .O(\DLX_IDinst_RegFile_31_5/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_16_2/LOGIC_ZERO_939  (
    .O(\DLX_IDinst_RegFile_16_2/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_552_940 (
    .IA(\DLX_IDinst_RegFile_16_2/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_16_2/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_627),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_552)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6271.INIT = 16'hDDF5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6271 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_579),
    .ADR1(DLX_IDinst_RegFile_17_2),
    .ADR2(DLX_IDinst_RegFile_16_2),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_627)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6281.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6281 (
    .ADR0(DLX_IDinst_RegFile_19_2),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_580),
    .ADR2(DLX_IDinst_RegFile_18_2),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_628)
  );
  X_BUF \DLX_IDinst_RegFile_16_2/COUTUSED  (
    .I(\DLX_IDinst_RegFile_16_2/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_553)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_553_941 (
    .IA(\DLX_IDinst_RegFile_16_2/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_552),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_628),
    .O(\DLX_IDinst_RegFile_16_2/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_16_2/CYINIT_942  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_551),
    .O(\DLX_IDinst_RegFile_16_2/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_24_2/LOGIC_ZERO_943  (
    .O(\DLX_IDinst_RegFile_24_2/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_44_944 (
    .IA(\DLX_IDinst_RegFile_24_2/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_24_2/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_103),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_44)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1031.INIT = 16'hCFAF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1031 (
    .ADR0(DLX_IDinst_RegFile_24_2),
    .ADR1(DLX_IDinst_RegFile_25_2),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_55),
    .ADR3(DLX_IDinst_jtarget[16]),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_103)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1041.INIT = 16'hCFAF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1041 (
    .ADR0(DLX_IDinst_RegFile_26_2),
    .ADR1(DLX_IDinst_RegFile_27_2),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_56),
    .ADR3(DLX_IDinst_jtarget[16]),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_104)
  );
  X_BUF \DLX_IDinst_RegFile_24_2/COUTUSED  (
    .I(\DLX_IDinst_RegFile_24_2/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_45)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_45_945 (
    .IA(\DLX_IDinst_RegFile_24_2/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_44),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_104),
    .O(\DLX_IDinst_RegFile_24_2/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_24_2/CYINIT_946  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_43),
    .O(\DLX_IDinst_RegFile_24_2/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_31_6/LOGIC_ZERO_947  (
    .O(\DLX_IDinst_RegFile_31_6/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_622_948 (
    .IA(\DLX_IDinst_RegFile_31_6/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_31_6/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_697),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_622)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6971.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6971 (
    .ADR0(DLX_IDinst_RegFile_29_6),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_585),
    .ADR2(DLX_IDinst_RegFile_28_6),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_697)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6981.INIT = 16'hF5DD;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6981 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_586),
    .ADR1(DLX_IDinst_RegFile_30_6),
    .ADR2(DLX_IDinst_RegFile_31_6),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_698)
  );
  X_BUF \DLX_IDinst_RegFile_31_6/COUTUSED  (
    .I(\DLX_IDinst_RegFile_31_6/CYMUXG ),
    .O(DLX_IDinst__n0620[6])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_623 (
    .IA(\DLX_IDinst_RegFile_31_6/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_622),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_698),
    .O(\DLX_IDinst_RegFile_31_6/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_31_6/CYINIT_949  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_621),
    .O(\DLX_IDinst_RegFile_31_6/CYINIT )
  );
  defparam DLX_IDinst_RegFile_19_21_950.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_19_21_950 (
    .I(DLX_IDinst_WB_data_eff[21]),
    .CE(DLX_IDinst__n0588),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_19_21)
  );
  X_ZERO \DLX_IDinst_RegFile_16_3/LOGIC_ZERO_951  (
    .O(\DLX_IDinst_RegFile_16_3/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_56_952 (
    .IA(\DLX_IDinst_RegFile_16_3/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_16_3/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_115),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_56)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1151.INIT = 16'hAFCF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1151 (
    .ADR0(DLX_IDinst_RegFile_17_3),
    .ADR1(DLX_IDinst_RegFile_16_3),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_51),
    .ADR3(DLX_IDinst_jtarget[16]),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_115)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1161.INIT = 16'hE2FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1161 (
    .ADR0(DLX_IDinst_RegFile_18_3),
    .ADR1(DLX_IDinst_jtarget[16]),
    .ADR2(DLX_IDinst_RegFile_19_3),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_52),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_116)
  );
  X_BUF \DLX_IDinst_RegFile_16_3/COUTUSED  (
    .I(\DLX_IDinst_RegFile_16_3/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_57)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_57_953 (
    .IA(\DLX_IDinst_RegFile_16_3/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_56),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_116),
    .O(\DLX_IDinst_RegFile_16_3/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_16_3/CYINIT_954  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_55),
    .O(\DLX_IDinst_RegFile_16_3/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_24_3/LOGIC_ZERO_955  (
    .O(\DLX_IDinst_RegFile_24_3/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_60_956 (
    .IA(\DLX_IDinst_RegFile_24_3/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_24_3/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_119),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_60)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1191.INIT = 16'hCFAF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1191 (
    .ADR0(DLX_IDinst_RegFile_24_3),
    .ADR1(DLX_IDinst_RegFile_25_3),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_55),
    .ADR3(DLX_IDinst_jtarget[16]),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_119)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1201.INIT = 16'hCFAF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1201 (
    .ADR0(DLX_IDinst_RegFile_26_3),
    .ADR1(DLX_IDinst_RegFile_27_3),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_56),
    .ADR3(DLX_IDinst_jtarget[16]),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_120)
  );
  X_BUF \DLX_IDinst_RegFile_24_3/COUTUSED  (
    .I(\DLX_IDinst_RegFile_24_3/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_61)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_61_957 (
    .IA(\DLX_IDinst_RegFile_24_3/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_60),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_120),
    .O(\DLX_IDinst_RegFile_24_3/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_24_3/CYINIT_958  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_59),
    .O(\DLX_IDinst_RegFile_24_3/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_31_7/LOGIC_ZERO_959  (
    .O(\DLX_IDinst_RegFile_31_7/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_638_960 (
    .IA(\DLX_IDinst_RegFile_31_7/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_31_7/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_713),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_638)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7131.INIT = 16'hDDF5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7131 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_585),
    .ADR1(DLX_IDinst_RegFile_29_7),
    .ADR2(DLX_IDinst_RegFile_28_7),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_713)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7141.INIT = 16'hF5DD;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7141 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_586),
    .ADR1(DLX_IDinst_RegFile_30_7),
    .ADR2(DLX_IDinst_RegFile_31_7),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_714)
  );
  X_BUF \DLX_IDinst_RegFile_31_7/COUTUSED  (
    .I(\DLX_IDinst_RegFile_31_7/CYMUXG ),
    .O(DLX_IDinst__n0620[7])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_639 (
    .IA(\DLX_IDinst_RegFile_31_7/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_638),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_714),
    .O(\DLX_IDinst_RegFile_31_7/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_31_7/CYINIT_961  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_637),
    .O(\DLX_IDinst_RegFile_31_7/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_16_4/LOGIC_ZERO_962  (
    .O(\DLX_IDinst_RegFile_16_4/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_72_963 (
    .IA(\DLX_IDinst_RegFile_16_4/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_16_4/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_131),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_72)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1311.INIT = 16'hFB73;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1311 (
    .ADR0(DLX_IDinst_jtarget[16]),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_51),
    .ADR2(DLX_IDinst_RegFile_16_4),
    .ADR3(DLX_IDinst_RegFile_17_4),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_131)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1321.INIT = 16'hE4FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1321 (
    .ADR0(DLX_IDinst_jtarget[16]),
    .ADR1(DLX_IDinst_RegFile_18_4),
    .ADR2(DLX_IDinst_RegFile_19_4),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_52),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_132)
  );
  X_BUF \DLX_IDinst_RegFile_16_4/COUTUSED  (
    .I(\DLX_IDinst_RegFile_16_4/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_73)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_73_964 (
    .IA(\DLX_IDinst_RegFile_16_4/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_72),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_132),
    .O(\DLX_IDinst_RegFile_16_4/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_16_4/CYINIT_965  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_71),
    .O(\DLX_IDinst_RegFile_16_4/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_17_0/LOGIC_ZERO_966  (
    .O(\DLX_IDinst_RegFile_17_0/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_520_967 (
    .IA(\DLX_IDinst_RegFile_17_0/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_17_0/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_595),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_520)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_5951.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_5951 (
    .ADR0(DLX_IDinst_RegFile_16_0),
    .ADR1(DLX_IDinst_RegFile_17_0),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_579),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_595)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_5961.INIT = 16'hDFD5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_5961 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_580),
    .ADR1(DLX_IDinst_RegFile_19_0),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR3(DLX_IDinst_RegFile_18_0),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_596)
  );
  X_BUF \DLX_IDinst_RegFile_17_0/COUTUSED  (
    .I(\DLX_IDinst_RegFile_17_0/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_521)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_521_968 (
    .IA(\DLX_IDinst_RegFile_17_0/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_520),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_596),
    .O(\DLX_IDinst_RegFile_17_0/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_17_0/CYINIT_969  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_519),
    .O(\DLX_IDinst_RegFile_17_0/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_24_4/LOGIC_ZERO_970  (
    .O(\DLX_IDinst_RegFile_24_4/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_76_971 (
    .IA(\DLX_IDinst_RegFile_24_4/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_24_4/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_135),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_76)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1351.INIT = 16'hDF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1351 (
    .ADR0(DLX_IDinst_jtarget[16]),
    .ADR1(DLX_IDinst_RegFile_25_4),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_55),
    .ADR3(DLX_IDinst_RegFile_24_4),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_135)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1361.INIT = 16'hF5DD;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1361 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_56),
    .ADR1(DLX_IDinst_RegFile_26_4),
    .ADR2(DLX_IDinst_RegFile_27_4),
    .ADR3(DLX_IDinst_jtarget[16]),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_136)
  );
  X_BUF \DLX_IDinst_RegFile_24_4/COUTUSED  (
    .I(\DLX_IDinst_RegFile_24_4/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_77)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_77_972 (
    .IA(\DLX_IDinst_RegFile_24_4/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_76),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_136),
    .O(\DLX_IDinst_RegFile_24_4/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_24_4/CYINIT_973  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_75),
    .O(\DLX_IDinst_RegFile_24_4/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_25_0/LOGIC_ZERO_974  (
    .O(\DLX_IDinst_RegFile_25_0/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_524_975 (
    .IA(\DLX_IDinst_RegFile_25_0/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_25_0/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_599),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_524)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_5991.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_5991 (
    .ADR0(DLX_IDinst_RegFile_24_0),
    .ADR1(DLX_IDinst_RegFile_25_0),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_583),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_599)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6001.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6001 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR1(DLX_IDinst_RegFile_26_0),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_584),
    .ADR3(DLX_IDinst_RegFile_27_0),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_600)
  );
  X_BUF \DLX_IDinst_RegFile_25_0/COUTUSED  (
    .I(\DLX_IDinst_RegFile_25_0/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_525)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_525_976 (
    .IA(\DLX_IDinst_RegFile_25_0/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_524),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_600),
    .O(\DLX_IDinst_RegFile_25_0/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_25_0/CYINIT_977  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_523),
    .O(\DLX_IDinst_RegFile_25_0/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_31_8/LOGIC_ZERO_978  (
    .O(\DLX_IDinst_RegFile_31_8/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_654_979 (
    .IA(\DLX_IDinst_RegFile_31_8/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_31_8/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_729),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_654)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7291.INIT = 16'hACFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7291 (
    .ADR0(DLX_IDinst_RegFile_29_8),
    .ADR1(DLX_IDinst_RegFile_28_8),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_585),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_729)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7301.INIT = 16'hB8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7301 (
    .ADR0(DLX_IDinst_RegFile_31_8),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR2(DLX_IDinst_RegFile_30_8),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_586),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_730)
  );
  X_BUF \DLX_IDinst_RegFile_31_8/COUTUSED  (
    .I(\DLX_IDinst_RegFile_31_8/CYMUXG ),
    .O(DLX_IDinst__n0620[8])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_655 (
    .IA(\DLX_IDinst_RegFile_31_8/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_654),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_730),
    .O(\DLX_IDinst_RegFile_31_8/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_31_8/CYINIT_980  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_653),
    .O(\DLX_IDinst_RegFile_31_8/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_16_5/LOGIC_ZERO_981  (
    .O(\DLX_IDinst_RegFile_16_5/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_88_982 (
    .IA(\DLX_IDinst_RegFile_16_5/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_16_5/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_147),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_88)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1471.INIT = 16'hFB3B;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1471 (
    .ADR0(DLX_IDinst_RegFile_16_5),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_51),
    .ADR2(DLX_IDinst_jtarget[16]),
    .ADR3(DLX_IDinst_RegFile_17_5),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_147)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1481.INIT = 16'hF7D5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1481 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_52),
    .ADR1(DLX_IDinst_jtarget[16]),
    .ADR2(DLX_IDinst_RegFile_19_5),
    .ADR3(DLX_IDinst_RegFile_18_5),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_148)
  );
  X_BUF \DLX_IDinst_RegFile_16_5/COUTUSED  (
    .I(\DLX_IDinst_RegFile_16_5/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_89)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_89_983 (
    .IA(\DLX_IDinst_RegFile_16_5/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_88),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_148),
    .O(\DLX_IDinst_RegFile_16_5/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_16_5/CYINIT_984  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_87),
    .O(\DLX_IDinst_RegFile_16_5/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_17_1/LOGIC_ZERO_985  (
    .O(\DLX_IDinst_RegFile_17_1/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_536_986 (
    .IA(\DLX_IDinst_RegFile_17_1/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_17_1/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_611),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_536)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6111.INIT = 16'hE4FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6111 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR1(DLX_IDinst_RegFile_16_1),
    .ADR2(DLX_IDinst_RegFile_17_1),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_579),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_611)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6121.INIT = 16'hFB3B;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6121 (
    .ADR0(DLX_IDinst_RegFile_18_1),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_580),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR3(DLX_IDinst_RegFile_19_1),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_612)
  );
  X_BUF \DLX_IDinst_RegFile_17_1/COUTUSED  (
    .I(\DLX_IDinst_RegFile_17_1/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_537)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_537_987 (
    .IA(\DLX_IDinst_RegFile_17_1/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_536),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_612),
    .O(\DLX_IDinst_RegFile_17_1/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_17_1/CYINIT_988  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_535),
    .O(\DLX_IDinst_RegFile_17_1/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_24_5/LOGIC_ZERO_989  (
    .O(\DLX_IDinst_RegFile_24_5/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_92_990 (
    .IA(\DLX_IDinst_RegFile_24_5/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_24_5/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_151),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_92)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1511.INIT = 16'hAFCF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1511 (
    .ADR0(DLX_IDinst_RegFile_25_5),
    .ADR1(DLX_IDinst_RegFile_24_5),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_55),
    .ADR3(DLX_IDinst_jtarget[16]),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_151)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1521.INIT = 16'hBFB3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1521 (
    .ADR0(DLX_IDinst_RegFile_27_5),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_56),
    .ADR2(DLX_IDinst_jtarget[16]),
    .ADR3(DLX_IDinst_RegFile_26_5),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_152)
  );
  X_BUF \DLX_IDinst_RegFile_24_5/COUTUSED  (
    .I(\DLX_IDinst_RegFile_24_5/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_93)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_93_991 (
    .IA(\DLX_IDinst_RegFile_24_5/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_92),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_152),
    .O(\DLX_IDinst_RegFile_24_5/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_24_5/CYINIT_992  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_91),
    .O(\DLX_IDinst_RegFile_24_5/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_25_1/LOGIC_ZERO_993  (
    .O(\DLX_IDinst_RegFile_25_1/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_540_994 (
    .IA(\DLX_IDinst_RegFile_25_1/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_25_1/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_615),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_540)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6151.INIT = 16'hCFAF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6151 (
    .ADR0(DLX_IDinst_RegFile_24_1),
    .ADR1(DLX_IDinst_RegFile_25_1),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_583),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_615)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6161.INIT = 16'hBFB3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6161 (
    .ADR0(DLX_IDinst_RegFile_27_1),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_584),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR3(DLX_IDinst_RegFile_26_1),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_616)
  );
  X_BUF \DLX_IDinst_RegFile_25_1/COUTUSED  (
    .I(\DLX_IDinst_RegFile_25_1/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_541)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_541_995 (
    .IA(\DLX_IDinst_RegFile_25_1/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_540),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_616),
    .O(\DLX_IDinst_RegFile_25_1/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_25_1/CYINIT_996  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_539),
    .O(\DLX_IDinst_RegFile_25_1/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_31_9/LOGIC_ZERO_997  (
    .O(\DLX_IDinst_RegFile_31_9/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_670_998 (
    .IA(\DLX_IDinst_RegFile_31_9/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_31_9/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_745),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_670)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7451.INIT = 16'hBF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7451 (
    .ADR0(DLX_IDinst_RegFile_29_9),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_585),
    .ADR3(DLX_IDinst_RegFile_28_9),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_745)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7461.INIT = 16'hBF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7461 (
    .ADR0(DLX_IDinst_RegFile_31_9),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_586),
    .ADR3(DLX_IDinst_RegFile_30_9),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_746)
  );
  X_BUF \DLX_IDinst_RegFile_31_9/COUTUSED  (
    .I(\DLX_IDinst_RegFile_31_9/CYMUXG ),
    .O(DLX_IDinst__n0620[9])
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_671 (
    .IA(\DLX_IDinst_RegFile_31_9/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_670),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_746),
    .O(\DLX_IDinst_RegFile_31_9/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_31_9/CYINIT_999  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_669),
    .O(\DLX_IDinst_RegFile_31_9/CYINIT )
  );
  defparam vga_top_vga1__n00084.INIT = 16'h8000;
  X_LUT4 vga_top_vga1__n00084 (
    .ADR0(vga_top_vga1_hcounter[4]),
    .ADR1(vga_top_vga1_hcounter[5]),
    .ADR2(vga_top_vga1_hcounter[7]),
    .ADR3(vga_top_vga1_hcounter[1]),
    .O(\CHOICE3139/GROM )
  );
  X_BUF \CHOICE3139/YUSED  (
    .I(\CHOICE3139/GROM ),
    .O(CHOICE3139)
  );
  X_ZERO \DLX_IDinst_RegFile_16_6/LOGIC_ZERO_1000  (
    .O(\DLX_IDinst_RegFile_16_6/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_104_1001 (
    .IA(\DLX_IDinst_RegFile_16_6/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_16_6/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_163),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_104)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1631.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1631 (
    .ADR0(DLX_IDinst_RegFile_17_6),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_51),
    .ADR2(DLX_IDinst_RegFile_16_6),
    .ADR3(DLX_IDinst_jtarget[16]),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_163)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1641.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1641 (
    .ADR0(DLX_IDinst_RegFile_18_6),
    .ADR1(DLX_IDinst_RegFile_19_6),
    .ADR2(DLX_IDinst_jtarget[16]),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_52),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_164)
  );
  X_BUF \DLX_IDinst_RegFile_16_6/COUTUSED  (
    .I(\DLX_IDinst_RegFile_16_6/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_105)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_105_1002 (
    .IA(\DLX_IDinst_RegFile_16_6/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_104),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_164),
    .O(\DLX_IDinst_RegFile_16_6/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_16_6/CYINIT_1003  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_103),
    .O(\DLX_IDinst_RegFile_16_6/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_24_6/LOGIC_ZERO_1004  (
    .O(\DLX_IDinst_RegFile_24_6/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_108_1005 (
    .IA(\DLX_IDinst_RegFile_24_6/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_24_6/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_167),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_108)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1671.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1671 (
    .ADR0(DLX_IDinst_RegFile_24_6),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_55),
    .ADR2(DLX_IDinst_RegFile_25_6),
    .ADR3(DLX_IDinst_jtarget[16]),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_167)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1681.INIT = 16'hDF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1681 (
    .ADR0(DLX_IDinst_jtarget[16]),
    .ADR1(DLX_IDinst_RegFile_27_6),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_56),
    .ADR3(DLX_IDinst_RegFile_26_6),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_168)
  );
  X_BUF \DLX_IDinst_RegFile_24_6/COUTUSED  (
    .I(\DLX_IDinst_RegFile_24_6/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_109)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_109_1006 (
    .IA(\DLX_IDinst_RegFile_24_6/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_108),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_168),
    .O(\DLX_IDinst_RegFile_24_6/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_24_6/CYINIT_1007  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_107),
    .O(\DLX_IDinst_RegFile_24_6/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_16_7/LOGIC_ZERO_1008  (
    .O(\DLX_IDinst_RegFile_16_7/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_632_1009 (
    .IA(\DLX_IDinst_RegFile_16_7/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_16_7/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_707),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_632)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7071.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7071 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_579),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR2(DLX_IDinst_RegFile_16_7),
    .ADR3(DLX_IDinst_RegFile_17_7),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_707)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7081.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7081 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_580),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR2(DLX_IDinst_RegFile_18_7),
    .ADR3(DLX_IDinst_RegFile_19_7),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_708)
  );
  X_BUF \DLX_IDinst_RegFile_16_7/COUTUSED  (
    .I(\DLX_IDinst_RegFile_16_7/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_633)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_633_1010 (
    .IA(\DLX_IDinst_RegFile_16_7/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_632),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_708),
    .O(\DLX_IDinst_RegFile_16_7/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_16_7/CYINIT_1011  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_631),
    .O(\DLX_IDinst_RegFile_16_7/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_17_3/LOGIC_ZERO_1012  (
    .O(\DLX_IDinst_RegFile_17_3/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_568_1013 (
    .IA(\DLX_IDinst_RegFile_17_3/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_17_3/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_643),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_568)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6431.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6431 (
    .ADR0(DLX_IDinst_RegFile_16_3),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_579),
    .ADR2(DLX_IDinst_RegFile_17_3),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_643)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6441.INIT = 16'hBF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6441 (
    .ADR0(DLX_IDinst_RegFile_19_3),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_580),
    .ADR3(DLX_IDinst_RegFile_18_3),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_644)
  );
  X_BUF \DLX_IDinst_RegFile_17_3/COUTUSED  (
    .I(\DLX_IDinst_RegFile_17_3/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_569)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_569_1014 (
    .IA(\DLX_IDinst_RegFile_17_3/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_568),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_644),
    .O(\DLX_IDinst_RegFile_17_3/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_17_3/CYINIT_1015  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_567),
    .O(\DLX_IDinst_RegFile_17_3/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_24_7/LOGIC_ZERO_1016  (
    .O(\DLX_IDinst_RegFile_24_7/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_124_1017 (
    .IA(\DLX_IDinst_RegFile_24_7/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_24_7/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_183),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_124)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1831.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1831 (
    .ADR0(DLX_IDinst_RegFile_24_7),
    .ADR1(DLX_IDinst_RegFile_25_7),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_55),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_183)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1841.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1841 (
    .ADR0(DLX_IDinst_RegFile_26_7),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_56),
    .ADR3(DLX_IDinst_RegFile_27_7),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_184)
  );
  X_BUF \DLX_IDinst_RegFile_24_7/COUTUSED  (
    .I(\DLX_IDinst_RegFile_24_7/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_125)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_125_1018 (
    .IA(\DLX_IDinst_RegFile_24_7/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_124),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_184),
    .O(\DLX_IDinst_RegFile_24_7/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_24_7/CYINIT_1019  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_123),
    .O(\DLX_IDinst_RegFile_24_7/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_25_3/LOGIC_ZERO_1020  (
    .O(\DLX_IDinst_RegFile_25_3/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_572_1021 (
    .IA(\DLX_IDinst_RegFile_25_3/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_25_3/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_647),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_572)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6471.INIT = 16'hE2FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6471 (
    .ADR0(DLX_IDinst_RegFile_24_3),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR2(DLX_IDinst_RegFile_25_3),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_583),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_647)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6481.INIT = 16'hF7D5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6481 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_584),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR2(DLX_IDinst_RegFile_27_3),
    .ADR3(DLX_IDinst_RegFile_26_3),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_648)
  );
  X_BUF \DLX_IDinst_RegFile_25_3/COUTUSED  (
    .I(\DLX_IDinst_RegFile_25_3/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_573)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_573_1022 (
    .IA(\DLX_IDinst_RegFile_25_3/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_572),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_648),
    .O(\DLX_IDinst_RegFile_25_3/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_25_3/CYINIT_1023  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_571),
    .O(\DLX_IDinst_RegFile_25_3/CYINIT )
  );
  defparam vga_top_vga1__n00094.INIT = 16'hFFFE;
  X_LUT4 vga_top_vga1__n00094 (
    .ADR0(vga_top_vga1_vcounter[4]),
    .ADR1(vga_top_vga1_vcounter[2]),
    .ADR2(vga_top_vga1_vcounter[5]),
    .ADR3(vga_top_vga1_vcounter[3]),
    .O(\CHOICE3455/GROM )
  );
  X_BUF \CHOICE3455/YUSED  (
    .I(\CHOICE3455/GROM ),
    .O(CHOICE3455)
  );
  X_ZERO \DLX_IDinst_RegFile_16_8/LOGIC_ZERO_1024  (
    .O(\DLX_IDinst_RegFile_16_8/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_136_1025 (
    .IA(\DLX_IDinst_RegFile_16_8/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_16_8/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_195),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_136)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1951.INIT = 16'hFB73;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1951 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_51),
    .ADR2(DLX_IDinst_RegFile_16_8),
    .ADR3(DLX_IDinst_RegFile_17_8),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_195)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1961.INIT = 16'hDFD5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1961 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_52),
    .ADR1(DLX_IDinst_RegFile_19_8),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR3(DLX_IDinst_RegFile_18_8),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_196)
  );
  X_BUF \DLX_IDinst_RegFile_16_8/COUTUSED  (
    .I(\DLX_IDinst_RegFile_16_8/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_137)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_137_1026 (
    .IA(\DLX_IDinst_RegFile_16_8/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_136),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_196),
    .O(\DLX_IDinst_RegFile_16_8/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_16_8/CYINIT_1027  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_135),
    .O(\DLX_IDinst_RegFile_16_8/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_17_4/LOGIC_ZERO_1028  (
    .O(\DLX_IDinst_RegFile_17_4/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_584_1029 (
    .IA(\DLX_IDinst_RegFile_17_4/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_17_4/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_659),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_584)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6591.INIT = 16'hDFD5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6591 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_579),
    .ADR1(DLX_IDinst_RegFile_17_4),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR3(DLX_IDinst_RegFile_16_4),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_659)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6601.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6601 (
    .ADR0(DLX_IDinst_RegFile_19_4),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_580),
    .ADR2(DLX_IDinst_RegFile_18_4),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_660)
  );
  X_BUF \DLX_IDinst_RegFile_17_4/COUTUSED  (
    .I(\DLX_IDinst_RegFile_17_4/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_585)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_585_1030 (
    .IA(\DLX_IDinst_RegFile_17_4/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_584),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_660),
    .O(\DLX_IDinst_RegFile_17_4/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_17_4/CYINIT_1031  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_583),
    .O(\DLX_IDinst_RegFile_17_4/CYINIT )
  );
  defparam DLX_IDinst_RegFile_19_13_1032.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_19_13_1032 (
    .I(DLX_IDinst_WB_data_eff[13]),
    .CE(DLX_IDinst__n0588),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_19_13)
  );
  X_ZERO \DLX_IDinst_RegFile_24_8/LOGIC_ZERO_1033  (
    .O(\DLX_IDinst_RegFile_24_8/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_140_1034 (
    .IA(\DLX_IDinst_RegFile_24_8/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_24_8/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_199),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_140)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1991.INIT = 16'hE2FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1991 (
    .ADR0(DLX_IDinst_RegFile_24_8),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR2(DLX_IDinst_RegFile_25_8),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_55),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_199)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2001.INIT = 16'hFB3B;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2001 (
    .ADR0(DLX_IDinst_RegFile_26_8),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_56),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR3(DLX_IDinst_RegFile_27_8),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_200)
  );
  X_BUF \DLX_IDinst_RegFile_24_8/COUTUSED  (
    .I(\DLX_IDinst_RegFile_24_8/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_141)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_141_1035 (
    .IA(\DLX_IDinst_RegFile_24_8/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_140),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_200),
    .O(\DLX_IDinst_RegFile_24_8/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_24_8/CYINIT_1036  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_139),
    .O(\DLX_IDinst_RegFile_24_8/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_25_4/LOGIC_ZERO_1037  (
    .O(\DLX_IDinst_RegFile_25_4/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_588_1038 (
    .IA(\DLX_IDinst_RegFile_25_4/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_25_4/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_663),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_588)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6631.INIT = 16'hDF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6631 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR1(DLX_IDinst_RegFile_25_4),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_583),
    .ADR3(DLX_IDinst_RegFile_24_4),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_663)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6641.INIT = 16'hDF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6641 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR1(DLX_IDinst_RegFile_27_4),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_584),
    .ADR3(DLX_IDinst_RegFile_26_4),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_664)
  );
  X_BUF \DLX_IDinst_RegFile_25_4/COUTUSED  (
    .I(\DLX_IDinst_RegFile_25_4/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_589)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_589_1039 (
    .IA(\DLX_IDinst_RegFile_25_4/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_588),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_664),
    .O(\DLX_IDinst_RegFile_25_4/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_25_4/CYINIT_1040  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_587),
    .O(\DLX_IDinst_RegFile_25_4/CYINIT )
  );
  defparam \DLX_IDinst__n0146<0>48 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst__n0146<0>48  (
    .ADR0(CHOICE3249),
    .ADR1(DLX_IDinst_N107105),
    .ADR2(N163574),
    .ADR3(N134590),
    .O(\CHOICE3251/FROM )
  );
  defparam \DLX_IDinst__n0146<31>48 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst__n0146<31>48  (
    .ADR0(CHOICE3230),
    .ADR1(DLX_IDinst_N107105),
    .ADR2(N134590),
    .ADR3(N163652),
    .O(\CHOICE3251/GROM )
  );
  X_BUF \CHOICE3251/XUSED  (
    .I(\CHOICE3251/FROM ),
    .O(CHOICE3251)
  );
  X_BUF \CHOICE3251/YUSED  (
    .I(\CHOICE3251/GROM ),
    .O(CHOICE3232)
  );
  X_ZERO \DLX_IDinst_RegFile_16_9/LOGIC_ZERO_1041  (
    .O(\DLX_IDinst_RegFile_16_9/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_152_1042 (
    .IA(\DLX_IDinst_RegFile_16_9/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_16_9/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_211),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_152)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2111.INIT = 16'hFB3B;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2111 (
    .ADR0(DLX_IDinst_RegFile_16_9),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_51),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR3(DLX_IDinst_RegFile_17_9),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_211)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2121.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2121 (
    .ADR0(DLX_IDinst_RegFile_18_9),
    .ADR1(DLX_IDinst_RegFile_19_9),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_52),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_212)
  );
  X_BUF \DLX_IDinst_RegFile_16_9/COUTUSED  (
    .I(\DLX_IDinst_RegFile_16_9/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_153)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_153_1043 (
    .IA(\DLX_IDinst_RegFile_16_9/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_152),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_212),
    .O(\DLX_IDinst_RegFile_16_9/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_16_9/CYINIT_1044  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_151),
    .O(\DLX_IDinst_RegFile_16_9/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_17_5/LOGIC_ZERO_1045  (
    .O(\DLX_IDinst_RegFile_17_5/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_600_1046 (
    .IA(\DLX_IDinst_RegFile_17_5/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_17_5/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_675),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_600)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6751.INIT = 16'hD8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6751 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR1(DLX_IDinst_RegFile_17_5),
    .ADR2(DLX_IDinst_RegFile_16_5),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_579),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_675)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6761.INIT = 16'hDF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6761 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR1(DLX_IDinst_RegFile_19_5),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_580),
    .ADR3(DLX_IDinst_RegFile_18_5),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_676)
  );
  X_BUF \DLX_IDinst_RegFile_17_5/COUTUSED  (
    .I(\DLX_IDinst_RegFile_17_5/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_601)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_601_1047 (
    .IA(\DLX_IDinst_RegFile_17_5/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_600),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_676),
    .O(\DLX_IDinst_RegFile_17_5/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_17_5/CYINIT_1048  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_599),
    .O(\DLX_IDinst_RegFile_17_5/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_24_9/LOGIC_ZERO_1049  (
    .O(\DLX_IDinst_RegFile_24_9/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_156_1050 (
    .IA(\DLX_IDinst_RegFile_24_9/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_24_9/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_215),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_156)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2151.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2151 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR1(DLX_IDinst_RegFile_24_9),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_55),
    .ADR3(DLX_IDinst_RegFile_25_9),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_215)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2161.INIT = 16'hCFAF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2161 (
    .ADR0(DLX_IDinst_RegFile_26_9),
    .ADR1(DLX_IDinst_RegFile_27_9),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_56),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_216)
  );
  X_BUF \DLX_IDinst_RegFile_24_9/COUTUSED  (
    .I(\DLX_IDinst_RegFile_24_9/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_157)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_157_1051 (
    .IA(\DLX_IDinst_RegFile_24_9/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_156),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_216),
    .O(\DLX_IDinst_RegFile_24_9/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_24_9/CYINIT_1052  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_155),
    .O(\DLX_IDinst_RegFile_24_9/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_25_5/LOGIC_ZERO_1053  (
    .O(\DLX_IDinst_RegFile_25_5/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_604_1054 (
    .IA(\DLX_IDinst_RegFile_25_5/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_25_5/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_679),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_604)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6791.INIT = 16'hFD5D;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6791 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_583),
    .ADR1(DLX_IDinst_RegFile_24_5),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR3(DLX_IDinst_RegFile_25_5),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_679)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6801.INIT = 16'hF7B3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6801 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_584),
    .ADR2(DLX_IDinst_RegFile_27_5),
    .ADR3(DLX_IDinst_RegFile_26_5),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_680)
  );
  X_BUF \DLX_IDinst_RegFile_25_5/COUTUSED  (
    .I(\DLX_IDinst_RegFile_25_5/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_605)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_605_1055 (
    .IA(\DLX_IDinst_RegFile_25_5/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_604),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_680),
    .O(\DLX_IDinst_RegFile_25_5/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_25_5/CYINIT_1056  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_603),
    .O(\DLX_IDinst_RegFile_25_5/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_17_6/LOGIC_ZERO_1057  (
    .O(\DLX_IDinst_RegFile_17_6/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_616_1058 (
    .IA(\DLX_IDinst_RegFile_17_6/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_17_6/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_691),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_616)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6911.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6911 (
    .ADR0(DLX_IDinst_RegFile_16_6),
    .ADR1(DLX_IDinst_RegFile_17_6),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_579),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_691)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6921.INIT = 16'hACFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6921 (
    .ADR0(DLX_IDinst_RegFile_19_6),
    .ADR1(DLX_IDinst_RegFile_18_6),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_580),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_692)
  );
  X_BUF \DLX_IDinst_RegFile_17_6/COUTUSED  (
    .I(\DLX_IDinst_RegFile_17_6/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_617)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_617_1059 (
    .IA(\DLX_IDinst_RegFile_17_6/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_616),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_692),
    .O(\DLX_IDinst_RegFile_17_6/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_17_6/CYINIT_1060  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_615),
    .O(\DLX_IDinst_RegFile_17_6/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_25_6/LOGIC_ZERO_1061  (
    .O(\DLX_IDinst_RegFile_25_6/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_620_1062 (
    .IA(\DLX_IDinst_RegFile_25_6/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_25_6/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_695),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_620)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6951.INIT = 16'hCFAF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6951 (
    .ADR0(DLX_IDinst_RegFile_24_6),
    .ADR1(DLX_IDinst_RegFile_25_6),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_583),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_695)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6961.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6961 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR1(DLX_IDinst_RegFile_26_6),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_584),
    .ADR3(DLX_IDinst_RegFile_27_6),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_696)
  );
  X_BUF \DLX_IDinst_RegFile_25_6/COUTUSED  (
    .I(\DLX_IDinst_RegFile_25_6/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_621)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_621_1063 (
    .IA(\DLX_IDinst_RegFile_25_6/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_620),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_696),
    .O(\DLX_IDinst_RegFile_25_6/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_25_6/CYINIT_1064  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_619),
    .O(\DLX_IDinst_RegFile_25_6/CYINIT )
  );
  defparam \vga_top_vga1_helpcounter_Madd__n0000_Mxor_Result<2>_Result1 .INIT = 16'h66CC;
  X_LUT4 \vga_top_vga1_helpcounter_Madd__n0000_Mxor_Result<2>_Result1  (
    .ADR0(vga_top_vga1_helpcounter[0]),
    .ADR1(vga_top_vga1_helpcounter[2]),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_helpcounter[1]),
    .O(vga_top_vga1_helpcounter__n0000[2])
  );
  defparam vga_top_vga1__n00521.INIT = 16'hC0FF;
  X_LUT4 vga_top_vga1__n00521 (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_helpcounter[2]),
    .ADR2(vga_top_vga1_helpcounter[1]),
    .ADR3(vga_top_vga1_clockcounter_FFd1),
    .O(\vga_top_vga1_helpcounter<2>/GROM )
  );
  X_BUF \vga_top_vga1_helpcounter<2>/YUSED  (
    .I(\vga_top_vga1_helpcounter<2>/GROM ),
    .O(vga_top_vga1__n0052)
  );
  X_ZERO \DLX_IDinst_RegFile_25_7/LOGIC_ZERO_1065  (
    .O(\DLX_IDinst_RegFile_25_7/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_636_1066 (
    .IA(\DLX_IDinst_RegFile_25_7/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_25_7/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_711),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_636)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7111.INIT = 16'hF7B3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7111 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_583),
    .ADR2(DLX_IDinst_RegFile_25_7),
    .ADR3(DLX_IDinst_RegFile_24_7),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_711)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7121.INIT = 16'hD8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7121 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR1(DLX_IDinst_RegFile_27_7),
    .ADR2(DLX_IDinst_RegFile_26_7),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_584),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_712)
  );
  X_BUF \DLX_IDinst_RegFile_25_7/COUTUSED  (
    .I(\DLX_IDinst_RegFile_25_7/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_637)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_637_1067 (
    .IA(\DLX_IDinst_RegFile_25_7/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_636),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_712),
    .O(\DLX_IDinst_RegFile_25_7/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_25_7/CYINIT_1068  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_635),
    .O(\DLX_IDinst_RegFile_25_7/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_25_8/LOGIC_ZERO_1069  (
    .O(\DLX_IDinst_RegFile_25_8/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_652_1070 (
    .IA(\DLX_IDinst_RegFile_25_8/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_25_8/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_727),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_652)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7271.INIT = 16'hF7D5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7271 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_583),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR2(DLX_IDinst_RegFile_25_8),
    .ADR3(DLX_IDinst_RegFile_24_8),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_727)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7281.INIT = 16'hF5DD;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7281 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_584),
    .ADR1(DLX_IDinst_RegFile_26_8),
    .ADR2(DLX_IDinst_RegFile_27_8),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_728)
  );
  X_BUF \DLX_IDinst_RegFile_25_8/COUTUSED  (
    .I(\DLX_IDinst_RegFile_25_8/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_653)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_653_1071 (
    .IA(\DLX_IDinst_RegFile_25_8/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_652),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_728),
    .O(\DLX_IDinst_RegFile_25_8/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_25_8/CYINIT_1072  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_651),
    .O(\DLX_IDinst_RegFile_25_8/CYINIT )
  );
  defparam vga_top_vga1__n00098.INIT = 16'hFFEE;
  X_LUT4 vga_top_vga1__n00098 (
    .ADR0(vga_top_vga1_vcounter[0]),
    .ADR1(vga_top_vga1_vcounter[1]),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_vcounter[8]),
    .O(\DLX_IFinst_IR_previous<22>/FROM )
  );
  defparam vga_top_vga1__n000910.INIT = 16'hFFFC;
  X_LUT4 vga_top_vga1__n000910 (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_vcounter[7]),
    .ADR2(vga_top_vga1_vcounter[6]),
    .ADR3(CHOICE3458),
    .O(\DLX_IFinst_IR_previous<22>/GROM )
  );
  X_BUF \DLX_IFinst_IR_previous<22>/XUSED  (
    .I(\DLX_IFinst_IR_previous<22>/FROM ),
    .O(CHOICE3458)
  );
  X_BUF \DLX_IFinst_IR_previous<22>/YUSED  (
    .I(\DLX_IFinst_IR_previous<22>/GROM ),
    .O(CHOICE3459)
  );
  defparam DLX_IDinst_RegFile_17_9_1073.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_17_9_1073 (
    .I(DLX_IDinst_WB_data_eff[9]),
    .CE(DLX_IDinst__n0584),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_17_9)
  );
  X_ZERO \DLX_IDinst_RegFile_17_9/LOGIC_ZERO_1074  (
    .O(\DLX_IDinst_RegFile_17_9/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_664_1075 (
    .IA(\DLX_IDinst_RegFile_17_9/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_17_9/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_739),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_664)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7391.INIT = 16'hDFD5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7391 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_579),
    .ADR1(DLX_IDinst_RegFile_17_9),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR3(DLX_IDinst_RegFile_16_9),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_739)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7401.INIT = 16'hDFD5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7401 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_580),
    .ADR1(DLX_IDinst_RegFile_19_9),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR3(DLX_IDinst_RegFile_18_9),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_740)
  );
  X_BUF \DLX_IDinst_RegFile_17_9/COUTUSED  (
    .I(\DLX_IDinst_RegFile_17_9/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_665)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_665_1076 (
    .IA(\DLX_IDinst_RegFile_17_9/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_664),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_740),
    .O(\DLX_IDinst_RegFile_17_9/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_17_9/CYINIT_1077  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_663),
    .O(\DLX_IDinst_RegFile_17_9/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_25_9/LOGIC_ZERO_1078  (
    .O(\DLX_IDinst_RegFile_25_9/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_668_1079 (
    .IA(\DLX_IDinst_RegFile_25_9/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_25_9/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_743),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_668)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7431.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7431 (
    .ADR0(DLX_IDinst_RegFile_24_9),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_583),
    .ADR2(DLX_IDinst_RegFile_25_9),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_743)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7441.INIT = 16'hDDF5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7441 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_584),
    .ADR1(DLX_IDinst_RegFile_27_9),
    .ADR2(DLX_IDinst_RegFile_26_9),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_744)
  );
  X_BUF \DLX_IDinst_RegFile_25_9/COUTUSED  (
    .I(\DLX_IDinst_RegFile_25_9/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_669)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_669_1080 (
    .IA(\DLX_IDinst_RegFile_25_9/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_668),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_744),
    .O(\DLX_IDinst_RegFile_25_9/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_25_9/CYINIT_1081  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_667),
    .O(\DLX_IDinst_RegFile_25_9/CYINIT )
  );
  defparam DLX_IDinst_RegFile_27_21_1082.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_27_21_1082 (
    .I(DLX_IDinst_WB_data_eff[21]),
    .CE(DLX_IDinst__n0604),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_27_21)
  );
  defparam DLX_IDinst_RegFile_26_29_1083.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_26_29_1083 (
    .I(DLX_IDinst_WB_data_eff[29]),
    .CE(DLX_IDinst__n0602),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_26_29)
  );
  defparam DLX_IDinst_RegFile_27_13_1084.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_27_13_1084 (
    .I(DLX_IDinst_WB_data_eff[13]),
    .CE(DLX_IDinst__n0604),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_27_13)
  );
  defparam DLX_IDinst_RegFile_19_22_1085.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_19_22_1085 (
    .I(DLX_IDinst_WB_data_eff[22]),
    .CE(DLX_IDinst__n0588),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_19_22)
  );
  defparam DLX_IFinst_IR_curr_N30871.INIT = 16'h0011;
  X_LUT4 DLX_IFinst_IR_curr_N30871 (
    .ADR0(DLX_IDinst_counter[1]),
    .ADR1(DLX_IDinst_counter[0]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_stall),
    .O(\DLX_IFinst_IR_curr_N3087/FROM )
  );
  defparam DLX_EXinst__n00061.INIT = 16'hFEFE;
  X_LUT4 DLX_EXinst__n00061 (
    .ADR0(DLX_IDinst_counter[1]),
    .ADR1(DLX_IDinst_counter[0]),
    .ADR2(reset_IBUF),
    .ADR3(VCC),
    .O(\DLX_IFinst_IR_curr_N3087/GROM )
  );
  X_BUF \DLX_IFinst_IR_curr_N3087/XUSED  (
    .I(\DLX_IFinst_IR_curr_N3087/FROM ),
    .O(DLX_IFinst_IR_curr_N3087)
  );
  X_BUF \DLX_IFinst_IR_curr_N3087/YUSED  (
    .I(\DLX_IFinst_IR_curr_N3087/GROM ),
    .O(DLX_EXinst__n0006)
  );
  defparam DLX_EXinst_Ker7495960.INIT = 16'h4400;
  X_LUT4 DLX_EXinst_Ker7495960 (
    .ADR0(DLX_IDinst_reg_out_B[5]),
    .ADR1(DLX_IDinst_reg_out_B_3_1),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[31]),
    .O(\DLX_IDinst_RegFile_6_9/FROM )
  );
  defparam DLX_EXinst__n00324.INIT = 16'hFFFE;
  X_LUT4 DLX_EXinst__n00324 (
    .ADR0(DLX_IDinst_reg_out_B[31]),
    .ADR1(DLX_IDinst_reg_out_B[5]),
    .ADR2(DLX_IDinst_reg_out_B[6]),
    .ADR3(DLX_IDinst_reg_out_B[7]),
    .O(\DLX_IDinst_RegFile_6_9/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_6_9/XUSED  (
    .I(\DLX_IDinst_RegFile_6_9/FROM ),
    .O(CHOICE1944)
  );
  X_BUF \DLX_IDinst_RegFile_6_9/YUSED  (
    .I(\DLX_IDinst_RegFile_6_9/GROM ),
    .O(CHOICE3570)
  );
  defparam \DLX_EXinst__n0007<4>106_SW0 .INIT = 16'hCCEC;
  X_LUT4 \DLX_EXinst__n0007<4>106_SW0  (
    .ADR0(DLX_EXinst_N76338),
    .ADR1(CHOICE4342),
    .ADR2(DLX_EXinst_N72898),
    .ADR3(DLX_IDinst_reg_out_B[3]),
    .O(\N163432/FROM )
  );
  defparam \DLX_EXinst__n0007<4>106 .INIT = 16'hD5C0;
  X_LUT4 \DLX_EXinst__n0007<4>106  (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(DLX_IDinst_reg_out_A[4]),
    .ADR2(DLX_EXinst_N74245),
    .ADR3(N163432),
    .O(\N163432/GROM )
  );
  X_BUF \N163432/XUSED  (
    .I(\N163432/FROM ),
    .O(N163432)
  );
  X_BUF \N163432/YUSED  (
    .I(\N163432/GROM ),
    .O(CHOICE4347)
  );
  defparam \DLX_EXinst__n0007<0>669 .INIT = 16'h0400;
  X_LUT4 \DLX_EXinst__n0007<0>669  (
    .ADR0(\DLX_IDinst_Imm[3] ),
    .ADR1(DLX_EXinst_N76318),
    .ADR2(\DLX_IDinst_Imm[2] ),
    .ADR3(\DLX_EXinst_Mshift__n0021_Sh[0] ),
    .O(\CHOICE6002/FROM )
  );
  defparam DLX_EXinst__n01405.INIT = 16'hAA80;
  X_LUT4 DLX_EXinst__n01405 (
    .ADR0(\DLX_IDinst_Imm[2] ),
    .ADR1(DLX_IDinst_IR_function_field[5]),
    .ADR2(\DLX_IDinst_Imm[0] ),
    .ADR3(\DLX_IDinst_Imm[3] ),
    .O(\CHOICE6002/GROM )
  );
  X_BUF \CHOICE6002/XUSED  (
    .I(\CHOICE6002/FROM ),
    .O(CHOICE6002)
  );
  X_BUF \CHOICE6002/YUSED  (
    .I(\CHOICE6002/GROM ),
    .O(CHOICE1299)
  );
  defparam DLX_EXinst__n00561.INIT = 16'h00C0;
  X_LUT4 DLX_EXinst__n00561 (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N76041),
    .ADR2(DLX_IDinst_IR_opcode_field[1]),
    .ADR3(DLX_IDinst_IR_opcode_field[0]),
    .O(\DLX_EXinst__n0056/FROM )
  );
  defparam \DLX_EXinst__n0007<27>75_SW0 .INIT = 16'hFAF0;
  X_LUT4 \DLX_EXinst__n0007<27>75_SW0  (
    .ADR0(\DLX_EXinst_Mshift__n0022_Sh[59] ),
    .ADR1(VCC),
    .ADR2(CHOICE4942),
    .ADR3(DLX_EXinst__n0056),
    .O(\DLX_EXinst__n0056/GROM )
  );
  X_BUF \DLX_EXinst__n0056/XUSED  (
    .I(\DLX_EXinst__n0056/FROM ),
    .O(DLX_EXinst__n0056)
  );
  X_BUF \DLX_EXinst__n0056/YUSED  (
    .I(\DLX_EXinst__n0056/GROM ),
    .O(N163530)
  );
  defparam DLX_EXinst__n01441.INIT = 16'h0033;
  X_LUT4 DLX_EXinst__n01441 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_counter[1]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_counter[0]),
    .O(\DLX_IDinst_RegFile_2_14/FROM )
  );
  defparam DLX_IDinst__n0164_SW0.INIT = 16'hCFAF;
  X_LUT4 DLX_IDinst__n0164_SW0 (
    .ADR0(DLX_IDinst_current_IR[28]),
    .ADR1(DLX_IFinst_IR_latched[28]),
    .ADR2(DLX_IDinst_IR_latched[26]),
    .ADR3(DLX_EXinst__n0144),
    .O(\DLX_IDinst_RegFile_2_14/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_2_14/XUSED  (
    .I(\DLX_IDinst_RegFile_2_14/FROM ),
    .O(DLX_EXinst__n0144)
  );
  X_BUF \DLX_IDinst_RegFile_2_14/YUSED  (
    .I(\DLX_IDinst_RegFile_2_14/GROM ),
    .O(N127043)
  );
  defparam DLX_EXinst__n00801.INIT = 16'h0100;
  X_LUT4 DLX_EXinst__n00801 (
    .ADR0(\DLX_IDinst_Imm[1] ),
    .ADR1(\DLX_IDinst_Imm[0] ),
    .ADR2(DLX_IDinst_IR_function_field[5]),
    .ADR3(DLX_EXinst_N76002),
    .O(\DLX_EXinst__n0080/FROM )
  );
  defparam \DLX_EXinst__n0007<23>272_SW0 .INIT = 16'hDCCC;
  X_LUT4 \DLX_EXinst__n0007<23>272_SW0  (
    .ADR0(N148323),
    .ADR1(CHOICE4051),
    .ADR2(CHOICE4037),
    .ADR3(DLX_EXinst__n0080),
    .O(\DLX_EXinst__n0080/GROM )
  );
  X_BUF \DLX_EXinst__n0080/XUSED  (
    .I(\DLX_EXinst__n0080/FROM ),
    .O(DLX_EXinst__n0080)
  );
  X_BUF \DLX_EXinst__n0080/YUSED  (
    .I(\DLX_EXinst__n0080/GROM ),
    .O(N163390)
  );
  defparam DLX_IDinst_RegFile_19_30_1086.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_19_30_1086 (
    .I(DLX_IDinst_WB_data_eff[30]),
    .CE(DLX_IDinst__n0588),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_19_30)
  );
  defparam DLX_EXinst__n00771.INIT = 16'h1000;
  X_LUT4 DLX_EXinst__n00771 (
    .ADR0(\DLX_IDinst_Imm[0] ),
    .ADR1(\DLX_IDinst_Imm[1] ),
    .ADR2(DLX_EXinst_N76002),
    .ADR3(DLX_IDinst_IR_function_field[5]),
    .O(\DLX_EXinst__n0077/FROM )
  );
  defparam \DLX_EXinst__n0007<31>45 .INIT = 16'hFECE;
  X_LUT4 \DLX_EXinst__n0007<31>45  (
    .ADR0(DLX_EXinst__n0079),
    .ADR1(N163931),
    .ADR2(DLX_IDinst_reg_out_B[31]),
    .ADR3(DLX_EXinst__n0077),
    .O(\DLX_EXinst__n0077/GROM )
  );
  X_BUF \DLX_EXinst__n0077/XUSED  (
    .I(\DLX_EXinst__n0077/FROM ),
    .O(DLX_EXinst__n0077)
  );
  X_BUF \DLX_EXinst__n0077/YUSED  (
    .I(\DLX_EXinst__n0077/GROM ),
    .O(CHOICE5779)
  );
  defparam DLX_EXinst__n00781.INIT = 16'h4000;
  X_LUT4 DLX_EXinst__n00781 (
    .ADR0(\DLX_IDinst_Imm[1] ),
    .ADR1(DLX_IDinst_IR_function_field[5]),
    .ADR2(DLX_EXinst_N76002),
    .ADR3(\DLX_IDinst_Imm[0] ),
    .O(\DLX_EXinst__n0078/FROM )
  );
  defparam \DLX_EXinst__n0007<28>196 .INIT = 16'hCC08;
  X_LUT4 \DLX_EXinst__n0007<28>196  (
    .ADR0(DLX_EXinst__n0079),
    .ADR1(DLX_IDinst_reg_out_B[28]),
    .ADR2(DLX_IDinst_reg_out_A[28]),
    .ADR3(DLX_EXinst__n0078),
    .O(\DLX_EXinst__n0078/GROM )
  );
  X_BUF \DLX_EXinst__n0078/XUSED  (
    .I(\DLX_EXinst__n0078/FROM ),
    .O(DLX_EXinst__n0078)
  );
  X_BUF \DLX_EXinst__n0078/YUSED  (
    .I(\DLX_EXinst__n0078/GROM ),
    .O(CHOICE4886)
  );
  defparam DLX_EXinst__n00791.INIT = 16'h0800;
  X_LUT4 DLX_EXinst__n00791 (
    .ADR0(\DLX_IDinst_Imm[1] ),
    .ADR1(DLX_EXinst_N76002),
    .ADR2(\DLX_IDinst_Imm[0] ),
    .ADR3(DLX_IDinst_IR_function_field[5]),
    .O(\DLX_IDinst_RegFile_0_21/FROM )
  );
  defparam \DLX_EXinst__n0007<4>72 .INIT = 16'hFCCC;
  X_LUT4 \DLX_EXinst__n0007<4>72  (
    .ADR0(VCC),
    .ADR1(CHOICE4341),
    .ADR2(DLX_IDinst_reg_out_A[4]),
    .ADR3(DLX_EXinst__n0079),
    .O(\DLX_IDinst_RegFile_0_21/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_0_21/XUSED  (
    .I(\DLX_IDinst_RegFile_0_21/FROM ),
    .O(DLX_EXinst__n0079)
  );
  X_BUF \DLX_IDinst_RegFile_0_21/YUSED  (
    .I(\DLX_IDinst_RegFile_0_21/GROM ),
    .O(CHOICE4342)
  );
  defparam DLX_IDinst_RegFile_19_14_1087.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_19_14_1087 (
    .I(DLX_IDinst_WB_data_eff[14]),
    .CE(DLX_IDinst__n0588),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_19_14)
  );
  defparam DLX_IDinst_RegFile_27_30_1088.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_27_30_1088 (
    .I(DLX_IDinst_WB_data_eff[30]),
    .CE(DLX_IDinst__n0604),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_27_30)
  );
  X_ZERO \DLX_IDinst_RegFile_4_10/LOGIC_ZERO_1089  (
    .O(\DLX_IDinst_RegFile_4_10/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_162_1090 (
    .IA(\DLX_IDinst_RegFile_4_10/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_4_10/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_221),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_162)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2211.INIT = 16'hFB73;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2211 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_45),
    .ADR2(DLX_IDinst_RegFile_4_10),
    .ADR3(DLX_IDinst_RegFile_5_10),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_221)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2221.INIT = 16'hD8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2221 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR1(DLX_IDinst_RegFile_7_10),
    .ADR2(DLX_IDinst_RegFile_6_10),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_46),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_222)
  );
  X_BUF \DLX_IDinst_RegFile_4_10/COUTUSED  (
    .I(\DLX_IDinst_RegFile_4_10/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_163)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_163_1091 (
    .IA(\DLX_IDinst_RegFile_4_10/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_162),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_222),
    .O(\DLX_IDinst_RegFile_4_10/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_4_10/CYINIT_1092  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_161),
    .O(\DLX_IDinst_RegFile_4_10/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_4_11/LOGIC_ZERO_1093  (
    .O(\DLX_IDinst_RegFile_4_11/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_178_1094 (
    .IA(\DLX_IDinst_RegFile_4_11/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_4_11/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_237),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_178)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2371.INIT = 16'hB8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2371 (
    .ADR0(DLX_IDinst_RegFile_5_11),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR2(DLX_IDinst_RegFile_4_11),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_45),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_237)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2381.INIT = 16'hBF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2381 (
    .ADR0(DLX_IDinst_RegFile_7_11),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_46),
    .ADR3(DLX_IDinst_RegFile_6_11),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_238)
  );
  X_BUF \DLX_IDinst_RegFile_4_11/COUTUSED  (
    .I(\DLX_IDinst_RegFile_4_11/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_179)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_179_1095 (
    .IA(\DLX_IDinst_RegFile_4_11/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_178),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_238),
    .O(\DLX_IDinst_RegFile_4_11/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_4_11/CYINIT_1096  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_177),
    .O(\DLX_IDinst_RegFile_4_11/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_4_12/LOGIC_ZERO_1097  (
    .O(\DLX_IDinst_RegFile_4_12/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_194_1098 (
    .IA(\DLX_IDinst_RegFile_4_12/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_4_12/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_253),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_194)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2531.INIT = 16'hBFB3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2531 (
    .ADR0(DLX_IDinst_RegFile_5_12),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_45),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR3(DLX_IDinst_RegFile_4_12),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_253)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2541.INIT = 16'hDDF5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2541 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_46),
    .ADR1(DLX_IDinst_RegFile_7_12),
    .ADR2(DLX_IDinst_RegFile_6_12),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_254)
  );
  X_BUF \DLX_IDinst_RegFile_4_12/COUTUSED  (
    .I(\DLX_IDinst_RegFile_4_12/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_195)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_195_1099 (
    .IA(\DLX_IDinst_RegFile_4_12/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_194),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_254),
    .O(\DLX_IDinst_RegFile_4_12/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_4_12/CYINIT_1100  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_193),
    .O(\DLX_IDinst_RegFile_4_12/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_4_20/LOGIC_ZERO_1101  (
    .O(\DLX_IDinst_RegFile_4_20/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_322_1102 (
    .IA(\DLX_IDinst_RegFile_4_20/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_4_20/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_381),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_322)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3811.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3811 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_45),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR2(DLX_IDinst_RegFile_4_20),
    .ADR3(DLX_IDinst_RegFile_5_20),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_381)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3821.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3821 (
    .ADR0(DLX_IDinst_RegFile_6_20),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_46),
    .ADR3(DLX_IDinst_RegFile_7_20),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_382)
  );
  X_BUF \DLX_IDinst_RegFile_4_20/COUTUSED  (
    .I(\DLX_IDinst_RegFile_4_20/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_323)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_323_1103 (
    .IA(\DLX_IDinst_RegFile_4_20/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_322),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_382),
    .O(\DLX_IDinst_RegFile_4_20/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_4_20/CYINIT_1104  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_321),
    .O(\DLX_IDinst_RegFile_4_20/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_4_13/LOGIC_ZERO_1105  (
    .O(\DLX_IDinst_RegFile_4_13/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_210_1106 (
    .IA(\DLX_IDinst_RegFile_4_13/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_4_13/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_269),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_210)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2691.INIT = 16'hBFB3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2691 (
    .ADR0(DLX_IDinst_RegFile_5_13),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_45),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR3(DLX_IDinst_RegFile_4_13),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_269)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2701.INIT = 16'hDFD5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2701 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_46),
    .ADR1(DLX_IDinst_RegFile_7_13),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR3(DLX_IDinst_RegFile_6_13),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_270)
  );
  X_BUF \DLX_IDinst_RegFile_4_13/COUTUSED  (
    .I(\DLX_IDinst_RegFile_4_13/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_211)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_211_1107 (
    .IA(\DLX_IDinst_RegFile_4_13/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_210),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_270),
    .O(\DLX_IDinst_RegFile_4_13/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_4_13/CYINIT_1108  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_209),
    .O(\DLX_IDinst_RegFile_4_13/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_4_21/LOGIC_ZERO_1109  (
    .O(\DLX_IDinst_RegFile_4_21/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_338_1110 (
    .IA(\DLX_IDinst_RegFile_4_21/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_4_21/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_397),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_338)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3971.INIT = 16'hAFCF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3971 (
    .ADR0(DLX_IDinst_RegFile_5_21),
    .ADR1(DLX_IDinst_RegFile_4_21),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_45),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_397)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3981.INIT = 16'hBF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3981 (
    .ADR0(DLX_IDinst_RegFile_7_21),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_46),
    .ADR3(DLX_IDinst_RegFile_6_21),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_398)
  );
  X_BUF \DLX_IDinst_RegFile_4_21/COUTUSED  (
    .I(\DLX_IDinst_RegFile_4_21/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_339)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_339_1111 (
    .IA(\DLX_IDinst_RegFile_4_21/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_338),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_398),
    .O(\DLX_IDinst_RegFile_4_21/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_4_21/CYINIT_1112  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_337),
    .O(\DLX_IDinst_RegFile_4_21/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_4_14/LOGIC_ZERO_1113  (
    .O(\DLX_IDinst_RegFile_4_14/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_226_1114 (
    .IA(\DLX_IDinst_RegFile_4_14/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_4_14/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_285),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_226)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2851.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2851 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_45),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR2(DLX_IDinst_RegFile_4_14),
    .ADR3(DLX_IDinst_RegFile_5_14),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_285)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2861.INIT = 16'hB8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2861 (
    .ADR0(DLX_IDinst_RegFile_7_14),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR2(DLX_IDinst_RegFile_6_14),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_46),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_286)
  );
  X_BUF \DLX_IDinst_RegFile_4_14/COUTUSED  (
    .I(\DLX_IDinst_RegFile_4_14/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_227)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_227_1115 (
    .IA(\DLX_IDinst_RegFile_4_14/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_226),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_286),
    .O(\DLX_IDinst_RegFile_4_14/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_4_14/CYINIT_1116  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_225),
    .O(\DLX_IDinst_RegFile_4_14/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_4_22/LOGIC_ZERO_1117  (
    .O(\DLX_IDinst_RegFile_4_22/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_354_1118 (
    .IA(\DLX_IDinst_RegFile_4_22/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_4_22/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_413),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_354)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4131.INIT = 16'hDF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4131 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR1(DLX_IDinst_RegFile_5_22),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_45),
    .ADR3(DLX_IDinst_RegFile_4_22),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_413)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4141.INIT = 16'hE4FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4141 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR1(DLX_IDinst_RegFile_6_22),
    .ADR2(DLX_IDinst_RegFile_7_22),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_46),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_414)
  );
  X_BUF \DLX_IDinst_RegFile_4_22/COUTUSED  (
    .I(\DLX_IDinst_RegFile_4_22/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_355)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_355_1119 (
    .IA(\DLX_IDinst_RegFile_4_22/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_354),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_414),
    .O(\DLX_IDinst_RegFile_4_22/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_4_22/CYINIT_1120  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_353),
    .O(\DLX_IDinst_RegFile_4_22/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_4_30/LOGIC_ZERO_1121  (
    .O(\DLX_IDinst_RegFile_4_30/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_994_1122 (
    .IA(\DLX_IDinst_RegFile_4_30/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_4_30/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1069),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_994)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10691.INIT = 16'hFD5D;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10691 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_573),
    .ADR1(DLX_IDinst_RegFile_4_30),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR3(DLX_IDinst_RegFile_5_30),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1069)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10701.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10701 (
    .ADR0(DLX_IDinst_RegFile_6_30),
    .ADR1(DLX_IDinst_RegFile_7_30),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_574),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1070)
  );
  X_BUF \DLX_IDinst_RegFile_4_30/COUTUSED  (
    .I(\DLX_IDinst_RegFile_4_30/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_995)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_995_1123 (
    .IA(\DLX_IDinst_RegFile_4_30/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_994),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1070),
    .O(\DLX_IDinst_RegFile_4_30/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_4_30/CYINIT_1124  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_993),
    .O(\DLX_IDinst_RegFile_4_30/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_4_31/LOGIC_ZERO_1125  (
    .O(\DLX_IDinst_RegFile_4_31/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_1010_1126 (
    .IA(\DLX_IDinst_RegFile_4_31/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_4_31/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1085),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_1010)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10851.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10851 (
    .ADR0(DLX_IDinst_RegFile_4_31),
    .ADR1(DLX_IDinst_RegFile_5_31),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_573),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1085)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10861.INIT = 16'hCFAF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10861 (
    .ADR0(DLX_IDinst_RegFile_6_31),
    .ADR1(DLX_IDinst_RegFile_7_31),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_574),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1086)
  );
  X_BUF \DLX_IDinst_RegFile_4_31/COUTUSED  (
    .I(\DLX_IDinst_RegFile_4_31/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_1011)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_1011_1127 (
    .IA(\DLX_IDinst_RegFile_4_31/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_1010),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1086),
    .O(\DLX_IDinst_RegFile_4_31/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_4_31/CYINIT_1128  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_1009),
    .O(\DLX_IDinst_RegFile_4_31/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_4_15/LOGIC_ZERO_1129  (
    .O(\DLX_IDinst_RegFile_4_15/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_242_1130 (
    .IA(\DLX_IDinst_RegFile_4_15/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_4_15/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_301),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_242)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3011.INIT = 16'hACFF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3011 (
    .ADR0(DLX_IDinst_RegFile_5_15),
    .ADR1(DLX_IDinst_RegFile_4_15),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_45),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_301)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3021.INIT = 16'hCFAF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3021 (
    .ADR0(DLX_IDinst_RegFile_6_15),
    .ADR1(DLX_IDinst_RegFile_7_15),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_46),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_302)
  );
  X_BUF \DLX_IDinst_RegFile_4_15/COUTUSED  (
    .I(\DLX_IDinst_RegFile_4_15/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_243)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_243_1131 (
    .IA(\DLX_IDinst_RegFile_4_15/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_242),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_302),
    .O(\DLX_IDinst_RegFile_4_15/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_4_15/CYINIT_1132  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_241),
    .O(\DLX_IDinst_RegFile_4_15/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_4_23/LOGIC_ZERO_1133  (
    .O(\DLX_IDinst_RegFile_4_23/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_370_1134 (
    .IA(\DLX_IDinst_RegFile_4_23/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_4_23/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_429),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_370)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4291.INIT = 16'hFB73;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4291 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_45),
    .ADR2(DLX_IDinst_RegFile_4_23),
    .ADR3(DLX_IDinst_RegFile_5_23),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_429)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4301.INIT = 16'hAFCF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4301 (
    .ADR0(DLX_IDinst_RegFile_7_23),
    .ADR1(DLX_IDinst_RegFile_6_23),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_46),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_430)
  );
  X_BUF \DLX_IDinst_RegFile_4_23/COUTUSED  (
    .I(\DLX_IDinst_RegFile_4_23/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_371)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_371_1135 (
    .IA(\DLX_IDinst_RegFile_4_23/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_370),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_430),
    .O(\DLX_IDinst_RegFile_4_23/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_4_23/CYINIT_1136  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_369),
    .O(\DLX_IDinst_RegFile_4_23/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_4_16/LOGIC_ZERO_1137  (
    .O(\DLX_IDinst_RegFile_4_16/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_258_1138 (
    .IA(\DLX_IDinst_RegFile_4_16/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_4_16/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_317),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_258)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3171.INIT = 16'hF5DD;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3171 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_45),
    .ADR1(DLX_IDinst_RegFile_4_16),
    .ADR2(DLX_IDinst_RegFile_5_16),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_317)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3181.INIT = 16'hFD5D;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3181 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_46),
    .ADR1(DLX_IDinst_RegFile_6_16),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR3(DLX_IDinst_RegFile_7_16),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_318)
  );
  X_BUF \DLX_IDinst_RegFile_4_16/COUTUSED  (
    .I(\DLX_IDinst_RegFile_4_16/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_259)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_259_1139 (
    .IA(\DLX_IDinst_RegFile_4_16/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_258),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_318),
    .O(\DLX_IDinst_RegFile_4_16/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_4_16/CYINIT_1140  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_257),
    .O(\DLX_IDinst_RegFile_4_16/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_4_24/LOGIC_ZERO_1141  (
    .O(\DLX_IDinst_RegFile_4_24/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_386_1142 (
    .IA(\DLX_IDinst_RegFile_4_24/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_4_24/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_445),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_386)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4451.INIT = 16'hF5DD;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4451 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_45),
    .ADR1(DLX_IDinst_RegFile_4_24),
    .ADR2(DLX_IDinst_RegFile_5_24),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_445)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4461.INIT = 16'hE2FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4461 (
    .ADR0(DLX_IDinst_RegFile_6_24),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR2(DLX_IDinst_RegFile_7_24),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_46),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_446)
  );
  X_BUF \DLX_IDinst_RegFile_4_24/COUTUSED  (
    .I(\DLX_IDinst_RegFile_4_24/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_387)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_387_1143 (
    .IA(\DLX_IDinst_RegFile_4_24/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_386),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_446),
    .O(\DLX_IDinst_RegFile_4_24/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_4_24/CYINIT_1144  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_385),
    .O(\DLX_IDinst_RegFile_4_24/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_4_17/LOGIC_ZERO_1145  (
    .O(\DLX_IDinst_RegFile_4_17/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_274_1146 (
    .IA(\DLX_IDinst_RegFile_4_17/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_4_17/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_333),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_274)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3331.INIT = 16'hF7D5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3331 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_45),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR2(DLX_IDinst_RegFile_5_17),
    .ADR3(DLX_IDinst_RegFile_4_17),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_333)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3341.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3341 (
    .ADR0(DLX_IDinst_RegFile_6_17),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_46),
    .ADR3(DLX_IDinst_RegFile_7_17),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_334)
  );
  X_BUF \DLX_IDinst_RegFile_4_17/COUTUSED  (
    .I(\DLX_IDinst_RegFile_4_17/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_275)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_275_1147 (
    .IA(\DLX_IDinst_RegFile_4_17/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_274),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_334),
    .O(\DLX_IDinst_RegFile_4_17/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_4_17/CYINIT_1148  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_273),
    .O(\DLX_IDinst_RegFile_4_17/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_4_25/LOGIC_ZERO_1149  (
    .O(\DLX_IDinst_RegFile_4_25/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_402_1150 (
    .IA(\DLX_IDinst_RegFile_4_25/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_4_25/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_461),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_402)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4611.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4611 (
    .ADR0(DLX_IDinst_RegFile_4_25),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_45),
    .ADR3(DLX_IDinst_RegFile_5_25),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_461)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4621.INIT = 16'hFD5D;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4621 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_46),
    .ADR1(DLX_IDinst_RegFile_6_25),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR3(DLX_IDinst_RegFile_7_25),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_462)
  );
  X_BUF \DLX_IDinst_RegFile_4_25/COUTUSED  (
    .I(\DLX_IDinst_RegFile_4_25/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_403)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_403_1151 (
    .IA(\DLX_IDinst_RegFile_4_25/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_402),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_462),
    .O(\DLX_IDinst_RegFile_4_25/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_4_25/CYINIT_1152  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_401),
    .O(\DLX_IDinst_RegFile_4_25/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_4_18/LOGIC_ZERO_1153  (
    .O(\DLX_IDinst_RegFile_4_18/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_290_1154 (
    .IA(\DLX_IDinst_RegFile_4_18/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_4_18/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_349),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_290)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3491.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3491 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR1(DLX_IDinst_RegFile_4_18),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_45),
    .ADR3(DLX_IDinst_RegFile_5_18),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_349)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3501.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3501 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_46),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR2(DLX_IDinst_RegFile_6_18),
    .ADR3(DLX_IDinst_RegFile_7_18),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_350)
  );
  X_BUF \DLX_IDinst_RegFile_4_18/COUTUSED  (
    .I(\DLX_IDinst_RegFile_4_18/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_291)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_291_1155 (
    .IA(\DLX_IDinst_RegFile_4_18/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_290),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_350),
    .O(\DLX_IDinst_RegFile_4_18/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_4_18/CYINIT_1156  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_289),
    .O(\DLX_IDinst_RegFile_4_18/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_4_26/LOGIC_ZERO_1157  (
    .O(\DLX_IDinst_RegFile_4_26/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_418_1158 (
    .IA(\DLX_IDinst_RegFile_4_26/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_4_26/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_477),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_418)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4771.INIT = 16'hBFB3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4771 (
    .ADR0(DLX_IDinst_RegFile_5_26),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_45),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR3(DLX_IDinst_RegFile_4_26),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_477)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4781.INIT = 16'hDDF5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4781 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_46),
    .ADR1(DLX_IDinst_RegFile_7_26),
    .ADR2(DLX_IDinst_RegFile_6_26),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_478)
  );
  X_BUF \DLX_IDinst_RegFile_4_26/COUTUSED  (
    .I(\DLX_IDinst_RegFile_4_26/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_419)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_419_1159 (
    .IA(\DLX_IDinst_RegFile_4_26/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_418),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_478),
    .O(\DLX_IDinst_RegFile_4_26/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_4_26/CYINIT_1160  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_417),
    .O(\DLX_IDinst_RegFile_4_26/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_5_10/LOGIC_ZERO_1161  (
    .O(\DLX_IDinst_RegFile_5_10/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_674_1162 (
    .IA(\DLX_IDinst_RegFile_5_10/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_5_10/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_749),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_674)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7491.INIT = 16'hD8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7491 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR1(DLX_IDinst_RegFile_5_10),
    .ADR2(DLX_IDinst_RegFile_4_10),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_573),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_749)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7501.INIT = 16'hD8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7501 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR1(DLX_IDinst_RegFile_7_10),
    .ADR2(DLX_IDinst_RegFile_6_10),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_574),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_750)
  );
  X_BUF \DLX_IDinst_RegFile_5_10/COUTUSED  (
    .I(\DLX_IDinst_RegFile_5_10/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_675)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_675_1163 (
    .IA(\DLX_IDinst_RegFile_5_10/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_674),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_750),
    .O(\DLX_IDinst_RegFile_5_10/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_5_10/CYINIT_1164  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_673),
    .O(\DLX_IDinst_RegFile_5_10/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_4_19/LOGIC_ZERO_1165  (
    .O(\DLX_IDinst_RegFile_4_19/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_306_1166 (
    .IA(\DLX_IDinst_RegFile_4_19/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_4_19/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_365),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_306)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3651.INIT = 16'hDFD5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3651 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_45),
    .ADR1(DLX_IDinst_RegFile_5_19),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR3(DLX_IDinst_RegFile_4_19),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_365)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3661.INIT = 16'hACFF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3661 (
    .ADR0(DLX_IDinst_RegFile_7_19),
    .ADR1(DLX_IDinst_RegFile_6_19),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_46),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_366)
  );
  X_BUF \DLX_IDinst_RegFile_4_19/COUTUSED  (
    .I(\DLX_IDinst_RegFile_4_19/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_307)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_307_1167 (
    .IA(\DLX_IDinst_RegFile_4_19/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_306),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_366),
    .O(\DLX_IDinst_RegFile_4_19/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_4_19/CYINIT_1168  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_305),
    .O(\DLX_IDinst_RegFile_4_19/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_4_27/LOGIC_ZERO_1169  (
    .O(\DLX_IDinst_RegFile_4_27/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_434_1170 (
    .IA(\DLX_IDinst_RegFile_4_27/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_4_27/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_493),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_434)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4931.INIT = 16'hBFB3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4931 (
    .ADR0(DLX_IDinst_RegFile_5_27),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_45),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR3(DLX_IDinst_RegFile_4_27),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_493)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4941.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4941 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR1(DLX_IDinst_RegFile_6_27),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_46),
    .ADR3(DLX_IDinst_RegFile_7_27),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_494)
  );
  X_BUF \DLX_IDinst_RegFile_4_27/COUTUSED  (
    .I(\DLX_IDinst_RegFile_4_27/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_435)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_435_1171 (
    .IA(\DLX_IDinst_RegFile_4_27/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_434),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_494),
    .O(\DLX_IDinst_RegFile_4_27/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_4_27/CYINIT_1172  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_433),
    .O(\DLX_IDinst_RegFile_4_27/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_5_11/LOGIC_ZERO_1173  (
    .O(\DLX_IDinst_RegFile_5_11/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_690_1174 (
    .IA(\DLX_IDinst_RegFile_5_11/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_5_11/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_765),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_690)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7651.INIT = 16'hF5DD;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7651 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_573),
    .ADR1(DLX_IDinst_RegFile_4_11),
    .ADR2(DLX_IDinst_RegFile_5_11),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_765)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7661.INIT = 16'hBFB3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7661 (
    .ADR0(DLX_IDinst_RegFile_7_11),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_574),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR3(DLX_IDinst_RegFile_6_11),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_766)
  );
  X_BUF \DLX_IDinst_RegFile_5_11/COUTUSED  (
    .I(\DLX_IDinst_RegFile_5_11/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_691)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_691_1175 (
    .IA(\DLX_IDinst_RegFile_5_11/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_690),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_766),
    .O(\DLX_IDinst_RegFile_5_11/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_5_11/CYINIT_1176  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_689),
    .O(\DLX_IDinst_RegFile_5_11/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_4_28/LOGIC_ZERO_1177  (
    .O(\DLX_IDinst_RegFile_4_28/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_962_1178 (
    .IA(\DLX_IDinst_RegFile_4_28/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_4_28/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1037),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_962)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10371.INIT = 16'hAFCF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10371 (
    .ADR0(DLX_IDinst_RegFile_5_28),
    .ADR1(DLX_IDinst_RegFile_4_28),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_573),
    .ADR3(DLX_IDinst_jtarget[21]),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1037)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10381.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10381 (
    .ADR0(DLX_IDinst_RegFile_7_28),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_574),
    .ADR2(DLX_IDinst_RegFile_6_28),
    .ADR3(DLX_IDinst_jtarget[21]),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1038)
  );
  X_BUF \DLX_IDinst_RegFile_4_28/COUTUSED  (
    .I(\DLX_IDinst_RegFile_4_28/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_963)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_963_1179 (
    .IA(\DLX_IDinst_RegFile_4_28/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_962),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1038),
    .O(\DLX_IDinst_RegFile_4_28/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_4_28/CYINIT_1180  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_961),
    .O(\DLX_IDinst_RegFile_4_28/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_5_20/LOGIC_ZERO_1181  (
    .O(\DLX_IDinst_RegFile_5_20/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_834_1182 (
    .IA(\DLX_IDinst_RegFile_5_20/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_5_20/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_909),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_834)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9091.INIT = 16'hF7B3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9091 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_573),
    .ADR2(DLX_IDinst_RegFile_5_20),
    .ADR3(DLX_IDinst_RegFile_4_20),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_909)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9101.INIT = 16'hDF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9101 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR1(DLX_IDinst_RegFile_7_20),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_574),
    .ADR3(DLX_IDinst_RegFile_6_20),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_910)
  );
  X_BUF \DLX_IDinst_RegFile_5_20/COUTUSED  (
    .I(\DLX_IDinst_RegFile_5_20/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_835)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_835_1183 (
    .IA(\DLX_IDinst_RegFile_5_20/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_834),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_910),
    .O(\DLX_IDinst_RegFile_5_20/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_5_20/CYINIT_1184  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_833),
    .O(\DLX_IDinst_RegFile_5_20/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_5_12/LOGIC_ZERO_1185  (
    .O(\DLX_IDinst_RegFile_5_12/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_706_1186 (
    .IA(\DLX_IDinst_RegFile_5_12/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_5_12/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_781),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_706)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7811.INIT = 16'hE4FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7811 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR1(DLX_IDinst_RegFile_4_12),
    .ADR2(DLX_IDinst_RegFile_5_12),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_573),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_781)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7821.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7821 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR1(DLX_IDinst_RegFile_6_12),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_574),
    .ADR3(DLX_IDinst_RegFile_7_12),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_782)
  );
  X_BUF \DLX_IDinst_RegFile_5_12/COUTUSED  (
    .I(\DLX_IDinst_RegFile_5_12/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_707)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_707_1187 (
    .IA(\DLX_IDinst_RegFile_5_12/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_706),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_782),
    .O(\DLX_IDinst_RegFile_5_12/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_5_12/CYINIT_1188  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_705),
    .O(\DLX_IDinst_RegFile_5_12/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_4_29/LOGIC_ZERO_1189  (
    .O(\DLX_IDinst_RegFile_4_29/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_978_1190 (
    .IA(\DLX_IDinst_RegFile_4_29/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_4_29/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1053),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_978)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10531.INIT = 16'hDF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10531 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR1(DLX_IDinst_RegFile_5_29),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_573),
    .ADR3(DLX_IDinst_RegFile_4_29),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1053)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10541.INIT = 16'hAFCF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10541 (
    .ADR0(DLX_IDinst_RegFile_7_29),
    .ADR1(DLX_IDinst_RegFile_6_29),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_574),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1054)
  );
  X_BUF \DLX_IDinst_RegFile_4_29/COUTUSED  (
    .I(\DLX_IDinst_RegFile_4_29/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_979)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_979_1191 (
    .IA(\DLX_IDinst_RegFile_4_29/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_978),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1054),
    .O(\DLX_IDinst_RegFile_4_29/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_4_29/CYINIT_1192  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_977),
    .O(\DLX_IDinst_RegFile_4_29/CYINIT )
  );
  defparam DLX_IDinst_RegFile_27_22_1193.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_27_22_1193 (
    .I(DLX_IDinst_WB_data_eff[22]),
    .CE(DLX_IDinst__n0604),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_27_22)
  );
  X_ZERO \DLX_IDinst_RegFile_5_21/LOGIC_ZERO_1194  (
    .O(\DLX_IDinst_RegFile_5_21/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_850_1195 (
    .IA(\DLX_IDinst_RegFile_5_21/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_5_21/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_925),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_850)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9251.INIT = 16'hE4FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9251 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR1(DLX_IDinst_RegFile_4_21),
    .ADR2(DLX_IDinst_RegFile_5_21),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_573),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_925)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9261.INIT = 16'hFB3B;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9261 (
    .ADR0(DLX_IDinst_RegFile_6_21),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_574),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR3(DLX_IDinst_RegFile_7_21),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_926)
  );
  X_BUF \DLX_IDinst_RegFile_5_21/COUTUSED  (
    .I(\DLX_IDinst_RegFile_5_21/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_851)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_851_1196 (
    .IA(\DLX_IDinst_RegFile_5_21/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_850),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_926),
    .O(\DLX_IDinst_RegFile_5_21/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_5_21/CYINIT_1197  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_849),
    .O(\DLX_IDinst_RegFile_5_21/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_5_13/LOGIC_ZERO_1198  (
    .O(\DLX_IDinst_RegFile_5_13/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_722_1199 (
    .IA(\DLX_IDinst_RegFile_5_13/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_5_13/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_797),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_722)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7971.INIT = 16'hF7B3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7971 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_573),
    .ADR2(DLX_IDinst_RegFile_5_13),
    .ADR3(DLX_IDinst_RegFile_4_13),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_797)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7981.INIT = 16'hDF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7981 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR1(DLX_IDinst_RegFile_7_13),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_574),
    .ADR3(DLX_IDinst_RegFile_6_13),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_798)
  );
  X_BUF \DLX_IDinst_RegFile_5_13/COUTUSED  (
    .I(\DLX_IDinst_RegFile_5_13/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_723)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_723_1200 (
    .IA(\DLX_IDinst_RegFile_5_13/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_722),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_798),
    .O(\DLX_IDinst_RegFile_5_13/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_5_13/CYINIT_1201  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_721),
    .O(\DLX_IDinst_RegFile_5_13/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_5_30/LOGIC_ZERO_1202  (
    .O(\DLX_IDinst_RegFile_5_30/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_482_1203 (
    .IA(\DLX_IDinst_RegFile_5_30/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_5_30/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_541),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_482)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5411.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5411 (
    .ADR0(DLX_IDinst_RegFile_5_30),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_45),
    .ADR2(DLX_IDinst_RegFile_4_30),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_541)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5421.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5421 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_46),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR2(DLX_IDinst_RegFile_6_30),
    .ADR3(DLX_IDinst_RegFile_7_30),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_542)
  );
  X_BUF \DLX_IDinst_RegFile_5_30/COUTUSED  (
    .I(\DLX_IDinst_RegFile_5_30/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_483)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_483_1204 (
    .IA(\DLX_IDinst_RegFile_5_30/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_482),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_542),
    .O(\DLX_IDinst_RegFile_5_30/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_5_30/CYINIT_1205  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_481),
    .O(\DLX_IDinst_RegFile_5_30/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_5_22/LOGIC_ZERO_1206  (
    .O(\DLX_IDinst_RegFile_5_22/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_866_1207 (
    .IA(\DLX_IDinst_RegFile_5_22/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_5_22/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_941),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_866)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9411.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9411 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_573),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR2(DLX_IDinst_RegFile_4_22),
    .ADR3(DLX_IDinst_RegFile_5_22),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_941)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9421.INIT = 16'hDDF5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9421 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_574),
    .ADR1(DLX_IDinst_RegFile_7_22),
    .ADR2(DLX_IDinst_RegFile_6_22),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_942)
  );
  X_BUF \DLX_IDinst_RegFile_5_22/COUTUSED  (
    .I(\DLX_IDinst_RegFile_5_22/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_867)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_867_1208 (
    .IA(\DLX_IDinst_RegFile_5_22/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_866),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_942),
    .O(\DLX_IDinst_RegFile_5_22/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_5_22/CYINIT_1209  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_865),
    .O(\DLX_IDinst_RegFile_5_22/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_5_14/LOGIC_ZERO_1210  (
    .O(\DLX_IDinst_RegFile_5_14/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_738_1211 (
    .IA(\DLX_IDinst_RegFile_5_14/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_5_14/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_813),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_738)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8131.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8131 (
    .ADR0(DLX_IDinst_RegFile_4_14),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_573),
    .ADR2(DLX_IDinst_RegFile_5_14),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_813)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8141.INIT = 16'hDDF5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8141 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_574),
    .ADR1(DLX_IDinst_RegFile_7_14),
    .ADR2(DLX_IDinst_RegFile_6_14),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_814)
  );
  X_BUF \DLX_IDinst_RegFile_5_14/COUTUSED  (
    .I(\DLX_IDinst_RegFile_5_14/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_739)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_739_1212 (
    .IA(\DLX_IDinst_RegFile_5_14/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_738),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_814),
    .O(\DLX_IDinst_RegFile_5_14/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_5_14/CYINIT_1213  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_737),
    .O(\DLX_IDinst_RegFile_5_14/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_5_31/LOGIC_ZERO_1214  (
    .O(\DLX_IDinst_RegFile_5_31/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_498_1215 (
    .IA(\DLX_IDinst_RegFile_5_31/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_5_31/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_557),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_498)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5571.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5571 (
    .ADR0(DLX_IDinst_RegFile_4_31),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_45),
    .ADR3(DLX_IDinst_RegFile_5_31),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_557)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5581.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5581 (
    .ADR0(DLX_IDinst_RegFile_6_31),
    .ADR1(DLX_IDinst_RegFile_7_31),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_46),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_558)
  );
  X_BUF \DLX_IDinst_RegFile_5_31/COUTUSED  (
    .I(\DLX_IDinst_RegFile_5_31/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_499)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_499_1216 (
    .IA(\DLX_IDinst_RegFile_5_31/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_498),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_558),
    .O(\DLX_IDinst_RegFile_5_31/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_5_31/CYINIT_1217  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_497),
    .O(\DLX_IDinst_RegFile_5_31/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_5_23/LOGIC_ZERO_1218  (
    .O(\DLX_IDinst_RegFile_5_23/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_882_1219 (
    .IA(\DLX_IDinst_RegFile_5_23/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_5_23/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_957),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_882)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9571.INIT = 16'hCFAF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9571 (
    .ADR0(DLX_IDinst_RegFile_4_23),
    .ADR1(DLX_IDinst_RegFile_5_23),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_573),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_957)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9581.INIT = 16'hAFCF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9581 (
    .ADR0(DLX_IDinst_RegFile_7_23),
    .ADR1(DLX_IDinst_RegFile_6_23),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_574),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_958)
  );
  X_BUF \DLX_IDinst_RegFile_5_23/COUTUSED  (
    .I(\DLX_IDinst_RegFile_5_23/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_883)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_883_1220 (
    .IA(\DLX_IDinst_RegFile_5_23/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_882),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_958),
    .O(\DLX_IDinst_RegFile_5_23/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_5_23/CYINIT_1221  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_881),
    .O(\DLX_IDinst_RegFile_5_23/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_5_15/LOGIC_ZERO_1222  (
    .O(\DLX_IDinst_RegFile_5_15/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_754_1223 (
    .IA(\DLX_IDinst_RegFile_5_15/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_5_15/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_829),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_754)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8291.INIT = 16'hCFAF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8291 (
    .ADR0(DLX_IDinst_RegFile_4_15),
    .ADR1(DLX_IDinst_RegFile_5_15),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_573),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_829)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8301.INIT = 16'hFB3B;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8301 (
    .ADR0(DLX_IDinst_RegFile_6_15),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_574),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR3(DLX_IDinst_RegFile_7_15),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_830)
  );
  X_BUF \DLX_IDinst_RegFile_5_15/COUTUSED  (
    .I(\DLX_IDinst_RegFile_5_15/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_755)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_755_1224 (
    .IA(\DLX_IDinst_RegFile_5_15/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_754),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_830),
    .O(\DLX_IDinst_RegFile_5_15/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_5_15/CYINIT_1225  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_753),
    .O(\DLX_IDinst_RegFile_5_15/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_5_24/LOGIC_ZERO_1226  (
    .O(\DLX_IDinst_RegFile_5_24/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_898_1227 (
    .IA(\DLX_IDinst_RegFile_5_24/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_5_24/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_973),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_898)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9731.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9731 (
    .ADR0(DLX_IDinst_RegFile_4_24),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_573),
    .ADR3(DLX_IDinst_RegFile_5_24),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_973)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9741.INIT = 16'hDF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9741 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR1(DLX_IDinst_RegFile_7_24),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_574),
    .ADR3(DLX_IDinst_RegFile_6_24),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_974)
  );
  X_BUF \DLX_IDinst_RegFile_5_24/COUTUSED  (
    .I(\DLX_IDinst_RegFile_5_24/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_899)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_899_1228 (
    .IA(\DLX_IDinst_RegFile_5_24/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_898),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_974),
    .O(\DLX_IDinst_RegFile_5_24/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_5_24/CYINIT_1229  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_897),
    .O(\DLX_IDinst_RegFile_5_24/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_5_16/LOGIC_ZERO_1230  (
    .O(\DLX_IDinst_RegFile_5_16/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_770_1231 (
    .IA(\DLX_IDinst_RegFile_5_16/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_5_16/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_845),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_770)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8451.INIT = 16'hFB3B;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8451 (
    .ADR0(DLX_IDinst_RegFile_4_16),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_573),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR3(DLX_IDinst_RegFile_5_16),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_845)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8461.INIT = 16'hBFB3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8461 (
    .ADR0(DLX_IDinst_RegFile_7_16),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_574),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR3(DLX_IDinst_RegFile_6_16),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_846)
  );
  X_BUF \DLX_IDinst_RegFile_5_16/COUTUSED  (
    .I(\DLX_IDinst_RegFile_5_16/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_771)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_771_1232 (
    .IA(\DLX_IDinst_RegFile_5_16/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_770),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_846),
    .O(\DLX_IDinst_RegFile_5_16/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_5_16/CYINIT_1233  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_769),
    .O(\DLX_IDinst_RegFile_5_16/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_5_25/LOGIC_ZERO_1234  (
    .O(\DLX_IDinst_RegFile_5_25/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_914_1235 (
    .IA(\DLX_IDinst_RegFile_5_25/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_5_25/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_989),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_914)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9891.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9891 (
    .ADR0(DLX_IDinst_RegFile_4_25),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_573),
    .ADR2(DLX_IDinst_RegFile_5_25),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_989)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9901.INIT = 16'hF5DD;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9901 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_574),
    .ADR1(DLX_IDinst_RegFile_6_25),
    .ADR2(DLX_IDinst_RegFile_7_25),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_990)
  );
  X_BUF \DLX_IDinst_RegFile_5_25/COUTUSED  (
    .I(\DLX_IDinst_RegFile_5_25/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_915)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_915_1236 (
    .IA(\DLX_IDinst_RegFile_5_25/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_914),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_990),
    .O(\DLX_IDinst_RegFile_5_25/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_5_25/CYINIT_1237  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_913),
    .O(\DLX_IDinst_RegFile_5_25/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_5_17/LOGIC_ZERO_1238  (
    .O(\DLX_IDinst_RegFile_5_17/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_786_1239 (
    .IA(\DLX_IDinst_RegFile_5_17/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_5_17/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_861),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_786)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8611.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8611 (
    .ADR0(DLX_IDinst_RegFile_4_17),
    .ADR1(DLX_IDinst_RegFile_5_17),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_573),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_861)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8621.INIT = 16'hDFD5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8621 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_574),
    .ADR1(DLX_IDinst_RegFile_7_17),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR3(DLX_IDinst_RegFile_6_17),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_862)
  );
  X_BUF \DLX_IDinst_RegFile_5_17/COUTUSED  (
    .I(\DLX_IDinst_RegFile_5_17/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_787)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_787_1240 (
    .IA(\DLX_IDinst_RegFile_5_17/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_786),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_862),
    .O(\DLX_IDinst_RegFile_5_17/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_5_17/CYINIT_1241  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_785),
    .O(\DLX_IDinst_RegFile_5_17/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_5_26/LOGIC_ZERO_1242  (
    .O(\DLX_IDinst_RegFile_5_26/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_930_1243 (
    .IA(\DLX_IDinst_RegFile_5_26/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_5_26/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1005),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_930)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10051.INIT = 16'hBFB3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10051 (
    .ADR0(DLX_IDinst_RegFile_5_26),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_573),
    .ADR2(DLX_IDinst_jtarget[21]),
    .ADR3(DLX_IDinst_RegFile_4_26),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1005)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10061.INIT = 16'hBFB3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10061 (
    .ADR0(DLX_IDinst_RegFile_7_26),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_574),
    .ADR2(DLX_IDinst_jtarget[21]),
    .ADR3(DLX_IDinst_RegFile_6_26),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1006)
  );
  X_BUF \DLX_IDinst_RegFile_5_26/COUTUSED  (
    .I(\DLX_IDinst_RegFile_5_26/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_931)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_931_1244 (
    .IA(\DLX_IDinst_RegFile_5_26/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_930),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1006),
    .O(\DLX_IDinst_RegFile_5_26/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_5_26/CYINIT_1245  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_929),
    .O(\DLX_IDinst_RegFile_5_26/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_5_18/LOGIC_ZERO_1246  (
    .O(\DLX_IDinst_RegFile_5_18/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_802_1247 (
    .IA(\DLX_IDinst_RegFile_5_18/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_5_18/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_877),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_802)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8771.INIT = 16'hF5DD;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8771 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_573),
    .ADR1(DLX_IDinst_RegFile_4_18),
    .ADR2(DLX_IDinst_RegFile_5_18),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_877)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8781.INIT = 16'hFB73;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8781 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_574),
    .ADR2(DLX_IDinst_RegFile_6_18),
    .ADR3(DLX_IDinst_RegFile_7_18),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_878)
  );
  X_BUF \DLX_IDinst_RegFile_5_18/COUTUSED  (
    .I(\DLX_IDinst_RegFile_5_18/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_803)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_803_1248 (
    .IA(\DLX_IDinst_RegFile_5_18/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_802),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_878),
    .O(\DLX_IDinst_RegFile_5_18/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_5_18/CYINIT_1249  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_801),
    .O(\DLX_IDinst_RegFile_5_18/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_5_27/LOGIC_ZERO_1250  (
    .O(\DLX_IDinst_RegFile_5_27/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_946_1251 (
    .IA(\DLX_IDinst_RegFile_5_27/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_5_27/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1021),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_946)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10211.INIT = 16'hAFCF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10211 (
    .ADR0(DLX_IDinst_RegFile_5_27),
    .ADR1(DLX_IDinst_RegFile_4_27),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_573),
    .ADR3(DLX_IDinst_jtarget[21]),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1021)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10221.INIT = 16'hE2FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10221 (
    .ADR0(DLX_IDinst_RegFile_6_27),
    .ADR1(DLX_IDinst_jtarget[21]),
    .ADR2(DLX_IDinst_RegFile_7_27),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_574),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1022)
  );
  X_BUF \DLX_IDinst_RegFile_5_27/COUTUSED  (
    .I(\DLX_IDinst_RegFile_5_27/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_947)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_947_1252 (
    .IA(\DLX_IDinst_RegFile_5_27/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_946),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1022),
    .O(\DLX_IDinst_RegFile_5_27/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_5_27/CYINIT_1253  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_945),
    .O(\DLX_IDinst_RegFile_5_27/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_5_19/LOGIC_ZERO_1254  (
    .O(\DLX_IDinst_RegFile_5_19/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_818_1255 (
    .IA(\DLX_IDinst_RegFile_5_19/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_5_19/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_893),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_818)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8931.INIT = 16'hF7B3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8931 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_573),
    .ADR2(DLX_IDinst_RegFile_5_19),
    .ADR3(DLX_IDinst_RegFile_4_19),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_893)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8941.INIT = 16'hDFD5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8941 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_574),
    .ADR1(DLX_IDinst_RegFile_7_19),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR3(DLX_IDinst_RegFile_6_19),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_894)
  );
  X_BUF \DLX_IDinst_RegFile_5_19/COUTUSED  (
    .I(\DLX_IDinst_RegFile_5_19/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_819)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_819_1256 (
    .IA(\DLX_IDinst_RegFile_5_19/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_818),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_894),
    .O(\DLX_IDinst_RegFile_5_19/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_5_19/CYINIT_1257  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_817),
    .O(\DLX_IDinst_RegFile_5_19/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_5_28/LOGIC_ZERO_1258  (
    .O(\DLX_IDinst_RegFile_5_28/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_450_1259 (
    .IA(\DLX_IDinst_RegFile_5_28/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_5_28/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_509),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_450)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5091.INIT = 16'hFD5D;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5091 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_45),
    .ADR1(DLX_IDinst_RegFile_4_28),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR3(DLX_IDinst_RegFile_5_28),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_509)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5101.INIT = 16'hE4FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5101 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR1(DLX_IDinst_RegFile_6_28),
    .ADR2(DLX_IDinst_RegFile_7_28),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_46),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_510)
  );
  X_BUF \DLX_IDinst_RegFile_5_28/COUTUSED  (
    .I(\DLX_IDinst_RegFile_5_28/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_451)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_451_1260 (
    .IA(\DLX_IDinst_RegFile_5_28/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_450),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_510),
    .O(\DLX_IDinst_RegFile_5_28/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_5_28/CYINIT_1261  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_449),
    .O(\DLX_IDinst_RegFile_5_28/CYINIT )
  );
  defparam DLX_IDinst_RegFile_19_23_1262.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_19_23_1262 (
    .I(DLX_IDinst_WB_data_eff[23]),
    .CE(DLX_IDinst__n0588),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_19_23)
  );
  defparam DLX_IDinst_RegFile_27_14_1263.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_27_14_1263 (
    .I(DLX_IDinst_WB_data_eff[14]),
    .CE(DLX_IDinst__n0604),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_27_14)
  );
  X_ZERO \DLX_IDinst_RegFile_8_10/LOGIC_ZERO_1264  (
    .O(\DLX_IDinst_RegFile_8_10/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_164_1265 (
    .IA(\DLX_IDinst_RegFile_8_10/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_8_10/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_223),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_164)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2231.INIT = 16'hFB3B;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2231 (
    .ADR0(DLX_IDinst_RegFile_8_10),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_47),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR3(DLX_IDinst_RegFile_9_10),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_223)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2241.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2241 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR1(DLX_IDinst_RegFile_10_10),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_48),
    .ADR3(DLX_IDinst_RegFile_11_10),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_224)
  );
  X_BUF \DLX_IDinst_RegFile_8_10/COUTUSED  (
    .I(\DLX_IDinst_RegFile_8_10/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_165)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_165_1266 (
    .IA(\DLX_IDinst_RegFile_8_10/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_164),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_224),
    .O(\DLX_IDinst_RegFile_8_10/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_8_10/CYINIT_1267  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_163),
    .O(\DLX_IDinst_RegFile_8_10/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_8_11/LOGIC_ZERO_1268  (
    .O(\DLX_IDinst_RegFile_8_11/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_180_1269 (
    .IA(\DLX_IDinst_RegFile_8_11/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_8_11/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_239),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_180)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2391.INIT = 16'hDDF5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2391 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_47),
    .ADR1(DLX_IDinst_RegFile_9_11),
    .ADR2(DLX_IDinst_RegFile_8_11),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_239)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2401.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2401 (
    .ADR0(DLX_IDinst_RegFile_10_11),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_48),
    .ADR2(DLX_IDinst_RegFile_11_11),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_240)
  );
  X_BUF \DLX_IDinst_RegFile_8_11/COUTUSED  (
    .I(\DLX_IDinst_RegFile_8_11/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_181)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_181_1270 (
    .IA(\DLX_IDinst_RegFile_8_11/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_180),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_240),
    .O(\DLX_IDinst_RegFile_8_11/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_8_11/CYINIT_1271  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_179),
    .O(\DLX_IDinst_RegFile_8_11/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_8_20/LOGIC_ZERO_1272  (
    .O(\DLX_IDinst_RegFile_8_20/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_324_1273 (
    .IA(\DLX_IDinst_RegFile_8_20/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_8_20/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_383),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_324)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3831.INIT = 16'hF7D5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3831 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_47),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR2(DLX_IDinst_RegFile_9_20),
    .ADR3(DLX_IDinst_RegFile_8_20),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_383)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3841.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3841 (
    .ADR0(DLX_IDinst_RegFile_10_20),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_48),
    .ADR2(DLX_IDinst_RegFile_11_20),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_384)
  );
  X_BUF \DLX_IDinst_RegFile_8_20/COUTUSED  (
    .I(\DLX_IDinst_RegFile_8_20/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_325)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_325_1274 (
    .IA(\DLX_IDinst_RegFile_8_20/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_324),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_384),
    .O(\DLX_IDinst_RegFile_8_20/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_8_20/CYINIT_1275  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_323),
    .O(\DLX_IDinst_RegFile_8_20/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_8_12/LOGIC_ZERO_1276  (
    .O(\DLX_IDinst_RegFile_8_12/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_196_1277 (
    .IA(\DLX_IDinst_RegFile_8_12/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_8_12/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_255),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_196)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2551.INIT = 16'hE4FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2551 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR1(DLX_IDinst_RegFile_8_12),
    .ADR2(DLX_IDinst_RegFile_9_12),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_47),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_255)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2561.INIT = 16'hBF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2561 (
    .ADR0(DLX_IDinst_RegFile_11_12),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_48),
    .ADR3(DLX_IDinst_RegFile_10_12),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_256)
  );
  X_BUF \DLX_IDinst_RegFile_8_12/COUTUSED  (
    .I(\DLX_IDinst_RegFile_8_12/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_197)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_197_1278 (
    .IA(\DLX_IDinst_RegFile_8_12/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_196),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_256),
    .O(\DLX_IDinst_RegFile_8_12/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_8_12/CYINIT_1279  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_195),
    .O(\DLX_IDinst_RegFile_8_12/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_8_21/LOGIC_ZERO_1280  (
    .O(\DLX_IDinst_RegFile_8_21/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_340_1281 (
    .IA(\DLX_IDinst_RegFile_8_21/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_8_21/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_399),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_340)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3991.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3991 (
    .ADR0(DLX_IDinst_RegFile_8_21),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_47),
    .ADR2(DLX_IDinst_RegFile_9_21),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_399)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4001.INIT = 16'hFB3B;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4001 (
    .ADR0(DLX_IDinst_RegFile_10_21),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_48),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR3(DLX_IDinst_RegFile_11_21),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_400)
  );
  X_BUF \DLX_IDinst_RegFile_8_21/COUTUSED  (
    .I(\DLX_IDinst_RegFile_8_21/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_341)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_341_1282 (
    .IA(\DLX_IDinst_RegFile_8_21/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_340),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_400),
    .O(\DLX_IDinst_RegFile_8_21/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_8_21/CYINIT_1283  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_339),
    .O(\DLX_IDinst_RegFile_8_21/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_8_13/LOGIC_ZERO_1284  (
    .O(\DLX_IDinst_RegFile_8_13/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_212_1285 (
    .IA(\DLX_IDinst_RegFile_8_13/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_8_13/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_271),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_212)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2711.INIT = 16'hE2FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2711 (
    .ADR0(DLX_IDinst_RegFile_8_13),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR2(DLX_IDinst_RegFile_9_13),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_47),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_271)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2721.INIT = 16'hBF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2721 (
    .ADR0(DLX_IDinst_RegFile_11_13),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_48),
    .ADR3(DLX_IDinst_RegFile_10_13),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_272)
  );
  X_BUF \DLX_IDinst_RegFile_8_13/COUTUSED  (
    .I(\DLX_IDinst_RegFile_8_13/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_213)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_213_1286 (
    .IA(\DLX_IDinst_RegFile_8_13/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_212),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_272),
    .O(\DLX_IDinst_RegFile_8_13/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_8_13/CYINIT_1287  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_211),
    .O(\DLX_IDinst_RegFile_8_13/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_8_30/LOGIC_ZERO_1288  (
    .O(\DLX_IDinst_RegFile_8_30/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_996_1289 (
    .IA(\DLX_IDinst_RegFile_8_30/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_8_30/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1071),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_996)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10711.INIT = 16'hFD5D;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10711 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_575),
    .ADR1(DLX_IDinst_RegFile_8_30),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR3(DLX_IDinst_RegFile_9_30),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1071)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10721.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10721 (
    .ADR0(DLX_IDinst_RegFile_11_30),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_576),
    .ADR2(DLX_IDinst_RegFile_10_30),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1072)
  );
  X_BUF \DLX_IDinst_RegFile_8_30/COUTUSED  (
    .I(\DLX_IDinst_RegFile_8_30/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_997)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_997_1290 (
    .IA(\DLX_IDinst_RegFile_8_30/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_996),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1072),
    .O(\DLX_IDinst_RegFile_8_30/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_8_30/CYINIT_1291  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_995),
    .O(\DLX_IDinst_RegFile_8_30/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_8_22/LOGIC_ZERO_1292  (
    .O(\DLX_IDinst_RegFile_8_22/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_356_1293 (
    .IA(\DLX_IDinst_RegFile_8_22/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_8_22/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_415),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_356)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4151.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4151 (
    .ADR0(DLX_IDinst_RegFile_8_22),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_47),
    .ADR3(DLX_IDinst_RegFile_9_22),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_415)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4161.INIT = 16'hBFB3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4161 (
    .ADR0(DLX_IDinst_RegFile_11_22),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_48),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR3(DLX_IDinst_RegFile_10_22),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_416)
  );
  X_BUF \DLX_IDinst_RegFile_8_22/COUTUSED  (
    .I(\DLX_IDinst_RegFile_8_22/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_357)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_357_1294 (
    .IA(\DLX_IDinst_RegFile_8_22/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_356),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_416),
    .O(\DLX_IDinst_RegFile_8_22/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_8_22/CYINIT_1295  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_355),
    .O(\DLX_IDinst_RegFile_8_22/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_8_14/LOGIC_ZERO_1296  (
    .O(\DLX_IDinst_RegFile_8_14/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_228_1297 (
    .IA(\DLX_IDinst_RegFile_8_14/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_8_14/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_287),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_228)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2871.INIT = 16'hDFD5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2871 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_47),
    .ADR1(DLX_IDinst_RegFile_9_14),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR3(DLX_IDinst_RegFile_8_14),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_287)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2881.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2881 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_48),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR2(DLX_IDinst_RegFile_10_14),
    .ADR3(DLX_IDinst_RegFile_11_14),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_288)
  );
  X_BUF \DLX_IDinst_RegFile_8_14/COUTUSED  (
    .I(\DLX_IDinst_RegFile_8_14/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_229)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_229_1298 (
    .IA(\DLX_IDinst_RegFile_8_14/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_228),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_288),
    .O(\DLX_IDinst_RegFile_8_14/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_8_14/CYINIT_1299  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_227),
    .O(\DLX_IDinst_RegFile_8_14/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_8_23/LOGIC_ZERO_1300  (
    .O(\DLX_IDinst_RegFile_8_23/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_372_1301 (
    .IA(\DLX_IDinst_RegFile_8_23/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_8_23/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_431),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_372)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4311.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4311 (
    .ADR0(DLX_IDinst_RegFile_8_23),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_47),
    .ADR2(DLX_IDinst_RegFile_9_23),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_431)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4321.INIT = 16'hDDF5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4321 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_48),
    .ADR1(DLX_IDinst_RegFile_11_23),
    .ADR2(DLX_IDinst_RegFile_10_23),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_432)
  );
  X_BUF \DLX_IDinst_RegFile_8_23/COUTUSED  (
    .I(\DLX_IDinst_RegFile_8_23/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_373)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_373_1302 (
    .IA(\DLX_IDinst_RegFile_8_23/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_372),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_432),
    .O(\DLX_IDinst_RegFile_8_23/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_8_23/CYINIT_1303  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_371),
    .O(\DLX_IDinst_RegFile_8_23/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_8_15/LOGIC_ZERO_1304  (
    .O(\DLX_IDinst_RegFile_8_15/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_244_1305 (
    .IA(\DLX_IDinst_RegFile_8_15/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_8_15/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_303),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_244)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3031.INIT = 16'hAFCF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3031 (
    .ADR0(DLX_IDinst_RegFile_9_15),
    .ADR1(DLX_IDinst_RegFile_8_15),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_47),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_303)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3041.INIT = 16'hACFF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3041 (
    .ADR0(DLX_IDinst_RegFile_11_15),
    .ADR1(DLX_IDinst_RegFile_10_15),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_48),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_304)
  );
  X_BUF \DLX_IDinst_RegFile_8_15/COUTUSED  (
    .I(\DLX_IDinst_RegFile_8_15/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_245)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_245_1306 (
    .IA(\DLX_IDinst_RegFile_8_15/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_244),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_304),
    .O(\DLX_IDinst_RegFile_8_15/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_8_15/CYINIT_1307  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_243),
    .O(\DLX_IDinst_RegFile_8_15/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_8_31/LOGIC_ZERO_1308  (
    .O(\DLX_IDinst_RegFile_8_31/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_1012_1309 (
    .IA(\DLX_IDinst_RegFile_8_31/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_8_31/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1087),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_1012)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10871.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10871 (
    .ADR0(DLX_IDinst_RegFile_9_31),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_575),
    .ADR2(DLX_IDinst_RegFile_8_31),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1087)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10881.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10881 (
    .ADR0(DLX_IDinst_RegFile_10_31),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_576),
    .ADR2(DLX_IDinst_RegFile_11_31),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1088)
  );
  X_BUF \DLX_IDinst_RegFile_8_31/COUTUSED  (
    .I(\DLX_IDinst_RegFile_8_31/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_1013)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_1013_1310 (
    .IA(\DLX_IDinst_RegFile_8_31/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_1012),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1088),
    .O(\DLX_IDinst_RegFile_8_31/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_8_31/CYINIT_1311  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_1011),
    .O(\DLX_IDinst_RegFile_8_31/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_8_24/LOGIC_ZERO_1312  (
    .O(\DLX_IDinst_RegFile_8_24/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_388_1313 (
    .IA(\DLX_IDinst_RegFile_8_24/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_8_24/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_447),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_388)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4471.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4471 (
    .ADR0(DLX_IDinst_RegFile_8_24),
    .ADR1(DLX_IDinst_RegFile_9_24),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_47),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_447)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4481.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4481 (
    .ADR0(DLX_IDinst_RegFile_10_24),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_48),
    .ADR2(DLX_IDinst_RegFile_11_24),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_448)
  );
  X_BUF \DLX_IDinst_RegFile_8_24/COUTUSED  (
    .I(\DLX_IDinst_RegFile_8_24/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_389)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_389_1314 (
    .IA(\DLX_IDinst_RegFile_8_24/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_388),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_448),
    .O(\DLX_IDinst_RegFile_8_24/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_8_24/CYINIT_1315  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_387),
    .O(\DLX_IDinst_RegFile_8_24/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_8_16/LOGIC_ZERO_1316  (
    .O(\DLX_IDinst_RegFile_8_16/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_260_1317 (
    .IA(\DLX_IDinst_RegFile_8_16/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_8_16/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_319),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_260)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3191.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3191 (
    .ADR0(DLX_IDinst_RegFile_8_16),
    .ADR1(DLX_IDinst_RegFile_9_16),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_47),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_319)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3201.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3201 (
    .ADR0(DLX_IDinst_RegFile_10_16),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_48),
    .ADR2(DLX_IDinst_RegFile_11_16),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_320)
  );
  X_BUF \DLX_IDinst_RegFile_8_16/COUTUSED  (
    .I(\DLX_IDinst_RegFile_8_16/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_261)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_261_1318 (
    .IA(\DLX_IDinst_RegFile_8_16/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_260),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_320),
    .O(\DLX_IDinst_RegFile_8_16/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_8_16/CYINIT_1319  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_259),
    .O(\DLX_IDinst_RegFile_8_16/CYINIT )
  );
  defparam DLX_IDinst_RegFile_19_15_1320.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_19_15_1320 (
    .I(DLX_IDinst_WB_data_eff[15]),
    .CE(DLX_IDinst__n0588),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_19_15)
  );
  X_ZERO \DLX_IDinst_RegFile_8_25/LOGIC_ZERO_1321  (
    .O(\DLX_IDinst_RegFile_8_25/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_404_1322 (
    .IA(\DLX_IDinst_RegFile_8_25/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_8_25/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_463),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_404)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4631.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4631 (
    .ADR0(DLX_IDinst_RegFile_8_25),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_47),
    .ADR2(DLX_IDinst_RegFile_9_25),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_463)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4641.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4641 (
    .ADR0(DLX_IDinst_RegFile_10_25),
    .ADR1(DLX_IDinst_RegFile_11_25),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_48),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_464)
  );
  X_BUF \DLX_IDinst_RegFile_8_25/COUTUSED  (
    .I(\DLX_IDinst_RegFile_8_25/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_405)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_405_1323 (
    .IA(\DLX_IDinst_RegFile_8_25/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_404),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_464),
    .O(\DLX_IDinst_RegFile_8_25/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_8_25/CYINIT_1324  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_403),
    .O(\DLX_IDinst_RegFile_8_25/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_8_17/LOGIC_ZERO_1325  (
    .O(\DLX_IDinst_RegFile_8_17/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_276_1326 (
    .IA(\DLX_IDinst_RegFile_8_17/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_8_17/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_335),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_276)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3351.INIT = 16'hB8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3351 (
    .ADR0(DLX_IDinst_RegFile_9_17),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR2(DLX_IDinst_RegFile_8_17),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_47),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_335)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3361.INIT = 16'hBFB3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3361 (
    .ADR0(DLX_IDinst_RegFile_11_17),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_48),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR3(DLX_IDinst_RegFile_10_17),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_336)
  );
  X_BUF \DLX_IDinst_RegFile_8_17/COUTUSED  (
    .I(\DLX_IDinst_RegFile_8_17/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_277)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_277_1327 (
    .IA(\DLX_IDinst_RegFile_8_17/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_276),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_336),
    .O(\DLX_IDinst_RegFile_8_17/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_8_17/CYINIT_1328  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_275),
    .O(\DLX_IDinst_RegFile_8_17/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_8_26/LOGIC_ZERO_1329  (
    .O(\DLX_IDinst_RegFile_8_26/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_420_1330 (
    .IA(\DLX_IDinst_RegFile_8_26/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_8_26/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_479),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_420)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4791.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4791 (
    .ADR0(DLX_IDinst_RegFile_8_26),
    .ADR1(DLX_IDinst_RegFile_9_26),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_47),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_479)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4801.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4801 (
    .ADR0(DLX_IDinst_RegFile_10_26),
    .ADR1(DLX_IDinst_RegFile_11_26),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_48),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_480)
  );
  X_BUF \DLX_IDinst_RegFile_8_26/COUTUSED  (
    .I(\DLX_IDinst_RegFile_8_26/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_421)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_421_1331 (
    .IA(\DLX_IDinst_RegFile_8_26/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_420),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_480),
    .O(\DLX_IDinst_RegFile_8_26/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_8_26/CYINIT_1332  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_419),
    .O(\DLX_IDinst_RegFile_8_26/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_8_18/LOGIC_ZERO_1333  (
    .O(\DLX_IDinst_RegFile_8_18/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_292_1334 (
    .IA(\DLX_IDinst_RegFile_8_18/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_8_18/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_351),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_292)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3511.INIT = 16'hDFD5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3511 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_47),
    .ADR1(DLX_IDinst_RegFile_9_18),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR3(DLX_IDinst_RegFile_8_18),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_351)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3521.INIT = 16'hCFAF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3521 (
    .ADR0(DLX_IDinst_RegFile_10_18),
    .ADR1(DLX_IDinst_RegFile_11_18),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_48),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_352)
  );
  X_BUF \DLX_IDinst_RegFile_8_18/COUTUSED  (
    .I(\DLX_IDinst_RegFile_8_18/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_293)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_293_1335 (
    .IA(\DLX_IDinst_RegFile_8_18/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_292),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_352),
    .O(\DLX_IDinst_RegFile_8_18/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_8_18/CYINIT_1336  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_291),
    .O(\DLX_IDinst_RegFile_8_18/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_9_10/LOGIC_ZERO_1337  (
    .O(\DLX_IDinst_RegFile_9_10/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_676_1338 (
    .IA(\DLX_IDinst_RegFile_9_10/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_9_10/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_751),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_676)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7511.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7511 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_575),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR2(DLX_IDinst_RegFile_8_10),
    .ADR3(DLX_IDinst_RegFile_9_10),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_751)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7521.INIT = 16'hCFAF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7521 (
    .ADR0(DLX_IDinst_RegFile_10_10),
    .ADR1(DLX_IDinst_RegFile_11_10),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_576),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_752)
  );
  X_BUF \DLX_IDinst_RegFile_9_10/COUTUSED  (
    .I(\DLX_IDinst_RegFile_9_10/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_677)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_677_1339 (
    .IA(\DLX_IDinst_RegFile_9_10/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_676),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_752),
    .O(\DLX_IDinst_RegFile_9_10/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_9_10/CYINIT_1340  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_675),
    .O(\DLX_IDinst_RegFile_9_10/CYINIT )
  );
  defparam \DLX_EXinst__n0007<4>216_SW0 .INIT = 16'h1400;
  X_LUT4 \DLX_EXinst__n0007<4>216_SW0  (
    .ADR0(DLX_IDinst_IR_opcode_field[0]),
    .ADR1(DLX_IDinst_reg_out_A[4]),
    .ADR2(DLX_IDinst_IR_opcode_field[1]),
    .ADR3(DLX_EXinst_N76011),
    .O(\N163827/FROM )
  );
  defparam \DLX_EXinst__n0007<4>216 .INIT = 16'hFFF8;
  X_LUT4 \DLX_EXinst__n0007<4>216  (
    .ADR0(\DLX_EXinst_Mshift__n0022_Sh[52] ),
    .ADR1(DLX_EXinst_N76441),
    .ADR2(CHOICE4371),
    .ADR3(N163827),
    .O(\N163827/GROM )
  );
  X_BUF \N163827/XUSED  (
    .I(\N163827/FROM ),
    .O(N163827)
  );
  X_BUF \N163827/YUSED  (
    .I(\N163827/GROM ),
    .O(CHOICE4373)
  );
  defparam DLX_IDinst_RegFile_19_31_1341.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_19_31_1341 (
    .I(DLX_IDinst_WB_data_eff[31]),
    .CE(DLX_IDinst__n0588),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_19_31)
  );
  X_ZERO \DLX_IDinst_RegFile_8_27/LOGIC_ZERO_1342  (
    .O(\DLX_IDinst_RegFile_8_27/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_436_1343 (
    .IA(\DLX_IDinst_RegFile_8_27/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_8_27/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_495),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_436)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4951.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4951 (
    .ADR0(DLX_IDinst_RegFile_8_27),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_47),
    .ADR3(DLX_IDinst_RegFile_9_27),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_495)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4961.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4961 (
    .ADR0(DLX_IDinst_RegFile_10_27),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_48),
    .ADR3(DLX_IDinst_RegFile_11_27),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_496)
  );
  X_BUF \DLX_IDinst_RegFile_8_27/COUTUSED  (
    .I(\DLX_IDinst_RegFile_8_27/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_437)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_437_1344 (
    .IA(\DLX_IDinst_RegFile_8_27/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_436),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_496),
    .O(\DLX_IDinst_RegFile_8_27/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_8_27/CYINIT_1345  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_435),
    .O(\DLX_IDinst_RegFile_8_27/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_8_19/LOGIC_ZERO_1346  (
    .O(\DLX_IDinst_RegFile_8_19/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_308_1347 (
    .IA(\DLX_IDinst_RegFile_8_19/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_8_19/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_367),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_308)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3671.INIT = 16'hE4FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3671 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR1(DLX_IDinst_RegFile_8_19),
    .ADR2(DLX_IDinst_RegFile_9_19),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_47),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_367)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3681.INIT = 16'hDF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3681 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR1(DLX_IDinst_RegFile_11_19),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_48),
    .ADR3(DLX_IDinst_RegFile_10_19),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_368)
  );
  X_BUF \DLX_IDinst_RegFile_8_19/COUTUSED  (
    .I(\DLX_IDinst_RegFile_8_19/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_309)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_309_1348 (
    .IA(\DLX_IDinst_RegFile_8_19/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_308),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_368),
    .O(\DLX_IDinst_RegFile_8_19/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_8_19/CYINIT_1349  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_307),
    .O(\DLX_IDinst_RegFile_8_19/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_9_11/LOGIC_ZERO_1350  (
    .O(\DLX_IDinst_RegFile_9_11/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_692_1351 (
    .IA(\DLX_IDinst_RegFile_9_11/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_9_11/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_767),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_692)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7671.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7671 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR1(DLX_IDinst_RegFile_8_11),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_575),
    .ADR3(DLX_IDinst_RegFile_9_11),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_767)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7681.INIT = 16'hDDF5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7681 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_576),
    .ADR1(DLX_IDinst_RegFile_11_11),
    .ADR2(DLX_IDinst_RegFile_10_11),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_768)
  );
  X_BUF \DLX_IDinst_RegFile_9_11/COUTUSED  (
    .I(\DLX_IDinst_RegFile_9_11/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_693)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_693_1352 (
    .IA(\DLX_IDinst_RegFile_9_11/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_692),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_768),
    .O(\DLX_IDinst_RegFile_9_11/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_9_11/CYINIT_1353  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_691),
    .O(\DLX_IDinst_RegFile_9_11/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_8_28/LOGIC_ZERO_1354  (
    .O(\DLX_IDinst_RegFile_8_28/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_964_1355 (
    .IA(\DLX_IDinst_RegFile_8_28/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_8_28/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1039),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_964)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10391.INIT = 16'hFB3B;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10391 (
    .ADR0(DLX_IDinst_RegFile_8_28),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_575),
    .ADR2(DLX_IDinst_jtarget[21]),
    .ADR3(DLX_IDinst_RegFile_9_28),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1039)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10401.INIT = 16'hF7D5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10401 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_576),
    .ADR1(DLX_IDinst_jtarget[21]),
    .ADR2(DLX_IDinst_RegFile_11_28),
    .ADR3(DLX_IDinst_RegFile_10_28),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1040)
  );
  X_BUF \DLX_IDinst_RegFile_8_28/COUTUSED  (
    .I(\DLX_IDinst_RegFile_8_28/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_965)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_965_1356 (
    .IA(\DLX_IDinst_RegFile_8_28/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_964),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1040),
    .O(\DLX_IDinst_RegFile_8_28/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_8_28/CYINIT_1357  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_963),
    .O(\DLX_IDinst_RegFile_8_28/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_9_20/LOGIC_ZERO_1358  (
    .O(\DLX_IDinst_RegFile_9_20/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_836_1359 (
    .IA(\DLX_IDinst_RegFile_9_20/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_9_20/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_911),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_836)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9111.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9111 (
    .ADR0(DLX_IDinst_RegFile_9_20),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_575),
    .ADR2(DLX_IDinst_RegFile_8_20),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_911)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9121.INIT = 16'hD8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9121 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR1(DLX_IDinst_RegFile_11_20),
    .ADR2(DLX_IDinst_RegFile_10_20),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_576),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_912)
  );
  X_BUF \DLX_IDinst_RegFile_9_20/COUTUSED  (
    .I(\DLX_IDinst_RegFile_9_20/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_837)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_837_1360 (
    .IA(\DLX_IDinst_RegFile_9_20/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_836),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_912),
    .O(\DLX_IDinst_RegFile_9_20/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_9_20/CYINIT_1361  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_835),
    .O(\DLX_IDinst_RegFile_9_20/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_9_12/LOGIC_ZERO_1362  (
    .O(\DLX_IDinst_RegFile_9_12/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_708_1363 (
    .IA(\DLX_IDinst_RegFile_9_12/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_9_12/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_783),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_708)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7831.INIT = 16'hD8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7831 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR1(DLX_IDinst_RegFile_9_12),
    .ADR2(DLX_IDinst_RegFile_8_12),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_575),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_783)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7841.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7841 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR1(DLX_IDinst_RegFile_10_12),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_576),
    .ADR3(DLX_IDinst_RegFile_11_12),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_784)
  );
  X_BUF \DLX_IDinst_RegFile_9_12/COUTUSED  (
    .I(\DLX_IDinst_RegFile_9_12/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_709)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_709_1364 (
    .IA(\DLX_IDinst_RegFile_9_12/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_708),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_784),
    .O(\DLX_IDinst_RegFile_9_12/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_9_12/CYINIT_1365  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_707),
    .O(\DLX_IDinst_RegFile_9_12/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_8_29/LOGIC_ZERO_1366  (
    .O(\DLX_IDinst_RegFile_8_29/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_980_1367 (
    .IA(\DLX_IDinst_RegFile_8_29/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_8_29/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1055),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_980)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10551.INIT = 16'hF7D5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10551 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_575),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR2(DLX_IDinst_RegFile_9_29),
    .ADR3(DLX_IDinst_RegFile_8_29),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1055)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10561.INIT = 16'hAFCF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10561 (
    .ADR0(DLX_IDinst_RegFile_11_29),
    .ADR1(DLX_IDinst_RegFile_10_29),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_576),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1056)
  );
  X_BUF \DLX_IDinst_RegFile_8_29/COUTUSED  (
    .I(\DLX_IDinst_RegFile_8_29/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_981)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_981_1368 (
    .IA(\DLX_IDinst_RegFile_8_29/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_980),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1056),
    .O(\DLX_IDinst_RegFile_8_29/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_8_29/CYINIT_1369  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_979),
    .O(\DLX_IDinst_RegFile_8_29/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_9_21/LOGIC_ZERO_1370  (
    .O(\DLX_IDinst_RegFile_9_21/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_852_1371 (
    .IA(\DLX_IDinst_RegFile_9_21/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_9_21/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_927),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_852)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9271.INIT = 16'hFB73;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9271 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_575),
    .ADR2(DLX_IDinst_RegFile_8_21),
    .ADR3(DLX_IDinst_RegFile_9_21),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_927)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9281.INIT = 16'hACFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9281 (
    .ADR0(DLX_IDinst_RegFile_11_21),
    .ADR1(DLX_IDinst_RegFile_10_21),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_576),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_928)
  );
  X_BUF \DLX_IDinst_RegFile_9_21/COUTUSED  (
    .I(\DLX_IDinst_RegFile_9_21/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_853)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_853_1372 (
    .IA(\DLX_IDinst_RegFile_9_21/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_852),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_928),
    .O(\DLX_IDinst_RegFile_9_21/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_9_21/CYINIT_1373  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_851),
    .O(\DLX_IDinst_RegFile_9_21/CYINIT )
  );
  defparam DLX_IDinst_RegFile_27_15_1374.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_27_15_1374 (
    .I(DLX_IDinst_WB_data_eff[15]),
    .CE(DLX_IDinst__n0604),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_27_15)
  );
  X_ZERO \DLX_IDinst_RegFile_9_13/LOGIC_ZERO_1375  (
    .O(\DLX_IDinst_RegFile_9_13/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_724_1376 (
    .IA(\DLX_IDinst_RegFile_9_13/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_9_13/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_799),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_724)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7991.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7991 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR1(DLX_IDinst_RegFile_8_13),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_575),
    .ADR3(DLX_IDinst_RegFile_9_13),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_799)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8001.INIT = 16'hDFD5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8001 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_576),
    .ADR1(DLX_IDinst_RegFile_11_13),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR3(DLX_IDinst_RegFile_10_13),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_800)
  );
  X_BUF \DLX_IDinst_RegFile_9_13/COUTUSED  (
    .I(\DLX_IDinst_RegFile_9_13/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_725)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_725_1377 (
    .IA(\DLX_IDinst_RegFile_9_13/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_724),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_800),
    .O(\DLX_IDinst_RegFile_9_13/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_9_13/CYINIT_1378  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_723),
    .O(\DLX_IDinst_RegFile_9_13/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_9_30/LOGIC_ZERO_1379  (
    .O(\DLX_IDinst_RegFile_9_30/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_484_1380 (
    .IA(\DLX_IDinst_RegFile_9_30/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_9_30/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_543),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_484)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5431.INIT = 16'hCFAF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5431 (
    .ADR0(DLX_IDinst_RegFile_8_30),
    .ADR1(DLX_IDinst_RegFile_9_30),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_47),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_543)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5441.INIT = 16'hDF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5441 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR1(DLX_IDinst_RegFile_11_30),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_48),
    .ADR3(DLX_IDinst_RegFile_10_30),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_544)
  );
  X_BUF \DLX_IDinst_RegFile_9_30/COUTUSED  (
    .I(\DLX_IDinst_RegFile_9_30/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_485)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_485_1381 (
    .IA(\DLX_IDinst_RegFile_9_30/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_484),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_544),
    .O(\DLX_IDinst_RegFile_9_30/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_9_30/CYINIT_1382  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_483),
    .O(\DLX_IDinst_RegFile_9_30/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_9_22/LOGIC_ZERO_1383  (
    .O(\DLX_IDinst_RegFile_9_22/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_868_1384 (
    .IA(\DLX_IDinst_RegFile_9_22/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_9_22/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_943),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_868)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9431.INIT = 16'hFB73;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9431 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_575),
    .ADR2(DLX_IDinst_RegFile_8_22),
    .ADR3(DLX_IDinst_RegFile_9_22),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_943)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9441.INIT = 16'hACFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9441 (
    .ADR0(DLX_IDinst_RegFile_11_22),
    .ADR1(DLX_IDinst_RegFile_10_22),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_576),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_944)
  );
  X_BUF \DLX_IDinst_RegFile_9_22/COUTUSED  (
    .I(\DLX_IDinst_RegFile_9_22/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_869)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_869_1385 (
    .IA(\DLX_IDinst_RegFile_9_22/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_868),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_944),
    .O(\DLX_IDinst_RegFile_9_22/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_9_22/CYINIT_1386  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_867),
    .O(\DLX_IDinst_RegFile_9_22/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_9_23/LOGIC_ZERO_1387  (
    .O(\DLX_IDinst_RegFile_9_23/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_884_1388 (
    .IA(\DLX_IDinst_RegFile_9_23/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_9_23/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_959),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_884)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9591.INIT = 16'hE2FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9591 (
    .ADR0(DLX_IDinst_RegFile_8_23),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR2(DLX_IDinst_RegFile_9_23),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_575),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_959)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9601.INIT = 16'hACFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9601 (
    .ADR0(DLX_IDinst_RegFile_11_23),
    .ADR1(DLX_IDinst_RegFile_10_23),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_576),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_960)
  );
  X_BUF \DLX_IDinst_RegFile_9_23/COUTUSED  (
    .I(\DLX_IDinst_RegFile_9_23/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_885)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_885_1389 (
    .IA(\DLX_IDinst_RegFile_9_23/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_884),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_960),
    .O(\DLX_IDinst_RegFile_9_23/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_9_23/CYINIT_1390  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_883),
    .O(\DLX_IDinst_RegFile_9_23/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_9_15/LOGIC_ZERO_1391  (
    .O(\DLX_IDinst_RegFile_9_15/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_756_1392 (
    .IA(\DLX_IDinst_RegFile_9_15/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_9_15/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_831),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_756)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8311.INIT = 16'hAFCF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8311 (
    .ADR0(DLX_IDinst_RegFile_9_15),
    .ADR1(DLX_IDinst_RegFile_8_15),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_575),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_831)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8321.INIT = 16'hAFCF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8321 (
    .ADR0(DLX_IDinst_RegFile_11_15),
    .ADR1(DLX_IDinst_RegFile_10_15),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_576),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_832)
  );
  X_BUF \DLX_IDinst_RegFile_9_15/COUTUSED  (
    .I(\DLX_IDinst_RegFile_9_15/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_757)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_757_1393 (
    .IA(\DLX_IDinst_RegFile_9_15/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_756),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_832),
    .O(\DLX_IDinst_RegFile_9_15/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_9_15/CYINIT_1394  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_755),
    .O(\DLX_IDinst_RegFile_9_15/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_9_31/LOGIC_ZERO_1395  (
    .O(\DLX_IDinst_RegFile_9_31/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_500_1396 (
    .IA(\DLX_IDinst_RegFile_9_31/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_9_31/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_559),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_500)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5591.INIT = 16'hDFD5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5591 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_47),
    .ADR1(DLX_IDinst_RegFile_9_31),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR3(DLX_IDinst_RegFile_8_31),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_559)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5601.INIT = 16'hD8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5601 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR1(DLX_IDinst_RegFile_11_31),
    .ADR2(DLX_IDinst_RegFile_10_31),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_48),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_560)
  );
  X_BUF \DLX_IDinst_RegFile_9_31/COUTUSED  (
    .I(\DLX_IDinst_RegFile_9_31/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_501)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_501_1397 (
    .IA(\DLX_IDinst_RegFile_9_31/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_500),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_560),
    .O(\DLX_IDinst_RegFile_9_31/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_9_31/CYINIT_1398  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_499),
    .O(\DLX_IDinst_RegFile_9_31/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_9_24/LOGIC_ZERO_1399  (
    .O(\DLX_IDinst_RegFile_9_24/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_900_1400 (
    .IA(\DLX_IDinst_RegFile_9_24/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_9_24/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_975),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_900)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9751.INIT = 16'hE2FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9751 (
    .ADR0(DLX_IDinst_RegFile_8_24),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR2(DLX_IDinst_RegFile_9_24),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_575),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_975)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9761.INIT = 16'hACFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9761 (
    .ADR0(DLX_IDinst_RegFile_11_24),
    .ADR1(DLX_IDinst_RegFile_10_24),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_576),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_976)
  );
  X_BUF \DLX_IDinst_RegFile_9_24/COUTUSED  (
    .I(\DLX_IDinst_RegFile_9_24/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_901)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_901_1401 (
    .IA(\DLX_IDinst_RegFile_9_24/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_900),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_976),
    .O(\DLX_IDinst_RegFile_9_24/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_9_24/CYINIT_1402  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_899),
    .O(\DLX_IDinst_RegFile_9_24/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_9_16/LOGIC_ZERO_1403  (
    .O(\DLX_IDinst_RegFile_9_16/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_772_1404 (
    .IA(\DLX_IDinst_RegFile_9_16/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_9_16/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_847),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_772)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8471.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8471 (
    .ADR0(DLX_IDinst_RegFile_9_16),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_575),
    .ADR2(DLX_IDinst_RegFile_8_16),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_847)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8481.INIT = 16'hF7B3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8481 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_576),
    .ADR2(DLX_IDinst_RegFile_11_16),
    .ADR3(DLX_IDinst_RegFile_10_16),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_848)
  );
  X_BUF \DLX_IDinst_RegFile_9_16/COUTUSED  (
    .I(\DLX_IDinst_RegFile_9_16/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_773)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_773_1405 (
    .IA(\DLX_IDinst_RegFile_9_16/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_772),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_848),
    .O(\DLX_IDinst_RegFile_9_16/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_9_16/CYINIT_1406  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_771),
    .O(\DLX_IDinst_RegFile_9_16/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_9_25/LOGIC_ZERO_1407  (
    .O(\DLX_IDinst_RegFile_9_25/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_916_1408 (
    .IA(\DLX_IDinst_RegFile_9_25/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_9_25/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_991),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_916)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9911.INIT = 16'hDFD5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9911 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_575),
    .ADR1(DLX_IDinst_RegFile_9_25),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR3(DLX_IDinst_RegFile_8_25),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_991)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9921.INIT = 16'hB8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9921 (
    .ADR0(DLX_IDinst_RegFile_11_25),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR2(DLX_IDinst_RegFile_10_25),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_576),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_992)
  );
  X_BUF \DLX_IDinst_RegFile_9_25/COUTUSED  (
    .I(\DLX_IDinst_RegFile_9_25/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_917)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_917_1409 (
    .IA(\DLX_IDinst_RegFile_9_25/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_916),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_992),
    .O(\DLX_IDinst_RegFile_9_25/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_9_25/CYINIT_1410  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_915),
    .O(\DLX_IDinst_RegFile_9_25/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_9_17/LOGIC_ZERO_1411  (
    .O(\DLX_IDinst_RegFile_9_17/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_788_1412 (
    .IA(\DLX_IDinst_RegFile_9_17/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_9_17/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_863),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_788)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8631.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8631 (
    .ADR0(DLX_IDinst_RegFile_8_17),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_575),
    .ADR3(DLX_IDinst_RegFile_9_17),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_863)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8641.INIT = 16'hF7B3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8641 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_576),
    .ADR2(DLX_IDinst_RegFile_11_17),
    .ADR3(DLX_IDinst_RegFile_10_17),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_864)
  );
  X_BUF \DLX_IDinst_RegFile_9_17/COUTUSED  (
    .I(\DLX_IDinst_RegFile_9_17/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_789)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_789_1413 (
    .IA(\DLX_IDinst_RegFile_9_17/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_788),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_864),
    .O(\DLX_IDinst_RegFile_9_17/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_9_17/CYINIT_1414  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_787),
    .O(\DLX_IDinst_RegFile_9_17/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_9_26/LOGIC_ZERO_1415  (
    .O(\DLX_IDinst_RegFile_9_26/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_932_1416 (
    .IA(\DLX_IDinst_RegFile_9_26/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_9_26/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1007),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_932)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10071.INIT = 16'hACFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10071 (
    .ADR0(DLX_IDinst_RegFile_9_26),
    .ADR1(DLX_IDinst_RegFile_8_26),
    .ADR2(DLX_IDinst_jtarget[21]),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_575),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1007)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10081.INIT = 16'hE4FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10081 (
    .ADR0(DLX_IDinst_jtarget[21]),
    .ADR1(DLX_IDinst_RegFile_10_26),
    .ADR2(DLX_IDinst_RegFile_11_26),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_576),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1008)
  );
  X_BUF \DLX_IDinst_RegFile_9_26/COUTUSED  (
    .I(\DLX_IDinst_RegFile_9_26/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_933)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_933_1417 (
    .IA(\DLX_IDinst_RegFile_9_26/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_932),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1008),
    .O(\DLX_IDinst_RegFile_9_26/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_9_26/CYINIT_1418  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_931),
    .O(\DLX_IDinst_RegFile_9_26/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_9_18/LOGIC_ZERO_1419  (
    .O(\DLX_IDinst_RegFile_9_18/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_804_1420 (
    .IA(\DLX_IDinst_RegFile_9_18/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_9_18/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_879),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_804)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8791.INIT = 16'hAFCF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8791 (
    .ADR0(DLX_IDinst_RegFile_9_18),
    .ADR1(DLX_IDinst_RegFile_8_18),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_575),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_879)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8801.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8801 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR1(DLX_IDinst_RegFile_10_18),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_576),
    .ADR3(DLX_IDinst_RegFile_11_18),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_880)
  );
  X_BUF \DLX_IDinst_RegFile_9_18/COUTUSED  (
    .I(\DLX_IDinst_RegFile_9_18/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_805)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_805_1421 (
    .IA(\DLX_IDinst_RegFile_9_18/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_804),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_880),
    .O(\DLX_IDinst_RegFile_9_18/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_9_18/CYINIT_1422  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_803),
    .O(\DLX_IDinst_RegFile_9_18/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_9_27/LOGIC_ZERO_1423  (
    .O(\DLX_IDinst_RegFile_9_27/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_948_1424 (
    .IA(\DLX_IDinst_RegFile_9_27/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_9_27/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1023),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_948)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10231.INIT = 16'hDF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10231 (
    .ADR0(DLX_IDinst_jtarget[21]),
    .ADR1(DLX_IDinst_RegFile_9_27),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_575),
    .ADR3(DLX_IDinst_RegFile_8_27),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1023)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10241.INIT = 16'hBFB3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10241 (
    .ADR0(DLX_IDinst_RegFile_11_27),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_576),
    .ADR2(DLX_IDinst_jtarget[21]),
    .ADR3(DLX_IDinst_RegFile_10_27),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1024)
  );
  X_BUF \DLX_IDinst_RegFile_9_27/COUTUSED  (
    .I(\DLX_IDinst_RegFile_9_27/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_949)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_949_1425 (
    .IA(\DLX_IDinst_RegFile_9_27/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_948),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1024),
    .O(\DLX_IDinst_RegFile_9_27/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_9_27/CYINIT_1426  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_947),
    .O(\DLX_IDinst_RegFile_9_27/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_9_19/LOGIC_ZERO_1427  (
    .O(\DLX_IDinst_RegFile_9_19/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_820_1428 (
    .IA(\DLX_IDinst_RegFile_9_19/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_9_19/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_895),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_820)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8951.INIT = 16'hFB3B;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8951 (
    .ADR0(DLX_IDinst_RegFile_8_19),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_575),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR3(DLX_IDinst_RegFile_9_19),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_895)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8961.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8961 (
    .ADR0(DLX_IDinst_RegFile_10_19),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_576),
    .ADR2(DLX_IDinst_RegFile_11_19),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_896)
  );
  X_BUF \DLX_IDinst_RegFile_9_19/COUTUSED  (
    .I(\DLX_IDinst_RegFile_9_19/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_821)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_821_1429 (
    .IA(\DLX_IDinst_RegFile_9_19/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_820),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_896),
    .O(\DLX_IDinst_RegFile_9_19/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_9_19/CYINIT_1430  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_819),
    .O(\DLX_IDinst_RegFile_9_19/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_9_28/LOGIC_ZERO_1431  (
    .O(\DLX_IDinst_RegFile_9_28/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_452_1432 (
    .IA(\DLX_IDinst_RegFile_9_28/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_9_28/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_511),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_452)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5111.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5111 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_47),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR2(DLX_IDinst_RegFile_8_28),
    .ADR3(DLX_IDinst_RegFile_9_28),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_511)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5121.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5121 (
    .ADR0(DLX_IDinst_RegFile_11_28),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_48),
    .ADR2(DLX_IDinst_RegFile_10_28),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_512)
  );
  X_BUF \DLX_IDinst_RegFile_9_28/COUTUSED  (
    .I(\DLX_IDinst_RegFile_9_28/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_453)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_453_1433 (
    .IA(\DLX_IDinst_RegFile_9_28/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_452),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_512),
    .O(\DLX_IDinst_RegFile_9_28/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_9_28/CYINIT_1434  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_451),
    .O(\DLX_IDinst_RegFile_9_28/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_9_29/LOGIC_ZERO_1435  (
    .O(\DLX_IDinst_RegFile_9_29/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_468_1436 (
    .IA(\DLX_IDinst_RegFile_9_29/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_9_29/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_527),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_468)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5271.INIT = 16'hF7D5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5271 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_47),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR2(DLX_IDinst_RegFile_9_29),
    .ADR3(DLX_IDinst_RegFile_8_29),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_527)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5281.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5281 (
    .ADR0(DLX_IDinst_RegFile_10_29),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_48),
    .ADR2(DLX_IDinst_RegFile_11_29),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_528)
  );
  X_BUF \DLX_IDinst_RegFile_9_29/COUTUSED  (
    .I(\DLX_IDinst_RegFile_9_29/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_469)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_469_1437 (
    .IA(\DLX_IDinst_RegFile_9_29/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_468),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_528),
    .O(\DLX_IDinst_RegFile_9_29/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_9_29/CYINIT_1438  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_467),
    .O(\DLX_IDinst_RegFile_9_29/CYINIT )
  );
  defparam vga_top_vga1_Ker112924_SW0.INIT = 16'hFFFE;
  X_LUT4 vga_top_vga1_Ker112924_SW0 (
    .ADR0(vga_top_vga1_hcounter[13]),
    .ADR1(vga_top_vga1_hcounter[10]),
    .ADR2(vga_top_vga1_hcounter[11]),
    .ADR3(vga_top_vga1_hcounter[12]),
    .O(\N136625/FROM )
  );
  defparam vga_top_vga1_Ker112924.INIT = 16'h0001;
  X_LUT4 vga_top_vga1_Ker112924 (
    .ADR0(vga_top_vga1_hcounter[15]),
    .ADR1(vga_top_vga1_hcounter[14]),
    .ADR2(vga_top_vga1_hcounter[6]),
    .ADR3(N136625),
    .O(\N136625/GROM )
  );
  X_BUF \N136625/XUSED  (
    .I(\N136625/FROM ),
    .O(N136625)
  );
  X_BUF \N136625/YUSED  (
    .I(\N136625/GROM ),
    .O(vga_top_vga1_N112926)
  );
  defparam DLX_IDinst__n01611.INIT = 16'h0100;
  X_LUT4 DLX_IDinst__n01611 (
    .ADR0(DLX_MEMinst_opcode_of_WB[4]),
    .ADR1(DLX_MEMinst_opcode_of_WB[3]),
    .ADR2(DLX_MEMinst_opcode_of_WB[1]),
    .ADR3(DLX_MEMinst_opcode_of_WB[5]),
    .O(\DLX_MEMinst_opcode_of_WB<1>/GROM )
  );
  X_BUF \DLX_MEMinst_opcode_of_WB<1>/YUSED  (
    .I(\DLX_MEMinst_opcode_of_WB<1>/GROM ),
    .O(DLX_IDinst__n0161)
  );
  defparam \Mshift__n0000_Sh<35>1 .INIT = 16'h2200;
  X_LUT4 \Mshift__n0000_Sh<35>1  (
    .ADR0(DLX_EXinst_ALU_result[13]),
    .ADR1(DLX_EXinst_ALU_result[14]),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_ALU_result[12]),
    .O(\DLX_IFinst_IR_previous<3>/FROM )
  );
  defparam Ker6303213.INIT = 16'hB1A0;
  X_LUT4 Ker6303213 (
    .ADR0(DLX_EXinst_ALU_result[14]),
    .ADR1(DLX_EXinst_ALU_result[13]),
    .ADR2(vram_out_cpu[4]),
    .ADR3(vram_out_cpu[0]),
    .O(\DLX_IFinst_IR_previous<3>/GROM )
  );
  X_BUF \DLX_IFinst_IR_previous<3>/XUSED  (
    .I(\DLX_IFinst_IR_previous<3>/FROM ),
    .O(Mshift__n0000_Sh[35])
  );
  X_BUF \DLX_IFinst_IR_previous<3>/YUSED  (
    .I(\DLX_IFinst_IR_previous<3>/GROM ),
    .O(CHOICE246)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5610.INIT = 16'h0080;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5610 (
    .ADR0(DLX_IDinst_jtarget[17]),
    .ADR1(DLX_IDinst_jtarget[19]),
    .ADR2(DLX_IDinst_jtarget[20]),
    .ADR3(DLX_IDinst_jtarget[18]),
    .O(\DLX_IDinst_RegFile_3_28/FROM )
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_571.INIT = 16'h0080;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_571 (
    .ADR0(DLX_IDinst_jtarget[18]),
    .ADR1(DLX_IDinst_jtarget[20]),
    .ADR2(DLX_IDinst_jtarget[19]),
    .ADR3(DLX_IDinst_jtarget[17]),
    .O(\DLX_IDinst_RegFile_3_28/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_3_28/XUSED  (
    .I(\DLX_IDinst_RegFile_3_28/FROM ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_56)
  );
  X_BUF \DLX_IDinst_RegFile_3_28/YUSED  (
    .I(\DLX_IDinst_RegFile_3_28/GROM ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_57)
  );
  defparam DLX_IFinst_IR_previous_9.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_9 (
    .I(DLX_IFinst_IR_latched[9]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[9])
  );
  defparam \Mshift__n0000_Sh<34>1 .INIT = 16'h1010;
  X_LUT4 \Mshift__n0000_Sh<34>1  (
    .ADR0(DLX_EXinst_ALU_result[12]),
    .ADR1(DLX_EXinst_ALU_result[14]),
    .ADR2(DLX_EXinst_ALU_result[13]),
    .ADR3(VCC),
    .O(\DLX_IFinst_IR_previous<9>/FROM )
  );
  defparam Ker6307113.INIT = 16'hCC0A;
  X_LUT4 Ker6307113 (
    .ADR0(RAM_read_data[0]),
    .ADR1(vram_out_cpu[3]),
    .ADR2(DLX_EXinst_ALU_result[13]),
    .ADR3(DLX_EXinst_ALU_result[14]),
    .O(\DLX_IFinst_IR_previous<9>/GROM )
  );
  X_BUF \DLX_IFinst_IR_previous<9>/XUSED  (
    .I(\DLX_IFinst_IR_previous<9>/FROM ),
    .O(Mshift__n0000_Sh[34])
  );
  X_BUF \DLX_IFinst_IR_previous<9>/YUSED  (
    .I(\DLX_IFinst_IR_previous<9>/GROM ),
    .O(CHOICE254)
  );
  defparam DLX_IDinst__n014940_SW0.INIT = 16'hB888;
  X_LUT4 DLX_IDinst__n014940_SW0 (
    .ADR0(DLX_IDinst__n0436),
    .ADR1(DLX_IDinst__n0434),
    .ADR2(DLX_IDinst__n0437),
    .ADR3(DLX_IDinst__n0439),
    .O(\N163210/FROM )
  );
  defparam DLX_IDinst__n014940.INIT = 16'h4540;
  X_LUT4 DLX_IDinst__n014940 (
    .ADR0(DLX_IDinst__n0166),
    .ADR1(DLX_IDinst__n0433),
    .ADR2(DLX_IDinst__n0167),
    .ADR3(N163210),
    .O(\N163210/GROM )
  );
  X_BUF \N163210/XUSED  (
    .I(\N163210/FROM ),
    .O(N163210)
  );
  X_BUF \N163210/YUSED  (
    .I(\N163210/GROM ),
    .O(CHOICE3487)
  );
  defparam \DLX_EXinst_Mshift__n0021_Sh<41>_SW0 .INIT = 16'h03CF;
  X_LUT4 \DLX_EXinst_Mshift__n0021_Sh<41>_SW0  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_Imm_3_1),
    .ADR2(\DLX_EXinst_Mshift__n0021_Sh[9] ),
    .ADR3(\DLX_EXinst_Mshift__n0021_Sh[1] ),
    .O(\DLX_IDinst_EPC<9>/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0021_Sh<41> .INIT = 16'h202F;
  X_LUT4 \DLX_EXinst_Mshift__n0021_Sh<41>  (
    .ADR0(\DLX_EXinst_Mshift__n0021_Sh[5] ),
    .ADR1(DLX_IDinst_Imm_3_1),
    .ADR2(DLX_IDinst_Imm_2_1),
    .ADR3(N131439),
    .O(\DLX_IDinst_EPC<9>/GROM )
  );
  X_BUF \DLX_IDinst_EPC<9>/XUSED  (
    .I(\DLX_IDinst_EPC<9>/FROM ),
    .O(N131439)
  );
  X_BUF \DLX_IDinst_EPC<9>/YUSED  (
    .I(\DLX_IDinst_EPC<9>/GROM ),
    .O(\DLX_EXinst_Mshift__n0021_Sh[41] )
  );
  defparam DLX_EXinst_Ker73996.INIT = 16'hAFA0;
  X_LUT4 DLX_EXinst_Ker73996 (
    .ADR0(\DLX_EXinst_Mshift__n0021_Sh[10] ),
    .ADR1(VCC),
    .ADR2(\DLX_IDinst_Imm[3] ),
    .ADR3(N130261),
    .O(\DLX_IDinst_RegFile_0_10/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0021_Sh<42>_SW0 .INIT = 16'h330F;
  X_LUT4 \DLX_EXinst_Mshift__n0021_Sh<42>_SW0  (
    .ADR0(VCC),
    .ADR1(\DLX_EXinst_Mshift__n0021_Sh[2] ),
    .ADR2(\DLX_EXinst_Mshift__n0021_Sh[10] ),
    .ADR3(DLX_IDinst_Imm_3_1),
    .O(\DLX_IDinst_RegFile_0_10/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_0_10/XUSED  (
    .I(\DLX_IDinst_RegFile_0_10/FROM ),
    .O(DLX_EXinst_N73998)
  );
  X_BUF \DLX_IDinst_RegFile_0_10/YUSED  (
    .I(\DLX_IDinst_RegFile_0_10/GROM ),
    .O(N131503)
  );
  defparam DLX_IDinst__n043141_SW0.INIT = 16'h75FE;
  X_LUT4 DLX_IDinst__n043141_SW0 (
    .ADR0(DLX_IDinst_IR_latched[31]),
    .ADR1(DLX_IDinst_IR_latched[26]),
    .ADR2(DLX_IDinst_IR_latched[27]),
    .ADR3(DLX_IDinst_IR_latched[29]),
    .O(\DLX_IDinst_RegFile_2_1/FROM )
  );
  defparam DLX_IDinst__n043141.INIT = 16'h0003;
  X_LUT4 DLX_IDinst__n043141 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_IR_latched[28]),
    .ADR2(DLX_IDinst_IR_latched[30]),
    .ADR3(N164562),
    .O(\DLX_IDinst_RegFile_2_1/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_2_1/XUSED  (
    .I(\DLX_IDinst_RegFile_2_1/FROM ),
    .O(N164562)
  );
  X_BUF \DLX_IDinst_RegFile_2_1/YUSED  (
    .I(\DLX_IDinst_RegFile_2_1/GROM ),
    .O(N137212)
  );
  defparam DLX_EXinst_Ker73991.INIT = 16'hF0AA;
  X_LUT4 DLX_EXinst_Ker73991 (
    .ADR0(N130209),
    .ADR1(VCC),
    .ADR2(\DLX_EXinst_Mshift__n0021_Sh[9] ),
    .ADR3(\DLX_IDinst_Imm[3] ),
    .O(\DLX_IDinst_RegFile_0_20/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0021_Sh<45>_SW0 .INIT = 16'hF5A0;
  X_LUT4 \DLX_EXinst_Mshift__n0021_Sh<45>_SW0  (
    .ADR0(DLX_IDinst_Imm_2_1),
    .ADR1(VCC),
    .ADR2(\DLX_EXinst_Mshift__n0021_Sh[9] ),
    .ADR3(\DLX_EXinst_Mshift__n0021_Sh[13] ),
    .O(\DLX_IDinst_RegFile_0_20/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_0_20/XUSED  (
    .I(\DLX_IDinst_RegFile_0_20/FROM ),
    .O(DLX_EXinst_N73993)
  );
  X_BUF \DLX_IDinst_RegFile_0_20/YUSED  (
    .I(\DLX_IDinst_RegFile_0_20/GROM ),
    .O(N130363)
  );
  defparam DLX_IDinst_RegFile_27_31_1439.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_27_31_1439 (
    .I(DLX_IDinst_WB_data_eff[31]),
    .CE(DLX_IDinst__n0604),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_27_31)
  );
  defparam vga_top_vga1__n000972_SW0.INIT = 16'hFFEA;
  X_LUT4 vga_top_vga1__n000972_SW0 (
    .ADR0(vga_top_vga1_helpme),
    .ADR1(vga_top_vga1_N112941),
    .ADR2(CHOICE3468),
    .ADR3(CHOICE3470),
    .O(\N163708/FROM )
  );
  defparam vga_top_vga1__n000972.INIT = 16'hFFA8;
  X_LUT4 vga_top_vga1__n000972 (
    .ADR0(vga_top_vga1_vcounter[9]),
    .ADR1(CHOICE3459),
    .ADR2(CHOICE3455),
    .ADR3(N163708),
    .O(\N163708/GROM )
  );
  X_BUF \N163708/XUSED  (
    .I(\N163708/FROM ),
    .O(N163708)
  );
  X_BUF \N163708/YUSED  (
    .I(\N163708/GROM ),
    .O(N147636)
  );
  defparam DLX_EXinst_Ker7437228.INIT = 16'h1AF0;
  X_LUT4 DLX_EXinst_Ker7437228 (
    .ADR0(DLX_IDinst_reg_out_B_2_1),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(DLX_IDinst_reg_out_B[5]),
    .ADR3(DLX_IDinst_reg_out_B[3]),
    .O(\DLX_IDinst_RegFile_30_31/FROM )
  );
  defparam DLX_EXinst_Ker74372107.INIT = 16'h00B8;
  X_LUT4 DLX_EXinst_Ker74372107 (
    .ADR0(\DLX_EXinst_Mshift__n0024_Sh[30] ),
    .ADR1(DLX_IDinst_reg_out_B[3]),
    .ADR2(\DLX_EXinst_Mshift__n0019_Sh[22] ),
    .ADR3(DLX_IDinst_reg_out_B_2_1),
    .O(\DLX_IDinst_RegFile_30_31/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_30_31/XUSED  (
    .I(\DLX_IDinst_RegFile_30_31/FROM ),
    .O(CHOICE3113)
  );
  X_BUF \DLX_IDinst_RegFile_30_31/YUSED  (
    .I(\DLX_IDinst_RegFile_30_31/GROM ),
    .O(CHOICE3130)
  );
  defparam DLX_IDinst_RegFile_19_24_1440.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_19_24_1440 (
    .I(DLX_IDinst_WB_data_eff[24]),
    .CE(DLX_IDinst__n0588),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_19_24)
  );
  defparam DLX_EXinst_Ker74372135.INIT = 16'hEEEC;
  X_LUT4 DLX_EXinst_Ker74372135 (
    .ADR0(DLX_EXinst_N76421),
    .ADR1(N163618),
    .ADR2(CHOICE3130),
    .ADR3(CHOICE3133),
    .O(\N145644/FROM )
  );
  defparam \DLX_EXinst__n0007<6>87 .INIT = 16'hECA0;
  X_LUT4 \DLX_EXinst__n0007<6>87  (
    .ADR0(DLX_EXinst_ALU_result[6]),
    .ADR1(DLX_IDinst_reg_out_B[4]),
    .ADR2(N134884),
    .ADR3(N145644),
    .O(\N145644/GROM )
  );
  X_BUF \N145644/XUSED  (
    .I(\N145644/FROM ),
    .O(N145644)
  );
  X_BUF \N145644/YUSED  (
    .I(\N145644/GROM ),
    .O(CHOICE3900)
  );
  defparam DLX_EXinst_Ker74367101.INIT = 16'hECA0;
  X_LUT4 DLX_EXinst_Ker74367101 (
    .ADR0(DLX_EXinst_N76421),
    .ADR1(CHOICE3036),
    .ADR2(CHOICE3043),
    .ADR3(N148609),
    .O(\N145073/FROM )
  );
  defparam \DLX_EXinst__n0007<5>87 .INIT = 16'hEAC0;
  X_LUT4 \DLX_EXinst__n0007<5>87  (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(DLX_EXinst_ALU_result[5]),
    .ADR2(N134884),
    .ADR3(N145073),
    .O(\N145073/GROM )
  );
  X_BUF \N145073/XUSED  (
    .I(\N145073/FROM ),
    .O(N145073)
  );
  X_BUF \N145073/YUSED  (
    .I(\N145073/GROM ),
    .O(CHOICE3959)
  );
  defparam DLX_EXinst_Ker7437715.INIT = 16'h5410;
  X_LUT4 DLX_EXinst_Ker7437715 (
    .ADR0(DLX_IDinst_reg_out_B_3_1),
    .ADR1(DLX_IDinst_reg_out_B_2_1),
    .ADR2(\DLX_EXinst_Mshift__n0019_Sh[23] ),
    .ADR3(\DLX_EXinst_Mshift__n0019_Sh[27] ),
    .O(\DLX_IDinst_RegFile_2_2/FROM )
  );
  defparam DLX_EXinst_Ker74377109.INIT = 16'h7250;
  X_LUT4 DLX_EXinst_Ker74377109 (
    .ADR0(DLX_IDinst_reg_out_B_2_1),
    .ADR1(DLX_IDinst_reg_out_B[3]),
    .ADR2(DLX_EXinst_N73103),
    .ADR3(\DLX_EXinst_Mshift__n0019_Sh[27] ),
    .O(\DLX_IDinst_RegFile_2_2/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_2_2/XUSED  (
    .I(\DLX_IDinst_RegFile_2_2/FROM ),
    .O(CHOICE3052)
  );
  X_BUF \DLX_IDinst_RegFile_2_2/YUSED  (
    .I(\DLX_IDinst_RegFile_2_2/GROM ),
    .O(CHOICE3072)
  );
  defparam DLX_EXinst_Ker74377118.INIT = 16'hEAC0;
  X_LUT4 DLX_EXinst_Ker74377118 (
    .ADR0(CHOICE3072),
    .ADR1(CHOICE3065),
    .ADR2(N148609),
    .ADR3(DLX_EXinst_N76421),
    .O(\N145258/FROM )
  );
  defparam \DLX_EXinst__n0007<7>87 .INIT = 16'hECA0;
  X_LUT4 \DLX_EXinst__n0007<7>87  (
    .ADR0(DLX_EXinst_ALU_result[7]),
    .ADR1(DLX_IDinst_reg_out_B[4]),
    .ADR2(N134884),
    .ADR3(N145258),
    .O(\N145258/GROM )
  );
  X_BUF \N145258/XUSED  (
    .I(\N145258/FROM ),
    .O(N145258)
  );
  X_BUF \N145258/YUSED  (
    .I(\N145258/GROM ),
    .O(CHOICE3841)
  );
  defparam DLX_EXinst_Ker74652107.INIT = 16'hECA0;
  X_LUT4 DLX_EXinst_Ker74652107 (
    .ADR0(CHOICE2938),
    .ADR1(CHOICE2945),
    .ADR2(N147520),
    .ADR3(DLX_EXinst_N76441),
    .O(\N144481/FROM )
  );
  defparam \DLX_EXinst__n0007<22>92 .INIT = 16'hD5C0;
  X_LUT4 \DLX_EXinst__n0007<22>92  (
    .ADR0(\DLX_IDinst_Imm[4] ),
    .ADR1(\DLX_IDinst_Imm[31] ),
    .ADR2(N163282),
    .ADR3(N144481),
    .O(\N144481/GROM )
  );
  X_BUF \N144481/XUSED  (
    .I(\N144481/FROM ),
    .O(N144481)
  );
  X_BUF \N144481/YUSED  (
    .I(\N144481/GROM ),
    .O(CHOICE4084)
  );
  defparam DLX_EXinst_Ker76181133.INIT = 16'h0001;
  X_LUT4 DLX_EXinst_Ker76181133 (
    .ADR0(DLX_IDinst_reg_out_B[7]),
    .ADR1(DLX_IDinst_reg_out_B[9]),
    .ADR2(DLX_IDinst_reg_out_B[8]),
    .ADR3(DLX_IDinst_reg_out_B[6]),
    .O(\DLX_IDinst_RegFile_2_3/FROM )
  );
  defparam DLX_EXinst_Ker76181134.INIT = 16'hCC00;
  X_LUT4 DLX_EXinst_Ker76181134 (
    .ADR0(VCC),
    .ADR1(CHOICE3639),
    .ADR2(VCC),
    .ADR3(CHOICE3646),
    .O(\DLX_IDinst_RegFile_2_3/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_2_3/XUSED  (
    .I(\DLX_IDinst_RegFile_2_3/FROM ),
    .O(CHOICE3646)
  );
  X_BUF \DLX_IDinst_RegFile_2_3/YUSED  (
    .I(\DLX_IDinst_RegFile_2_3/GROM ),
    .O(CHOICE3647)
  );
  defparam DLX_EXinst_Ker74647108.INIT = 16'hF888;
  X_LUT4 DLX_EXinst_Ker74647108 (
    .ADR0(CHOICE2972),
    .ADR1(DLX_EXinst_N76441),
    .ADR2(CHOICE2965),
    .ADR3(N147520),
    .O(\N144646/FROM )
  );
  defparam \DLX_EXinst__n0007<21>92 .INIT = 16'hB3A0;
  X_LUT4 \DLX_EXinst__n0007<21>92  (
    .ADR0(\DLX_IDinst_Imm[31] ),
    .ADR1(\DLX_IDinst_Imm[4] ),
    .ADR2(N163704),
    .ADR3(N144646),
    .O(\N144646/GROM )
  );
  X_BUF \N144646/XUSED  (
    .I(\N144646/FROM ),
    .O(N144646)
  );
  X_BUF \N144646/YUSED  (
    .I(\N144646/GROM ),
    .O(CHOICE4149)
  );
  defparam DLX_EXinst_Ker76159129.INIT = 16'h0001;
  X_LUT4 DLX_EXinst_Ker76159129 (
    .ADR0(\DLX_IDinst_Imm[8] ),
    .ADR1(\DLX_IDinst_Imm[9] ),
    .ADR2(\DLX_IDinst_Imm[7] ),
    .ADR3(\DLX_IDinst_Imm[10] ),
    .O(\CHOICE3449/FROM )
  );
  defparam DLX_EXinst_Ker76159153.INIT = 16'h1000;
  X_LUT4 DLX_EXinst_Ker76159153 (
    .ADR0(\DLX_IDinst_Imm[31] ),
    .ADR1(\DLX_IDinst_Imm[15] ),
    .ADR2(CHOICE3442),
    .ADR3(CHOICE3449),
    .O(\CHOICE3449/GROM )
  );
  X_BUF \CHOICE3449/XUSED  (
    .I(\CHOICE3449/FROM ),
    .O(CHOICE3449)
  );
  X_BUF \CHOICE3449/YUSED  (
    .I(\CHOICE3449/GROM ),
    .O(CHOICE3451)
  );
  defparam DLX_EXinst_Ker7464713.INIT = 16'hA820;
  X_LUT4 DLX_EXinst_Ker7464713 (
    .ADR0(DLX_IDinst_Imm_2_1),
    .ADR1(DLX_IDinst_Imm_3_1),
    .ADR2(\DLX_EXinst_Mshift__n0020_Sh[25] ),
    .ADR3(DLX_IDinst_reg_out_A[31]),
    .O(\DLX_IDinst_RegFile_2_4/FROM )
  );
  defparam DLX_EXinst_Ker74657109.INIT = 16'h7250;
  X_LUT4 DLX_EXinst_Ker74657109 (
    .ADR0(DLX_IDinst_Imm_2_1),
    .ADR1(DLX_IDinst_Imm_3_1),
    .ADR2(DLX_EXinst_N73168),
    .ADR3(\DLX_EXinst_Mshift__n0020_Sh[27] ),
    .O(\DLX_IDinst_RegFile_2_4/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_2_4/XUSED  (
    .I(\DLX_IDinst_RegFile_2_4/FROM ),
    .O(CHOICE2953)
  );
  X_BUF \DLX_IDinst_RegFile_2_4/YUSED  (
    .I(\DLX_IDinst_RegFile_2_4/GROM ),
    .O(CHOICE3101)
  );
  defparam DLX_EXinst_Ker74657118.INIT = 16'hF888;
  X_LUT4 DLX_EXinst_Ker74657118 (
    .ADR0(N147520),
    .ADR1(CHOICE3094),
    .ADR2(CHOICE3101),
    .ADR3(DLX_EXinst_N76441),
    .O(\N145443/FROM )
  );
  defparam \DLX_EXinst__n0007<23>92 .INIT = 16'hB3A0;
  X_LUT4 \DLX_EXinst__n0007<23>92  (
    .ADR0(N163460),
    .ADR1(\DLX_IDinst_Imm[4] ),
    .ADR2(\DLX_IDinst_Imm[31] ),
    .ADR3(N145443),
    .O(\N145443/GROM )
  );
  X_BUF \N145443/XUSED  (
    .I(\N145443/FROM ),
    .O(N145443)
  );
  X_BUF \N145443/YUSED  (
    .I(\N145443/GROM ),
    .O(CHOICE4019)
  );
  defparam DLX_EXinst_ALU_result_7.INIT = 1'b0;
  X_SFF DLX_EXinst_ALU_result_7 (
    .I(N162807),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(N136886),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_ALU_result[7])
  );
  defparam DLX_IDinst__n01161.INIT = 16'hC0EA;
  X_LUT4 DLX_IDinst__n01161 (
    .ADR0(DLX_EXinst__n0144),
    .ADR1(DLX_IDinst_delay_slot),
    .ADR2(DLX_IDinst_slot_num_FFd2),
    .ADR3(DLX_IDinst_stall),
    .O(\DLX_IDinst_RegFile_31_13/FROM )
  );
  defparam DLX_IDinst__n06371.INIT = 16'hAAFF;
  X_LUT4 DLX_IDinst__n06371 (
    .ADR0(DLX_IDinst__n0387),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst__n0116),
    .O(\DLX_IDinst_RegFile_31_13/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_31_13/XUSED  (
    .I(\DLX_IDinst_RegFile_31_13/FROM ),
    .O(DLX_IDinst__n0116)
  );
  X_BUF \DLX_IDinst_RegFile_31_13/YUSED  (
    .I(\DLX_IDinst_RegFile_31_13/GROM ),
    .O(DLX_IDinst__n0637)
  );
  defparam DLX_IDinst__n03111.INIT = 16'h0008;
  X_LUT4 DLX_IDinst__n03111 (
    .ADR0(DLX_IDinst_IR_latched[30]),
    .ADR1(DLX_IDinst_IR_latched[27]),
    .ADR2(DLX_IDinst_IR_latched[28]),
    .ADR3(DLX_IDinst_IR_latched[26]),
    .O(\DLX_IDinst__n0311/FROM )
  );
  defparam DLX_IDinst__n011715.INIT = 16'hCC80;
  X_LUT4 DLX_IDinst__n011715 (
    .ADR0(DLX_IDinst__n0462),
    .ADR1(DLX_IDinst_N108443),
    .ADR2(DLX_IDinst_N108221),
    .ADR3(DLX_IDinst__n0311),
    .O(\DLX_IDinst__n0311/GROM )
  );
  X_BUF \DLX_IDinst__n0311/XUSED  (
    .I(\DLX_IDinst__n0311/FROM ),
    .O(DLX_IDinst__n0311)
  );
  X_BUF \DLX_IDinst__n0311/YUSED  (
    .I(\DLX_IDinst__n0311/GROM ),
    .O(CHOICE3352)
  );
  defparam DLX_IDinst__n01519.INIT = 16'hFFFE;
  X_LUT4 DLX_IDinst__n01519 (
    .ADR0(DLX_IDinst_IR_latched[29]),
    .ADR1(DLX_IDinst_IR_latched[31]),
    .ADR2(DLX_IDinst_IR_latched[28]),
    .ADR3(DLX_IDinst_IR_latched[27]),
    .O(\CHOICE3321/FROM )
  );
  defparam DLX_IDinst__n015119.INIT = 16'hF0D0;
  X_LUT4 DLX_IDinst__n015119 (
    .ADR0(DLX_IDinst_IR_latched[30]),
    .ADR1(DLX_IDinst_IR_latched[26]),
    .ADR2(DLX_IDinst_delay_slot),
    .ADR3(CHOICE3321),
    .O(\CHOICE3321/GROM )
  );
  X_BUF \CHOICE3321/XUSED  (
    .I(\CHOICE3321/FROM ),
    .O(CHOICE3321)
  );
  X_BUF \CHOICE3321/YUSED  (
    .I(\CHOICE3321/GROM ),
    .O(CHOICE3323)
  );
  defparam DLX_IDinst_Ker107607_SW0.INIT = 16'hF000;
  X_LUT4 DLX_IDinst_Ker107607_SW0 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_N108165),
    .ADR3(DLX_IDinst_IR_latched[27]),
    .O(\DLX_IDinst_RegFile_31_22/FROM )
  );
  defparam DLX_IDinst__n01631.INIT = 16'hFEFF;
  X_LUT4 DLX_IDinst__n01631 (
    .ADR0(DLX_IDinst_IR_latched[28]),
    .ADR1(DLX_IDinst_IR_latched[29]),
    .ADR2(DLX_IDinst_IR_latched[31]),
    .ADR3(DLX_IDinst_IR_latched[27]),
    .O(\DLX_IDinst_RegFile_31_22/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_31_22/XUSED  (
    .I(\DLX_IDinst_RegFile_31_22/FROM ),
    .O(N136696)
  );
  X_BUF \DLX_IDinst_RegFile_31_22/YUSED  (
    .I(\DLX_IDinst_RegFile_31_22/GROM ),
    .O(DLX_IDinst__n0163)
  );
  defparam DLX_IDinst__n04341.INIT = 16'hCCC4;
  X_LUT4 DLX_IDinst__n04341 (
    .ADR0(DLX_IDinst_N108244),
    .ADR1(DLX_IDinst__n0104),
    .ADR2(DLX_IDinst_jtarget[21]),
    .ADR3(DLX_IDinst_jtarget[22]),
    .O(\DLX_IDinst_RegFile_15_31/FROM )
  );
  defparam DLX_IDinst__n01661.INIT = 16'hF0D0;
  X_LUT4 DLX_IDinst__n01661 (
    .ADR0(DLX_IDinst_N108244),
    .ADR1(DLX_IDinst_jtarget[22]),
    .ADR2(DLX_IDinst__n0100),
    .ADR3(DLX_IDinst_jtarget[21]),
    .O(\DLX_IDinst_RegFile_15_31/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_15_31/XUSED  (
    .I(\DLX_IDinst_RegFile_15_31/FROM ),
    .O(DLX_IDinst__n0434)
  );
  X_BUF \DLX_IDinst_RegFile_15_31/YUSED  (
    .I(\DLX_IDinst_RegFile_15_31/GROM ),
    .O(DLX_IDinst__n0166)
  );
  defparam DLX_IDinst__n01671.INIT = 16'h00F0;
  X_LUT4 DLX_IDinst__n01671 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IDinst__n0102),
    .ADR3(DLX_IDinst__n0381),
    .O(\DLX_IDinst_RegFile_31_16/FROM )
  );
  defparam DLX_IDinst_Ker1081501.INIT = 16'h000B;
  X_LUT4 DLX_IDinst_Ker1081501 (
    .ADR0(DLX_IDinst__n0382),
    .ADR1(DLX_IDinst__n0100),
    .ADR2(DLX_IDinst__n0434),
    .ADR3(DLX_IDinst__n0167),
    .O(\DLX_IDinst_RegFile_31_16/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_31_16/XUSED  (
    .I(\DLX_IDinst_RegFile_31_16/FROM ),
    .O(DLX_IDinst__n0167)
  );
  X_BUF \DLX_IDinst_RegFile_31_16/YUSED  (
    .I(\DLX_IDinst_RegFile_31_16/GROM ),
    .O(DLX_IDinst_N108152)
  );
  defparam DLX_IDinst__n01751.INIT = 16'h0088;
  X_LUT4 DLX_IDinst__n01751 (
    .ADR0(DLX_IDinst__n0367),
    .ADR1(DLX_MEMinst_reg_write_MEM),
    .ADR2(VCC),
    .ADR3(DLX_IDinst__n0382),
    .O(\DLX_IDinst_RegFile_15_18/FROM )
  );
  defparam \DLX_IDinst_Mmux_regA_eff_Result<27>1 .INIT = 16'hF0AA;
  X_LUT4 \DLX_IDinst_Mmux_regA_eff_Result<27>1  (
    .ADR0(DLX_IDinst__n0620[27]),
    .ADR1(VCC),
    .ADR2(DLX_MEMinst_RF_data_in[27]),
    .ADR3(DLX_IDinst__n0175),
    .O(\DLX_IDinst_RegFile_15_18/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_15_18/XUSED  (
    .I(\DLX_IDinst_RegFile_15_18/FROM ),
    .O(DLX_IDinst__n0175)
  );
  X_BUF \DLX_IDinst_RegFile_15_18/YUSED  (
    .I(\DLX_IDinst_RegFile_15_18/GROM ),
    .O(\DLX_IDinst_regA_eff[27] )
  );
  defparam DLX_IDinst_Ker10707436.INIT = 16'h5511;
  X_LUT4 DLX_IDinst_Ker10707436 (
    .ADR0(DLX_IDinst__n0434),
    .ADR1(DLX_IDinst__n0102),
    .ADR2(VCC),
    .ADR3(DLX_IDinst__n0381),
    .O(\DLX_IDinst_RegFile_15_19/FROM )
  );
  defparam DLX_IDinst__n01761.INIT = 16'h5000;
  X_LUT4 DLX_IDinst__n01761 (
    .ADR0(DLX_IDinst__n0381),
    .ADR1(VCC),
    .ADR2(DLX_IDinst__n0368),
    .ADR3(DLX_MEMinst_reg_write_MEM),
    .O(\DLX_IDinst_RegFile_15_19/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_15_19/XUSED  (
    .I(\DLX_IDinst_RegFile_15_19/FROM ),
    .O(CHOICE2118)
  );
  X_BUF \DLX_IDinst_RegFile_15_19/YUSED  (
    .I(\DLX_IDinst_RegFile_15_19/GROM ),
    .O(DLX_IDinst__n0176)
  );
  defparam DLX_IDinst__n05841.INIT = 16'h0500;
  X_LUT4 DLX_IDinst__n05841 (
    .ADR0(DLX_MEMinst_reg_dst_out[3]),
    .ADR1(VCC),
    .ADR2(DLX_MEMinst_reg_dst_out[1]),
    .ADR3(DLX_IDinst_N108531),
    .O(\DLX_IDinst_RegFile_19_0/FROM )
  );
  defparam DLX_IDinst__n06001.INIT = 16'h0A00;
  X_LUT4 DLX_IDinst__n06001 (
    .ADR0(DLX_IDinst_N108531),
    .ADR1(VCC),
    .ADR2(DLX_MEMinst_reg_dst_out[1]),
    .ADR3(DLX_MEMinst_reg_dst_out[3]),
    .O(\DLX_IDinst_RegFile_19_0/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_19_0/XUSED  (
    .I(\DLX_IDinst_RegFile_19_0/FROM ),
    .O(DLX_IDinst__n0584)
  );
  X_BUF \DLX_IDinst_RegFile_19_0/YUSED  (
    .I(\DLX_IDinst_RegFile_19_0/GROM ),
    .O(DLX_IDinst__n0600)
  );
  defparam DLX_IDinst__n00971.INIT = 16'h0080;
  X_LUT4 DLX_IDinst__n00971 (
    .ADR0(DLX_IDinst_IR_latched[26]),
    .ADR1(DLX_IDinst_IR_latched[30]),
    .ADR2(DLX_IDinst_N108165),
    .ADR3(DLX_IDinst_IR_latched[27]),
    .O(\DLX_IDinst__n0097/FROM )
  );
  defparam DLX_IDinst__n04531.INIT = 16'hFF04;
  X_LUT4 DLX_IDinst__n04531 (
    .ADR0(DLX_IDinst_CLI),
    .ADR1(INT_IBUF),
    .ADR2(DLX_IDinst_delay_slot),
    .ADR3(DLX_IDinst__n0097),
    .O(\DLX_IDinst__n0097/GROM )
  );
  X_BUF \DLX_IDinst__n0097/XUSED  (
    .I(\DLX_IDinst__n0097/FROM ),
    .O(DLX_IDinst__n0097)
  );
  X_BUF \DLX_IDinst__n0097/YUSED  (
    .I(\DLX_IDinst__n0097/GROM ),
    .O(DLX_IDinst__n0453)
  );
  defparam DLX_IDinst__n01951.INIT = 16'h0010;
  X_LUT4 DLX_IDinst__n01951 (
    .ADR0(DLX_IDinst_IR_latched[26]),
    .ADR1(DLX_IDinst_IR_latched[27]),
    .ADR2(DLX_IDinst_N108165),
    .ADR3(DLX_IDinst_IR_latched[30]),
    .O(\DLX_IDinst__n0629<1>/FROM )
  );
  defparam DLX_IDinst_Ker10720631.INIT = 16'hC0EA;
  X_LUT4 DLX_IDinst_Ker10720631 (
    .ADR0(N163562),
    .ADR1(CHOICE2103),
    .ADR2(DLX_IDinst_N108496),
    .ADR3(DLX_IDinst__n0629[1]),
    .O(\DLX_IDinst__n0629<1>/GROM )
  );
  X_BUF \DLX_IDinst__n0629<1>/XUSED  (
    .I(\DLX_IDinst__n0629<1>/FROM ),
    .O(DLX_IDinst__n0629[1])
  );
  X_BUF \DLX_IDinst__n0629<1>/YUSED  (
    .I(\DLX_IDinst__n0629<1>/GROM ),
    .O(N139563)
  );
  defparam DLX_IDinst__n04361.INIT = 16'hFEF0;
  X_LUT4 DLX_IDinst__n04361 (
    .ADR0(CHOICE1989),
    .ADR1(CHOICE1994),
    .ADR2(N135272),
    .ADR3(DLX_IDinst_N108254),
    .O(\DLX_IDinst__n0436/GROM )
  );
  X_BUF \DLX_IDinst__n0436/YUSED  (
    .I(\DLX_IDinst__n0436/GROM ),
    .O(DLX_IDinst__n0436)
  );
  defparam DLX_IDinst__n04371.INIT = 16'h00AA;
  X_LUT4 DLX_IDinst__n04371 (
    .ADR0(DLX_IDinst__n0105),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst__n0381),
    .O(\DLX_IFinst_IR_curr<13>/FROM )
  );
  defparam DLX_IDinst_Ker1084631.INIT = 16'h0700;
  X_LUT4 DLX_IDinst_Ker1084631 (
    .ADR0(N137212),
    .ADR1(DLX_IDinst_N108254),
    .ADR2(N135272),
    .ADR3(DLX_IDinst__n0437),
    .O(\DLX_IFinst_IR_curr<13>/GROM )
  );
  X_BUF \DLX_IFinst_IR_curr<13>/XUSED  (
    .I(\DLX_IFinst_IR_curr<13>/FROM ),
    .O(DLX_IDinst__n0437)
  );
  X_BUF \DLX_IFinst_IR_curr<13>/YUSED  (
    .I(\DLX_IFinst_IR_curr<13>/GROM ),
    .O(DLX_IDinst_N108465)
  );
  defparam DLX_IDinst_RegFile_24_30_1441.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_24_30_1441 (
    .I(DLX_IDinst_WB_data_eff[30]),
    .CE(DLX_IDinst__n0598),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_24_30)
  );
  defparam DLX_IDinst__n05661.INIT = 16'h2020;
  X_LUT4 DLX_IDinst__n05661 (
    .ADR0(DLX_MEMinst_reg_dst_out[3]),
    .ADR1(DLX_MEMinst_reg_dst_out[1]),
    .ADR2(DLX_IDinst_N108517),
    .ADR3(VCC),
    .O(\DLX_IDinst_RegFile_24_30/FROM )
  );
  defparam DLX_IDinst__n05501.INIT = 16'h1100;
  X_LUT4 DLX_IDinst__n05501 (
    .ADR0(DLX_MEMinst_reg_dst_out[3]),
    .ADR1(DLX_MEMinst_reg_dst_out[1]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_N108517),
    .O(\DLX_IDinst_RegFile_24_30/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_24_30/XUSED  (
    .I(\DLX_IDinst_RegFile_24_30/FROM ),
    .O(DLX_IDinst__n0566)
  );
  X_BUF \DLX_IDinst_RegFile_24_30/YUSED  (
    .I(\DLX_IDinst_RegFile_24_30/GROM ),
    .O(DLX_IDinst__n0550)
  );
  defparam DLX_IDinst__n05901.INIT = 16'h0202;
  X_LUT4 DLX_IDinst__n05901 (
    .ADR0(DLX_IDinst_N108545),
    .ADR1(DLX_MEMinst_reg_dst_out[3]),
    .ADR2(DLX_MEMinst_reg_dst_out[1]),
    .ADR3(VCC),
    .O(\DLX_IFinst_IR_curr<30>/FROM )
  );
  defparam DLX_IDinst__n06061.INIT = 16'h2020;
  X_LUT4 DLX_IDinst__n06061 (
    .ADR0(DLX_IDinst_N108545),
    .ADR1(DLX_MEMinst_reg_dst_out[1]),
    .ADR2(DLX_MEMinst_reg_dst_out[3]),
    .ADR3(VCC),
    .O(\DLX_IFinst_IR_curr<30>/GROM )
  );
  X_BUF \DLX_IFinst_IR_curr<30>/XUSED  (
    .I(\DLX_IFinst_IR_curr<30>/FROM ),
    .O(DLX_IDinst__n0590)
  );
  X_BUF \DLX_IFinst_IR_curr<30>/YUSED  (
    .I(\DLX_IFinst_IR_curr<30>/GROM ),
    .O(DLX_IDinst__n0606)
  );
  defparam DLX_IDinst_RegFile_17_17_1442.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_17_17_1442 (
    .I(DLX_IDinst_WB_data_eff[17]),
    .CE(DLX_IDinst__n0584),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_17_17)
  );
  defparam DLX_IDinst_Ker107171_SW0.INIT = 16'hDDDD;
  X_LUT4 DLX_IDinst_Ker107171_SW0 (
    .ADR0(DLX_IDinst__n0116),
    .ADR1(DLX_IDinst__n0387),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IDinst_RegFile_17_17/FROM )
  );
  defparam DLX_IDinst__n06141.INIT = 16'hFFBB;
  X_LUT4 DLX_IDinst__n06141 (
    .ADR0(DLX_IDinst_N108249),
    .ADR1(DLX_IDinst__n0387),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_stall),
    .O(\DLX_IDinst_RegFile_17_17/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_17_17/XUSED  (
    .I(\DLX_IDinst_RegFile_17_17/FROM ),
    .O(N127094)
  );
  X_BUF \DLX_IDinst_RegFile_17_17/YUSED  (
    .I(\DLX_IDinst_RegFile_17_17/GROM ),
    .O(DLX_IDinst__n0614)
  );
  defparam DLX_IDinst__n05561.INIT = 16'h2200;
  X_LUT4 DLX_IDinst__n05561 (
    .ADR0(DLX_MEMinst_reg_dst_out[1]),
    .ADR1(DLX_MEMinst_reg_dst_out[3]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_N108510),
    .O(\DLX_IFinst_IR_curr<22>/FROM )
  );
  defparam DLX_IDinst__n05521.INIT = 16'h0500;
  X_LUT4 DLX_IDinst__n05521 (
    .ADR0(DLX_MEMinst_reg_dst_out[1]),
    .ADR1(VCC),
    .ADR2(DLX_MEMinst_reg_dst_out[3]),
    .ADR3(DLX_IDinst_N108510),
    .O(\DLX_IFinst_IR_curr<22>/GROM )
  );
  X_BUF \DLX_IFinst_IR_curr<22>/XUSED  (
    .I(\DLX_IFinst_IR_curr<22>/FROM ),
    .O(DLX_IDinst__n0556)
  );
  X_BUF \DLX_IFinst_IR_curr<22>/YUSED  (
    .I(\DLX_IFinst_IR_curr<22>/GROM ),
    .O(DLX_IDinst__n0552)
  );
  defparam DLX_IDinst__n05641.INIT = 16'h5000;
  X_LUT4 DLX_IDinst__n05641 (
    .ADR0(DLX_MEMinst_reg_dst_out[3]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_N108538),
    .ADR3(DLX_MEMinst_reg_dst_out[1]),
    .O(\DLX_IFinst_IR_curr<14>/FROM )
  );
  defparam DLX_IDinst__n05601.INIT = 16'h0050;
  X_LUT4 DLX_IDinst__n05601 (
    .ADR0(DLX_MEMinst_reg_dst_out[3]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_N108538),
    .ADR3(DLX_MEMinst_reg_dst_out[1]),
    .O(\DLX_IFinst_IR_curr<14>/GROM )
  );
  X_BUF \DLX_IFinst_IR_curr<14>/XUSED  (
    .I(\DLX_IFinst_IR_curr<14>/FROM ),
    .O(DLX_IDinst__n0564)
  );
  X_BUF \DLX_IFinst_IR_curr<14>/YUSED  (
    .I(\DLX_IFinst_IR_curr<14>/GROM ),
    .O(DLX_IDinst__n0560)
  );
  defparam DLX_IFinst_IR_curr_23.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_23 (
    .I(IR[23]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[23])
  );
  defparam DLX_IDinst__n05921.INIT = 16'h0202;
  X_LUT4 DLX_IDinst__n05921 (
    .ADR0(DLX_IDinst_N108524),
    .ADR1(DLX_MEMinst_reg_dst_out[1]),
    .ADR2(DLX_MEMinst_reg_dst_out[3]),
    .ADR3(VCC),
    .O(\DLX_IFinst_IR_curr<23>/FROM )
  );
  defparam DLX_IDinst__n06081.INIT = 16'h0808;
  X_LUT4 DLX_IDinst__n06081 (
    .ADR0(DLX_MEMinst_reg_dst_out[3]),
    .ADR1(DLX_IDinst_N108524),
    .ADR2(DLX_MEMinst_reg_dst_out[1]),
    .ADR3(VCC),
    .O(\DLX_IFinst_IR_curr<23>/GROM )
  );
  X_BUF \DLX_IFinst_IR_curr<23>/XUSED  (
    .I(\DLX_IFinst_IR_curr<23>/FROM ),
    .O(DLX_IDinst__n0592)
  );
  X_BUF \DLX_IFinst_IR_curr<23>/YUSED  (
    .I(\DLX_IFinst_IR_curr<23>/GROM ),
    .O(DLX_IDinst__n0608)
  );
  defparam DLX_IDinst_RegFile_19_29_1443.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_19_29_1443 (
    .I(DLX_IDinst_WB_data_eff[29]),
    .CE(DLX_IDinst__n0588),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_19_29)
  );
  defparam DLX_IDinst__n05581.INIT = 16'h0202;
  X_LUT4 DLX_IDinst__n05581 (
    .ADR0(DLX_IDinst_N108559),
    .ADR1(DLX_MEMinst_reg_dst_out[3]),
    .ADR2(DLX_MEMinst_reg_dst_out[1]),
    .ADR3(VCC),
    .O(\DLX_IDinst_RegFile_19_29/FROM )
  );
  defparam DLX_IDinst__n05701.INIT = 16'h8080;
  X_LUT4 DLX_IDinst__n05701 (
    .ADR0(DLX_IDinst_N108517),
    .ADR1(DLX_MEMinst_reg_dst_out[3]),
    .ADR2(DLX_MEMinst_reg_dst_out[1]),
    .ADR3(VCC),
    .O(\DLX_IDinst_RegFile_19_29/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_19_29/XUSED  (
    .I(\DLX_IDinst_RegFile_19_29/FROM ),
    .O(DLX_IDinst__n0558)
  );
  X_BUF \DLX_IDinst_RegFile_19_29/YUSED  (
    .I(\DLX_IDinst_RegFile_19_29/GROM ),
    .O(DLX_IDinst__n0570)
  );
  defparam DLX_IDinst_RegFile_19_16_1444.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_19_16_1444 (
    .I(DLX_IDinst_WB_data_eff[16]),
    .CE(DLX_IDinst__n0588),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_19_16)
  );
  defparam DLX_IDinst__n05741.INIT = 16'h2020;
  X_LUT4 DLX_IDinst__n05741 (
    .ADR0(DLX_IDinst_N108559),
    .ADR1(DLX_MEMinst_reg_dst_out[1]),
    .ADR2(DLX_MEMinst_reg_dst_out[3]),
    .ADR3(VCC),
    .O(\DLX_IDinst_RegFile_0_3/FROM )
  );
  defparam DLX_IDinst__n05621.INIT = 16'h0808;
  X_LUT4 DLX_IDinst__n05621 (
    .ADR0(DLX_IDinst_N108559),
    .ADR1(DLX_MEMinst_reg_dst_out[1]),
    .ADR2(DLX_MEMinst_reg_dst_out[3]),
    .ADR3(VCC),
    .O(\DLX_IDinst_RegFile_0_3/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_0_3/XUSED  (
    .I(\DLX_IDinst_RegFile_0_3/FROM ),
    .O(DLX_IDinst__n0574)
  );
  X_BUF \DLX_IDinst_RegFile_0_3/YUSED  (
    .I(\DLX_IDinst_RegFile_0_3/GROM ),
    .O(DLX_IDinst__n0562)
  );
  defparam DLX_IDinst_Ker108226114.INIT = 16'h3313;
  X_LUT4 DLX_IDinst_Ker108226114 (
    .ADR0(DLX_IDinst_N108503),
    .ADR1(DLX_IDinst__n0097),
    .ADR2(DLX_IDinst_IR_latched[27]),
    .ADR3(DLX_IDinst_IR_latched[30]),
    .O(\DLX_EXinst_ALU_result<5>/FROM )
  );
  defparam DLX_IDinst__n06351.INIT = 16'h00EA;
  X_LUT4 DLX_IDinst__n06351 (
    .ADR0(DLX_IDinst_Ker1084541_1),
    .ADR1(DLX_IDinst_IR_latched[27]),
    .ADR2(DLX_IDinst_N108503),
    .ADR3(DLX_IDinst_IR_latched[30]),
    .O(\DLX_EXinst_ALU_result<5>/GROM )
  );
  X_BUF \DLX_EXinst_ALU_result<5>/XUSED  (
    .I(\DLX_EXinst_ALU_result<5>/FROM ),
    .O(CHOICE3396)
  );
  X_BUF \DLX_EXinst_ALU_result<5>/YUSED  (
    .I(\DLX_EXinst_ALU_result<5>/GROM ),
    .O(DLX_IDinst__n0635)
  );
  defparam DLX_IDinst__n05861.INIT = 16'h3000;
  X_LUT4 DLX_IDinst__n05861 (
    .ADR0(VCC),
    .ADR1(DLX_MEMinst_reg_dst_out[3]),
    .ADR2(DLX_IDinst_N108552),
    .ADR3(DLX_MEMinst_reg_dst_out[1]),
    .O(\DLX_IDinst_RegFile_23_1/FROM )
  );
  defparam DLX_IDinst__n05821.INIT = 16'h1010;
  X_LUT4 DLX_IDinst__n05821 (
    .ADR0(DLX_MEMinst_reg_dst_out[1]),
    .ADR1(DLX_MEMinst_reg_dst_out[3]),
    .ADR2(DLX_IDinst_N108552),
    .ADR3(VCC),
    .O(\DLX_IDinst_RegFile_23_1/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_23_1/XUSED  (
    .I(\DLX_IDinst_RegFile_23_1/FROM ),
    .O(DLX_IDinst__n0586)
  );
  X_BUF \DLX_IDinst_RegFile_23_1/YUSED  (
    .I(\DLX_IDinst_RegFile_23_1/GROM ),
    .O(DLX_IDinst__n0582)
  );
  defparam DLX_IDinst__n05761.INIT = 16'h2200;
  X_LUT4 DLX_IDinst__n05761 (
    .ADR0(DLX_MEMinst_reg_dst_out[3]),
    .ADR1(DLX_MEMinst_reg_dst_out[1]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_N108538),
    .O(\DLX_IDinst_RegFile_14_6/FROM )
  );
  defparam DLX_IDinst__n05681.INIT = 16'h00A0;
  X_LUT4 DLX_IDinst__n05681 (
    .ADR0(DLX_IDinst_N108510),
    .ADR1(VCC),
    .ADR2(DLX_MEMinst_reg_dst_out[3]),
    .ADR3(DLX_MEMinst_reg_dst_out[1]),
    .O(\DLX_IDinst_RegFile_14_6/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_14_6/XUSED  (
    .I(\DLX_IDinst_RegFile_14_6/FROM ),
    .O(DLX_IDinst__n0576)
  );
  X_BUF \DLX_IDinst_RegFile_14_6/YUSED  (
    .I(\DLX_IDinst_RegFile_14_6/GROM ),
    .O(DLX_IDinst__n0568)
  );
  defparam DLX_IDinst__n05881.INIT = 16'h0088;
  X_LUT4 DLX_IDinst__n05881 (
    .ADR0(DLX_IDinst_N108531),
    .ADR1(DLX_MEMinst_reg_dst_out[1]),
    .ADR2(VCC),
    .ADR3(DLX_MEMinst_reg_dst_out[3]),
    .O(\DLX_IDinst_RegFile_0_5/FROM )
  );
  defparam DLX_IDinst__n05941.INIT = 16'h00A0;
  X_LUT4 DLX_IDinst__n05941 (
    .ADR0(DLX_IDinst_N108545),
    .ADR1(VCC),
    .ADR2(DLX_MEMinst_reg_dst_out[1]),
    .ADR3(DLX_MEMinst_reg_dst_out[3]),
    .O(\DLX_IDinst_RegFile_0_5/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_0_5/XUSED  (
    .I(\DLX_IDinst_RegFile_0_5/FROM ),
    .O(DLX_IDinst__n0588)
  );
  X_BUF \DLX_IDinst_RegFile_0_5/YUSED  (
    .I(\DLX_IDinst_RegFile_0_5/GROM ),
    .O(DLX_IDinst__n0594)
  );
  defparam DLX_IDinst__n05981.INIT = 16'h0088;
  X_LUT4 DLX_IDinst__n05981 (
    .ADR0(DLX_IDinst_N108552),
    .ADR1(DLX_MEMinst_reg_dst_out[3]),
    .ADR2(VCC),
    .ADR3(DLX_MEMinst_reg_dst_out[1]),
    .O(\DLX_IFinst_IR_curr<17>/FROM )
  );
  defparam DLX_IDinst__n05961.INIT = 16'h5000;
  X_LUT4 DLX_IDinst__n05961 (
    .ADR0(DLX_MEMinst_reg_dst_out[3]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_N108524),
    .ADR3(DLX_MEMinst_reg_dst_out[1]),
    .O(\DLX_IFinst_IR_curr<17>/GROM )
  );
  X_BUF \DLX_IFinst_IR_curr<17>/XUSED  (
    .I(\DLX_IFinst_IR_curr<17>/FROM ),
    .O(DLX_IDinst__n0598)
  );
  X_BUF \DLX_IFinst_IR_curr<17>/YUSED  (
    .I(\DLX_IFinst_IR_curr<17>/GROM ),
    .O(DLX_IDinst__n0596)
  );
  defparam \DLX_EXinst__n0007<10>51 .INIT = 16'hFCEE;
  X_LUT4 \DLX_EXinst__n0007<10>51  (
    .ADR0(DLX_EXinst__n0079),
    .ADR1(DLX_EXinst_N74245),
    .ADR2(DLX_EXinst__n0077),
    .ADR3(DLX_IDinst_reg_out_B[10]),
    .O(\DLX_IFinst_IR_curr<26>/FROM )
  );
  defparam \DLX_EXinst__n0007<10>12 .INIT = 16'hA0A8;
  X_LUT4 \DLX_EXinst__n0007<10>12  (
    .ADR0(DLX_IDinst_reg_out_B[10]),
    .ADR1(DLX_EXinst__n0079),
    .ADR2(DLX_EXinst__n0078),
    .ADR3(DLX_IDinst_reg_out_A[10]),
    .O(\DLX_IFinst_IR_curr<26>/GROM )
  );
  X_BUF \DLX_IFinst_IR_curr<26>/XUSED  (
    .I(\DLX_IFinst_IR_curr<26>/FROM ),
    .O(CHOICE4459)
  );
  X_BUF \DLX_IFinst_IR_curr<26>/YUSED  (
    .I(\DLX_IFinst_IR_curr<26>/GROM ),
    .O(CHOICE4445)
  );
  defparam DLX_IFinst_IR_curr_18.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_18 (
    .I(IR[18]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[18])
  );
  defparam \DLX_EXinst__n0007<11>25 .INIT = 16'hD080;
  X_LUT4 \DLX_EXinst__n0007<11>25  (
    .ADR0(DLX_IDinst_reg_out_B[2]),
    .ADR1(DLX_EXinst_N74686),
    .ADR2(DLX_EXinst_N76457),
    .ADR3(DLX_EXinst_N74991),
    .O(\DLX_IFinst_IR_curr<18>/FROM )
  );
  defparam \DLX_EXinst__n0007<10>25 .INIT = 16'hE200;
  X_LUT4 \DLX_EXinst__n0007<10>25  (
    .ADR0(DLX_EXinst_N74681),
    .ADR1(DLX_IDinst_reg_out_B[2]),
    .ADR2(DLX_EXinst_N74441),
    .ADR3(DLX_EXinst_N76457),
    .O(\DLX_IFinst_IR_curr<18>/GROM )
  );
  X_BUF \DLX_IFinst_IR_curr<18>/XUSED  (
    .I(\DLX_IFinst_IR_curr<18>/FROM ),
    .O(CHOICE4390)
  );
  X_BUF \DLX_IFinst_IR_curr<18>/YUSED  (
    .I(\DLX_IFinst_IR_curr<18>/GROM ),
    .O(CHOICE4450)
  );
  defparam DLX_IDinst_RegFile_14_7_1445.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_14_7_1445 (
    .I(DLX_MEMinst_RF_data_in[7]),
    .CE(DLX_IDinst__n0578),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_14_7)
  );
  defparam \DLX_EXinst__n0007<11>51 .INIT = 16'hFEF4;
  X_LUT4 \DLX_EXinst__n0007<11>51  (
    .ADR0(DLX_IDinst_reg_out_B[11]),
    .ADR1(DLX_EXinst__n0079),
    .ADR2(DLX_EXinst_N74245),
    .ADR3(DLX_EXinst__n0077),
    .O(\DLX_IDinst_RegFile_14_7/FROM )
  );
  defparam \DLX_EXinst__n0007<11>12 .INIT = 16'hC4C0;
  X_LUT4 \DLX_EXinst__n0007<11>12  (
    .ADR0(DLX_IDinst_reg_out_A[11]),
    .ADR1(DLX_IDinst_reg_out_B[11]),
    .ADR2(DLX_EXinst__n0078),
    .ADR3(DLX_EXinst__n0079),
    .O(\DLX_IDinst_RegFile_14_7/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_14_7/XUSED  (
    .I(\DLX_IDinst_RegFile_14_7/FROM ),
    .O(CHOICE4399)
  );
  X_BUF \DLX_IDinst_RegFile_14_7/YUSED  (
    .I(\DLX_IDinst_RegFile_14_7/GROM ),
    .O(CHOICE4385)
  );
  defparam \DLX_EXinst__n0007<12>62 .INIT = 16'hFFE4;
  X_LUT4 \DLX_EXinst__n0007<12>62  (
    .ADR0(DLX_IDinst_reg_out_B[12]),
    .ADR1(DLX_EXinst__n0079),
    .ADR2(DLX_EXinst__n0077),
    .ADR3(DLX_EXinst_N74245),
    .O(\DLX_IDinst_RegFile_11_20/FROM )
  );
  defparam \DLX_EXinst__n0007<12>13 .INIT = 16'hBA00;
  X_LUT4 \DLX_EXinst__n0007<12>13  (
    .ADR0(DLX_EXinst__n0078),
    .ADR1(DLX_IDinst_reg_out_A[12]),
    .ADR2(DLX_EXinst__n0079),
    .ADR3(DLX_IDinst_reg_out_B[12]),
    .O(\DLX_IDinst_RegFile_11_20/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_11_20/XUSED  (
    .I(\DLX_IDinst_RegFile_11_20/FROM ),
    .O(CHOICE3782)
  );
  X_BUF \DLX_IDinst_RegFile_11_20/YUSED  (
    .I(\DLX_IDinst_RegFile_11_20/GROM ),
    .O(CHOICE3766)
  );
  defparam \DLX_EXinst__n0007<4>207 .INIT = 16'hEECC;
  X_LUT4 \DLX_EXinst__n0007<4>207  (
    .ADR0(DLX_EXinst_N75154),
    .ADR1(DLX_EXinst__n0053),
    .ADR2(VCC),
    .ADR3(N147520),
    .O(\DLX_IDinst_RegFile_11_30/FROM )
  );
  defparam \DLX_EXinst__n0007<20>51 .INIT = 16'hAE0C;
  X_LUT4 \DLX_EXinst__n0007<20>51  (
    .ADR0(DLX_EXinst_N75154),
    .ADR1(N163526),
    .ADR2(N146478),
    .ADR3(N147520),
    .O(\DLX_IDinst_RegFile_11_30/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_11_30/XUSED  (
    .I(\DLX_IDinst_RegFile_11_30/FROM ),
    .O(CHOICE4371)
  );
  X_BUF \DLX_IDinst_RegFile_11_30/YUSED  (
    .I(\DLX_IDinst_RegFile_11_30/GROM ),
    .O(CHOICE4647)
  );
  defparam \DLX_EXinst__n0007<20>29 .INIT = 16'hA280;
  X_LUT4 \DLX_EXinst__n0007<20>29  (
    .ADR0(DLX_EXinst__n0055),
    .ADR1(\DLX_IDinst_Imm[3] ),
    .ADR2(DLX_EXinst_N74223),
    .ADR3(DLX_EXinst_N75377),
    .O(\DLX_IDinst_RegFile_11_15/FROM )
  );
  defparam \DLX_EXinst__n0007<20>51_SW0 .INIT = 16'hFF88;
  X_LUT4 \DLX_EXinst__n0007<20>51_SW0  (
    .ADR0(\DLX_EXinst_Mshift__n0022_Sh[52] ),
    .ADR1(DLX_EXinst__n0056),
    .ADR2(VCC),
    .ADR3(CHOICE4642),
    .O(\DLX_IDinst_RegFile_11_15/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_11_15/XUSED  (
    .I(\DLX_IDinst_RegFile_11_15/FROM ),
    .O(CHOICE4642)
  );
  X_BUF \DLX_IDinst_RegFile_11_15/YUSED  (
    .I(\DLX_IDinst_RegFile_11_15/GROM ),
    .O(N163526)
  );
  defparam \DLX_EXinst__n0007<12>71 .INIT = 16'hECA0;
  X_LUT4 \DLX_EXinst__n0007<12>71  (
    .ADR0(DLX_IDinst_reg_out_A[12]),
    .ADR1(DLX_EXinst_ALU_result[12]),
    .ADR2(CHOICE3782),
    .ADR3(N134884),
    .O(\CHOICE3784/FROM )
  );
  defparam \DLX_EXinst__n0007<12>80 .INIT = 16'hFF32;
  X_LUT4 \DLX_EXinst__n0007<12>80  (
    .ADR0(CHOICE3773),
    .ADR1(DLX_IDinst_reg_out_B[4]),
    .ADR2(CHOICE3774),
    .ADR3(CHOICE3784),
    .O(\CHOICE3784/GROM )
  );
  X_BUF \CHOICE3784/XUSED  (
    .I(\CHOICE3784/FROM ),
    .O(CHOICE3784)
  );
  X_BUF \CHOICE3784/YUSED  (
    .I(\CHOICE3784/GROM ),
    .O(CHOICE3785)
  );
  defparam \DLX_EXinst__n0007<15>39 .INIT = 16'hA030;
  X_LUT4 \DLX_EXinst__n0007<15>39  (
    .ADR0(DLX_EXinst_N72913),
    .ADR1(N130157),
    .ADR2(DLX_EXinst_N76338),
    .ADR3(DLX_IDinst_reg_out_B[3]),
    .O(\DLX_IDinst_RegFile_11_25/FROM )
  );
  defparam \DLX_EXinst__n0007<13>34 .INIT = 16'hD100;
  X_LUT4 \DLX_EXinst__n0007<13>34  (
    .ADR0(N130051),
    .ADR1(DLX_IDinst_reg_out_B[3]),
    .ADR2(DLX_EXinst_N72903),
    .ADR3(DLX_EXinst_N76338),
    .O(\DLX_IDinst_RegFile_11_25/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_11_25/XUSED  (
    .I(\DLX_IDinst_RegFile_11_25/FROM ),
    .O(CHOICE4274)
  );
  X_BUF \DLX_IDinst_RegFile_11_25/YUSED  (
    .I(\DLX_IDinst_RegFile_11_25/GROM ),
    .O(CHOICE3719)
  );
  defparam \DLX_EXinst__n0007<8>113_SW0 .INIT = 16'hEAC0;
  X_LUT4 \DLX_EXinst__n0007<8>113_SW0  (
    .ADR0(CHOICE5139),
    .ADR1(N148609),
    .ADR2(CHOICE5146),
    .ADR3(DLX_IDinst_reg_out_A[8]),
    .O(\N163538/FROM )
  );
  defparam \DLX_EXinst__n0007<8>113 .INIT = 16'hFFEA;
  X_LUT4 \DLX_EXinst__n0007<8>113  (
    .ADR0(CHOICE5154),
    .ADR1(DLX_EXinst_ALU_result[8]),
    .ADR2(N134884),
    .ADR3(N163538),
    .O(\N163538/GROM )
  );
  X_BUF \N163538/XUSED  (
    .I(\N163538/FROM ),
    .O(N163538)
  );
  X_BUF \N163538/YUSED  (
    .I(\N163538/GROM ),
    .O(CHOICE5156)
  );
  defparam \DLX_EXinst__n0007<0>165 .INIT = 16'hFFE4;
  X_LUT4 \DLX_EXinst__n0007<0>165  (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(DLX_EXinst__n0079),
    .ADR2(DLX_EXinst__n0077),
    .ADR3(DLX_EXinst_N74245),
    .O(\DLX_IDinst_RegFile_1_24/FROM )
  );
  defparam \DLX_EXinst__n0007<13>62 .INIT = 16'hFFE4;
  X_LUT4 \DLX_EXinst__n0007<13>62  (
    .ADR0(DLX_IDinst_reg_out_B[13]),
    .ADR1(DLX_EXinst__n0079),
    .ADR2(DLX_EXinst__n0077),
    .ADR3(DLX_EXinst_N74245),
    .O(\DLX_IDinst_RegFile_1_24/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_1_24/XUSED  (
    .I(\DLX_IDinst_RegFile_1_24/FROM ),
    .O(CHOICE5901)
  );
  X_BUF \DLX_IDinst_RegFile_1_24/YUSED  (
    .I(\DLX_IDinst_RegFile_1_24/GROM ),
    .O(CHOICE3727)
  );
  defparam \DLX_EXinst__n0007<13>71 .INIT = 16'hECA0;
  X_LUT4 \DLX_EXinst__n0007<13>71  (
    .ADR0(DLX_EXinst_ALU_result[13]),
    .ADR1(DLX_IDinst_reg_out_A[13]),
    .ADR2(N134884),
    .ADR3(CHOICE3727),
    .O(\CHOICE3729/FROM )
  );
  defparam \DLX_EXinst__n0007<13>80 .INIT = 16'hFF54;
  X_LUT4 \DLX_EXinst__n0007<13>80  (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(CHOICE3718),
    .ADR2(CHOICE3719),
    .ADR3(CHOICE3729),
    .O(\CHOICE3729/GROM )
  );
  X_BUF \CHOICE3729/XUSED  (
    .I(\CHOICE3729/FROM ),
    .O(CHOICE3729)
  );
  X_BUF \CHOICE3729/YUSED  (
    .I(\CHOICE3729/GROM ),
    .O(CHOICE3730)
  );
  defparam DLX_EXinst_Ker729011.INIT = 16'hB8B8;
  X_LUT4 DLX_EXinst_Ker729011 (
    .ADR0(\DLX_EXinst_Mshift__n0023_Sh[1] ),
    .ADR1(DLX_IDinst_reg_out_B[2]),
    .ADR2(\DLX_EXinst_Mshift__n0023_Sh[5] ),
    .ADR3(VCC),
    .O(\DLX_IDinst_RegFile_23_3/FROM )
  );
  defparam \DLX_EXinst__n0007<14>33 .INIT = 16'hAC00;
  X_LUT4 \DLX_EXinst__n0007<14>33  (
    .ADR0(DLX_EXinst_N74731),
    .ADR1(DLX_EXinst_N74441),
    .ADR2(DLX_IDinst_reg_out_B[2]),
    .ADR3(DLX_EXinst_N72710),
    .O(\DLX_IDinst_RegFile_23_3/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_23_3/XUSED  (
    .I(\DLX_IDinst_RegFile_23_3/FROM ),
    .O(DLX_EXinst_N72903)
  );
  X_BUF \DLX_IDinst_RegFile_23_3/YUSED  (
    .I(\DLX_IDinst_RegFile_23_3/GROM ),
    .O(CHOICE3663)
  );
  defparam DLX_EXinst_Ker73851.INIT = 16'hCCF0;
  X_LUT4 DLX_EXinst_Ker73851 (
    .ADR0(VCC),
    .ADR1(\DLX_EXinst_Mshift__n0023_Sh[10] ),
    .ADR2(N130001),
    .ADR3(DLX_IDinst_reg_out_B[3]),
    .O(\DLX_IDinst_RegFile_14_8/FROM )
  );
  defparam \DLX_EXinst__n0007<14>34 .INIT = 16'h808A;
  X_LUT4 \DLX_EXinst__n0007<14>34  (
    .ADR0(DLX_EXinst_N76338),
    .ADR1(DLX_EXinst_N72908),
    .ADR2(DLX_IDinst_reg_out_B[3]),
    .ADR3(N130105),
    .O(\DLX_IDinst_RegFile_14_8/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_14_8/XUSED  (
    .I(\DLX_IDinst_RegFile_14_8/FROM ),
    .O(DLX_EXinst_N73853)
  );
  X_BUF \DLX_IDinst_RegFile_14_8/YUSED  (
    .I(\DLX_IDinst_RegFile_14_8/GROM ),
    .O(CHOICE3664)
  );
  defparam \DLX_EXinst__n0007<27>21 .INIT = 16'hECA0;
  X_LUT4 \DLX_EXinst__n0007<27>21  (
    .ADR0(DLX_EXinst__n0012[27]),
    .ADR1(\DLX_IDinst_Imm[11] ),
    .ADR2(DLX_EXinst__n0109),
    .ADR3(DLX_EXinst__n0051),
    .O(\DLX_IDinst_RegFile_3_2/FROM )
  );
  defparam \DLX_EXinst__n0007<22>70 .INIT = 16'hECA0;
  X_LUT4 \DLX_EXinst__n0007<22>70  (
    .ADR0(DLX_EXinst__n0012[22]),
    .ADR1(DLX_EXinst__n0051),
    .ADR2(DLX_EXinst__n0109),
    .ADR3(\DLX_IDinst_Imm[6] ),
    .O(\DLX_IDinst_RegFile_3_2/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_3_2/XUSED  (
    .I(\DLX_IDinst_RegFile_3_2/FROM ),
    .O(CHOICE4929)
  );
  X_BUF \DLX_IDinst_RegFile_3_2/YUSED  (
    .I(\DLX_IDinst_RegFile_3_2/GROM ),
    .O(CHOICE4075)
  );
  defparam \DLX_EXinst__n0007<3>165 .INIT = 16'hA0A8;
  X_LUT4 \DLX_EXinst__n0007<3>165  (
    .ADR0(DLX_IDinst_reg_out_B[3]),
    .ADR1(DLX_EXinst__n0079),
    .ADR2(DLX_EXinst__n0078),
    .ADR3(DLX_IDinst_reg_out_A[3]),
    .O(\DLX_IDinst_RegFile_3_3/FROM )
  );
  defparam \DLX_EXinst__n0007<14>62 .INIT = 16'hFCFA;
  X_LUT4 \DLX_EXinst__n0007<14>62  (
    .ADR0(DLX_EXinst__n0079),
    .ADR1(DLX_EXinst__n0077),
    .ADR2(DLX_EXinst_N74245),
    .ADR3(DLX_IDinst_reg_out_B[14]),
    .O(\DLX_IDinst_RegFile_3_3/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_3_3/XUSED  (
    .I(\DLX_IDinst_RegFile_3_3/FROM ),
    .O(CHOICE5469)
  );
  X_BUF \DLX_IDinst_RegFile_3_3/YUSED  (
    .I(\DLX_IDinst_RegFile_3_3/GROM ),
    .O(CHOICE3672)
  );
  defparam DLX_IDinst_RegFile_27_16_1446.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_27_16_1446 (
    .I(DLX_IDinst_WB_data_eff[16]),
    .CE(DLX_IDinst__n0604),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_27_16)
  );
  defparam \DLX_EXinst__n0007<14>71 .INIT = 16'hF888;
  X_LUT4 \DLX_EXinst__n0007<14>71  (
    .ADR0(DLX_EXinst_ALU_result[14]),
    .ADR1(N134884),
    .ADR2(CHOICE3672),
    .ADR3(DLX_IDinst_reg_out_A[14]),
    .O(\CHOICE3674/FROM )
  );
  defparam \DLX_EXinst__n0007<14>80 .INIT = 16'hFF54;
  X_LUT4 \DLX_EXinst__n0007<14>80  (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(CHOICE3663),
    .ADR2(CHOICE3664),
    .ADR3(CHOICE3674),
    .O(\CHOICE3674/GROM )
  );
  X_BUF \CHOICE3674/XUSED  (
    .I(\CHOICE3674/FROM ),
    .O(CHOICE3674)
  );
  X_BUF \CHOICE3674/YUSED  (
    .I(\CHOICE3674/GROM ),
    .O(CHOICE3675)
  );
  defparam \DLX_EXinst__n0007<25>21 .INIT = 16'hEAC0;
  X_LUT4 \DLX_EXinst__n0007<25>21  (
    .ADR0(DLX_EXinst__n0051),
    .ADR1(DLX_EXinst__n0012[25]),
    .ADR2(DLX_EXinst__n0109),
    .ADR3(\DLX_IDinst_Imm[9] ),
    .O(\DLX_IDinst_RegFile_22_9/FROM )
  );
  defparam \DLX_EXinst__n0007<23>70 .INIT = 16'hF888;
  X_LUT4 \DLX_EXinst__n0007<23>70  (
    .ADR0(\DLX_IDinst_Imm[7] ),
    .ADR1(DLX_EXinst__n0051),
    .ADR2(DLX_EXinst__n0109),
    .ADR3(DLX_EXinst__n0012[23]),
    .O(\DLX_IDinst_RegFile_22_9/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_22_9/XUSED  (
    .I(\DLX_IDinst_RegFile_22_9/FROM ),
    .O(CHOICE5063)
  );
  X_BUF \DLX_IDinst_RegFile_22_9/YUSED  (
    .I(\DLX_IDinst_RegFile_22_9/GROM ),
    .O(CHOICE4010)
  );
  defparam \DLX_EXinst__n0007<2>165 .INIT = 16'hC4C0;
  X_LUT4 \DLX_EXinst__n0007<2>165  (
    .ADR0(DLX_IDinst_reg_out_A[2]),
    .ADR1(DLX_IDinst_reg_out_B[2]),
    .ADR2(DLX_EXinst__n0078),
    .ADR3(DLX_EXinst__n0079),
    .O(\DLX_IDinst_RegFile_7_5/FROM )
  );
  defparam \DLX_EXinst__n0007<0>207 .INIT = 16'h88A8;
  X_LUT4 \DLX_EXinst__n0007<0>207  (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(DLX_EXinst__n0078),
    .ADR2(DLX_EXinst__n0079),
    .ADR3(DLX_IDinst_reg_out_A[0]),
    .O(\DLX_IDinst_RegFile_7_5/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_7_5/XUSED  (
    .I(\DLX_IDinst_RegFile_7_5/FROM ),
    .O(CHOICE5545)
  );
  X_BUF \DLX_IDinst_RegFile_7_5/YUSED  (
    .I(\DLX_IDinst_RegFile_7_5/GROM ),
    .O(CHOICE5908)
  );
  defparam DLX_IDinst_RegFile_27_24_1447.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_27_24_1447 (
    .I(DLX_IDinst_WB_data_eff[24]),
    .CE(DLX_IDinst__n0604),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_27_24)
  );
  defparam DLX_EXinst_Ker7551825.INIT = 16'h2028;
  X_LUT4 DLX_EXinst_Ker7551825 (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(DLX_IDinst_reg_out_B[5]),
    .ADR2(DLX_EXinst_N72822),
    .ADR3(DLX_IDinst_reg_out_B[1]),
    .O(\DLX_IDinst_RegFile_2_8/FROM )
  );
  defparam \DLX_EXinst__n0007<0>208 .INIT = 16'h8800;
  X_LUT4 \DLX_EXinst__n0007<0>208  (
    .ADR0(DLX_IDinst_reg_out_B[5]),
    .ADR1(N148609),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[31]),
    .O(\DLX_IDinst_RegFile_2_8/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_2_8/XUSED  (
    .I(\DLX_IDinst_RegFile_2_8/FROM ),
    .O(CHOICE2049)
  );
  X_BUF \DLX_IDinst_RegFile_2_8/YUSED  (
    .I(\DLX_IDinst_RegFile_2_8/GROM ),
    .O(CHOICE5909)
  );
  defparam DLX_EXinst_Ker759711.INIT = 16'h2200;
  X_LUT4 DLX_EXinst_Ker759711 (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(N148323),
    .ADR2(VCC),
    .ADR3(DLX_EXinst__n0080),
    .O(\DLX_IDinst_RegFile_23_7/FROM )
  );
  defparam \DLX_EXinst__n0007<0>225 .INIT = 16'h0040;
  X_LUT4 \DLX_EXinst__n0007<0>225  (
    .ADR0(DLX_EXinst_N72822),
    .ADR1(DLX_EXinst_N76268),
    .ADR2(\DLX_EXinst_Mshift__n0023_Sh[0] ),
    .ADR3(N148323),
    .O(\DLX_IDinst_RegFile_23_7/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_23_7/XUSED  (
    .I(\DLX_IDinst_RegFile_23_7/FROM ),
    .O(DLX_EXinst_N75973)
  );
  X_BUF \DLX_IDinst_RegFile_23_7/YUSED  (
    .I(\DLX_IDinst_RegFile_23_7/GROM ),
    .O(CHOICE5915)
  );
  defparam \DLX_EXinst__n0007<15>67 .INIT = 16'hEFEA;
  X_LUT4 \DLX_EXinst__n0007<15>67  (
    .ADR0(DLX_EXinst_N74245),
    .ADR1(DLX_EXinst__n0077),
    .ADR2(DLX_IDinst_reg_out_B[15]),
    .ADR3(DLX_EXinst__n0079),
    .O(\CHOICE4282/FROM )
  );
  defparam \DLX_EXinst__n0007<15>76 .INIT = 16'hEAC0;
  X_LUT4 \DLX_EXinst__n0007<15>76  (
    .ADR0(DLX_IDinst_reg_out_A[15]),
    .ADR1(DLX_EXinst_ALU_result[15]),
    .ADR2(N134884),
    .ADR3(CHOICE4282),
    .O(\CHOICE4282/GROM )
  );
  X_BUF \CHOICE4282/XUSED  (
    .I(\CHOICE4282/FROM ),
    .O(CHOICE4282)
  );
  X_BUF \CHOICE4282/YUSED  (
    .I(\CHOICE4282/GROM ),
    .O(CHOICE4284)
  );
  defparam \DLX_EXinst__n0007<15>85 .INIT = 16'hFF0E;
  X_LUT4 \DLX_EXinst__n0007<15>85  (
    .ADR0(CHOICE4274),
    .ADR1(CHOICE4273),
    .ADR2(DLX_IDinst_reg_out_B[4]),
    .ADR3(CHOICE4284),
    .O(\CHOICE4285/FROM )
  );
  defparam \DLX_EXinst__n0007<15>110 .INIT = 16'hAAA8;
  X_LUT4 \DLX_EXinst__n0007<15>110  (
    .ADR0(DLX_EXinst__n0036),
    .ADR1(CHOICE4266),
    .ADR2(CHOICE4263),
    .ADR3(CHOICE4285),
    .O(\CHOICE4285/GROM )
  );
  X_BUF \CHOICE4285/XUSED  (
    .I(\CHOICE4285/FROM ),
    .O(CHOICE4285)
  );
  X_BUF \CHOICE4285/YUSED  (
    .I(\CHOICE4285/GROM ),
    .O(CHOICE4287)
  );
  defparam DLX_EXinst_Ker7445415.INIT = 16'h0C0A;
  X_LUT4 DLX_EXinst_Ker7445415 (
    .ADR0(\DLX_EXinst_Mshift__n0019_Sh[27] ),
    .ADR1(DLX_IDinst_reg_out_A[31]),
    .ADR2(DLX_IDinst_reg_out_B_2_1),
    .ADR3(DLX_IDinst_reg_out_B[5]),
    .O(\DLX_IDinst_RegFile_27_23/FROM )
  );
  defparam \DLX_EXinst__n0007<24>45 .INIT = 16'h22B8;
  X_LUT4 \DLX_EXinst__n0007<24>45  (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(N163790),
    .ADR2(DLX_EXinst_N73369),
    .ADR3(DLX_IDinst_reg_out_B[5]),
    .O(\DLX_IDinst_RegFile_27_23/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_27_23/XUSED  (
    .I(\DLX_IDinst_RegFile_27_23/FROM ),
    .O(CHOICE1830)
  );
  X_BUF \DLX_IDinst_RegFile_27_23/YUSED  (
    .I(\DLX_IDinst_RegFile_27_23/GROM ),
    .O(CHOICE5598)
  );
  defparam \DLX_EXinst__n0007<0>335 .INIT = 16'h4000;
  X_LUT4 \DLX_EXinst__n0007<0>335  (
    .ADR0(\DLX_IDinst_Imm[4] ),
    .ADR1(\DLX_IDinst_Imm[3] ),
    .ADR2(CHOICE5939),
    .ADR3(DLX_IDinst_IR_function_field[5]),
    .O(\DLX_IDinst_RegFile_3_5/FROM )
  );
  defparam \DLX_EXinst__n0007<0>390_SW0_SW0 .INIT = 16'hFFEE;
  X_LUT4 \DLX_EXinst__n0007<0>390_SW0_SW0  (
    .ADR0(CHOICE5909),
    .ADR1(CHOICE5915),
    .ADR2(VCC),
    .ADR3(CHOICE5941),
    .O(\DLX_IDinst_RegFile_3_5/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_3_5/XUSED  (
    .I(\DLX_IDinst_RegFile_3_5/FROM ),
    .O(CHOICE5941)
  );
  X_BUF \DLX_IDinst_RegFile_3_5/YUSED  (
    .I(\DLX_IDinst_RegFile_3_5/GROM ),
    .O(N164591)
  );
  defparam \DLX_EXinst__n0007<18>27 .INIT = 16'hEAC0;
  X_LUT4 \DLX_EXinst__n0007<18>27  (
    .ADR0(DLX_EXinst__n0109),
    .ADR1(DLX_EXinst__n0051),
    .ADR2(\DLX_IDinst_Imm[2] ),
    .ADR3(DLX_EXinst__n0012[18]),
    .O(\DLX_IFinst_IR_previous<11>/FROM )
  );
  defparam \DLX_EXinst__n0007<17>27 .INIT = 16'hF888;
  X_LUT4 \DLX_EXinst__n0007<17>27  (
    .ADR0(DLX_EXinst__n0012[17]),
    .ADR1(DLX_EXinst__n0109),
    .ADR2(DLX_EXinst__n0051),
    .ADR3(\DLX_IDinst_Imm[1] ),
    .O(\DLX_IFinst_IR_previous<11>/GROM )
  );
  X_BUF \DLX_IFinst_IR_previous<11>/XUSED  (
    .I(\DLX_IFinst_IR_previous<11>/FROM ),
    .O(CHOICE5203)
  );
  X_BUF \DLX_IFinst_IR_previous<11>/YUSED  (
    .I(\DLX_IFinst_IR_previous<11>/GROM ),
    .O(CHOICE5361)
  );
  defparam \DLX_EXinst__n0007<1>221 .INIT = 16'hFDEC;
  X_LUT4 \DLX_EXinst__n0007<1>221  (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(DLX_EXinst_N74245),
    .ADR2(DLX_EXinst__n0077),
    .ADR3(DLX_EXinst__n0079),
    .O(\CHOICE5741/FROM )
  );
  defparam \DLX_EXinst__n0007<1>261_SW0 .INIT = 16'hF888;
  X_LUT4 \DLX_EXinst__n0007<1>261_SW0  (
    .ADR0(N137859),
    .ADR1(DLX_EXinst_N75983),
    .ADR2(CHOICE5741),
    .ADR3(DLX_IDinst_reg_out_A[1]),
    .O(\CHOICE5741/GROM )
  );
  X_BUF \CHOICE5741/XUSED  (
    .I(\CHOICE5741/FROM ),
    .O(CHOICE5741)
  );
  X_BUF \CHOICE5741/YUSED  (
    .I(\CHOICE5741/GROM ),
    .O(N163648)
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<24>1 .INIT = 16'hE4E4;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<24>1  (
    .ADR0(DLX_EXinst_mem_to_reg_EX),
    .ADR1(DLX_EXinst_ALU_result[24]),
    .ADR2(DM_read_data[24]),
    .ADR3(VCC),
    .O(DLX_MEMinst__n0000[24])
  );
  defparam \DLX_EXinst__n0007<24>85 .INIT = 16'hECA0;
  X_LUT4 \DLX_EXinst__n0007<24>85  (
    .ADR0(DLX_EXinst__n0012[24]),
    .ADR1(DLX_EXinst_ALU_result[24]),
    .ADR2(DLX_EXinst__n0127),
    .ADR3(N134884),
    .O(\DLX_MEMinst_RF_data_in<24>/GROM )
  );
  X_BUF \DLX_MEMinst_RF_data_in<24>/YUSED  (
    .I(\DLX_MEMinst_RF_data_in<24>/GROM ),
    .O(CHOICE5603)
  );
  defparam \DLX_EXinst__n0007<0>471 .INIT = 16'h0503;
  X_LUT4 \DLX_EXinst__n0007<0>471  (
    .ADR0(N164614),
    .ADR1(N164612),
    .ADR2(DLX_IDinst_IR_opcode_field[2]),
    .ADR3(DLX_IDinst_IR_opcode_field[0]),
    .O(\CHOICE5967/FROM )
  );
  defparam \DLX_EXinst__n0007<0>477 .INIT = 16'hFF54;
  X_LUT4 \DLX_EXinst__n0007<0>477  (
    .ADR0(DLX_IDinst_IR_opcode_field[1]),
    .ADR1(CHOICE5952),
    .ADR2(CHOICE5958),
    .ADR3(CHOICE5967),
    .O(\CHOICE5967/GROM )
  );
  X_BUF \CHOICE5967/XUSED  (
    .I(\CHOICE5967/FROM ),
    .O(CHOICE5967)
  );
  X_BUF \CHOICE5967/YUSED  (
    .I(\CHOICE5967/GROM ),
    .O(CHOICE5968)
  );
  defparam \DLX_EXinst__n0007<24>96 .INIT = 16'hFBEA;
  X_LUT4 \DLX_EXinst__n0007<24>96  (
    .ADR0(DLX_EXinst_N74245),
    .ADR1(DLX_IDinst_reg_out_B[24]),
    .ADR2(DLX_EXinst__n0077),
    .ADR3(DLX_EXinst__n0079),
    .O(\DLX_IDinst_RegFile_2_9/FROM )
  );
  defparam \DLX_EXinst__n0007<24>206 .INIT = 16'hFCCC;
  X_LUT4 \DLX_EXinst__n0007<24>206  (
    .ADR0(VCC),
    .ADR1(CHOICE5630),
    .ADR2(DLX_IDinst_reg_out_A[24]),
    .ADR3(CHOICE5608),
    .O(\DLX_IDinst_RegFile_2_9/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_2_9/XUSED  (
    .I(\DLX_IDinst_RegFile_2_9/FROM ),
    .O(CHOICE5608)
  );
  X_BUF \DLX_IDinst_RegFile_2_9/YUSED  (
    .I(\DLX_IDinst_RegFile_2_9/GROM ),
    .O(CHOICE5631)
  );
  defparam \DLX_EXinst__n0007<17>136_SW0 .INIT = 16'h0A28;
  X_LUT4 \DLX_EXinst__n0007<17>136_SW0  (
    .ADR0(DLX_EXinst_N76011),
    .ADR1(DLX_IDinst_reg_out_A[17]),
    .ADR2(DLX_IDinst_IR_opcode_field[1]),
    .ADR3(DLX_IDinst_IR_opcode_field[0]),
    .O(\DLX_IFinst_IR_previous<23>/FROM )
  );
  defparam \DLX_EXinst__n0007<0>529 .INIT = 16'h0A28;
  X_LUT4 \DLX_EXinst__n0007<0>529  (
    .ADR0(DLX_EXinst_N76011),
    .ADR1(DLX_IDinst_IR_opcode_field[0]),
    .ADR2(DLX_IDinst_IR_opcode_field[1]),
    .ADR3(DLX_IDinst_reg_out_A[0]),
    .O(\DLX_IFinst_IR_previous<23>/GROM )
  );
  X_BUF \DLX_IFinst_IR_previous<23>/XUSED  (
    .I(\DLX_IFinst_IR_previous<23>/FROM ),
    .O(N163631)
  );
  X_BUF \DLX_IFinst_IR_previous<23>/YUSED  (
    .I(\DLX_IFinst_IR_previous<23>/GROM ),
    .O(CHOICE5976)
  );
  defparam DLX_IDinst_RegFile_10_1_1448.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_10_1_1448 (
    .I(DLX_MEMinst_RF_data_in[1]),
    .CE(DLX_IDinst__n0570),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_10_1)
  );
  defparam \DLX_EXinst__n0007<3>234 .INIT = 16'hD080;
  X_LUT4 \DLX_EXinst__n0007<3>234  (
    .ADR0(DLX_IDinst_reg_out_B[2]),
    .ADR1(DLX_EXinst_N73103),
    .ADR2(DLX_EXinst_N76431),
    .ADR3(DLX_EXinst_N74976),
    .O(\DLX_IDinst_RegFile_10_1/FROM )
  );
  defparam \DLX_EXinst__n0007<1>234 .INIT = 16'hD080;
  X_LUT4 \DLX_EXinst__n0007<1>234  (
    .ADR0(DLX_IDinst_reg_out_B[2]),
    .ADR1(DLX_EXinst_N73093),
    .ADR2(DLX_EXinst_N76431),
    .ADR3(DLX_EXinst_N74726),
    .O(\DLX_IDinst_RegFile_10_1/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_10_1/XUSED  (
    .I(\DLX_IDinst_RegFile_10_1/FROM ),
    .O(CHOICE5492)
  );
  X_BUF \DLX_IDinst_RegFile_10_1/YUSED  (
    .I(\DLX_IDinst_RegFile_10_1/GROM ),
    .O(CHOICE5747)
  );
  defparam DLX_EXinst_Ker7618111.INIT = 16'h4000;
  X_LUT4 DLX_EXinst_Ker7618111 (
    .ADR0(DLX_IDinst_IR_function_field[5]),
    .ADR1(DLX_IDinst_Imm_1_1),
    .ADR2(\DLX_IDinst_Imm[0] ),
    .ADR3(DLX_EXinst_N76002),
    .O(\DLX_IDinst_RegFile_10_2/FROM )
  );
  defparam \DLX_EXinst__n0007<0>538 .INIT = 16'hECA0;
  X_LUT4 \DLX_EXinst__n0007<0>538  (
    .ADR0(CHOICE5976),
    .ADR1(DLX_EXinst__n0109),
    .ADR2(\DLX_IDinst_Imm[0] ),
    .ADR3(DLX_EXinst__n0012[0]),
    .O(\DLX_IDinst_RegFile_10_2/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_10_2/XUSED  (
    .I(\DLX_IDinst_RegFile_10_2/FROM ),
    .O(CHOICE3600)
  );
  X_BUF \DLX_IDinst_RegFile_10_2/YUSED  (
    .I(\DLX_IDinst_RegFile_10_2/GROM ),
    .O(CHOICE5978)
  );
  defparam \DLX_EXinst__n0007<25>75 .INIT = 16'h8F88;
  X_LUT4 \DLX_EXinst__n0007<25>75  (
    .ADR0(N147520),
    .ADR1(N138481),
    .ADR2(N146478),
    .ADR3(N163610),
    .O(\CHOICE5081/FROM )
  );
  defparam \DLX_EXinst__n0007<25>97 .INIT = 16'hB3A0;
  X_LUT4 \DLX_EXinst__n0007<25>97  (
    .ADR0(N163606),
    .ADR1(\DLX_IDinst_Imm[4] ),
    .ADR2(\DLX_IDinst_Imm[31] ),
    .ADR3(CHOICE5081),
    .O(\CHOICE5081/GROM )
  );
  X_BUF \CHOICE5081/XUSED  (
    .I(\CHOICE5081/FROM ),
    .O(CHOICE5081)
  );
  X_BUF \CHOICE5081/YUSED  (
    .I(\CHOICE5081/GROM ),
    .O(CHOICE5083)
  );
  defparam \DLX_EXinst__n0007<0>299 .INIT = 16'h0503;
  X_LUT4 \DLX_EXinst__n0007<0>299  (
    .ADR0(N164620),
    .ADR1(N164618),
    .ADR2(\DLX_IDinst_Imm[2] ),
    .ADR3(\DLX_IDinst_Imm[0] ),
    .O(\CHOICE5938/FROM )
  );
  defparam \DLX_EXinst__n0007<0>305 .INIT = 16'hFF0E;
  X_LUT4 \DLX_EXinst__n0007<0>305  (
    .ADR0(CHOICE5929),
    .ADR1(CHOICE5923),
    .ADR2(\DLX_IDinst_Imm[1] ),
    .ADR3(CHOICE5938),
    .O(\CHOICE5938/GROM )
  );
  X_BUF \CHOICE5938/XUSED  (
    .I(\CHOICE5938/FROM ),
    .O(CHOICE5938)
  );
  X_BUF \CHOICE5938/YUSED  (
    .I(\CHOICE5938/GROM ),
    .O(CHOICE5939)
  );
  defparam DLX_EXinst_Ker746941.INIT = 16'hEE44;
  X_LUT4 DLX_EXinst_Ker746941 (
    .ADR0(DLX_IDinst_reg_out_B_3_1),
    .ADR1(\DLX_EXinst_Mshift__n0019_Sh[9] ),
    .ADR2(VCC),
    .ADR3(\DLX_EXinst_Mshift__n0019_Sh[17] ),
    .O(\DLX_IDinst_RegFile_10_4/FROM )
  );
  defparam \DLX_EXinst__n0007<1>172 .INIT = 16'hCC50;
  X_LUT4 \DLX_EXinst__n0007<1>172  (
    .ADR0(DLX_EXinst_N73239),
    .ADR1(\DLX_EXinst_Mshift__n0019_Sh[9] ),
    .ADR2(DLX_IDinst_reg_out_A[1]),
    .ADR3(DLX_IDinst_reg_out_B[3]),
    .O(\DLX_IDinst_RegFile_10_4/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_10_4/XUSED  (
    .I(\DLX_IDinst_RegFile_10_4/FROM ),
    .O(DLX_EXinst_N74696)
  );
  X_BUF \DLX_IDinst_RegFile_10_4/YUSED  (
    .I(\DLX_IDinst_RegFile_10_4/GROM ),
    .O(CHOICE5729)
  );
  defparam \DLX_EXinst__n0007<0>708 .INIT = 16'h88C8;
  X_LUT4 \DLX_EXinst__n0007<0>708  (
    .ADR0(DLX_EXinst__n0053),
    .ADR1(DLX_IDinst_reg_out_A[0]),
    .ADR2(DLX_EXinst__n0054),
    .ADR3(\DLX_IDinst_Imm[0] ),
    .O(\CHOICE6008/FROM )
  );
  defparam \DLX_EXinst__n0007<0>712 .INIT = 16'hFF54;
  X_LUT4 \DLX_EXinst__n0007<0>712  (
    .ADR0(\DLX_IDinst_Imm[4] ),
    .ADR1(CHOICE5999),
    .ADR2(CHOICE6002),
    .ADR3(CHOICE6008),
    .O(\CHOICE6008/GROM )
  );
  X_BUF \CHOICE6008/XUSED  (
    .I(\CHOICE6008/FROM ),
    .O(CHOICE6008)
  );
  X_BUF \CHOICE6008/YUSED  (
    .I(\CHOICE6008/GROM ),
    .O(CHOICE6009)
  );
  defparam \DLX_EXinst__n0007<1>261 .INIT = 16'hFEFC;
  X_LUT4 \DLX_EXinst__n0007<1>261  (
    .ADR0(DLX_EXinst_ALU_result[1]),
    .ADR1(N163648),
    .ADR2(CHOICE5749),
    .ADR3(N134884),
    .O(\CHOICE5751/FROM )
  );
  defparam \DLX_EXinst__n0007<1>3321_SW0_SW0 .INIT = 16'hAAA8;
  X_LUT4 \DLX_EXinst__n0007<1>3321_SW0_SW0  (
    .ADR0(DLX_EXinst__n0036),
    .ADR1(CHOICE5732),
    .ADR2(CHOICE5724),
    .ADR3(CHOICE5751),
    .O(\CHOICE5751/GROM )
  );
  X_BUF \CHOICE5751/XUSED  (
    .I(\CHOICE5751/FROM ),
    .O(CHOICE5751)
  );
  X_BUF \CHOICE5751/YUSED  (
    .I(\CHOICE5751/GROM ),
    .O(N164573)
  );
  defparam \DLX_EXinst__n0007<0>581 .INIT = 16'h8D88;
  X_LUT4 \DLX_EXinst__n0007<0>581  (
    .ADR0(\DLX_IDinst_Imm[0] ),
    .ADR1(N164636),
    .ADR2(\DLX_IDinst_Imm[1] ),
    .ADR3(DLX_IDinst_reg_out_A[0]),
    .O(\DLX_IDinst_RegFile_10_5/FROM )
  );
  defparam \DLX_EXinst__n0007<0>590 .INIT = 16'hFF20;
  X_LUT4 \DLX_EXinst__n0007<0>590  (
    .ADR0(DLX_IDinst_reg_out_A[2]),
    .ADR1(\DLX_IDinst_Imm[0] ),
    .ADR2(\DLX_IDinst_Imm[1] ),
    .ADR3(CHOICE5993),
    .O(\DLX_IDinst_RegFile_10_5/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_10_5/XUSED  (
    .I(\DLX_IDinst_RegFile_10_5/FROM ),
    .O(CHOICE5993)
  );
  X_BUF \DLX_IDinst_RegFile_10_5/YUSED  (
    .I(\DLX_IDinst_RegFile_10_5/GROM ),
    .O(CHOICE5994)
  );
  defparam \DLX_EXinst__n0007<3>318 .INIT = 16'hECA0;
  X_LUT4 \DLX_EXinst__n0007<3>318  (
    .ADR0(DLX_IDinst_reg_out_A[5]),
    .ADR1(DLX_IDinst_reg_out_A[6]),
    .ADR2(DLX_EXinst_N74347),
    .ADR3(DLX_EXinst_N74625),
    .O(\DLX_IDinst_RegFile_11_1/FROM )
  );
  defparam \DLX_EXinst__n0007<1>318 .INIT = 16'hF888;
  X_LUT4 \DLX_EXinst__n0007<1>318  (
    .ADR0(DLX_EXinst_N74347),
    .ADR1(DLX_IDinst_reg_out_A[3]),
    .ADR2(DLX_IDinst_reg_out_A[4]),
    .ADR3(DLX_EXinst_N74625),
    .O(\DLX_IDinst_RegFile_11_1/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_11_1/XUSED  (
    .I(\DLX_IDinst_RegFile_11_1/FROM ),
    .O(CHOICE5503)
  );
  X_BUF \DLX_IDinst_RegFile_11_1/YUSED  (
    .I(\DLX_IDinst_RegFile_11_1/GROM ),
    .O(CHOICE5758)
  );
  defparam \DLX_EXinst__n0007<6>143 .INIT = 16'hF888;
  X_LUT4 \DLX_EXinst__n0007<6>143  (
    .ADR0(N144481),
    .ADR1(\DLX_IDinst_Imm[4] ),
    .ADR2(CHOICE3910),
    .ADR3(\DLX_IDinst_Imm[6] ),
    .O(\DLX_IFinst_IR_previous<28>/FROM )
  );
  defparam \DLX_EXinst__n0007<0>728 .INIT = 16'hEAAA;
  X_LUT4 \DLX_EXinst__n0007<0>728  (
    .ADR0(N163953),
    .ADR1(DLX_EXinst_N73267),
    .ADR2(\DLX_EXinst_Mshift__n0020_Sh[80] ),
    .ADR3(\DLX_IDinst_Imm[4] ),
    .O(\DLX_IFinst_IR_previous<28>/GROM )
  );
  X_BUF \DLX_IFinst_IR_previous<28>/XUSED  (
    .I(\DLX_IFinst_IR_previous<28>/FROM ),
    .O(CHOICE3912)
  );
  X_BUF \DLX_IFinst_IR_previous<28>/YUSED  (
    .I(\DLX_IFinst_IR_previous<28>/GROM ),
    .O(CHOICE6013)
  );
  defparam \DLX_EXinst__n0007<26>84 .INIT = 16'h00CC;
  X_LUT4 \DLX_EXinst__n0007<26>84  (
    .ADR0(VCC),
    .ADR1(CHOICE5014),
    .ADR2(VCC),
    .ADR3(\DLX_IDinst_Imm[4] ),
    .O(\DLX_IFinst_IR_previous<29>/FROM )
  );
  defparam \DLX_EXinst__n0007<26>110 .INIT = 16'hFFEA;
  X_LUT4 \DLX_EXinst__n0007<26>110  (
    .ADR0(N163242),
    .ADR1(DLX_EXinst__n0012[26]),
    .ADR2(DLX_EXinst__n0109),
    .ADR3(CHOICE5015),
    .O(\DLX_IFinst_IR_previous<29>/GROM )
  );
  X_BUF \DLX_IFinst_IR_previous<29>/XUSED  (
    .I(\DLX_IFinst_IR_previous<29>/FROM ),
    .O(CHOICE5015)
  );
  X_BUF \DLX_IFinst_IR_previous<29>/YUSED  (
    .I(\DLX_IFinst_IR_previous<29>/GROM ),
    .O(CHOICE5017)
  );
  defparam \DLX_EXinst__n0007<2>221 .INIT = 16'hFBEA;
  X_LUT4 \DLX_EXinst__n0007<2>221  (
    .ADR0(DLX_EXinst_N74245),
    .ADR1(DLX_IDinst_reg_out_B[2]),
    .ADR2(DLX_EXinst__n0077),
    .ADR3(DLX_EXinst__n0079),
    .O(\CHOICE5562/FROM )
  );
  defparam \DLX_EXinst__n0007<2>261_SW0 .INIT = 16'hF888;
  X_LUT4 \DLX_EXinst__n0007<2>261_SW0  (
    .ADR0(DLX_EXinst_N75983),
    .ADR1(N137372),
    .ADR2(DLX_IDinst_reg_out_A[2]),
    .ADR3(CHOICE5562),
    .O(\CHOICE5562/GROM )
  );
  X_BUF \CHOICE5562/XUSED  (
    .I(\CHOICE5562/FROM ),
    .O(CHOICE5562)
  );
  X_BUF \CHOICE5562/YUSED  (
    .I(\CHOICE5562/GROM ),
    .O(N163394)
  );
  defparam \DLX_EXinst__n0007<27>75 .INIT = 16'hC0EA;
  X_LUT4 \DLX_EXinst__n0007<27>75  (
    .ADR0(N163530),
    .ADR1(N137774),
    .ADR2(N147520),
    .ADR3(N146478),
    .O(\CHOICE4947/FROM )
  );
  defparam \DLX_EXinst__n0007<27>97 .INIT = 16'hD5C0;
  X_LUT4 \DLX_EXinst__n0007<27>97  (
    .ADR0(\DLX_IDinst_Imm[4] ),
    .ADR1(\DLX_IDinst_Imm[31] ),
    .ADR2(N163518),
    .ADR3(CHOICE4947),
    .O(\CHOICE4947/GROM )
  );
  X_BUF \CHOICE4947/XUSED  (
    .I(\CHOICE4947/FROM ),
    .O(CHOICE4947)
  );
  X_BUF \CHOICE4947/YUSED  (
    .I(\CHOICE4947/GROM ),
    .O(CHOICE4949)
  );
  defparam \DLX_EXinst__n0007<2>261 .INIT = 16'hFFEA;
  X_LUT4 \DLX_EXinst__n0007<2>261  (
    .ADR0(N163394),
    .ADR1(DLX_EXinst_ALU_result[2]),
    .ADR2(N134884),
    .ADR3(CHOICE5570),
    .O(\CHOICE5572/FROM )
  );
  defparam \DLX_EXinst__n0007<2>3321_SW0_SW0 .INIT = 16'hCCC8;
  X_LUT4 \DLX_EXinst__n0007<2>3321_SW0_SW0  (
    .ADR0(CHOICE5545),
    .ADR1(DLX_EXinst__n0036),
    .ADR2(CHOICE5553),
    .ADR3(CHOICE5572),
    .O(\CHOICE5572/GROM )
  );
  X_BUF \CHOICE5572/XUSED  (
    .I(\CHOICE5572/FROM ),
    .O(CHOICE5572)
  );
  X_BUF \CHOICE5572/YUSED  (
    .I(\CHOICE5572/GROM ),
    .O(N164587)
  );
  defparam \DLX_EXinst__n0007<29>29 .INIT = 16'hA0AC;
  X_LUT4 \DLX_EXinst__n0007<29>29  (
    .ADR0(\DLX_EXinst_Mshift__n0021_Sh[21] ),
    .ADR1(DLX_IDinst_reg_out_A[29]),
    .ADR2(\DLX_IDinst_Imm[3] ),
    .ADR3(DLX_EXinst_N73211),
    .O(\DLX_IDinst_RegFile_10_7/FROM )
  );
  defparam \DLX_EXinst__n0007<28>39 .INIT = 16'hBA10;
  X_LUT4 \DLX_EXinst__n0007<28>39  (
    .ADR0(\DLX_IDinst_Imm[2] ),
    .ADR1(DLX_EXinst_N73211),
    .ADR2(DLX_IDinst_reg_out_A[28]),
    .ADR3(\DLX_EXinst_Mshift__n0021_Sh[24] ),
    .O(\DLX_IDinst_RegFile_10_7/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_10_7/XUSED  (
    .I(\DLX_IDinst_RegFile_10_7/FROM ),
    .O(CHOICE4787)
  );
  X_BUF \DLX_IDinst_RegFile_10_7/YUSED  (
    .I(\DLX_IDinst_RegFile_10_7/GROM ),
    .O(CHOICE4861)
  );
  defparam DLX_IDinst_RegFile_19_25_1449.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_19_25_1449 (
    .I(DLX_IDinst_WB_data_eff[25]),
    .CE(DLX_IDinst__n0588),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_19_25)
  );
  defparam \DLX_EXinst__n0007<3>221 .INIT = 16'hFFAC;
  X_LUT4 \DLX_EXinst__n0007<3>221  (
    .ADR0(DLX_EXinst__n0077),
    .ADR1(DLX_EXinst__n0079),
    .ADR2(DLX_IDinst_reg_out_B[3]),
    .ADR3(DLX_EXinst_N74245),
    .O(\CHOICE5486/FROM )
  );
  defparam \DLX_EXinst__n0007<3>261_SW0 .INIT = 16'hEAC0;
  X_LUT4 \DLX_EXinst__n0007<3>261_SW0  (
    .ADR0(DLX_IDinst_reg_out_A[3]),
    .ADR1(N138371),
    .ADR2(DLX_EXinst_N75983),
    .ADR3(CHOICE5486),
    .O(\CHOICE5486/GROM )
  );
  X_BUF \CHOICE5486/XUSED  (
    .I(\CHOICE5486/FROM ),
    .O(CHOICE5486)
  );
  X_BUF \CHOICE5486/YUSED  (
    .I(\CHOICE5486/GROM ),
    .O(N163493)
  );
  defparam \DLX_EXinst__n0007<3>261 .INIT = 16'hFFF8;
  X_LUT4 \DLX_EXinst__n0007<3>261  (
    .ADR0(DLX_EXinst_ALU_result[3]),
    .ADR1(N134884),
    .ADR2(CHOICE5494),
    .ADR3(N163493),
    .O(\CHOICE5496/FROM )
  );
  defparam \DLX_EXinst__n0007<3>3321_SW0_SW0 .INIT = 16'hCCC8;
  X_LUT4 \DLX_EXinst__n0007<3>3321_SW0_SW0  (
    .ADR0(CHOICE5477),
    .ADR1(DLX_EXinst__n0036),
    .ADR2(CHOICE5469),
    .ADR3(CHOICE5496),
    .O(\CHOICE5496/GROM )
  );
  X_BUF \CHOICE5496/XUSED  (
    .I(\CHOICE5496/FROM ),
    .O(CHOICE5496)
  );
  X_BUF \CHOICE5496/YUSED  (
    .I(\CHOICE5496/GROM ),
    .O(N164601)
  );
  defparam \DLX_EXinst__n0007<4>233 .INIT = 16'hECA0;
  X_LUT4 \DLX_EXinst__n0007<4>233  (
    .ADR0(\DLX_IDinst_Imm[4] ),
    .ADR1(DLX_IDinst_reg_out_A[4]),
    .ADR2(CHOICE4373),
    .ADR3(DLX_EXinst__n0053),
    .O(\DLX_IDinst_RegFile_6_10/FROM )
  );
  defparam \DLX_EXinst__n0007<4>261 .INIT = 16'h0F04;
  X_LUT4 \DLX_EXinst__n0007<4>261  (
    .ADR0(\DLX_IDinst_Imm[4] ),
    .ADR1(CHOICE4362),
    .ADR2(DLX_EXinst__n0036),
    .ADR3(CHOICE4375),
    .O(\DLX_IDinst_RegFile_6_10/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_6_10/XUSED  (
    .I(\DLX_IDinst_RegFile_6_10/FROM ),
    .O(CHOICE4375)
  );
  X_BUF \DLX_IDinst_RegFile_6_10/YUSED  (
    .I(\DLX_IDinst_RegFile_6_10/GROM ),
    .O(CHOICE4377)
  );
  defparam DLX_IFinst_IR_previous_2.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_2 (
    .I(DLX_IFinst_IR_latched[2]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[2])
  );
  defparam DLX_IDinst_RegFile_10_8_1450.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_10_8_1450 (
    .I(DLX_IDinst_WB_data_eff[8]),
    .CE(DLX_IDinst__n0570),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_10_8)
  );
  defparam \DLX_EXinst__n0007<4>165 .INIT = 16'hF8F8;
  X_LUT4 \DLX_EXinst__n0007<4>165  (
    .ADR0(DLX_IDinst_reg_out_A[4]),
    .ADR1(DLX_EXinst__n0054),
    .ADR2(CHOICE4360),
    .ADR3(VCC),
    .O(\DLX_IDinst_RegFile_10_8/FROM )
  );
  defparam \DLX_EXinst__n0007<4>174 .INIT = 16'hFF40;
  X_LUT4 \DLX_EXinst__n0007<4>174  (
    .ADR0(\DLX_IDinst_Imm[3] ),
    .ADR1(DLX_EXinst_N76318),
    .ADR2(DLX_EXinst_N72983),
    .ADR3(CHOICE4361),
    .O(\DLX_IDinst_RegFile_10_8/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_10_8/XUSED  (
    .I(\DLX_IDinst_RegFile_10_8/FROM ),
    .O(CHOICE4361)
  );
  X_BUF \DLX_IDinst_RegFile_10_8/YUSED  (
    .I(\DLX_IDinst_RegFile_10_8/GROM ),
    .O(CHOICE4362)
  );
  defparam DLX_IDinst_RegFile_27_17_1451.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_27_17_1451 (
    .I(DLX_IDinst_WB_data_eff[17]),
    .CE(DLX_IDinst__n0604),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_27_17)
  );
  defparam DLX_IFinst_IR_previous_7.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_7 (
    .I(DLX_IFinst_IR_latched[7]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[7])
  );
  defparam DLX_EXinst_ALU_result_4_1_1452.INIT = 1'b0;
  X_SFF DLX_EXinst_ALU_result_4_1_1452 (
    .I(\DLX_EXinst_ALU_result<4>/GROM ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(N136886),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_ALU_result_4_1)
  );
  defparam \DLX_EXinst__n0007<4>273 .INIT = 16'hFFA8;
  X_LUT4 \DLX_EXinst__n0007<4>273  (
    .ADR0(DLX_EXinst__n0036),
    .ADR1(CHOICE4347),
    .ADR2(CHOICE4332),
    .ADR3(CHOICE4377),
    .O(\DLX_EXinst_ALU_result<4>/FROM )
  );
  defparam \DLX_EXinst__n0007<4>2851 .INIT = 16'hFFA0;
  X_LUT4 \DLX_EXinst__n0007<4>2851  (
    .ADR0(DLX_EXinst_N73959),
    .ADR1(VCC),
    .ADR2(DLX_EXinst__n0012[4]),
    .ADR3(CHOICE4378),
    .O(\DLX_EXinst_ALU_result<4>/GROM )
  );
  X_BUF \DLX_EXinst_ALU_result<4>/XUSED  (
    .I(\DLX_EXinst_ALU_result<4>/FROM ),
    .O(CHOICE4378)
  );
  X_BUF \DLX_EXinst_ALU_result<4>/YUSED  (
    .I(\DLX_EXinst_ALU_result<4>/GROM ),
    .O(N162850)
  );
  defparam DLX_IFinst_IR_previous_8.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_8 (
    .I(DLX_IFinst_IR_latched[8]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[8])
  );
  defparam DLX_IDinst_RegFile_6_11_1453.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_6_11_1453 (
    .I(DLX_IDinst_WB_data_eff[11]),
    .CE(DLX_IDinst__n0562),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_6_11)
  );
  defparam DLX_EXinst_Ker7515711.INIT = 16'h40C0;
  X_LUT4 DLX_EXinst_Ker7515711 (
    .ADR0(DLX_IDinst_Imm_1_1),
    .ADR1(\DLX_IDinst_Imm[5] ),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(DLX_IDinst_Imm_2_1),
    .O(\DLX_IDinst_RegFile_6_11/FROM )
  );
  defparam \DLX_EXinst__n0007<5>143 .INIT = 16'hF888;
  X_LUT4 \DLX_EXinst__n0007<5>143  (
    .ADR0(CHOICE3969),
    .ADR1(\DLX_IDinst_Imm[5] ),
    .ADR2(\DLX_IDinst_Imm[4] ),
    .ADR3(N144646),
    .O(\DLX_IDinst_RegFile_6_11/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_6_11/XUSED  (
    .I(\DLX_IDinst_RegFile_6_11/FROM ),
    .O(CHOICE1859)
  );
  X_BUF \DLX_IDinst_RegFile_6_11/YUSED  (
    .I(\DLX_IDinst_RegFile_6_11/GROM ),
    .O(CHOICE3971)
  );
  defparam \DLX_EXinst__n0007<6>168 .INIT = 16'h0040;
  X_LUT4 \DLX_EXinst__n0007<6>168  (
    .ADR0(N146478),
    .ADR1(DLX_EXinst_N72993),
    .ADR2(DLX_EXinst__n0055),
    .ADR3(\DLX_IDinst_Imm[3] ),
    .O(\DLX_IFinst_PC<11>/FROM )
  );
  defparam \DLX_EXinst__n0007<5>168 .INIT = 16'h0040;
  X_LUT4 \DLX_EXinst__n0007<5>168  (
    .ADR0(N146478),
    .ADR1(DLX_EXinst_N72988),
    .ADR2(DLX_EXinst__n0055),
    .ADR3(\DLX_IDinst_Imm[3] ),
    .O(\DLX_IFinst_PC<11>/GROM )
  );
  X_BUF \DLX_IFinst_PC<11>/XUSED  (
    .I(\DLX_IFinst_PC<11>/FROM ),
    .O(CHOICE3921)
  );
  X_BUF \DLX_IFinst_PC<11>/YUSED  (
    .I(\DLX_IFinst_PC<11>/GROM ),
    .O(CHOICE3980)
  );
  defparam \DLX_EXinst__n0007<5>198 .INIT = 16'h8C88;
  X_LUT4 \DLX_EXinst__n0007<5>198  (
    .ADR0(DLX_EXinst__n0053),
    .ADR1(DLX_IDinst_reg_out_A[5]),
    .ADR2(\DLX_IDinst_Imm[5] ),
    .ADR3(DLX_EXinst__n0054),
    .O(\CHOICE3986/FROM )
  );
  defparam \DLX_EXinst__n0007<5>202 .INIT = 16'hFF32;
  X_LUT4 \DLX_EXinst__n0007<5>202  (
    .ADR0(CHOICE3977),
    .ADR1(\DLX_IDinst_Imm[4] ),
    .ADR2(CHOICE3980),
    .ADR3(CHOICE3986),
    .O(\CHOICE3986/GROM )
  );
  X_BUF \CHOICE3986/XUSED  (
    .I(\CHOICE3986/FROM ),
    .O(CHOICE3986)
  );
  X_BUF \CHOICE3986/YUSED  (
    .I(\CHOICE3986/GROM ),
    .O(CHOICE3987)
  );
  defparam \DLX_EXinst__n0007<3>98_SW0 .INIT = 16'hB080;
  X_LUT4 \DLX_EXinst__n0007<3>98_SW0  (
    .ADR0(N133984),
    .ADR1(\DLX_IDinst_Imm[2] ),
    .ADR2(DLX_EXinst_N76473),
    .ADR3(CHOICE5447),
    .O(\DLX_IDinst_RegFile_14_31/FROM )
  );
  defparam \DLX_EXinst__n0007<6>162 .INIT = 16'hE200;
  X_LUT4 \DLX_EXinst__n0007<6>162  (
    .ADR0(N134056),
    .ADR1(\DLX_IDinst_Imm[2] ),
    .ADR2(DLX_EXinst_N74936),
    .ADR3(DLX_EXinst_N73267),
    .O(\DLX_IDinst_RegFile_14_31/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_14_31/XUSED  (
    .I(\DLX_IDinst_RegFile_14_31/FROM ),
    .O(N163542)
  );
  X_BUF \DLX_IDinst_RegFile_14_31/YUSED  (
    .I(\DLX_IDinst_RegFile_14_31/GROM ),
    .O(CHOICE3918)
  );
  defparam DLX_IDinst_RegFile_19_17_1454.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_19_17_1454 (
    .I(DLX_IDinst_WB_data_eff[17]),
    .CE(DLX_IDinst__n0588),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_19_17)
  );
  defparam \DLX_EXinst__n0007<6>198 .INIT = 16'hC4C0;
  X_LUT4 \DLX_EXinst__n0007<6>198  (
    .ADR0(\DLX_IDinst_Imm[6] ),
    .ADR1(DLX_IDinst_reg_out_A[6]),
    .ADR2(DLX_EXinst__n0053),
    .ADR3(DLX_EXinst__n0054),
    .O(\CHOICE3927/FROM )
  );
  defparam \DLX_EXinst__n0007<6>202 .INIT = 16'hFF32;
  X_LUT4 \DLX_EXinst__n0007<6>202  (
    .ADR0(CHOICE3918),
    .ADR1(\DLX_IDinst_Imm[4] ),
    .ADR2(CHOICE3921),
    .ADR3(CHOICE3927),
    .O(\CHOICE3927/GROM )
  );
  X_BUF \CHOICE3927/XUSED  (
    .I(\CHOICE3927/FROM ),
    .O(CHOICE3927)
  );
  X_BUF \CHOICE3927/YUSED  (
    .I(\CHOICE3927/GROM ),
    .O(CHOICE3928)
  );
  defparam \DLX_EXinst__n0007<7>134 .INIT = 16'h5600;
  X_LUT4 \DLX_EXinst__n0007<7>134  (
    .ADR0(DLX_IDinst_IR_opcode_field[1]),
    .ADR1(DLX_IDinst_reg_out_A[7]),
    .ADR2(DLX_IDinst_IR_opcode_field[0]),
    .ADR3(DLX_EXinst_N76011),
    .O(\CHOICE3851/FROM )
  );
  defparam \DLX_EXinst__n0007<7>143 .INIT = 16'hECA0;
  X_LUT4 \DLX_EXinst__n0007<7>143  (
    .ADR0(N145443),
    .ADR1(\DLX_IDinst_Imm[7] ),
    .ADR2(\DLX_IDinst_Imm[4] ),
    .ADR3(CHOICE3851),
    .O(\CHOICE3851/GROM )
  );
  X_BUF \CHOICE3851/XUSED  (
    .I(\CHOICE3851/FROM ),
    .O(CHOICE3851)
  );
  X_BUF \CHOICE3851/YUSED  (
    .I(\CHOICE3851/GROM ),
    .O(CHOICE3853)
  );
  defparam DLX_EXinst_Ker730161.INIT = 16'hF5A0;
  X_LUT4 DLX_EXinst_Ker730161 (
    .ADR0(\DLX_IDinst_Imm[3] ),
    .ADR1(VCC),
    .ADR2(\DLX_EXinst_Mshift__n0020_Sh[30] ),
    .ADR3(\DLX_EXinst_Mshift__n0022_Sh[22] ),
    .O(\DLX_IDinst_RegFile_30_16/FROM )
  );
  defparam \DLX_EXinst__n0007<7>168 .INIT = 16'h1000;
  X_LUT4 \DLX_EXinst__n0007<7>168  (
    .ADR0(\DLX_IDinst_Imm[3] ),
    .ADR1(N146478),
    .ADR2(DLX_EXinst_N72998),
    .ADR3(DLX_EXinst__n0055),
    .O(\DLX_IDinst_RegFile_30_16/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_30_16/XUSED  (
    .I(\DLX_IDinst_RegFile_30_16/FROM ),
    .O(DLX_EXinst_N73018)
  );
  X_BUF \DLX_IDinst_RegFile_30_16/YUSED  (
    .I(\DLX_IDinst_RegFile_30_16/GROM ),
    .O(CHOICE3862)
  );
  defparam DLX_IDinst_Ker10822633.INIT = 16'h00FA;
  X_LUT4 DLX_IDinst_Ker10822633 (
    .ADR0(DLX_IDinst__n0105),
    .ADR1(VCC),
    .ADR2(DLX_IDinst__n0102),
    .ADR3(DLX_IDinst__n0381),
    .O(\DLX_IDinst_RegFile_22_17/FROM )
  );
  defparam \DLX_IDinst__n0142<3>_SW0_SW0 .INIT = 16'h33B3;
  X_LUT4 \DLX_IDinst__n0142<3>_SW0_SW0  (
    .ADR0(DLX_IDinst__n0439),
    .ADR1(DLX_IDinst_N108152),
    .ADR2(DLX_IDinst__n0105),
    .ADR3(DLX_IDinst__n0381),
    .O(\DLX_IDinst_RegFile_22_17/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_22_17/XUSED  (
    .I(\DLX_IDinst_RegFile_22_17/FROM ),
    .O(CHOICE3377)
  );
  X_BUF \DLX_IDinst_RegFile_22_17/YUSED  (
    .I(\DLX_IDinst_RegFile_22_17/GROM ),
    .O(N164150)
  );
  defparam \DLX_EXinst__n0007<7>198 .INIT = 16'hCE00;
  X_LUT4 \DLX_EXinst__n0007<7>198  (
    .ADR0(DLX_EXinst__n0054),
    .ADR1(DLX_EXinst__n0053),
    .ADR2(\DLX_IDinst_Imm[7] ),
    .ADR3(DLX_IDinst_reg_out_A[7]),
    .O(\CHOICE3868/FROM )
  );
  defparam \DLX_EXinst__n0007<7>202 .INIT = 16'hFF0E;
  X_LUT4 \DLX_EXinst__n0007<7>202  (
    .ADR0(CHOICE3859),
    .ADR1(CHOICE3862),
    .ADR2(\DLX_IDinst_Imm[4] ),
    .ADR3(CHOICE3868),
    .O(\CHOICE3868/GROM )
  );
  X_BUF \CHOICE3868/XUSED  (
    .I(\CHOICE3868/FROM ),
    .O(CHOICE3868)
  );
  X_BUF \CHOICE3868/YUSED  (
    .I(\CHOICE3868/GROM ),
    .O(CHOICE3869)
  );
  defparam \DLX_EXinst__n0007<8>163 .INIT = 16'hECA0;
  X_LUT4 \DLX_EXinst__n0007<8>163  (
    .ADR0(DLX_EXinst_N76285),
    .ADR1(DLX_EXinst_N76463),
    .ADR2(N164155),
    .ADR3(\DLX_EXinst_Mshift__n0021_Sh[40] ),
    .O(\CHOICE5165/GROM )
  );
  X_BUF \CHOICE5165/YUSED  (
    .I(\CHOICE5165/GROM ),
    .O(CHOICE5165)
  );
  defparam \DLX_EXinst__n0007<9>178 .INIT = 16'h1E00;
  X_LUT4 \DLX_EXinst__n0007<9>178  (
    .ADR0(DLX_IDinst_IR_opcode_field[0]),
    .ADR1(DLX_IDinst_reg_out_A[9]),
    .ADR2(DLX_IDinst_IR_opcode_field[1]),
    .ADR3(DLX_EXinst_N76011),
    .O(\DLX_IDinst_RegFile_14_18/FROM )
  );
  defparam \DLX_EXinst__n0007<9>179 .INIT = 16'hAA00;
  X_LUT4 \DLX_EXinst__n0007<9>179  (
    .ADR0(\DLX_IDinst_Imm[9] ),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(CHOICE4552),
    .O(\DLX_IDinst_RegFile_14_18/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_14_18/XUSED  (
    .I(\DLX_IDinst_RegFile_14_18/FROM ),
    .O(CHOICE4552)
  );
  X_BUF \DLX_IDinst_RegFile_14_18/YUSED  (
    .I(\DLX_IDinst_RegFile_14_18/GROM ),
    .O(CHOICE4553)
  );
  defparam \DLX_EXinst__n0007<9>187 .INIT = 16'hEAAA;
  X_LUT4 \DLX_EXinst__n0007<9>187  (
    .ADR0(CHOICE4553),
    .ADR1(\DLX_IDinst_Imm[4] ),
    .ADR2(N138481),
    .ADR3(N147520),
    .O(\DLX_IDinst_RegFile_6_21/FROM )
  );
  defparam \DLX_EXinst__n0007<9>194 .INIT = 16'hFFF0;
  X_LUT4 \DLX_EXinst__n0007<9>194  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(CHOICE4545),
    .ADR3(CHOICE4554),
    .O(\DLX_IDinst_RegFile_6_21/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_6_21/XUSED  (
    .I(\DLX_IDinst_RegFile_6_21/FROM ),
    .O(CHOICE4554)
  );
  X_BUF \DLX_IDinst_RegFile_6_21/YUSED  (
    .I(\DLX_IDinst_RegFile_6_21/GROM ),
    .O(CHOICE4555)
  );
  defparam \DLX_EXinst__n0007<8>244_SW0 .INIT = 16'hA0C0;
  X_LUT4 \DLX_EXinst__n0007<8>244_SW0  (
    .ADR0(DLX_EXinst_N74706),
    .ADR1(DLX_EXinst_N74946),
    .ADR2(DLX_EXinst_N76473),
    .ADR3(\DLX_IDinst_Imm[2] ),
    .O(\N163489/FROM )
  );
  defparam \DLX_EXinst__n0007<8>244 .INIT = 16'hFFF8;
  X_LUT4 \DLX_EXinst__n0007<8>244  (
    .ADR0(CHOICE5181),
    .ADR1(\DLX_IDinst_Imm[8] ),
    .ADR2(CHOICE5186),
    .ADR3(N163489),
    .O(\N163489/GROM )
  );
  X_BUF \N163489/XUSED  (
    .I(\N163489/FROM ),
    .O(N163489)
  );
  X_BUF \N163489/YUSED  (
    .I(\N163489/GROM ),
    .O(CHOICE5188)
  );
  defparam DLX_EXinst__n000545_SW0.INIT = 16'h0040;
  X_LUT4 DLX_EXinst__n000545_SW0 (
    .ADR0(\DLX_IDinst_Imm[0] ),
    .ADR1(CHOICE2089),
    .ADR2(DLX_EXinst__n0036),
    .ADR3(DLX_IDinst_IR_function_field[5]),
    .O(\N164119/FROM )
  );
  defparam DLX_EXinst__n000545.INIT = 16'hFFFE;
  X_LUT4 DLX_EXinst__n000545 (
    .ADR0(reset_IBUF),
    .ADR1(DLX_IDinst_counter[0]),
    .ADR2(DLX_IDinst_counter[1]),
    .ADR3(N164119),
    .O(\N164119/GROM )
  );
  X_BUF \N164119/XUSED  (
    .I(\N164119/FROM ),
    .O(N164119)
  );
  X_BUF \N164119/YUSED  (
    .I(\N164119/GROM ),
    .O(N139488)
  );
  defparam \Mshift__n0000_Sh<37>1 .INIT = 16'h4400;
  X_LUT4 \Mshift__n0000_Sh<37>1  (
    .ADR0(DLX_EXinst_ALU_result[13]),
    .ADR1(DLX_EXinst_ALU_result[12]),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_ALU_result[14]),
    .O(\DLX_IDinst_RegFile_23_10/FROM )
  );
  defparam \DM_read_data<10>1 .INIT = 16'hAA10;
  X_LUT4 \DM_read_data<10>1  (
    .ADR0(DLX_EXinst_ALU_result[13]),
    .ADR1(DLX_EXinst_ALU_result[12]),
    .ADR2(RAM_read_data[10]),
    .ADR3(DLX_EXinst_ALU_result[14]),
    .O(\DLX_IDinst_RegFile_23_10/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_23_10/XUSED  (
    .I(\DLX_IDinst_RegFile_23_10/FROM ),
    .O(Mshift__n0000_Sh[37])
  );
  X_BUF \DLX_IDinst_RegFile_23_10/YUSED  (
    .I(\DLX_IDinst_RegFile_23_10/GROM ),
    .O(DM_read_data[10])
  );
  defparam \Mshift__n0000_Sh<33>1 .INIT = 16'h1100;
  X_LUT4 \Mshift__n0000_Sh<33>1  (
    .ADR0(DLX_EXinst_ALU_result[13]),
    .ADR1(DLX_EXinst_ALU_result[14]),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_ALU_result[12]),
    .O(\DLX_IDinst_RegFile_5_29/FROM )
  );
  defparam \DM_read_data<11>1 .INIT = 16'h8988;
  X_LUT4 \DM_read_data<11>1  (
    .ADR0(DLX_EXinst_ALU_result[13]),
    .ADR1(DLX_EXinst_ALU_result[14]),
    .ADR2(DLX_EXinst_ALU_result[12]),
    .ADR3(RAM_read_data[11]),
    .O(\DLX_IDinst_RegFile_5_29/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_5_29/XUSED  (
    .I(\DLX_IDinst_RegFile_5_29/FROM ),
    .O(Mshift__n0000_Sh[33])
  );
  X_BUF \DLX_IDinst_RegFile_5_29/YUSED  (
    .I(\DLX_IDinst_RegFile_5_29/GROM ),
    .O(DM_read_data[11])
  );
  defparam \Mshift__n0000_Sh<36>1 .INIT = 16'h0044;
  X_LUT4 \Mshift__n0000_Sh<36>1  (
    .ADR0(DLX_EXinst_ALU_result[13]),
    .ADR1(DLX_EXinst_ALU_result[14]),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_ALU_result[12]),
    .O(\DLX_IDinst_RegFile_14_27/FROM )
  );
  defparam \DM_read_data<12>1 .INIT = 16'hAA04;
  X_LUT4 \DM_read_data<12>1  (
    .ADR0(DLX_EXinst_ALU_result[13]),
    .ADR1(RAM_read_data[12]),
    .ADR2(DLX_EXinst_ALU_result[12]),
    .ADR3(DLX_EXinst_ALU_result[14]),
    .O(\DLX_IDinst_RegFile_14_27/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_14_27/XUSED  (
    .I(\DLX_IDinst_RegFile_14_27/FROM ),
    .O(Mshift__n0000_Sh[36])
  );
  X_BUF \DLX_IDinst_RegFile_14_27/YUSED  (
    .I(\DLX_IDinst_RegFile_14_27/GROM ),
    .O(DM_read_data[12])
  );
  defparam \DM_read_data<24>1 .INIT = 16'hCC10;
  X_LUT4 \DM_read_data<24>1  (
    .ADR0(DLX_EXinst_ALU_result[12]),
    .ADR1(DLX_EXinst_ALU_result[13]),
    .ADR2(RAM_read_data[24]),
    .ADR3(DLX_EXinst_ALU_result[14]),
    .O(\DLX_IDinst_RegFile_6_22/FROM )
  );
  defparam \DM_read_data<20>1 .INIT = 16'hAA04;
  X_LUT4 \DM_read_data<20>1  (
    .ADR0(DLX_EXinst_ALU_result[13]),
    .ADR1(RAM_read_data[20]),
    .ADR2(DLX_EXinst_ALU_result[12]),
    .ADR3(DLX_EXinst_ALU_result[14]),
    .O(\DLX_IDinst_RegFile_6_22/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_6_22/XUSED  (
    .I(\DLX_IDinst_RegFile_6_22/FROM ),
    .O(DM_read_data[24])
  );
  X_BUF \DLX_IDinst_RegFile_6_22/YUSED  (
    .I(\DLX_IDinst_RegFile_6_22/GROM ),
    .O(DM_read_data[20])
  );
  defparam \DM_read_data<25>1 .INIT = 16'hAA10;
  X_LUT4 \DM_read_data<25>1  (
    .ADR0(DLX_EXinst_ALU_result[14]),
    .ADR1(DLX_EXinst_ALU_result[12]),
    .ADR2(RAM_read_data[25]),
    .ADR3(DLX_EXinst_ALU_result[13]),
    .O(\DLX_IDinst_RegFile_22_19/FROM )
  );
  defparam \DM_read_data<13>1 .INIT = 16'hAA04;
  X_LUT4 \DM_read_data<13>1  (
    .ADR0(DLX_EXinst_ALU_result[14]),
    .ADR1(RAM_read_data[13]),
    .ADR2(DLX_EXinst_ALU_result[12]),
    .ADR3(DLX_EXinst_ALU_result[13]),
    .O(\DLX_IDinst_RegFile_22_19/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_22_19/XUSED  (
    .I(\DLX_IDinst_RegFile_22_19/FROM ),
    .O(DM_read_data[25])
  );
  X_BUF \DLX_IDinst_RegFile_22_19/YUSED  (
    .I(\DLX_IDinst_RegFile_22_19/GROM ),
    .O(DM_read_data[13])
  );
  defparam \DM_read_data<26>1 .INIT = 16'hA0A4;
  X_LUT4 \DM_read_data<26>1  (
    .ADR0(DLX_EXinst_ALU_result[14]),
    .ADR1(RAM_read_data[26]),
    .ADR2(DLX_EXinst_ALU_result[13]),
    .ADR3(DLX_EXinst_ALU_result[12]),
    .O(\DLX_IDinst_RegFile_6_14/FROM )
  );
  defparam \DM_read_data<21>1 .INIT = 16'h8988;
  X_LUT4 \DM_read_data<21>1  (
    .ADR0(DLX_EXinst_ALU_result[14]),
    .ADR1(DLX_EXinst_ALU_result[13]),
    .ADR2(DLX_EXinst_ALU_result[12]),
    .ADR3(RAM_read_data[21]),
    .O(\DLX_IDinst_RegFile_6_14/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_6_14/XUSED  (
    .I(\DLX_IDinst_RegFile_6_14/FROM ),
    .O(DM_read_data[26])
  );
  X_BUF \DLX_IDinst_RegFile_6_14/YUSED  (
    .I(\DLX_IDinst_RegFile_6_14/GROM ),
    .O(DM_read_data[21])
  );
  defparam \DM_read_data<27>1 .INIT = 16'hAA10;
  X_LUT4 \DM_read_data<27>1  (
    .ADR0(DLX_EXinst_ALU_result[13]),
    .ADR1(DLX_EXinst_ALU_result[12]),
    .ADR2(RAM_read_data[27]),
    .ADR3(DLX_EXinst_ALU_result[14]),
    .O(\DLX_IDinst_RegFile_6_30/FROM )
  );
  defparam \DM_read_data<30>1 .INIT = 16'hCC10;
  X_LUT4 \DM_read_data<30>1  (
    .ADR0(DLX_EXinst_ALU_result[12]),
    .ADR1(DLX_EXinst_ALU_result[13]),
    .ADR2(RAM_read_data[30]),
    .ADR3(DLX_EXinst_ALU_result[14]),
    .O(\DLX_IDinst_RegFile_6_30/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_6_30/XUSED  (
    .I(\DLX_IDinst_RegFile_6_30/FROM ),
    .O(DM_read_data[27])
  );
  X_BUF \DLX_IDinst_RegFile_6_30/YUSED  (
    .I(\DLX_IDinst_RegFile_6_30/GROM ),
    .O(DM_read_data[30])
  );
  defparam \DM_read_data<28>1 .INIT = 16'hF004;
  X_LUT4 \DM_read_data<28>1  (
    .ADR0(DLX_EXinst_ALU_result[12]),
    .ADR1(RAM_read_data[28]),
    .ADR2(DLX_EXinst_ALU_result[14]),
    .ADR3(DLX_EXinst_ALU_result[13]),
    .O(\DLX_IDinst_RegFile_6_31/FROM )
  );
  defparam \DM_read_data<14>1 .INIT = 16'hC1C0;
  X_LUT4 \DM_read_data<14>1  (
    .ADR0(DLX_EXinst_ALU_result[12]),
    .ADR1(DLX_EXinst_ALU_result[13]),
    .ADR2(DLX_EXinst_ALU_result[14]),
    .ADR3(RAM_read_data[14]),
    .O(\DLX_IDinst_RegFile_6_31/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_6_31/XUSED  (
    .I(\DLX_IDinst_RegFile_6_31/FROM ),
    .O(DM_read_data[28])
  );
  X_BUF \DLX_IDinst_RegFile_6_31/YUSED  (
    .I(\DLX_IDinst_RegFile_6_31/GROM ),
    .O(DM_read_data[14])
  );
  defparam \DM_read_data<29>1 .INIT = 16'h8898;
  X_LUT4 \DM_read_data<29>1  (
    .ADR0(DLX_EXinst_ALU_result[14]),
    .ADR1(DLX_EXinst_ALU_result[13]),
    .ADR2(RAM_read_data[29]),
    .ADR3(DLX_EXinst_ALU_result[12]),
    .O(\DLX_IDinst_RegFile_6_15/FROM )
  );
  defparam \DM_read_data<22>1 .INIT = 16'h8988;
  X_LUT4 \DM_read_data<22>1  (
    .ADR0(DLX_EXinst_ALU_result[14]),
    .ADR1(DLX_EXinst_ALU_result[13]),
    .ADR2(DLX_EXinst_ALU_result[12]),
    .ADR3(RAM_read_data[22]),
    .O(\DLX_IDinst_RegFile_6_15/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_6_15/XUSED  (
    .I(\DLX_IDinst_RegFile_6_15/FROM ),
    .O(DM_read_data[29])
  );
  X_BUF \DLX_IDinst_RegFile_6_15/YUSED  (
    .I(\DLX_IDinst_RegFile_6_15/GROM ),
    .O(DM_read_data[22])
  );
  defparam \DM_read_data<1>1 .INIT = 16'hC0C2;
  X_LUT4 \DM_read_data<1>1  (
    .ADR0(RAM_read_data[1]),
    .ADR1(DLX_EXinst_ALU_result[14]),
    .ADR2(DLX_EXinst_ALU_result[13]),
    .ADR3(DLX_EXinst_ALU_result[12]),
    .O(\DM_read_data<1>/FROM )
  );
  defparam \DM_read_data<31>1 .INIT = 16'hA1A0;
  X_LUT4 \DM_read_data<31>1  (
    .ADR0(DLX_EXinst_ALU_result[13]),
    .ADR1(DLX_EXinst_ALU_result[12]),
    .ADR2(DLX_EXinst_ALU_result[14]),
    .ADR3(RAM_read_data[31]),
    .O(\DM_read_data<1>/GROM )
  );
  X_BUF \DM_read_data<1>/XUSED  (
    .I(\DM_read_data<1>/FROM ),
    .O(DM_read_data[1])
  );
  X_BUF \DM_read_data<1>/YUSED  (
    .I(\DM_read_data<1>/GROM ),
    .O(DM_read_data[31])
  );
  defparam \DM_read_data<2>1 .INIT = 16'hCC10;
  X_LUT4 \DM_read_data<2>1  (
    .ADR0(DLX_EXinst_ALU_result[12]),
    .ADR1(DLX_EXinst_ALU_result[13]),
    .ADR2(RAM_read_data[2]),
    .ADR3(DLX_EXinst_ALU_result[14]),
    .O(\DM_read_data<2>/FROM )
  );
  defparam \DM_read_data<15>1 .INIT = 16'hCC10;
  X_LUT4 \DM_read_data<15>1  (
    .ADR0(DLX_EXinst_ALU_result[12]),
    .ADR1(DLX_EXinst_ALU_result[13]),
    .ADR2(RAM_read_data[15]),
    .ADR3(DLX_EXinst_ALU_result[14]),
    .O(\DM_read_data<2>/GROM )
  );
  X_BUF \DM_read_data<2>/XUSED  (
    .I(\DM_read_data<2>/FROM ),
    .O(DM_read_data[2])
  );
  X_BUF \DM_read_data<2>/YUSED  (
    .I(\DM_read_data<2>/GROM ),
    .O(DM_read_data[15])
  );
  defparam \DM_read_data<3>1 .INIT = 16'hAA10;
  X_LUT4 \DM_read_data<3>1  (
    .ADR0(DLX_EXinst_ALU_result[14]),
    .ADR1(DLX_EXinst_ALU_result[12]),
    .ADR2(RAM_read_data[3]),
    .ADR3(DLX_EXinst_ALU_result[13]),
    .O(\DLX_IDinst_RegFile_6_24/FROM )
  );
  defparam \DM_read_data<23>1 .INIT = 16'hCC10;
  X_LUT4 \DM_read_data<23>1  (
    .ADR0(DLX_EXinst_ALU_result[12]),
    .ADR1(DLX_EXinst_ALU_result[14]),
    .ADR2(RAM_read_data[23]),
    .ADR3(DLX_EXinst_ALU_result[13]),
    .O(\DLX_IDinst_RegFile_6_24/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_6_24/XUSED  (
    .I(\DLX_IDinst_RegFile_6_24/FROM ),
    .O(DM_read_data[3])
  );
  X_BUF \DLX_IDinst_RegFile_6_24/YUSED  (
    .I(\DLX_IDinst_RegFile_6_24/GROM ),
    .O(DM_read_data[23])
  );
  defparam \DM_read_data<4>1 .INIT = 16'hF004;
  X_LUT4 \DM_read_data<4>1  (
    .ADR0(DLX_EXinst_ALU_result[12]),
    .ADR1(RAM_read_data[4]),
    .ADR2(DLX_EXinst_ALU_result[13]),
    .ADR3(DLX_EXinst_ALU_result[14]),
    .O(\DLX_IDinst_RegFile_6_17/FROM )
  );
  defparam \DM_read_data<16>1 .INIT = 16'hF004;
  X_LUT4 \DM_read_data<16>1  (
    .ADR0(DLX_EXinst_ALU_result[12]),
    .ADR1(RAM_read_data[16]),
    .ADR2(DLX_EXinst_ALU_result[14]),
    .ADR3(DLX_EXinst_ALU_result[13]),
    .O(\DLX_IDinst_RegFile_6_17/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_6_17/XUSED  (
    .I(\DLX_IDinst_RegFile_6_17/FROM ),
    .O(DM_read_data[4])
  );
  X_BUF \DLX_IDinst_RegFile_6_17/YUSED  (
    .I(\DLX_IDinst_RegFile_6_17/GROM ),
    .O(DM_read_data[16])
  );
  defparam \DM_read_data<5>1 .INIT = 16'h8898;
  X_LUT4 \DM_read_data<5>1  (
    .ADR0(DLX_EXinst_ALU_result[13]),
    .ADR1(DLX_EXinst_ALU_result[14]),
    .ADR2(RAM_read_data[5]),
    .ADR3(DLX_EXinst_ALU_result[12]),
    .O(\DLX_IDinst_RegFile_6_25/FROM )
  );
  defparam \DM_read_data<17>1 .INIT = 16'hCC10;
  X_LUT4 \DM_read_data<17>1  (
    .ADR0(DLX_EXinst_ALU_result[12]),
    .ADR1(DLX_EXinst_ALU_result[13]),
    .ADR2(RAM_read_data[17]),
    .ADR3(DLX_EXinst_ALU_result[14]),
    .O(\DLX_IDinst_RegFile_6_25/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_6_25/XUSED  (
    .I(\DLX_IDinst_RegFile_6_25/FROM ),
    .O(DM_read_data[5])
  );
  X_BUF \DLX_IDinst_RegFile_6_25/YUSED  (
    .I(\DLX_IDinst_RegFile_6_25/GROM ),
    .O(DM_read_data[17])
  );
  defparam \DM_read_data<6>1 .INIT = 16'hF002;
  X_LUT4 \DM_read_data<6>1  (
    .ADR0(RAM_read_data[6]),
    .ADR1(DLX_EXinst_ALU_result[12]),
    .ADR2(DLX_EXinst_ALU_result[13]),
    .ADR3(DLX_EXinst_ALU_result[14]),
    .O(\DLX_IDinst_RegFile_7_10/FROM )
  );
  defparam \DM_read_data<18>1 .INIT = 16'hC0C2;
  X_LUT4 \DM_read_data<18>1  (
    .ADR0(RAM_read_data[18]),
    .ADR1(DLX_EXinst_ALU_result[13]),
    .ADR2(DLX_EXinst_ALU_result[14]),
    .ADR3(DLX_EXinst_ALU_result[12]),
    .O(\DLX_IDinst_RegFile_7_10/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_7_10/XUSED  (
    .I(\DLX_IDinst_RegFile_7_10/FROM ),
    .O(DM_read_data[6])
  );
  X_BUF \DLX_IDinst_RegFile_7_10/YUSED  (
    .I(\DLX_IDinst_RegFile_7_10/GROM ),
    .O(DM_read_data[18])
  );
  defparam DLX_EXinst__n001480_SW0.INIT = 16'hFEFE;
  X_LUT4 DLX_EXinst__n001480_SW0 (
    .ADR0(CHOICE3010),
    .ADR1(DLX_IDinst_IR_opcode_field[2]),
    .ADR2(DLX_IDinst_IR_opcode_field[1]),
    .ADR3(VCC),
    .O(\DLX_IDinst_RegFile_6_18/FROM )
  );
  defparam DLX_EXinst__n001480.INIT = 16'hFBF8;
  X_LUT4 DLX_EXinst__n001480 (
    .ADR0(N163158),
    .ADR1(DLX_IDinst_IR_opcode_field[5]),
    .ADR2(DLX_IDinst_IR_opcode_field[4]),
    .ADR3(N163156),
    .O(\DLX_IDinst_RegFile_6_18/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_6_18/XUSED  (
    .I(\DLX_IDinst_RegFile_6_18/FROM ),
    .O(N163156)
  );
  X_BUF \DLX_IDinst_RegFile_6_18/YUSED  (
    .I(\DLX_IDinst_RegFile_6_18/GROM ),
    .O(N144912)
  );
  defparam DLX_EXinst_Ker7621812.INIT = 16'h0002;
  X_LUT4 DLX_EXinst_Ker7621812 (
    .ADR0(DLX_IDinst_IR_opcode_field[3]),
    .ADR1(DLX_IDinst_IR_opcode_field[0]),
    .ADR2(DLX_IDinst_IR_opcode_field[5]),
    .ADR3(DLX_IDinst_IR_opcode_field[2]),
    .O(\CHOICE1669/FROM )
  );
  defparam DLX_EXinst__n001480_SW1.INIT = 16'hFA30;
  X_LUT4 DLX_EXinst__n001480_SW1 (
    .ADR0(DLX_IDinst_IR_opcode_field[3]),
    .ADR1(DLX_IDinst_IR_opcode_field[0]),
    .ADR2(DLX_IDinst_IR_opcode_field[1]),
    .ADR3(DLX_IDinst_IR_opcode_field[2]),
    .O(\CHOICE1669/GROM )
  );
  X_BUF \CHOICE1669/XUSED  (
    .I(\CHOICE1669/FROM ),
    .O(CHOICE1669)
  );
  X_BUF \CHOICE1669/YUSED  (
    .I(\CHOICE1669/GROM ),
    .O(N163158)
  );
  defparam \DM_read_data<7>1 .INIT = 16'hC1C0;
  X_LUT4 \DM_read_data<7>1  (
    .ADR0(DLX_EXinst_ALU_result[12]),
    .ADR1(DLX_EXinst_ALU_result[13]),
    .ADR2(DLX_EXinst_ALU_result[14]),
    .ADR3(RAM_read_data[7]),
    .O(\DLX_IDinst_RegFile_15_17/FROM )
  );
  defparam \DM_read_data<19>1 .INIT = 16'h8988;
  X_LUT4 \DM_read_data<19>1  (
    .ADR0(DLX_EXinst_ALU_result[13]),
    .ADR1(DLX_EXinst_ALU_result[14]),
    .ADR2(DLX_EXinst_ALU_result[12]),
    .ADR3(RAM_read_data[19]),
    .O(\DLX_IDinst_RegFile_15_17/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_15_17/XUSED  (
    .I(\DLX_IDinst_RegFile_15_17/FROM ),
    .O(DM_read_data[7])
  );
  X_BUF \DLX_IDinst_RegFile_15_17/YUSED  (
    .I(\DLX_IDinst_RegFile_15_17/GROM ),
    .O(DM_read_data[19])
  );
  defparam \DLX_EXinst__n0007<10>194_SW0 .INIT = 16'hCA00;
  X_LUT4 \DLX_EXinst__n0007<10>194_SW0  (
    .ADR0(DLX_EXinst_N74936),
    .ADR1(DLX_EXinst_N74701),
    .ADR2(\DLX_IDinst_Imm[2] ),
    .ADR3(DLX_EXinst_N76473),
    .O(\N163688/FROM )
  );
  defparam \DLX_EXinst__n0007<10>194 .INIT = 16'hFFEC;
  X_LUT4 \DLX_EXinst__n0007<10>194  (
    .ADR0(\DLX_IDinst_Imm[10] ),
    .ADR1(CHOICE4493),
    .ADR2(CHOICE4490),
    .ADR3(N163688),
    .O(\N163688/GROM )
  );
  X_BUF \N163688/XUSED  (
    .I(\N163688/FROM ),
    .O(N163688)
  );
  X_BUF \N163688/YUSED  (
    .I(\N163688/GROM ),
    .O(CHOICE4495)
  );
  defparam DLX_IDinst_Ker108231_SW0.INIT = 16'h2F2A;
  X_LUT4 DLX_IDinst_Ker108231_SW0 (
    .ADR0(DLX_IDinst_stall),
    .ADR1(DLX_IDinst_slot_num_FFd2),
    .ADR2(DLX_IDinst_delay_slot),
    .ADR3(FREEZE_IBUF),
    .O(\N132648/FROM )
  );
  defparam DLX_IDinst__n06171.INIT = 16'h0001;
  X_LUT4 DLX_IDinst__n06171 (
    .ADR0(reset_IBUF),
    .ADR1(DLX_IDinst_N108100),
    .ADR2(DLX_IDinst__n0376),
    .ADR3(N132648),
    .O(\N132648/GROM )
  );
  X_BUF \N132648/XUSED  (
    .I(\N132648/FROM ),
    .O(N132648)
  );
  X_BUF \N132648/YUSED  (
    .I(\N132648/GROM ),
    .O(DLX_IDinst__n0617)
  );
  defparam DLX_IFinst__n00001.INIT = 16'hFFFC;
  X_LUT4 DLX_IFinst__n00001 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_counter[1]),
    .ADR2(DLX_IDinst_counter[0]),
    .ADR3(DLX_IDinst_stall),
    .O(\DLX_IFinst_stalled/FROM )
  );
  defparam DLX_IFinst_PC_ClkEn_INV1.INIT = 16'h0001;
  X_LUT4 DLX_IFinst_PC_ClkEn_INV1 (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(DLX_IDinst_stall),
    .ADR2(DLX_IDinst_counter[1]),
    .ADR3(DLX_IDinst_counter[0]),
    .O(\DLX_IFinst_stalled/GROM )
  );
  X_INV \DLX_IFinst_stalled/CEMUX  (
    .I(DLX_IDinst_branch_sig),
    .O(\DLX_IFinst_stalled/CEMUXNOT )
  );
  X_BUF \DLX_IFinst_stalled/XUSED  (
    .I(\DLX_IFinst_stalled/FROM ),
    .O(DLX_IFinst__n0000)
  );
  X_BUF \DLX_IFinst_stalled/YUSED  (
    .I(\DLX_IFinst_stalled/GROM ),
    .O(DLX_IFinst_PC_N3087)
  );
  defparam DLX_IDinst_Ker107570_SW0.INIT = 16'h0200;
  X_LUT4 DLX_IDinst_Ker107570_SW0 (
    .ADR0(DLX_IDinst__n0629[1]),
    .ADR1(DLX_IDinst__n0381),
    .ADR2(DLX_IDinst__n0439),
    .ADR3(DLX_IDinst__n0105),
    .O(\N127012/FROM )
  );
  defparam DLX_IDinst_Ker107570.INIT = 16'hFF08;
  X_LUT4 DLX_IDinst_Ker107570 (
    .ADR0(DLX_IDinst__n0313),
    .ADR1(DLX_IDinst_N108443),
    .ADR2(DLX_IDinst__n0437),
    .ADR3(N127012),
    .O(\N127012/GROM )
  );
  X_BUF \N127012/XUSED  (
    .I(\N127012/FROM ),
    .O(N127012)
  );
  X_BUF \N127012/YUSED  (
    .I(\N127012/GROM ),
    .O(DLX_IDinst_N107572)
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<6>_SW0 .INIT = 16'hCFC0;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<6>_SW0  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[3]),
    .ADR2(DLX_IDinst_reg_out_B[1]),
    .ADR3(DLX_IDinst_reg_out_A[5]),
    .O(\DLX_IDinst_RegFile_6_27/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<6> .INIT = 16'hEE44;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<6>  (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(DLX_EXinst_N73599),
    .ADR2(VCC),
    .ADR3(N130977),
    .O(\DLX_IDinst_RegFile_6_27/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_6_27/XUSED  (
    .I(\DLX_IDinst_RegFile_6_27/FROM ),
    .O(N130977)
  );
  X_BUF \DLX_IDinst_RegFile_6_27/YUSED  (
    .I(\DLX_IDinst_RegFile_6_27/GROM ),
    .O(\DLX_EXinst_Mshift__n0023_Sh[6] )
  );
  defparam \DLX_EXinst__n0007<11>194_SW0 .INIT = 16'hAC00;
  X_LUT4 \DLX_EXinst__n0007<11>194_SW0  (
    .ADR0(DLX_EXinst_N75139),
    .ADR1(DLX_EXinst_N74941),
    .ADR2(\DLX_IDinst_Imm[2] ),
    .ADR3(DLX_EXinst_N76473),
    .O(\N163230/FROM )
  );
  defparam \DLX_EXinst__n0007<11>194 .INIT = 16'hFFF8;
  X_LUT4 \DLX_EXinst__n0007<11>194  (
    .ADR0(CHOICE4430),
    .ADR1(\DLX_IDinst_Imm[11] ),
    .ADR2(CHOICE4433),
    .ADR3(N163230),
    .O(\N163230/GROM )
  );
  X_BUF \N163230/XUSED  (
    .I(\N163230/FROM ),
    .O(N163230)
  );
  X_BUF \N163230/YUSED  (
    .I(\N163230/GROM ),
    .O(CHOICE4435)
  );
  defparam \DLX_EXinst_Mshift__n0020_Sh<27> .INIT = 16'hFC0C;
  X_LUT4 \DLX_EXinst_Mshift__n0020_Sh<27>  (
    .ADR0(VCC),
    .ADR1(N130467),
    .ADR2(DLX_IDinst_Imm_1_1),
    .ADR3(DLX_EXinst_N72791),
    .O(\DLX_IDinst_RegFile_31_18/FROM )
  );
  defparam DLX_EXinst_Ker753501.INIT = 16'hEE22;
  X_LUT4 DLX_EXinst_Ker753501 (
    .ADR0(\DLX_EXinst_Mshift__n0022_Sh[19] ),
    .ADR1(DLX_IDinst_Imm_3_1),
    .ADR2(VCC),
    .ADR3(\DLX_EXinst_Mshift__n0020_Sh[27] ),
    .O(\DLX_IDinst_RegFile_31_18/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_31_18/XUSED  (
    .I(\DLX_IDinst_RegFile_31_18/FROM ),
    .O(\DLX_EXinst_Mshift__n0020_Sh[27] )
  );
  X_BUF \DLX_IDinst_RegFile_31_18/YUSED  (
    .I(\DLX_IDinst_RegFile_31_18/GROM ),
    .O(DLX_EXinst_N75352)
  );
  defparam \DLX_IDinst__n0146<20>36_SW0 .INIT = 16'hBB5F;
  X_LUT4 \DLX_IDinst__n0146<20>36_SW0  (
    .ADR0(DLX_IDinst_jtarget[22]),
    .ADR1(\DLX_IDinst_Cause_Reg[31] ),
    .ADR2(DLX_IDinst_EPC[20]),
    .ADR3(DLX_IDinst_jtarget[21]),
    .O(\N163664/FROM )
  );
  defparam \DLX_IDinst__n0146<20>36 .INIT = 16'hC0EA;
  X_LUT4 \DLX_IDinst__n0146<20>36  (
    .ADR0(DLX_IDinst_N107105),
    .ADR1(\DLX_IDinst_regA_eff[20] ),
    .ADR2(N134590),
    .ADR3(N163664),
    .O(\N163664/GROM )
  );
  X_BUF \N163664/XUSED  (
    .I(\N163664/FROM ),
    .O(N163664)
  );
  X_BUF \N163664/YUSED  (
    .I(\N163664/GROM ),
    .O(CHOICE2723)
  );
  defparam reset_IBUF_1_1455.INIT = 16'hAAAA;
  X_LUT4 reset_IBUF_1_1455 (
    .ADR0(reset_IBUF),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IDinst_RegFile_7_20/FROM )
  );
  defparam vga_top_vga1__n0014_1456.INIT = 16'hFF51;
  X_LUT4 vga_top_vga1__n0014_1456 (
    .ADR0(N132456),
    .ADR1(vga_top_vga1_vcounter[5]),
    .ADR2(vga_top_vga1_N112921),
    .ADR3(reset_IBUF_1),
    .O(\DLX_IDinst_RegFile_7_20/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_7_20/XUSED  (
    .I(\DLX_IDinst_RegFile_7_20/FROM ),
    .O(reset_IBUF_1)
  );
  X_BUF \DLX_IDinst_RegFile_7_20/YUSED  (
    .I(\DLX_IDinst_RegFile_7_20/GROM ),
    .O(vga_top_vga1__n0014)
  );
  defparam DLX_IDinst_RegFile_19_26_1457.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_19_26_1457 (
    .I(DLX_IDinst_WB_data_eff[26]),
    .CE(DLX_IDinst__n0588),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_19_26)
  );
  defparam reset_IBUF_8_1458.INIT = 16'hFF00;
  X_LUT4 reset_IBUF_8_1458 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(reset_IBUF),
    .O(\DLX_IDinst_RegFile_23_27/FROM )
  );
  defparam reset_IBUF_2_1459.INIT = 16'hFF00;
  X_LUT4 reset_IBUF_2_1459 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(reset_IBUF),
    .O(\DLX_IDinst_RegFile_23_27/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_23_27/XUSED  (
    .I(\DLX_IDinst_RegFile_23_27/FROM ),
    .O(reset_IBUF_8)
  );
  X_BUF \DLX_IDinst_RegFile_23_27/YUSED  (
    .I(\DLX_IDinst_RegFile_23_27/GROM ),
    .O(reset_IBUF_2)
  );
  defparam reset_IBUF_7_1460.INIT = 16'hFF00;
  X_LUT4 reset_IBUF_7_1460 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(reset_IBUF),
    .O(\DLX_IDinst_RegFile_7_12/FROM )
  );
  defparam reset_IBUF_3_1461.INIT = 16'hFF00;
  X_LUT4 reset_IBUF_3_1461 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(reset_IBUF),
    .O(\DLX_IDinst_RegFile_7_12/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_7_12/XUSED  (
    .I(\DLX_IDinst_RegFile_7_12/FROM ),
    .O(reset_IBUF_7)
  );
  X_BUF \DLX_IDinst_RegFile_7_12/YUSED  (
    .I(\DLX_IDinst_RegFile_7_12/GROM ),
    .O(reset_IBUF_3)
  );
  defparam reset_IBUF_6_1462.INIT = 16'hAAAA;
  X_LUT4 reset_IBUF_6_1462 (
    .ADR0(reset_IBUF),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IDinst_RegFile_31_19/FROM )
  );
  defparam reset_IBUF_4_1463.INIT = 16'hFF00;
  X_LUT4 reset_IBUF_4_1463 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(reset_IBUF),
    .O(\DLX_IDinst_RegFile_31_19/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_31_19/XUSED  (
    .I(\DLX_IDinst_RegFile_31_19/FROM ),
    .O(reset_IBUF_6)
  );
  X_BUF \DLX_IDinst_RegFile_31_19/YUSED  (
    .I(\DLX_IDinst_RegFile_31_19/GROM ),
    .O(reset_IBUF_4)
  );
  defparam reset_IBUF_5_1464.INIT = 16'hAAAA;
  X_LUT4 reset_IBUF_5_1464 (
    .ADR0(reset_IBUF),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\reset_IBUF_5/GROM )
  );
  X_BUF \reset_IBUF_5/YUSED  (
    .I(\reset_IBUF_5/GROM ),
    .O(reset_IBUF_5)
  );
  defparam DLX_IDinst_Ker10707415.INIT = 16'h0057;
  X_LUT4 DLX_IDinst_Ker10707415 (
    .ADR0(DLX_IDinst_N108443),
    .ADR1(DLX_IDinst_N108221),
    .ADR2(DLX_IDinst__n0311),
    .ADR3(DLX_IDinst__n0437),
    .O(\CHOICE2112/FROM )
  );
  defparam DLX_IDinst_Ker107835_SW0.INIT = 16'h0080;
  X_LUT4 DLX_IDinst_Ker107835_SW0 (
    .ADR0(DLX_IDinst_N107033),
    .ADR1(DLX_IDinst_N108443),
    .ADR2(DLX_IDinst__n0311),
    .ADR3(DLX_IDinst__n0453),
    .O(\CHOICE2112/GROM )
  );
  X_BUF \CHOICE2112/XUSED  (
    .I(\CHOICE2112/FROM ),
    .O(CHOICE2112)
  );
  X_BUF \CHOICE2112/YUSED  (
    .I(\CHOICE2112/GROM ),
    .O(N137086)
  );
  defparam \DLX_EXinst_Mshift__n0021_Sh<0>1 .INIT = 16'h0022;
  X_LUT4 \DLX_EXinst_Mshift__n0021_Sh<0>1  (
    .ADR0(DLX_IDinst_reg_out_A[0]),
    .ADR1(DLX_IDinst_Imm_1_1),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_Imm_0_1),
    .O(\DLX_EXinst_Mshift__n0021_Sh<0>/FROM )
  );
  defparam DLX_EXinst_Ker729811.INIT = 16'hFA0A;
  X_LUT4 DLX_EXinst_Ker729811 (
    .ADR0(\DLX_EXinst_Mshift__n0021_Sh[4] ),
    .ADR1(VCC),
    .ADR2(\DLX_IDinst_Imm[2] ),
    .ADR3(\DLX_EXinst_Mshift__n0021_Sh[0] ),
    .O(\DLX_EXinst_Mshift__n0021_Sh<0>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0021_Sh<0>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0021_Sh<0>/FROM ),
    .O(\DLX_EXinst_Mshift__n0021_Sh[0] )
  );
  X_BUF \DLX_EXinst_Mshift__n0021_Sh<0>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0021_Sh<0>/GROM ),
    .O(DLX_EXinst_N72983)
  );
  defparam DLX_IDinst_RegFile_19_18_1465.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_19_18_1465 (
    .I(DLX_IDinst_WB_data_eff[18]),
    .CE(DLX_IDinst__n0588),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_19_18)
  );
  defparam \DLX_EXinst_Mshift__n0021_Sh<40> .INIT = 16'h11B1;
  X_LUT4 \DLX_EXinst_Mshift__n0021_Sh<40>  (
    .ADR0(DLX_IDinst_Imm_2_1),
    .ADR1(N131375),
    .ADR2(\DLX_EXinst_Mshift__n0021_Sh[4] ),
    .ADR3(DLX_IDinst_Imm_3_1),
    .O(\DLX_EXinst_Mshift__n0021_Sh<40>/FROM )
  );
  defparam \DLX_EXinst__n0007<24>380 .INIT = 16'hFE0E;
  X_LUT4 \DLX_EXinst__n0007<24>380  (
    .ADR0(CHOICE5667),
    .ADR1(CHOICE5668),
    .ADR2(\DLX_IDinst_Imm[4] ),
    .ADR3(\DLX_EXinst_Mshift__n0021_Sh[40] ),
    .O(\DLX_EXinst_Mshift__n0021_Sh<40>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0021_Sh<40>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0021_Sh<40>/FROM ),
    .O(\DLX_EXinst_Mshift__n0021_Sh[40] )
  );
  X_BUF \DLX_EXinst_Mshift__n0021_Sh<40>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0021_Sh<40>/GROM ),
    .O(CHOICE5671)
  );
  defparam \DLX_EXinst_Mshift__n0021_Sh<1>1 .INIT = 16'h5140;
  X_LUT4 \DLX_EXinst_Mshift__n0021_Sh<1>1  (
    .ADR0(DLX_IDinst_Imm_1_1),
    .ADR1(DLX_IDinst_Imm_0_1),
    .ADR2(DLX_IDinst_reg_out_A[0]),
    .ADR3(DLX_IDinst_reg_out_A[1]),
    .O(\DLX_EXinst_Mshift__n0021_Sh<1>/FROM )
  );
  defparam DLX_EXinst_Ker729861.INIT = 16'hEE44;
  X_LUT4 DLX_EXinst_Ker729861 (
    .ADR0(\DLX_IDinst_Imm[2] ),
    .ADR1(\DLX_EXinst_Mshift__n0021_Sh[5] ),
    .ADR2(VCC),
    .ADR3(\DLX_EXinst_Mshift__n0021_Sh[1] ),
    .O(\DLX_EXinst_Mshift__n0021_Sh<1>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0021_Sh<1>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0021_Sh<1>/FROM ),
    .O(\DLX_EXinst_Mshift__n0021_Sh[1] )
  );
  X_BUF \DLX_EXinst_Mshift__n0021_Sh<1>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0021_Sh<1>/GROM ),
    .O(DLX_EXinst_N72988)
  );
  defparam \DLX_EXinst_Mshift__n0021_Sh<42> .INIT = 16'h5303;
  X_LUT4 \DLX_EXinst_Mshift__n0021_Sh<42>  (
    .ADR0(DLX_IDinst_Imm_3_1),
    .ADR1(N131503),
    .ADR2(DLX_IDinst_Imm_2_1),
    .ADR3(\DLX_EXinst_Mshift__n0021_Sh[6] ),
    .O(\DLX_EXinst_Mshift__n0021_Sh<42>/FROM )
  );
  defparam \DLX_EXinst__n0007<26>10 .INIT = 16'h0800;
  X_LUT4 \DLX_EXinst__n0007<26>10  (
    .ADR0(DLX_EXinst__n0055),
    .ADR1(\DLX_IDinst_Imm[4] ),
    .ADR2(N146478),
    .ADR3(\DLX_EXinst_Mshift__n0021_Sh[42] ),
    .O(\DLX_EXinst_Mshift__n0021_Sh<42>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0021_Sh<42>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0021_Sh<42>/FROM ),
    .O(\DLX_EXinst_Mshift__n0021_Sh[42] )
  );
  X_BUF \DLX_EXinst_Mshift__n0021_Sh<42>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0021_Sh<42>/GROM ),
    .O(CHOICE4992)
  );
  defparam \DLX_IDinst__n0146<21>36_SW0 .INIT = 16'hF53F;
  X_LUT4 \DLX_IDinst__n0146<21>36_SW0  (
    .ADR0(\DLX_IDinst_Cause_Reg[31] ),
    .ADR1(DLX_IDinst_EPC[21]),
    .ADR2(DLX_IDinst_jtarget[22]),
    .ADR3(DLX_IDinst_jtarget[21]),
    .O(\N163442/FROM )
  );
  defparam \DLX_IDinst__n0146<21>36 .INIT = 16'h88F8;
  X_LUT4 \DLX_IDinst__n0146<21>36  (
    .ADR0(\DLX_IDinst_regA_eff[21] ),
    .ADR1(N134590),
    .ADR2(DLX_IDinst_N107105),
    .ADR3(N163442),
    .O(\N163442/GROM )
  );
  X_BUF \N163442/XUSED  (
    .I(\N163442/FROM ),
    .O(N163442)
  );
  X_BUF \N163442/YUSED  (
    .I(\N163442/GROM ),
    .O(CHOICE2738)
  );
  defparam \DLX_EXinst_Mshift__n0021_Sh<8>1 .INIT = 16'hF0AA;
  X_LUT4 \DLX_EXinst_Mshift__n0021_Sh<8>1  (
    .ADR0(DLX_EXinst_N73509),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N72933),
    .ADR3(DLX_IDinst_Imm_0_1),
    .O(\DLX_EXinst_Mshift__n0021_Sh<8>/FROM )
  );
  defparam DLX_EXinst_Ker742211.INIT = 16'hEE22;
  X_LUT4 DLX_EXinst_Ker742211 (
    .ADR0(\DLX_EXinst_Mshift__n0021_Sh[12] ),
    .ADR1(DLX_IDinst_Imm_2_1),
    .ADR2(VCC),
    .ADR3(\DLX_EXinst_Mshift__n0021_Sh[8] ),
    .O(\DLX_EXinst_Mshift__n0021_Sh<8>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0021_Sh<8>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0021_Sh<8>/FROM ),
    .O(\DLX_EXinst_Mshift__n0021_Sh[8] )
  );
  X_BUF \DLX_EXinst_Mshift__n0021_Sh<8>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0021_Sh<8>/GROM ),
    .O(DLX_EXinst_N74223)
  );
  defparam DLX_IDinst_Mmux__n0162_inst_lut3_961.INIT = 16'hE4E4;
  X_LUT4 DLX_IDinst_Mmux__n0162_inst_lut3_961 (
    .ADR0(DLX_MEMinst_opcode_of_WB[0]),
    .ADR1(DLX_MEMinst_RF_data_in[7]),
    .ADR2(DLX_MEMinst_RF_data_in[15]),
    .ADR3(VCC),
    .O(\DLX_IDinst_RegFile_10_30/FROM )
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<30>1 .INIT = 16'h7430;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<30>1  (
    .ADR0(DLX_MEMinst_opcode_of_WB[2]),
    .ADR1(DLX_IDinst__n0161),
    .ADR2(DLX_MEMinst_RF_data_in[30]),
    .ADR3(DLX_IDinst_Mmux__n0162__net105),
    .O(\DLX_IDinst_RegFile_10_30/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_10_30/XUSED  (
    .I(\DLX_IDinst_RegFile_10_30/FROM ),
    .O(DLX_IDinst_Mmux__n0162__net105)
  );
  X_BUF \DLX_IDinst_RegFile_10_30/YUSED  (
    .I(\DLX_IDinst_RegFile_10_30/GROM ),
    .O(DLX_IDinst_WB_data_eff[30])
  );
  defparam \DLX_IDinst__n0114<30>6 .INIT = 16'hECA0;
  X_LUT4 \DLX_IDinst__n0114<30>6  (
    .ADR0(DLX_IDinst__n0098),
    .ADR1(DLX_IDinst_branch_address[30]),
    .ADR2(DLX_IDinst_EPC[30]),
    .ADR3(DLX_IDinst_N108305),
    .O(\DLX_IDinst_EPC<10>/FROM )
  );
  defparam \DLX_IDinst__n0114<10>6 .INIT = 16'hECA0;
  X_LUT4 \DLX_IDinst__n0114<10>6  (
    .ADR0(DLX_IDinst_EPC[10]),
    .ADR1(DLX_IDinst_branch_address[10]),
    .ADR2(DLX_IDinst__n0098),
    .ADR3(DLX_IDinst_N108305),
    .O(\DLX_IDinst_EPC<10>/GROM )
  );
  X_BUF \DLX_IDinst_EPC<10>/XUSED  (
    .I(\DLX_IDinst_EPC<10>/FROM ),
    .O(CHOICE2386)
  );
  X_BUF \DLX_IDinst_EPC<10>/YUSED  (
    .I(\DLX_IDinst_EPC<10>/GROM ),
    .O(CHOICE2231)
  );
  defparam \DLX_IDinst__n0114<23>6 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst__n0114<23>6  (
    .ADR0(DLX_IDinst__n0098),
    .ADR1(DLX_IDinst_EPC[23]),
    .ADR2(DLX_IDinst_branch_address[23]),
    .ADR3(DLX_IDinst_N108305),
    .O(\DLX_IDinst_EPC<11>/FROM )
  );
  defparam \DLX_IDinst__n0114<11>6 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst__n0114<11>6  (
    .ADR0(DLX_IDinst_EPC[11]),
    .ADR1(DLX_IDinst__n0098),
    .ADR2(DLX_IDinst_N108305),
    .ADR3(DLX_IDinst_branch_address[11]),
    .O(\DLX_IDinst_EPC<11>/GROM )
  );
  X_BUF \DLX_IDinst_EPC<11>/XUSED  (
    .I(\DLX_IDinst_EPC<11>/FROM ),
    .O(CHOICE2463)
  );
  X_BUF \DLX_IDinst_EPC<11>/YUSED  (
    .I(\DLX_IDinst_EPC<11>/GROM ),
    .O(CHOICE2242)
  );
  defparam \DLX_IDinst__n0114<5>6 .INIT = 16'hEAC0;
  X_LUT4 \DLX_IDinst__n0114<5>6  (
    .ADR0(DLX_IDinst__n0098),
    .ADR1(DLX_IDinst_N108305),
    .ADR2(DLX_IDinst_branch_address[5]),
    .ADR3(DLX_IDinst_EPC[5]),
    .O(\DLX_IDinst_EPC<20>/FROM )
  );
  defparam \DLX_IDinst__n0114<20>6 .INIT = 16'hEAC0;
  X_LUT4 \DLX_IDinst__n0114<20>6  (
    .ADR0(DLX_IDinst_N108305),
    .ADR1(DLX_IDinst_EPC[20]),
    .ADR2(DLX_IDinst__n0098),
    .ADR3(DLX_IDinst_branch_address[20]),
    .O(\DLX_IDinst_EPC<20>/GROM )
  );
  X_BUF \DLX_IDinst_EPC<20>/XUSED  (
    .I(\DLX_IDinst_EPC<20>/FROM ),
    .O(CHOICE2188)
  );
  X_BUF \DLX_IDinst_EPC<20>/YUSED  (
    .I(\DLX_IDinst_EPC<20>/GROM ),
    .O(CHOICE2353)
  );
  defparam \DLX_IDinst__n0114<17>6 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst__n0114<17>6  (
    .ADR0(DLX_IDinst_branch_address[17]),
    .ADR1(DLX_IDinst_N108305),
    .ADR2(DLX_IDinst__n0098),
    .ADR3(DLX_IDinst_EPC[17]),
    .O(\DLX_IDinst_EPC<12>/FROM )
  );
  defparam \DLX_IDinst__n0114<12>6 .INIT = 16'hEAC0;
  X_LUT4 \DLX_IDinst__n0114<12>6  (
    .ADR0(DLX_IDinst_N108305),
    .ADR1(DLX_IDinst__n0098),
    .ADR2(DLX_IDinst_EPC[12]),
    .ADR3(DLX_IDinst_branch_address[12]),
    .O(\DLX_IDinst_EPC<12>/GROM )
  );
  X_BUF \DLX_IDinst_EPC<12>/XUSED  (
    .I(\DLX_IDinst_EPC<12>/FROM ),
    .O(CHOICE2320)
  );
  X_BUF \DLX_IDinst_EPC<12>/YUSED  (
    .I(\DLX_IDinst_EPC<12>/GROM ),
    .O(CHOICE2253)
  );
  defparam \DLX_IDinst__n0114<27>6 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst__n0114<27>6  (
    .ADR0(DLX_IDinst_EPC[27]),
    .ADR1(DLX_IDinst__n0098),
    .ADR2(DLX_IDinst_N108305),
    .ADR3(DLX_IDinst_branch_address[27]),
    .O(\DLX_IDinst_EPC<21>/FROM )
  );
  defparam \DLX_IDinst__n0114<21>6 .INIT = 16'hECA0;
  X_LUT4 \DLX_IDinst__n0114<21>6  (
    .ADR0(DLX_IDinst__n0098),
    .ADR1(DLX_IDinst_branch_address[21]),
    .ADR2(DLX_IDinst_EPC[21]),
    .ADR3(DLX_IDinst_N108305),
    .O(\DLX_IDinst_EPC<21>/GROM )
  );
  X_BUF \DLX_IDinst_EPC<21>/XUSED  (
    .I(\DLX_IDinst_EPC<21>/FROM ),
    .O(CHOICE2419)
  );
  X_BUF \DLX_IDinst_EPC<21>/YUSED  (
    .I(\DLX_IDinst_EPC<21>/GROM ),
    .O(CHOICE2364)
  );
  defparam \DLX_IDinst__n0114<4>6 .INIT = 16'hECA0;
  X_LUT4 \DLX_IDinst__n0114<4>6  (
    .ADR0(DLX_IDinst_branch_address[4]),
    .ADR1(DLX_IDinst__n0098),
    .ADR2(DLX_IDinst_N108305),
    .ADR3(DLX_IDinst_EPC[4]),
    .O(\DLX_IDinst_EPC<13>/FROM )
  );
  defparam \DLX_IDinst__n0114<13>6 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst__n0114<13>6  (
    .ADR0(DLX_IDinst_EPC[13]),
    .ADR1(DLX_IDinst__n0098),
    .ADR2(DLX_IDinst_N108305),
    .ADR3(DLX_IDinst_branch_address[13]),
    .O(\DLX_IDinst_EPC<13>/GROM )
  );
  X_BUF \DLX_IDinst_EPC<13>/XUSED  (
    .I(\DLX_IDinst_EPC<13>/FROM ),
    .O(CHOICE2177)
  );
  X_BUF \DLX_IDinst_EPC<13>/YUSED  (
    .I(\DLX_IDinst_EPC<13>/GROM ),
    .O(CHOICE2264)
  );
  defparam \DLX_IDinst__n0114<15>6 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst__n0114<15>6  (
    .ADR0(DLX_IDinst_branch_address[15]),
    .ADR1(DLX_IDinst_N108305),
    .ADR2(DLX_IDinst__n0098),
    .ADR3(DLX_IDinst_EPC[15]),
    .O(\DLX_IDinst_EPC<22>/FROM )
  );
  defparam \DLX_IDinst__n0114<22>6 .INIT = 16'hEAC0;
  X_LUT4 \DLX_IDinst__n0114<22>6  (
    .ADR0(DLX_IDinst_EPC[22]),
    .ADR1(DLX_IDinst_N108305),
    .ADR2(DLX_IDinst_branch_address[22]),
    .ADR3(DLX_IDinst__n0098),
    .O(\DLX_IDinst_EPC<22>/GROM )
  );
  X_BUF \DLX_IDinst_EPC<22>/XUSED  (
    .I(\DLX_IDinst_EPC<22>/FROM ),
    .O(CHOICE2286)
  );
  X_BUF \DLX_IDinst_EPC<22>/YUSED  (
    .I(\DLX_IDinst_EPC<22>/GROM ),
    .O(CHOICE2375)
  );
  defparam \DLX_IDinst__n0114<24>6 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst__n0114<24>6  (
    .ADR0(DLX_IDinst__n0098),
    .ADR1(DLX_IDinst_EPC[24]),
    .ADR2(DLX_IDinst_branch_address[24]),
    .ADR3(DLX_IDinst_N108305),
    .O(\DLX_IDinst_EPC<14>/FROM )
  );
  defparam \DLX_IDinst__n0114<14>6 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst__n0114<14>6  (
    .ADR0(DLX_IDinst_branch_address[14]),
    .ADR1(DLX_IDinst_N108305),
    .ADR2(DLX_IDinst_EPC[14]),
    .ADR3(DLX_IDinst__n0098),
    .O(\DLX_IDinst_EPC<14>/GROM )
  );
  X_BUF \DLX_IDinst_EPC<14>/XUSED  (
    .I(\DLX_IDinst_EPC<14>/FROM ),
    .O(CHOICE2452)
  );
  X_BUF \DLX_IDinst_EPC<14>/YUSED  (
    .I(\DLX_IDinst_EPC<14>/GROM ),
    .O(CHOICE2275)
  );
  defparam \DLX_IDinst__n0114<31>5 .INIT = 16'hFF88;
  X_LUT4 \DLX_IDinst__n0114<31>5  (
    .ADR0(DLX_IDinst__n0098),
    .ADR1(DLX_IDinst_EPC[31]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst__n0453),
    .O(\DLX_IDinst_EPC<31>/FROM )
  );
  defparam \DLX_IDinst__n0114<31>13 .INIT = 16'h5540;
  X_LUT4 \DLX_IDinst__n0114<31>13  (
    .ADR0(DLX_IDinst_N108456),
    .ADR1(DLX_IDinst_branch_address[31]),
    .ADR2(DLX_IDinst_N108305),
    .ADR3(CHOICE3171),
    .O(\DLX_IDinst_EPC<31>/GROM )
  );
  X_BUF \DLX_IDinst_EPC<31>/XUSED  (
    .I(\DLX_IDinst_EPC<31>/FROM ),
    .O(CHOICE3171)
  );
  X_BUF \DLX_IDinst_EPC<31>/YUSED  (
    .I(\DLX_IDinst_EPC<31>/GROM ),
    .O(CHOICE3173)
  );
  defparam \DLX_IDinst__n0114<0>6 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst__n0114<0>6  (
    .ADR0(DLX_IDinst__n0098),
    .ADR1(DLX_IDinst_EPC[0]),
    .ADR2(DLX_IDinst_N108305),
    .ADR3(DLX_IDinst_branch_address[0]),
    .O(\DLX_IDinst_EPC<16>/FROM )
  );
  defparam \DLX_IDinst__n0114<16>6 .INIT = 16'hECA0;
  X_LUT4 \DLX_IDinst__n0114<16>6  (
    .ADR0(DLX_IDinst_branch_address[16]),
    .ADR1(DLX_IDinst__n0098),
    .ADR2(DLX_IDinst_N108305),
    .ADR3(DLX_IDinst_EPC[16]),
    .O(\DLX_IDinst_EPC<16>/GROM )
  );
  X_BUF \DLX_IDinst_EPC<16>/XUSED  (
    .I(\DLX_IDinst_EPC<16>/FROM ),
    .O(CHOICE3156)
  );
  X_BUF \DLX_IDinst_EPC<16>/YUSED  (
    .I(\DLX_IDinst_EPC<16>/GROM ),
    .O(CHOICE2309)
  );
  defparam \DLX_IDinst__n0114<3>6 .INIT = 16'hECA0;
  X_LUT4 \DLX_IDinst__n0114<3>6  (
    .ADR0(DLX_IDinst_N108305),
    .ADR1(DLX_IDinst__n0098),
    .ADR2(DLX_IDinst_branch_address[3]),
    .ADR3(DLX_IDinst_EPC[3]),
    .O(\DLX_IDinst_EPC<25>/FROM )
  );
  defparam \DLX_IDinst__n0114<25>6 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst__n0114<25>6  (
    .ADR0(DLX_IDinst_N108305),
    .ADR1(DLX_IDinst_branch_address[25]),
    .ADR2(DLX_IDinst_EPC[25]),
    .ADR3(DLX_IDinst__n0098),
    .O(\DLX_IDinst_EPC<25>/GROM )
  );
  X_BUF \DLX_IDinst_EPC<25>/XUSED  (
    .I(\DLX_IDinst_EPC<25>/FROM ),
    .O(CHOICE2166)
  );
  X_BUF \DLX_IDinst_EPC<25>/YUSED  (
    .I(\DLX_IDinst_EPC<25>/GROM ),
    .O(CHOICE2441)
  );
  defparam \DLX_IDinst__n0114<29>6 .INIT = 16'hEAC0;
  X_LUT4 \DLX_IDinst__n0114<29>6  (
    .ADR0(DLX_IDinst_EPC[29]),
    .ADR1(DLX_IDinst_N108305),
    .ADR2(DLX_IDinst_branch_address[29]),
    .ADR3(DLX_IDinst__n0098),
    .O(\DLX_IDinst_EPC<18>/FROM )
  );
  defparam \DLX_IDinst__n0114<18>6 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst__n0114<18>6  (
    .ADR0(DLX_IDinst__n0098),
    .ADR1(DLX_IDinst_EPC[18]),
    .ADR2(DLX_IDinst_N108305),
    .ADR3(DLX_IDinst_branch_address[18]),
    .O(\DLX_IDinst_EPC<18>/GROM )
  );
  X_BUF \DLX_IDinst_EPC<18>/XUSED  (
    .I(\DLX_IDinst_EPC<18>/FROM ),
    .O(CHOICE2397)
  );
  X_BUF \DLX_IDinst_EPC<18>/YUSED  (
    .I(\DLX_IDinst_EPC<18>/GROM ),
    .O(CHOICE2331)
  );
  defparam \DLX_IDinst__n0114<9>6 .INIT = 16'hEAC0;
  X_LUT4 \DLX_IDinst__n0114<9>6  (
    .ADR0(DLX_IDinst_branch_address[9]),
    .ADR1(DLX_IDinst_EPC[9]),
    .ADR2(DLX_IDinst__n0098),
    .ADR3(DLX_IDinst_N108305),
    .O(\DLX_IDinst_EPC<19>/FROM )
  );
  defparam \DLX_IDinst__n0114<19>6 .INIT = 16'hEAC0;
  X_LUT4 \DLX_IDinst__n0114<19>6  (
    .ADR0(DLX_IDinst_branch_address[19]),
    .ADR1(DLX_IDinst_EPC[19]),
    .ADR2(DLX_IDinst__n0098),
    .ADR3(DLX_IDinst_N108305),
    .O(\DLX_IDinst_EPC<19>/GROM )
  );
  X_BUF \DLX_IDinst_EPC<19>/XUSED  (
    .I(\DLX_IDinst_EPC<19>/FROM ),
    .O(CHOICE2220)
  );
  X_BUF \DLX_IDinst_EPC<19>/YUSED  (
    .I(\DLX_IDinst_EPC<19>/GROM ),
    .O(CHOICE2342)
  );
  defparam \DLX_IDinst__n0114<2>6 .INIT = 16'hEAC0;
  X_LUT4 \DLX_IDinst__n0114<2>6  (
    .ADR0(DLX_IDinst_branch_address[2]),
    .ADR1(DLX_IDinst_EPC[2]),
    .ADR2(DLX_IDinst__n0098),
    .ADR3(DLX_IDinst_N108305),
    .O(\DLX_IDinst_EPC<28>/FROM )
  );
  defparam \DLX_IDinst__n0114<28>6 .INIT = 16'hECA0;
  X_LUT4 \DLX_IDinst__n0114<28>6  (
    .ADR0(DLX_IDinst_EPC[28]),
    .ADR1(DLX_IDinst_branch_address[28]),
    .ADR2(DLX_IDinst__n0098),
    .ADR3(DLX_IDinst_N108305),
    .O(\DLX_IDinst_EPC<28>/GROM )
  );
  X_BUF \DLX_IDinst_EPC<28>/XUSED  (
    .I(\DLX_IDinst_EPC<28>/FROM ),
    .O(CHOICE2155)
  );
  X_BUF \DLX_IDinst_EPC<28>/YUSED  (
    .I(\DLX_IDinst_EPC<28>/GROM ),
    .O(CHOICE2408)
  );
  defparam \DLX_EXinst__n0007<21>131_SW0 .INIT = 16'hFFFA;
  X_LUT4 \DLX_EXinst__n0007<21>131_SW0  (
    .ADR0(CHOICE4125),
    .ADR1(VCC),
    .ADR2(CHOICE4140),
    .ADR3(CHOICE4149),
    .O(\N163680/FROM )
  );
  defparam \DLX_EXinst__n0007<21>131 .INIT = 16'h0F08;
  X_LUT4 \DLX_EXinst__n0007<21>131  (
    .ADR0(CHOICE4135),
    .ADR1(DLX_EXinst_N76318),
    .ADR2(DLX_EXinst__n0036),
    .ADR3(N163680),
    .O(\N163680/GROM )
  );
  X_BUF \N163680/XUSED  (
    .I(\N163680/FROM ),
    .O(N163680)
  );
  X_BUF \N163680/YUSED  (
    .I(\N163680/GROM ),
    .O(CHOICE4153)
  );
  defparam DLX_IDinst_RegFile_27_26_1466.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_27_26_1466 (
    .I(DLX_IDinst_WB_data_eff[26]),
    .CE(DLX_IDinst__n0604),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_27_26)
  );
  defparam \DLX_IDinst__n0146<22>36_SW0 .INIT = 16'hBB5F;
  X_LUT4 \DLX_IDinst__n0146<22>36_SW0  (
    .ADR0(DLX_IDinst_jtarget[22]),
    .ADR1(\DLX_IDinst_Cause_Reg[31] ),
    .ADR2(DLX_IDinst_EPC[22]),
    .ADR3(DLX_IDinst_jtarget[21]),
    .O(\N163700/FROM )
  );
  defparam \DLX_IDinst__n0146<22>36 .INIT = 16'hC0EA;
  X_LUT4 \DLX_IDinst__n0146<22>36  (
    .ADR0(DLX_IDinst_N107105),
    .ADR1(N134590),
    .ADR2(\DLX_IDinst_regA_eff[22] ),
    .ADR3(N163700),
    .O(\N163700/GROM )
  );
  X_BUF \N163700/XUSED  (
    .I(\N163700/FROM ),
    .O(N163700)
  );
  X_BUF \N163700/YUSED  (
    .I(\N163700/GROM ),
    .O(CHOICE2753)
  );
  defparam \DLX_IDinst__n0146<30>36_SW0 .INIT = 16'h9BDF;
  X_LUT4 \DLX_IDinst__n0146<30>36_SW0  (
    .ADR0(DLX_IDinst_jtarget[21]),
    .ADR1(DLX_IDinst_jtarget[22]),
    .ADR2(\DLX_IDinst_Cause_Reg[31] ),
    .ADR3(DLX_IDinst_EPC[30]),
    .O(\N163325/FROM )
  );
  defparam \DLX_IDinst__n0146<30>36 .INIT = 16'h88F8;
  X_LUT4 \DLX_IDinst__n0146<30>36  (
    .ADR0(\DLX_IDinst_regA_eff[30] ),
    .ADR1(N134590),
    .ADR2(DLX_IDinst_N107105),
    .ADR3(N163325),
    .O(\N163325/GROM )
  );
  X_BUF \N163325/XUSED  (
    .I(\N163325/FROM ),
    .O(N163325)
  );
  X_BUF \N163325/YUSED  (
    .I(\N163325/GROM ),
    .O(CHOICE2873)
  );
  defparam vga_top_vga1_Ker1129021.INIT = 16'h0004;
  X_LUT4 vga_top_vga1_Ker1129021 (
    .ADR0(vga_top_vga1_hcounter[7]),
    .ADR1(vga_top_vga1_N112926),
    .ADR2(vga_top_vga1_hcounter[4]),
    .ADR3(vga_top_vga1_hcounter[1]),
    .O(\vga_top_vga1_N112904/FROM )
  );
  defparam vga_top_vga1_Ker1129341.INIT = 16'hA000;
  X_LUT4 vga_top_vga1_Ker1129341 (
    .ADR0(vga_top_vga1_hcounter[5]),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_hcounter[2]),
    .ADR3(vga_top_vga1_N112904),
    .O(\vga_top_vga1_N112904/GROM )
  );
  X_BUF \vga_top_vga1_N112904/XUSED  (
    .I(\vga_top_vga1_N112904/FROM ),
    .O(vga_top_vga1_N112904)
  );
  X_BUF \vga_top_vga1_N112904/YUSED  (
    .I(\vga_top_vga1_N112904/GROM ),
    .O(vga_top_vga1_N112936)
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<0>1 .INIT = 16'h1010;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<0>1  (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(DLX_IDinst_reg_out_A[0]),
    .ADR3(VCC),
    .O(\DLX_EXinst_Mshift__n0023_Sh<0>/FROM )
  );
  defparam \DLX_EXinst__n0007<16>44 .INIT = 16'hF4F0;
  X_LUT4 \DLX_EXinst__n0007<16>44  (
    .ADR0(DLX_EXinst_N72822),
    .ADR1(DLX_IDinst_reg_out_B[4]),
    .ADR2(CHOICE4573),
    .ADR3(\DLX_EXinst_Mshift__n0023_Sh[0] ),
    .O(\DLX_EXinst_Mshift__n0023_Sh<0>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0023_Sh<0>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0023_Sh<0>/FROM ),
    .O(\DLX_EXinst_Mshift__n0023_Sh[0] )
  );
  X_BUF \DLX_EXinst_Mshift__n0023_Sh<0>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0023_Sh<0>/GROM ),
    .O(CHOICE4574)
  );
  defparam vga_top_vga1_Ker1129081.INIT = 16'h1100;
  X_LUT4 vga_top_vga1_Ker1129081 (
    .ADR0(vga_top_vga1_vcounter[4]),
    .ADR1(vga_top_vga1_vcounter[5]),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_N112941),
    .O(\vga_top_vga1_N112910/FROM )
  );
  defparam vga_top_vga1__n000819.INIT = 16'h7F00;
  X_LUT4 vga_top_vga1__n000819 (
    .ADR0(vga_top_vga1_vcounter[1]),
    .ADR1(vga_top_vga1_vcounter[2]),
    .ADR2(vga_top_vga1_vcounter[3]),
    .ADR3(vga_top_vga1_N112910),
    .O(\vga_top_vga1_N112910/GROM )
  );
  X_BUF \vga_top_vga1_N112910/XUSED  (
    .I(\vga_top_vga1_N112910/FROM ),
    .O(vga_top_vga1_N112910)
  );
  X_BUF \vga_top_vga1_N112910/YUSED  (
    .I(\vga_top_vga1_N112910/GROM ),
    .O(CHOICE3146)
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<1>1 .INIT = 16'h00E4;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<1>1  (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(DLX_IDinst_reg_out_A[1]),
    .ADR2(DLX_IDinst_reg_out_A[0]),
    .ADR3(DLX_IDinst_reg_out_B[1]),
    .O(\DLX_EXinst_Mshift__n0023_Sh<1>/FROM )
  );
  defparam \DLX_EXinst__n0007<17>367_SW0 .INIT = 16'hF4F0;
  X_LUT4 \DLX_EXinst__n0007<17>367_SW0  (
    .ADR0(DLX_EXinst_N72822),
    .ADR1(DLX_EXinst_N75973),
    .ADR2(CHOICE5424),
    .ADR3(\DLX_EXinst_Mshift__n0023_Sh[1] ),
    .O(\DLX_EXinst_Mshift__n0023_Sh<1>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0023_Sh<1>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0023_Sh<1>/FROM ),
    .O(\DLX_EXinst_Mshift__n0023_Sh[1] )
  );
  X_BUF \DLX_EXinst_Mshift__n0023_Sh<1>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0023_Sh<1>/GROM ),
    .O(N163584)
  );
  defparam vga_top_vga1_Ker1129191.INIT = 16'h0003;
  X_LUT4 vga_top_vga1_Ker1129191 (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_vcounter[3]),
    .ADR2(vga_top_vga1_vcounter[4]),
    .ADR3(vga_top_vga1_vcounter[2]),
    .O(\vga_top_vga1_N112921/FROM )
  );
  defparam vga_top_vga1__n000954.INIT = 16'h1311;
  X_LUT4 vga_top_vga1__n000954 (
    .ADR0(vga_top_vga1_vcounter[5]),
    .ADR1(vga_top_vga1_vcounter[9]),
    .ADR2(vga_top_vga1_vcounter[1]),
    .ADR3(vga_top_vga1_N112921),
    .O(\vga_top_vga1_N112921/GROM )
  );
  X_BUF \vga_top_vga1_N112921/XUSED  (
    .I(\vga_top_vga1_N112921/FROM ),
    .O(vga_top_vga1_N112921)
  );
  X_BUF \vga_top_vga1_N112921/YUSED  (
    .I(\vga_top_vga1_N112921/GROM ),
    .O(CHOICE3468)
  );
  defparam vga_top_vga1_Ker1129441.INIT = 16'h0001;
  X_LUT4 vga_top_vga1_Ker1129441 (
    .ADR0(vga_top_vga1_hcounter[3]),
    .ADR1(vga_top_vga1_hcounter[2]),
    .ADR2(vga_top_vga1_hcounter[8]),
    .ADR3(vga_top_vga1_hcounter[0]),
    .O(\vga_top_vga1_N112946/FROM )
  );
  defparam vga_top_vga1__n000835.INIT = 16'hAA00;
  X_LUT4 vga_top_vga1__n000835 (
    .ADR0(vga_top_vga1_N112926),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_N112946),
    .O(\vga_top_vga1_N112946/GROM )
  );
  X_BUF \vga_top_vga1_N112946/XUSED  (
    .I(\vga_top_vga1_N112946/FROM ),
    .O(vga_top_vga1_N112946)
  );
  X_BUF \vga_top_vga1_N112946/YUSED  (
    .I(\vga_top_vga1_N112946/GROM ),
    .O(CHOICE3149)
  );
  defparam vga_top_vga1_Ker1129391.INIT = 16'h0011;
  X_LUT4 vga_top_vga1_Ker1129391 (
    .ADR0(vga_top_vga1_vcounter[6]),
    .ADR1(vga_top_vga1_vcounter[7]),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_vcounter[8]),
    .O(\vga_top_vga1_N112941/GROM )
  );
  X_BUF \vga_top_vga1_N112941/YUSED  (
    .I(\vga_top_vga1_N112941/GROM ),
    .O(vga_top_vga1_N112941)
  );
  defparam \DLX_IDinst__n0146<23>36_SW0 .INIT = 16'hF53F;
  X_LUT4 \DLX_IDinst__n0146<23>36_SW0  (
    .ADR0(\DLX_IDinst_Cause_Reg[31] ),
    .ADR1(DLX_IDinst_EPC[23]),
    .ADR2(DLX_IDinst_jtarget[22]),
    .ADR3(DLX_IDinst_jtarget[21]),
    .O(\N163510/FROM )
  );
  defparam \DLX_IDinst__n0146<23>36 .INIT = 16'h88F8;
  X_LUT4 \DLX_IDinst__n0146<23>36  (
    .ADR0(\DLX_IDinst_regA_eff[23] ),
    .ADR1(N134590),
    .ADR2(DLX_IDinst_N107105),
    .ADR3(N163510),
    .O(\N163510/GROM )
  );
  X_BUF \N163510/XUSED  (
    .I(\N163510/FROM ),
    .O(N163510)
  );
  X_BUF \N163510/YUSED  (
    .I(\N163510/GROM ),
    .O(CHOICE2768)
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<7>1 .INIT = 16'hF5A0;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<7>1  (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N73599),
    .ADR3(DLX_EXinst_N72848),
    .O(\DLX_EXinst_Mshift__n0023_Sh<7>/FROM )
  );
  defparam DLX_EXinst_Ker729111.INIT = 16'hAFA0;
  X_LUT4 DLX_EXinst_Ker729111 (
    .ADR0(\DLX_EXinst_Mshift__n0023_Sh[3] ),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[2]),
    .ADR3(\DLX_EXinst_Mshift__n0023_Sh[7] ),
    .O(\DLX_EXinst_Mshift__n0023_Sh<7>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0023_Sh<7>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0023_Sh<7>/FROM ),
    .O(\DLX_EXinst_Mshift__n0023_Sh[7] )
  );
  X_BUF \DLX_EXinst_Mshift__n0023_Sh<7>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0023_Sh<7>/GROM ),
    .O(DLX_EXinst_N72913)
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<8>1 .INIT = 16'hFC0C;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<8>1  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N73604),
    .ADR2(DLX_IDinst_reg_out_B[0]),
    .ADR3(DLX_EXinst_N72848),
    .O(\DLX_EXinst_Mshift__n0023_Sh<8>/FROM )
  );
  defparam DLX_EXinst_Ker740491.INIT = 16'hEE44;
  X_LUT4 DLX_EXinst_Ker740491 (
    .ADR0(DLX_IDinst_reg_out_B[2]),
    .ADR1(\DLX_EXinst_Mshift__n0023_Sh[12] ),
    .ADR2(VCC),
    .ADR3(\DLX_EXinst_Mshift__n0023_Sh[8] ),
    .O(\DLX_EXinst_Mshift__n0023_Sh<8>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0023_Sh<8>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0023_Sh<8>/FROM ),
    .O(\DLX_EXinst_Mshift__n0023_Sh[8] )
  );
  X_BUF \DLX_EXinst_Mshift__n0023_Sh<8>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0023_Sh<8>/GROM ),
    .O(DLX_EXinst_N74051)
  );
  defparam DLX_EXinst_Ker730211.INIT = 16'hEE44;
  X_LUT4 DLX_EXinst_Ker730211 (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(DLX_IDinst_reg_out_A[5]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[7]),
    .O(\DLX_EXinst_N73023/FROM )
  );
  defparam DLX_EXinst_Ker7443439_SW0.INIT = 16'hD800;
  X_LUT4 DLX_EXinst_Ker7443439_SW0 (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(DLX_IDinst_reg_out_A[7]),
    .ADR2(DLX_IDinst_reg_out_A[5]),
    .ADR3(DLX_IDinst_reg_out_B[0]),
    .O(\DLX_EXinst_N73023/GROM )
  );
  X_BUF \DLX_EXinst_N73023/XUSED  (
    .I(\DLX_EXinst_N73023/FROM ),
    .O(DLX_EXinst_N73023)
  );
  X_BUF \DLX_EXinst_N73023/YUSED  (
    .I(\DLX_EXinst_N73023/GROM ),
    .O(N163136)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_cy_261_1467.INIT = 16'hDD44;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_cy_261_1467 (
    .ADR0(DLX_IDinst_reg_out_B[31]),
    .ADR1(DLX_IDinst_reg_out_A[31]),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_Mcompar__n0095_inst_cy_260),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_261/FROM )
  );
  defparam \DLX_EXinst__n0007<0>242 .INIT = 16'h20E0;
  X_LUT4 \DLX_EXinst__n0007<0>242  (
    .ADR0(DLX_EXinst__n0087),
    .ADR1(\DLX_IDinst_Imm[2] ),
    .ADR2(\DLX_IDinst_Imm[0] ),
    .ADR3(DLX_EXinst_Mcompar__n0095_inst_cy_261),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_261/GROM )
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_261/XUSED  (
    .I(\DLX_EXinst_Mcompar__n0095_inst_cy_261/FROM ),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_261)
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_261/YUSED  (
    .I(\DLX_EXinst_Mcompar__n0095_inst_cy_261/GROM ),
    .O(CHOICE5923)
  );
  defparam \DLX_EXinst__n0007<21>272_SW0 .INIT = 16'hFF08;
  X_LUT4 \DLX_EXinst__n0007<21>272_SW0  (
    .ADR0(CHOICE4167),
    .ADR1(DLX_EXinst__n0080),
    .ADR2(N148323),
    .ADR3(CHOICE4181),
    .O(\N163639/GROM )
  );
  X_BUF \N163639/YUSED  (
    .I(\N163639/GROM ),
    .O(N163639)
  );
  defparam \DLX_IDinst__n0114<0>37 .INIT = 16'hCCDC;
  X_LUT4 \DLX_IDinst__n0114<0>37  (
    .ADR0(DLX_IDinst__n0453),
    .ADR1(CHOICE3164),
    .ADR2(CHOICE3156),
    .ADR3(DLX_IDinst_N108456),
    .O(\DLX_IDinst_branch_address<0>/FROM )
  );
  defparam \DLX_IDinst__n0114<0>47 .INIT = 16'hFFA0;
  X_LUT4 \DLX_IDinst__n0114<0>47  (
    .ADR0(N137082),
    .ADR1(VCC),
    .ADR2(DLX_IDinst__n0157[0]),
    .ADR3(CHOICE3165),
    .O(N145826)
  );
  X_BUF \DLX_IDinst_branch_address<0>/XUSED  (
    .I(\DLX_IDinst_branch_address<0>/FROM ),
    .O(CHOICE3165)
  );
  defparam \DLX_IDinst__n0114<1>25 .INIT = 16'hAAAE;
  X_LUT4 \DLX_IDinst__n0114<1>25  (
    .ADR0(CHOICE2148),
    .ADR1(CHOICE2144),
    .ADR2(DLX_IDinst__n0453),
    .ADR3(DLX_IDinst_N108456),
    .O(\DLX_IDinst_branch_address<1>/FROM )
  );
  defparam \DLX_IDinst__n0114<1>31 .INIT = 16'hFFA0;
  X_LUT4 \DLX_IDinst__n0114<1>31  (
    .ADR0(N137082),
    .ADR1(VCC),
    .ADR2(DLX_IDinst__n0157[1]),
    .ADR3(CHOICE2149),
    .O(N139826)
  );
  X_BUF \DLX_IDinst_branch_address<1>/XUSED  (
    .I(\DLX_IDinst_branch_address<1>/FROM ),
    .O(CHOICE2149)
  );
  defparam \DLX_IDinst__n0114<2>25 .INIT = 16'hFF10;
  X_LUT4 \DLX_IDinst__n0114<2>25  (
    .ADR0(DLX_IDinst__n0453),
    .ADR1(DLX_IDinst_N108456),
    .ADR2(CHOICE2155),
    .ADR3(CHOICE2159),
    .O(\DLX_IDinst_branch_address<2>/FROM )
  );
  defparam \DLX_IDinst__n0114<2>31 .INIT = 16'hFFA0;
  X_LUT4 \DLX_IDinst__n0114<2>31  (
    .ADR0(DLX_IDinst__n0157[2]),
    .ADR1(VCC),
    .ADR2(N137082),
    .ADR3(CHOICE2160),
    .O(N139889)
  );
  X_BUF \DLX_IDinst_branch_address<2>/XUSED  (
    .I(\DLX_IDinst_branch_address<2>/FROM ),
    .O(CHOICE2160)
  );
  defparam \DLX_EXinst__n0007<22>131_SW0 .INIT = 16'hFFFC;
  X_LUT4 \DLX_EXinst__n0007<22>131_SW0  (
    .ADR0(VCC),
    .ADR1(CHOICE4084),
    .ADR2(CHOICE4075),
    .ADR3(CHOICE4060),
    .O(\N163278/FROM )
  );
  defparam \DLX_EXinst__n0007<22>131 .INIT = 16'h5540;
  X_LUT4 \DLX_EXinst__n0007<22>131  (
    .ADR0(DLX_EXinst__n0036),
    .ADR1(CHOICE4070),
    .ADR2(DLX_EXinst_N76318),
    .ADR3(N163278),
    .O(\N163278/GROM )
  );
  X_BUF \N163278/XUSED  (
    .I(\N163278/FROM ),
    .O(N163278)
  );
  X_BUF \N163278/YUSED  (
    .I(\N163278/GROM ),
    .O(CHOICE4088)
  );
  defparam \DLX_EXinst_Mshift__n0024_Sh<50> .INIT = 16'hFC30;
  X_LUT4 \DLX_EXinst_Mshift__n0024_Sh<50>  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_B_2_1),
    .ADR2(DLX_EXinst_N74731),
    .ADR3(N131027),
    .O(\DLX_EXinst_Mshift__n0024_Sh<50>/FROM )
  );
  defparam \DLX_EXinst__n0007<18>298_SW0 .INIT = 16'hEEAA;
  X_LUT4 \DLX_EXinst__n0007<18>298_SW0  (
    .ADR0(CHOICE5258),
    .ADR1(DLX_EXinst__n0081),
    .ADR2(VCC),
    .ADR3(\DLX_EXinst_Mshift__n0024_Sh[50] ),
    .O(\DLX_EXinst_Mshift__n0024_Sh<50>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0024_Sh<50>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0024_Sh<50>/FROM ),
    .O(\DLX_EXinst_Mshift__n0024_Sh[50] )
  );
  X_BUF \DLX_EXinst_Mshift__n0024_Sh<50>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0024_Sh<50>/GROM ),
    .O(N163302)
  );
  defparam \DLX_IDinst__n0114<3>25 .INIT = 16'hFF10;
  X_LUT4 \DLX_IDinst__n0114<3>25  (
    .ADR0(DLX_IDinst_N108456),
    .ADR1(DLX_IDinst__n0453),
    .ADR2(CHOICE2166),
    .ADR3(CHOICE2170),
    .O(\DLX_IDinst_branch_address<3>/FROM )
  );
  defparam \DLX_IDinst__n0114<3>31 .INIT = 16'hFF88;
  X_LUT4 \DLX_IDinst__n0114<3>31  (
    .ADR0(DLX_IDinst__n0157[3]),
    .ADR1(N137082),
    .ADR2(VCC),
    .ADR3(CHOICE2171),
    .O(N139952)
  );
  X_BUF \DLX_IDinst_branch_address<3>/XUSED  (
    .I(\DLX_IDinst_branch_address<3>/FROM ),
    .O(CHOICE2171)
  );
  defparam DLX_IDinst_RegFile_28_10_1468.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_28_10_1468 (
    .I(DLX_IDinst_WB_data_eff[10]),
    .CE(DLX_IDinst__n0606),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_28_10)
  );
  defparam \DLX_IDinst__n0114<4>25 .INIT = 16'hCCCE;
  X_LUT4 \DLX_IDinst__n0114<4>25  (
    .ADR0(CHOICE2177),
    .ADR1(CHOICE2181),
    .ADR2(DLX_IDinst_N108456),
    .ADR3(DLX_IDinst__n0453),
    .O(\DLX_IDinst_branch_address<4>/FROM )
  );
  defparam \DLX_IDinst__n0114<4>31 .INIT = 16'hFFA0;
  X_LUT4 \DLX_IDinst__n0114<4>31  (
    .ADR0(DLX_IDinst__n0157[4]),
    .ADR1(VCC),
    .ADR2(N137082),
    .ADR3(CHOICE2182),
    .O(N140015)
  );
  X_BUF \DLX_IDinst_branch_address<4>/XUSED  (
    .I(\DLX_IDinst_branch_address<4>/FROM ),
    .O(CHOICE2182)
  );
  defparam \DLX_IDinst__n0146<16>36_SW0 .INIT = 16'h9DBF;
  X_LUT4 \DLX_IDinst__n0146<16>36_SW0  (
    .ADR0(DLX_IDinst_jtarget[21]),
    .ADR1(DLX_IDinst_jtarget[22]),
    .ADR2(DLX_IDinst_EPC[16]),
    .ADR3(\DLX_IDinst_Cause_Reg[31] ),
    .O(\N163447/FROM )
  );
  defparam \DLX_IDinst__n0146<16>36 .INIT = 16'h8F88;
  X_LUT4 \DLX_IDinst__n0146<16>36  (
    .ADR0(\DLX_IDinst_regA_eff[16] ),
    .ADR1(N134590),
    .ADR2(N163447),
    .ADR3(DLX_IDinst_N107105),
    .O(\N163447/GROM )
  );
  X_BUF \N163447/XUSED  (
    .I(\N163447/FROM ),
    .O(N163447)
  );
  X_BUF \N163447/YUSED  (
    .I(\N163447/GROM ),
    .O(CHOICE2663)
  );
  defparam \DLX_IDinst__n0146<24>36_SW0 .INIT = 16'h9BDF;
  X_LUT4 \DLX_IDinst__n0146<24>36_SW0  (
    .ADR0(DLX_IDinst_jtarget[22]),
    .ADR1(DLX_IDinst_jtarget[21]),
    .ADR2(DLX_IDinst_EPC[24]),
    .ADR3(\DLX_IDinst_Cause_Reg[31] ),
    .O(\N163262/FROM )
  );
  defparam \DLX_IDinst__n0146<24>36 .INIT = 16'h88F8;
  X_LUT4 \DLX_IDinst__n0146<24>36  (
    .ADR0(\DLX_IDinst_regA_eff[24] ),
    .ADR1(N134590),
    .ADR2(DLX_IDinst_N107105),
    .ADR3(N163262),
    .O(\N163262/GROM )
  );
  X_BUF \N163262/XUSED  (
    .I(\N163262/FROM ),
    .O(N163262)
  );
  X_BUF \N163262/YUSED  (
    .I(\N163262/GROM ),
    .O(CHOICE2783)
  );
  defparam DLX_IDinst_RegFile_27_18_1469.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_27_18_1469 (
    .I(DLX_IDinst_WB_data_eff[18]),
    .CE(DLX_IDinst__n0604),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_27_18)
  );
  defparam \DLX_IDinst__n0114<5>25 .INIT = 16'hF0F2;
  X_LUT4 \DLX_IDinst__n0114<5>25  (
    .ADR0(CHOICE2188),
    .ADR1(DLX_IDinst__n0453),
    .ADR2(CHOICE2192),
    .ADR3(DLX_IDinst_N108456),
    .O(\DLX_IDinst_EPC<0>/FROM )
  );
  defparam \DLX_IDinst__n0114<5>31 .INIT = 16'hFF88;
  X_LUT4 \DLX_IDinst__n0114<5>31  (
    .ADR0(DLX_IDinst__n0157[5]),
    .ADR1(N137082),
    .ADR2(VCC),
    .ADR3(CHOICE2193),
    .O(N140078)
  );
  X_BUF \DLX_IDinst_EPC<0>/XUSED  (
    .I(\DLX_IDinst_EPC<0>/FROM ),
    .O(CHOICE2193)
  );
  defparam \DLX_IDinst__n0114<6>37 .INIT = 16'hF0F2;
  X_LUT4 \DLX_IDinst__n0114<6>37  (
    .ADR0(CHOICE3185),
    .ADR1(DLX_IDinst__n0453),
    .ADR2(CHOICE3193),
    .ADR3(DLX_IDinst_N108456),
    .O(\DLX_IDinst_branch_address<6>/FROM )
  );
  defparam \DLX_IDinst__n0114<6>47 .INIT = 16'hFF88;
  X_LUT4 \DLX_IDinst__n0114<6>47  (
    .ADR0(N137082),
    .ADR1(DLX_IDinst__n0157[6]),
    .ADR2(VCC),
    .ADR3(CHOICE3194),
    .O(N145997)
  );
  X_BUF \DLX_IDinst_branch_address<6>/XUSED  (
    .I(\DLX_IDinst_branch_address<6>/FROM ),
    .O(CHOICE3194)
  );
  defparam \DLX_IDinst__n0114<7>19 .INIT = 16'hECA0;
  X_LUT4 \DLX_IDinst__n0114<7>19  (
    .ADR0(DLX_IDinst__n0157[7]),
    .ADR1(DLX_IDinst_N107870),
    .ADR2(DLX_IDinst_N107609),
    .ADR3(\DLX_IDinst_regA_eff[7] ),
    .O(\DLX_IDinst_branch_address<7>/FROM )
  );
  defparam \DLX_IDinst__n0114<7>20 .INIT = 16'hFFF0;
  X_LUT4 \DLX_IDinst__n0114<7>20  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(CHOICE2200),
    .ADR3(CHOICE2203),
    .O(N140126)
  );
  X_BUF \DLX_IDinst_branch_address<7>/XUSED  (
    .I(\DLX_IDinst_branch_address<7>/FROM ),
    .O(CHOICE2203)
  );
  defparam \DLX_IDinst__n0114<8>25 .INIT = 16'hF0F2;
  X_LUT4 \DLX_IDinst__n0114<8>25  (
    .ADR0(CHOICE2209),
    .ADR1(DLX_IDinst__n0453),
    .ADR2(CHOICE2213),
    .ADR3(DLX_IDinst_N108456),
    .O(\DLX_IDinst_branch_address<8>/FROM )
  );
  defparam \DLX_IDinst__n0114<8>31 .INIT = 16'hFF88;
  X_LUT4 \DLX_IDinst__n0114<8>31  (
    .ADR0(DLX_IDinst__n0157[8]),
    .ADR1(N137082),
    .ADR2(VCC),
    .ADR3(CHOICE2214),
    .O(N140193)
  );
  X_BUF \DLX_IDinst_branch_address<8>/XUSED  (
    .I(\DLX_IDinst_branch_address<8>/FROM ),
    .O(CHOICE2214)
  );
  defparam \DLX_IDinst__n0114<9>25 .INIT = 16'hF1F0;
  X_LUT4 \DLX_IDinst__n0114<9>25  (
    .ADR0(DLX_IDinst_N108456),
    .ADR1(DLX_IDinst__n0453),
    .ADR2(CHOICE2224),
    .ADR3(CHOICE2220),
    .O(\DLX_IDinst_branch_address<9>/FROM )
  );
  defparam \DLX_IDinst__n0114<9>31 .INIT = 16'hFFA0;
  X_LUT4 \DLX_IDinst__n0114<9>31  (
    .ADR0(N137082),
    .ADR1(VCC),
    .ADR2(DLX_IDinst__n0157[9]),
    .ADR3(CHOICE2225),
    .O(N140256)
  );
  X_BUF \DLX_IDinst_branch_address<9>/XUSED  (
    .I(\DLX_IDinst_branch_address<9>/FROM ),
    .O(CHOICE2225)
  );
  defparam \DLX_IDinst__n0146<25>36_SW0 .INIT = 16'hDD3F;
  X_LUT4 \DLX_IDinst__n0146<25>36_SW0  (
    .ADR0(\DLX_IDinst_Cause_Reg[31] ),
    .ADR1(DLX_IDinst_jtarget[22]),
    .ADR2(DLX_IDinst_EPC[25]),
    .ADR3(DLX_IDinst_jtarget[21]),
    .O(\N163622/FROM )
  );
  defparam \DLX_IDinst__n0146<25>36 .INIT = 16'hA0EC;
  X_LUT4 \DLX_IDinst__n0146<25>36  (
    .ADR0(\DLX_IDinst_regA_eff[25] ),
    .ADR1(DLX_IDinst_N107105),
    .ADR2(N134590),
    .ADR3(N163622),
    .O(\N163622/GROM )
  );
  X_BUF \N163622/XUSED  (
    .I(\N163622/FROM ),
    .O(N163622)
  );
  X_BUF \N163622/YUSED  (
    .I(\N163622/GROM ),
    .O(CHOICE2798)
  );
  defparam \DLX_IDinst__n0146<17>36_SW0 .INIT = 16'hDD3F;
  X_LUT4 \DLX_IDinst__n0146<17>36_SW0  (
    .ADR0(\DLX_IDinst_Cause_Reg[31] ),
    .ADR1(DLX_IDinst_jtarget[22]),
    .ADR2(DLX_IDinst_EPC[17]),
    .ADR3(DLX_IDinst_jtarget[21]),
    .O(\N163588/FROM )
  );
  defparam \DLX_IDinst__n0146<17>36 .INIT = 16'h88F8;
  X_LUT4 \DLX_IDinst__n0146<17>36  (
    .ADR0(\DLX_IDinst_regA_eff[17] ),
    .ADR1(N134590),
    .ADR2(DLX_IDinst_N107105),
    .ADR3(N163588),
    .O(\N163588/GROM )
  );
  X_BUF \N163588/XUSED  (
    .I(\N163588/FROM ),
    .O(N163588)
  );
  X_BUF \N163588/YUSED  (
    .I(\N163588/GROM ),
    .O(CHOICE2678)
  );
  defparam \DLX_IDinst__n0145<0>40 .INIT = 16'hA800;
  X_LUT4 \DLX_IDinst__n0145<0>40  (
    .ADR0(DLX_IDinst_N107223),
    .ADR1(N135079),
    .ADR2(CHOICE2911),
    .ADR3(CHOICE2918),
    .O(\DLX_IDinst_counter<0>/FROM )
  );
  defparam \DLX_IDinst__n0145<0>52 .INIT = 16'hFF0C;
  X_LUT4 \DLX_IDinst__n0145<0>52  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst__n0387),
    .ADR2(DLX_IDinst_counter[0]),
    .ADR3(CHOICE2919),
    .O(N144314)
  );
  X_BUF \DLX_IDinst_counter<0>/XUSED  (
    .I(\DLX_IDinst_counter<0>/FROM ),
    .O(CHOICE2919)
  );
  defparam \DLX_EXinst__n0007<23>131_SW0 .INIT = 16'hFFFA;
  X_LUT4 \DLX_EXinst__n0007<23>131_SW0  (
    .ADR0(CHOICE3995),
    .ADR1(VCC),
    .ADR2(CHOICE4019),
    .ADR3(CHOICE4010),
    .O(\N163456/FROM )
  );
  defparam \DLX_EXinst__n0007<23>131 .INIT = 16'h0F08;
  X_LUT4 \DLX_EXinst__n0007<23>131  (
    .ADR0(DLX_EXinst_N76318),
    .ADR1(CHOICE4005),
    .ADR2(DLX_EXinst__n0036),
    .ADR3(N163456),
    .O(\N163456/GROM )
  );
  X_BUF \N163456/XUSED  (
    .I(\N163456/FROM ),
    .O(N163456)
  );
  X_BUF \N163456/YUSED  (
    .I(\N163456/GROM ),
    .O(CHOICE4023)
  );
  defparam \DLX_EXinst__n0007<15>220_SW0 .INIT = 16'hBBBA;
  X_LUT4 \DLX_EXinst__n0007<15>220_SW0  (
    .ADR0(CHOICE4312),
    .ADR1(\DLX_IDinst_Imm[4] ),
    .ADR2(CHOICE4301),
    .ADR3(CHOICE4302),
    .O(\N163477/FROM )
  );
  defparam \DLX_EXinst__n0007<15>220 .INIT = 16'hFFEA;
  X_LUT4 \DLX_EXinst__n0007<15>220  (
    .ADR0(CHOICE4308),
    .ADR1(CHOICE4294),
    .ADR2(\DLX_IDinst_Imm[15] ),
    .ADR3(N163477),
    .O(\N163477/GROM )
  );
  X_BUF \N163477/XUSED  (
    .I(\N163477/FROM ),
    .O(N163477)
  );
  X_BUF \N163477/YUSED  (
    .I(\N163477/GROM ),
    .O(CHOICE4314)
  );
  defparam \DLX_IDinst__n0146<26>36_SW0 .INIT = 16'hAF77;
  X_LUT4 \DLX_IDinst__n0146<26>36_SW0  (
    .ADR0(DLX_IDinst_jtarget[21]),
    .ADR1(\DLX_IDinst_Cause_Reg[31] ),
    .ADR2(DLX_IDinst_EPC[26]),
    .ADR3(DLX_IDinst_jtarget[22]),
    .O(\N163465/FROM )
  );
  defparam \DLX_IDinst__n0146<26>36 .INIT = 16'hA0EC;
  X_LUT4 \DLX_IDinst__n0146<26>36  (
    .ADR0(N134590),
    .ADR1(DLX_IDinst_N107105),
    .ADR2(\DLX_IDinst_regA_eff[26] ),
    .ADR3(N163465),
    .O(\N163465/GROM )
  );
  X_BUF \N163465/XUSED  (
    .I(\N163465/FROM ),
    .O(N163465)
  );
  X_BUF \N163465/YUSED  (
    .I(\N163465/GROM ),
    .O(CHOICE2813)
  );
  defparam \DLX_IDinst__n0146<18>36_SW0 .INIT = 16'h9DBF;
  X_LUT4 \DLX_IDinst__n0146<18>36_SW0  (
    .ADR0(DLX_IDinst_jtarget[21]),
    .ADR1(DLX_IDinst_jtarget[22]),
    .ADR2(DLX_IDinst_EPC[18]),
    .ADR3(\DLX_IDinst_Cause_Reg[31] ),
    .O(\N163452/FROM )
  );
  defparam \DLX_IDinst__n0146<18>36 .INIT = 16'hA0EC;
  X_LUT4 \DLX_IDinst__n0146<18>36  (
    .ADR0(\DLX_IDinst_regA_eff[18] ),
    .ADR1(DLX_IDinst_N107105),
    .ADR2(N134590),
    .ADR3(N163452),
    .O(\N163452/GROM )
  );
  X_BUF \N163452/XUSED  (
    .I(\N163452/FROM ),
    .O(N163452)
  );
  X_BUF \N163452/YUSED  (
    .I(\N163452/GROM ),
    .O(CHOICE2708)
  );
  defparam \DLX_EXinst_Mshift__n0022_Sh<24>_SW0 .INIT = 16'hD8D8;
  X_LUT4 \DLX_EXinst_Mshift__n0022_Sh<24>_SW0  (
    .ADR0(DLX_IDinst_Imm_1_1),
    .ADR1(DLX_IDinst_reg_out_A[27]),
    .ADR2(DLX_IDinst_reg_out_A[25]),
    .ADR3(VCC),
    .O(\N131077/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0022_Sh<24> .INIT = 16'hFA0A;
  X_LUT4 \DLX_EXinst_Mshift__n0022_Sh<24>  (
    .ADR0(DLX_EXinst_N73897),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_Imm_0_1),
    .ADR3(N131077),
    .O(\N131077/GROM )
  );
  X_BUF \N131077/XUSED  (
    .I(\N131077/FROM ),
    .O(N131077)
  );
  X_BUF \N131077/YUSED  (
    .I(\N131077/GROM ),
    .O(\DLX_EXinst_Mshift__n0022_Sh[24] )
  );
  defparam \DLX_IDinst__n0146<10>36_SW0 .INIT = 16'hD3DF;
  X_LUT4 \DLX_IDinst__n0146<10>36_SW0  (
    .ADR0(DLX_IDinst_EPC[10]),
    .ADR1(DLX_IDinst_jtarget[21]),
    .ADR2(DLX_IDinst_jtarget[22]),
    .ADR3(\DLX_IDinst_Cause_Reg[10] ),
    .O(\DLX_IDinst_Cause_Reg<10>/FROM )
  );
  defparam \DLX_IDinst__n0146<10>36 .INIT = 16'hA0EC;
  X_LUT4 \DLX_IDinst__n0146<10>36  (
    .ADR0(N134590),
    .ADR1(DLX_IDinst_N107105),
    .ADR2(\DLX_IDinst_regA_eff[10] ),
    .ADR3(N163578),
    .O(\DLX_IDinst_Cause_Reg<10>/GROM )
  );
  X_BUF \DLX_IDinst_Cause_Reg<10>/XUSED  (
    .I(\DLX_IDinst_Cause_Reg<10>/FROM ),
    .O(N163578)
  );
  X_BUF \DLX_IDinst_Cause_Reg<10>/YUSED  (
    .I(\DLX_IDinst_Cause_Reg<10>/GROM ),
    .O(CHOICE2573)
  );
  defparam \DLX_IDinst__n0146<11>36_SW0 .INIT = 16'h9DBF;
  X_LUT4 \DLX_IDinst__n0146<11>36_SW0  (
    .ADR0(DLX_IDinst_jtarget[22]),
    .ADR1(DLX_IDinst_jtarget[21]),
    .ADR2(\DLX_IDinst_Cause_Reg[11] ),
    .ADR3(DLX_IDinst_EPC[11]),
    .O(\DLX_IDinst_Cause_Reg<11>/FROM )
  );
  defparam \DLX_IDinst__n0146<11>36 .INIT = 16'h88F8;
  X_LUT4 \DLX_IDinst__n0146<11>36  (
    .ADR0(N134590),
    .ADR1(\DLX_IDinst_regA_eff[11] ),
    .ADR2(DLX_IDinst_N107105),
    .ADR3(N163234),
    .O(\DLX_IDinst_Cause_Reg<11>/GROM )
  );
  X_BUF \DLX_IDinst_Cause_Reg<11>/XUSED  (
    .I(\DLX_IDinst_Cause_Reg<11>/FROM ),
    .O(N163234)
  );
  X_BUF \DLX_IDinst_Cause_Reg<11>/YUSED  (
    .I(\DLX_IDinst_Cause_Reg<11>/GROM ),
    .O(CHOICE2588)
  );
  defparam \DLX_IDinst__n0146<12>36_SW0 .INIT = 16'hCF77;
  X_LUT4 \DLX_IDinst__n0146<12>36_SW0  (
    .ADR0(DLX_IDinst_EPC[12]),
    .ADR1(DLX_IDinst_jtarget[22]),
    .ADR2(\DLX_IDinst_Cause_Reg[12] ),
    .ADR3(DLX_IDinst_jtarget[21]),
    .O(\DLX_IDinst_Cause_Reg<12>/FROM )
  );
  defparam \DLX_IDinst__n0146<12>36 .INIT = 16'hA0EC;
  X_LUT4 \DLX_IDinst__n0146<12>36  (
    .ADR0(N134590),
    .ADR1(DLX_IDinst_N107105),
    .ADR2(\DLX_IDinst_regA_eff[12] ),
    .ADR3(N163361),
    .O(\DLX_IDinst_Cause_Reg<12>/GROM )
  );
  X_BUF \DLX_IDinst_Cause_Reg<12>/XUSED  (
    .I(\DLX_IDinst_Cause_Reg<12>/FROM ),
    .O(N163361)
  );
  X_BUF \DLX_IDinst_Cause_Reg<12>/YUSED  (
    .I(\DLX_IDinst_Cause_Reg<12>/GROM ),
    .O(CHOICE2603)
  );
  defparam \DLX_IDinst__n0146<13>36_SW0 .INIT = 16'hD3DF;
  X_LUT4 \DLX_IDinst__n0146<13>36_SW0  (
    .ADR0(DLX_IDinst_EPC[13]),
    .ADR1(DLX_IDinst_jtarget[21]),
    .ADR2(DLX_IDinst_jtarget[22]),
    .ADR3(\DLX_IDinst_Cause_Reg[13] ),
    .O(\DLX_IDinst_Cause_Reg<13>/FROM )
  );
  defparam \DLX_IDinst__n0146<13>36 .INIT = 16'hC0EA;
  X_LUT4 \DLX_IDinst__n0146<13>36  (
    .ADR0(DLX_IDinst_N107105),
    .ADR1(\DLX_IDinst_regA_eff[13] ),
    .ADR2(N134590),
    .ADR3(N163566),
    .O(\DLX_IDinst_Cause_Reg<13>/GROM )
  );
  X_BUF \DLX_IDinst_Cause_Reg<13>/XUSED  (
    .I(\DLX_IDinst_Cause_Reg<13>/FROM ),
    .O(N163566)
  );
  X_BUF \DLX_IDinst_Cause_Reg<13>/YUSED  (
    .I(\DLX_IDinst_Cause_Reg<13>/GROM ),
    .O(CHOICE2618)
  );
  defparam \DLX_IDinst__n0146<14>36_SW0 .INIT = 16'hB5BF;
  X_LUT4 \DLX_IDinst__n0146<14>36_SW0  (
    .ADR0(DLX_IDinst_jtarget[22]),
    .ADR1(\DLX_IDinst_Cause_Reg[14] ),
    .ADR2(DLX_IDinst_jtarget[21]),
    .ADR3(DLX_IDinst_EPC[14]),
    .O(\DLX_IDinst_Cause_Reg<14>/FROM )
  );
  defparam \DLX_IDinst__n0146<14>36 .INIT = 16'hC0EA;
  X_LUT4 \DLX_IDinst__n0146<14>36  (
    .ADR0(DLX_IDinst_N107105),
    .ADR1(N134590),
    .ADR2(\DLX_IDinst_regA_eff[14] ),
    .ADR3(N163382),
    .O(\DLX_IDinst_Cause_Reg<14>/GROM )
  );
  X_BUF \DLX_IDinst_Cause_Reg<14>/XUSED  (
    .I(\DLX_IDinst_Cause_Reg<14>/FROM ),
    .O(N163382)
  );
  X_BUF \DLX_IDinst_Cause_Reg<14>/YUSED  (
    .I(\DLX_IDinst_Cause_Reg<14>/GROM ),
    .O(CHOICE2633)
  );
  defparam \DLX_IDinst__n0146<15>36_SW0 .INIT = 16'h9BDF;
  X_LUT4 \DLX_IDinst__n0146<15>36_SW0  (
    .ADR0(DLX_IDinst_jtarget[22]),
    .ADR1(DLX_IDinst_jtarget[21]),
    .ADR2(DLX_IDinst_EPC[15]),
    .ADR3(\DLX_IDinst_Cause_Reg[15] ),
    .O(\DLX_IDinst_Cause_Reg<15>/FROM )
  );
  defparam \DLX_IDinst__n0146<15>36 .INIT = 16'h88F8;
  X_LUT4 \DLX_IDinst__n0146<15>36  (
    .ADR0(N134590),
    .ADR1(\DLX_IDinst_regA_eff[15] ),
    .ADR2(DLX_IDinst_N107105),
    .ADR3(N163329),
    .O(\DLX_IDinst_Cause_Reg<15>/GROM )
  );
  X_BUF \DLX_IDinst_Cause_Reg<15>/XUSED  (
    .I(\DLX_IDinst_Cause_Reg<15>/FROM ),
    .O(N163329)
  );
  X_BUF \DLX_IDinst_Cause_Reg<15>/YUSED  (
    .I(\DLX_IDinst_Cause_Reg<15>/GROM ),
    .O(CHOICE2648)
  );
  defparam \DLX_IDinst__n0146<27>36_SW0 .INIT = 16'hC7F7;
  X_LUT4 \DLX_IDinst__n0146<27>36_SW0  (
    .ADR0(\DLX_IDinst_Cause_Reg[31] ),
    .ADR1(DLX_IDinst_jtarget[21]),
    .ADR2(DLX_IDinst_jtarget[22]),
    .ADR3(DLX_IDinst_EPC[27]),
    .O(\DLX_IDinst_Cause_Reg<31>/FROM )
  );
  defparam \DLX_IDinst__n0146<27>36 .INIT = 16'hA0EC;
  X_LUT4 \DLX_IDinst__n0146<27>36  (
    .ADR0(N134590),
    .ADR1(DLX_IDinst_N107105),
    .ADR2(\DLX_IDinst_regA_eff[27] ),
    .ADR3(N163254),
    .O(\DLX_IDinst_Cause_Reg<31>/GROM )
  );
  X_BUF \DLX_IDinst_Cause_Reg<31>/XUSED  (
    .I(\DLX_IDinst_Cause_Reg<31>/FROM ),
    .O(N163254)
  );
  X_BUF \DLX_IDinst_Cause_Reg<31>/YUSED  (
    .I(\DLX_IDinst_Cause_Reg<31>/GROM ),
    .O(CHOICE2828)
  );
  defparam \DLX_EXinst_Mshift__n0019_Sh<23> .INIT = 16'hCCAA;
  X_LUT4 \DLX_EXinst_Mshift__n0019_Sh<23>  (
    .ADR0(DLX_EXinst_N73068),
    .ADR1(N130927),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[0]),
    .O(\DLX_EXinst_Mshift__n0019_Sh<23>/FROM )
  );
  defparam DLX_EXinst_Ker731011.INIT = 16'h4F40;
  X_LUT4 DLX_EXinst_Ker731011 (
    .ADR0(DLX_EXinst_N73239),
    .ADR1(DLX_IDinst_reg_out_A[31]),
    .ADR2(DLX_IDinst_reg_out_B[3]),
    .ADR3(\DLX_EXinst_Mshift__n0019_Sh[23] ),
    .O(\DLX_EXinst_Mshift__n0019_Sh<23>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0019_Sh<23>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0019_Sh<23>/FROM ),
    .O(\DLX_EXinst_Mshift__n0019_Sh[23] )
  );
  X_BUF \DLX_EXinst_Mshift__n0019_Sh<23>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0019_Sh<23>/GROM ),
    .O(DLX_EXinst_N73103)
  );
  defparam \vga_top_vga1_helpcounter_Madd__n0000_Mxor_Result<1>_Result1 .INIT = 16'h33CC;
  X_LUT4 \vga_top_vga1_helpcounter_Madd__n0000_Mxor_Result<1>_Result1  (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_helpcounter[1]),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_helpcounter[0]),
    .O(vga_top_vga1_helpcounter__n0000[1])
  );
  X_INV \vga_top_vga1_helpcounter<0>/BXMUX  (
    .I(vga_top_vga1_helpcounter[0]),
    .O(\vga_top_vga1_helpcounter<0>/BXMUXNOT )
  );
  defparam \DLX_IDinst__n0146<19>36_SW0 .INIT = 16'hDD3F;
  X_LUT4 \DLX_IDinst__n0146<19>36_SW0  (
    .ADR0(\DLX_IDinst_Cause_Reg[31] ),
    .ADR1(DLX_IDinst_jtarget[22]),
    .ADR2(DLX_IDinst_EPC[19]),
    .ADR3(DLX_IDinst_jtarget[21]),
    .O(\N163737/FROM )
  );
  defparam \DLX_IDinst__n0146<19>36 .INIT = 16'h88F8;
  X_LUT4 \DLX_IDinst__n0146<19>36  (
    .ADR0(N134590),
    .ADR1(\DLX_IDinst_regA_eff[19] ),
    .ADR2(DLX_IDinst_N107105),
    .ADR3(N163737),
    .O(\N163737/GROM )
  );
  X_BUF \N163737/XUSED  (
    .I(\N163737/FROM ),
    .O(N163737)
  );
  X_BUF \N163737/YUSED  (
    .I(\N163737/GROM ),
    .O(CHOICE2693)
  );
  defparam \DLX_EXinst__n0007<31>261_SW0 .INIT = 16'hFEFC;
  X_LUT4 \DLX_EXinst__n0007<31>261_SW0  (
    .ADR0(CHOICE5779),
    .ADR1(CHOICE5807),
    .ADR2(N164729),
    .ADR3(DLX_IDinst_reg_out_A[31]),
    .O(\N163550/FROM )
  );
  defparam \DLX_EXinst__n0007<31>261 .INIT = 16'hCCC8;
  X_LUT4 \DLX_EXinst__n0007<31>261  (
    .ADR0(CHOICE5764),
    .ADR1(DLX_EXinst__n0036),
    .ADR2(CHOICE5771),
    .ADR3(N163550),
    .O(\N163550/GROM )
  );
  X_BUF \N163550/XUSED  (
    .I(\N163550/FROM ),
    .O(N163550)
  );
  X_BUF \N163550/YUSED  (
    .I(\N163550/GROM ),
    .O(CHOICE5811)
  );
  defparam DLX_EXinst_Ker7437769_SW0.INIT = 16'hECEC;
  X_LUT4 DLX_EXinst_Ker7437769_SW0 (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(CHOICE3052),
    .ADR2(DLX_IDinst_reg_out_B_3_1),
    .ADR3(VCC),
    .O(\N163178/FROM )
  );
  defparam DLX_EXinst_Ker7437769.INIT = 16'h8F80;
  X_LUT4 DLX_EXinst_Ker7437769 (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(CHOICE3062),
    .ADR2(DLX_IDinst_reg_out_B[5]),
    .ADR3(N163178),
    .O(\N163178/GROM )
  );
  X_BUF \N163178/XUSED  (
    .I(\N163178/FROM ),
    .O(N163178)
  );
  X_BUF \N163178/YUSED  (
    .I(\N163178/GROM ),
    .O(CHOICE3065)
  );
  defparam \DLX_EXinst__n0007<1>98_SW0 .INIT = 16'hB800;
  X_LUT4 \DLX_EXinst__n0007<1>98_SW0  (
    .ADR0(N134488),
    .ADR1(\DLX_IDinst_Imm[2] ),
    .ADR2(CHOICE5702),
    .ADR3(DLX_EXinst_N76473),
    .O(\N163668/GROM )
  );
  X_BUF \N163668/YUSED  (
    .I(\N163668/GROM ),
    .O(N163668)
  );
  defparam DLX_IDinst_RegFile_19_27_1470.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_19_27_1470 (
    .I(DLX_IDinst_WB_data_eff[27]),
    .CE(DLX_IDinst__n0588),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_19_27)
  );
  defparam \DLX_IDinst__n0146<28>36_SW0 .INIT = 16'h9BDF;
  X_LUT4 \DLX_IDinst__n0146<28>36_SW0  (
    .ADR0(DLX_IDinst_jtarget[21]),
    .ADR1(DLX_IDinst_jtarget[22]),
    .ADR2(\DLX_IDinst_Cause_Reg[31] ),
    .ADR3(DLX_IDinst_EPC[28]),
    .O(\N163643/FROM )
  );
  defparam \DLX_IDinst__n0146<28>36 .INIT = 16'hA0EC;
  X_LUT4 \DLX_IDinst__n0146<28>36  (
    .ADR0(\DLX_IDinst_regA_eff[28] ),
    .ADR1(DLX_IDinst_N107105),
    .ADR2(N134590),
    .ADR3(N163643),
    .O(\N163643/GROM )
  );
  X_BUF \N163643/XUSED  (
    .I(\N163643/FROM ),
    .O(N163643)
  );
  X_BUF \N163643/YUSED  (
    .I(\N163643/GROM ),
    .O(CHOICE2843)
  );
  defparam DLX_EXinst_Ker730111.INIT = 16'hD8D8;
  X_LUT4 DLX_EXinst_Ker730111 (
    .ADR0(\DLX_IDinst_Imm[3] ),
    .ADR1(\DLX_EXinst_Mshift__n0020_Sh[29] ),
    .ADR2(\DLX_EXinst_Mshift__n0022_Sh[21] ),
    .ADR3(VCC),
    .O(\DLX_EXinst_N73013/FROM )
  );
  defparam \DLX_EXinst__n0007<31>382_SW0 .INIT = 16'hDDD8;
  X_LUT4 \DLX_EXinst__n0007<31>382_SW0  (
    .ADR0(\DLX_IDinst_Imm[3] ),
    .ADR1(\DLX_EXinst_Mshift__n0021_Sh[23] ),
    .ADR2(CHOICE5829),
    .ADR3(CHOICE5824),
    .O(\DLX_EXinst_N73013/GROM )
  );
  X_BUF \DLX_EXinst_N73013/XUSED  (
    .I(\DLX_EXinst_N73013/FROM ),
    .O(DLX_EXinst_N73013)
  );
  X_BUF \DLX_EXinst_N73013/YUSED  (
    .I(\DLX_EXinst_N73013/GROM ),
    .O(N163186)
  );
  defparam DLX_EXinst_Ker734221.INIT = 16'hAACC;
  X_LUT4 DLX_EXinst_Ker734221 (
    .ADR0(DLX_IDinst_reg_out_A[8]),
    .ADR1(DLX_IDinst_reg_out_A[6]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[1]),
    .O(\DLX_EXinst_N73424/FROM )
  );
  defparam DLX_EXinst_Ker7443415.INIT = 16'h00CA;
  X_LUT4 DLX_EXinst_Ker7443415 (
    .ADR0(DLX_IDinst_reg_out_A[4]),
    .ADR1(DLX_IDinst_reg_out_A[6]),
    .ADR2(DLX_IDinst_reg_out_B[1]),
    .ADR3(DLX_IDinst_reg_out_B[0]),
    .O(\DLX_EXinst_N73424/GROM )
  );
  X_BUF \DLX_EXinst_N73424/XUSED  (
    .I(\DLX_EXinst_N73424/FROM ),
    .O(DLX_EXinst_N73424)
  );
  X_BUF \DLX_EXinst_N73424/YUSED  (
    .I(\DLX_EXinst_N73424/GROM ),
    .O(CHOICE1749)
  );
  defparam DLX_EXinst_Ker7516254.INIT = 16'h30B8;
  X_LUT4 DLX_EXinst_Ker7516254 (
    .ADR0(\DLX_EXinst_Mshift__n0019_Sh[23] ),
    .ADR1(DLX_IDinst_reg_out_B_2_1),
    .ADR2(DLX_EXinst_N74976),
    .ADR3(DLX_IDinst_reg_out_B_3_1),
    .O(\CHOICE1907/FROM )
  );
  defparam DLX_EXinst_Ker7516264.INIT = 16'hD5C0;
  X_LUT4 DLX_EXinst_Ker7516264 (
    .ADR0(DLX_IDinst_reg_out_B[5]),
    .ADR1(DLX_IDinst_reg_out_A[31]),
    .ADR2(CHOICE1899),
    .ADR3(CHOICE1907),
    .O(\CHOICE1907/GROM )
  );
  X_BUF \CHOICE1907/XUSED  (
    .I(\CHOICE1907/FROM ),
    .O(CHOICE1907)
  );
  X_BUF \CHOICE1907/YUSED  (
    .I(\CHOICE1907/GROM ),
    .O(N138371)
  );
  defparam DLX_EXinst_Ker7514728.INIT = 16'h00B8;
  X_LUT4 DLX_EXinst_Ker7514728 (
    .ADR0(\DLX_EXinst_Mshift__n0020_Sh[29] ),
    .ADR1(DLX_IDinst_Imm_2_1),
    .ADR2(\DLX_EXinst_Mshift__n0020_Sh[25] ),
    .ADR3(\DLX_IDinst_Imm[5] ),
    .O(\CHOICE1921/FROM )
  );
  defparam DLX_EXinst_Ker7514764.INIT = 16'hCFCE;
  X_LUT4 DLX_EXinst_Ker7514764 (
    .ADR0(CHOICE1915),
    .ADR1(CHOICE1926),
    .ADR2(DLX_IDinst_Imm_3_1),
    .ADR3(CHOICE1921),
    .O(\CHOICE1921/GROM )
  );
  X_BUF \CHOICE1921/XUSED  (
    .I(\CHOICE1921/FROM ),
    .O(CHOICE1921)
  );
  X_BUF \CHOICE1921/YUSED  (
    .I(\CHOICE1921/GROM ),
    .O(N138481)
  );
  defparam DLX_EXinst_Ker7534054.INIT = 16'h50D8;
  X_LUT4 DLX_EXinst_Ker7534054 (
    .ADR0(DLX_IDinst_Imm_2_1),
    .ADR1(\DLX_EXinst_Mshift__n0022_Sh[23] ),
    .ADR2(DLX_EXinst_N75352),
    .ADR3(DLX_IDinst_Imm_3_1),
    .O(\CHOICE1963/FROM )
  );
  defparam DLX_EXinst_Ker7534064.INIT = 16'hB3A0;
  X_LUT4 DLX_EXinst_Ker7534064 (
    .ADR0(CHOICE1955),
    .ADR1(\DLX_IDinst_Imm[5] ),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(CHOICE1963),
    .O(\CHOICE1963/GROM )
  );
  X_BUF \CHOICE1963/XUSED  (
    .I(\CHOICE1963/FROM ),
    .O(CHOICE1963)
  );
  X_BUF \CHOICE1963/YUSED  (
    .I(\CHOICE1963/GROM ),
    .O(N138713)
  );
  defparam DLX_IDinst_Ker1085291.INIT = 16'h4000;
  X_LUT4 DLX_IDinst_Ker1085291 (
    .ADR0(DLX_MEMinst_reg_dst_out[2]),
    .ADR1(DLX_MEMinst_reg_write_MEM),
    .ADR2(DLX_MEMinst_reg_dst_out[0]),
    .ADR3(DLX_MEMinst_reg_dst_out[4]),
    .O(\DLX_MEMinst_reg_dst_out<0>/FROM )
  );
  defparam DLX_IDinst__n06041.INIT = 16'hC000;
  X_LUT4 DLX_IDinst__n06041 (
    .ADR0(VCC),
    .ADR1(DLX_MEMinst_reg_dst_out[1]),
    .ADR2(DLX_MEMinst_reg_dst_out[3]),
    .ADR3(DLX_IDinst_N108531),
    .O(\DLX_MEMinst_reg_dst_out<0>/GROM )
  );
  X_BUF \DLX_MEMinst_reg_dst_out<0>/XUSED  (
    .I(\DLX_MEMinst_reg_dst_out<0>/FROM ),
    .O(DLX_IDinst_N108531)
  );
  X_BUF \DLX_MEMinst_reg_dst_out<0>/YUSED  (
    .I(\DLX_MEMinst_reg_dst_out<0>/GROM ),
    .O(DLX_IDinst__n0604)
  );
  defparam DLX_IDinst_Ker1085221.INIT = 16'h8000;
  X_LUT4 DLX_IDinst_Ker1085221 (
    .ADR0(DLX_MEMinst_reg_write_MEM),
    .ADR1(DLX_MEMinst_reg_dst_out[4]),
    .ADR2(DLX_MEMinst_reg_dst_out[2]),
    .ADR3(DLX_MEMinst_reg_dst_out[0]),
    .O(\DLX_MEMinst_reg_dst_out<1>/FROM )
  );
  defparam DLX_IDinst__n06121.INIT = 16'h8800;
  X_LUT4 DLX_IDinst__n06121 (
    .ADR0(DLX_MEMinst_reg_dst_out[1]),
    .ADR1(DLX_MEMinst_reg_dst_out[3]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_N108524),
    .O(\DLX_MEMinst_reg_dst_out<1>/GROM )
  );
  X_BUF \DLX_MEMinst_reg_dst_out<1>/XUSED  (
    .I(\DLX_MEMinst_reg_dst_out<1>/FROM ),
    .O(DLX_IDinst_N108524)
  );
  X_BUF \DLX_MEMinst_reg_dst_out<1>/YUSED  (
    .I(\DLX_MEMinst_reg_dst_out<1>/GROM ),
    .O(DLX_IDinst__n0612)
  );
  defparam DLX_IDinst_Ker1085081.INIT = 16'h1000;
  X_LUT4 DLX_IDinst_Ker1085081 (
    .ADR0(DLX_MEMinst_reg_dst_out[2]),
    .ADR1(DLX_MEMinst_reg_dst_out[4]),
    .ADR2(DLX_MEMinst_reg_dst_out[0]),
    .ADR3(DLX_MEMinst_reg_write_MEM),
    .O(\DLX_MEMinst_reg_dst_out<2>/FROM )
  );
  defparam DLX_IDinst__n05721.INIT = 16'h8800;
  X_LUT4 DLX_IDinst__n05721 (
    .ADR0(DLX_MEMinst_reg_dst_out[1]),
    .ADR1(DLX_MEMinst_reg_dst_out[3]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_N108510),
    .O(\DLX_MEMinst_reg_dst_out<2>/GROM )
  );
  X_BUF \DLX_MEMinst_reg_dst_out<2>/XUSED  (
    .I(\DLX_MEMinst_reg_dst_out<2>/FROM ),
    .O(DLX_IDinst_N108510)
  );
  X_BUF \DLX_MEMinst_reg_dst_out<2>/YUSED  (
    .I(\DLX_MEMinst_reg_dst_out<2>/GROM ),
    .O(DLX_IDinst__n0572)
  );
  defparam DLX_EXinst_Ker7437256.INIT = 16'h0A0A;
  X_LUT4 DLX_EXinst_Ker7437256 (
    .ADR0(CHOICE3121),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[5]),
    .ADR3(VCC),
    .O(\CHOICE3122/FROM )
  );
  defparam DLX_EXinst_Ker74372135_SW0.INIT = 16'hCC80;
  X_LUT4 DLX_EXinst_Ker74372135_SW0 (
    .ADR0(CHOICE3113),
    .ADR1(N148609),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(CHOICE3122),
    .O(\CHOICE3122/GROM )
  );
  X_BUF \CHOICE3122/XUSED  (
    .I(\CHOICE3122/FROM ),
    .O(CHOICE3122)
  );
  X_BUF \CHOICE3122/YUSED  (
    .I(\CHOICE3122/GROM ),
    .O(N163618)
  );
  defparam DLX_EXinst_Ker763861.INIT = 16'h5500;
  X_LUT4 DLX_EXinst_Ker763861 (
    .ADR0(DLX_IDinst_reg_out_B_3_1),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[31]),
    .O(\DLX_EXinst_N76388/FROM )
  );
  defparam DLX_EXinst_Ker7436713.INIT = 16'hA808;
  X_LUT4 DLX_EXinst_Ker7436713 (
    .ADR0(DLX_IDinst_reg_out_B[2]),
    .ADR1(\DLX_EXinst_Mshift__n0019_Sh[25] ),
    .ADR2(DLX_IDinst_reg_out_B[3]),
    .ADR3(DLX_IDinst_reg_out_A[31]),
    .O(\DLX_EXinst_N76388/GROM )
  );
  X_BUF \DLX_EXinst_N76388/XUSED  (
    .I(\DLX_EXinst_N76388/FROM ),
    .O(DLX_EXinst_N76388)
  );
  X_BUF \DLX_EXinst_N76388/YUSED  (
    .I(\DLX_EXinst_N76388/GROM ),
    .O(CHOICE3026)
  );
  defparam DLX_IDinst_Ker1085431.INIT = 16'h4000;
  X_LUT4 DLX_IDinst_Ker1085431 (
    .ADR0(DLX_MEMinst_reg_dst_out[0]),
    .ADR1(DLX_MEMinst_reg_dst_out[2]),
    .ADR2(DLX_MEMinst_reg_write_MEM),
    .ADR3(DLX_MEMinst_reg_dst_out[4]),
    .O(\DLX_MEMinst_reg_dst_out<3>/FROM )
  );
  defparam DLX_IDinst__n06101.INIT = 16'hA000;
  X_LUT4 DLX_IDinst__n06101 (
    .ADR0(DLX_MEMinst_reg_dst_out[1]),
    .ADR1(VCC),
    .ADR2(DLX_MEMinst_reg_dst_out[3]),
    .ADR3(DLX_IDinst_N108545),
    .O(\DLX_MEMinst_reg_dst_out<3>/GROM )
  );
  X_BUF \DLX_MEMinst_reg_dst_out<3>/XUSED  (
    .I(\DLX_MEMinst_reg_dst_out<3>/FROM ),
    .O(DLX_IDinst_N108545)
  );
  X_BUF \DLX_MEMinst_reg_dst_out<3>/YUSED  (
    .I(\DLX_MEMinst_reg_dst_out<3>/GROM ),
    .O(DLX_IDinst__n0610)
  );
  X_ZERO \DLX_MEMinst_reg_dst_out<4>/LOGIC_ZERO_1471  (
    .O(\DLX_MEMinst_reg_dst_out<4>/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mcompar__n0368_inst_cy_264 (
    .IA(\DLX_MEMinst_reg_dst_out<4>/LOGIC_ZERO ),
    .IB(\DLX_MEMinst_reg_dst_out<4>/CYINIT ),
    .SEL(DLX_IDinst_Mcompar__n0368_inst_lut4_42),
    .O(\DLX_MEMinst_reg_dst_out<4>/CYMUXF )
  );
  defparam DLX_IDinst_Mcompar__n0368_inst_lut4_421.INIT = 16'hB487;
  X_LUT4 DLX_IDinst_Mcompar__n0368_inst_lut4_421 (
    .ADR0(DLX_IFinst_IR_latched[20]),
    .ADR1(DLX_EXinst__n0144),
    .ADR2(DLX_MEMinst_reg_dst_out[4]),
    .ADR3(DLX_IDinst_current_IR[20]),
    .O(DLX_IDinst_Mcompar__n0368_inst_lut4_42)
  );
  X_BUF \DLX_MEMinst_reg_dst_out<4>/XBUSED  (
    .I(\DLX_MEMinst_reg_dst_out<4>/CYMUXF ),
    .O(DLX_IDinst__n0368)
  );
  X_BUF \DLX_MEMinst_reg_dst_out<4>/CYINIT_1472  (
    .I(DLX_IDinst_Mcompar__n0368_inst_cy_263),
    .O(\DLX_MEMinst_reg_dst_out<4>/CYINIT )
  );
  defparam DLX_EXinst_Ker7515756.INIT = 16'h2020;
  X_LUT4 DLX_EXinst_Ker7515756 (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(\DLX_IDinst_Imm[5] ),
    .ADR2(DLX_IDinst_Imm_3_1),
    .ADR3(VCC),
    .O(\CHOICE1870/FROM )
  );
  defparam DLX_EXinst_Ker7515760.INIT = 16'hFF54;
  X_LUT4 DLX_EXinst_Ker7515760 (
    .ADR0(DLX_IDinst_Imm_3_1),
    .ADR1(CHOICE1859),
    .ADR2(CHOICE1865),
    .ADR3(CHOICE1870),
    .O(\CHOICE1870/GROM )
  );
  X_BUF \CHOICE1870/XUSED  (
    .I(\CHOICE1870/FROM ),
    .O(CHOICE1870)
  );
  X_BUF \CHOICE1870/YUSED  (
    .I(\CHOICE1870/GROM ),
    .O(N138143)
  );
  defparam DLX_EXinst_Ker7551832.INIT = 16'h0004;
  X_LUT4 DLX_EXinst_Ker7551832 (
    .ADR0(DLX_IDinst_reg_out_B[5]),
    .ADR1(\DLX_EXinst_Mshift__n0019_Sh[30] ),
    .ADR2(DLX_IDinst_reg_out_B_2_1),
    .ADR3(DLX_IDinst_reg_out_B_3_1),
    .O(\CHOICE2053/FROM )
  );
  defparam DLX_EXinst_Ker7551320.INIT = 16'h0008;
  X_LUT4 DLX_EXinst_Ker7551320 (
    .ADR0(DLX_IDinst_reg_out_B[5]),
    .ADR1(\DLX_EXinst_Mshift__n0019_Sh[61] ),
    .ADR2(DLX_IDinst_reg_out_B_2_1),
    .ADR3(DLX_IDinst_reg_out_B_3_1),
    .O(\CHOICE2053/GROM )
  );
  X_BUF \CHOICE2053/XUSED  (
    .I(\CHOICE2053/FROM ),
    .O(CHOICE2053)
  );
  X_BUF \CHOICE2053/YUSED  (
    .I(\CHOICE2053/GROM ),
    .O(CHOICE2035)
  );
  defparam DLX_IDinst_RegFile_19_19_1473.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_19_19_1473 (
    .I(DLX_IDinst_WB_data_eff[19]),
    .CE(DLX_IDinst__n0588),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_19_19)
  );
  defparam \DLX_EXinst__n0007<16>128_SW0 .INIT = 16'hA088;
  X_LUT4 \DLX_EXinst__n0007<16>128_SW0  (
    .ADR0(DLX_EXinst_N76457),
    .ADR1(DLX_EXinst_N74721),
    .ADR2(DLX_EXinst_N72809),
    .ADR3(DLX_IDinst_reg_out_B[2]),
    .O(\N164172/FROM )
  );
  defparam \DLX_EXinst__n0007<16>128 .INIT = 16'hFFF8;
  X_LUT4 \DLX_EXinst__n0007<16>128  (
    .ADR0(N134884),
    .ADR1(DLX_EXinst_ALU_result[16]),
    .ADR2(CHOICE4589),
    .ADR3(N164172),
    .O(\N164172/GROM )
  );
  X_BUF \N164172/XUSED  (
    .I(\N164172/FROM ),
    .O(N164172)
  );
  X_BUF \N164172/YUSED  (
    .I(\N164172/GROM ),
    .O(CHOICE4591)
  );
  defparam DLX_EXinst_Ker7550847.INIT = 16'h0008;
  X_LUT4 DLX_EXinst_Ker7550847 (
    .ADR0(DLX_EXinst_N76421),
    .ADR1(\DLX_EXinst_Mshift__n0019_Sh[28] ),
    .ADR2(DLX_IDinst_reg_out_B_2_1),
    .ADR3(DLX_IDinst_reg_out_B_3_1),
    .O(\CHOICE1280/FROM )
  );
  defparam DLX_EXinst_Ker7437750.INIT = 16'h01FF;
  X_LUT4 DLX_EXinst_Ker7437750 (
    .ADR0(DLX_IDinst_reg_out_B_2_1),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(DLX_IDinst_reg_out_B[0]),
    .ADR3(DLX_IDinst_reg_out_B_3_1),
    .O(\CHOICE1280/GROM )
  );
  X_BUF \CHOICE1280/XUSED  (
    .I(\CHOICE1280/FROM ),
    .O(CHOICE1280)
  );
  X_BUF \CHOICE1280/YUSED  (
    .I(\CHOICE1280/GROM ),
    .O(CHOICE3062)
  );
  defparam DLX_IDinst_RegFile_27_27_1474.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_27_27_1474 (
    .I(DLX_IDinst_WB_data_eff[27]),
    .CE(DLX_IDinst__n0604),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_27_27)
  );
  defparam DLX_EXinst_Ker7551350.INIT = 16'hFFE0;
  X_LUT4 DLX_EXinst_Ker7551350 (
    .ADR0(CHOICE2032),
    .ADR1(CHOICE2035),
    .ADR2(N148609),
    .ADR3(CHOICE2040),
    .O(\N139189/FROM )
  );
  defparam \DLX_EXinst__n0007<29>273 .INIT = 16'hEFEE;
  X_LUT4 \DLX_EXinst__n0007<29>273  (
    .ADR0(CHOICE4812),
    .ADR1(CHOICE4834),
    .ADR2(DLX_IDinst_reg_out_B[4]),
    .ADR3(N139189),
    .O(\N139189/GROM )
  );
  X_BUF \N139189/XUSED  (
    .I(\N139189/FROM ),
    .O(N139189)
  );
  X_BUF \N139189/YUSED  (
    .I(\N139189/GROM ),
    .O(CHOICE4835)
  );
  defparam DLX_EXinst_Ker7621835.INIT = 16'h000E;
  X_LUT4 DLX_EXinst_Ker7621835 (
    .ADR0(CHOICE1669),
    .ADR1(CHOICE1670),
    .ADR2(DLX_IDinst_IR_opcode_field[4]),
    .ADR3(DLX_EXinst__n0036),
    .O(\N136960/FROM )
  );
  defparam \DLX_EXinst__n0013<16>1 .INIT = 16'hECA0;
  X_LUT4 \DLX_EXinst__n0013<16>1  (
    .ADR0(DLX_IDinst_reg_out_B[16]),
    .ADR1(\DLX_IDinst_Imm[31] ),
    .ADR2(DLX_EXinst__n0036),
    .ADR3(N136960),
    .O(\N136960/GROM )
  );
  X_BUF \N136960/XUSED  (
    .I(\N136960/FROM ),
    .O(N136960)
  );
  X_BUF \N136960/YUSED  (
    .I(\N136960/GROM ),
    .O(DLX_EXinst__n0013[16])
  );
  defparam DLX_EXinst_Ker7465298.INIT = 16'h4E44;
  X_LUT4 DLX_EXinst_Ker7465298 (
    .ADR0(DLX_IDinst_Imm_2_1),
    .ADR1(DLX_EXinst_N73163),
    .ADR2(DLX_IDinst_Imm_3_1),
    .ADR3(\DLX_EXinst_Mshift__n0020_Sh[26] ),
    .O(\CHOICE2945/FROM )
  );
  defparam DLX_EXinst_Ker7465213.INIT = 16'h88A0;
  X_LUT4 DLX_EXinst_Ker7465213 (
    .ADR0(DLX_IDinst_Imm_2_1),
    .ADR1(DLX_IDinst_reg_out_A[31]),
    .ADR2(\DLX_EXinst_Mshift__n0020_Sh[26] ),
    .ADR3(DLX_IDinst_Imm_3_1),
    .O(\CHOICE2945/GROM )
  );
  X_BUF \CHOICE2945/XUSED  (
    .I(\CHOICE2945/FROM ),
    .O(CHOICE2945)
  );
  X_BUF \CHOICE2945/YUSED  (
    .I(\CHOICE2945/GROM ),
    .O(CHOICE2926)
  );
  defparam \DLX_EXinst__n0008<26>1 .INIT = 16'h8888;
  X_LUT4 \DLX_EXinst__n0008<26>1  (
    .ADR0(DLX_EXinst_N72746),
    .ADR1(DLX_IDinst_reg_out_B[26]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst__n0008[26])
  );
  defparam DLX_EXinst_Ker7618131.INIT = 16'h0001;
  X_LUT4 DLX_EXinst_Ker7618131 (
    .ADR0(DLX_IDinst_reg_out_B[28]),
    .ADR1(DLX_IDinst_reg_out_B[27]),
    .ADR2(DLX_IDinst_reg_out_B[26]),
    .ADR3(DLX_IDinst_reg_out_B[29]),
    .O(\DLX_EXinst_reg_out_B_EX<26>/GROM )
  );
  X_BUF \DLX_EXinst_reg_out_B_EX<26>/YUSED  (
    .I(\DLX_EXinst_reg_out_B_EX<26>/GROM ),
    .O(CHOICE3608)
  );
  defparam DLX_EXinst_Ker7618144.INIT = 16'h0001;
  X_LUT4 DLX_EXinst_Ker7618144 (
    .ADR0(DLX_IDinst_reg_out_B[23]),
    .ADR1(DLX_IDinst_reg_out_B[22]),
    .ADR2(DLX_IDinst_reg_out_B[24]),
    .ADR3(DLX_IDinst_reg_out_B[25]),
    .O(\CHOICE3615/FROM )
  );
  defparam DLX_EXinst_Ker7618145.INIT = 16'hF000;
  X_LUT4 DLX_EXinst_Ker7618145 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(CHOICE3608),
    .ADR3(CHOICE3615),
    .O(\CHOICE3615/GROM )
  );
  X_BUF \CHOICE3615/XUSED  (
    .I(\CHOICE3615/FROM ),
    .O(CHOICE3615)
  );
  X_BUF \CHOICE3615/YUSED  (
    .I(\CHOICE3615/GROM ),
    .O(CHOICE3616)
  );
  defparam DLX_EXinst_Ker7550849.INIT = 16'hFFC0;
  X_LUT4 DLX_EXinst_Ker7550849 (
    .ADR0(VCC),
    .ADR1(CHOICE1276),
    .ADR2(N148609),
    .ADR3(CHOICE1280),
    .O(\N134683/FROM )
  );
  defparam \DLX_EXinst__n0007<28>325 .INIT = 16'hFBFA;
  X_LUT4 \DLX_EXinst__n0007<28>325  (
    .ADR0(CHOICE4886),
    .ADR1(DLX_IDinst_reg_out_B[4]),
    .ADR2(CHOICE4911),
    .ADR3(N134683),
    .O(\N134683/GROM )
  );
  X_BUF \N134683/XUSED  (
    .I(\N134683/FROM ),
    .O(N134683)
  );
  X_BUF \N134683/YUSED  (
    .I(\N134683/GROM ),
    .O(CHOICE4912)
  );
  defparam \DLX_EXinst__n0008<18>1 .INIT = 16'h8888;
  X_LUT4 \DLX_EXinst__n0008<18>1  (
    .ADR0(DLX_EXinst_N72746),
    .ADR1(DLX_IDinst_reg_out_B[18]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst__n0008[18])
  );
  defparam DLX_EXinst_Ker7618183.INIT = 16'h0001;
  X_LUT4 DLX_EXinst_Ker7618183 (
    .ADR0(DLX_IDinst_reg_out_B[20]),
    .ADR1(DLX_IDinst_reg_out_B[19]),
    .ADR2(DLX_IDinst_reg_out_B[18]),
    .ADR3(DLX_IDinst_reg_out_B[21]),
    .O(\DLX_EXinst_reg_out_B_EX<18>/GROM )
  );
  X_BUF \DLX_EXinst_reg_out_B_EX<18>/YUSED  (
    .I(\DLX_EXinst_reg_out_B_EX<18>/GROM ),
    .O(CHOICE3624)
  );
  defparam DLX_EXinst_Ker7551866.INIT = 16'hFCEC;
  X_LUT4 DLX_EXinst_Ker7551866 (
    .ADR0(CHOICE2049),
    .ADR1(CHOICE2058),
    .ADR2(N148609),
    .ADR3(CHOICE2053),
    .O(\N139297/FROM )
  );
  defparam \DLX_EXinst__n0007<30>273 .INIT = 16'hFDFC;
  X_LUT4 \DLX_EXinst__n0007<30>273  (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(CHOICE4763),
    .ADR2(CHOICE4741),
    .ADR3(N139297),
    .O(\N139297/GROM )
  );
  X_BUF \N139297/XUSED  (
    .I(\N139297/FROM ),
    .O(N139297)
  );
  X_BUF \N139297/YUSED  (
    .I(\N139297/GROM ),
    .O(CHOICE4764)
  );
  defparam DLX_EXinst_Ker7465715.INIT = 16'h3202;
  X_LUT4 DLX_EXinst_Ker7465715 (
    .ADR0(\DLX_EXinst_Mshift__n0022_Sh[23] ),
    .ADR1(DLX_IDinst_Imm_3_1),
    .ADR2(DLX_IDinst_Imm_2_1),
    .ADR3(\DLX_EXinst_Mshift__n0020_Sh[27] ),
    .O(\CHOICE3081/FROM )
  );
  defparam DLX_EXinst_Ker7465769_SW0.INIT = 16'hFFA0;
  X_LUT4 DLX_EXinst_Ker7465769_SW0 (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_Imm_3_1),
    .ADR3(CHOICE3081),
    .O(\CHOICE3081/GROM )
  );
  X_BUF \CHOICE3081/XUSED  (
    .I(\CHOICE3081/FROM ),
    .O(CHOICE3081)
  );
  X_BUF \CHOICE3081/YUSED  (
    .I(\CHOICE3081/GROM ),
    .O(N163140)
  );
  defparam DLX_EXinst_Ker7465750.INIT = 16'h3337;
  X_LUT4 DLX_EXinst_Ker7465750 (
    .ADR0(DLX_IDinst_Imm_1_1),
    .ADR1(DLX_IDinst_Imm_3_1),
    .ADR2(\DLX_IDinst_Imm[0] ),
    .ADR3(DLX_IDinst_Imm_2_1),
    .O(\CHOICE3091/FROM )
  );
  defparam DLX_EXinst_Ker7465769.INIT = 16'hE444;
  X_LUT4 DLX_EXinst_Ker7465769 (
    .ADR0(\DLX_IDinst_Imm[5] ),
    .ADR1(N163140),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(CHOICE3091),
    .O(\CHOICE3091/GROM )
  );
  X_BUF \CHOICE3091/XUSED  (
    .I(\CHOICE3091/FROM ),
    .O(CHOICE3091)
  );
  X_BUF \CHOICE3091/YUSED  (
    .I(\CHOICE3091/GROM ),
    .O(CHOICE3094)
  );
  defparam DLX_EXinst_Ker7565247.INIT = 16'h1000;
  X_LUT4 DLX_EXinst_Ker7565247 (
    .ADR0(DLX_IDinst_Imm_3_1),
    .ADR1(DLX_IDinst_Imm_2_1),
    .ADR2(DLX_EXinst_N76441),
    .ADR3(\DLX_EXinst_Mshift__n0020_Sh[28] ),
    .O(\CHOICE1295/FROM )
  );
  defparam \DLX_EXinst__n0007<12>134 .INIT = 16'hCC80;
  X_LUT4 \DLX_EXinst__n0007<12>134  (
    .ADR0(CHOICE1291),
    .ADR1(\DLX_IDinst_Imm[4] ),
    .ADR2(N147520),
    .ADR3(CHOICE1295),
    .O(\CHOICE1295/GROM )
  );
  X_BUF \CHOICE1295/XUSED  (
    .I(\CHOICE1295/FROM ),
    .O(CHOICE1295)
  );
  X_BUF \CHOICE1295/YUSED  (
    .I(\CHOICE1295/GROM ),
    .O(CHOICE3795)
  );
  defparam DLX_EXinst_Ker7565720.INIT = 16'h0040;
  X_LUT4 DLX_EXinst_Ker7565720 (
    .ADR0(DLX_IDinst_Imm_3_1),
    .ADR1(\DLX_EXinst_Mshift__n0020_Sh[61] ),
    .ADR2(\DLX_IDinst_Imm[5] ),
    .ADR3(DLX_IDinst_Imm_2_1),
    .O(\CHOICE2020/FROM )
  );
  defparam DLX_EXinst_Ker7566232.INIT = 16'h0002;
  X_LUT4 DLX_EXinst_Ker7566232 (
    .ADR0(\DLX_EXinst_Mshift__n0020_Sh[30] ),
    .ADR1(DLX_IDinst_Imm_3_1),
    .ADR2(DLX_IDinst_Imm_2_1),
    .ADR3(\DLX_IDinst_Imm[5] ),
    .O(\CHOICE2020/GROM )
  );
  X_BUF \CHOICE2020/XUSED  (
    .I(\CHOICE2020/FROM ),
    .O(CHOICE2020)
  );
  X_BUF \CHOICE2020/YUSED  (
    .I(\CHOICE2020/GROM ),
    .O(CHOICE2071)
  );
  defparam DLX_EXinst_Ker735471.INIT = 16'hF5A0;
  X_LUT4 DLX_EXinst_Ker735471 (
    .ADR0(DLX_IDinst_Imm_1_1),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[8]),
    .ADR3(DLX_IDinst_reg_out_A[6]),
    .O(\DLX_EXinst_N73549/FROM )
  );
  defparam DLX_EXinst_Ker7566225.INIT = 16'h0A20;
  X_LUT4 DLX_EXinst_Ker7566225 (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(DLX_IDinst_Imm_1_1),
    .ADR2(\DLX_IDinst_Imm[5] ),
    .ADR3(DLX_EXinst_N72815),
    .O(\DLX_EXinst_N73549/GROM )
  );
  X_BUF \DLX_EXinst_N73549/XUSED  (
    .I(\DLX_EXinst_N73549/FROM ),
    .O(DLX_EXinst_N73549)
  );
  X_BUF \DLX_EXinst_N73549/YUSED  (
    .I(\DLX_EXinst_N73549/GROM ),
    .O(CHOICE2067)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5410.INIT = 16'h2000;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5410 (
    .ADR0(DLX_IDinst_jtarget[20]),
    .ADR1(DLX_IDinst_jtarget[19]),
    .ADR2(DLX_IDinst_jtarget[18]),
    .ADR3(DLX_IDinst_jtarget[17]),
    .O(\DLX_IDinst_Mmux__COND_4_inst_lut4_54/FROM )
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5010.INIT = 16'h2000;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5010 (
    .ADR0(DLX_IDinst_jtarget[19]),
    .ADR1(DLX_IDinst_jtarget[20]),
    .ADR2(DLX_IDinst_jtarget[17]),
    .ADR3(DLX_IDinst_jtarget[18]),
    .O(\DLX_IDinst_Mmux__COND_4_inst_lut4_54/GROM )
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_lut4_54/XUSED  (
    .I(\DLX_IDinst_Mmux__COND_4_inst_lut4_54/FROM ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_54)
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_lut4_54/YUSED  (
    .I(\DLX_IDinst_Mmux__COND_4_inst_lut4_54/GROM ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_50)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5310.INIT = 16'h0040;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5310 (
    .ADR0(DLX_IDinst_jtarget[19]),
    .ADR1(DLX_IDinst_jtarget[18]),
    .ADR2(DLX_IDinst_jtarget[20]),
    .ADR3(DLX_IDinst_jtarget[17]),
    .O(\DLX_IDinst_Mmux__COND_4_inst_lut4_53/FROM )
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4310.INIT = 16'h0001;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4310 (
    .ADR0(DLX_IDinst_jtarget[17]),
    .ADR1(DLX_IDinst_jtarget[19]),
    .ADR2(DLX_IDinst_jtarget[20]),
    .ADR3(DLX_IDinst_jtarget[18]),
    .O(\DLX_IDinst_Mmux__COND_4_inst_lut4_53/GROM )
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_lut4_53/XUSED  (
    .I(\DLX_IDinst_Mmux__COND_4_inst_lut4_53/FROM ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_53)
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_lut4_53/YUSED  (
    .I(\DLX_IDinst_Mmux__COND_4_inst_lut4_53/GROM ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_43)
  );
  defparam DLX_EXinst_Ker7565747.INIT = 16'h0400;
  X_LUT4 DLX_EXinst_Ker7565747 (
    .ADR0(DLX_IDinst_Imm_3_1),
    .ADR1(DLX_EXinst_N76441),
    .ADR2(DLX_IDinst_Imm_2_1),
    .ADR3(\DLX_EXinst_Mshift__n0022_Sh[29] ),
    .O(\CHOICE2025/FROM )
  );
  defparam DLX_EXinst_Ker7566263.INIT = 16'h0400;
  X_LUT4 DLX_EXinst_Ker7566263 (
    .ADR0(DLX_IDinst_Imm_3_1),
    .ADR1(DLX_EXinst_N76441),
    .ADR2(DLX_IDinst_Imm_2_1),
    .ADR3(\DLX_EXinst_Mshift__n0022_Sh[30] ),
    .O(\CHOICE2025/GROM )
  );
  X_BUF \CHOICE2025/XUSED  (
    .I(\CHOICE2025/FROM ),
    .O(CHOICE2025)
  );
  X_BUF \CHOICE2025/YUSED  (
    .I(\CHOICE2025/GROM ),
    .O(CHOICE2076)
  );
  defparam DLX_EXinst_Ker7566266.INIT = 16'hFFE0;
  X_LUT4 DLX_EXinst_Ker7566266 (
    .ADR0(CHOICE2071),
    .ADR1(CHOICE2067),
    .ADR2(N147520),
    .ADR3(CHOICE2076),
    .O(\N139405/FROM )
  );
  defparam \DLX_EXinst__n0007<30>116 .INIT = 16'hFDFC;
  X_LUT4 \DLX_EXinst__n0007<30>116  (
    .ADR0(\DLX_IDinst_Imm[4] ),
    .ADR1(CHOICE4730),
    .ADR2(CHOICE4708),
    .ADR3(N139405),
    .O(\N139405/GROM )
  );
  X_BUF \N139405/XUSED  (
    .I(\N139405/FROM ),
    .O(N139405)
  );
  X_BUF \N139405/YUSED  (
    .I(\N139405/GROM ),
    .O(CHOICE4731)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4910.INIT = 16'h0020;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4910 (
    .ADR0(DLX_IDinst_jtarget[19]),
    .ADR1(DLX_IDinst_jtarget[17]),
    .ADR2(DLX_IDinst_jtarget[18]),
    .ADR3(DLX_IDinst_jtarget[20]),
    .O(\DLX_IDinst_Mmux__COND_4_inst_lut4_49/FROM )
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5210.INIT = 16'h0400;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5210 (
    .ADR0(DLX_IDinst_jtarget[18]),
    .ADR1(DLX_IDinst_jtarget[17]),
    .ADR2(DLX_IDinst_jtarget[19]),
    .ADR3(DLX_IDinst_jtarget[20]),
    .O(\DLX_IDinst_Mmux__COND_4_inst_lut4_49/GROM )
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_lut4_49/XUSED  (
    .I(\DLX_IDinst_Mmux__COND_4_inst_lut4_49/FROM ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_49)
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_lut4_49/YUSED  (
    .I(\DLX_IDinst_Mmux__COND_4_inst_lut4_49/GROM ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_52)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4810.INIT = 16'h0020;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4810 (
    .ADR0(DLX_IDinst_jtarget[17]),
    .ADR1(DLX_IDinst_jtarget[18]),
    .ADR2(DLX_IDinst_jtarget[19]),
    .ADR3(DLX_IDinst_jtarget[20]),
    .O(\DLX_IDinst_Mmux__COND_4_inst_lut4_48/FROM )
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4410.INIT = 16'h0010;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4410 (
    .ADR0(DLX_IDinst_jtarget[20]),
    .ADR1(DLX_IDinst_jtarget[18]),
    .ADR2(DLX_IDinst_jtarget[17]),
    .ADR3(DLX_IDinst_jtarget[19]),
    .O(\DLX_IDinst_Mmux__COND_4_inst_lut4_48/GROM )
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_lut4_48/XUSED  (
    .I(\DLX_IDinst_Mmux__COND_4_inst_lut4_48/FROM ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_48)
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_lut4_48/YUSED  (
    .I(\DLX_IDinst_Mmux__COND_4_inst_lut4_48/GROM ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_44)
  );
  defparam DLX_EXinst_Ker730561.INIT = 16'hAAF0;
  X_LUT4 DLX_EXinst_Ker730561 (
    .ADR0(DLX_IDinst_reg_out_A[21]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[19]),
    .ADR3(DLX_IDinst_reg_out_B[1]),
    .O(\DLX_EXinst_N73058/FROM )
  );
  defparam DLX_EXinst_Ker7495411.INIT = 16'h20A0;
  X_LUT4 DLX_EXinst_Ker7495411 (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(DLX_IDinst_reg_out_B_2_1),
    .ADR2(DLX_IDinst_reg_out_B[5]),
    .ADR3(DLX_IDinst_reg_out_B[1]),
    .O(\DLX_EXinst_N73058/GROM )
  );
  X_BUF \DLX_EXinst_N73058/XUSED  (
    .I(\DLX_EXinst_N73058/FROM ),
    .O(DLX_EXinst_N73058)
  );
  X_BUF \DLX_EXinst_N73058/YUSED  (
    .I(\DLX_EXinst_N73058/GROM ),
    .O(CHOICE1877)
  );
  defparam \DLX_IDinst__n0146<29>36_SW0 .INIT = 16'hD3DF;
  X_LUT4 \DLX_IDinst__n0146<29>36_SW0  (
    .ADR0(\DLX_IDinst_Cause_Reg[31] ),
    .ADR1(DLX_IDinst_jtarget[22]),
    .ADR2(DLX_IDinst_jtarget[21]),
    .ADR3(DLX_IDinst_EPC[29]),
    .O(\N163506/FROM )
  );
  defparam \DLX_IDinst__n0146<29>36 .INIT = 16'hA0EC;
  X_LUT4 \DLX_IDinst__n0146<29>36  (
    .ADR0(N134590),
    .ADR1(DLX_IDinst_N107105),
    .ADR2(\DLX_IDinst_regA_eff[29] ),
    .ADR3(N163506),
    .O(\N163506/GROM )
  );
  X_BUF \N163506/XUSED  (
    .I(\N163506/FROM ),
    .O(N163506)
  );
  X_BUF \N163506/YUSED  (
    .I(\N163506/GROM ),
    .O(CHOICE2858)
  );
  defparam DLX_EXinst_Ker7565750.INIT = 16'hFFA8;
  X_LUT4 DLX_EXinst_Ker7565750 (
    .ADR0(N147520),
    .ADR1(CHOICE2020),
    .ADR2(CHOICE2017),
    .ADR3(CHOICE2025),
    .O(\N139100/FROM )
  );
  defparam \DLX_EXinst__n0007<29>116 .INIT = 16'hEFEE;
  X_LUT4 \DLX_EXinst__n0007<29>116  (
    .ADR0(CHOICE4801),
    .ADR1(CHOICE4779),
    .ADR2(\DLX_IDinst_Imm[4] ),
    .ADR3(N139100),
    .O(\N139100/GROM )
  );
  X_BUF \N139100/XUSED  (
    .I(\N139100/FROM ),
    .O(N139100)
  );
  X_BUF \N139100/YUSED  (
    .I(\N139100/GROM ),
    .O(CHOICE4802)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4710.INIT = 16'h0010;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4710 (
    .ADR0(DLX_IDinst_jtarget[18]),
    .ADR1(DLX_IDinst_jtarget[17]),
    .ADR2(DLX_IDinst_jtarget[19]),
    .ADR3(DLX_IDinst_jtarget[20]),
    .O(\DLX_IDinst_Mmux__COND_4_inst_lut4_47/FROM )
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4510.INIT = 16'h0004;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4510 (
    .ADR0(DLX_IDinst_jtarget[17]),
    .ADR1(DLX_IDinst_jtarget[18]),
    .ADR2(DLX_IDinst_jtarget[20]),
    .ADR3(DLX_IDinst_jtarget[19]),
    .O(\DLX_IDinst_Mmux__COND_4_inst_lut4_47/GROM )
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_lut4_47/XUSED  (
    .I(\DLX_IDinst_Mmux__COND_4_inst_lut4_47/FROM ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_47)
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_lut4_47/YUSED  (
    .I(\DLX_IDinst_Mmux__COND_4_inst_lut4_47/GROM ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_45)
  );
  defparam \DLX_IDinst__n0135<4> .INIT = 16'h00C8;
  X_LUT4 \DLX_IDinst__n0135<4>  (
    .ADR0(DLX_IDinst__n0453),
    .ADR1(DLX_IDinst_jtarget[20]),
    .ADR2(N127400),
    .ADR3(DLX_IDinst_N108456),
    .O(DLX_IDinst__n0135[4])
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4610.INIT = 16'h1000;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4610 (
    .ADR0(DLX_IDinst_jtarget[19]),
    .ADR1(DLX_IDinst_jtarget[20]),
    .ADR2(DLX_IDinst_jtarget[17]),
    .ADR3(DLX_IDinst_jtarget[18]),
    .O(\DLX_IDinst_rt_addr<4>/GROM )
  );
  X_BUF \DLX_IDinst_rt_addr<4>/YUSED  (
    .I(\DLX_IDinst_rt_addr<4>/GROM ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_46)
  );
  defparam DLX_EXinst_Ker7495456.INIT = 16'h0A00;
  X_LUT4 DLX_EXinst_Ker7495456 (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[5]),
    .ADR3(DLX_IDinst_reg_out_B_3_1),
    .O(\CHOICE1888/FROM )
  );
  defparam DLX_EXinst_Ker7495460.INIT = 16'hFF54;
  X_LUT4 DLX_EXinst_Ker7495460 (
    .ADR0(DLX_IDinst_reg_out_B_3_1),
    .ADR1(CHOICE1877),
    .ADR2(CHOICE1883),
    .ADR3(CHOICE1888),
    .O(\CHOICE1888/GROM )
  );
  X_BUF \CHOICE1888/XUSED  (
    .I(\CHOICE1888/FROM ),
    .O(CHOICE1888)
  );
  X_BUF \CHOICE1888/YUSED  (
    .I(\CHOICE1888/GROM ),
    .O(N138249)
  );
  defparam DLX_EXinst_Ker7495928.INIT = 16'h5404;
  X_LUT4 DLX_EXinst_Ker7495928 (
    .ADR0(DLX_IDinst_reg_out_B[5]),
    .ADR1(\DLX_EXinst_Mshift__n0019_Sh[25] ),
    .ADR2(DLX_IDinst_reg_out_B_2_1),
    .ADR3(\DLX_EXinst_Mshift__n0019_Sh[29] ),
    .O(\CHOICE1939/FROM )
  );
  defparam DLX_EXinst_Ker7495964.INIT = 16'hAFAE;
  X_LUT4 DLX_EXinst_Ker7495964 (
    .ADR0(CHOICE1944),
    .ADR1(CHOICE1933),
    .ADR2(DLX_IDinst_reg_out_B_3_1),
    .ADR3(CHOICE1939),
    .O(\CHOICE1939/GROM )
  );
  X_BUF \CHOICE1939/XUSED  (
    .I(\CHOICE1939/FROM ),
    .O(CHOICE1939)
  );
  X_BUF \CHOICE1939/YUSED  (
    .I(\CHOICE1939/GROM ),
    .O(N138591)
  );
  defparam \DLX_EXinst__n0007<31>567_SW0 .INIT = 16'hAAFE;
  X_LUT4 \DLX_EXinst__n0007<31>567_SW0  (
    .ADR0(CHOICE5864),
    .ADR1(CHOICE5841),
    .ADR2(CHOICE5838),
    .ADR3(N146478),
    .O(\DLX_EXinst_ALU_result<31>/FROM )
  );
  defparam \DLX_EXinst__n0007<31>567 .INIT = 16'h0F0E;
  X_LUT4 \DLX_EXinst__n0007<31>567  (
    .ADR0(CHOICE5846),
    .ADR1(CHOICE5850),
    .ADR2(DLX_EXinst__n0036),
    .ADR3(N163497),
    .O(CHOICE5867)
  );
  X_BUF \DLX_EXinst_ALU_result<31>/XUSED  (
    .I(\DLX_EXinst_ALU_result<31>/FROM ),
    .O(N163497)
  );
  defparam \DLX_EXinst__n0007<24>247_SW0 .INIT = 16'hFCCC;
  X_LUT4 \DLX_EXinst__n0007<24>247_SW0  (
    .ADR0(VCC),
    .ADR1(CHOICE5631),
    .ADR2(N148609),
    .ADR3(CHOICE5598),
    .O(\N163246/FROM )
  );
  defparam \DLX_EXinst__n0007<24>247 .INIT = 16'hCCC8;
  X_LUT4 \DLX_EXinst__n0007<24>247  (
    .ADR0(CHOICE5603),
    .ADR1(DLX_EXinst__n0036),
    .ADR2(CHOICE5585),
    .ADR3(N163246),
    .O(\N163246/GROM )
  );
  X_BUF \N163246/XUSED  (
    .I(\N163246/FROM ),
    .O(N163246)
  );
  X_BUF \N163246/YUSED  (
    .I(\N163246/GROM ),
    .O(CHOICE5634)
  );
  defparam DLX_IDinst_Ker108226127.INIT = 16'h0010;
  X_LUT4 DLX_IDinst_Ker108226127 (
    .ADR0(N163124),
    .ADR1(DLX_IDinst_Ker1084541_1),
    .ADR2(CHOICE3396),
    .ADR3(DLX_IDinst__n0098),
    .O(\N147200/FROM )
  );
  defparam \DLX_IDinst_slot_num_FFd4-In30_SW0 .INIT = 16'hFBF0;
  X_LUT4 \DLX_IDinst_slot_num_FFd4-In30_SW0  (
    .ADR0(DLX_IDinst_CLI),
    .ADR1(INT_IBUF),
    .ADR2(FREEZE_IBUF),
    .ADR3(N147200),
    .O(\N147200/GROM )
  );
  X_BUF \N147200/XUSED  (
    .I(\N147200/FROM ),
    .O(N147200)
  );
  X_BUF \N147200/YUSED  (
    .I(\N147200/GROM ),
    .O(N164719)
  );
  defparam DLX_IDinst__n0381_1475.INIT = 16'h0001;
  X_LUT4 DLX_IDinst__n0381_1475 (
    .ADR0(DLX_IDinst_jtarget[20]),
    .ADR1(DLX_IDinst_jtarget[19]),
    .ADR2(N126925),
    .ADR3(DLX_IDinst_jtarget[18]),
    .O(\DLX_IDinst__n0381/FROM )
  );
  defparam DLX_IDinst_Ker1084941.INIT = 16'hCC44;
  X_LUT4 DLX_IDinst_Ker1084941 (
    .ADR0(DLX_IDinst__n0105),
    .ADR1(DLX_IDinst_N108152),
    .ADR2(VCC),
    .ADR3(DLX_IDinst__n0381),
    .O(\DLX_IDinst__n0381/GROM )
  );
  X_BUF \DLX_IDinst__n0381/XUSED  (
    .I(\DLX_IDinst__n0381/FROM ),
    .O(DLX_IDinst__n0381)
  );
  X_BUF \DLX_IDinst__n0381/YUSED  (
    .I(\DLX_IDinst__n0381/GROM ),
    .O(DLX_IDinst_N108496)
  );
  defparam DLX_IDinst_Ker107397112.INIT = 16'h5450;
  X_LUT4 DLX_IDinst_Ker107397112 (
    .ADR0(DLX_IDinst_IR_opcode_field[5]),
    .ADR1(CHOICE1338),
    .ADR2(CHOICE1346),
    .ADR3(DLX_IDinst_IR_opcode_field[3]),
    .O(\CHOICE1348/FROM )
  );
  defparam DLX_IDinst_Ker107397126.INIT = 16'hFF54;
  X_LUT4 DLX_IDinst_Ker107397126 (
    .ADR0(DLX_IDinst_IR_opcode_field[3]),
    .ADR1(CHOICE1327),
    .ADR2(CHOICE1320),
    .ADR3(CHOICE1348),
    .O(\CHOICE1348/GROM )
  );
  X_BUF \CHOICE1348/XUSED  (
    .I(\CHOICE1348/FROM ),
    .O(CHOICE1348)
  );
  X_BUF \CHOICE1348/YUSED  (
    .I(\CHOICE1348/GROM ),
    .O(N135079)
  );
  X_ONE \vga_top_vga1_videoon/LOGIC_ONE_1476  (
    .O(\vga_top_vga1_videoon/LOGIC_ONE )
  );
  defparam \vga_top_vga1_blueout<1>1 .INIT = 16'h0404;
  X_LUT4 \vga_top_vga1_blueout<1>1  (
    .ADR0(reset_IBUF_1),
    .ADR1(vga_top_vga1_videoon),
    .ADR2(vram_out_vga_eff),
    .ADR3(VCC),
    .O(\vga_top_vga1_videoon/FROM )
  );
  defparam \vga_top_vga1_greenout<1>1 .INIT = 16'h0404;
  X_LUT4 \vga_top_vga1_greenout<1>1  (
    .ADR0(reset_IBUF_1),
    .ADR1(vga_top_vga1_videoon),
    .ADR2(vram_out_vga_eff),
    .ADR3(VCC),
    .O(\vga_top_vga1_videoon/GROM )
  );
  X_BUF \vga_top_vga1_videoon/XUSED  (
    .I(\vga_top_vga1_videoon/FROM ),
    .O(blue_1_OBUF)
  );
  X_BUF \vga_top_vga1_videoon/YUSED  (
    .I(\vga_top_vga1_videoon/GROM ),
    .O(green_1_OBUF)
  );
  defparam \DLX_EXinst__n0007<25>223_SW0 .INIT = 16'hFCF0;
  X_LUT4 \DLX_EXinst__n0007<25>223_SW0  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst__n0081),
    .ADR2(CHOICE5108),
    .ADR3(\DLX_EXinst_Mshift__n0024_Sh[57] ),
    .O(\N163534/FROM )
  );
  defparam \DLX_EXinst__n0007<25>223 .INIT = 16'hD5C0;
  X_LUT4 \DLX_EXinst__n0007<25>223  (
    .ADR0(N148323),
    .ADR1(N148609),
    .ADR2(N138591),
    .ADR3(N163534),
    .O(\N163534/GROM )
  );
  X_BUF \N163534/XUSED  (
    .I(\N163534/FROM ),
    .O(N163534)
  );
  X_BUF \N163534/YUSED  (
    .I(\N163534/GROM ),
    .O(CHOICE5113)
  );
  defparam DLX_IDinst_Ker1084541_1_1477.INIT = 16'h8800;
  X_LUT4 DLX_IDinst_Ker1084541_1_1477 (
    .ADR0(DLX_IDinst_IR_latched[26]),
    .ADR1(DLX_IDinst_N108165),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_IR_latched[27]),
    .O(\DLX_IDinst_Ker1084541_1/FROM )
  );
  defparam \DLX_IDinst__n0145<0>37 .INIT = 16'h0032;
  X_LUT4 \DLX_IDinst__n0145<0>37  (
    .ADR0(DLX_IDinst__n0167),
    .ADR1(DLX_IDinst__n0387),
    .ADR2(DLX_IDinst__n0166),
    .ADR3(DLX_IDinst_Ker1084541_1),
    .O(\DLX_IDinst_Ker1084541_1/GROM )
  );
  X_BUF \DLX_IDinst_Ker1084541_1/XUSED  (
    .I(\DLX_IDinst_Ker1084541_1/FROM ),
    .O(DLX_IDinst_Ker1084541_1)
  );
  X_BUF \DLX_IDinst_Ker1084541_1/YUSED  (
    .I(\DLX_IDinst_Ker1084541_1/GROM ),
    .O(CHOICE2918)
  );
  defparam DLX_IDinst_RegFile_27_19_1478.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_27_19_1478 (
    .I(DLX_IDinst_WB_data_eff[19]),
    .CE(DLX_IDinst__n0604),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_27_19)
  );
  defparam \DLX_EXinst__n0007<25>139_SW0 .INIT = 16'hFFFA;
  X_LUT4 \DLX_EXinst__n0007<25>139_SW0  (
    .ADR0(CHOICE5058),
    .ADR1(VCC),
    .ADR2(CHOICE5063),
    .ADR3(CHOICE5083),
    .O(\N163602/FROM )
  );
  defparam \DLX_EXinst__n0007<25>139 .INIT = 16'h0F08;
  X_LUT4 \DLX_EXinst__n0007<25>139  (
    .ADR0(\DLX_EXinst_Mshift__n0021_Sh[41] ),
    .ADR1(DLX_EXinst_N75993),
    .ADR2(DLX_EXinst__n0036),
    .ADR3(N163602),
    .O(\N163602/GROM )
  );
  X_BUF \N163602/XUSED  (
    .I(\N163602/FROM ),
    .O(N163602)
  );
  X_BUF \N163602/YUSED  (
    .I(\N163602/GROM ),
    .O(CHOICE5087)
  );
  defparam \DM_read_data<9>1 .INIT = 16'hAA04;
  X_LUT4 \DM_read_data<9>1  (
    .ADR0(DLX_EXinst_ALU_result[13]),
    .ADR1(RAM_read_data[9]),
    .ADR2(DLX_EXinst_ALU_result[12]),
    .ADR3(DLX_EXinst_ALU_result[14]),
    .O(\DM_read_data<9>/FROM )
  );
  defparam \DM_read_data<8>1 .INIT = 16'hC0C2;
  X_LUT4 \DM_read_data<8>1  (
    .ADR0(RAM_read_data[8]),
    .ADR1(DLX_EXinst_ALU_result[14]),
    .ADR2(DLX_EXinst_ALU_result[13]),
    .ADR3(DLX_EXinst_ALU_result[12]),
    .O(\DM_read_data<9>/GROM )
  );
  X_BUF \DM_read_data<9>/XUSED  (
    .I(\DM_read_data<9>/FROM ),
    .O(DM_read_data[9])
  );
  X_BUF \DM_read_data<9>/YUSED  (
    .I(\DM_read_data<9>/GROM ),
    .O(DM_read_data[8])
  );
  defparam \DLX_EXinst__n0007<17>179_SW0 .INIT = 16'hAEAA;
  X_LUT4 \DLX_EXinst__n0007<17>179_SW0  (
    .ADR0(CHOICE5354),
    .ADR1(\DLX_EXinst_Mshift__n0021_Sh[1] ),
    .ADR2(DLX_EXinst_N72815),
    .ADR3(DLX_EXinst_N75993),
    .O(\N163627/FROM )
  );
  defparam \DLX_EXinst__n0007<17>179 .INIT = 16'h3332;
  X_LUT4 \DLX_EXinst__n0007<17>179  (
    .ADR0(CHOICE5361),
    .ADR1(DLX_EXinst__n0036),
    .ADR2(CHOICE5385),
    .ADR3(N163627),
    .O(\N163627/GROM )
  );
  X_BUF \N163627/XUSED  (
    .I(\N163627/FROM ),
    .O(N163627)
  );
  X_BUF \N163627/YUSED  (
    .I(\N163627/GROM ),
    .O(CHOICE5389)
  );
  defparam \DLX_EXinst__n0007<26>223_SW0 .INIT = 16'hFCF0;
  X_LUT4 \DLX_EXinst__n0007<26>223_SW0  (
    .ADR0(VCC),
    .ADR1(\DLX_EXinst_Mshift__n0024_Sh[58] ),
    .ADR2(CHOICE5041),
    .ADR3(DLX_EXinst__n0081),
    .O(\N163692/FROM )
  );
  defparam \DLX_EXinst__n0007<26>223 .INIT = 16'hD5C0;
  X_LUT4 \DLX_EXinst__n0007<26>223  (
    .ADR0(N148323),
    .ADR1(N138249),
    .ADR2(N148609),
    .ADR3(N163692),
    .O(\N163692/GROM )
  );
  X_BUF \N163692/XUSED  (
    .I(\N163692/FROM ),
    .O(N163692)
  );
  X_BUF \N163692/YUSED  (
    .I(\N163692/GROM ),
    .O(CHOICE5046)
  );
  defparam \DLX_IDinst__n0114<6>6 .INIT = 16'hEAC0;
  X_LUT4 \DLX_IDinst__n0114<6>6  (
    .ADR0(DLX_IDinst__n0098),
    .ADR1(DLX_IDinst_N108305),
    .ADR2(DLX_IDinst_branch_address[6]),
    .ADR3(DLX_IDinst_EPC[6]),
    .O(\DLX_IDinst_EPC<1>/FROM )
  );
  defparam \DLX_IDinst__n0114<1>6 .INIT = 16'hECA0;
  X_LUT4 \DLX_IDinst__n0114<1>6  (
    .ADR0(DLX_IDinst_N108305),
    .ADR1(DLX_IDinst__n0098),
    .ADR2(DLX_IDinst_branch_address[1]),
    .ADR3(DLX_IDinst_EPC[1]),
    .O(\DLX_IDinst_EPC<1>/GROM )
  );
  X_BUF \DLX_IDinst_EPC<1>/XUSED  (
    .I(\DLX_IDinst_EPC<1>/FROM ),
    .O(CHOICE3185)
  );
  X_BUF \DLX_IDinst_EPC<1>/YUSED  (
    .I(\DLX_IDinst_EPC<1>/GROM ),
    .O(CHOICE2144)
  );
  defparam \DLX_IDinst__n0114<7>4 .INIT = 16'hFF88;
  X_LUT4 \DLX_IDinst__n0114<7>4  (
    .ADR0(DLX_IDinst__n0098),
    .ADR1(DLX_IDinst_EPC[7]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst__n0453),
    .O(\DLX_IDinst_EPC<7>/FROM )
  );
  defparam \DLX_IDinst__n0114<7>12 .INIT = 16'h3320;
  X_LUT4 \DLX_IDinst__n0114<7>12  (
    .ADR0(DLX_IDinst_branch_address[7]),
    .ADR1(DLX_IDinst_N108456),
    .ADR2(DLX_IDinst_N108305),
    .ADR3(CHOICE2198),
    .O(\DLX_IDinst_EPC<7>/GROM )
  );
  X_BUF \DLX_IDinst_EPC<7>/XUSED  (
    .I(\DLX_IDinst_EPC<7>/FROM ),
    .O(CHOICE2198)
  );
  X_BUF \DLX_IDinst_EPC<7>/YUSED  (
    .I(\DLX_IDinst_EPC<7>/GROM ),
    .O(CHOICE2200)
  );
  defparam DLX_IDinst_RegFile_28_11_1479.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_28_11_1479 (
    .I(DLX_IDinst_WB_data_eff[11]),
    .CE(DLX_IDinst__n0606),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_28_11)
  );
  defparam DLX_IDinst__n0137152_SW0.INIT = 16'hCCF0;
  X_LUT4 DLX_IDinst__n0137152_SW0 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst__n0629[1]),
    .ADR2(DLX_IDinst__n0098),
    .ADR3(DLX_IDinst__n0453),
    .O(\DLX_IDinst_EPC<8>/FROM )
  );
  defparam \DLX_IDinst__n0114<8>6 .INIT = 16'hF888;
  X_LUT4 \DLX_IDinst__n0114<8>6  (
    .ADR0(DLX_IDinst_branch_address[8]),
    .ADR1(DLX_IDinst_N108305),
    .ADR2(DLX_IDinst__n0098),
    .ADR3(DLX_IDinst_EPC[8]),
    .O(\DLX_IDinst_EPC<8>/GROM )
  );
  X_BUF \DLX_IDinst_EPC<8>/XUSED  (
    .I(\DLX_IDinst_EPC<8>/FROM ),
    .O(N163190)
  );
  X_BUF \DLX_IDinst_EPC<8>/YUSED  (
    .I(\DLX_IDinst_EPC<8>/GROM ),
    .O(CHOICE2209)
  );
  defparam \DLX_EXinst__n0007<1>3321_SW0 .INIT = 16'hFEEE;
  X_LUT4 \DLX_EXinst__n0007<1>3321_SW0  (
    .ADR0(CHOICE5758),
    .ADR1(N164573),
    .ADR2(DLX_IDinst_reg_out_A[2]),
    .ADR3(DLX_EXinst_N74136),
    .O(\DLX_EXinst_ALU_result<1>/FROM )
  );
  defparam \DLX_EXinst__n0007<1>3321 .INIT = 16'hFFEA;
  X_LUT4 \DLX_EXinst__n0007<1>3321  (
    .ADR0(N136886),
    .ADR1(DLX_EXinst__n0012[1]),
    .ADR2(DLX_EXinst_N73959),
    .ADR3(N163270),
    .O(\DLX_EXinst_ALU_result<1>/GROM )
  );
  X_BUF \DLX_EXinst_ALU_result<1>/XUSED  (
    .I(\DLX_EXinst_ALU_result<1>/FROM ),
    .O(N163270)
  );
  X_BUF \DLX_EXinst_ALU_result<1>/YUSED  (
    .I(\DLX_EXinst_ALU_result<1>/GROM ),
    .O(N162854)
  );
  defparam vga_top_vga1_Ker112929.INIT = 16'h1000;
  X_LUT4 vga_top_vga1_Ker112929 (
    .ADR0(N136748),
    .ADR1(vga_top_vga1_vcounter[0]),
    .ADR2(vga_top_vga1_N112936),
    .ADR3(vga_top_vga1_vcounter[1]),
    .O(\vga_top_vga1_N112931/FROM )
  );
  defparam vga_top_vga1__n0014_SW0.INIT = 16'hF3FF;
  X_LUT4 vga_top_vga1__n0014_SW0 (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_N112941),
    .ADR2(vga_top_vga1_vcounter[9]),
    .ADR3(vga_top_vga1_N112931),
    .O(\vga_top_vga1_N112931/GROM )
  );
  X_BUF \vga_top_vga1_N112931/XUSED  (
    .I(\vga_top_vga1_N112931/FROM ),
    .O(vga_top_vga1_N112931)
  );
  X_BUF \vga_top_vga1_N112931/YUSED  (
    .I(\vga_top_vga1_N112931/GROM ),
    .O(N132456)
  );
  defparam \DLX_EXinst__n0007<18>179_SW0 .INIT = 16'hF2F0;
  X_LUT4 \DLX_EXinst__n0007<18>179_SW0  (
    .ADR0(\DLX_EXinst_Mshift__n0021_Sh[2] ),
    .ADR1(DLX_EXinst_N72815),
    .ADR2(CHOICE5196),
    .ADR3(DLX_EXinst_N75993),
    .O(\N163407/FROM )
  );
  defparam \DLX_EXinst__n0007<18>179 .INIT = 16'h0F0E;
  X_LUT4 \DLX_EXinst__n0007<18>179  (
    .ADR0(CHOICE5203),
    .ADR1(CHOICE5227),
    .ADR2(DLX_EXinst__n0036),
    .ADR3(N163407),
    .O(\N163407/GROM )
  );
  X_BUF \N163407/XUSED  (
    .I(\N163407/FROM ),
    .O(N163407)
  );
  X_BUF \N163407/YUSED  (
    .I(\N163407/GROM ),
    .O(CHOICE5231)
  );
  defparam \DLX_IDinst__n0018<0>1 .INIT = 16'hEC00;
  X_LUT4 \DLX_IDinst__n0018<0>1  (
    .ADR0(N139656),
    .ADR1(DLX_IDinst__n0453),
    .ADR2(DLX_IDinst_N107033),
    .ADR3(DLX_IDinst_jtarget[11]),
    .O(\DLX_IDinst_rd_addr<0>/FROM )
  );
  defparam \DLX_IDinst__n0136<0>1 .INIT = 16'hFF80;
  X_LUT4 \DLX_IDinst__n0136<0>1  (
    .ADR0(DLX_IDinst_IR_latched[26]),
    .ADR1(DLX_IDinst_IR_latched[27]),
    .ADR2(DLX_IDinst_N108165),
    .ADR3(DLX_IDinst__n0018[0]),
    .O(DLX_IDinst__n0136[0])
  );
  X_BUF \DLX_IDinst_rd_addr<0>/XUSED  (
    .I(\DLX_IDinst_rd_addr<0>/FROM ),
    .O(DLX_IDinst__n0018[0])
  );
  defparam \DLX_IDinst__n0018<1>1 .INIT = 16'hC888;
  X_LUT4 \DLX_IDinst__n0018<1>1  (
    .ADR0(DLX_IDinst__n0453),
    .ADR1(DLX_IDinst_jtarget[12]),
    .ADR2(N139656),
    .ADR3(DLX_IDinst_N107033),
    .O(\DLX_IDinst_rd_addr<1>/FROM )
  );
  defparam \DLX_IDinst__n0136<1>1 .INIT = 16'hFF80;
  X_LUT4 \DLX_IDinst__n0136<1>1  (
    .ADR0(DLX_IDinst_N108165),
    .ADR1(DLX_IDinst_IR_latched[27]),
    .ADR2(DLX_IDinst_IR_latched[26]),
    .ADR3(DLX_IDinst__n0018[1]),
    .O(DLX_IDinst__n0136[1])
  );
  X_BUF \DLX_IDinst_rd_addr<1>/XUSED  (
    .I(\DLX_IDinst_rd_addr<1>/FROM ),
    .O(DLX_IDinst__n0018[1])
  );
  defparam \DLX_IDinst__n0025<5>1 .INIT = 16'hA8A0;
  X_LUT4 \DLX_IDinst__n0025<5>1  (
    .ADR0(DLX_IDinst_jtarget[5]),
    .ADR1(DLX_IDinst_N107033),
    .ADR2(DLX_IDinst__n0453),
    .ADR3(N139656),
    .O(\DLX_IDinst_Imm<5>/FROM )
  );
  defparam DLX_IDinst__n01291.INIT = 16'h7F00;
  X_LUT4 DLX_IDinst__n01291 (
    .ADR0(DLX_IDinst_IR_latched[27]),
    .ADR1(DLX_IDinst_N108165),
    .ADR2(DLX_IDinst_IR_latched[26]),
    .ADR3(DLX_IDinst__n0025[5]),
    .O(DLX_IDinst__n0129)
  );
  X_BUF \DLX_IDinst_Imm<5>/XUSED  (
    .I(\DLX_IDinst_Imm<5>/FROM ),
    .O(DLX_IDinst__n0025[5])
  );
  defparam \DLX_IDinst__n0018<2>1 .INIT = 16'hA8A0;
  X_LUT4 \DLX_IDinst__n0018<2>1  (
    .ADR0(DLX_IDinst_jtarget[13]),
    .ADR1(N139656),
    .ADR2(DLX_IDinst__n0453),
    .ADR3(DLX_IDinst_N107033),
    .O(\DLX_IDinst_rd_addr<2>/FROM )
  );
  defparam \DLX_IDinst__n0136<2>1 .INIT = 16'hFF80;
  X_LUT4 \DLX_IDinst__n0136<2>1  (
    .ADR0(DLX_IDinst_N108165),
    .ADR1(DLX_IDinst_IR_latched[26]),
    .ADR2(DLX_IDinst_IR_latched[27]),
    .ADR3(DLX_IDinst__n0018[2]),
    .O(DLX_IDinst__n0136[2])
  );
  X_BUF \DLX_IDinst_rd_addr<2>/XUSED  (
    .I(\DLX_IDinst_rd_addr<2>/FROM ),
    .O(DLX_IDinst__n0018[2])
  );
  defparam DLX_EXinst_Ker760001.INIT = 16'h0044;
  X_LUT4 DLX_EXinst_Ker760001 (
    .ADR0(DLX_IDinst_Imm_3_1),
    .ADR1(DLX_IDinst_Imm_2_1),
    .ADR2(VCC),
    .ADR3(\DLX_IDinst_Imm[4] ),
    .O(\DLX_EXinst_N76002/FROM )
  );
  defparam DLX_EXinst__n00811.INIT = 16'h0400;
  X_LUT4 DLX_EXinst__n00811 (
    .ADR0(\DLX_IDinst_Imm[0] ),
    .ADR1(\DLX_IDinst_Imm[1] ),
    .ADR2(DLX_IDinst_IR_function_field[5]),
    .ADR3(DLX_EXinst_N76002),
    .O(\DLX_EXinst_N76002/GROM )
  );
  X_BUF \DLX_EXinst_N76002/XUSED  (
    .I(\DLX_EXinst_N76002/FROM ),
    .O(DLX_EXinst_N76002)
  );
  X_BUF \DLX_EXinst_N76002/YUSED  (
    .I(\DLX_EXinst_N76002/GROM ),
    .O(DLX_EXinst__n0081)
  );
  defparam DLX_EXinst_Ker738951.INIT = 16'hACAC;
  X_LUT4 DLX_EXinst_Ker738951 (
    .ADR0(DLX_IDinst_reg_out_A[26]),
    .ADR1(DLX_IDinst_reg_out_A[24]),
    .ADR2(DLX_IDinst_Imm_1_1),
    .ADR3(VCC),
    .O(\DLX_EXinst_N73897/FROM )
  );
  defparam DLX_EXinst_Ker733521.INIT = 16'hCACA;
  X_LUT4 DLX_EXinst_Ker733521 (
    .ADR0(DLX_IDinst_reg_out_A[26]),
    .ADR1(DLX_IDinst_reg_out_A[24]),
    .ADR2(DLX_IDinst_reg_out_B[1]),
    .ADR3(VCC),
    .O(\DLX_EXinst_N73897/GROM )
  );
  X_BUF \DLX_EXinst_N73897/XUSED  (
    .I(\DLX_EXinst_N73897/FROM ),
    .O(DLX_EXinst_N73897)
  );
  X_BUF \DLX_EXinst_N73897/YUSED  (
    .I(\DLX_EXinst_N73897/GROM ),
    .O(DLX_EXinst_N73354)
  );
  defparam DLX_EXinst_Ker732651.INIT = 16'hFF0A;
  X_LUT4 DLX_EXinst_Ker732651 (
    .ADR0(N147520),
    .ADR1(VCC),
    .ADR2(\DLX_IDinst_Imm[5] ),
    .ADR3(DLX_EXinst_N76441),
    .O(\DLX_EXinst_N73267/FROM )
  );
  defparam \DLX_EXinst__n0007<4>163 .INIT = 16'hAC00;
  X_LUT4 \DLX_EXinst__n0007<4>163  (
    .ADR0(DLX_EXinst_N74946),
    .ADR1(N137680),
    .ADR2(\DLX_IDinst_Imm[2] ),
    .ADR3(DLX_EXinst_N73267),
    .O(\DLX_EXinst_N73267/GROM )
  );
  X_BUF \DLX_EXinst_N73267/XUSED  (
    .I(\DLX_EXinst_N73267/FROM ),
    .O(DLX_EXinst_N73267)
  );
  X_BUF \DLX_EXinst_N73267/YUSED  (
    .I(\DLX_EXinst_N73267/GROM ),
    .O(CHOICE4360)
  );
  defparam DLX_EXinst_Ker728011.INIT = 16'hFC30;
  X_LUT4 DLX_EXinst_Ker728011 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_B[0]),
    .ADR2(DLX_IDinst_reg_out_A[29]),
    .ADR3(DLX_IDinst_reg_out_A[30]),
    .O(\DLX_EXinst_N72803/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0024_Sh<29>1 .INIT = 16'h4F40;
  X_LUT4 \DLX_EXinst_Mshift__n0024_Sh<29>1  (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(DLX_IDinst_reg_out_A[31]),
    .ADR2(DLX_IDinst_reg_out_B[1]),
    .ADR3(DLX_EXinst_N72803),
    .O(\DLX_EXinst_N72803/GROM )
  );
  X_BUF \DLX_EXinst_N72803/XUSED  (
    .I(\DLX_EXinst_N72803/FROM ),
    .O(DLX_EXinst_N72803)
  );
  X_BUF \DLX_EXinst_N72803/YUSED  (
    .I(\DLX_EXinst_N72803/GROM ),
    .O(\DLX_EXinst_Mshift__n0024_Sh[29] )
  );
  defparam DLX_EXinst_Ker736021.INIT = 16'hF5A0;
  X_LUT4 DLX_EXinst_Ker736021 (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[6]),
    .ADR3(DLX_IDinst_reg_out_A[8]),
    .O(\DLX_EXinst_N73604/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<9>1 .INIT = 16'hEE44;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<9>1  (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(DLX_EXinst_N72853),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N73604),
    .O(\DLX_EXinst_N73604/GROM )
  );
  X_BUF \DLX_EXinst_N73604/XUSED  (
    .I(\DLX_EXinst_N73604/FROM ),
    .O(DLX_EXinst_N73604)
  );
  X_BUF \DLX_EXinst_N73604/YUSED  (
    .I(\DLX_EXinst_N73604/GROM ),
    .O(\DLX_EXinst_Mshift__n0023_Sh[9] )
  );
  defparam DLX_EXinst_Ker735221.INIT = 16'hBB88;
  X_LUT4 DLX_EXinst_Ker735221 (
    .ADR0(DLX_IDinst_reg_out_A[16]),
    .ADR1(DLX_IDinst_Imm_1_1),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[14]),
    .O(\DLX_EXinst_N73524/FROM )
  );
  defparam DLX_EXinst_Ker74709_SW0.INIT = 16'hFC30;
  X_LUT4 DLX_EXinst_Ker74709_SW0 (
    .ADR0(VCC),
    .ADR1(\DLX_IDinst_Imm[0] ),
    .ADR2(DLX_EXinst_N73128),
    .ADR3(DLX_EXinst_N73524),
    .O(\DLX_EXinst_N73524/GROM )
  );
  X_BUF \DLX_EXinst_N73524/XUSED  (
    .I(\DLX_EXinst_N73524/FROM ),
    .O(DLX_EXinst_N73524)
  );
  X_BUF \DLX_EXinst_N73524/YUSED  (
    .I(\DLX_EXinst_N73524/GROM ),
    .O(N130773)
  );
  defparam DLX_EXinst_Ker742431.INIT = 16'hFFAA;
  X_LUT4 DLX_EXinst_Ker742431 (
    .ADR0(DLX_EXinst__n0078),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_EXinst__n0083),
    .O(\DLX_EXinst_N74245/FROM )
  );
  defparam \DLX_EXinst__n0007<29>242 .INIT = 16'hFFB8;
  X_LUT4 \DLX_EXinst__n0007<29>242  (
    .ADR0(DLX_EXinst__n0077),
    .ADR1(DLX_IDinst_reg_out_B[29]),
    .ADR2(DLX_EXinst__n0079),
    .ADR3(DLX_EXinst_N74245),
    .O(\DLX_EXinst_N74245/GROM )
  );
  X_BUF \DLX_EXinst_N74245/XUSED  (
    .I(\DLX_EXinst_N74245/FROM ),
    .O(DLX_EXinst_N74245)
  );
  X_BUF \DLX_EXinst_N74245/YUSED  (
    .I(\DLX_EXinst_N74245/GROM ),
    .O(CHOICE4831)
  );
  defparam DLX_EXinst_Ker735521.INIT = 16'hE4E4;
  X_LUT4 DLX_EXinst_Ker735521 (
    .ADR0(DLX_IDinst_Imm_1_1),
    .ADR1(DLX_IDinst_reg_out_A[8]),
    .ADR2(DLX_IDinst_reg_out_A[10]),
    .ADR3(VCC),
    .O(\DLX_EXinst_N73554/FROM )
  );
  defparam DLX_EXinst_Ker734271.INIT = 16'hFA0A;
  X_LUT4 DLX_EXinst_Ker734271 (
    .ADR0(DLX_IDinst_reg_out_A[8]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[1]),
    .ADR3(DLX_IDinst_reg_out_A[10]),
    .O(\DLX_EXinst_N73554/GROM )
  );
  X_BUF \DLX_EXinst_N73554/XUSED  (
    .I(\DLX_EXinst_N73554/FROM ),
    .O(DLX_EXinst_N73554)
  );
  X_BUF \DLX_EXinst_N73554/YUSED  (
    .I(\DLX_EXinst_N73554/GROM ),
    .O(DLX_EXinst_N73429)
  );
  defparam DLX_EXinst_Ker735071.INIT = 16'hFC30;
  X_LUT4 DLX_EXinst_Ker735071 (
    .ADR0(VCC),
    .ADR1(\DLX_IDinst_Imm[1] ),
    .ADR2(DLX_IDinst_reg_out_A[8]),
    .ADR3(DLX_IDinst_reg_out_A[6]),
    .O(\DLX_EXinst_N73509/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0021_Sh<9>1 .INIT = 16'hEE44;
  X_LUT4 \DLX_EXinst_Mshift__n0021_Sh<9>1  (
    .ADR0(DLX_IDinst_Imm_0_1),
    .ADR1(DLX_EXinst_N72938),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N73509),
    .O(\DLX_EXinst_N73509/GROM )
  );
  X_BUF \DLX_EXinst_N73509/XUSED  (
    .I(\DLX_EXinst_N73509/FROM ),
    .O(DLX_EXinst_N73509)
  );
  X_BUF \DLX_EXinst_N73509/YUSED  (
    .I(\DLX_EXinst_N73509/GROM ),
    .O(\DLX_EXinst_Mshift__n0021_Sh[9] )
  );
  defparam DLX_EXinst_Ker728201.INIT = 16'hFAFA;
  X_LUT4 DLX_EXinst_Ker728201 (
    .ADR0(DLX_IDinst_reg_out_B[2]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[3]),
    .ADR3(VCC),
    .O(\DLX_EXinst_N72822/FROM )
  );
  defparam DLX_EXinst_Ker7550830.INIT = 16'h30E2;
  X_LUT4 DLX_EXinst_Ker7550830 (
    .ADR0(\DLX_EXinst_Mshift__n0019_Sh[28] ),
    .ADR1(DLX_IDinst_reg_out_B[5]),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(DLX_EXinst_N72822),
    .O(\DLX_EXinst_N72822/GROM )
  );
  X_BUF \DLX_EXinst_N72822/XUSED  (
    .I(\DLX_EXinst_N72822/FROM ),
    .O(DLX_EXinst_N72822)
  );
  X_BUF \DLX_EXinst_N72822/YUSED  (
    .I(\DLX_EXinst_N72822/GROM ),
    .O(CHOICE1276)
  );
  defparam DLX_EXinst_Ker727081.INIT = 16'hAAEE;
  X_LUT4 DLX_EXinst_Ker727081 (
    .ADR0(DLX_EXinst_N76421),
    .ADR1(N148609),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[5]),
    .O(\DLX_EXinst_N72710/FROM )
  );
  defparam \DLX_EXinst__n0007<4>70 .INIT = 16'hD800;
  X_LUT4 \DLX_EXinst__n0007<4>70  (
    .ADR0(DLX_IDinst_reg_out_B[2]),
    .ADR1(DLX_EXinst_N74691),
    .ADR2(N137448),
    .ADR3(DLX_EXinst_N72710),
    .O(\DLX_EXinst_N72710/GROM )
  );
  X_BUF \DLX_EXinst_N72710/XUSED  (
    .I(\DLX_EXinst_N72710/FROM ),
    .O(DLX_EXinst_N72710)
  );
  X_BUF \DLX_EXinst_N72710/YUSED  (
    .I(\DLX_EXinst_N72710/GROM ),
    .O(CHOICE4341)
  );
  defparam DLX_EXinst_Ker734621.INIT = 16'hAFA0;
  X_LUT4 DLX_EXinst_Ker734621 (
    .ADR0(DLX_IDinst_reg_out_A[8]),
    .ADR1(VCC),
    .ADR2(\DLX_IDinst_Imm[1] ),
    .ADR3(DLX_IDinst_reg_out_A[10]),
    .O(\DLX_EXinst_N73464/FROM )
  );
  defparam DLX_EXinst_Ker733721.INIT = 16'hFA0A;
  X_LUT4 DLX_EXinst_Ker733721 (
    .ADR0(DLX_IDinst_reg_out_A[26]),
    .ADR1(VCC),
    .ADR2(\DLX_IDinst_Imm[1] ),
    .ADR3(DLX_IDinst_reg_out_A[24]),
    .O(\DLX_EXinst_N73464/GROM )
  );
  X_BUF \DLX_EXinst_N73464/XUSED  (
    .I(\DLX_EXinst_N73464/FROM ),
    .O(DLX_EXinst_N73464)
  );
  X_BUF \DLX_EXinst_N73464/YUSED  (
    .I(\DLX_EXinst_N73464/GROM ),
    .O(DLX_EXinst_N73374)
  );
  defparam DLX_EXinst_Ker735171.INIT = 16'hFA0A;
  X_LUT4 DLX_EXinst_Ker735171 (
    .ADR0(DLX_IDinst_reg_out_A[12]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_Imm_1_1),
    .ADR3(DLX_IDinst_reg_out_A[14]),
    .O(\DLX_EXinst_N73519/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0022_Sh<11>1 .INIT = 16'hFA0A;
  X_LUT4 \DLX_EXinst_Mshift__n0022_Sh<11>1  (
    .ADR0(DLX_EXinst_N73123),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_Imm_0_1),
    .ADR3(DLX_EXinst_N73519),
    .O(\DLX_EXinst_N73519/GROM )
  );
  X_BUF \DLX_EXinst_N73519/XUSED  (
    .I(\DLX_EXinst_N73519/FROM ),
    .O(DLX_EXinst_N73519)
  );
  X_BUF \DLX_EXinst_N73519/YUSED  (
    .I(\DLX_EXinst_N73519/GROM ),
    .O(\DLX_EXinst_Mshift__n0022_Sh[11] )
  );
  defparam DLX_EXinst_Ker728131.INIT = 16'hEEEE;
  X_LUT4 DLX_EXinst_Ker728131 (
    .ADR0(\DLX_IDinst_Imm[2] ),
    .ADR1(\DLX_IDinst_Imm[3] ),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_EXinst_N72815/FROM )
  );
  defparam DLX_EXinst_Ker7565230.INIT = 16'h7610;
  X_LUT4 DLX_EXinst_Ker7565230 (
    .ADR0(\DLX_IDinst_Imm[5] ),
    .ADR1(DLX_EXinst_N72815),
    .ADR2(\DLX_EXinst_Mshift__n0020_Sh[28] ),
    .ADR3(DLX_IDinst_reg_out_A[31]),
    .O(\DLX_EXinst_N72815/GROM )
  );
  X_BUF \DLX_EXinst_N72815/XUSED  (
    .I(\DLX_EXinst_N72815/FROM ),
    .O(DLX_EXinst_N72815)
  );
  X_BUF \DLX_EXinst_N72815/YUSED  (
    .I(\DLX_EXinst_N72815/GROM ),
    .O(CHOICE1291)
  );
  defparam DLX_EXinst_Ker735421.INIT = 16'hFC0C;
  X_LUT4 DLX_EXinst_Ker735421 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[22]),
    .ADR2(DLX_IDinst_Imm_1_1),
    .ADR3(DLX_IDinst_reg_out_A[24]),
    .O(\DLX_EXinst_N73544/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0022_Sh<21>1 .INIT = 16'hFC0C;
  X_LUT4 \DLX_EXinst_Mshift__n0022_Sh<21>1  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N73148),
    .ADR2(DLX_IDinst_Imm_0_1),
    .ADR3(DLX_EXinst_N73544),
    .O(\DLX_EXinst_N73544/GROM )
  );
  X_BUF \DLX_EXinst_N73544/XUSED  (
    .I(\DLX_EXinst_N73544/FROM ),
    .O(DLX_EXinst_N73544)
  );
  X_BUF \DLX_EXinst_N73544/YUSED  (
    .I(\DLX_EXinst_N73544/GROM ),
    .O(\DLX_EXinst_Mshift__n0022_Sh[21] )
  );
  defparam DLX_EXinst_Ker733821.INIT = 16'hCCAA;
  X_LUT4 DLX_EXinst_Ker733821 (
    .ADR0(DLX_IDinst_reg_out_A[10]),
    .ADR1(DLX_IDinst_reg_out_A[12]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[1]),
    .O(\DLX_EXinst_N73384/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0019_Sh<9>1 .INIT = 16'hFC0C;
  X_LUT4 \DLX_EXinst_Mshift__n0019_Sh<9>1  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N73033),
    .ADR2(DLX_IDinst_reg_out_B[0]),
    .ADR3(DLX_EXinst_N73384),
    .O(\DLX_EXinst_N73384/GROM )
  );
  X_BUF \DLX_EXinst_N73384/XUSED  (
    .I(\DLX_EXinst_N73384/FROM ),
    .O(DLX_EXinst_N73384)
  );
  X_BUF \DLX_EXinst_N73384/YUSED  (
    .I(\DLX_EXinst_N73384/GROM ),
    .O(\DLX_EXinst_Mshift__n0019_Sh[9] )
  );
  defparam DLX_EXinst_Ker728071.INIT = 16'hCACA;
  X_LUT4 DLX_EXinst_Ker728071 (
    .ADR0(\DLX_EXinst_Mshift__n0019_Sh[20] ),
    .ADR1(\DLX_EXinst_Mshift__n0019_Sh[28] ),
    .ADR2(DLX_IDinst_reg_out_B[3]),
    .ADR3(VCC),
    .O(\DLX_EXinst_N72809/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0024_Sh<52>1 .INIT = 16'h7340;
  X_LUT4 \DLX_EXinst_Mshift__n0024_Sh<52>1  (
    .ADR0(DLX_IDinst_reg_out_B_3_1),
    .ADR1(DLX_IDinst_reg_out_B_2_1),
    .ADR2(\DLX_EXinst_Mshift__n0019_Sh[24] ),
    .ADR3(DLX_EXinst_N72809),
    .O(\DLX_EXinst_N72809/GROM )
  );
  X_BUF \DLX_EXinst_N72809/XUSED  (
    .I(\DLX_EXinst_N72809/FROM ),
    .O(DLX_EXinst_N72809)
  );
  X_BUF \DLX_EXinst_N72809/YUSED  (
    .I(\DLX_EXinst_N72809/GROM ),
    .O(\DLX_EXinst_Mshift__n0024_Sh[52] )
  );
  defparam DLX_IDinst_RegFile_28_12_1480.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_28_12_1480 (
    .I(DLX_IDinst_WB_data_eff[12]),
    .CE(DLX_IDinst__n0606),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_28_12)
  );
  defparam DLX_EXinst_Ker735271.INIT = 16'hF0AA;
  X_LUT4 DLX_EXinst_Ker735271 (
    .ADR0(DLX_IDinst_reg_out_A[16]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[18]),
    .ADR3(DLX_IDinst_Imm_1_1),
    .O(\DLX_EXinst_N73529/FROM )
  );
  defparam DLX_EXinst_Ker75137_SW0.INIT = 16'hFC30;
  X_LUT4 DLX_EXinst_Ker75137_SW0 (
    .ADR0(VCC),
    .ADR1(\DLX_IDinst_Imm[0] ),
    .ADR2(DLX_EXinst_N73133),
    .ADR3(DLX_EXinst_N73529),
    .O(\DLX_EXinst_N73529/GROM )
  );
  X_BUF \DLX_EXinst_N73529/XUSED  (
    .I(\DLX_EXinst_N73529/FROM ),
    .O(DLX_EXinst_N73529)
  );
  X_BUF \DLX_EXinst_N73529/YUSED  (
    .I(\DLX_EXinst_N73529/GROM ),
    .O(N130875)
  );
  defparam DLX_EXinst_Ker733671.INIT = 16'hACAC;
  X_LUT4 DLX_EXinst_Ker733671 (
    .ADR0(\DLX_EXinst_Mshift__n0019_Sh[28] ),
    .ADR1(\DLX_EXinst_Mshift__n0019_Sh[24] ),
    .ADR2(DLX_IDinst_reg_out_B[2]),
    .ADR3(VCC),
    .O(\DLX_EXinst_N73369/FROM )
  );
  defparam \DLX_EXinst__n0007<24>175 .INIT = 16'h1000;
  X_LUT4 \DLX_EXinst__n0007<24>175  (
    .ADR0(DLX_IDinst_reg_out_B[3]),
    .ADR1(DLX_IDinst_reg_out_B[4]),
    .ADR2(DLX_EXinst__n0081),
    .ADR3(DLX_EXinst_N73369),
    .O(\DLX_EXinst_N73369/GROM )
  );
  X_BUF \DLX_EXinst_N73369/XUSED  (
    .I(\DLX_EXinst_N73369/FROM ),
    .O(DLX_EXinst_N73369)
  );
  X_BUF \DLX_EXinst_N73369/YUSED  (
    .I(\DLX_EXinst_N73369/GROM ),
    .O(CHOICE5628)
  );
  defparam DLX_EXinst_Ker734721.INIT = 16'hFA50;
  X_LUT4 DLX_EXinst_Ker734721 (
    .ADR0(\DLX_IDinst_Imm[1] ),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[14]),
    .ADR3(DLX_IDinst_reg_out_A[12]),
    .O(\DLX_EXinst_N73474/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0021_Sh<15>1 .INIT = 16'hEE22;
  X_LUT4 \DLX_EXinst_Mshift__n0021_Sh<15>1  (
    .ADR0(DLX_EXinst_N72953),
    .ADR1(DLX_IDinst_Imm_0_1),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N73474),
    .O(\DLX_EXinst_N73474/GROM )
  );
  X_BUF \DLX_EXinst_N73474/XUSED  (
    .I(\DLX_EXinst_N73474/FROM ),
    .O(DLX_EXinst_N73474)
  );
  X_BUF \DLX_EXinst_N73474/YUSED  (
    .I(\DLX_EXinst_N73474/GROM ),
    .O(\DLX_EXinst_Mshift__n0021_Sh[15] )
  );
  defparam DLX_EXinst_Ker733921.INIT = 16'hF5A0;
  X_LUT4 DLX_EXinst_Ker733921 (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[16]),
    .ADR3(DLX_IDinst_reg_out_A[14]),
    .O(\DLX_EXinst_N73394/FROM )
  );
  defparam DLX_EXinst_Ker74449_SW0.INIT = 16'hEE44;
  X_LUT4 DLX_EXinst_Ker74449_SW0 (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(DLX_EXinst_N73043),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N73394),
    .O(\DLX_EXinst_N73394/GROM )
  );
  X_BUF \DLX_EXinst_N73394/XUSED  (
    .I(\DLX_EXinst_N73394/FROM ),
    .O(DLX_EXinst_N73394)
  );
  X_BUF \DLX_EXinst_N73394/YUSED  (
    .I(\DLX_EXinst_N73394/GROM ),
    .O(N130519)
  );
  defparam DLX_EXinst_Ker727441.INIT = 16'hFBFF;
  X_LUT4 DLX_EXinst_Ker727441 (
    .ADR0(DLX_IDinst_reg_dst),
    .ADR1(DLX_EXinst_N76047),
    .ADR2(DLX_IDinst_IR_opcode_field[2]),
    .ADR3(DLX_IDinst_IR_opcode_field[3]),
    .O(\DLX_EXinst_reg_out_B_EX<0>/FROM )
  );
  defparam \DLX_EXinst__n0008<31>1 .INIT = 16'hF000;
  X_LUT4 \DLX_EXinst__n0008<31>1  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[31]),
    .ADR3(DLX_EXinst_N72746),
    .O(DLX_EXinst__n0008[31])
  );
  X_BUF \DLX_EXinst_reg_out_B_EX<0>/XUSED  (
    .I(\DLX_EXinst_reg_out_B_EX<0>/FROM ),
    .O(DLX_EXinst_N72746)
  );
  defparam DLX_EXinst_Ker735371.INIT = 16'hDD88;
  X_LUT4 DLX_EXinst_Ker735371 (
    .ADR0(DLX_IDinst_Imm_1_1),
    .ADR1(DLX_IDinst_reg_out_A[22]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[20]),
    .O(\DLX_EXinst_N73539/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0022_Sh<19>1 .INIT = 16'hFA50;
  X_LUT4 \DLX_EXinst_Mshift__n0022_Sh<19>1  (
    .ADR0(DLX_IDinst_Imm_0_1),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N73143),
    .ADR3(DLX_EXinst_N73539),
    .O(\DLX_EXinst_N73539/GROM )
  );
  X_BUF \DLX_EXinst_N73539/XUSED  (
    .I(\DLX_EXinst_N73539/FROM ),
    .O(DLX_EXinst_N73539)
  );
  X_BUF \DLX_EXinst_N73539/YUSED  (
    .I(\DLX_EXinst_N73539/GROM ),
    .O(\DLX_EXinst_Mshift__n0022_Sh[19] )
  );
  defparam DLX_EXinst_Ker760091.INIT = 16'h0200;
  X_LUT4 DLX_EXinst_Ker760091 (
    .ADR0(DLX_IDinst_IR_opcode_field[3]),
    .ADR1(DLX_IDinst_IR_opcode_field[5]),
    .ADR2(DLX_IDinst_IR_opcode_field[4]),
    .ADR3(DLX_IDinst_IR_opcode_field[2]),
    .O(\DLX_EXinst_N76011/FROM )
  );
  defparam DLX_EXinst__n00531.INIT = 16'h0A00;
  X_LUT4 DLX_EXinst__n00531 (
    .ADR0(DLX_IDinst_IR_opcode_field[0]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_IR_opcode_field[1]),
    .ADR3(DLX_EXinst_N76011),
    .O(\DLX_EXinst_N76011/GROM )
  );
  X_BUF \DLX_EXinst_N76011/XUSED  (
    .I(\DLX_EXinst_N76011/FROM ),
    .O(DLX_EXinst_N76011)
  );
  X_BUF \DLX_EXinst_N76011/YUSED  (
    .I(\DLX_EXinst_N76011/GROM ),
    .O(DLX_EXinst__n0053)
  );
  defparam DLX_EXinst_Ker733771.INIT = 16'hFC30;
  X_LUT4 DLX_EXinst_Ker733771 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_Imm_2_1),
    .ADR2(\DLX_EXinst_Mshift__n0022_Sh[24] ),
    .ADR3(\DLX_EXinst_Mshift__n0020_Sh[28] ),
    .O(\DLX_EXinst_N73379/GROM )
  );
  X_BUF \DLX_EXinst_N73379/YUSED  (
    .I(\DLX_EXinst_N73379/GROM ),
    .O(DLX_EXinst_N73379)
  );
  defparam DLX_EXinst_Ker735621.INIT = 16'hCFC0;
  X_LUT4 DLX_EXinst_Ker735621 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[10]),
    .ADR2(DLX_IDinst_reg_out_B[1]),
    .ADR3(DLX_IDinst_reg_out_A[12]),
    .O(\DLX_EXinst_N73564/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<13>1 .INIT = 16'hFA0A;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<13>1  (
    .ADR0(DLX_EXinst_N72863),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[0]),
    .ADR3(DLX_EXinst_N73564),
    .O(\DLX_EXinst_N73564/GROM )
  );
  X_BUF \DLX_EXinst_N73564/XUSED  (
    .I(\DLX_EXinst_N73564/FROM ),
    .O(DLX_EXinst_N73564)
  );
  X_BUF \DLX_EXinst_N73564/YUSED  (
    .I(\DLX_EXinst_N73564/GROM ),
    .O(\DLX_EXinst_Mshift__n0023_Sh[13] )
  );
  defparam DLX_EXinst_Ker741941.INIT = 16'hF3C0;
  X_LUT4 DLX_EXinst_Ker741941 (
    .ADR0(VCC),
    .ADR1(\DLX_IDinst_Imm[3] ),
    .ADR2(\DLX_EXinst_Mshift__n0021_Sh[13] ),
    .ADR3(\DLX_EXinst_Mshift__n0021_Sh[21] ),
    .O(\DLX_EXinst_N74196/FROM )
  );
  defparam \DLX_EXinst__n0007<25>53 .INIT = 16'hC808;
  X_LUT4 \DLX_EXinst__n0007<25>53  (
    .ADR0(N133768),
    .ADR1(DLX_EXinst__n0055),
    .ADR2(\DLX_IDinst_Imm[2] ),
    .ADR3(DLX_EXinst_N74196),
    .O(\DLX_EXinst_N74196/GROM )
  );
  X_BUF \DLX_EXinst_N74196/XUSED  (
    .I(\DLX_EXinst_N74196/FROM ),
    .O(DLX_EXinst_N74196)
  );
  X_BUF \DLX_EXinst_N74196/YUSED  (
    .I(\DLX_EXinst_N74196/GROM ),
    .O(CHOICE5076)
  );
  defparam DLX_EXinst_Ker735771.INIT = 16'hF3C0;
  X_LUT4 DLX_EXinst_Ker735771 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(DLX_IDinst_reg_out_A[16]),
    .ADR3(DLX_IDinst_reg_out_A[18]),
    .O(\DLX_EXinst_N73579/FROM )
  );
  defparam DLX_EXinst_Ker734821.INIT = 16'hF0AA;
  X_LUT4 DLX_EXinst_Ker734821 (
    .ADR0(DLX_IDinst_reg_out_A[18]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[16]),
    .ADR3(\DLX_IDinst_Imm[1] ),
    .O(\DLX_EXinst_N73579/GROM )
  );
  X_BUF \DLX_EXinst_N73579/XUSED  (
    .I(\DLX_EXinst_N73579/FROM ),
    .O(DLX_EXinst_N73579)
  );
  X_BUF \DLX_EXinst_N73579/YUSED  (
    .I(\DLX_EXinst_N73579/GROM ),
    .O(DLX_EXinst_N73484)
  );
  defparam DLX_EXinst_Ker728511.INIT = 16'hAACC;
  X_LUT4 DLX_EXinst_Ker728511 (
    .ADR0(DLX_IDinst_reg_out_A[7]),
    .ADR1(DLX_IDinst_reg_out_A[9]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[1]),
    .O(\DLX_EXinst_N72853/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<10>1 .INIT = 16'hFC30;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<10>1  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_B[0]),
    .ADR2(DLX_EXinst_N73559),
    .ADR3(DLX_EXinst_N72853),
    .O(\DLX_EXinst_N72853/GROM )
  );
  X_BUF \DLX_EXinst_N72853/XUSED  (
    .I(\DLX_EXinst_N72853/FROM ),
    .O(DLX_EXinst_N72853)
  );
  X_BUF \DLX_EXinst_N72853/YUSED  (
    .I(\DLX_EXinst_N72853/GROM ),
    .O(\DLX_EXinst_Mshift__n0023_Sh[10] )
  );
  defparam DLX_EXinst_Ker733871.INIT = 16'hAFA0;
  X_LUT4 DLX_EXinst_Ker733871 (
    .ADR0(DLX_IDinst_reg_out_A[14]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[1]),
    .ADR3(DLX_IDinst_reg_out_A[12]),
    .O(\DLX_EXinst_N73389/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0019_Sh<11>1 .INIT = 16'hFC30;
  X_LUT4 \DLX_EXinst_Mshift__n0019_Sh<11>1  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_B[0]),
    .ADR2(DLX_EXinst_N73038),
    .ADR3(DLX_EXinst_N73389),
    .O(\DLX_EXinst_N73389/GROM )
  );
  X_BUF \DLX_EXinst_N73389/XUSED  (
    .I(\DLX_EXinst_N73389/FROM ),
    .O(DLX_EXinst_N73389)
  );
  X_BUF \DLX_EXinst_N73389/YUSED  (
    .I(\DLX_EXinst_N73389/GROM ),
    .O(\DLX_EXinst_Mshift__n0019_Sh[11] )
  );
  defparam DLX_EXinst_Ker734671.INIT = 16'hCACA;
  X_LUT4 DLX_EXinst_Ker734671 (
    .ADR0(DLX_IDinst_reg_out_A[12]),
    .ADR1(DLX_IDinst_reg_out_A[10]),
    .ADR2(\DLX_IDinst_Imm[1] ),
    .ADR3(VCC),
    .O(\DLX_EXinst_N73469/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0021_Sh<13>1 .INIT = 16'hEE44;
  X_LUT4 \DLX_EXinst_Mshift__n0021_Sh<13>1  (
    .ADR0(DLX_IDinst_Imm_0_1),
    .ADR1(DLX_EXinst_N72948),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N73469),
    .O(\DLX_EXinst_N73469/GROM )
  );
  X_BUF \DLX_EXinst_N73469/XUSED  (
    .I(\DLX_EXinst_N73469/FROM ),
    .O(DLX_EXinst_N73469)
  );
  X_BUF \DLX_EXinst_N73469/YUSED  (
    .I(\DLX_EXinst_N73469/GROM ),
    .O(\DLX_EXinst_Mshift__n0021_Sh[13] )
  );
  defparam DLX_EXinst_Ker734921.INIT = 16'hAFA0;
  X_LUT4 DLX_EXinst_Ker734921 (
    .ADR0(DLX_IDinst_reg_out_A[20]),
    .ADR1(VCC),
    .ADR2(\DLX_IDinst_Imm[1] ),
    .ADR3(DLX_IDinst_reg_out_A[22]),
    .O(\DLX_EXinst_N73494/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0021_Sh<23>1 .INIT = 16'hFC0C;
  X_LUT4 \DLX_EXinst_Mshift__n0021_Sh<23>1  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N72973),
    .ADR2(DLX_IDinst_Imm_0_1),
    .ADR3(DLX_EXinst_N73494),
    .O(\DLX_EXinst_N73494/GROM )
  );
  X_BUF \DLX_EXinst_N73494/XUSED  (
    .I(\DLX_EXinst_N73494/FROM ),
    .O(DLX_EXinst_N73494)
  );
  X_BUF \DLX_EXinst_N73494/YUSED  (
    .I(\DLX_EXinst_N73494/GROM ),
    .O(\DLX_EXinst_Mshift__n0021_Sh[23] )
  );
  defparam DLX_EXinst_Ker735721.INIT = 16'hAFA0;
  X_LUT4 DLX_EXinst_Ker735721 (
    .ADR0(DLX_IDinst_reg_out_A[14]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[1]),
    .ADR3(DLX_IDinst_reg_out_A[16]),
    .O(\DLX_EXinst_N73574/FROM )
  );
  defparam DLX_EXinst_Ker73846_SW0.INIT = 16'hFA50;
  X_LUT4 DLX_EXinst_Ker73846_SW0 (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N72873),
    .ADR3(DLX_EXinst_N73574),
    .O(\DLX_EXinst_N73574/GROM )
  );
  X_BUF \DLX_EXinst_N73574/XUSED  (
    .I(\DLX_EXinst_N73574/FROM ),
    .O(DLX_EXinst_N73574)
  );
  X_BUF \DLX_EXinst_N73574/YUSED  (
    .I(\DLX_EXinst_N73574/GROM ),
    .O(N129951)
  );
  defparam DLX_EXinst_Ker74684.INIT = 16'hE2E2;
  X_LUT4 DLX_EXinst_Ker74684 (
    .ADR0(N130621),
    .ADR1(DLX_IDinst_reg_out_B_3_1),
    .ADR2(\DLX_EXinst_Mshift__n0019_Sh[23] ),
    .ADR3(VCC),
    .O(\DLX_EXinst_N74686/FROM )
  );
  defparam DLX_EXinst_Ker744441.INIT = 16'hE2E2;
  X_LUT4 DLX_EXinst_Ker744441 (
    .ADR0(\DLX_EXinst_Mshift__n0019_Sh[12] ),
    .ADR1(DLX_IDinst_reg_out_B_3_1),
    .ADR2(\DLX_EXinst_Mshift__n0019_Sh[20] ),
    .ADR3(VCC),
    .O(\DLX_EXinst_N74686/GROM )
  );
  X_BUF \DLX_EXinst_N74686/XUSED  (
    .I(\DLX_EXinst_N74686/FROM ),
    .O(DLX_EXinst_N74686)
  );
  X_BUF \DLX_EXinst_N74686/YUSED  (
    .I(\DLX_EXinst_N74686/GROM ),
    .O(DLX_EXinst_N74446)
  );
  defparam DLX_EXinst_Ker729411.INIT = 16'hEE22;
  X_LUT4 DLX_EXinst_Ker729411 (
    .ADR0(DLX_IDinst_reg_out_A[11]),
    .ADR1(\DLX_IDinst_Imm[1] ),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[9]),
    .O(\DLX_EXinst_N72943/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0021_Sh<12>1 .INIT = 16'hFA50;
  X_LUT4 \DLX_EXinst_Mshift__n0021_Sh<12>1  (
    .ADR0(DLX_IDinst_Imm_0_1),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N73469),
    .ADR3(DLX_EXinst_N72943),
    .O(\DLX_EXinst_N72943/GROM )
  );
  X_BUF \DLX_EXinst_N72943/XUSED  (
    .I(\DLX_EXinst_N72943/FROM ),
    .O(DLX_EXinst_N72943)
  );
  X_BUF \DLX_EXinst_N72943/YUSED  (
    .I(\DLX_EXinst_N72943/GROM ),
    .O(\DLX_EXinst_Mshift__n0021_Sh[12] )
  );
  defparam DLX_IDinst_RegFile_28_13_1481.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_28_13_1481 (
    .I(DLX_IDinst_WB_data_eff[13]),
    .CE(DLX_IDinst__n0606),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_28_13)
  );
  defparam DLX_EXinst_Ker728611.INIT = 16'hAACC;
  X_LUT4 DLX_EXinst_Ker728611 (
    .ADR0(DLX_IDinst_reg_out_A[11]),
    .ADR1(DLX_IDinst_reg_out_A[13]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[1]),
    .O(\DLX_EXinst_N72863/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<14>1 .INIT = 16'hFC0C;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<14>1  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N73569),
    .ADR2(DLX_IDinst_reg_out_B[0]),
    .ADR3(DLX_EXinst_N72863),
    .O(\DLX_EXinst_N72863/GROM )
  );
  X_BUF \DLX_EXinst_N72863/XUSED  (
    .I(\DLX_EXinst_N72863/FROM ),
    .O(DLX_EXinst_N72863)
  );
  X_BUF \DLX_EXinst_N72863/YUSED  (
    .I(\DLX_EXinst_N72863/GROM ),
    .O(\DLX_EXinst_Mshift__n0023_Sh[14] )
  );
  defparam DLX_EXinst_Ker733971.INIT = 16'hD8D8;
  X_LUT4 DLX_EXinst_Ker733971 (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(DLX_IDinst_reg_out_A[18]),
    .ADR2(DLX_IDinst_reg_out_A[16]),
    .ADR3(VCC),
    .O(\DLX_EXinst_N73399/FROM )
  );
  defparam DLX_EXinst_Ker74684_SW0.INIT = 16'hEE44;
  X_LUT4 DLX_EXinst_Ker74684_SW0 (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(DLX_EXinst_N73048),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N73399),
    .O(\DLX_EXinst_N73399/GROM )
  );
  X_BUF \DLX_EXinst_N73399/XUSED  (
    .I(\DLX_EXinst_N73399/FROM ),
    .O(DLX_EXinst_N73399)
  );
  X_BUF \DLX_EXinst_N73399/YUSED  (
    .I(\DLX_EXinst_N73399/GROM ),
    .O(N130621)
  );
  defparam DLX_EXinst_Ker760451.INIT = 16'h0500;
  X_LUT4 DLX_EXinst_Ker760451 (
    .ADR0(DLX_IDinst_IR_opcode_field[4]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_IR_opcode_field[1]),
    .ADR3(DLX_IDinst_IR_opcode_field[5]),
    .O(\DLX_EXinst_word/FROM )
  );
  defparam DLX_EXinst__n00111.INIT = 16'h2A00;
  X_LUT4 DLX_EXinst__n00111 (
    .ADR0(DLX_IDinst_IR_opcode_field[0]),
    .ADR1(DLX_IDinst_IR_opcode_field[3]),
    .ADR2(DLX_IDinst_IR_opcode_field[2]),
    .ADR3(DLX_EXinst_N76047),
    .O(DLX_EXinst__n0011)
  );
  X_BUF \DLX_EXinst_word/XUSED  (
    .I(\DLX_EXinst_word/FROM ),
    .O(DLX_EXinst_N76047)
  );
  defparam DLX_IDinst_RegFile_28_21_1482.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_28_21_1482 (
    .I(DLX_IDinst_WB_data_eff[21]),
    .CE(DLX_IDinst__n0606),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_28_21)
  );
  defparam DLX_EXinst_Ker734771.INIT = 16'hAFA0;
  X_LUT4 DLX_EXinst_Ker734771 (
    .ADR0(DLX_IDinst_reg_out_A[14]),
    .ADR1(VCC),
    .ADR2(\DLX_IDinst_Imm[1] ),
    .ADR3(DLX_IDinst_reg_out_A[16]),
    .O(\DLX_EXinst_N73479/FROM )
  );
  defparam DLX_EXinst_Ker73991_SW0.INIT = 16'hFC30;
  X_LUT4 DLX_EXinst_Ker73991_SW0 (
    .ADR0(VCC),
    .ADR1(\DLX_IDinst_Imm[0] ),
    .ADR2(DLX_EXinst_N72958),
    .ADR3(DLX_EXinst_N73479),
    .O(\DLX_EXinst_N73479/GROM )
  );
  X_BUF \DLX_EXinst_N73479/XUSED  (
    .I(\DLX_EXinst_N73479/FROM ),
    .O(DLX_EXinst_N73479)
  );
  X_BUF \DLX_EXinst_N73479/YUSED  (
    .I(\DLX_EXinst_N73479/GROM ),
    .O(N130209)
  );
  defparam DLX_EXinst_Ker735571.INIT = 16'hAAF0;
  X_LUT4 DLX_EXinst_Ker735571 (
    .ADR0(DLX_IDinst_reg_out_A[8]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[10]),
    .ADR3(DLX_IDinst_reg_out_B[1]),
    .O(\DLX_EXinst_N73559/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<11>1 .INIT = 16'hFA50;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<11>1  (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N72858),
    .ADR3(DLX_EXinst_N73559),
    .O(\DLX_EXinst_N73559/GROM )
  );
  X_BUF \DLX_EXinst_N73559/XUSED  (
    .I(\DLX_EXinst_N73559/FROM ),
    .O(DLX_EXinst_N73559)
  );
  X_BUF \DLX_EXinst_N73559/YUSED  (
    .I(\DLX_EXinst_N73559/GROM ),
    .O(\DLX_EXinst_Mshift__n0023_Sh[11] )
  );
  defparam DLX_EXinst__n00101.INIT = 16'h1030;
  X_LUT4 DLX_EXinst__n00101 (
    .ADR0(DLX_IDinst_IR_opcode_field[3]),
    .ADR1(DLX_IDinst_IR_opcode_field[0]),
    .ADR2(DLX_EXinst_N76047),
    .ADR3(DLX_IDinst_IR_opcode_field[2]),
    .O(DLX_EXinst__n0010)
  );
  defparam DLX_EXinst_Ker763101.INIT = 16'h5500;
  X_LUT4 DLX_EXinst_Ker763101 (
    .ADR0(DLX_IDinst_IR_opcode_field[5]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_IR_opcode_field[3]),
    .O(\DLX_EXinst_byte/GROM )
  );
  X_BUF \DLX_EXinst_byte/YUSED  (
    .I(\DLX_EXinst_byte/GROM ),
    .O(DLX_EXinst_N76312)
  );
  defparam DLX_EXinst_Ker735821.INIT = 16'hE2E2;
  X_LUT4 DLX_EXinst_Ker735821 (
    .ADR0(DLX_IDinst_reg_out_A[20]),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(DLX_IDinst_reg_out_A[18]),
    .ADR3(VCC),
    .O(\DLX_EXinst_N73584/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<21>1 .INIT = 16'hFA0A;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<21>1  (
    .ADR0(DLX_EXinst_N72883),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[0]),
    .ADR3(DLX_EXinst_N73584),
    .O(\DLX_EXinst_N73584/GROM )
  );
  X_BUF \DLX_EXinst_N73584/XUSED  (
    .I(\DLX_EXinst_N73584/FROM ),
    .O(DLX_EXinst_N73584)
  );
  X_BUF \DLX_EXinst_N73584/YUSED  (
    .I(\DLX_EXinst_N73584/GROM ),
    .O(\DLX_EXinst_Mshift__n0023_Sh[21] )
  );
  defparam DLX_EXinst_Ker728711.INIT = 16'hCFC0;
  X_LUT4 DLX_EXinst_Ker728711 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[15]),
    .ADR2(DLX_IDinst_reg_out_B[1]),
    .ADR3(DLX_IDinst_reg_out_A[17]),
    .O(\DLX_EXinst_N72873/FROM )
  );
  defparam DLX_EXinst_Ker73851_SW0.INIT = 16'hEE22;
  X_LUT4 DLX_EXinst_Ker73851_SW0 (
    .ADR0(DLX_EXinst_N73579),
    .ADR1(DLX_IDinst_reg_out_B[0]),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N72873),
    .O(\DLX_EXinst_N72873/GROM )
  );
  X_BUF \DLX_EXinst_N72873/XUSED  (
    .I(\DLX_EXinst_N72873/FROM ),
    .O(DLX_EXinst_N72873)
  );
  X_BUF \DLX_EXinst_N72873/YUSED  (
    .I(\DLX_EXinst_N72873/GROM ),
    .O(N130001)
  );
  defparam DLX_EXinst_Ker735671.INIT = 16'hFA50;
  X_LUT4 DLX_EXinst_Ker735671 (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[14]),
    .ADR3(DLX_IDinst_reg_out_A[12]),
    .O(\DLX_EXinst_N73569/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<15>1 .INIT = 16'hEE22;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<15>1  (
    .ADR0(DLX_EXinst_N72868),
    .ADR1(DLX_IDinst_reg_out_B[0]),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N73569),
    .O(\DLX_EXinst_N73569/GROM )
  );
  X_BUF \DLX_EXinst_N73569/XUSED  (
    .I(\DLX_EXinst_N73569/FROM ),
    .O(DLX_EXinst_N73569)
  );
  X_BUF \DLX_EXinst_N73569/YUSED  (
    .I(\DLX_EXinst_N73569/GROM ),
    .O(\DLX_EXinst_Mshift__n0023_Sh[15] )
  );
  defparam DLX_EXinst_Ker734871.INIT = 16'hAACC;
  X_LUT4 DLX_EXinst_Ker734871 (
    .ADR0(DLX_IDinst_reg_out_A[18]),
    .ADR1(DLX_IDinst_reg_out_A[20]),
    .ADR2(VCC),
    .ADR3(\DLX_IDinst_Imm[1] ),
    .O(\DLX_EXinst_N73489/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0021_Sh<21>1 .INIT = 16'hFA0A;
  X_LUT4 \DLX_EXinst_Mshift__n0021_Sh<21>1  (
    .ADR0(DLX_EXinst_N72968),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_Imm_0_1),
    .ADR3(DLX_EXinst_N73489),
    .O(\DLX_EXinst_N73489/GROM )
  );
  X_BUF \DLX_EXinst_N73489/XUSED  (
    .I(\DLX_EXinst_N73489/FROM ),
    .O(DLX_EXinst_N73489)
  );
  X_BUF \DLX_EXinst_N73489/YUSED  (
    .I(\DLX_EXinst_N73489/GROM ),
    .O(\DLX_EXinst_Mshift__n0021_Sh[21] )
  );
  defparam DLX_EXinst_Ker741991.INIT = 16'hFC0C;
  X_LUT4 DLX_EXinst_Ker741991 (
    .ADR0(VCC),
    .ADR1(\DLX_EXinst_Mshift__n0021_Sh[22] ),
    .ADR2(\DLX_IDinst_Imm[3] ),
    .ADR3(\DLX_EXinst_Mshift__n0021_Sh[14] ),
    .O(\DLX_EXinst_N74201/FROM )
  );
  defparam \DLX_EXinst__n0007<26>53 .INIT = 16'hE040;
  X_LUT4 \DLX_EXinst__n0007<26>53  (
    .ADR0(\DLX_IDinst_Imm[2] ),
    .ADR1(N134128),
    .ADR2(DLX_EXinst__n0055),
    .ADR3(DLX_EXinst_N74201),
    .O(\DLX_EXinst_N74201/GROM )
  );
  X_BUF \DLX_EXinst_N74201/XUSED  (
    .I(\DLX_EXinst_N74201/FROM ),
    .O(DLX_EXinst_N74201)
  );
  X_BUF \DLX_EXinst_N74201/YUSED  (
    .I(\DLX_EXinst_N74201/GROM ),
    .O(CHOICE5009)
  );
  defparam DLX_EXinst_Ker760391.INIT = 16'h0008;
  X_LUT4 DLX_EXinst_Ker760391 (
    .ADR0(DLX_IDinst_IR_opcode_field[2]),
    .ADR1(DLX_IDinst_IR_opcode_field[4]),
    .ADR2(DLX_IDinst_IR_opcode_field[3]),
    .ADR3(DLX_IDinst_IR_opcode_field[5]),
    .O(\DLX_EXinst_N76041/FROM )
  );
  defparam DLX_EXinst__n00551.INIT = 16'h1100;
  X_LUT4 DLX_EXinst__n00551 (
    .ADR0(DLX_IDinst_IR_opcode_field[0]),
    .ADR1(DLX_IDinst_IR_opcode_field[1]),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N76041),
    .O(\DLX_EXinst_N76041/GROM )
  );
  X_BUF \DLX_EXinst_N76041/XUSED  (
    .I(\DLX_EXinst_N76041/FROM ),
    .O(DLX_EXinst_N76041)
  );
  X_BUF \DLX_EXinst_N76041/YUSED  (
    .I(\DLX_EXinst_N76041/GROM ),
    .O(DLX_EXinst__n0055)
  );
  defparam DLX_EXinst_Ker728561.INIT = 16'hACAC;
  X_LUT4 DLX_EXinst_Ker728561 (
    .ADR0(DLX_IDinst_reg_out_A[9]),
    .ADR1(DLX_IDinst_reg_out_A[11]),
    .ADR2(DLX_IDinst_reg_out_B[1]),
    .ADR3(VCC),
    .O(\DLX_EXinst_N72858/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<12>1 .INIT = 16'hEE22;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<12>1  (
    .ADR0(DLX_EXinst_N73564),
    .ADR1(DLX_IDinst_reg_out_B[0]),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N72858),
    .O(\DLX_EXinst_N72858/GROM )
  );
  X_BUF \DLX_EXinst_N72858/XUSED  (
    .I(\DLX_EXinst_N72858/FROM ),
    .O(DLX_EXinst_N72858)
  );
  X_BUF \DLX_EXinst_N72858/YUSED  (
    .I(\DLX_EXinst_N72858/GROM ),
    .O(\DLX_EXinst_Mshift__n0023_Sh[12] )
  );
  defparam DLX_EXinst_Ker75137.INIT = 16'hFC30;
  X_LUT4 DLX_EXinst_Ker75137 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_Imm_3_1),
    .ADR2(N130875),
    .ADR3(\DLX_EXinst_Mshift__n0022_Sh[23] ),
    .O(\DLX_EXinst_N75139/FROM )
  );
  defparam DLX_EXinst_Ker747041.INIT = 16'hEE44;
  X_LUT4 DLX_EXinst_Ker747041 (
    .ADR0(DLX_IDinst_Imm_3_1),
    .ADR1(\DLX_EXinst_Mshift__n0022_Sh[12] ),
    .ADR2(VCC),
    .ADR3(\DLX_EXinst_Mshift__n0022_Sh[20] ),
    .O(\DLX_EXinst_N75139/GROM )
  );
  X_BUF \DLX_EXinst_N75139/XUSED  (
    .I(\DLX_EXinst_N75139/FROM ),
    .O(DLX_EXinst_N75139)
  );
  X_BUF \DLX_EXinst_N75139/YUSED  (
    .I(\DLX_EXinst_N75139/GROM ),
    .O(DLX_EXinst_N74706)
  );
  defparam DLX_EXinst_Ker729611.INIT = 16'hFA0A;
  X_LUT4 DLX_EXinst_Ker729611 (
    .ADR0(DLX_IDinst_reg_out_A[19]),
    .ADR1(VCC),
    .ADR2(\DLX_IDinst_Imm[1] ),
    .ADR3(DLX_IDinst_reg_out_A[17]),
    .O(\DLX_EXinst_N72963/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0021_Sh<20>1 .INIT = 16'hFA0A;
  X_LUT4 \DLX_EXinst_Mshift__n0021_Sh<20>1  (
    .ADR0(DLX_EXinst_N73489),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_Imm_0_1),
    .ADR3(DLX_EXinst_N72963),
    .O(\DLX_EXinst_N72963/GROM )
  );
  X_BUF \DLX_EXinst_N72963/XUSED  (
    .I(\DLX_EXinst_N72963/FROM ),
    .O(DLX_EXinst_N72963)
  );
  X_BUF \DLX_EXinst_N72963/YUSED  (
    .I(\DLX_EXinst_N72963/GROM ),
    .O(\DLX_EXinst_Mshift__n0021_Sh[20] )
  );
  defparam DLX_EXinst_Ker728811.INIT = 16'hFA50;
  X_LUT4 DLX_EXinst_Ker728811 (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[21]),
    .ADR3(DLX_IDinst_reg_out_A[19]),
    .O(\DLX_EXinst_N72883/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<22>1 .INIT = 16'hFA50;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<22>1  (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N73589),
    .ADR3(DLX_EXinst_N72883),
    .O(\DLX_EXinst_N72883/GROM )
  );
  X_BUF \DLX_EXinst_N72883/XUSED  (
    .I(\DLX_EXinst_N72883/FROM ),
    .O(DLX_EXinst_N72883)
  );
  X_BUF \DLX_EXinst_N72883/YUSED  (
    .I(\DLX_EXinst_N72883/GROM ),
    .O(\DLX_EXinst_Mshift__n0023_Sh[22] )
  );
  defparam DLX_EXinst_Ker729461.INIT = 16'hACAC;
  X_LUT4 DLX_EXinst_Ker729461 (
    .ADR0(DLX_IDinst_reg_out_A[11]),
    .ADR1(DLX_IDinst_reg_out_A[13]),
    .ADR2(\DLX_IDinst_Imm[1] ),
    .ADR3(VCC),
    .O(\DLX_EXinst_N72948/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0021_Sh<14>1 .INIT = 16'hFA50;
  X_LUT4 \DLX_EXinst_Mshift__n0021_Sh<14>1  (
    .ADR0(DLX_IDinst_Imm_0_1),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N73474),
    .ADR3(DLX_EXinst_N72948),
    .O(\DLX_EXinst_N72948/GROM )
  );
  X_BUF \DLX_EXinst_N72948/XUSED  (
    .I(\DLX_EXinst_N72948/FROM ),
    .O(DLX_EXinst_N72948)
  );
  X_BUF \DLX_EXinst_N72948/YUSED  (
    .I(\DLX_EXinst_N72948/GROM ),
    .O(\DLX_EXinst_Mshift__n0021_Sh[14] )
  );
  defparam DLX_EXinst_Ker728861.INIT = 16'hB8B8;
  X_LUT4 DLX_EXinst_Ker728861 (
    .ADR0(DLX_IDinst_reg_out_A[21]),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(DLX_IDinst_reg_out_A[23]),
    .ADR3(VCC),
    .O(\DLX_EXinst_N72888/FROM )
  );
  defparam DLX_EXinst_Ker728911.INIT = 16'hF3C0;
  X_LUT4 DLX_EXinst_Ker728911 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(DLX_IDinst_reg_out_A[23]),
    .ADR3(DLX_IDinst_reg_out_A[25]),
    .O(\DLX_EXinst_N72888/GROM )
  );
  X_BUF \DLX_EXinst_N72888/XUSED  (
    .I(\DLX_EXinst_N72888/FROM ),
    .O(DLX_EXinst_N72888)
  );
  X_BUF \DLX_EXinst_N72888/YUSED  (
    .I(\DLX_EXinst_N72888/GROM ),
    .O(DLX_EXinst_N72893)
  );
  defparam DLX_EXinst_Ker727951.INIT = 16'hEE22;
  X_LUT4 DLX_EXinst_Ker727951 (
    .ADR0(\DLX_EXinst_Mshift__n0022_Sh[20] ),
    .ADR1(\DLX_IDinst_Imm[3] ),
    .ADR2(VCC),
    .ADR3(\DLX_EXinst_Mshift__n0020_Sh[28] ),
    .O(\DLX_EXinst_N72797/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0022_Sh<52>1 .INIT = 16'h5D08;
  X_LUT4 \DLX_EXinst_Mshift__n0022_Sh<52>1  (
    .ADR0(DLX_IDinst_Imm_2_1),
    .ADR1(\DLX_EXinst_Mshift__n0022_Sh[24] ),
    .ADR2(DLX_IDinst_Imm_3_1),
    .ADR3(DLX_EXinst_N72797),
    .O(\DLX_EXinst_N72797/GROM )
  );
  X_BUF \DLX_EXinst_N72797/XUSED  (
    .I(\DLX_EXinst_N72797/FROM ),
    .O(DLX_EXinst_N72797)
  );
  X_BUF \DLX_EXinst_N72797/YUSED  (
    .I(\DLX_EXinst_N72797/GROM ),
    .O(\DLX_EXinst_Mshift__n0022_Sh[52] )
  );
  defparam DLX_EXinst_Ker735871.INIT = 16'hDD88;
  X_LUT4 DLX_EXinst_Ker735871 (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(DLX_IDinst_reg_out_A[20]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[22]),
    .O(\DLX_EXinst_N73589/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<23>1 .INIT = 16'hFC0C;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<23>1  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N72888),
    .ADR2(DLX_IDinst_reg_out_B[0]),
    .ADR3(DLX_EXinst_N73589),
    .O(\DLX_EXinst_N73589/GROM )
  );
  X_BUF \DLX_EXinst_N73589/XUSED  (
    .I(\DLX_EXinst_N73589/FROM ),
    .O(DLX_EXinst_N73589)
  );
  X_BUF \DLX_EXinst_N73589/YUSED  (
    .I(\DLX_EXinst_N73589/GROM ),
    .O(\DLX_EXinst_Mshift__n0023_Sh[23] )
  );
  defparam DLX_EXinst_Ker763161.INIT = 16'h0100;
  X_LUT4 DLX_EXinst_Ker763161 (
    .ADR0(DLX_IDinst_IR_opcode_field[0]),
    .ADR1(DLX_IDinst_IR_opcode_field[1]),
    .ADR2(N146478),
    .ADR3(DLX_EXinst_N76041),
    .O(\DLX_EXinst_N76318/FROM )
  );
  defparam \DLX_EXinst__n0007<15>165 .INIT = 16'hB800;
  X_LUT4 \DLX_EXinst__n0007<15>165  (
    .ADR0(DLX_EXinst_N72998),
    .ADR1(\DLX_IDinst_Imm[3] ),
    .ADR2(N130415),
    .ADR3(DLX_EXinst_N76318),
    .O(\DLX_EXinst_N76318/GROM )
  );
  X_BUF \DLX_EXinst_N76318/XUSED  (
    .I(\DLX_EXinst_N76318/FROM ),
    .O(DLX_EXinst_N76318)
  );
  X_BUF \DLX_EXinst_N76318/YUSED  (
    .I(\DLX_EXinst_N76318/GROM ),
    .O(CHOICE4302)
  );
  defparam DLX_EXinst_Ker729561.INIT = 16'hACAC;
  X_LUT4 DLX_EXinst_Ker729561 (
    .ADR0(DLX_IDinst_reg_out_A[15]),
    .ADR1(DLX_IDinst_reg_out_A[17]),
    .ADR2(\DLX_IDinst_Imm[1] ),
    .ADR3(VCC),
    .O(\DLX_EXinst_N72958/FROM )
  );
  defparam DLX_EXinst_Ker73996_SW0.INIT = 16'hEE22;
  X_LUT4 DLX_EXinst_Ker73996_SW0 (
    .ADR0(DLX_EXinst_N73484),
    .ADR1(\DLX_IDinst_Imm[0] ),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N72958),
    .O(\DLX_EXinst_N72958/GROM )
  );
  X_BUF \DLX_EXinst_N72958/XUSED  (
    .I(\DLX_EXinst_N72958/FROM ),
    .O(DLX_EXinst_N72958)
  );
  X_BUF \DLX_EXinst_N72958/YUSED  (
    .I(\DLX_EXinst_N72958/GROM ),
    .O(N130261)
  );
  defparam DLX_EXinst_Ker728761.INIT = 16'hE2E2;
  X_LUT4 DLX_EXinst_Ker728761 (
    .ADR0(DLX_IDinst_reg_out_A[19]),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(DLX_IDinst_reg_out_A[17]),
    .ADR3(VCC),
    .O(\DLX_EXinst_N72878/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<20>1 .INIT = 16'hFC0C;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<20>1  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N73584),
    .ADR2(DLX_IDinst_reg_out_B[0]),
    .ADR3(DLX_EXinst_N72878),
    .O(\DLX_EXinst_N72878/GROM )
  );
  X_BUF \DLX_EXinst_N72878/XUSED  (
    .I(\DLX_EXinst_N72878/FROM ),
    .O(DLX_EXinst_N72878)
  );
  X_BUF \DLX_EXinst_N72878/YUSED  (
    .I(\DLX_EXinst_N72878/GROM ),
    .O(\DLX_EXinst_Mshift__n0023_Sh[20] )
  );
  defparam DLX_EXinst_Ker727891.INIT = 16'hEE44;
  X_LUT4 DLX_EXinst_Ker727891 (
    .ADR0(\DLX_IDinst_Imm[0] ),
    .ADR1(DLX_IDinst_reg_out_A[29]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[30]),
    .O(\DLX_EXinst_N72791/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0022_Sh<29>1 .INIT = 16'h7520;
  X_LUT4 \DLX_EXinst_Mshift__n0022_Sh<29>1  (
    .ADR0(DLX_IDinst_Imm_1_1),
    .ADR1(DLX_IDinst_Imm_0_1),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(DLX_EXinst_N72791),
    .O(\DLX_EXinst_N72791/GROM )
  );
  X_BUF \DLX_EXinst_N72791/XUSED  (
    .I(\DLX_EXinst_N72791/FROM ),
    .O(DLX_EXinst_N72791)
  );
  X_BUF \DLX_EXinst_N72791/YUSED  (
    .I(\DLX_EXinst_N72791/GROM ),
    .O(\DLX_EXinst_Mshift__n0022_Sh[29] )
  );
  defparam DLX_EXinst_Ker729661.INIT = 16'hCCAA;
  X_LUT4 DLX_EXinst_Ker729661 (
    .ADR0(DLX_IDinst_reg_out_A[21]),
    .ADR1(DLX_IDinst_reg_out_A[19]),
    .ADR2(VCC),
    .ADR3(\DLX_IDinst_Imm[1] ),
    .O(\DLX_EXinst_N72968/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0021_Sh<22>1 .INIT = 16'hEE22;
  X_LUT4 \DLX_EXinst_Mshift__n0021_Sh<22>1  (
    .ADR0(DLX_EXinst_N73494),
    .ADR1(DLX_IDinst_Imm_0_1),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N72968),
    .O(\DLX_EXinst_N72968/GROM )
  );
  X_BUF \DLX_EXinst_N72968/XUSED  (
    .I(\DLX_EXinst_N72968/FROM ),
    .O(DLX_EXinst_N72968)
  );
  X_BUF \DLX_EXinst_N72968/YUSED  (
    .I(\DLX_EXinst_N72968/GROM ),
    .O(\DLX_EXinst_Mshift__n0021_Sh[22] )
  );
  defparam DLX_IDinst_Ker10720623.INIT = 16'h01FF;
  X_LUT4 DLX_IDinst_Ker10720623 (
    .ADR0(DLX_IDinst__n0313),
    .ADR1(DLX_IDinst_N108221),
    .ADR2(DLX_IDinst__n0311),
    .ADR3(DLX_IDinst_N108443),
    .O(\CHOICE2103/GROM )
  );
  X_BUF \CHOICE2103/YUSED  (
    .I(\CHOICE2103/GROM ),
    .O(CHOICE2103)
  );
  defparam DLX_EXinst_Ker749891.INIT = 16'hF3C0;
  X_LUT4 DLX_EXinst_Ker749891 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_B_3_1),
    .ADR2(\DLX_EXinst_Mshift__n0019_Sh[19] ),
    .ADR3(\DLX_EXinst_Mshift__n0019_Sh[11] ),
    .O(\DLX_EXinst_N74991/FROM )
  );
  defparam DLX_EXinst_Ker747191.INIT = 16'hCCAA;
  X_LUT4 DLX_EXinst_Ker747191 (
    .ADR0(\DLX_EXinst_Mshift__n0019_Sh[16] ),
    .ADR1(\DLX_EXinst_Mshift__n0019_Sh[24] ),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B_3_1),
    .O(\DLX_EXinst_N74991/GROM )
  );
  X_BUF \DLX_EXinst_N74991/XUSED  (
    .I(\DLX_EXinst_N74991/FROM ),
    .O(DLX_EXinst_N74991)
  );
  X_BUF \DLX_EXinst_N74991/YUSED  (
    .I(\DLX_EXinst_N74991/GROM ),
    .O(DLX_EXinst_N74721)
  );
  defparam DLX_EXinst_Ker763361.INIT = 16'h0004;
  X_LUT4 DLX_EXinst_Ker763361 (
    .ADR0(CHOICE3576),
    .ADR1(DLX_EXinst__n0080),
    .ADR2(CHOICE3570),
    .ADR3(CHOICE3592),
    .O(\DLX_EXinst_N76338/FROM )
  );
  defparam \DLX_EXinst__n0007<12>34 .INIT = 16'hCA00;
  X_LUT4 \DLX_EXinst__n0007<12>34  (
    .ADR0(DLX_EXinst_N74051),
    .ADR1(DLX_EXinst_N72898),
    .ADR2(DLX_IDinst_reg_out_B[3]),
    .ADR3(DLX_EXinst_N76338),
    .O(\DLX_EXinst_N76338/GROM )
  );
  X_BUF \DLX_EXinst_N76338/XUSED  (
    .I(\DLX_EXinst_N76338/FROM ),
    .O(DLX_EXinst_N76338)
  );
  X_BUF \DLX_EXinst_N76338/YUSED  (
    .I(\DLX_EXinst_N76338/GROM ),
    .O(CHOICE3774)
  );
  defparam DLX_EXinst_Ker728961.INIT = 16'hEE22;
  X_LUT4 DLX_EXinst_Ker728961 (
    .ADR0(\DLX_EXinst_Mshift__n0023_Sh[4] ),
    .ADR1(DLX_IDinst_reg_out_B[2]),
    .ADR2(VCC),
    .ADR3(\DLX_EXinst_Mshift__n0023_Sh[0] ),
    .O(\DLX_EXinst_N72898/FROM )
  );
  defparam \DLX_EXinst__n0007<20>310_SW0 .INIT = 16'hDCCC;
  X_LUT4 \DLX_EXinst__n0007<20>310_SW0  (
    .ADR0(DLX_IDinst_reg_out_B[3]),
    .ADR1(CHOICE4696),
    .ADR2(DLX_EXinst_N75973),
    .ADR3(DLX_EXinst_N72898),
    .O(\DLX_EXinst_N72898/GROM )
  );
  X_BUF \DLX_EXinst_N72898/XUSED  (
    .I(\DLX_EXinst_N72898/FROM ),
    .O(DLX_EXinst_N72898)
  );
  X_BUF \DLX_EXinst_N72898/YUSED  (
    .I(\DLX_EXinst_N72898/GROM ),
    .O(N163473)
  );
  defparam DLX_EXinst_Ker73846.INIT = 16'hE4E4;
  X_LUT4 DLX_EXinst_Ker73846 (
    .ADR0(DLX_IDinst_reg_out_B[3]),
    .ADR1(N129951),
    .ADR2(\DLX_EXinst_Mshift__n0023_Sh[9] ),
    .ADR3(VCC),
    .O(\DLX_EXinst_N73848/FROM )
  );
  defparam DLX_EXinst_Ker738561.INIT = 16'hEE44;
  X_LUT4 DLX_EXinst_Ker738561 (
    .ADR0(DLX_IDinst_reg_out_B[3]),
    .ADR1(\DLX_EXinst_Mshift__n0023_Sh[19] ),
    .ADR2(VCC),
    .ADR3(\DLX_EXinst_Mshift__n0023_Sh[11] ),
    .O(\DLX_EXinst_N73848/GROM )
  );
  X_BUF \DLX_EXinst_N73848/XUSED  (
    .I(\DLX_EXinst_N73848/FROM ),
    .O(DLX_EXinst_N73848)
  );
  X_BUF \DLX_EXinst_N73848/YUSED  (
    .I(\DLX_EXinst_N73848/GROM ),
    .O(DLX_EXinst_N73858)
  );
  defparam DLX_IDinst_RegFile_28_30_1483.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_28_30_1483 (
    .I(DLX_IDinst_WB_data_eff[30]),
    .CE(DLX_IDinst__n0606),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_28_30)
  );
  defparam DLX_EXinst_Ker762831.INIT = 16'h0080;
  X_LUT4 DLX_EXinst_Ker762831 (
    .ADR0(DLX_IDinst_IR_opcode_field[1]),
    .ADR1(\DLX_IDinst_Imm[4] ),
    .ADR2(DLX_EXinst_N76041),
    .ADR3(DLX_IDinst_IR_opcode_field[0]),
    .O(\DLX_EXinst_N76285/GROM )
  );
  X_BUF \DLX_EXinst_N76285/YUSED  (
    .I(\DLX_EXinst_N76285/GROM ),
    .O(DLX_EXinst_N76285)
  );
  defparam DLX_EXinst_Ker764291.INIT = 16'hA0A0;
  X_LUT4 DLX_EXinst_Ker764291 (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst__n0081),
    .ADR3(VCC),
    .O(\DLX_EXinst_N76431/FROM )
  );
  defparam \DLX_EXinst__n0007<2>234 .INIT = 16'hE200;
  X_LUT4 \DLX_EXinst__n0007<2>234  (
    .ADR0(DLX_EXinst_N74731),
    .ADR1(DLX_IDinst_reg_out_B[2]),
    .ADR2(N131027),
    .ADR3(DLX_EXinst_N76431),
    .O(\DLX_EXinst_N76431/GROM )
  );
  X_BUF \DLX_EXinst_N76431/XUSED  (
    .I(\DLX_EXinst_N76431/FROM ),
    .O(DLX_EXinst_N76431)
  );
  X_BUF \DLX_EXinst_N76431/YUSED  (
    .I(\DLX_EXinst_N76431/GROM ),
    .O(CHOICE5568)
  );
  defparam DLX_EXinst_Ker739571.INIT = 16'hACAC;
  X_LUT4 DLX_EXinst_Ker739571 (
    .ADR0(DLX_EXinst__n0127),
    .ADR1(DLX_EXinst__n0109),
    .ADR2(DLX_EXinst__n0036),
    .ADR3(VCC),
    .O(\DLX_EXinst_ALU_result<9>/FROM )
  );
  defparam \DLX_EXinst__n0007<9>2491 .INIT = 16'hEECC;
  X_LUT4 \DLX_EXinst__n0007<9>2491  (
    .ADR0(DLX_EXinst__n0012[9]),
    .ADR1(CHOICE4558),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N73959),
    .O(\DLX_EXinst_ALU_result<9>/GROM )
  );
  X_BUF \DLX_EXinst_ALU_result<9>/XUSED  (
    .I(\DLX_EXinst_ALU_result<9>/FROM ),
    .O(DLX_EXinst_N73959)
  );
  X_BUF \DLX_EXinst_ALU_result<9>/YUSED  (
    .I(\DLX_EXinst_ALU_result<9>/GROM ),
    .O(N162810)
  );
  defparam DLX_EXinst_Ker764611.INIT = 16'h0004;
  X_LUT4 DLX_EXinst_Ker764611 (
    .ADR0(\DLX_IDinst_Imm[4] ),
    .ADR1(DLX_EXinst_N76041),
    .ADR2(DLX_IDinst_IR_opcode_field[1]),
    .ADR3(DLX_IDinst_IR_opcode_field[0]),
    .O(\DLX_EXinst_N76463/FROM )
  );
  defparam \DLX_EXinst__n0007<11>126 .INIT = 16'hEAC0;
  X_LUT4 \DLX_EXinst__n0007<11>126  (
    .ADR0(\DLX_EXinst_Mshift__n0021_Sh[43] ),
    .ADR1(DLX_EXinst_N76285),
    .ADR2(\DLX_EXinst_Mshift__n0022_Sh[59] ),
    .ADR3(DLX_EXinst_N76463),
    .O(\DLX_EXinst_N76463/GROM )
  );
  X_BUF \DLX_EXinst_N76463/XUSED  (
    .I(\DLX_EXinst_N76463/FROM ),
    .O(DLX_EXinst_N76463)
  );
  X_BUF \DLX_EXinst_N76463/YUSED  (
    .I(\DLX_EXinst_N76463/GROM ),
    .O(CHOICE4414)
  );
  defparam DLX_EXinst_Ker74699.INIT = 16'hF0AA;
  X_LUT4 DLX_EXinst_Ker74699 (
    .ADR0(N130825),
    .ADR1(VCC),
    .ADR2(\DLX_EXinst_Mshift__n0022_Sh[22] ),
    .ADR3(DLX_IDinst_Imm_3_1),
    .O(\DLX_EXinst_N74701/FROM )
  );
  defparam DLX_EXinst_Ker749341.INIT = 16'hFC0C;
  X_LUT4 DLX_EXinst_Ker749341 (
    .ADR0(VCC),
    .ADR1(\DLX_EXinst_Mshift__n0022_Sh[10] ),
    .ADR2(DLX_IDinst_Imm_3_1),
    .ADR3(\DLX_EXinst_Mshift__n0022_Sh[18] ),
    .O(\DLX_EXinst_N74701/GROM )
  );
  X_BUF \DLX_EXinst_N74701/XUSED  (
    .I(\DLX_EXinst_N74701/FROM ),
    .O(DLX_EXinst_N74701)
  );
  X_BUF \DLX_EXinst_N74701/YUSED  (
    .I(\DLX_EXinst_N74701/GROM ),
    .O(DLX_EXinst_N74936)
  );
  defparam DLX_IDinst_Ker10707440.INIT = 16'h00E0;
  X_LUT4 DLX_IDinst_Ker10707440 (
    .ADR0(CHOICE2112),
    .ADR1(DLX_IDinst_N108465),
    .ADR2(CHOICE2118),
    .ADR3(DLX_IDinst__n0166),
    .O(\CHOICE2119/FROM )
  );
  defparam DLX_IDinst__n011823_SW0.INIT = 16'hEEEA;
  X_LUT4 DLX_IDinst__n011823_SW0 (
    .ADR0(DLX_IDinst__n0453),
    .ADR1(DLX_IDinst_N107033),
    .ADR2(DLX_IDinst_N107405),
    .ADR3(CHOICE2119),
    .O(\CHOICE2119/GROM )
  );
  X_BUF \CHOICE2119/XUSED  (
    .I(\CHOICE2119/FROM ),
    .O(CHOICE2119)
  );
  X_BUF \CHOICE2119/YUSED  (
    .I(\CHOICE2119/GROM ),
    .O(N164702)
  );
  defparam DLX_EXinst_Ker764551.INIT = 16'h5054;
  X_LUT4 DLX_EXinst_Ker764551 (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(N148609),
    .ADR2(DLX_EXinst_N76421),
    .ADR3(DLX_IDinst_reg_out_B[5]),
    .O(\DLX_EXinst_N76457/FROM )
  );
  defparam \DLX_EXinst__n0007<2>189 .INIT = 16'hB800;
  X_LUT4 \DLX_EXinst__n0007<2>189  (
    .ADR0(N133408),
    .ADR1(DLX_IDinst_reg_out_B[2]),
    .ADR2(CHOICE5550),
    .ADR3(DLX_EXinst_N76457),
    .O(\DLX_EXinst_N76457/GROM )
  );
  X_BUF \DLX_EXinst_N76457/XUSED  (
    .I(\DLX_EXinst_N76457/FROM ),
    .O(DLX_EXinst_N76457)
  );
  X_BUF \DLX_EXinst_N76457/YUSED  (
    .I(\DLX_EXinst_N76457/GROM ),
    .O(CHOICE5553)
  );
  defparam DLX_EXinst_Ker764711.INIT = 16'h00CE;
  X_LUT4 DLX_EXinst_Ker764711 (
    .ADR0(N147520),
    .ADR1(DLX_EXinst_N76441),
    .ADR2(\DLX_IDinst_Imm[5] ),
    .ADR3(\DLX_IDinst_Imm[4] ),
    .O(\DLX_EXinst_N76473/FROM )
  );
  defparam \DLX_EXinst__n0007<2>65 .INIT = 16'hAC00;
  X_LUT4 \DLX_EXinst__n0007<2>65  (
    .ADR0(N134056),
    .ADR1(CHOICE5523),
    .ADR2(\DLX_IDinst_Imm[2] ),
    .ADR3(DLX_EXinst_N76473),
    .O(\DLX_EXinst_N76473/GROM )
  );
  X_BUF \DLX_EXinst_N76473/XUSED  (
    .I(\DLX_EXinst_N76473/FROM ),
    .O(DLX_EXinst_N76473)
  );
  X_BUF \DLX_EXinst_N76473/YUSED  (
    .I(\DLX_EXinst_N76473/GROM ),
    .O(CHOICE5526)
  );
  defparam DLX_EXinst_Ker746791.INIT = 16'hCFC0;
  X_LUT4 DLX_EXinst_Ker746791 (
    .ADR0(VCC),
    .ADR1(\DLX_EXinst_Mshift__n0019_Sh[18] ),
    .ADR2(DLX_IDinst_reg_out_B_3_1),
    .ADR3(\DLX_EXinst_Mshift__n0019_Sh[10] ),
    .O(\DLX_EXinst_N74681/GROM )
  );
  X_BUF \DLX_EXinst_N74681/YUSED  (
    .I(\DLX_EXinst_N74681/GROM ),
    .O(DLX_EXinst_N74681)
  );
  defparam DLX_EXinst_Ker74709.INIT = 16'hAACC;
  X_LUT4 DLX_EXinst_Ker74709 (
    .ADR0(\DLX_EXinst_Mshift__n0022_Sh[21] ),
    .ADR1(N130773),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_Imm_3_1),
    .O(\DLX_EXinst_N74711/FROM )
  );
  defparam DLX_EXinst_Ker749391.INIT = 16'hAFA0;
  X_LUT4 DLX_EXinst_Ker749391 (
    .ADR0(\DLX_EXinst_Mshift__n0022_Sh[19] ),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_Imm_3_1),
    .ADR3(\DLX_EXinst_Mshift__n0022_Sh[11] ),
    .O(\DLX_EXinst_N74711/GROM )
  );
  X_BUF \DLX_EXinst_N74711/XUSED  (
    .I(\DLX_EXinst_N74711/FROM ),
    .O(DLX_EXinst_N74711)
  );
  X_BUF \DLX_EXinst_N74711/YUSED  (
    .I(\DLX_EXinst_N74711/GROM ),
    .O(DLX_EXinst_N74941)
  );
  defparam DLX_IDinst_Ker10707449.INIT = 16'hFAFA;
  X_LUT4 DLX_IDinst_Ker10707449 (
    .ADR0(DLX_IDinst_N107405),
    .ADR1(VCC),
    .ADR2(CHOICE2119),
    .ADR3(VCC),
    .O(\N139656/GROM )
  );
  X_BUF \N139656/YUSED  (
    .I(\N139656/GROM ),
    .O(N139656)
  );
  defparam DLX_EXinst_Ker749491.INIT = 16'hF0CC;
  X_LUT4 DLX_EXinst_Ker749491 (
    .ADR0(VCC),
    .ADR1(\DLX_EXinst_Mshift__n0022_Sh[9] ),
    .ADR2(\DLX_EXinst_Mshift__n0022_Sh[17] ),
    .ADR3(DLX_IDinst_Imm_3_1),
    .O(\DLX_EXinst_N74951/GROM )
  );
  X_BUF \DLX_EXinst_N74951/YUSED  (
    .I(\DLX_EXinst_N74951/GROM ),
    .O(DLX_EXinst_N74951)
  );
  defparam DLX_EXinst_Ker764941.INIT = 16'h8080;
  X_LUT4 DLX_EXinst_Ker764941 (
    .ADR0(DLX_EXinst_N72710),
    .ADR1(DLX_EXinst_N75964),
    .ADR2(DLX_IDinst_reg_out_B[0]),
    .ADR3(VCC),
    .O(\DLX_EXinst_N76496/FROM )
  );
  defparam DLX_EXinst_Ker74134.INIT = 16'h8F88;
  X_LUT4 DLX_EXinst_Ker74134 (
    .ADR0(\DLX_IDinst_Imm[0] ),
    .ADR1(N131955),
    .ADR2(DLX_IDinst_reg_out_B[1]),
    .ADR3(DLX_EXinst_N76496),
    .O(\DLX_EXinst_N76496/GROM )
  );
  X_BUF \DLX_EXinst_N76496/XUSED  (
    .I(\DLX_EXinst_N76496/FROM ),
    .O(DLX_EXinst_N76496)
  );
  X_BUF \DLX_EXinst_N76496/YUSED  (
    .I(\DLX_EXinst_N76496/GROM ),
    .O(DLX_EXinst_N74136)
  );
  defparam DLX_EXinst_Ker764881.INIT = 16'h4040;
  X_LUT4 DLX_EXinst_Ker764881 (
    .ADR0(N146478),
    .ADR1(DLX_EXinst_N76412),
    .ADR2(DLX_EXinst__n0055),
    .ADR3(VCC),
    .O(\DLX_EXinst_N76490/FROM )
  );
  defparam DLX_EXinst_Ker74128_SW0.INIT = 16'h3000;
  X_LUT4 DLX_EXinst_Ker74128_SW0 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_Imm_1_1),
    .ADR2(\DLX_IDinst_Imm[0] ),
    .ADR3(DLX_EXinst_N76490),
    .O(\DLX_EXinst_N76490/GROM )
  );
  X_BUF \DLX_EXinst_N76490/XUSED  (
    .I(\DLX_EXinst_N76490/FROM ),
    .O(DLX_EXinst_N76490)
  );
  X_BUF \DLX_EXinst_N76490/YUSED  (
    .I(\DLX_EXinst_N76490/GROM ),
    .O(N131996)
  );
  defparam DLX_EXinst_Ker749691.INIT = 16'hAACC;
  X_LUT4 DLX_EXinst_Ker749691 (
    .ADR0(\DLX_EXinst_Mshift__n0022_Sh[24] ),
    .ADR1(\DLX_EXinst_Mshift__n0022_Sh[16] ),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_Imm_3_1),
    .O(\DLX_EXinst_N74971/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0020_Sh<80>1 .INIT = 16'hF3C0;
  X_LUT4 \DLX_EXinst_Mshift__n0020_Sh<80>1  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_Imm_2_1),
    .ADR2(DLX_EXinst_N72797),
    .ADR3(DLX_EXinst_N74971),
    .O(\DLX_EXinst_N74971/GROM )
  );
  X_BUF \DLX_EXinst_N74971/XUSED  (
    .I(\DLX_EXinst_N74971/FROM ),
    .O(DLX_EXinst_N74971)
  );
  X_BUF \DLX_EXinst_N74971/YUSED  (
    .I(\DLX_EXinst_N74971/GROM ),
    .O(\DLX_EXinst_Mshift__n0020_Sh[80] )
  );
  defparam \DLX_EXinst__n0007<6>241_SW0_SW0 .INIT = 16'hF5F4;
  X_LUT4 \DLX_EXinst__n0007<6>241_SW0_SW0  (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(CHOICE3889),
    .ADR2(CHOICE3900),
    .ADR3(CHOICE3886),
    .O(\N164607/FROM )
  );
  defparam \DLX_EXinst__n0007<6>241_SW0 .INIT = 16'hFFEA;
  X_LUT4 \DLX_EXinst__n0007<6>241_SW0  (
    .ADR0(CHOICE3897),
    .ADR1(CHOICE3880),
    .ADR2(DLX_IDinst_reg_out_A[6]),
    .ADR3(N164607),
    .O(\N164607/GROM )
  );
  X_BUF \N164607/XUSED  (
    .I(\N164607/FROM ),
    .O(N164607)
  );
  X_BUF \N164607/YUSED  (
    .I(\N164607/GROM ),
    .O(N163198)
  );
  defparam DLX_EXinst_Ker759911.INIT = 16'h0088;
  X_LUT4 DLX_EXinst_Ker759911 (
    .ADR0(DLX_EXinst__n0055),
    .ADR1(\DLX_IDinst_Imm[4] ),
    .ADR2(VCC),
    .ADR3(N146478),
    .O(\DLX_EXinst_N75993/FROM )
  );
  defparam \DLX_EXinst__n0007<19>14 .INIT = 16'h1000;
  X_LUT4 \DLX_EXinst__n0007<19>14  (
    .ADR0(\DLX_IDinst_Imm[3] ),
    .ADR1(\DLX_IDinst_Imm[2] ),
    .ADR2(\DLX_EXinst_Mshift__n0021_Sh[3] ),
    .ADR3(DLX_EXinst_N75993),
    .O(\DLX_EXinst_N75993/GROM )
  );
  X_BUF \DLX_EXinst_N75993/XUSED  (
    .I(\DLX_EXinst_N75993/FROM ),
    .O(DLX_EXinst_N75993)
  );
  X_BUF \DLX_EXinst_N75993/YUSED  (
    .I(\DLX_EXinst_N75993/GROM ),
    .O(CHOICE5278)
  );
  defparam DLX_IDinst_Ker10735446.INIT = 16'h3035;
  X_LUT4 DLX_IDinst_Ker10735446 (
    .ADR0(DLX_IDinst_Ker1084541_1),
    .ADR1(N163838),
    .ADR2(DLX_IDinst__n0637),
    .ADR3(N163836),
    .O(\N134590/FROM )
  );
  defparam \DLX_IDinst__n0146<6>48 .INIT = 16'hECA0;
  X_LUT4 \DLX_IDinst__n0146<6>48  (
    .ADR0(CHOICE3211),
    .ADR1(N163724),
    .ADR2(DLX_IDinst_N107105),
    .ADR3(N134590),
    .O(\N134590/GROM )
  );
  X_BUF \N134590/XUSED  (
    .I(\N134590/FROM ),
    .O(N134590)
  );
  X_BUF \N134590/YUSED  (
    .I(\N134590/GROM ),
    .O(CHOICE3213)
  );
  defparam DLX_IDinst_Ker10822663.INIT = 16'hCFCE;
  X_LUT4 DLX_IDinst_Ker10822663 (
    .ADR0(DLX_IDinst__n0104),
    .ADR1(N163831),
    .ADR2(DLX_IDinst__n0382),
    .ADR3(DLX_IDinst__n0100),
    .O(\CHOICE3386/FROM )
  );
  defparam DLX_IDinst_Ker108226127_SW0.INIT = 16'h000D;
  X_LUT4 DLX_IDinst_Ker108226127_SW0 (
    .ADR0(CHOICE3373),
    .ADR1(DLX_IDinst__n0106),
    .ADR2(CHOICE3377),
    .ADR3(CHOICE3386),
    .O(\CHOICE3386/GROM )
  );
  X_BUF \CHOICE3386/XUSED  (
    .I(\CHOICE3386/FROM ),
    .O(CHOICE3386)
  );
  X_BUF \CHOICE3386/YUSED  (
    .I(\CHOICE3386/GROM ),
    .O(N163124)
  );
  defparam DLX_IDinst_Ker10825782.INIT = 16'hCC04;
  X_LUT4 DLX_IDinst_Ker10825782 (
    .ADR0(DLX_IDinst__n0104),
    .ADR1(CHOICE3300),
    .ADR2(DLX_IDinst__n0100),
    .ADR3(DLX_IDinst__n0382),
    .O(\CHOICE3301/FROM )
  );
  defparam DLX_IDinst_Ker108257139.INIT = 16'h0302;
  X_LUT4 DLX_IDinst_Ker108257139 (
    .ADR0(N163258),
    .ADR1(DLX_IFinst_IR_latched[29]),
    .ADR2(DLX_IFinst_IR_latched[31]),
    .ADR3(CHOICE3301),
    .O(\CHOICE3301/GROM )
  );
  X_BUF \CHOICE3301/XUSED  (
    .I(\CHOICE3301/FROM ),
    .O(CHOICE3301)
  );
  X_BUF \CHOICE3301/YUSED  (
    .I(\CHOICE3301/GROM ),
    .O(N146700)
  );
  defparam DLX_EXinst_Mcompar__n0069_inst_cy_261_1484.INIT = 16'h8E8E;
  X_LUT4 DLX_EXinst_Mcompar__n0069_inst_cy_261_1484 (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(DLX_EXinst_Mcompar__n0069_inst_cy_260),
    .ADR2(DLX_IDinst_Imm_31_1),
    .ADR3(VCC),
    .O(\DLX_EXinst_Mcompar__n0069_inst_cy_261/FROM )
  );
  defparam \DLX_EXinst__n0007<0>414 .INIT = 16'h08C8;
  X_LUT4 \DLX_EXinst__n0007<0>414  (
    .ADR0(DLX_EXinst__n0061),
    .ADR1(DLX_IDinst_IR_opcode_field[0]),
    .ADR2(DLX_IDinst_IR_opcode_field[2]),
    .ADR3(DLX_EXinst_Mcompar__n0069_inst_cy_261),
    .O(\DLX_EXinst_Mcompar__n0069_inst_cy_261/GROM )
  );
  X_BUF \DLX_EXinst_Mcompar__n0069_inst_cy_261/XUSED  (
    .I(\DLX_EXinst_Mcompar__n0069_inst_cy_261/FROM ),
    .O(DLX_EXinst_Mcompar__n0069_inst_cy_261)
  );
  X_BUF \DLX_EXinst_Mcompar__n0069_inst_cy_261/YUSED  (
    .I(\DLX_EXinst_Mcompar__n0069_inst_cy_261/GROM ),
    .O(CHOICE5952)
  );
  defparam DLX_IDinst_RegFile_28_14_1485.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_28_14_1485 (
    .I(DLX_IDinst_WB_data_eff[14]),
    .CE(DLX_IDinst__n0606),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_28_14)
  );
  defparam DLX_IDinst_Ker10739725.INIT = 16'h00CC;
  X_LUT4 DLX_IDinst_Ker10739725 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_IR_opcode_field[5]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_IR_opcode_field[4]),
    .O(\CHOICE1326/FROM )
  );
  defparam DLX_IDinst_Ker10739730.INIT = 16'h5D00;
  X_LUT4 DLX_IDinst_Ker10739730 (
    .ADR0(DLX_IDinst_IR_opcode_field[1]),
    .ADR1(DLX_IDinst_IR_opcode_field[0]),
    .ADR2(DLX_IDinst_IR_opcode_field[2]),
    .ADR3(CHOICE1326),
    .O(\CHOICE1326/GROM )
  );
  X_BUF \CHOICE1326/XUSED  (
    .I(\CHOICE1326/FROM ),
    .O(CHOICE1326)
  );
  X_BUF \CHOICE1326/YUSED  (
    .I(\CHOICE1326/GROM ),
    .O(CHOICE1327)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_cy_229_1486.INIT = 16'hB2B2;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_cy_229_1486 (
    .ADR0(DLX_EXinst_Mcompar__n0093_inst_cy_228),
    .ADR1(DLX_IDinst_reg_out_A[31]),
    .ADR2(DLX_IDinst_reg_out_B[31]),
    .ADR3(VCC),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_229/FROM )
  );
  defparam \DLX_EXinst__n0007<0>257 .INIT = 16'h0454;
  X_LUT4 \DLX_EXinst__n0007<0>257  (
    .ADR0(\DLX_IDinst_Imm[0] ),
    .ADR1(DLX_EXinst__n0085),
    .ADR2(\DLX_IDinst_Imm[2] ),
    .ADR3(DLX_EXinst_Mcompar__n0093_inst_cy_229),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_229/GROM )
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_229/XUSED  (
    .I(\DLX_EXinst_Mcompar__n0093_inst_cy_229/FROM ),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_229)
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_229/YUSED  (
    .I(\DLX_EXinst_Mcompar__n0093_inst_cy_229/GROM ),
    .O(CHOICE5929)
  );
  defparam DLX_IDinst_Ker10757422.INIT = 16'h0C00;
  X_LUT4 DLX_IDinst_Ker10757422 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_N108574),
    .ADR2(DLX_IDinst__n0453),
    .ADR3(DLX_IDinst_N108221),
    .O(\CHOICE1693/FROM )
  );
  defparam DLX_IDinst_Ker10757425.INIT = 16'hFF0C;
  X_LUT4 DLX_IDinst_Ker10757425 (
    .ADR0(VCC),
    .ADR1(CHOICE1689),
    .ADR2(DLX_IDinst_IR_latched[30]),
    .ADR3(CHOICE1693),
    .O(\CHOICE1693/GROM )
  );
  X_BUF \CHOICE1693/XUSED  (
    .I(\CHOICE1693/FROM ),
    .O(CHOICE1693)
  );
  X_BUF \CHOICE1693/YUSED  (
    .I(\CHOICE1693/GROM ),
    .O(N137082)
  );
  defparam DLX_IDinst_RegFile_28_22_1487.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_28_22_1487 (
    .I(DLX_IDinst_WB_data_eff[22]),
    .CE(DLX_IDinst__n0606),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_28_22)
  );
  defparam \DLX_EXinst__n0007<2>3321_SW0 .INIT = 16'hFFEA;
  X_LUT4 \DLX_EXinst__n0007<2>3321_SW0  (
    .ADR0(CHOICE5579),
    .ADR1(DLX_EXinst_N74136),
    .ADR2(DLX_IDinst_reg_out_A[3]),
    .ADR3(N164587),
    .O(\DLX_EXinst_ALU_result<2>/FROM )
  );
  defparam \DLX_EXinst__n0007<2>3321 .INIT = 16'hFFF8;
  X_LUT4 \DLX_EXinst__n0007<2>3321  (
    .ADR0(DLX_EXinst__n0012[2]),
    .ADR1(DLX_EXinst_N73959),
    .ADR2(N136886),
    .ADR3(N163266),
    .O(\DLX_EXinst_ALU_result<2>/GROM )
  );
  X_BUF \DLX_EXinst_ALU_result<2>/XUSED  (
    .I(\DLX_EXinst_ALU_result<2>/FROM ),
    .O(N163266)
  );
  X_BUF \DLX_EXinst_ALU_result<2>/YUSED  (
    .I(\DLX_EXinst_ALU_result<2>/GROM ),
    .O(N162841)
  );
  defparam DLX_IDinst__n0115_SW0.INIT = 16'hAAEE;
  X_LUT4 DLX_IDinst__n0115_SW0 (
    .ADR0(DLX_IDinst_intr_slot),
    .ADR1(FREEZE_IBUF),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_delay_slot),
    .O(\N132148/FROM )
  );
  defparam DLX_IDinst__n0115_1488.INIT = 16'hFFEF;
  X_LUT4 DLX_IDinst__n0115_1488 (
    .ADR0(reset_IBUF),
    .ADR1(DLX_IDinst__n0376),
    .ADR2(DLX_EXinst__n0144),
    .ADR3(N132148),
    .O(\N132148/GROM )
  );
  X_BUF \N132148/XUSED  (
    .I(\N132148/FROM ),
    .O(N132148)
  );
  X_BUF \N132148/YUSED  (
    .I(\N132148/GROM ),
    .O(DLX_IDinst__n0115)
  );
  defparam DLX_IDinst_mem_write_1489.INIT = 1'b0;
  X_SFF DLX_IDinst_mem_write_1489 (
    .I(DLX_IDinst__n0141),
    .CE(DLX_IDinst__n0116),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_IDinst__n0115),
    .O(DLX_IDinst_mem_write)
  );
  defparam DLX_IDinst__n0141_SW0.INIT = 16'h5FFF;
  X_LUT4 DLX_IDinst__n0141_SW0 (
    .ADR0(DLX_IDinst__n0163),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_N107223),
    .ADR3(N139563),
    .O(\DLX_IDinst_mem_write/FROM )
  );
  defparam DLX_IDinst__n0141_1490.INIT = 16'h0020;
  X_LUT4 DLX_IDinst__n0141_1490 (
    .ADR0(DLX_IDinst__n0427),
    .ADR1(DLX_IDinst_N108456),
    .ADR2(DLX_IDinst_N108476),
    .ADR3(N132422),
    .O(DLX_IDinst__n0141)
  );
  X_BUF \DLX_IDinst_mem_write/XUSED  (
    .I(\DLX_IDinst_mem_write/FROM ),
    .O(N132422)
  );
  defparam \DLX_IDinst_slot_num_FFd2-In17_SW0 .INIT = 16'hFFFC;
  X_LUT4 \DLX_IDinst_slot_num_FFd2-In17_SW0  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_slot_num_FFd1),
    .ADR2(DLX_IDinst_slot_num_FFd4),
    .ADR3(DLX_IDinst_slot_num_FFd3),
    .O(\N163222/GROM )
  );
  X_BUF \N163222/YUSED  (
    .I(\N163222/GROM ),
    .O(N163222)
  );
  defparam DLX_IDinst__n0139_SW0.INIT = 16'hA3AF;
  X_LUT4 DLX_IDinst__n0139_SW0 (
    .ADR0(DLX_IDinst__n0629[1]),
    .ADR1(N139563),
    .ADR2(DLX_IDinst__n0453),
    .ADR3(DLX_IDinst_N107033),
    .O(\DLX_IDinst_mem_to_reg/FROM )
  );
  defparam DLX_IDinst__n0139_1491.INIT = 16'h0040;
  X_LUT4 DLX_IDinst__n0139_1491 (
    .ADR0(DLX_IDinst_N108456),
    .ADR1(DLX_IDinst__n0163),
    .ADR2(DLX_IDinst__n0164),
    .ADR3(N136962),
    .O(DLX_IDinst__n0139)
  );
  X_BUF \DLX_IDinst_mem_to_reg/XUSED  (
    .I(\DLX_IDinst_mem_to_reg/FROM ),
    .O(N136962)
  );
  defparam DLX_IDinst__n0530_SW1.INIT = 16'hEEE0;
  X_LUT4 DLX_IDinst__n0530_SW1 (
    .ADR0(DLX_IDinst_delay_slot),
    .ADR1(DLX_IDinst_intr_slot),
    .ADR2(DLX_IDinst_slot_num_FFd1),
    .ADR3(DLX_IDinst_slot_num_FFd3),
    .O(\N164089/FROM )
  );
  defparam DLX_IDinst__n0530_1492.INIT = 16'h0F05;
  X_LUT4 DLX_IDinst__n0530_1492 (
    .ADR0(DLX_IDinst__n0387),
    .ADR1(VCC),
    .ADR2(DLX_IDinst__n0391),
    .ADR3(N164089),
    .O(\N164089/GROM )
  );
  X_BUF \N164089/XUSED  (
    .I(\N164089/FROM ),
    .O(N164089)
  );
  X_BUF \N164089/YUSED  (
    .I(\N164089/GROM ),
    .O(DLX_IDinst__n0530)
  );
  defparam DLX_EXinst_Ker74128.INIT = 16'hDCCC;
  X_LUT4 DLX_EXinst_Ker74128 (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(N131996),
    .ADR2(DLX_EXinst_N76479),
    .ADR3(DLX_IDinst_reg_out_B[0]),
    .O(\DLX_EXinst_N74130/FROM )
  );
  defparam \DLX_EXinst__n0007<29>315 .INIT = 16'hECA0;
  X_LUT4 \DLX_EXinst__n0007<29>315  (
    .ADR0(DLX_EXinst_N73794),
    .ADR1(DLX_IDinst_reg_out_A[28]),
    .ADR2(DLX_IDinst_reg_out_A[27]),
    .ADR3(DLX_EXinst_N74130),
    .O(\DLX_EXinst_N74130/GROM )
  );
  X_BUF \DLX_EXinst_N74130/XUSED  (
    .I(\DLX_EXinst_N74130/FROM ),
    .O(DLX_EXinst_N74130)
  );
  X_BUF \DLX_EXinst_N74130/YUSED  (
    .I(\DLX_EXinst_N74130/GROM ),
    .O(CHOICE4841)
  );
  defparam DLX_EXinst_Ker73285.INIT = 16'hF8F0;
  X_LUT4 DLX_EXinst_Ker73285 (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(N132064),
    .ADR3(DLX_EXinst_N76479),
    .O(\DLX_EXinst_N73287/FROM )
  );
  defparam \DLX_EXinst__n0007<29>297 .INIT = 16'hF000;
  X_LUT4 \DLX_EXinst__n0007<29>297  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[26]),
    .ADR3(DLX_EXinst_N73287),
    .O(\DLX_EXinst_N73287/GROM )
  );
  X_BUF \DLX_EXinst_N73287/XUSED  (
    .I(\DLX_EXinst_N73287/FROM ),
    .O(DLX_EXinst_N73287)
  );
  X_BUF \DLX_EXinst_N73287/YUSED  (
    .I(\DLX_EXinst_N73287/GROM ),
    .O(CHOICE4837)
  );
  defparam DLX_EXinst_Ker72763.INIT = 16'hFFEF;
  X_LUT4 DLX_EXinst_Ker72763 (
    .ADR0(DLX_IDinst_IR_opcode_field[1]),
    .ADR1(N164077),
    .ADR2(DLX_IDinst_IR_opcode_field[3]),
    .ADR3(DLX_IDinst_IR_opcode_field[0]),
    .O(\DLX_EXinst_reg_out_B_EX<2>/FROM )
  );
  defparam \DLX_EXinst__n0008<15>1 .INIT = 16'hCC00;
  X_LUT4 \DLX_EXinst__n0008<15>1  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_B[15]),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N72765),
    .O(DLX_EXinst__n0008[15])
  );
  X_BUF \DLX_EXinst_reg_out_B_EX<2>/XUSED  (
    .I(\DLX_EXinst_reg_out_B_EX<2>/FROM ),
    .O(DLX_EXinst_N72765)
  );
  defparam DLX_IDinst__n0616_SW0.INIT = 16'hBBFF;
  X_LUT4 DLX_IDinst__n0616_SW0 (
    .ADR0(DLX_IDinst_delay_slot),
    .ADR1(DLX_IDinst_intr_slot),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_slot_num_FFd3),
    .O(\N132193/FROM )
  );
  defparam DLX_IDinst__n0616_1493.INIT = 16'h0515;
  X_LUT4 DLX_IDinst__n0616_1493 (
    .ADR0(DLX_IDinst__n0391),
    .ADR1(DLX_IDinst_slot_num_FFd1),
    .ADR2(DLX_IDinst__n0387),
    .ADR3(N132193),
    .O(\N132193/GROM )
  );
  X_BUF \N132193/XUSED  (
    .I(\N132193/FROM ),
    .O(N132193)
  );
  X_BUF \N132193/YUSED  (
    .I(\N132193/GROM ),
    .O(DLX_IDinst__n0616)
  );
  defparam DLX_EXinst_Ker74623.INIT = 16'hF888;
  X_LUT4 DLX_EXinst_Ker74623 (
    .ADR0(DLX_EXinst_N76496),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(N132037),
    .ADR3(\DLX_IDinst_Imm[0] ),
    .O(\DLX_EXinst_N74625/FROM )
  );
  defparam \DLX_EXinst__n0007<2>318 .INIT = 16'hF888;
  X_LUT4 \DLX_EXinst__n0007<2>318  (
    .ADR0(DLX_EXinst_N74347),
    .ADR1(DLX_IDinst_reg_out_A[4]),
    .ADR2(DLX_IDinst_reg_out_A[5]),
    .ADR3(DLX_EXinst_N74625),
    .O(\DLX_EXinst_N74625/GROM )
  );
  X_BUF \DLX_EXinst_N74625/XUSED  (
    .I(\DLX_EXinst_N74625/FROM ),
    .O(DLX_EXinst_N74625)
  );
  X_BUF \DLX_EXinst_N74625/YUSED  (
    .I(\DLX_EXinst_N74625/GROM ),
    .O(CHOICE5579)
  );
  defparam DLX_IDinst_Mmux__n0162_inst_mux_f5_201.INIT = 16'hCC0A;
  X_LUT4 DLX_IDinst_Mmux__n0162_inst_mux_f5_201 (
    .ADR0(DLX_MEMinst_RF_data_in[7]),
    .ADR1(DLX_MEMinst_RF_data_in[11]),
    .ADR2(DLX_MEMinst_opcode_of_WB[2]),
    .ADR3(DLX_MEMinst_opcode_of_WB[0]),
    .O(\DLX_IDinst_RegFile_10_11/FROM )
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<11>1 .INIT = 16'hEE22;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<11>1  (
    .ADR0(DLX_MEMinst_RF_data_in[11]),
    .ADR1(DLX_IDinst__n0161),
    .ADR2(VCC),
    .ADR3(DLX_IDinst__n0618[43]),
    .O(\DLX_IDinst_RegFile_10_11/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_10_11/XUSED  (
    .I(\DLX_IDinst_RegFile_10_11/FROM ),
    .O(DLX_IDinst__n0618[43])
  );
  X_BUF \DLX_IDinst_RegFile_10_11/YUSED  (
    .I(\DLX_IDinst_RegFile_10_11/GROM ),
    .O(DLX_IDinst_WB_data_eff[11])
  );
  defparam DLX_IDinst_Mmux__n0162_inst_mux_f5_211.INIT = 16'hDC10;
  X_LUT4 DLX_IDinst_Mmux__n0162_inst_mux_f5_211 (
    .ADR0(DLX_MEMinst_opcode_of_WB[2]),
    .ADR1(DLX_MEMinst_opcode_of_WB[0]),
    .ADR2(DLX_MEMinst_RF_data_in[7]),
    .ADR3(DLX_MEMinst_RF_data_in[12]),
    .O(\DLX_IDinst_RegFile_10_12/FROM )
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<12>1 .INIT = 16'hFA50;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<12>1  (
    .ADR0(DLX_IDinst__n0161),
    .ADR1(VCC),
    .ADR2(DLX_MEMinst_RF_data_in[12]),
    .ADR3(DLX_IDinst__n0618[44]),
    .O(\DLX_IDinst_RegFile_10_12/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_10_12/XUSED  (
    .I(\DLX_IDinst_RegFile_10_12/FROM ),
    .O(DLX_IDinst__n0618[44])
  );
  X_BUF \DLX_IDinst_RegFile_10_12/YUSED  (
    .I(\DLX_IDinst_RegFile_10_12/GROM ),
    .O(DLX_IDinst_WB_data_eff[12])
  );
  defparam DLX_IDinst_Mmux__n0162_inst_mux_f5_221.INIT = 16'hCC0A;
  X_LUT4 DLX_IDinst_Mmux__n0162_inst_mux_f5_221 (
    .ADR0(DLX_MEMinst_RF_data_in[7]),
    .ADR1(DLX_MEMinst_RF_data_in[13]),
    .ADR2(DLX_MEMinst_opcode_of_WB[2]),
    .ADR3(DLX_MEMinst_opcode_of_WB[0]),
    .O(\DLX_IDinst_RegFile_10_13/FROM )
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<13>1 .INIT = 16'hFC0C;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<13>1  (
    .ADR0(VCC),
    .ADR1(DLX_MEMinst_RF_data_in[13]),
    .ADR2(DLX_IDinst__n0161),
    .ADR3(DLX_IDinst__n0618[45]),
    .O(\DLX_IDinst_RegFile_10_13/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_10_13/XUSED  (
    .I(\DLX_IDinst_RegFile_10_13/FROM ),
    .O(DLX_IDinst__n0618[45])
  );
  X_BUF \DLX_IDinst_RegFile_10_13/YUSED  (
    .I(\DLX_IDinst_RegFile_10_13/GROM ),
    .O(DLX_IDinst_WB_data_eff[13])
  );
  defparam DLX_IDinst_Mmux__n0162_inst_mux_f5_231.INIT = 16'hBA10;
  X_LUT4 DLX_IDinst_Mmux__n0162_inst_mux_f5_231 (
    .ADR0(DLX_MEMinst_opcode_of_WB[0]),
    .ADR1(DLX_MEMinst_opcode_of_WB[2]),
    .ADR2(DLX_MEMinst_RF_data_in[7]),
    .ADR3(DLX_MEMinst_RF_data_in[14]),
    .O(\DLX_IDinst_RegFile_10_14/FROM )
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<14>1 .INIT = 16'hEE22;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<14>1  (
    .ADR0(DLX_MEMinst_RF_data_in[14]),
    .ADR1(DLX_IDinst__n0161),
    .ADR2(VCC),
    .ADR3(DLX_IDinst__n0618[46]),
    .O(\DLX_IDinst_RegFile_10_14/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_10_14/XUSED  (
    .I(\DLX_IDinst_RegFile_10_14/FROM ),
    .O(DLX_IDinst__n0618[46])
  );
  X_BUF \DLX_IDinst_RegFile_10_14/YUSED  (
    .I(\DLX_IDinst_RegFile_10_14/GROM ),
    .O(DLX_IDinst_WB_data_eff[14])
  );
  defparam DLX_IDinst_Mmux__n0162_inst_mux_f5_241.INIT = 16'h88B8;
  X_LUT4 DLX_IDinst_Mmux__n0162_inst_mux_f5_241 (
    .ADR0(DLX_MEMinst_RF_data_in[15]),
    .ADR1(DLX_MEMinst_opcode_of_WB[0]),
    .ADR2(DLX_MEMinst_RF_data_in[7]),
    .ADR3(DLX_MEMinst_opcode_of_WB[2]),
    .O(\DLX_IDinst_RegFile_10_15/FROM )
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<15>1 .INIT = 16'hEE44;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<15>1  (
    .ADR0(DLX_IDinst__n0161),
    .ADR1(DLX_MEMinst_RF_data_in[15]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst__n0618[47]),
    .O(\DLX_IDinst_RegFile_10_15/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_10_15/XUSED  (
    .I(\DLX_IDinst_RegFile_10_15/FROM ),
    .O(DLX_IDinst__n0618[47])
  );
  X_BUF \DLX_IDinst_RegFile_10_15/YUSED  (
    .I(\DLX_IDinst_RegFile_10_15/GROM ),
    .O(DLX_IDinst_WB_data_eff[15])
  );
  defparam DLX_IDinst_Mmux__n0162_inst_mux_f5_171.INIT = 16'hF022;
  X_LUT4 DLX_IDinst_Mmux__n0162_inst_mux_f5_171 (
    .ADR0(DLX_MEMinst_RF_data_in[7]),
    .ADR1(DLX_MEMinst_opcode_of_WB[2]),
    .ADR2(DLX_MEMinst_RF_data_in[8]),
    .ADR3(DLX_MEMinst_opcode_of_WB[0]),
    .O(\DLX_IDinst_RegFile_0_8/FROM )
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<8>1 .INIT = 16'hFC30;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<8>1  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst__n0161),
    .ADR2(DLX_MEMinst_RF_data_in[8]),
    .ADR3(DLX_IDinst__n0618[40]),
    .O(\DLX_IDinst_RegFile_0_8/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_0_8/XUSED  (
    .I(\DLX_IDinst_RegFile_0_8/FROM ),
    .O(DLX_IDinst__n0618[40])
  );
  X_BUF \DLX_IDinst_RegFile_0_8/YUSED  (
    .I(\DLX_IDinst_RegFile_0_8/GROM ),
    .O(DLX_IDinst_WB_data_eff[8])
  );
  defparam DLX_IDinst__n0387_SW1.INIT = 16'hFEFE;
  X_LUT4 DLX_IDinst__n0387_SW1 (
    .ADR0(DLX_IDinst_intr_slot),
    .ADR1(DLX_IDinst_counter[1]),
    .ADR2(DLX_IDinst__n0376),
    .ADR3(VCC),
    .O(\N164094/FROM )
  );
  defparam DLX_IDinst__n0387_1494.INIT = 16'hFFF4;
  X_LUT4 DLX_IDinst__n0387_1494 (
    .ADR0(DLX_IDinst_delay_slot),
    .ADR1(FREEZE_IBUF),
    .ADR2(DLX_IDinst_counter[0]),
    .ADR3(N164094),
    .O(\N164094/GROM )
  );
  X_BUF \N164094/XUSED  (
    .I(\N164094/FROM ),
    .O(N164094)
  );
  X_BUF \N164094/YUSED  (
    .I(\N164094/GROM ),
    .O(DLX_IDinst__n0387)
  );
  defparam DLX_IDinst_Mmux__n0162_inst_mux_f5_181.INIT = 16'hCE02;
  X_LUT4 DLX_IDinst_Mmux__n0162_inst_mux_f5_181 (
    .ADR0(DLX_MEMinst_RF_data_in[7]),
    .ADR1(DLX_MEMinst_opcode_of_WB[0]),
    .ADR2(DLX_MEMinst_opcode_of_WB[2]),
    .ADR3(DLX_MEMinst_RF_data_in[9]),
    .O(\DLX_IDinst_RegFile_0_9/FROM )
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<9>1 .INIT = 16'hFC30;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<9>1  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst__n0161),
    .ADR2(DLX_MEMinst_RF_data_in[9]),
    .ADR3(DLX_IDinst__n0618[41]),
    .O(\DLX_IDinst_RegFile_0_9/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_0_9/XUSED  (
    .I(\DLX_IDinst_RegFile_0_9/FROM ),
    .O(DLX_IDinst__n0618[41])
  );
  X_BUF \DLX_IDinst_RegFile_0_9/YUSED  (
    .I(\DLX_IDinst_RegFile_0_9/GROM ),
    .O(DLX_IDinst_WB_data_eff[9])
  );
  defparam DLX_IDinst_Mmux__n0162_inst_mux_f5_191.INIT = 16'hD1C0;
  X_LUT4 DLX_IDinst_Mmux__n0162_inst_mux_f5_191 (
    .ADR0(DLX_MEMinst_opcode_of_WB[2]),
    .ADR1(DLX_MEMinst_opcode_of_WB[0]),
    .ADR2(DLX_MEMinst_RF_data_in[10]),
    .ADR3(DLX_MEMinst_RF_data_in[7]),
    .O(\DLX_IDinst_RegFile_10_10/FROM )
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<10>1 .INIT = 16'hEE22;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<10>1  (
    .ADR0(DLX_MEMinst_RF_data_in[10]),
    .ADR1(DLX_IDinst__n0161),
    .ADR2(VCC),
    .ADR3(DLX_IDinst__n0618[42]),
    .O(\DLX_IDinst_RegFile_10_10/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_10_10/XUSED  (
    .I(\DLX_IDinst_RegFile_10_10/FROM ),
    .O(DLX_IDinst__n0618[42])
  );
  X_BUF \DLX_IDinst_RegFile_10_10/YUSED  (
    .I(\DLX_IDinst_RegFile_10_10/GROM ),
    .O(DLX_IDinst_WB_data_eff[10])
  );
  defparam DLX_IDinst__n0549_SW0.INIT = 16'hF3F0;
  X_LUT4 DLX_IDinst__n0549_SW0 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_delay_slot),
    .ADR2(DLX_IDinst__n0376),
    .ADR3(FREEZE_IBUF),
    .O(\N132252/FROM )
  );
  defparam DLX_IDinst__n0549_1495.INIT = 16'h0313;
  X_LUT4 DLX_IDinst__n0549_1495 (
    .ADR0(DLX_IDinst_intr_slot),
    .ADR1(DLX_IDinst__n0391),
    .ADR2(DLX_EXinst__n0144),
    .ADR3(N132252),
    .O(\N132252/GROM )
  );
  X_BUF \N132252/XUSED  (
    .I(\N132252/FROM ),
    .O(N132252)
  );
  X_BUF \N132252/YUSED  (
    .I(\N132252/GROM ),
    .O(DLX_IDinst__n0549)
  );
  defparam \DLX_EXinst__n0007<3>3321_SW0 .INIT = 16'hFFEC;
  X_LUT4 \DLX_EXinst__n0007<3>3321_SW0  (
    .ADR0(DLX_EXinst_N74136),
    .ADR1(CHOICE5503),
    .ADR2(DLX_IDinst_reg_out_A[4]),
    .ADR3(N164601),
    .O(\DLX_EXinst_ALU_result<3>/FROM )
  );
  defparam \DLX_EXinst__n0007<3>3321 .INIT = 16'hFFF8;
  X_LUT4 \DLX_EXinst__n0007<3>3321  (
    .ADR0(DLX_EXinst_N73959),
    .ADR1(DLX_EXinst__n0012[3]),
    .ADR2(N136886),
    .ADR3(N163274),
    .O(\DLX_EXinst_ALU_result<3>/GROM )
  );
  X_BUF \DLX_EXinst_ALU_result<3>/XUSED  (
    .I(\DLX_EXinst_ALU_result<3>/FROM ),
    .O(N163274)
  );
  X_BUF \DLX_EXinst_ALU_result<3>/YUSED  (
    .I(\DLX_EXinst_ALU_result<3>/GROM ),
    .O(N162860)
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<41>_SW0 .INIT = 16'h0C3F;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<41>_SW0  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_B_2_1),
    .ADR2(\DLX_EXinst_Mshift__n0023_Sh[5] ),
    .ADR3(\DLX_EXinst_Mshift__n0023_Sh[9] ),
    .O(\N131191/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<41> .INIT = 16'h2075;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<41>  (
    .ADR0(DLX_IDinst_reg_out_B_3_1),
    .ADR1(DLX_IDinst_reg_out_B_2_1),
    .ADR2(\DLX_EXinst_Mshift__n0023_Sh[1] ),
    .ADR3(N131191),
    .O(\N131191/GROM )
  );
  X_BUF \N131191/XUSED  (
    .I(\N131191/FROM ),
    .O(N131191)
  );
  X_BUF \N131191/YUSED  (
    .I(\N131191/GROM ),
    .O(\DLX_EXinst_Mshift__n0023_Sh[41] )
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<42>_SW0 .INIT = 16'h5533;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<42>_SW0  (
    .ADR0(\DLX_EXinst_Mshift__n0023_Sh[6] ),
    .ADR1(\DLX_EXinst_Mshift__n0023_Sh[10] ),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B_2_1),
    .O(\N131255/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<42> .INIT = 16'h4073;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<42>  (
    .ADR0(DLX_IDinst_reg_out_B_2_1),
    .ADR1(DLX_IDinst_reg_out_B_3_1),
    .ADR2(\DLX_EXinst_Mshift__n0023_Sh[2] ),
    .ADR3(N131255),
    .O(\N131255/GROM )
  );
  X_BUF \N131255/XUSED  (
    .I(\N131255/FROM ),
    .O(N131255)
  );
  X_BUF \N131255/YUSED  (
    .I(\N131255/GROM ),
    .O(\DLX_EXinst_Mshift__n0023_Sh[42] )
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<43>_SW0 .INIT = 16'h0F55;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<43>_SW0  (
    .ADR0(\DLX_EXinst_Mshift__n0023_Sh[11] ),
    .ADR1(VCC),
    .ADR2(\DLX_EXinst_Mshift__n0023_Sh[7] ),
    .ADR3(DLX_IDinst_reg_out_B_2_1),
    .O(\N131315/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<43> .INIT = 16'h085D;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<43>  (
    .ADR0(DLX_IDinst_reg_out_B_3_1),
    .ADR1(\DLX_EXinst_Mshift__n0023_Sh[3] ),
    .ADR2(DLX_IDinst_reg_out_B_2_1),
    .ADR3(N131315),
    .O(\N131315/GROM )
  );
  X_BUF \N131315/XUSED  (
    .I(\N131315/FROM ),
    .O(N131315)
  );
  X_BUF \N131315/YUSED  (
    .I(\N131315/GROM ),
    .O(\DLX_EXinst_Mshift__n0023_Sh[43] )
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<46>_SW0 .INIT = 16'h03F3;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<46>_SW0  (
    .ADR0(VCC),
    .ADR1(\DLX_EXinst_Mshift__n0023_Sh[14] ),
    .ADR2(DLX_IDinst_reg_out_B_2_1),
    .ADR3(\DLX_EXinst_Mshift__n0023_Sh[10] ),
    .O(\N130105/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<45>_SW0 .INIT = 16'h03F3;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<45>_SW0  (
    .ADR0(VCC),
    .ADR1(\DLX_EXinst_Mshift__n0023_Sh[13] ),
    .ADR2(DLX_IDinst_reg_out_B_2_1),
    .ADR3(\DLX_EXinst_Mshift__n0023_Sh[9] ),
    .O(\N130105/GROM )
  );
  X_BUF \N130105/XUSED  (
    .I(\N130105/FROM ),
    .O(N130105)
  );
  X_BUF \N130105/YUSED  (
    .I(\N130105/GROM ),
    .O(N130051)
  );
  defparam DLX_IDinst_RegFile_28_23_1496.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_28_23_1496 (
    .I(DLX_IDinst_WB_data_eff[23]),
    .CE(DLX_IDinst__n0606),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_28_23)
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<47>_SW0 .INIT = 16'h3355;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<47>_SW0  (
    .ADR0(\DLX_EXinst_Mshift__n0023_Sh[15] ),
    .ADR1(\DLX_EXinst_Mshift__n0023_Sh[11] ),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B_2_1),
    .O(\N130157/FROM )
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<47> .INIT = 16'hC0F3;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<47>  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_B_3_1),
    .ADR2(DLX_EXinst_N72913),
    .ADR3(N130157),
    .O(\N130157/GROM )
  );
  X_BUF \N130157/XUSED  (
    .I(\N130157/FROM ),
    .O(N130157)
  );
  X_BUF \N130157/YUSED  (
    .I(\N130157/GROM ),
    .O(\DLX_EXinst_Mshift__n0023_Sh[47] )
  );
  defparam \DLX_EXinst_Mshift__n0021_Sh<2> .INIT = 16'h3055;
  X_LUT4 \DLX_EXinst_Mshift__n0021_Sh<2>  (
    .ADR0(N131693),
    .ADR1(DLX_IDinst_Imm_0_1),
    .ADR2(DLX_IDinst_reg_out_A[0]),
    .ADR3(DLX_IDinst_Imm_1_1),
    .O(\DLX_EXinst_Mshift__n0021_Sh<2>/FROM )
  );
  defparam DLX_EXinst_Ker729911.INIT = 16'hFC30;
  X_LUT4 DLX_EXinst_Ker729911 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_Imm_2_1),
    .ADR2(\DLX_EXinst_Mshift__n0021_Sh[6] ),
    .ADR3(\DLX_EXinst_Mshift__n0021_Sh[2] ),
    .O(\DLX_EXinst_Mshift__n0021_Sh<2>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0021_Sh<2>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0021_Sh<2>/FROM ),
    .O(\DLX_EXinst_Mshift__n0021_Sh[2] )
  );
  X_BUF \DLX_EXinst_Mshift__n0021_Sh<2>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0021_Sh<2>/GROM ),
    .O(DLX_EXinst_N72993)
  );
  defparam \DLX_EXinst_Mshift__n0021_Sh<7> .INIT = 16'hAAF0;
  X_LUT4 \DLX_EXinst_Mshift__n0021_Sh<7>  (
    .ADR0(N130725),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N72933),
    .ADR3(DLX_IDinst_Imm_0_1),
    .O(\DLX_EXinst_Mshift__n0021_Sh<7>/FROM )
  );
  defparam DLX_EXinst_Ker729961.INIT = 16'hBB88;
  X_LUT4 DLX_EXinst_Ker729961 (
    .ADR0(\DLX_EXinst_Mshift__n0021_Sh[3] ),
    .ADR1(DLX_IDinst_Imm_2_1),
    .ADR2(VCC),
    .ADR3(\DLX_EXinst_Mshift__n0021_Sh[7] ),
    .O(\DLX_EXinst_Mshift__n0021_Sh<7>/GROM )
  );
  X_BUF \DLX_EXinst_Mshift__n0021_Sh<7>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0021_Sh<7>/FROM ),
    .O(\DLX_EXinst_Mshift__n0021_Sh[7] )
  );
  X_BUF \DLX_EXinst_Mshift__n0021_Sh<7>/YUSED  (
    .I(\DLX_EXinst_Mshift__n0021_Sh<7>/GROM ),
    .O(DLX_EXinst_N72998)
  );
  defparam DLX_IDinst_Ker1074218.INIT = 16'h2222;
  X_LUT4 DLX_IDinst_Ker1074218 (
    .ADR0(DLX_EXinst_opcode_of_EX_reg[4]),
    .ADR1(DLX_EXinst_opcode_of_EX_reg[5]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_EXinst_opcode_of_EX_reg<0>/FROM )
  );
  defparam DLX_IDinst_Ker10742112.INIT = 16'h8C00;
  X_LUT4 DLX_IDinst_Ker10742112 (
    .ADR0(DLX_EXinst_opcode_of_EX_reg[1]),
    .ADR1(DLX_EXinst_opcode_of_EX_reg[2]),
    .ADR2(DLX_EXinst_opcode_of_EX_reg[0]),
    .ADR3(CHOICE1354),
    .O(\DLX_EXinst_opcode_of_EX_reg<0>/GROM )
  );
  X_BUF \DLX_EXinst_opcode_of_EX_reg<0>/XUSED  (
    .I(\DLX_EXinst_opcode_of_EX_reg<0>/FROM ),
    .O(CHOICE1354)
  );
  X_BUF \DLX_EXinst_opcode_of_EX_reg<0>/YUSED  (
    .I(\DLX_EXinst_opcode_of_EX_reg<0>/GROM ),
    .O(CHOICE1355)
  );
  defparam DLX_IDinst_Ker1082521.INIT = 16'h0050;
  X_LUT4 DLX_IDinst_Ker1082521 (
    .ADR0(DLX_EXinst_opcode_of_EX_reg[1]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_opcode_of_EX_reg[3]),
    .ADR3(DLX_EXinst_opcode_of_EX_reg[5]),
    .O(\DLX_EXinst_opcode_of_EX_reg<1>/FROM )
  );
  defparam DLX_IDinst__n04391.INIT = 16'hEEAA;
  X_LUT4 DLX_IDinst__n04391 (
    .ADR0(N135272),
    .ADR1(N137212),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_N108254),
    .O(\DLX_EXinst_opcode_of_EX_reg<1>/GROM )
  );
  X_BUF \DLX_EXinst_opcode_of_EX_reg<1>/XUSED  (
    .I(\DLX_EXinst_opcode_of_EX_reg<1>/FROM ),
    .O(DLX_IDinst_N108254)
  );
  X_BUF \DLX_EXinst_opcode_of_EX_reg<1>/YUSED  (
    .I(\DLX_EXinst_opcode_of_EX_reg<1>/GROM ),
    .O(DLX_IDinst__n0439)
  );
  defparam DLX_IDinst_Ker10742125.INIT = 16'h3030;
  X_LUT4 DLX_IDinst_Ker10742125 (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_opcode_of_EX_reg[4]),
    .ADR2(DLX_EXinst_opcode_of_EX_reg[5]),
    .ADR3(VCC),
    .O(\DLX_EXinst_opcode_of_EX_reg<2>/FROM )
  );
  defparam DLX_IDinst_Ker10742130.INIT = 16'h7300;
  X_LUT4 DLX_IDinst_Ker10742130 (
    .ADR0(DLX_EXinst_opcode_of_EX_reg[2]),
    .ADR1(DLX_EXinst_opcode_of_EX_reg[1]),
    .ADR2(DLX_EXinst_opcode_of_EX_reg[0]),
    .ADR3(CHOICE1361),
    .O(\DLX_EXinst_opcode_of_EX_reg<2>/GROM )
  );
  X_BUF \DLX_EXinst_opcode_of_EX_reg<2>/XUSED  (
    .I(\DLX_EXinst_opcode_of_EX_reg<2>/FROM ),
    .O(CHOICE1361)
  );
  X_BUF \DLX_EXinst_opcode_of_EX_reg<2>/YUSED  (
    .I(\DLX_EXinst_opcode_of_EX_reg<2>/GROM ),
    .O(CHOICE1362)
  );
  defparam DLX_IDinst_RegFile_28_31_1497.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_28_31_1497 (
    .I(DLX_IDinst_WB_data_eff[31]),
    .CE(DLX_IDinst__n0606),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_28_31)
  );
  defparam DLX_IDinst_Ker107421112.INIT = 16'h00EA;
  X_LUT4 DLX_IDinst_Ker107421112 (
    .ADR0(CHOICE1381),
    .ADR1(CHOICE1373),
    .ADR2(DLX_EXinst_opcode_of_EX_reg[3]),
    .ADR3(DLX_EXinst_opcode_of_EX_reg[5]),
    .O(\DLX_EXinst_opcode_of_EX_reg<3>/FROM )
  );
  defparam DLX_IDinst_Ker107421126.INIT = 16'hFF32;
  X_LUT4 DLX_IDinst_Ker107421126 (
    .ADR0(CHOICE1355),
    .ADR1(DLX_EXinst_opcode_of_EX_reg[3]),
    .ADR2(CHOICE1362),
    .ADR3(CHOICE1383),
    .O(\DLX_EXinst_opcode_of_EX_reg<3>/GROM )
  );
  X_BUF \DLX_EXinst_opcode_of_EX_reg<3>/XUSED  (
    .I(\DLX_EXinst_opcode_of_EX_reg<3>/FROM ),
    .O(CHOICE1383)
  );
  X_BUF \DLX_EXinst_opcode_of_EX_reg<3>/YUSED  (
    .I(\DLX_EXinst_opcode_of_EX_reg<3>/GROM ),
    .O(N135272)
  );
  defparam DLX_IDinst_Ker10742196.INIT = 16'h0001;
  X_LUT4 DLX_IDinst_Ker10742196 (
    .ADR0(DLX_EXinst_opcode_of_EX_reg[2]),
    .ADR1(DLX_EXinst_opcode_of_EX_reg[0]),
    .ADR2(DLX_EXinst_opcode_of_EX_reg[4]),
    .ADR3(DLX_EXinst_opcode_of_EX_reg[1]),
    .O(\DLX_EXinst_opcode_of_EX_reg<4>/FROM )
  );
  defparam DLX_IDinst_Ker10742177.INIT = 16'h37FF;
  X_LUT4 DLX_IDinst_Ker10742177 (
    .ADR0(DLX_EXinst_opcode_of_EX_reg[0]),
    .ADR1(DLX_EXinst_opcode_of_EX_reg[4]),
    .ADR2(DLX_EXinst_opcode_of_EX_reg[1]),
    .ADR3(DLX_EXinst_opcode_of_EX_reg[2]),
    .O(\DLX_EXinst_opcode_of_EX_reg<4>/GROM )
  );
  X_BUF \DLX_EXinst_opcode_of_EX_reg<4>/XUSED  (
    .I(\DLX_EXinst_opcode_of_EX_reg<4>/FROM ),
    .O(CHOICE1381)
  );
  X_BUF \DLX_EXinst_opcode_of_EX_reg<4>/YUSED  (
    .I(\DLX_EXinst_opcode_of_EX_reg<4>/GROM ),
    .O(CHOICE1373)
  );
  X_OPAD \DM_write/PAD  (
    .PAD(DM_write)
  );
  X_TRI DM_write_OBUF (
    .I(\DM_write/OUTMUX ),
    .CTL(\DM_write/ENABLE ),
    .O(DM_write)
  );
  X_INV \DM_write/ENABLEINV  (
    .I(\DM_write/TORGTS ),
    .O(\DM_write/ENABLE )
  );
  X_BUF \DM_write/GTS_OR  (
    .I(GTS),
    .O(\DM_write/TORGTS )
  );
  X_BUF \DM_write/OUTMUX_1498  (
    .I(DLX_EXinst_mem_write_EX_1),
    .O(\DM_write/OUTMUX )
  );
  X_BUF \DM_write/OMUX  (
    .I(DLX_IDinst_mem_write),
    .O(\DM_write/OD )
  );
  X_OPAD \CLI/PAD  (
    .PAD(CLI)
  );
  X_TRI CLI_OBUF (
    .I(\CLI/OUTMUX ),
    .CTL(\CLI/ENABLE ),
    .O(CLI)
  );
  X_INV \CLI/ENABLEINV  (
    .I(\CLI/TORGTS ),
    .O(\CLI/ENABLE )
  );
  X_BUF \CLI/GTS_OR  (
    .I(GTS),
    .O(\CLI/TORGTS )
  );
  X_BUF \CLI/OUTMUX_1499  (
    .I(DLX_IDinst_CLI_1),
    .O(\CLI/OUTMUX )
  );
  X_BUF \CLI/OMUX  (
    .I(DLX_IDinst__n0153),
    .O(\CLI/OD )
  );
  X_IPAD \INT/PAD  (
    .PAD(INT)
  );
  X_BUF \INT/IMUX  (
    .I(\INT/IBUF ),
    .O(INT_IBUF)
  );
  X_BUF INT_IBUF_1500 (
    .I(INT),
    .O(\INT/IBUF )
  );
  X_OPAD \NPC_eff<0>/PAD  (
    .PAD(NPC_eff[0])
  );
  X_TRI NPC_eff_0_OBUF (
    .I(\NPC_eff<0>/OUTMUX ),
    .CTL(\NPC_eff<0>/ENABLE ),
    .O(NPC_eff[0])
  );
  X_INV \NPC_eff<0>/ENABLEINV  (
    .I(\NPC_eff<0>/TORGTS ),
    .O(\NPC_eff<0>/ENABLE )
  );
  X_BUF \NPC_eff<0>/GTS_OR  (
    .I(GTS),
    .O(\NPC_eff<0>/TORGTS )
  );
  X_BUF \NPC_eff<0>/OUTMUX_1501  (
    .I(DLX_IFinst_NPC_0_1),
    .O(\NPC_eff<0>/OUTMUX )
  );
  X_BUF \NPC_eff<0>/OMUX  (
    .I(DLX_IFinst__n0001[0]),
    .O(\NPC_eff<0>/OD )
  );
  X_OPAD \NPC_eff<1>/PAD  (
    .PAD(NPC_eff[1])
  );
  X_TRI NPC_eff_1_OBUF (
    .I(\NPC_eff<1>/OUTMUX ),
    .CTL(\NPC_eff<1>/ENABLE ),
    .O(NPC_eff[1])
  );
  X_INV \NPC_eff<1>/ENABLEINV  (
    .I(\NPC_eff<1>/TORGTS ),
    .O(\NPC_eff<1>/ENABLE )
  );
  X_BUF \NPC_eff<1>/GTS_OR  (
    .I(GTS),
    .O(\NPC_eff<1>/TORGTS )
  );
  X_BUF \NPC_eff<1>/OUTMUX_1502  (
    .I(DLX_IFinst_NPC_1_1),
    .O(\NPC_eff<1>/OUTMUX )
  );
  X_BUF \NPC_eff<1>/OMUX  (
    .I(DLX_IFinst__n0001[1]),
    .O(\NPC_eff<1>/OD )
  );
  defparam DLX_IDinst_RegFile_28_15_1503.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_28_15_1503 (
    .I(DLX_IDinst_WB_data_eff[15]),
    .CE(DLX_IDinst__n0606),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_28_15)
  );
  X_OPAD \NPC_eff<2>/PAD  (
    .PAD(NPC_eff[2])
  );
  X_TRI NPC_eff_2_OBUF (
    .I(\NPC_eff<2>/OUTMUX ),
    .CTL(\NPC_eff<2>/ENABLE ),
    .O(NPC_eff[2])
  );
  X_INV \NPC_eff<2>/ENABLEINV  (
    .I(\NPC_eff<2>/TORGTS ),
    .O(\NPC_eff<2>/ENABLE )
  );
  X_BUF \NPC_eff<2>/GTS_OR  (
    .I(GTS),
    .O(\NPC_eff<2>/TORGTS )
  );
  X_BUF \NPC_eff<2>/OUTMUX_1504  (
    .I(DLX_IFinst_NPC_2_1),
    .O(\NPC_eff<2>/OUTMUX )
  );
  X_BUF \NPC_eff<2>/OMUX  (
    .I(DLX_IFinst__n0001[2]),
    .O(\NPC_eff<2>/OD )
  );
  X_OPAD \NPC_eff<3>/PAD  (
    .PAD(NPC_eff[3])
  );
  X_TRI NPC_eff_3_OBUF (
    .I(\NPC_eff<3>/OUTMUX ),
    .CTL(\NPC_eff<3>/ENABLE ),
    .O(NPC_eff[3])
  );
  X_INV \NPC_eff<3>/ENABLEINV  (
    .I(\NPC_eff<3>/TORGTS ),
    .O(\NPC_eff<3>/ENABLE )
  );
  X_BUF \NPC_eff<3>/GTS_OR  (
    .I(GTS),
    .O(\NPC_eff<3>/TORGTS )
  );
  X_BUF \NPC_eff<3>/OUTMUX_1505  (
    .I(DLX_IFinst_NPC_3_1),
    .O(\NPC_eff<3>/OUTMUX )
  );
  X_BUF \NPC_eff<3>/OMUX  (
    .I(DLX_IFinst__n0001[3]),
    .O(\NPC_eff<3>/OD )
  );
  X_OPAD \NPC_eff<4>/PAD  (
    .PAD(NPC_eff[4])
  );
  X_TRI NPC_eff_4_OBUF (
    .I(\NPC_eff<4>/OUTMUX ),
    .CTL(\NPC_eff<4>/ENABLE ),
    .O(NPC_eff[4])
  );
  X_INV \NPC_eff<4>/ENABLEINV  (
    .I(\NPC_eff<4>/TORGTS ),
    .O(\NPC_eff<4>/ENABLE )
  );
  X_BUF \NPC_eff<4>/GTS_OR  (
    .I(GTS),
    .O(\NPC_eff<4>/TORGTS )
  );
  X_BUF \NPC_eff<4>/OUTMUX_1506  (
    .I(DLX_IFinst_NPC_4_1),
    .O(\NPC_eff<4>/OUTMUX )
  );
  X_BUF \NPC_eff<4>/OMUX  (
    .I(DLX_IFinst__n0001[4]),
    .O(\NPC_eff<4>/OD )
  );
  X_OPAD \NPC_eff<5>/PAD  (
    .PAD(NPC_eff[5])
  );
  X_TRI NPC_eff_5_OBUF (
    .I(\NPC_eff<5>/OUTMUX ),
    .CTL(\NPC_eff<5>/ENABLE ),
    .O(NPC_eff[5])
  );
  X_INV \NPC_eff<5>/ENABLEINV  (
    .I(\NPC_eff<5>/TORGTS ),
    .O(\NPC_eff<5>/ENABLE )
  );
  X_BUF \NPC_eff<5>/GTS_OR  (
    .I(GTS),
    .O(\NPC_eff<5>/TORGTS )
  );
  X_BUF \NPC_eff<5>/OUTMUX_1507  (
    .I(DLX_IFinst_NPC_5_1),
    .O(\NPC_eff<5>/OUTMUX )
  );
  X_BUF \NPC_eff<5>/OMUX  (
    .I(DLX_IFinst__n0001[5]),
    .O(\NPC_eff<5>/OD )
  );
  X_OPAD \NPC_eff<6>/PAD  (
    .PAD(NPC_eff[6])
  );
  X_TRI NPC_eff_6_OBUF (
    .I(\NPC_eff<6>/OUTMUX ),
    .CTL(\NPC_eff<6>/ENABLE ),
    .O(NPC_eff[6])
  );
  X_INV \NPC_eff<6>/ENABLEINV  (
    .I(\NPC_eff<6>/TORGTS ),
    .O(\NPC_eff<6>/ENABLE )
  );
  X_BUF \NPC_eff<6>/GTS_OR  (
    .I(GTS),
    .O(\NPC_eff<6>/TORGTS )
  );
  X_BUF \NPC_eff<6>/OUTMUX_1508  (
    .I(DLX_IFinst_NPC_6_1),
    .O(\NPC_eff<6>/OUTMUX )
  );
  X_BUF \NPC_eff<6>/OMUX  (
    .I(DLX_IFinst__n0001[6]),
    .O(\NPC_eff<6>/OD )
  );
  X_OPAD \NPC_eff<7>/PAD  (
    .PAD(NPC_eff[7])
  );
  X_TRI NPC_eff_7_OBUF (
    .I(\NPC_eff<7>/OUTMUX ),
    .CTL(\NPC_eff<7>/ENABLE ),
    .O(NPC_eff[7])
  );
  X_INV \NPC_eff<7>/ENABLEINV  (
    .I(\NPC_eff<7>/TORGTS ),
    .O(\NPC_eff<7>/ENABLE )
  );
  X_BUF \NPC_eff<7>/GTS_OR  (
    .I(GTS),
    .O(\NPC_eff<7>/TORGTS )
  );
  X_BUF \NPC_eff<7>/OUTMUX_1509  (
    .I(DLX_IFinst_NPC_7_1),
    .O(\NPC_eff<7>/OUTMUX )
  );
  X_BUF \NPC_eff<7>/OMUX  (
    .I(DLX_IFinst__n0001[7]),
    .O(\NPC_eff<7>/OD )
  );
  X_OPAD \NPC_eff<8>/PAD  (
    .PAD(NPC_eff[8])
  );
  X_TRI NPC_eff_8_OBUF (
    .I(\NPC_eff<8>/OUTMUX ),
    .CTL(\NPC_eff<8>/ENABLE ),
    .O(NPC_eff[8])
  );
  X_INV \NPC_eff<8>/ENABLEINV  (
    .I(\NPC_eff<8>/TORGTS ),
    .O(\NPC_eff<8>/ENABLE )
  );
  X_BUF \NPC_eff<8>/GTS_OR  (
    .I(GTS),
    .O(\NPC_eff<8>/TORGTS )
  );
  X_BUF \NPC_eff<8>/OUTMUX_1510  (
    .I(DLX_IFinst_NPC_8_1),
    .O(\NPC_eff<8>/OUTMUX )
  );
  X_BUF \NPC_eff<8>/OMUX  (
    .I(DLX_IFinst__n0001[8]),
    .O(\NPC_eff<8>/OD )
  );
  X_OPAD \NPC_eff<9>/PAD  (
    .PAD(NPC_eff[9])
  );
  X_TRI NPC_eff_9_OBUF (
    .I(\NPC_eff<9>/OUTMUX ),
    .CTL(\NPC_eff<9>/ENABLE ),
    .O(NPC_eff[9])
  );
  X_INV \NPC_eff<9>/ENABLEINV  (
    .I(\NPC_eff<9>/TORGTS ),
    .O(\NPC_eff<9>/ENABLE )
  );
  X_BUF \NPC_eff<9>/GTS_OR  (
    .I(GTS),
    .O(\NPC_eff<9>/TORGTS )
  );
  X_BUF \NPC_eff<9>/OUTMUX_1511  (
    .I(DLX_IFinst_NPC_9_1),
    .O(\NPC_eff<9>/OUTMUX )
  );
  X_BUF \NPC_eff<9>/OMUX  (
    .I(DLX_IFinst__n0001[9]),
    .O(\NPC_eff<9>/OD )
  );
  X_OPAD \mask<0>/PAD  (
    .PAD(mask[0])
  );
  X_TRI mask_0_OBUF_1512 (
    .I(\mask<0>/OUTMUX ),
    .CTL(\mask<0>/ENABLE ),
    .O(mask[0])
  );
  X_INV \mask<0>/ENABLEINV  (
    .I(\mask<0>/TORGTS ),
    .O(\mask<0>/ENABLE )
  );
  X_BUF \mask<0>/GTS_OR  (
    .I(GTS),
    .O(\mask<0>/TORGTS )
  );
  X_BUF \mask<0>/OUTMUX_1513  (
    .I(mask_0_OBUF),
    .O(\mask<0>/OUTMUX )
  );
  X_OPAD \mask<3>/PAD  (
    .PAD(mask[3])
  );
  X_TRI mask_3_OBUF_1514 (
    .I(\mask<3>/OUTMUX ),
    .CTL(\mask<3>/ENABLE ),
    .O(mask[3])
  );
  X_INV \mask<3>/ENABLEINV  (
    .I(\mask<3>/TORGTS ),
    .O(\mask<3>/ENABLE )
  );
  X_BUF \mask<3>/GTS_OR  (
    .I(GTS),
    .O(\mask<3>/TORGTS )
  );
  X_BUF \mask<3>/OUTMUX_1515  (
    .I(mask_3_OBUF),
    .O(\mask<3>/OUTMUX )
  );
  X_OPAD \NPC_eff<10>/PAD  (
    .PAD(NPC_eff[10])
  );
  X_TRI NPC_eff_10_OBUF (
    .I(\NPC_eff<10>/OUTMUX ),
    .CTL(\NPC_eff<10>/ENABLE ),
    .O(NPC_eff[10])
  );
  X_INV \NPC_eff<10>/ENABLEINV  (
    .I(\NPC_eff<10>/TORGTS ),
    .O(\NPC_eff<10>/ENABLE )
  );
  X_BUF \NPC_eff<10>/GTS_OR  (
    .I(GTS),
    .O(\NPC_eff<10>/TORGTS )
  );
  X_BUF \NPC_eff<10>/OUTMUX_1516  (
    .I(DLX_IFinst_NPC_10_1),
    .O(\NPC_eff<10>/OUTMUX )
  );
  X_BUF \NPC_eff<10>/OMUX  (
    .I(DLX_IFinst__n0001[10]),
    .O(\NPC_eff<10>/OD )
  );
  X_OPAD \NPC_eff<11>/PAD  (
    .PAD(NPC_eff[11])
  );
  X_TRI NPC_eff_11_OBUF (
    .I(\NPC_eff<11>/OUTMUX ),
    .CTL(\NPC_eff<11>/ENABLE ),
    .O(NPC_eff[11])
  );
  X_INV \NPC_eff<11>/ENABLEINV  (
    .I(\NPC_eff<11>/TORGTS ),
    .O(\NPC_eff<11>/ENABLE )
  );
  X_BUF \NPC_eff<11>/GTS_OR  (
    .I(GTS),
    .O(\NPC_eff<11>/TORGTS )
  );
  X_BUF \NPC_eff<11>/OUTMUX_1517  (
    .I(DLX_IFinst_NPC_11_1),
    .O(\NPC_eff<11>/OUTMUX )
  );
  X_BUF \NPC_eff<11>/OMUX  (
    .I(DLX_IFinst__n0001[11]),
    .O(\NPC_eff<11>/OD )
  );
  X_OPAD \NPC_eff<12>/PAD  (
    .PAD(NPC_eff[12])
  );
  X_TRI NPC_eff_12_OBUF (
    .I(\NPC_eff<12>/OUTMUX ),
    .CTL(\NPC_eff<12>/ENABLE ),
    .O(NPC_eff[12])
  );
  X_INV \NPC_eff<12>/ENABLEINV  (
    .I(\NPC_eff<12>/TORGTS ),
    .O(\NPC_eff<12>/ENABLE )
  );
  X_BUF \NPC_eff<12>/GTS_OR  (
    .I(GTS),
    .O(\NPC_eff<12>/TORGTS )
  );
  X_BUF \NPC_eff<12>/OUTMUX_1518  (
    .I(DLX_IFinst_NPC_12_1),
    .O(\NPC_eff<12>/OUTMUX )
  );
  X_BUF \NPC_eff<12>/OMUX  (
    .I(DLX_IFinst__n0001[12]),
    .O(\NPC_eff<12>/OD )
  );
  X_OPAD \NPC_eff<13>/PAD  (
    .PAD(NPC_eff[13])
  );
  X_TRI NPC_eff_13_OBUF (
    .I(\NPC_eff<13>/OUTMUX ),
    .CTL(\NPC_eff<13>/ENABLE ),
    .O(NPC_eff[13])
  );
  X_INV \NPC_eff<13>/ENABLEINV  (
    .I(\NPC_eff<13>/TORGTS ),
    .O(\NPC_eff<13>/ENABLE )
  );
  X_BUF \NPC_eff<13>/GTS_OR  (
    .I(GTS),
    .O(\NPC_eff<13>/TORGTS )
  );
  X_BUF \NPC_eff<13>/OUTMUX_1519  (
    .I(DLX_IFinst_NPC_13_1),
    .O(\NPC_eff<13>/OUTMUX )
  );
  X_BUF \NPC_eff<13>/OMUX  (
    .I(DLX_IFinst__n0001[13]),
    .O(\NPC_eff<13>/OD )
  );
  X_OPAD \NPC_eff<14>/PAD  (
    .PAD(NPC_eff[14])
  );
  X_TRI NPC_eff_14_OBUF (
    .I(\NPC_eff<14>/OUTMUX ),
    .CTL(\NPC_eff<14>/ENABLE ),
    .O(NPC_eff[14])
  );
  X_INV \NPC_eff<14>/ENABLEINV  (
    .I(\NPC_eff<14>/TORGTS ),
    .O(\NPC_eff<14>/ENABLE )
  );
  X_BUF \NPC_eff<14>/GTS_OR  (
    .I(GTS),
    .O(\NPC_eff<14>/TORGTS )
  );
  X_BUF \NPC_eff<14>/OUTMUX_1520  (
    .I(DLX_IFinst_NPC_14_1),
    .O(\NPC_eff<14>/OUTMUX )
  );
  X_BUF \NPC_eff<14>/OMUX  (
    .I(DLX_IFinst__n0001[14]),
    .O(\NPC_eff<14>/OD )
  );
  X_OPAD \NPC_eff<15>/PAD  (
    .PAD(NPC_eff[15])
  );
  X_TRI NPC_eff_15_OBUF (
    .I(\NPC_eff<15>/OUTMUX ),
    .CTL(\NPC_eff<15>/ENABLE ),
    .O(NPC_eff[15])
  );
  X_INV \NPC_eff<15>/ENABLEINV  (
    .I(\NPC_eff<15>/TORGTS ),
    .O(\NPC_eff<15>/ENABLE )
  );
  X_BUF \NPC_eff<15>/GTS_OR  (
    .I(GTS),
    .O(\NPC_eff<15>/TORGTS )
  );
  X_BUF \NPC_eff<15>/OUTMUX_1521  (
    .I(DLX_IFinst_NPC_15_1),
    .O(\NPC_eff<15>/OUTMUX )
  );
  X_BUF \NPC_eff<15>/OMUX  (
    .I(DLX_IFinst__n0001[15]),
    .O(\NPC_eff<15>/OD )
  );
  X_OPAD \DM_write_data<0>/PAD  (
    .PAD(DM_write_data[0])
  );
  X_TRI DM_write_data_0_OBUF (
    .I(\DM_write_data<0>/OUTMUX ),
    .CTL(\DM_write_data<0>/ENABLE ),
    .O(DM_write_data[0])
  );
  X_INV \DM_write_data<0>/ENABLEINV  (
    .I(\DM_write_data<0>/TORGTS ),
    .O(\DM_write_data<0>/ENABLE )
  );
  X_BUF \DM_write_data<0>/GTS_OR  (
    .I(GTS),
    .O(\DM_write_data<0>/TORGTS )
  );
  X_BUF \DM_write_data<0>/OUTMUX_1522  (
    .I(DLX_EXinst_reg_out_B_EX_0_1),
    .O(\DM_write_data<0>/OUTMUX )
  );
  X_BUF \DM_write_data<0>/OMUX  (
    .I(DLX_IDinst_reg_out_B[0]),
    .O(\DM_write_data<0>/OD )
  );
  X_OPAD \blue<0>/PAD  (
    .PAD(blue[0])
  );
  X_TRI blue_0_OBUF_1523 (
    .I(\blue<0>/OUTMUX ),
    .CTL(\blue<0>/ENABLE ),
    .O(blue[0])
  );
  X_INV \blue<0>/ENABLEINV  (
    .I(\blue<0>/TORGTS ),
    .O(\blue<0>/ENABLE )
  );
  X_BUF \blue<0>/GTS_OR  (
    .I(GTS),
    .O(\blue<0>/TORGTS )
  );
  X_BUF \blue<0>/OUTMUX_1524  (
    .I(blue_0_OBUF),
    .O(\blue<0>/OUTMUX )
  );
  X_OPAD \blue<1>/PAD  (
    .PAD(blue[1])
  );
  X_TRI blue_1_OBUF_1525 (
    .I(\blue<1>/OUTMUX ),
    .CTL(\blue<1>/ENABLE ),
    .O(blue[1])
  );
  X_INV \blue<1>/ENABLEINV  (
    .I(\blue<1>/TORGTS ),
    .O(\blue<1>/ENABLE )
  );
  X_BUF \blue<1>/GTS_OR  (
    .I(GTS),
    .O(\blue<1>/TORGTS )
  );
  X_BUF \blue<1>/OUTMUX_1526  (
    .I(blue_1_OBUF),
    .O(\blue<1>/OUTMUX )
  );
  X_OPAD \blue<2>/PAD  (
    .PAD(blue[2])
  );
  X_TRI blue_2_OBUF_1527 (
    .I(\blue<2>/OUTMUX ),
    .CTL(\blue<2>/ENABLE ),
    .O(blue[2])
  );
  X_INV \blue<2>/ENABLEINV  (
    .I(\blue<2>/TORGTS ),
    .O(\blue<2>/ENABLE )
  );
  X_BUF \blue<2>/GTS_OR  (
    .I(GTS),
    .O(\blue<2>/TORGTS )
  );
  X_BUF \blue<2>/OUTMUX_1528  (
    .I(blue_2_OBUF),
    .O(\blue<2>/OUTMUX )
  );
  X_OPAD \mask<1>/PAD  (
    .PAD(mask[1])
  );
  X_TRI mask_1_OBUF_1529 (
    .I(\mask<1>/OUTMUX ),
    .CTL(\mask<1>/ENABLE ),
    .O(mask[1])
  );
  X_INV \mask<1>/ENABLEINV  (
    .I(\mask<1>/TORGTS ),
    .O(\mask<1>/ENABLE )
  );
  X_BUF \mask<1>/GTS_OR  (
    .I(GTS),
    .O(\mask<1>/TORGTS )
  );
  X_BUF \mask<1>/OUTMUX_1530  (
    .I(mask_1_OBUF),
    .O(\mask<1>/OUTMUX )
  );
  X_OPAD \mask<2>/PAD  (
    .PAD(mask[2])
  );
  X_TRI mask_2_OBUF_1531 (
    .I(\mask<2>/OUTMUX ),
    .CTL(\mask<2>/ENABLE ),
    .O(mask[2])
  );
  X_INV \mask<2>/ENABLEINV  (
    .I(\mask<2>/TORGTS ),
    .O(\mask<2>/ENABLE )
  );
  X_BUF \mask<2>/GTS_OR  (
    .I(GTS),
    .O(\mask<2>/TORGTS )
  );
  X_BUF \mask<2>/OUTMUX_1532  (
    .I(mask_2_OBUF),
    .O(\mask<2>/OUTMUX )
  );
  X_ZERO \hsync/LOGIC_ZERO_1533  (
    .O(\hsync/LOGIC_ZERO )
  );
  X_OPAD \hsync/PAD  (
    .PAD(hsync)
  );
  X_TRI hsync_OBUF (
    .I(\hsync/OUTMUX ),
    .CTL(\hsync/ENABLE ),
    .O(hsync)
  );
  X_INV \hsync/ENABLEINV  (
    .I(\hsync/TORGTS ),
    .O(\hsync/ENABLE )
  );
  X_BUF \hsync/GTS_OR  (
    .I(GTS),
    .O(\hsync/TORGTS )
  );
  X_BUF \hsync/OUTMUX_1534  (
    .I(vga_top_vga1_hsyncout),
    .O(\hsync/OUTMUX )
  );
  X_IPAD \reset/PAD  (
    .PAD(reset)
  );
  X_BUF \reset/IMUX  (
    .I(\reset/IBUF ),
    .O(reset_IBUF)
  );
  X_BUF reset_IBUF_1535 (
    .I(reset),
    .O(\reset/IBUF )
  );
  X_OPAD \stall/PAD  (
    .PAD(stall)
  );
  X_TRI stall_OBUF (
    .I(\stall/OUTMUX ),
    .CTL(\stall/ENABLE ),
    .O(stall)
  );
  X_INV \stall/ENABLEINV  (
    .I(\stall/TORGTS ),
    .O(\stall/ENABLE )
  );
  X_BUF \stall/GTS_OR  (
    .I(GTS),
    .O(\stall/TORGTS )
  );
  X_BUF \stall/OUTMUX_1536  (
    .I(DLX_IDinst_stall_1),
    .O(\stall/OUTMUX )
  );
  X_BUF \stall/OMUX  (
    .I(N147786),
    .O(\stall/OD )
  );
  X_ZERO \vsync/LOGIC_ZERO_1537  (
    .O(\vsync/LOGIC_ZERO )
  );
  X_OPAD \vsync/PAD  (
    .PAD(vsync)
  );
  X_TRI vsync_OBUF (
    .I(\vsync/OUTMUX ),
    .CTL(\vsync/ENABLE ),
    .O(vsync)
  );
  X_INV \vsync/ENABLEINV  (
    .I(\vsync/TORGTS ),
    .O(\vsync/ENABLE )
  );
  X_BUF \vsync/GTS_OR  (
    .I(GTS),
    .O(\vsync/TORGTS )
  );
  X_BUF \vsync/OUTMUX_1538  (
    .I(vga_top_vga1_vsyncout),
    .O(\vsync/OUTMUX )
  );
  X_IPAD \FREEZE/PAD  (
    .PAD(FREEZE)
  );
  X_BUF \FREEZE/IMUX  (
    .I(\FREEZE/IBUF ),
    .O(FREEZE_IBUF)
  );
  X_BUF FREEZE_IBUF_1539 (
    .I(FREEZE),
    .O(\FREEZE/IBUF )
  );
  X_OPAD \branch_sig/PAD  (
    .PAD(branch_sig)
  );
  X_TRI branch_sig_OBUF (
    .I(\branch_sig/OUTMUX ),
    .CTL(\branch_sig/ENABLE ),
    .O(branch_sig)
  );
  X_INV \branch_sig/ENABLEINV  (
    .I(\branch_sig/TORGTS ),
    .O(\branch_sig/ENABLE )
  );
  X_BUF \branch_sig/GTS_OR  (
    .I(GTS),
    .O(\branch_sig/TORGTS )
  );
  X_BUF \branch_sig/OUTMUX_1540  (
    .I(DLX_IDinst_branch_sig_1),
    .O(\branch_sig/OUTMUX )
  );
  X_BUF \branch_sig/OMUX  (
    .I(N146990),
    .O(\branch_sig/OD )
  );
  X_OPAD \red<0>/PAD  (
    .PAD(red[0])
  );
  X_TRI red_0_OBUF_1541 (
    .I(\red<0>/OUTMUX ),
    .CTL(\red<0>/ENABLE ),
    .O(red[0])
  );
  X_INV \red<0>/ENABLEINV  (
    .I(\red<0>/TORGTS ),
    .O(\red<0>/ENABLE )
  );
  X_BUF \red<0>/GTS_OR  (
    .I(GTS),
    .O(\red<0>/TORGTS )
  );
  X_BUF \red<0>/OUTMUX_1542  (
    .I(red_0_OBUF),
    .O(\red<0>/OUTMUX )
  );
  X_OPAD \red<1>/PAD  (
    .PAD(red[1])
  );
  X_TRI red_1_OBUF_1543 (
    .I(\red<1>/OUTMUX ),
    .CTL(\red<1>/ENABLE ),
    .O(red[1])
  );
  X_INV \red<1>/ENABLEINV  (
    .I(\red<1>/TORGTS ),
    .O(\red<1>/ENABLE )
  );
  X_BUF \red<1>/GTS_OR  (
    .I(GTS),
    .O(\red<1>/TORGTS )
  );
  X_BUF \red<1>/OUTMUX_1544  (
    .I(red_1_OBUF),
    .O(\red<1>/OUTMUX )
  );
  X_OPAD \green<0>/PAD  (
    .PAD(green[0])
  );
  X_TRI green_0_OBUF_1545 (
    .I(\green<0>/OUTMUX ),
    .CTL(\green<0>/ENABLE ),
    .O(green[0])
  );
  X_INV \green<0>/ENABLEINV  (
    .I(\green<0>/TORGTS ),
    .O(\green<0>/ENABLE )
  );
  X_BUF \green<0>/GTS_OR  (
    .I(GTS),
    .O(\green<0>/TORGTS )
  );
  X_BUF \green<0>/OUTMUX_1546  (
    .I(green_0_OBUF),
    .O(\green<0>/OUTMUX )
  );
  X_OPAD \green<1>/PAD  (
    .PAD(green[1])
  );
  X_TRI green_1_OBUF_1547 (
    .I(\green<1>/OUTMUX ),
    .CTL(\green<1>/ENABLE ),
    .O(green[1])
  );
  X_INV \green<1>/ENABLEINV  (
    .I(\green<1>/TORGTS ),
    .O(\green<1>/ENABLE )
  );
  X_BUF \green<1>/GTS_OR  (
    .I(GTS),
    .O(\green<1>/TORGTS )
  );
  X_BUF \green<1>/OUTMUX_1548  (
    .I(green_1_OBUF),
    .O(\green<1>/OUTMUX )
  );
  X_OPAD \green<2>/PAD  (
    .PAD(green[2])
  );
  X_TRI green_2_OBUF_1549 (
    .I(\green<2>/OUTMUX ),
    .CTL(\green<2>/ENABLE ),
    .O(green[2])
  );
  X_INV \green<2>/ENABLEINV  (
    .I(\green<2>/TORGTS ),
    .O(\green<2>/ENABLE )
  );
  X_BUF \green<2>/GTS_OR  (
    .I(GTS),
    .O(\green<2>/TORGTS )
  );
  X_BUF \green<2>/OUTMUX_1550  (
    .I(green_2_OBUF),
    .O(\green<2>/OUTMUX )
  );
  X_OPAD \DM_addr_eff<10>/PAD  (
    .PAD(DM_addr_eff[10])
  );
  X_TRI DM_addr_eff_10_OBUF (
    .I(\DM_addr_eff<10>/OUTMUX ),
    .CTL(\DM_addr_eff<10>/ENABLE ),
    .O(DM_addr_eff[10])
  );
  X_INV \DM_addr_eff<10>/ENABLEINV  (
    .I(\DM_addr_eff<10>/TORGTS ),
    .O(\DM_addr_eff<10>/ENABLE )
  );
  X_BUF \DM_addr_eff<10>/GTS_OR  (
    .I(GTS),
    .O(\DM_addr_eff<10>/TORGTS )
  );
  X_BUF \DM_addr_eff<10>/OUTMUX_1551  (
    .I(DLX_EXinst_ALU_result_10_1),
    .O(\DM_addr_eff<10>/OUTMUX )
  );
  X_OPAD \DM_addr_eff<11>/PAD  (
    .PAD(DM_addr_eff[11])
  );
  X_TRI DM_addr_eff_11_OBUF (
    .I(\DM_addr_eff<11>/OUTMUX ),
    .CTL(\DM_addr_eff<11>/ENABLE ),
    .O(DM_addr_eff[11])
  );
  X_INV \DM_addr_eff<11>/ENABLEINV  (
    .I(\DM_addr_eff<11>/TORGTS ),
    .O(\DM_addr_eff<11>/ENABLE )
  );
  X_BUF \DM_addr_eff<11>/GTS_OR  (
    .I(GTS),
    .O(\DM_addr_eff<11>/TORGTS )
  );
  X_BUF \DM_addr_eff<11>/OUTMUX_1552  (
    .I(DLX_EXinst_ALU_result_11_1),
    .O(\DM_addr_eff<11>/OUTMUX )
  );
  X_OPAD \DM_addr_eff<12>/PAD  (
    .PAD(DM_addr_eff[12])
  );
  X_TRI DM_addr_eff_12_OBUF (
    .I(\DM_addr_eff<12>/OUTMUX ),
    .CTL(\DM_addr_eff<12>/ENABLE ),
    .O(DM_addr_eff[12])
  );
  X_INV \DM_addr_eff<12>/ENABLEINV  (
    .I(\DM_addr_eff<12>/TORGTS ),
    .O(\DM_addr_eff<12>/ENABLE )
  );
  X_BUF \DM_addr_eff<12>/GTS_OR  (
    .I(GTS),
    .O(\DM_addr_eff<12>/TORGTS )
  );
  X_BUF \DM_addr_eff<12>/OUTMUX_1553  (
    .I(DLX_EXinst_ALU_result_12_1),
    .O(\DM_addr_eff<12>/OUTMUX )
  );
  X_OPAD \DM_addr_eff<13>/PAD  (
    .PAD(DM_addr_eff[13])
  );
  X_TRI DM_addr_eff_13_OBUF (
    .I(\DM_addr_eff<13>/OUTMUX ),
    .CTL(\DM_addr_eff<13>/ENABLE ),
    .O(DM_addr_eff[13])
  );
  X_INV \DM_addr_eff<13>/ENABLEINV  (
    .I(\DM_addr_eff<13>/TORGTS ),
    .O(\DM_addr_eff<13>/ENABLE )
  );
  X_BUF \DM_addr_eff<13>/GTS_OR  (
    .I(GTS),
    .O(\DM_addr_eff<13>/TORGTS )
  );
  X_BUF \DM_addr_eff<13>/OUTMUX_1554  (
    .I(DLX_EXinst_ALU_result_13_1),
    .O(\DM_addr_eff<13>/OUTMUX )
  );
  defparam DLX_IDinst_RegFile_28_24_1555.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_28_24_1555 (
    .I(DLX_IDinst_WB_data_eff[24]),
    .CE(DLX_IDinst__n0606),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_28_24)
  );
  X_OPAD \DM_addr_eff<14>/PAD  (
    .PAD(DM_addr_eff[14])
  );
  X_TRI DM_addr_eff_14_OBUF (
    .I(\DM_addr_eff<14>/OUTMUX ),
    .CTL(\DM_addr_eff<14>/ENABLE ),
    .O(DM_addr_eff[14])
  );
  X_INV \DM_addr_eff<14>/ENABLEINV  (
    .I(\DM_addr_eff<14>/TORGTS ),
    .O(\DM_addr_eff<14>/ENABLE )
  );
  X_BUF \DM_addr_eff<14>/GTS_OR  (
    .I(GTS),
    .O(\DM_addr_eff<14>/TORGTS )
  );
  X_BUF \DM_addr_eff<14>/OUTMUX_1556  (
    .I(DLX_EXinst_ALU_result_14_1),
    .O(\DM_addr_eff<14>/OUTMUX )
  );
  X_OPAD \DM_addr_eff<0>/PAD  (
    .PAD(DM_addr_eff[0])
  );
  X_TRI DM_addr_eff_0_OBUF (
    .I(\DM_addr_eff<0>/OUTMUX ),
    .CTL(\DM_addr_eff<0>/ENABLE ),
    .O(DM_addr_eff[0])
  );
  X_INV \DM_addr_eff<0>/ENABLEINV  (
    .I(\DM_addr_eff<0>/TORGTS ),
    .O(\DM_addr_eff<0>/ENABLE )
  );
  X_BUF \DM_addr_eff<0>/GTS_OR  (
    .I(GTS),
    .O(\DM_addr_eff<0>/TORGTS )
  );
  X_BUF \DM_addr_eff<0>/OUTMUX_1557  (
    .I(DLX_EXinst_ALU_result_0_1),
    .O(\DM_addr_eff<0>/OUTMUX )
  );
  X_OPAD \DM_addr_eff<1>/PAD  (
    .PAD(DM_addr_eff[1])
  );
  X_TRI DM_addr_eff_1_OBUF (
    .I(\DM_addr_eff<1>/OUTMUX ),
    .CTL(\DM_addr_eff<1>/ENABLE ),
    .O(DM_addr_eff[1])
  );
  X_INV \DM_addr_eff<1>/ENABLEINV  (
    .I(\DM_addr_eff<1>/TORGTS ),
    .O(\DM_addr_eff<1>/ENABLE )
  );
  X_BUF \DM_addr_eff<1>/GTS_OR  (
    .I(GTS),
    .O(\DM_addr_eff<1>/TORGTS )
  );
  X_BUF \DM_addr_eff<1>/OUTMUX_1558  (
    .I(DLX_EXinst_ALU_result_1_1),
    .O(\DM_addr_eff<1>/OUTMUX )
  );
  X_OPAD \DM_addr_eff<2>/PAD  (
    .PAD(DM_addr_eff[2])
  );
  X_TRI DM_addr_eff_2_OBUF (
    .I(\DM_addr_eff<2>/OUTMUX ),
    .CTL(\DM_addr_eff<2>/ENABLE ),
    .O(DM_addr_eff[2])
  );
  X_INV \DM_addr_eff<2>/ENABLEINV  (
    .I(\DM_addr_eff<2>/TORGTS ),
    .O(\DM_addr_eff<2>/ENABLE )
  );
  X_BUF \DM_addr_eff<2>/GTS_OR  (
    .I(GTS),
    .O(\DM_addr_eff<2>/TORGTS )
  );
  X_BUF \DM_addr_eff<2>/OUTMUX_1559  (
    .I(DLX_EXinst_ALU_result_2_1),
    .O(\DM_addr_eff<2>/OUTMUX )
  );
  X_OPAD \DM_addr_eff<3>/PAD  (
    .PAD(DM_addr_eff[3])
  );
  X_TRI DM_addr_eff_3_OBUF (
    .I(\DM_addr_eff<3>/OUTMUX ),
    .CTL(\DM_addr_eff<3>/ENABLE ),
    .O(DM_addr_eff[3])
  );
  X_INV \DM_addr_eff<3>/ENABLEINV  (
    .I(\DM_addr_eff<3>/TORGTS ),
    .O(\DM_addr_eff<3>/ENABLE )
  );
  X_BUF \DM_addr_eff<3>/GTS_OR  (
    .I(GTS),
    .O(\DM_addr_eff<3>/TORGTS )
  );
  X_BUF \DM_addr_eff<3>/OUTMUX_1560  (
    .I(DLX_EXinst_ALU_result_3_1),
    .O(\DM_addr_eff<3>/OUTMUX )
  );
  X_OPAD \DM_addr_eff<4>/PAD  (
    .PAD(DM_addr_eff[4])
  );
  X_TRI DM_addr_eff_4_OBUF (
    .I(\DM_addr_eff<4>/OUTMUX ),
    .CTL(\DM_addr_eff<4>/ENABLE ),
    .O(DM_addr_eff[4])
  );
  X_INV \DM_addr_eff<4>/ENABLEINV  (
    .I(\DM_addr_eff<4>/TORGTS ),
    .O(\DM_addr_eff<4>/ENABLE )
  );
  X_BUF \DM_addr_eff<4>/GTS_OR  (
    .I(GTS),
    .O(\DM_addr_eff<4>/TORGTS )
  );
  X_BUF \DM_addr_eff<4>/OUTMUX_1561  (
    .I(DLX_EXinst_ALU_result_4_1),
    .O(\DM_addr_eff<4>/OUTMUX )
  );
  defparam DLX_IDinst_RegFile_28_16_1562.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_28_16_1562 (
    .I(DLX_IDinst_WB_data_eff[16]),
    .CE(DLX_IDinst__n0606),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_28_16)
  );
  X_OPAD \DM_addr_eff<5>/PAD  (
    .PAD(DM_addr_eff[5])
  );
  X_TRI DM_addr_eff_5_OBUF (
    .I(\DM_addr_eff<5>/OUTMUX ),
    .CTL(\DM_addr_eff<5>/ENABLE ),
    .O(DM_addr_eff[5])
  );
  X_INV \DM_addr_eff<5>/ENABLEINV  (
    .I(\DM_addr_eff<5>/TORGTS ),
    .O(\DM_addr_eff<5>/ENABLE )
  );
  X_BUF \DM_addr_eff<5>/GTS_OR  (
    .I(GTS),
    .O(\DM_addr_eff<5>/TORGTS )
  );
  X_BUF \DM_addr_eff<5>/OUTMUX_1563  (
    .I(DLX_EXinst_ALU_result_5_1),
    .O(\DM_addr_eff<5>/OUTMUX )
  );
  X_OPAD \DM_addr_eff<6>/PAD  (
    .PAD(DM_addr_eff[6])
  );
  X_TRI DM_addr_eff_6_OBUF (
    .I(\DM_addr_eff<6>/OUTMUX ),
    .CTL(\DM_addr_eff<6>/ENABLE ),
    .O(DM_addr_eff[6])
  );
  X_INV \DM_addr_eff<6>/ENABLEINV  (
    .I(\DM_addr_eff<6>/TORGTS ),
    .O(\DM_addr_eff<6>/ENABLE )
  );
  X_BUF \DM_addr_eff<6>/GTS_OR  (
    .I(GTS),
    .O(\DM_addr_eff<6>/TORGTS )
  );
  X_BUF \DM_addr_eff<6>/OUTMUX_1564  (
    .I(DLX_EXinst_ALU_result_6_1),
    .O(\DM_addr_eff<6>/OUTMUX )
  );
  X_OPAD \DM_addr_eff<7>/PAD  (
    .PAD(DM_addr_eff[7])
  );
  X_TRI DM_addr_eff_7_OBUF (
    .I(\DM_addr_eff<7>/OUTMUX ),
    .CTL(\DM_addr_eff<7>/ENABLE ),
    .O(DM_addr_eff[7])
  );
  X_INV \DM_addr_eff<7>/ENABLEINV  (
    .I(\DM_addr_eff<7>/TORGTS ),
    .O(\DM_addr_eff<7>/ENABLE )
  );
  X_BUF \DM_addr_eff<7>/GTS_OR  (
    .I(GTS),
    .O(\DM_addr_eff<7>/TORGTS )
  );
  X_BUF \DM_addr_eff<7>/OUTMUX_1565  (
    .I(DLX_EXinst_ALU_result_7_1),
    .O(\DM_addr_eff<7>/OUTMUX )
  );
  X_OPAD \DM_addr_eff<8>/PAD  (
    .PAD(DM_addr_eff[8])
  );
  X_TRI DM_addr_eff_8_OBUF (
    .I(\DM_addr_eff<8>/OUTMUX ),
    .CTL(\DM_addr_eff<8>/ENABLE ),
    .O(DM_addr_eff[8])
  );
  X_INV \DM_addr_eff<8>/ENABLEINV  (
    .I(\DM_addr_eff<8>/TORGTS ),
    .O(\DM_addr_eff<8>/ENABLE )
  );
  X_BUF \DM_addr_eff<8>/GTS_OR  (
    .I(GTS),
    .O(\DM_addr_eff<8>/TORGTS )
  );
  X_BUF \DM_addr_eff<8>/OUTMUX_1566  (
    .I(DLX_EXinst_ALU_result_8_1),
    .O(\DM_addr_eff<8>/OUTMUX )
  );
  X_OPAD \DM_addr_eff<9>/PAD  (
    .PAD(DM_addr_eff[9])
  );
  X_TRI DM_addr_eff_9_OBUF (
    .I(\DM_addr_eff<9>/OUTMUX ),
    .CTL(\DM_addr_eff<9>/ENABLE ),
    .O(DM_addr_eff[9])
  );
  X_INV \DM_addr_eff<9>/ENABLEINV  (
    .I(\DM_addr_eff<9>/TORGTS ),
    .O(\DM_addr_eff<9>/ENABLE )
  );
  X_BUF \DM_addr_eff<9>/GTS_OR  (
    .I(GTS),
    .O(\DM_addr_eff<9>/TORGTS )
  );
  X_BUF \DM_addr_eff<9>/OUTMUX_1567  (
    .I(DLX_EXinst_ALU_result_9_1),
    .O(\DM_addr_eff<9>/OUTMUX )
  );
  X_OPAD \PIPEEMPTY/PAD  (
    .PAD(PIPEEMPTY)
  );
  X_TRI PIPEEMPTY_OBUF_1568 (
    .I(\PIPEEMPTY/OUTMUX ),
    .CTL(\PIPEEMPTY/ENABLE ),
    .O(PIPEEMPTY)
  );
  X_INV \PIPEEMPTY/ENABLEINV  (
    .I(\PIPEEMPTY/TORGTS ),
    .O(\PIPEEMPTY/ENABLE )
  );
  X_BUF \PIPEEMPTY/GTS_OR  (
    .I(GTS),
    .O(\PIPEEMPTY/TORGTS )
  );
  X_BUF \PIPEEMPTY/OUTMUX_1569  (
    .I(PIPEEMPTY_OBUF),
    .O(\PIPEEMPTY/OUTMUX )
  );
  X_OPAD \DM_read/PAD  (
    .PAD(DM_read)
  );
  X_TRI DM_read_OBUF (
    .I(\DM_read/OUTMUX ),
    .CTL(\DM_read/ENABLE ),
    .O(DM_read)
  );
  X_INV \DM_read/ENABLEINV  (
    .I(\DM_read/TORGTS ),
    .O(\DM_read/ENABLE )
  );
  X_BUF \DM_read/GTS_OR  (
    .I(GTS),
    .O(\DM_read/TORGTS )
  );
  X_BUF \DM_read/OUTMUX_1570  (
    .I(DLX_EXinst_mem_read_EX),
    .O(\DM_read/OUTMUX )
  );
  X_BUF \DM_read/OMUX  (
    .I(DLX_IDinst_mem_read),
    .O(\DM_read/OD )
  );
  X_OPAD \IR_MSB<0>/PAD  (
    .PAD(IR_MSB[0])
  );
  X_TRI IR_MSB_0_OBUF_1571 (
    .I(\IR_MSB<0>/OUTMUX ),
    .CTL(\IR_MSB<0>/ENABLE ),
    .O(IR_MSB[0])
  );
  X_INV \IR_MSB<0>/ENABLEINV  (
    .I(\IR_MSB<0>/TORGTS ),
    .O(\IR_MSB<0>/ENABLE )
  );
  X_BUF \IR_MSB<0>/GTS_OR  (
    .I(GTS),
    .O(\IR_MSB<0>/TORGTS )
  );
  X_BUF \IR_MSB<0>/OUTMUX_1572  (
    .I(IR_MSB_0_OBUF),
    .O(\IR_MSB<0>/OUTMUX )
  );
  X_OPAD \IR_MSB<1>/PAD  (
    .PAD(IR_MSB[1])
  );
  X_TRI IR_MSB_1_OBUF_1573 (
    .I(\IR_MSB<1>/OUTMUX ),
    .CTL(\IR_MSB<1>/ENABLE ),
    .O(IR_MSB[1])
  );
  X_INV \IR_MSB<1>/ENABLEINV  (
    .I(\IR_MSB<1>/TORGTS ),
    .O(\IR_MSB<1>/ENABLE )
  );
  X_BUF \IR_MSB<1>/GTS_OR  (
    .I(GTS),
    .O(\IR_MSB<1>/TORGTS )
  );
  X_BUF \IR_MSB<1>/OUTMUX_1574  (
    .I(IR_MSB_1_OBUF),
    .O(\IR_MSB<1>/OUTMUX )
  );
  X_OPAD \IR_MSB<2>/PAD  (
    .PAD(IR_MSB[2])
  );
  X_TRI IR_MSB_2_OBUF_1575 (
    .I(\IR_MSB<2>/OUTMUX ),
    .CTL(\IR_MSB<2>/ENABLE ),
    .O(IR_MSB[2])
  );
  X_INV \IR_MSB<2>/ENABLEINV  (
    .I(\IR_MSB<2>/TORGTS ),
    .O(\IR_MSB<2>/ENABLE )
  );
  X_BUF \IR_MSB<2>/GTS_OR  (
    .I(GTS),
    .O(\IR_MSB<2>/TORGTS )
  );
  X_BUF \IR_MSB<2>/OUTMUX_1576  (
    .I(IR_MSB_2_OBUF),
    .O(\IR_MSB<2>/OUTMUX )
  );
  X_OPAD \IR_MSB<3>/PAD  (
    .PAD(IR_MSB[3])
  );
  X_TRI IR_MSB_3_OBUF_1577 (
    .I(\IR_MSB<3>/OUTMUX ),
    .CTL(\IR_MSB<3>/ENABLE ),
    .O(IR_MSB[3])
  );
  X_INV \IR_MSB<3>/ENABLEINV  (
    .I(\IR_MSB<3>/TORGTS ),
    .O(\IR_MSB<3>/ENABLE )
  );
  X_BUF \IR_MSB<3>/GTS_OR  (
    .I(GTS),
    .O(\IR_MSB<3>/TORGTS )
  );
  X_BUF \IR_MSB<3>/OUTMUX_1578  (
    .I(IR_MSB_3_OBUF),
    .O(\IR_MSB<3>/OUTMUX )
  );
  X_OPAD \IR_MSB<4>/PAD  (
    .PAD(IR_MSB[4])
  );
  X_TRI IR_MSB_4_OBUF_1579 (
    .I(\IR_MSB<4>/OUTMUX ),
    .CTL(\IR_MSB<4>/ENABLE ),
    .O(IR_MSB[4])
  );
  X_INV \IR_MSB<4>/ENABLEINV  (
    .I(\IR_MSB<4>/TORGTS ),
    .O(\IR_MSB<4>/ENABLE )
  );
  X_BUF \IR_MSB<4>/GTS_OR  (
    .I(GTS),
    .O(\IR_MSB<4>/TORGTS )
  );
  X_BUF \IR_MSB<4>/OUTMUX_1580  (
    .I(IR_MSB_4_OBUF),
    .O(\IR_MSB<4>/OUTMUX )
  );
  X_OPAD \IR_MSB<5>/PAD  (
    .PAD(IR_MSB[5])
  );
  X_TRI IR_MSB_5_OBUF_1581 (
    .I(\IR_MSB<5>/OUTMUX ),
    .CTL(\IR_MSB<5>/ENABLE ),
    .O(IR_MSB[5])
  );
  X_INV \IR_MSB<5>/ENABLEINV  (
    .I(\IR_MSB<5>/TORGTS ),
    .O(\IR_MSB<5>/ENABLE )
  );
  X_BUF \IR_MSB<5>/GTS_OR  (
    .I(GTS),
    .O(\IR_MSB<5>/TORGTS )
  );
  X_BUF \IR_MSB<5>/OUTMUX_1582  (
    .I(IR_MSB_5_OBUF),
    .O(\IR_MSB<5>/OUTMUX )
  );
  X_OPAD \IR_MSB<6>/PAD  (
    .PAD(IR_MSB[6])
  );
  X_TRI IR_MSB_6_OBUF_1583 (
    .I(\IR_MSB<6>/OUTMUX ),
    .CTL(\IR_MSB<6>/ENABLE ),
    .O(IR_MSB[6])
  );
  X_INV \IR_MSB<6>/ENABLEINV  (
    .I(\IR_MSB<6>/TORGTS ),
    .O(\IR_MSB<6>/ENABLE )
  );
  X_BUF \IR_MSB<6>/GTS_OR  (
    .I(GTS),
    .O(\IR_MSB<6>/TORGTS )
  );
  X_BUF \IR_MSB<6>/OUTMUX_1584  (
    .I(IR_MSB_6_OBUF),
    .O(\IR_MSB<6>/OUTMUX )
  );
  X_OPAD \IR_MSB<7>/PAD  (
    .PAD(IR_MSB[7])
  );
  X_TRI IR_MSB_7_OBUF_1585 (
    .I(\IR_MSB<7>/OUTMUX ),
    .CTL(\IR_MSB<7>/ENABLE ),
    .O(IR_MSB[7])
  );
  X_INV \IR_MSB<7>/ENABLEINV  (
    .I(\IR_MSB<7>/TORGTS ),
    .O(\IR_MSB<7>/ENABLE )
  );
  X_BUF \IR_MSB<7>/GTS_OR  (
    .I(GTS),
    .O(\IR_MSB<7>/TORGTS )
  );
  X_BUF \IR_MSB<7>/OUTMUX_1586  (
    .I(IR_MSB_7_OBUF),
    .O(\IR_MSB<7>/OUTMUX )
  );
  X_ZERO \clkdivider/LOGIC_ZERO_1587  (
    .O(\clkdivider/LOGIC_ZERO )
  );
  defparam clkdivider.CLKDV_DIVIDE = 2.0;
  defparam clkdivider.DUTY_CYCLE_CORRECTION = "TRUE";
  defparam clkdivider.MAXPERCLKIN = 40000;
  X_CLKDLLE clkdivider (
    .CLKIN(\clk/new_buffer ),
    .CLKFB(clk0buf),
    .RST(\clkdivider/LOGIC_ZERO ),
    .CLK0(clk0),
    .CLK90(\clkdivider/CLK90 ),
    .CLK180(\clkdivider/CLK180 ),
    .CLK270(\clkdivider/CLK270 ),
    .CLK2X(\clkdivider/CLK2X ),
    .CLK2X180(\clkdivider/CLK2X180 ),
    .CLKDV(clkdivub),
    .LOCKED(\clkdivider/LOCKED )
  );
  X_ZERO \vga0/LOGIC_ZERO_1588  (
    .O(\vga0/LOGIC_ZERO )
  );
  X_ONE \vga0/LOGIC_ONE_1589  (
    .O(\vga0/LOGIC_ONE )
  );
  X_INV \vga0/CLKAMUX  (
    .I(clkdiv),
    .O(\vga0/CLKA_INTNOT )
  );
  defparam vga0.INIT_00 = 256'h000000000000000000001CE080F000008003FF00000000000000000000007F00;
  defparam vga0.INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga0.INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga0.INIT_03 = 256'h0000000000000000000000000000000000000000000000000000007000000000;
  defparam vga0.INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga0.INIT_05 = 256'h0000000000000000000000380000000000000000000000000000000000000070;
  defparam vga0.INIT_06 = 256'h0000E06000000000000000000000000000000000000000300000000000000000;
  defparam vga0.INIT_07 = 256'h00000000000001C000000000186060600000000000000000000001C000000000;
  defparam vga0.INIT_08 = 256'h00000000000080208000000000000000000000C0000000000000C02000000000;
  defparam vga0.INIT_09 = 256'h8000000000000000000000C000000000000080208000000000000000000000C0;
  defparam vga0.INIT_0A = 256'h000000C000000000000080208000000000000000000000800000000000008000;
  defparam vga0.INIT_0B = 256'h0000800080000000000000000000008000000000000080008000000000000000;
  defparam vga0.INIT_0C = 256'h0000000000000080000000000000800000000000000000000000008000000000;
  defparam vga0.INIT_0D = 256'h00000000000080008000000000000000000000C0000000000000802080000000;
  defparam vga0.INIT_0E = 256'h0000000000000008000000400000300000000000800000000000000000000080;
  defparam vga0.INIT_0F = 256'h0000003000001800000000000000000000000004000000600000300000000000;
  defparam vga0.SETUP_ALL = 2701;
  X_RAMB4_S1_S1 vga0 (
    .CLKA(\vga0/CLKA_INTNOT ),
    .CLKB(clkdiv),
    .ENA(Mshift__n0000_Sh[33]),
    .ENB(\vga0/LOGIC_ONE ),
    .RSTA(reset_IBUF_1),
    .RSTB(reset_IBUF_1),
    .WEA(DLX_EXinst_mem_write_EX),
    .WEB(\vga0/LOGIC_ZERO ),
    .GSR(GSR),
    .ADDRA({DLX_EXinst_ALU_result[11], DLX_EXinst_ALU_result[10], DLX_EXinst_ALU_result[9], DLX_EXinst_ALU_result[8], DLX_EXinst_ALU_result[7], 
DLX_EXinst_ALU_result[6], DLX_EXinst_ALU_result[5], DLX_EXinst_ALU_result[4], DLX_EXinst_ALU_result[3], DLX_EXinst_ALU_result[2], 
DLX_EXinst_ALU_result[1], DLX_EXinst_ALU_result[0]}),
    .ADDRB({vga_address[11], vga_address[10], vga_address[9], vga_address[8], vga_address[7], vga_address[6], 
vga_top_vga1_Madd_addressout_inst_lut2_331, vga_top_vga1_gridhcounter[4], vga_top_vga1_gridhcounter[3], vga_top_vga1_gridhcounter[2], 
vga_top_vga1_gridhcounter[1], vga_top_vga1_gridhcounter[0]}),
    .DIA({DLX_EXinst_reg_out_B_EX[0]}),
    .DIB({\vga0/DIB0 }),
    .DOA({vram_out_cpu[0]}),
    .DOB({vram_out_vga[0]})
  );
  X_ZERO \vga1/LOGIC_ZERO_1590  (
    .O(\vga1/LOGIC_ZERO )
  );
  X_ONE \vga1/LOGIC_ONE_1591  (
    .O(\vga1/LOGIC_ONE )
  );
  X_INV \vga1/CLKAMUX  (
    .I(clkdiv),
    .O(\vga1/CLKA_INTNOT )
  );
  defparam vga1.INIT_00 = 256'h000000010000000001400000000000300000180000000000000000000180001C;
  defparam vga1.INIT_01 = 256'h0000000000000018000010000000000100000000010000000000001800401000;
  defparam vga1.INIT_02 = 256'h0040100000000011000000000000000000000018004010000000000100000000;
  defparam vga1.INIT_03 = 256'h0000000000000000000000180040000000000001000000000000000000000008;
  defparam vga1.INIT_04 = 256'h0000000800000000000000000000000000000000000000180040000000000000;
  defparam vga1.INIT_05 = 256'h00000000C0000000C00000000000001000000000000000000000000000000000;
  defparam vga1.INIT_06 = 256'h00000000000000100000000000000000C0000000000000000000001000000000;
  defparam vga1.INIT_07 = 256'h0000000000000000C000000000000000000000000000000000000000C0000000;
  defparam vga1.INIT_08 = 256'h0000000000000000038000000000000000000000C00000000000000000000000;
  defparam vga1.INIT_09 = 256'h0380000000000000000000000000000000000000038000000000000000000000;
  defparam vga1.INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga1.INIT_0B = 256'h00000000C000000000000000000000000000000000000000C000000000000000;
  defparam vga1.INIT_0C = 256'h00000000000000000000000000000000C0000000000000000000000000000000;
  defparam vga1.INIT_0D = 256'h00000000000000000000000000000000000000000000000000000000C0000000;
  defparam vga1.INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga1.INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga1.SETUP_ALL = 2701;
  X_RAMB4_S1_S1 vga1 (
    .CLKA(\vga1/CLKA_INTNOT ),
    .CLKB(clkdiv),
    .ENA(Mshift__n0000_Sh[34]),
    .ENB(\vga1/LOGIC_ONE ),
    .RSTA(reset_IBUF_1),
    .RSTB(reset_IBUF_1),
    .WEA(DLX_EXinst_mem_write_EX),
    .WEB(\vga1/LOGIC_ZERO ),
    .GSR(GSR),
    .ADDRA({DLX_EXinst_ALU_result[11], DLX_EXinst_ALU_result[10], DLX_EXinst_ALU_result[9], DLX_EXinst_ALU_result[8], DLX_EXinst_ALU_result[7], 
DLX_EXinst_ALU_result[6], DLX_EXinst_ALU_result[5], DLX_EXinst_ALU_result[4], DLX_EXinst_ALU_result[3], DLX_EXinst_ALU_result[2], 
DLX_EXinst_ALU_result[1], DLX_EXinst_ALU_result[0]}),
    .ADDRB({vga_address[11], vga_address[10], vga_address[9], vga_address[8], vga_address[7], vga_address[6], 
vga_top_vga1_Madd_addressout_inst_lut2_331, vga_top_vga1_gridhcounter[4], vga_top_vga1_gridhcounter[3], vga_top_vga1_gridhcounter[2], 
vga_top_vga1_gridhcounter[1], vga_top_vga1_gridhcounter[0]}),
    .DIA({DLX_EXinst_reg_out_B_EX[0]}),
    .DIB({\vga1/DIB0 }),
    .DOA({vram_out_cpu[1]}),
    .DOB({vram_out_vga[1]})
  );
  X_ZERO \vga2/LOGIC_ZERO_1592  (
    .O(\vga2/LOGIC_ZERO )
  );
  X_ONE \vga2/LOGIC_ONE_1593  (
    .O(\vga2/LOGIC_ONE )
  );
  X_INV \vga2/CLKAMUX  (
    .I(clkdiv),
    .O(\vga2/CLKA_INTNOT )
  );
  defparam vga2.INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga2.INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga2.INIT_02 = 256'h0000000000000000000000000000001C00000000800000008000000000000000;
  defparam vga2.INIT_03 = 256'h000000000000001C000000000000000000000000000000000000001C00000000;
  defparam vga2.INIT_04 = 256'h0000000080000000800000000000000000000000000000000000000000000000;
  defparam vga2.INIT_05 = 256'h8000000000000000000000000000000080000000800000000000000000000000;
  defparam vga2.INIT_06 = 256'h0000000000000000800000008000000000000000000000000000000080000000;
  defparam vga2.INIT_07 = 256'h0000000000000000000000000000000000000000800000000000000000000000;
  defparam vga2.INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga2.INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga2.INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga2.INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga2.INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga2.INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga2.INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga2.INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga2.SETUP_ALL = 2701;
  X_RAMB4_S1_S1 vga2 (
    .CLKA(\vga2/CLKA_INTNOT ),
    .CLKB(clkdiv),
    .ENA(Mshift__n0000_Sh[35]),
    .ENB(\vga2/LOGIC_ONE ),
    .RSTA(reset_IBUF_1),
    .RSTB(reset_IBUF_1),
    .WEA(DLX_EXinst_mem_write_EX),
    .WEB(\vga2/LOGIC_ZERO ),
    .GSR(GSR),
    .ADDRA({DLX_EXinst_ALU_result[11], DLX_EXinst_ALU_result[10], DLX_EXinst_ALU_result[9], DLX_EXinst_ALU_result[8], DLX_EXinst_ALU_result[7], 
DLX_EXinst_ALU_result[6], DLX_EXinst_ALU_result[5], DLX_EXinst_ALU_result[4], DLX_EXinst_ALU_result[3], DLX_EXinst_ALU_result[2], 
DLX_EXinst_ALU_result[1], DLX_EXinst_ALU_result[0]}),
    .ADDRB({vga_address[11], vga_address[10], vga_address[9], vga_address[8], vga_address[7], vga_address[6], 
vga_top_vga1_Madd_addressout_inst_lut2_331, vga_top_vga1_gridhcounter[4], vga_top_vga1_gridhcounter[3], vga_top_vga1_gridhcounter[2], 
vga_top_vga1_gridhcounter[1], vga_top_vga1_gridhcounter[0]}),
    .DIA({DLX_EXinst_reg_out_B_EX[0]}),
    .DIB({\vga2/DIB0 }),
    .DOA({vram_out_cpu[2]}),
    .DOB({vram_out_vga[2]})
  );
  X_ZERO \vga3/LOGIC_ZERO_1594  (
    .O(\vga3/LOGIC_ZERO )
  );
  X_ONE \vga3/LOGIC_ONE_1595  (
    .O(\vga3/LOGIC_ONE )
  );
  X_INV \vga3/CLKAMUX  (
    .I(clkdiv),
    .O(\vga3/CLKA_INTNOT )
  );
  defparam vga3.INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga3.INIT_01 = 256'h0000000000000000000000000000000000000400000000000000000000000000;
  defparam vga3.INIT_02 = 256'h0000000000000000000012000000000000000000000000000000000000000C00;
  defparam vga3.INIT_03 = 256'h0000000000000000000000000000000000001800000000000000000000000000;
  defparam vga3.INIT_04 = 256'h0000000000000000000008000000000000003FF0000000000000000000000800;
  defparam vga3.INIT_05 = 256'h0000038000000000000000000000000000000000000000000000000000000000;
  defparam vga3.INIT_06 = 256'h0000000000000000000000000000008000000000000000000000000000000000;
  defparam vga3.INIT_07 = 256'h01C000000000000000000000000000000000000000000000010000000003FF00;
  defparam vga3.INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga3.INIT_09 = 256'h0000E00000000000000000000000000000000000000080000000000000000000;
  defparam vga3.INIT_0A = 256'h0000000000000000000000000000004000000000000000000000000000000000;
  defparam vga3.INIT_0B = 256'h00000000000001F000000000000000000000000000000000000000E000000000;
  defparam vga3.INIT_0C = 256'h00000000000000000000000000000000000003F8000000000000000000000000;
  defparam vga3.INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga3.INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga3.INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga3.SETUP_ALL = 2701;
  X_RAMB4_S1_S1 vga3 (
    .CLKA(\vga3/CLKA_INTNOT ),
    .CLKB(clkdiv),
    .ENA(Mshift__n0000_Sh[36]),
    .ENB(\vga3/LOGIC_ONE ),
    .RSTA(reset_IBUF_1),
    .RSTB(reset_IBUF_1),
    .WEA(DLX_EXinst_mem_write_EX),
    .WEB(\vga3/LOGIC_ZERO ),
    .GSR(GSR),
    .ADDRA({DLX_EXinst_ALU_result[11], DLX_EXinst_ALU_result[10], DLX_EXinst_ALU_result[9], DLX_EXinst_ALU_result[8], DLX_EXinst_ALU_result[7], 
DLX_EXinst_ALU_result[6], DLX_EXinst_ALU_result[5], DLX_EXinst_ALU_result[4], DLX_EXinst_ALU_result[3], DLX_EXinst_ALU_result[2], 
DLX_EXinst_ALU_result[1], DLX_EXinst_ALU_result[0]}),
    .ADDRB({vga_address[11], vga_address[10], vga_address[9], vga_address[8], vga_address[7], vga_address[6], 
vga_top_vga1_Madd_addressout_inst_lut2_331, vga_top_vga1_gridhcounter[4], vga_top_vga1_gridhcounter[3], vga_top_vga1_gridhcounter[2], 
vga_top_vga1_gridhcounter[1], vga_top_vga1_gridhcounter[0]}),
    .DIA({DLX_EXinst_reg_out_B_EX[0]}),
    .DIB({\vga3/DIB0 }),
    .DOA({vram_out_cpu[3]}),
    .DOB({vram_out_vga[3]})
  );
  X_ZERO \vga4/LOGIC_ZERO_1596  (
    .O(\vga4/LOGIC_ZERO )
  );
  X_ONE \vga4/LOGIC_ONE_1597  (
    .O(\vga4/LOGIC_ONE )
  );
  X_INV \vga4/CLKAMUX  (
    .I(clkdiv),
    .O(\vga4/CLKA_INTNOT )
  );
  defparam vga4.INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga4.INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga4.INIT_02 = 256'h00000000000000000003E000000000000000000000000000000000000003E000;
  defparam vga4.INIT_03 = 256'h0003E000000000000000000000000000000000000003E0000000000000000000;
  defparam vga4.INIT_04 = 256'h0000000000000000000000000003E00000000000000000000000000000000000;
  defparam vga4.INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga4.INIT_06 = 256'h0000000000000000006000000000000000700000000000000000000000C00000;
  defparam vga4.INIT_07 = 256'h000C00000000000000100000001E000000000000003000000000000000700000;
  defparam vga4.INIT_08 = 256'h0000000000000000000000000006000000000000000000000000000000000000;
  defparam vga4.INIT_09 = 256'h0000000000060000000000000000000000000000000000000006000000000000;
  defparam vga4.INIT_0A = 256'h00000000000000000000000000000000000600F0000000000000000000000000;
  defparam vga4.INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga4.INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga4.INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga4.INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga4.INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam vga4.SETUP_ALL = 2701;
  X_RAMB4_S1_S1 vga4 (
    .CLKA(\vga4/CLKA_INTNOT ),
    .CLKB(clkdiv),
    .ENA(Mshift__n0000_Sh[37]),
    .ENB(\vga4/LOGIC_ONE ),
    .RSTA(reset_IBUF_1),
    .RSTB(reset_IBUF_1),
    .WEA(DLX_EXinst_mem_write_EX),
    .WEB(\vga4/LOGIC_ZERO ),
    .GSR(GSR),
    .ADDRA({DLX_EXinst_ALU_result[11], DLX_EXinst_ALU_result[10], DLX_EXinst_ALU_result[9], DLX_EXinst_ALU_result[8], DLX_EXinst_ALU_result[7], 
DLX_EXinst_ALU_result[6], DLX_EXinst_ALU_result[5], DLX_EXinst_ALU_result[4], DLX_EXinst_ALU_result[3], DLX_EXinst_ALU_result[2], 
DLX_EXinst_ALU_result[1], DLX_EXinst_ALU_result[0]}),
    .ADDRB({vga_address[11], vga_address[10], vga_address[9], vga_address[8], vga_address[7], vga_address[6], 
vga_top_vga1_Madd_addressout_inst_lut2_331, vga_top_vga1_gridhcounter[4], vga_top_vga1_gridhcounter[3], vga_top_vga1_gridhcounter[2], 
vga_top_vga1_gridhcounter[1], vga_top_vga1_gridhcounter[0]}),
    .DIA({DLX_EXinst_reg_out_B_EX[0]}),
    .DIB({\vga4/DIB0 }),
    .DOA({vram_out_cpu[4]}),
    .DOB({vram_out_vga[4]})
  );
  X_ONE \block0/LOGIC_ONE_1598  (
    .O(\block0/LOGIC_ONE )
  );
  X_ZERO \block0/LOGIC_ZERO_1599  (
    .O(\block0/LOGIC_ZERO )
  );
  X_INV \block0/CLKAMUX  (
    .I(clkdiv),
    .O(\block0/CLKA_INTNOT )
  );
  defparam block0.INIT_00 = 256'h0000000000000000000000000000000000000000000000000000E80000000000;
  defparam block0.INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block0.INIT_02 = 256'hD0140001A000E8000001A00000280020203C00F4000000F00100200000E80000;
  defparam block0.INIT_03 = 256'h0205A02000003C001020280000244440A0000000C47801A000B4005CA0000000;
  defparam block0.INIT_04 = 256'h0028004C2020A0100C080400000000B401010021212101000820240006001F21;
  defparam block0.INIT_05 = 256'h008461FF603F9FA0A101002C0090202000002000C0010100250006001F200205;
  defparam block0.INIT_06 = 256'h019FA001002C009077002861605FA1A09F01010050019FC16061A09F01002C9F;
  defparam block0.INIT_07 = 256'hA0002C00905F606101019FA0A100B8FF6061773F01A0A1002C9F00EC5F60C19F;
  defparam block0.INIT_08 = 256'h0004A1A09F01019FA0A1002C013F9FA09F01A0A1002C9F00603F9F01A1A0019F;
  defparam block0.INIT_09 = 256'h0008000100080001000800010008000100080001000800010008000100080020;
  defparam block0.INIT_0A = 256'h0000000000EC0401001405200000010008202404010020010008200300200001;
  defparam block0.INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block0.INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block0.INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block0.INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block0.INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block0.SETUP_ALL = 2701;
  X_RAMB4_S8_S8 block0 (
    .CLKA(\block0/CLKA_INTNOT ),
    .CLKB(clkdiv),
    .ENA(mask_0_OBUF),
    .ENB(\block0/LOGIC_ONE ),
    .RSTA(\block0/LOGIC_ZERO ),
    .RSTB(\block0/LOGIC_ZERO ),
    .WEA(DLX_EXinst_mem_write_EX),
    .WEB(\block0/LOGIC_ZERO ),
    .GSR(GSR),
    .ADDRA({DLX_EXinst_ALU_result[10], DLX_EXinst_ALU_result[9], DLX_EXinst_ALU_result[8], DLX_EXinst_ALU_result[7], DLX_EXinst_ALU_result[6], 
DLX_EXinst_ALU_result[5], DLX_EXinst_ALU_result[4], DLX_EXinst_ALU_result[3], DLX_EXinst_ALU_result[2]}),
    .ADDRB({DLX_IFinst_NPC[10], DLX_IFinst_NPC[9], DLX_IFinst_NPC[8], DLX_IFinst_NPC[7], DLX_IFinst_NPC[6], DLX_IFinst_NPC[5], DLX_IFinst_NPC[4], 
DLX_IFinst_NPC[3], DLX_IFinst_NPC[2]}),
    .DIA({DLX_EXinst_reg_out_B_EX[7], DLX_EXinst_reg_out_B_EX[6], DLX_EXinst_reg_out_B_EX[5], DLX_EXinst_reg_out_B_EX[4], DLX_EXinst_reg_out_B_EX[3], 
DLX_EXinst_reg_out_B_EX[2], DLX_EXinst_reg_out_B_EX[1], DLX_EXinst_reg_out_B_EX[0]}),
    .DIB({\block0/DIB7 , \block0/DIB6 , \block0/DIB5 , \block0/DIB4 , \block0/DIB3 , \block0/DIB2 , \block0/DIB1 , \block0/DIB0 }),
    .DOA({RAM_read_data[7], RAM_read_data[6], RAM_read_data[5], RAM_read_data[4], RAM_read_data[3], RAM_read_data[2], RAM_read_data[1], 
RAM_read_data[0]}),
    .DOB({IR[7], IR[6], IR[5], IR[4], IR[3], IR[2], IR[1], IR[0]})
  );
  X_ONE \block1/LOGIC_ONE_1600  (
    .O(\block1/LOGIC_ONE )
  );
  X_ZERO \block1/LOGIC_ZERO_1601  (
    .O(\block1/LOGIC_ZERO )
  );
  X_INV \block1/CLKAMUX  (
    .I(clkdiv),
    .O(\block1/CLKA_INTNOT )
  );
  defparam block1.INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block1.INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block1.INIT_02 = 256'h00080000000000080000000001080088800800FF000000FF0000000000031000;
  defparam block1.INIT_03 = 256'h000000B80000080000C008000000080800080000FF0000000003000000080000;
  defparam block1.INIT_04 = 256'h000000006068000000000000000000FF000000A0A0A0000000A89800A08000B0;
  defparam block1.INIT_05 = 256'h00014A4A4A010000000000000000D0D00000F800FF000000B000B88000C80000;
  defparam block1.INIT_06 = 256'h00000000000000000000014A4A4A000000000000010000494A4A000000000000;
  defparam block1.INIT_07 = 256'h00000000004A4A4A000000000000004A4A4A000100000000000000004A4A4900;
  defparam block1.INIT_08 = 256'h0000000000000000000000000001000000000000000000000001000000000000;
  defparam block1.INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000040;
  defparam block1.INIT_0A = 256'h0000000000FF0000080800C8000000000008A000000000000000080000000000;
  defparam block1.INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block1.INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block1.INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block1.INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block1.INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block1.SETUP_ALL = 2701;
  X_RAMB4_S8_S8 block1 (
    .CLKA(\block1/CLKA_INTNOT ),
    .CLKB(clkdiv),
    .ENA(mask_1_OBUF),
    .ENB(\block1/LOGIC_ONE ),
    .RSTA(\block1/LOGIC_ZERO ),
    .RSTB(\block1/LOGIC_ZERO ),
    .WEA(DLX_EXinst_mem_write_EX),
    .WEB(\block1/LOGIC_ZERO ),
    .GSR(GSR),
    .ADDRA({DLX_EXinst_ALU_result[10], DLX_EXinst_ALU_result[9], DLX_EXinst_ALU_result[8], DLX_EXinst_ALU_result[7], DLX_EXinst_ALU_result[6], 
DLX_EXinst_ALU_result[5], DLX_EXinst_ALU_result[4], DLX_EXinst_ALU_result[3], DLX_EXinst_ALU_result[2]}),
    .ADDRB({DLX_IFinst_NPC[10], DLX_IFinst_NPC[9], DLX_IFinst_NPC[8], DLX_IFinst_NPC[7], DLX_IFinst_NPC[6], DLX_IFinst_NPC[5], DLX_IFinst_NPC[4], 
DLX_IFinst_NPC[3], DLX_IFinst_NPC[2]}),
    .DIA({DLX_EXinst_reg_out_B_EX[15], DLX_EXinst_reg_out_B_EX[14], DLX_EXinst_reg_out_B_EX[13], DLX_EXinst_reg_out_B_EX[12], 
DLX_EXinst_reg_out_B_EX[11], DLX_EXinst_reg_out_B_EX[10], DLX_EXinst_reg_out_B_EX[9], DLX_EXinst_reg_out_B_EX[8]}),
    .DIB({\block1/DIB7 , \block1/DIB6 , \block1/DIB5 , \block1/DIB4 , \block1/DIB3 , \block1/DIB2 , \block1/DIB1 , \block1/DIB0 }),
    .DOA({RAM_read_data[15], RAM_read_data[14], RAM_read_data[13], RAM_read_data[12], RAM_read_data[11], RAM_read_data[10], RAM_read_data[9], 
RAM_read_data[8]}),
    .DOB({IR[15], IR[14], IR[13], IR[12], IR[11], IR[10], IR[9], IR[8]})
  );
  X_ONE \block2/LOGIC_ONE_1602  (
    .O(\block2/LOGIC_ONE )
  );
  X_ZERO \block2/LOGIC_ZERO_1603  (
    .O(\block2/LOGIC_ZERO )
  );
  X_INV \block2/CLKAMUX  (
    .I(clkdiv),
    .O(\block2/CLKA_INTNOT )
  );
  defparam block2.INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block2.INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block2.INIT_02 = 256'h00EF0F31100000EF0F31100000EF0F00001F00FF000000FF2900000000096303;
  defparam block2.INIT_03 = 256'hD6F6120000E01F00000039190000181018391900A02531100000000018391900;
  defparam block2.INIT_04 = 256'h002000001F000EE0E0E0E0E000E0004052F795839817B500600074D39514F5D9;
  defparam block2.INIT_05 = 256'h0000575958545653525500A000204D7000E00C00C0CEAD36D736F817B82F39B9;
  defparam block2.INIT_06 = 256'h5957585500A000203900005758595253545556000052555758595354560020B9;
  defparam block2.INIT_07 = 256'h5800A000005253545556575859000052535455575658590020B9000052535456;
  defparam block2.INIT_08 = 256'h00005253545556575859000054575553545658590020B9000054565952535557;
  defparam block2.INIT_09 = 256'h00605B0800607B0800609B080060BB080060DB080060FB0800601B0800603B00;
  defparam block2.INIT_0A = 256'h000000E0000039183737180000E0010080009818140000010000000800C05608;
  defparam block2.INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block2.INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block2.INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block2.INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block2.INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block2.SETUP_ALL = 2701;
  X_RAMB4_S8_S8 block2 (
    .CLKA(\block2/CLKA_INTNOT ),
    .CLKB(clkdiv),
    .ENA(mask_2_OBUF),
    .ENB(\block2/LOGIC_ONE ),
    .RSTA(\block2/LOGIC_ZERO ),
    .RSTB(\block2/LOGIC_ZERO ),
    .WEA(DLX_EXinst_mem_write_EX),
    .WEB(\block2/LOGIC_ZERO ),
    .GSR(GSR),
    .ADDRA({DLX_EXinst_ALU_result[10], DLX_EXinst_ALU_result[9], DLX_EXinst_ALU_result[8], DLX_EXinst_ALU_result[7], DLX_EXinst_ALU_result[6], 
DLX_EXinst_ALU_result[5], DLX_EXinst_ALU_result[4], DLX_EXinst_ALU_result[3], DLX_EXinst_ALU_result[2]}),
    .ADDRB({DLX_IFinst_NPC[10], DLX_IFinst_NPC[9], DLX_IFinst_NPC[8], DLX_IFinst_NPC[7], DLX_IFinst_NPC[6], DLX_IFinst_NPC[5], DLX_IFinst_NPC[4], 
DLX_IFinst_NPC[3], DLX_IFinst_NPC[2]}),
    .DIA({DLX_EXinst_reg_out_B_EX[23], DLX_EXinst_reg_out_B_EX[22], DLX_EXinst_reg_out_B_EX[21], DLX_EXinst_reg_out_B_EX[20], 
DLX_EXinst_reg_out_B_EX[19], DLX_EXinst_reg_out_B_EX[18], DLX_EXinst_reg_out_B_EX[17], DLX_EXinst_reg_out_B_EX[16]}),
    .DIB({\block2/DIB7 , \block2/DIB6 , \block2/DIB5 , \block2/DIB4 , \block2/DIB3 , \block2/DIB2 , \block2/DIB1 , \block2/DIB0 }),
    .DOA({RAM_read_data[23], RAM_read_data[22], RAM_read_data[21], RAM_read_data[20], RAM_read_data[19], RAM_read_data[18], RAM_read_data[17], 
RAM_read_data[16]}),
    .DOB({IR[23], IR[22], IR[21], IR[20], IR[19], IR[18], IR[17], IR[16]})
  );
  X_ONE \block3/LOGIC_ONE_1604  (
    .O(\block3/LOGIC_ONE )
  );
  X_ZERO \block3/LOGIC_ZERO_1605  (
    .O(\block3/LOGIC_ZERO )
  );
  X_INV \block3/CLKAMUX  (
    .I(clkdiv),
    .O(\block3/CLKA_INTNOT )
  );
  defparam block3.INIT_00 = 256'h0000000000000000000000000000000000000000000000000054085454545454;
  defparam block3.INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block3.INIT_02 = 256'h0C253C2622540C253C2622540C253C0000AC540B5454540F2D540C545420243C;
  defparam block3.INIT_03 = 256'h525A2000544B8C540C00273C540CACAC2E273C54142E2626540C540C2E273C54;
  defparam block3.INIT_04 = 256'h5410540C000020ADADADADAD544B54162E26A202020026541200028E023C3202;
  defparam block3.INIT_05 = 256'h54082727272727272727541554160300544B0054152D25AF028F023C31035359;
  defparam block3.INIT_06 = 256'h2F2F2F27541554172E5408272727272727272F5408272F27272727272F54172D;
  defparam block3.INIT_07 = 256'h2F541554082F2F2F272F2F2F2F54082F2F2F2F2F2F2F2F54172D54082F2F2F27;
  defparam block3.INIT_08 = 256'h5408272727272F2F2F2F5408272F2F27272F2F2F54172D540827272F2727272F;
  defparam block3.INIT_09 = 256'h5413822554138225541382255413822554138225541382255413832554138300;
  defparam block3.INIT_0A = 256'h0000544B5417272FAF8F2000544B2054120002696D5408245415002D54168325;
  defparam block3.INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block3.INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block3.INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block3.INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block3.INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam block3.SETUP_ALL = 2701;
  X_RAMB4_S8_S8 block3 (
    .CLKA(\block3/CLKA_INTNOT ),
    .CLKB(clkdiv),
    .ENA(mask_3_OBUF),
    .ENB(\block3/LOGIC_ONE ),
    .RSTA(\block3/LOGIC_ZERO ),
    .RSTB(\block3/LOGIC_ZERO ),
    .WEA(DLX_EXinst_mem_write_EX),
    .WEB(\block3/LOGIC_ZERO ),
    .GSR(GSR),
    .ADDRA({DLX_EXinst_ALU_result[10], DLX_EXinst_ALU_result[9], DLX_EXinst_ALU_result[8], DLX_EXinst_ALU_result[7], DLX_EXinst_ALU_result[6], 
DLX_EXinst_ALU_result[5], DLX_EXinst_ALU_result[4], DLX_EXinst_ALU_result[3], DLX_EXinst_ALU_result[2]}),
    .ADDRB({DLX_IFinst_NPC[10], DLX_IFinst_NPC[9], DLX_IFinst_NPC[8], DLX_IFinst_NPC[7], DLX_IFinst_NPC[6], DLX_IFinst_NPC[5], DLX_IFinst_NPC[4], 
DLX_IFinst_NPC[3], DLX_IFinst_NPC[2]}),
    .DIA({DLX_EXinst_reg_out_B_EX[31], DLX_EXinst_reg_out_B_EX[30], DLX_EXinst_reg_out_B_EX[29], DLX_EXinst_reg_out_B_EX[28], 
DLX_EXinst_reg_out_B_EX[27], DLX_EXinst_reg_out_B_EX[26], DLX_EXinst_reg_out_B_EX[25], DLX_EXinst_reg_out_B_EX[24]}),
    .DIB({\block3/DIB7 , \block3/DIB6 , \block3/DIB5 , \block3/DIB4 , \block3/DIB3 , \block3/DIB2 , \block3/DIB1 , \block3/DIB0 }),
    .DOA({RAM_read_data[31], RAM_read_data[30], RAM_read_data[29], RAM_read_data[28], RAM_read_data[27], RAM_read_data[26], RAM_read_data[25], 
RAM_read_data[24]}),
    .DOB({IR_MSB_7_OBUF, IR_MSB_6_OBUF, IR_MSB_5_OBUF, IR_MSB_4_OBUF, IR_MSB_3_OBUF, IR_MSB_2_OBUF, IR_MSB_1_OBUF, IR_MSB_0_OBUF})
  );
  defparam DLX_IDinst_RegFile_28_25_1606.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_28_25_1606 (
    .I(DLX_IDinst_WB_data_eff[25]),
    .CE(DLX_IDinst__n0606),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_28_25)
  );
  X_MUX2 \DLX_EXinst_Mshift__n0019_Sh<24>281  (
    .IA(N165606),
    .IB(N165608),
    .SEL(DLX_IDinst_reg_out_B[0]),
    .O(\DLX_EXinst_Mshift__n0019_Sh<24>/F5MUX )
  );
  defparam \DLX_EXinst_Mshift__n0019_Sh<24>281_G .INIT = 16'hCFC0;
  X_LUT4 \DLX_EXinst_Mshift__n0019_Sh<24>281_G  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[27]),
    .ADR2(DLX_IDinst_reg_out_B[1]),
    .ADR3(DLX_IDinst_reg_out_A[25]),
    .O(N165608)
  );
  defparam \DLX_EXinst_Mshift__n0019_Sh<24>281_F .INIT = 16'hF0CC;
  X_LUT4 \DLX_EXinst_Mshift__n0019_Sh<24>281_F  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[24]),
    .ADR2(DLX_IDinst_reg_out_A[26]),
    .ADR3(DLX_IDinst_reg_out_B[1]),
    .O(N165606)
  );
  X_BUF \DLX_EXinst_Mshift__n0019_Sh<24>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0019_Sh<24>/F5MUX ),
    .O(\DLX_EXinst_Mshift__n0019_Sh[24] )
  );
  X_MUX2 \DLX_EXinst_Mshift__n0019_Sh<25>281  (
    .IA(N165526),
    .IB(N165528),
    .SEL(DLX_IDinst_reg_out_B[1]),
    .O(\DLX_EXinst_Mshift__n0019_Sh<25>/F5MUX )
  );
  defparam \DLX_EXinst_Mshift__n0019_Sh<25>281_G .INIT = 16'hAAF0;
  X_LUT4 \DLX_EXinst_Mshift__n0019_Sh<25>281_G  (
    .ADR0(DLX_IDinst_reg_out_A[28]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[27]),
    .ADR3(DLX_IDinst_reg_out_B[0]),
    .O(N165528)
  );
  defparam \DLX_EXinst_Mshift__n0019_Sh<25>281_F .INIT = 16'hB8B8;
  X_LUT4 \DLX_EXinst_Mshift__n0019_Sh<25>281_F  (
    .ADR0(DLX_IDinst_reg_out_A[26]),
    .ADR1(DLX_IDinst_reg_out_B[0]),
    .ADR2(DLX_IDinst_reg_out_A[25]),
    .ADR3(VCC),
    .O(N165526)
  );
  X_BUF \DLX_EXinst_Mshift__n0019_Sh<25>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0019_Sh<25>/F5MUX ),
    .O(\DLX_EXinst_Mshift__n0019_Sh[25] )
  );
  X_MUX2 \DLX_EXinst_Mshift__n0019_Sh<26>281  (
    .IA(N165336),
    .IB(N165338),
    .SEL(DLX_IDinst_reg_out_B[0]),
    .O(\DLX_EXinst_Mshift__n0019_Sh<26>/F5MUX )
  );
  defparam \DLX_EXinst_Mshift__n0019_Sh<26>281_G .INIT = 16'hF5A0;
  X_LUT4 \DLX_EXinst_Mshift__n0019_Sh<26>281_G  (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[29]),
    .ADR3(DLX_IDinst_reg_out_A[27]),
    .O(N165338)
  );
  defparam \DLX_EXinst_Mshift__n0019_Sh<26>281_F .INIT = 16'hEE44;
  X_LUT4 \DLX_EXinst_Mshift__n0019_Sh<26>281_F  (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(DLX_IDinst_reg_out_A[26]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[28]),
    .O(N165336)
  );
  X_BUF \DLX_EXinst_Mshift__n0019_Sh<26>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0019_Sh<26>/F5MUX ),
    .O(\DLX_EXinst_Mshift__n0019_Sh[26] )
  );
  X_MUX2 \DLX_EXinst_Mshift__n0019_Sh<28>281  (
    .IA(N165586),
    .IB(N165588),
    .SEL(DLX_IDinst_reg_out_B[1]),
    .O(\DLX_EXinst_Mshift__n0019_Sh<28>/F5MUX )
  );
  defparam \DLX_EXinst_Mshift__n0019_Sh<28>281_G .INIT = 16'hCACA;
  X_LUT4 \DLX_EXinst_Mshift__n0019_Sh<28>281_G  (
    .ADR0(DLX_IDinst_reg_out_A[30]),
    .ADR1(DLX_IDinst_reg_out_A[31]),
    .ADR2(DLX_IDinst_reg_out_B[0]),
    .ADR3(VCC),
    .O(N165588)
  );
  defparam \DLX_EXinst_Mshift__n0019_Sh<28>281_F .INIT = 16'hACAC;
  X_LUT4 \DLX_EXinst_Mshift__n0019_Sh<28>281_F  (
    .ADR0(DLX_IDinst_reg_out_A[29]),
    .ADR1(DLX_IDinst_reg_out_A[28]),
    .ADR2(DLX_IDinst_reg_out_B[0]),
    .ADR3(VCC),
    .O(N165586)
  );
  X_BUF \DLX_EXinst_Mshift__n0019_Sh<28>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0019_Sh<28>/F5MUX ),
    .O(\DLX_EXinst_Mshift__n0019_Sh[28] )
  );
  X_MUX2 \DLX_EXinst_Mshift__n0021_Sh<43>1  (
    .IA(N165511),
    .IB(N165513),
    .SEL(DLX_IDinst_Imm_2_1),
    .O(\DLX_EXinst_Mshift__n0021_Sh<43>/F5MUX )
  );
  defparam \DLX_EXinst_Mshift__n0021_Sh<43>1_G .INIT = 16'h00E2;
  X_LUT4 \DLX_EXinst_Mshift__n0021_Sh<43>1_G  (
    .ADR0(DLX_EXinst_N72933),
    .ADR1(DLX_IDinst_Imm_0_1),
    .ADR2(N130725),
    .ADR3(DLX_IDinst_Imm_3_1),
    .O(N165513)
  );
  defparam \DLX_EXinst_Mshift__n0021_Sh<43>1_F .INIT = 16'hE2E2;
  X_LUT4 \DLX_EXinst_Mshift__n0021_Sh<43>1_F  (
    .ADR0(\DLX_EXinst_Mshift__n0021_Sh[11] ),
    .ADR1(DLX_IDinst_Imm_3_1),
    .ADR2(\DLX_EXinst_Mshift__n0021_Sh[3] ),
    .ADR3(VCC),
    .O(N165511)
  );
  X_BUF \DLX_EXinst_Mshift__n0021_Sh<43>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0021_Sh<43>/F5MUX ),
    .O(\DLX_EXinst_Mshift__n0021_Sh[43] )
  );
  X_MUX2 \DLX_EXinst_Mshift__n0022_Sh<59>1  (
    .IA(N165941),
    .IB(N165943),
    .SEL(DLX_IDinst_Imm_2_1),
    .O(\DLX_EXinst_Mshift__n0022_Sh<59>/F5MUX )
  );
  defparam \DLX_EXinst_Mshift__n0022_Sh<59>1_G .INIT = 16'h0010;
  X_LUT4 \DLX_EXinst_Mshift__n0022_Sh<59>1_G  (
    .ADR0(DLX_IDinst_Imm_0_1),
    .ADR1(DLX_IDinst_Imm_3_1),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(DLX_IDinst_Imm_1_1),
    .O(N165943)
  );
  defparam \DLX_EXinst_Mshift__n0022_Sh<59>1_F .INIT = 16'h4540;
  X_LUT4 \DLX_EXinst_Mshift__n0022_Sh<59>1_F  (
    .ADR0(DLX_IDinst_Imm_3_1),
    .ADR1(DLX_EXinst_N72791),
    .ADR2(DLX_IDinst_Imm_1_1),
    .ADR3(N130467),
    .O(N165941)
  );
  X_BUF \DLX_EXinst_Mshift__n0022_Sh<59>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0022_Sh<59>/F5MUX ),
    .O(\DLX_EXinst_Mshift__n0022_Sh[59] )
  );
  X_MUX2 \DLX_EXinst_Mshift__n0023_Sh<40>1  (
    .IA(N165771),
    .IB(N165773),
    .SEL(DLX_IDinst_reg_out_B_3_1),
    .O(\DLX_EXinst_Mshift__n0023_Sh<40>/F5MUX )
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<40>1_G .INIT = 16'h0010;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<40>1_G  (
    .ADR0(DLX_IDinst_reg_out_B_2_1),
    .ADR1(DLX_IDinst_reg_out_B[0]),
    .ADR2(DLX_IDinst_reg_out_A[0]),
    .ADR3(DLX_IDinst_reg_out_B[1]),
    .O(N165773)
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<40>1_F .INIT = 16'hFA0A;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<40>1_F  (
    .ADR0(\DLX_EXinst_Mshift__n0023_Sh[8] ),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B_2_1),
    .ADR3(\DLX_EXinst_Mshift__n0023_Sh[4] ),
    .O(N165771)
  );
  X_BUF \DLX_EXinst_Mshift__n0023_Sh<40>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0023_Sh<40>/F5MUX ),
    .O(\DLX_EXinst_Mshift__n0023_Sh[40] )
  );
  X_MUX2 \DLX_EXinst_Mshift__n0021_Sh<3>281  (
    .IA(N165371),
    .IB(N165373),
    .SEL(DLX_IDinst_Imm_1_1),
    .O(\DLX_EXinst_Mshift__n0021_Sh<3>/F5MUX )
  );
  defparam \DLX_EXinst_Mshift__n0021_Sh<3>281_G .INIT = 16'hFA0A;
  X_LUT4 \DLX_EXinst_Mshift__n0021_Sh<3>281_G  (
    .ADR0(DLX_IDinst_reg_out_A[1]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_Imm_0_1),
    .ADR3(DLX_IDinst_reg_out_A[0]),
    .O(N165373)
  );
  defparam \DLX_EXinst_Mshift__n0021_Sh<3>281_F .INIT = 16'hF0CC;
  X_LUT4 \DLX_EXinst_Mshift__n0021_Sh<3>281_F  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[3]),
    .ADR2(DLX_IDinst_reg_out_A[2]),
    .ADR3(DLX_IDinst_Imm_0_1),
    .O(N165371)
  );
  X_BUF \DLX_EXinst_Mshift__n0021_Sh<3>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0021_Sh<3>/F5MUX ),
    .O(\DLX_EXinst_Mshift__n0021_Sh[3] )
  );
  X_MUX2 \DLX_EXinst_Mshift__n0021_Sh<4>281  (
    .IA(N165331),
    .IB(N165333),
    .SEL(DLX_IDinst_Imm_1_1),
    .O(\DLX_EXinst_Mshift__n0021_Sh<4>/F5MUX )
  );
  defparam \DLX_EXinst_Mshift__n0021_Sh<4>281_G .INIT = 16'hE4E4;
  X_LUT4 \DLX_EXinst_Mshift__n0021_Sh<4>281_G  (
    .ADR0(DLX_IDinst_Imm_0_1),
    .ADR1(DLX_IDinst_reg_out_A[2]),
    .ADR2(DLX_IDinst_reg_out_A[1]),
    .ADR3(VCC),
    .O(N165333)
  );
  defparam \DLX_EXinst_Mshift__n0021_Sh<4>281_F .INIT = 16'hD8D8;
  X_LUT4 \DLX_EXinst_Mshift__n0021_Sh<4>281_F  (
    .ADR0(DLX_IDinst_Imm_0_1),
    .ADR1(DLX_IDinst_reg_out_A[3]),
    .ADR2(DLX_IDinst_reg_out_A[4]),
    .ADR3(VCC),
    .O(N165331)
  );
  X_BUF \DLX_EXinst_Mshift__n0021_Sh<4>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0021_Sh<4>/F5MUX ),
    .O(\DLX_EXinst_Mshift__n0021_Sh[4] )
  );
  X_MUX2 \DLX_EXinst_Mshift__n0021_Sh<5>281  (
    .IA(N165636),
    .IB(N165638),
    .SEL(DLX_IDinst_Imm_0_1),
    .O(\DLX_EXinst_Mshift__n0021_Sh<5>/F5MUX )
  );
  defparam \DLX_EXinst_Mshift__n0021_Sh<5>281_G .INIT = 16'hACAC;
  X_LUT4 \DLX_EXinst_Mshift__n0021_Sh<5>281_G  (
    .ADR0(DLX_IDinst_reg_out_A[2]),
    .ADR1(DLX_IDinst_reg_out_A[4]),
    .ADR2(DLX_IDinst_Imm_1_1),
    .ADR3(VCC),
    .O(N165638)
  );
  defparam \DLX_EXinst_Mshift__n0021_Sh<5>281_F .INIT = 16'hACAC;
  X_LUT4 \DLX_EXinst_Mshift__n0021_Sh<5>281_F  (
    .ADR0(DLX_IDinst_reg_out_A[3]),
    .ADR1(DLX_IDinst_reg_out_A[5]),
    .ADR2(DLX_IDinst_Imm_1_1),
    .ADR3(VCC),
    .O(N165636)
  );
  X_BUF \DLX_EXinst_Mshift__n0021_Sh<5>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0021_Sh<5>/F5MUX ),
    .O(\DLX_EXinst_Mshift__n0021_Sh[5] )
  );
  X_MUX2 \DLX_EXinst_Mshift__n0021_Sh<6>281  (
    .IA(N165341),
    .IB(N165343),
    .SEL(DLX_IDinst_Imm_0_1),
    .O(\DLX_EXinst_Mshift__n0021_Sh<6>/F5MUX )
  );
  defparam \DLX_EXinst_Mshift__n0021_Sh<6>281_G .INIT = 16'hBB88;
  X_LUT4 \DLX_EXinst_Mshift__n0021_Sh<6>281_G  (
    .ADR0(DLX_IDinst_reg_out_A[3]),
    .ADR1(DLX_IDinst_Imm_1_1),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[5]),
    .O(N165343)
  );
  defparam \DLX_EXinst_Mshift__n0021_Sh<6>281_F .INIT = 16'hFC0C;
  X_LUT4 \DLX_EXinst_Mshift__n0021_Sh<6>281_F  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[6]),
    .ADR2(DLX_IDinst_Imm_1_1),
    .ADR3(DLX_IDinst_reg_out_A[4]),
    .O(N165341)
  );
  X_BUF \DLX_EXinst_Mshift__n0021_Sh<6>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0021_Sh<6>/F5MUX ),
    .O(\DLX_EXinst_Mshift__n0021_Sh[6] )
  );
  X_MUX2 \DLX_EXinst__n0007<21>341  (
    .IA(N165366),
    .IB(N165368),
    .SEL(\DLX_IDinst_Imm[2] ),
    .O(\CHOICE4135/F5MUX )
  );
  defparam \DLX_EXinst__n0007<21>341_G .INIT = 16'h2F20;
  X_LUT4 \DLX_EXinst__n0007<21>341_G  (
    .ADR0(\DLX_EXinst_Mshift__n0021_Sh[1] ),
    .ADR1(\DLX_IDinst_Imm[3] ),
    .ADR2(\DLX_IDinst_Imm[4] ),
    .ADR3(DLX_EXinst_N73993),
    .O(N165368)
  );
  defparam \DLX_EXinst__n0007<21>341_F .INIT = 16'h5C0C;
  X_LUT4 \DLX_EXinst__n0007<21>341_F  (
    .ADR0(\DLX_IDinst_Imm[3] ),
    .ADR1(DLX_EXinst_N74196),
    .ADR2(\DLX_IDinst_Imm[4] ),
    .ADR3(\DLX_EXinst_Mshift__n0021_Sh[5] ),
    .O(N165366)
  );
  X_BUF \CHOICE4135/XUSED  (
    .I(\CHOICE4135/F5MUX ),
    .O(CHOICE4135)
  );
  X_MUX2 \DLX_EXinst__n0007<22>341  (
    .IA(N165361),
    .IB(N165363),
    .SEL(\DLX_IDinst_Imm[2] ),
    .O(\CHOICE4070/F5MUX )
  );
  defparam \DLX_EXinst__n0007<22>341_G .INIT = 16'h7250;
  X_LUT4 \DLX_EXinst__n0007<22>341_G  (
    .ADR0(\DLX_IDinst_Imm[4] ),
    .ADR1(\DLX_IDinst_Imm[3] ),
    .ADR2(DLX_EXinst_N73998),
    .ADR3(\DLX_EXinst_Mshift__n0021_Sh[2] ),
    .O(N165363)
  );
  defparam \DLX_EXinst__n0007<22>341_F .INIT = 16'h7250;
  X_LUT4 \DLX_EXinst__n0007<22>341_F  (
    .ADR0(\DLX_IDinst_Imm[4] ),
    .ADR1(\DLX_IDinst_Imm[3] ),
    .ADR2(DLX_EXinst_N74201),
    .ADR3(\DLX_EXinst_Mshift__n0021_Sh[6] ),
    .O(N165361)
  );
  X_BUF \CHOICE4070/XUSED  (
    .I(\CHOICE4070/F5MUX ),
    .O(CHOICE4070)
  );
  X_MUX2 \DLX_EXinst__n0007<30>641  (
    .IA(N165496),
    .IB(N165498),
    .SEL(\DLX_IDinst_Imm[4] ),
    .O(\CHOICE4721/F5MUX )
  );
  defparam \DLX_EXinst__n0007<30>641_G .INIT = 16'hA088;
  X_LUT4 \DLX_EXinst__n0007<30>641_G  (
    .ADR0(DLX_EXinst_N76318),
    .ADR1(N130311),
    .ADR2(DLX_EXinst_N72993),
    .ADR3(\DLX_IDinst_Imm[3] ),
    .O(N165498)
  );
  defparam \DLX_EXinst__n0007<30>641_F .INIT = 16'hA820;
  X_LUT4 \DLX_EXinst__n0007<30>641_F  (
    .ADR0(DLX_EXinst_N76318),
    .ADR1(\DLX_IDinst_Imm[2] ),
    .ADR2(CHOICE4716),
    .ADR3(N134128),
    .O(N165496)
  );
  X_BUF \CHOICE4721/XUSED  (
    .I(\CHOICE4721/F5MUX ),
    .O(CHOICE4721)
  );
  X_MUX2 \DLX_EXinst__n0007<23>341  (
    .IA(N165531),
    .IB(N165533),
    .SEL(\DLX_IDinst_Imm[2] ),
    .O(\CHOICE4005/F5MUX )
  );
  defparam \DLX_EXinst__n0007<23>341_G .INIT = 16'h0ACC;
  X_LUT4 \DLX_EXinst__n0007<23>341_G  (
    .ADR0(\DLX_EXinst_Mshift__n0021_Sh[3] ),
    .ADR1(DLX_EXinst_N74003),
    .ADR2(\DLX_IDinst_Imm[3] ),
    .ADR3(\DLX_IDinst_Imm[4] ),
    .O(N165533)
  );
  defparam \DLX_EXinst__n0007<23>341_F .INIT = 16'h22F0;
  X_LUT4 \DLX_EXinst__n0007<23>341_F  (
    .ADR0(\DLX_EXinst_Mshift__n0021_Sh[7] ),
    .ADR1(\DLX_IDinst_Imm[3] ),
    .ADR2(DLX_EXinst_N74206),
    .ADR3(\DLX_IDinst_Imm[4] ),
    .O(N165531)
  );
  X_BUF \CHOICE4005/XUSED  (
    .I(\CHOICE4005/F5MUX ),
    .O(CHOICE4005)
  );
  X_MUX2 \DLX_EXinst__n0007<30>941  (
    .IA(N165846),
    .IB(N165848),
    .SEL(DLX_IDinst_IR_opcode_field[0]),
    .O(\CHOICE4729/F5MUX )
  );
  defparam \DLX_EXinst__n0007<30>941_G .INIT = 16'hE200;
  X_LUT4 \DLX_EXinst__n0007<30>941_G  (
    .ADR0(\DLX_IDinst_Imm[31] ),
    .ADR1(DLX_IDinst_IR_opcode_field[1]),
    .ADR2(\DLX_IDinst_Imm[14] ),
    .ADR3(DLX_EXinst_N76011),
    .O(N165848)
  );
  defparam \DLX_EXinst__n0007<30>941_F .INIT = 16'h2800;
  X_LUT4 \DLX_EXinst__n0007<30>941_F  (
    .ADR0(\DLX_IDinst_Imm[31] ),
    .ADR1(DLX_IDinst_IR_opcode_field[1]),
    .ADR2(DLX_IDinst_reg_out_A[30]),
    .ADR3(DLX_EXinst_N76011),
    .O(N165846)
  );
  X_BUF \CHOICE4729/XUSED  (
    .I(\CHOICE4729/F5MUX ),
    .O(CHOICE4729)
  );
  X_MUX2 \DLX_EXinst__n0007<0>1431  (
    .IA(N165521),
    .IB(N165523),
    .SEL(DLX_IDinst_reg_out_B[4]),
    .O(\CHOICE5896/F5MUX )
  );
  defparam \DLX_EXinst__n0007<0>1431_G .INIT = 16'hA0C0;
  X_LUT4 \DLX_EXinst__n0007<0>1431_G  (
    .ADR0(DLX_EXinst_N72809),
    .ADR1(DLX_EXinst_N74721),
    .ADR2(DLX_EXinst_N72710),
    .ADR3(DLX_IDinst_reg_out_B[2]),
    .O(N165523)
  );
  defparam \DLX_EXinst__n0007<0>1431_F .INIT = 16'hC480;
  X_LUT4 \DLX_EXinst__n0007<0>1431_F  (
    .ADR0(DLX_IDinst_reg_out_B[2]),
    .ADR1(DLX_EXinst_N72710),
    .ADR2(N137448),
    .ADR3(CHOICE5890),
    .O(N165521)
  );
  X_BUF \CHOICE5896/XUSED  (
    .I(\CHOICE5896/F5MUX ),
    .O(CHOICE5896)
  );
  X_MUX2 \DLX_EXinst__n0007<16>351  (
    .IA(N165631),
    .IB(N165633),
    .SEL(DLX_IDinst_reg_out_B[2]),
    .O(\CHOICE4573/F5MUX )
  );
  defparam \DLX_EXinst__n0007<16>351_G .INIT = 16'h00E2;
  X_LUT4 \DLX_EXinst__n0007<16>351_G  (
    .ADR0(\DLX_EXinst_Mshift__n0023_Sh[12] ),
    .ADR1(DLX_IDinst_reg_out_B[3]),
    .ADR2(\DLX_EXinst_Mshift__n0023_Sh[4] ),
    .ADR3(DLX_IDinst_reg_out_B[4]),
    .O(N165633)
  );
  defparam \DLX_EXinst__n0007<16>351_F .INIT = 16'h5410;
  X_LUT4 \DLX_EXinst__n0007<16>351_F  (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(DLX_IDinst_reg_out_B[3]),
    .ADR2(\DLX_EXinst_Mshift__n0023_Sh[16] ),
    .ADR3(\DLX_EXinst_Mshift__n0023_Sh[8] ),
    .O(N165631)
  );
  X_BUF \CHOICE4573/XUSED  (
    .I(\CHOICE4573/F5MUX ),
    .O(CHOICE4573)
  );
  X_MUX2 \DLX_EXinst__n0007<31>851  (
    .IA(N165516),
    .IB(N165518),
    .SEL(DLX_IDinst_reg_out_B[0]),
    .O(\CHOICE5791/F5MUX )
  );
  defparam \DLX_EXinst__n0007<31>851_G .INIT = 16'hFACA;
  X_LUT4 \DLX_EXinst__n0007<31>851_G  (
    .ADR0(DLX_IDinst_reg_out_A[30]),
    .ADR1(DLX_IDinst_reg_out_A[28]),
    .ADR2(DLX_IDinst_reg_out_B[1]),
    .ADR3(\DLX_EXinst_Mshift__n0024_Sh[31] ),
    .O(N165518)
  );
  defparam \DLX_EXinst__n0007<31>851_F .INIT = 16'hF5A0;
  X_LUT4 \DLX_EXinst__n0007<31>851_F  (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[29]),
    .ADR3(DLX_IDinst_reg_out_A[31]),
    .O(N165516)
  );
  X_BUF \CHOICE5791/XUSED  (
    .I(\CHOICE5791/F5MUX ),
    .O(CHOICE5791)
  );
  X_MUX2 \DLX_EXinst__n0007<17>741  (
    .IA(N165591),
    .IB(N165593),
    .SEL(\DLX_IDinst_Imm[3] ),
    .O(\CHOICE5378/F5MUX )
  );
  defparam \DLX_EXinst__n0007<17>741_G .INIT = 16'hE020;
  X_LUT4 \DLX_EXinst__n0007<17>741_G  (
    .ADR0(\DLX_EXinst_Mshift__n0021_Sh[9] ),
    .ADR1(\DLX_IDinst_Imm[2] ),
    .ADR2(DLX_EXinst__n0055),
    .ADR3(\DLX_EXinst_Mshift__n0021_Sh[5] ),
    .O(N165593)
  );
  defparam \DLX_EXinst__n0007<17>741_F .INIT = 16'hAC00;
  X_LUT4 \DLX_EXinst__n0007<17>741_F  (
    .ADR0(\DLX_EXinst_Mshift__n0021_Sh[13] ),
    .ADR1(N130209),
    .ADR2(\DLX_IDinst_Imm[2] ),
    .ADR3(DLX_EXinst__n0055),
    .O(N165591)
  );
  X_BUF \CHOICE5378/XUSED  (
    .I(\CHOICE5378/F5MUX ),
    .O(CHOICE5378)
  );
  X_MUX2 \DLX_EXinst__n0007<0>6531  (
    .IA(N165416),
    .IB(N165418),
    .SEL(\DLX_IDinst_Imm[2] ),
    .O(\CHOICE5999/F5MUX )
  );
  defparam \DLX_EXinst__n0007<0>6531_G .INIT = 16'hE0A0;
  X_LUT4 \DLX_EXinst__n0007<0>6531_G  (
    .ADR0(CHOICE1791),
    .ADR1(\DLX_EXinst_Mshift__n0022_Sh[12] ),
    .ADR2(DLX_EXinst_N73267),
    .ADR3(\DLX_IDinst_Imm[3] ),
    .O(N165418)
  );
  defparam \DLX_EXinst__n0007<0>6531_F .INIT = 16'hC0A0;
  X_LUT4 \DLX_EXinst__n0007<0>6531_F  (
    .ADR0(CHOICE5994),
    .ADR1(\DLX_EXinst_Mshift__n0022_Sh[8] ),
    .ADR2(DLX_EXinst_N73267),
    .ADR3(\DLX_IDinst_Imm[3] ),
    .O(N165416)
  );
  X_BUF \CHOICE5999/XUSED  (
    .I(\CHOICE5999/F5MUX ),
    .O(CHOICE5999)
  );
  defparam DLX_IDinst_RegFile_28_26_1607.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_28_26_1607 (
    .I(DLX_IDinst_WB_data_eff[26]),
    .CE(DLX_IDinst__n0606),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_28_26)
  );
  X_MUX2 \DLX_EXinst__n0007<18>741  (
    .IA(N165451),
    .IB(N165453),
    .SEL(\DLX_IDinst_Imm[3] ),
    .O(\CHOICE5220/F5MUX )
  );
  defparam \DLX_EXinst__n0007<18>741_G .INIT = 16'hA280;
  X_LUT4 \DLX_EXinst__n0007<18>741_G  (
    .ADR0(DLX_EXinst__n0055),
    .ADR1(\DLX_IDinst_Imm[2] ),
    .ADR2(\DLX_EXinst_Mshift__n0021_Sh[6] ),
    .ADR3(\DLX_EXinst_Mshift__n0021_Sh[10] ),
    .O(N165453)
  );
  defparam \DLX_EXinst__n0007<18>741_F .INIT = 16'h88A0;
  X_LUT4 \DLX_EXinst__n0007<18>741_F  (
    .ADR0(DLX_EXinst__n0055),
    .ADR1(\DLX_EXinst_Mshift__n0021_Sh[14] ),
    .ADR2(N130261),
    .ADR3(\DLX_IDinst_Imm[2] ),
    .O(N165451)
  );
  X_BUF \CHOICE5220/XUSED  (
    .I(\CHOICE5220/F5MUX ),
    .O(CHOICE5220)
  );
  X_MUX2 \DLX_EXinst__n0007<19>741  (
    .IA(N165411),
    .IB(N165413),
    .SEL(\DLX_IDinst_Imm[3] ),
    .O(\CHOICE5299/F5MUX )
  );
  defparam \DLX_EXinst__n0007<19>741_G .INIT = 16'hB080;
  X_LUT4 \DLX_EXinst__n0007<19>741_G  (
    .ADR0(\DLX_EXinst_Mshift__n0021_Sh[7] ),
    .ADR1(\DLX_IDinst_Imm[2] ),
    .ADR2(DLX_EXinst__n0055),
    .ADR3(\DLX_EXinst_Mshift__n0021_Sh[11] ),
    .O(N165413)
  );
  defparam \DLX_EXinst__n0007<19>741_F .INIT = 16'hC840;
  X_LUT4 \DLX_EXinst__n0007<19>741_F  (
    .ADR0(\DLX_IDinst_Imm[2] ),
    .ADR1(DLX_EXinst__n0055),
    .ADR2(\DLX_EXinst_Mshift__n0021_Sh[19] ),
    .ADR3(\DLX_EXinst_Mshift__n0021_Sh[15] ),
    .O(N165411)
  );
  X_BUF \CHOICE5299/XUSED  (
    .I(\CHOICE5299/F5MUX ),
    .O(CHOICE5299)
  );
  X_MUX2 \DLX_EXinst__n0007<28>861  (
    .IA(N165421),
    .IB(N165423),
    .SEL(\DLX_IDinst_Imm[3] ),
    .O(\CHOICE4866/F5MUX )
  );
  defparam \DLX_EXinst__n0007<28>861_G .INIT = 16'hE200;
  X_LUT4 \DLX_EXinst__n0007<28>861_G  (
    .ADR0(DLX_EXinst_N75377),
    .ADR1(\DLX_IDinst_Imm[4] ),
    .ADR2(DLX_EXinst_N72983),
    .ADR3(DLX_EXinst_N76318),
    .O(N165423)
  );
  defparam \DLX_EXinst__n0007<28>861_F .INIT = 16'hE200;
  X_LUT4 \DLX_EXinst__n0007<28>861_F  (
    .ADR0(CHOICE4861),
    .ADR1(\DLX_IDinst_Imm[4] ),
    .ADR2(DLX_EXinst_N74223),
    .ADR3(DLX_EXinst_N76318),
    .O(N165421)
  );
  X_BUF \CHOICE4866/XUSED  (
    .I(\CHOICE4866/F5MUX ),
    .O(CHOICE4866)
  );
  defparam DLX_IDinst_RegFile_28_17_1608.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_28_17_1608 (
    .I(DLX_IDinst_WB_data_eff[17]),
    .CE(DLX_IDinst__n0606),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_28_17)
  );
  X_MUX2 \DLX_EXinst__n0007<29>641  (
    .IA(N165491),
    .IB(N165493),
    .SEL(\DLX_IDinst_Imm[4] ),
    .O(\CHOICE4792/F5MUX )
  );
  defparam \DLX_EXinst__n0007<29>641_G .INIT = 16'hB080;
  X_LUT4 \DLX_EXinst__n0007<29>641_G  (
    .ADR0(DLX_EXinst_N72988),
    .ADR1(\DLX_IDinst_Imm[3] ),
    .ADR2(DLX_EXinst_N76318),
    .ADR3(N130363),
    .O(N165493)
  );
  defparam \DLX_EXinst__n0007<29>641_F .INIT = 16'hC808;
  X_LUT4 \DLX_EXinst__n0007<29>641_F  (
    .ADR0(CHOICE4787),
    .ADR1(DLX_EXinst_N76318),
    .ADR2(\DLX_IDinst_Imm[2] ),
    .ADR3(N133768),
    .O(N165491)
  );
  X_BUF \CHOICE4792/XUSED  (
    .I(\CHOICE4792/F5MUX ),
    .O(CHOICE4792)
  );
  X_MUX2 \DLX_EXinst_Mshift__n0019_Sh<27>1  (
    .IA(N165571),
    .IB(N165573),
    .SEL(DLX_IDinst_reg_out_B[1]),
    .O(\DLX_EXinst_Mshift__n0019_Sh<27>/F5MUX )
  );
  defparam \DLX_EXinst_Mshift__n0019_Sh<27>1_G .INIT = 16'hCCAA;
  X_LUT4 \DLX_EXinst_Mshift__n0019_Sh<27>1_G  (
    .ADR0(DLX_IDinst_reg_out_A[29]),
    .ADR1(DLX_IDinst_reg_out_A[30]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[0]),
    .O(N165573)
  );
  defparam \DLX_EXinst_Mshift__n0019_Sh<27>1_F .INIT = 16'hFC30;
  X_LUT4 \DLX_EXinst_Mshift__n0019_Sh<27>1_F  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_B[0]),
    .ADR2(DLX_IDinst_reg_out_A[27]),
    .ADR3(DLX_IDinst_reg_out_A[28]),
    .O(N165571)
  );
  X_BUF \DLX_EXinst_Mshift__n0019_Sh<27>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0019_Sh<27>/F5MUX ),
    .O(\DLX_EXinst_Mshift__n0019_Sh[27] )
  );
  X_MUX2 \DLX_EXinst__n0007<29>941  (
    .IA(N165916),
    .IB(N165918),
    .SEL(DLX_IDinst_IR_opcode_field[0]),
    .O(\CHOICE4800/F5MUX )
  );
  defparam \DLX_EXinst__n0007<29>941_G .INIT = 16'h8A80;
  X_LUT4 \DLX_EXinst__n0007<29>941_G  (
    .ADR0(DLX_EXinst_N76011),
    .ADR1(\DLX_IDinst_Imm[13] ),
    .ADR2(DLX_IDinst_IR_opcode_field[1]),
    .ADR3(\DLX_IDinst_Imm[31] ),
    .O(N165918)
  );
  defparam \DLX_EXinst__n0007<29>941_F .INIT = 16'h2800;
  X_LUT4 \DLX_EXinst__n0007<29>941_F  (
    .ADR0(DLX_EXinst_N76011),
    .ADR1(DLX_IDinst_reg_out_A[29]),
    .ADR2(DLX_IDinst_IR_opcode_field[1]),
    .ADR3(\DLX_IDinst_Imm[31] ),
    .O(N165916)
  );
  X_BUF \CHOICE4800/XUSED  (
    .I(\CHOICE4800/F5MUX ),
    .O(CHOICE4800)
  );
  X_MUX2 \DLX_EXinst__n0007<8>2861  (
    .IA(N165786),
    .IB(N165788),
    .SEL(DLX_EXinst__n0036),
    .O(\CHOICE5191/F5MUX )
  );
  defparam \DLX_EXinst__n0007<8>2861_G .INIT = 16'hFFFA;
  X_LUT4 \DLX_EXinst__n0007<8>2861_G  (
    .ADR0(CHOICE5132),
    .ADR1(VCC),
    .ADR2(CHOICE5127),
    .ADR3(CHOICE5156),
    .O(N165788)
  );
  defparam \DLX_EXinst__n0007<8>2861_F .INIT = 16'hEEFE;
  X_LUT4 \DLX_EXinst__n0007<8>2861_F  (
    .ADR0(CHOICE5170),
    .ADR1(CHOICE5188),
    .ADR2(CHOICE5165),
    .ADR3(N146478),
    .O(N165786)
  );
  X_BUF \CHOICE5191/XUSED  (
    .I(\CHOICE5191/F5MUX ),
    .O(CHOICE5191)
  );
  X_MUX2 \DLX_EXinst__n0007<9>2341  (
    .IA(N165681),
    .IB(N165683),
    .SEL(DLX_EXinst__n0036),
    .O(\CHOICE4558/F5MUX )
  );
  defparam \DLX_EXinst__n0007<9>2341_G .INIT = 16'hFFFC;
  X_LUT4 \DLX_EXinst__n0007<9>2341_G  (
    .ADR0(VCC),
    .ADR1(CHOICE4505),
    .ADR2(CHOICE4510),
    .ADR3(CHOICE4527),
    .O(N165683)
  );
  defparam \DLX_EXinst__n0007<9>2341_F .INIT = 16'hEFEE;
  X_LUT4 \DLX_EXinst__n0007<9>2341_F  (
    .ADR0(CHOICE4555),
    .ADR1(CHOICE4539),
    .ADR2(N146478),
    .ADR3(CHOICE4534),
    .O(N165681)
  );
  X_BUF \CHOICE4558/XUSED  (
    .I(\CHOICE4558/F5MUX ),
    .O(CHOICE4558)
  );
  X_MUX2 \DLX_EXinst_Mshift__n0020_Sh<25>281  (
    .IA(N165621),
    .IB(N165623),
    .SEL(DLX_IDinst_Imm_0_1),
    .O(\DLX_EXinst_Mshift__n0020_Sh<25>/F5MUX )
  );
  defparam \DLX_EXinst_Mshift__n0020_Sh<25>281_G .INIT = 16'hEE22;
  X_LUT4 \DLX_EXinst_Mshift__n0020_Sh<25>281_G  (
    .ADR0(DLX_IDinst_reg_out_A[26]),
    .ADR1(DLX_IDinst_Imm_1_1),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[28]),
    .O(N165623)
  );
  defparam \DLX_EXinst_Mshift__n0020_Sh<25>281_F .INIT = 16'hF0CC;
  X_LUT4 \DLX_EXinst_Mshift__n0020_Sh<25>281_F  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[25]),
    .ADR2(DLX_IDinst_reg_out_A[27]),
    .ADR3(DLX_IDinst_Imm_1_1),
    .O(N165621)
  );
  X_BUF \DLX_EXinst_Mshift__n0020_Sh<25>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0020_Sh<25>/F5MUX ),
    .O(\DLX_EXinst_Mshift__n0020_Sh[25] )
  );
  X_MUX2 \DLX_EXinst_Mshift__n0020_Sh<26>281  (
    .IA(N165446),
    .IB(N165448),
    .SEL(DLX_IDinst_Imm_0_1),
    .O(\DLX_EXinst_Mshift__n0020_Sh<26>/F5MUX )
  );
  defparam \DLX_EXinst_Mshift__n0020_Sh<26>281_G .INIT = 16'hEE22;
  X_LUT4 \DLX_EXinst_Mshift__n0020_Sh<26>281_G  (
    .ADR0(DLX_IDinst_reg_out_A[27]),
    .ADR1(DLX_IDinst_Imm_1_1),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[29]),
    .O(N165448)
  );
  defparam \DLX_EXinst_Mshift__n0020_Sh<26>281_F .INIT = 16'hF0CC;
  X_LUT4 \DLX_EXinst_Mshift__n0020_Sh<26>281_F  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[26]),
    .ADR2(DLX_IDinst_reg_out_A[28]),
    .ADR3(DLX_IDinst_Imm_1_1),
    .O(N165446)
  );
  X_BUF \DLX_EXinst_Mshift__n0020_Sh<26>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0020_Sh<26>/F5MUX ),
    .O(\DLX_EXinst_Mshift__n0020_Sh[26] )
  );
  X_MUX2 \DLX_EXinst_Mshift__n0020_Sh<28>281  (
    .IA(N165471),
    .IB(N165473),
    .SEL(DLX_IDinst_Imm_1_1),
    .O(\DLX_EXinst_Mshift__n0020_Sh<28>/F5MUX )
  );
  defparam \DLX_EXinst_Mshift__n0020_Sh<28>281_G .INIT = 16'hFA50;
  X_LUT4 \DLX_EXinst_Mshift__n0020_Sh<28>281_G  (
    .ADR0(DLX_IDinst_Imm_0_1),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[30]),
    .ADR3(DLX_IDinst_reg_out_A[31]),
    .O(N165473)
  );
  defparam \DLX_EXinst_Mshift__n0020_Sh<28>281_F .INIT = 16'hCCAA;
  X_LUT4 \DLX_EXinst_Mshift__n0020_Sh<28>281_F  (
    .ADR0(DLX_IDinst_reg_out_A[28]),
    .ADR1(DLX_IDinst_reg_out_A[29]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_Imm_0_1),
    .O(N165471)
  );
  X_BUF \DLX_EXinst_Mshift__n0020_Sh<28>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0020_Sh<28>/F5MUX ),
    .O(\DLX_EXinst_Mshift__n0020_Sh[28] )
  );
  X_MUX2 \DLX_EXinst_Mshift__n0023_Sh<3>281  (
    .IA(N165616),
    .IB(N165618),
    .SEL(DLX_IDinst_reg_out_B[0]),
    .O(\DLX_EXinst_Mshift__n0023_Sh<3>/F5MUX )
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<3>281_G .INIT = 16'hCCF0;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<3>281_G  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[0]),
    .ADR2(DLX_IDinst_reg_out_A[2]),
    .ADR3(DLX_IDinst_reg_out_B[1]),
    .O(N165618)
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<3>281_F .INIT = 16'hE4E4;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<3>281_F  (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(DLX_IDinst_reg_out_A[3]),
    .ADR2(DLX_IDinst_reg_out_A[1]),
    .ADR3(VCC),
    .O(N165616)
  );
  X_BUF \DLX_EXinst_Mshift__n0023_Sh<3>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0023_Sh<3>/F5MUX ),
    .O(\DLX_EXinst_Mshift__n0023_Sh[3] )
  );
  X_MUX2 \DLX_EXinst_Mshift__n0023_Sh<4>281  (
    .IA(N165601),
    .IB(N165603),
    .SEL(DLX_IDinst_reg_out_B[1]),
    .O(\DLX_EXinst_Mshift__n0023_Sh<4>/F5MUX )
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<4>281_G .INIT = 16'hF3C0;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<4>281_G  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_B[0]),
    .ADR2(DLX_IDinst_reg_out_A[1]),
    .ADR3(DLX_IDinst_reg_out_A[2]),
    .O(N165603)
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<4>281_F .INIT = 16'hBB88;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<4>281_F  (
    .ADR0(DLX_IDinst_reg_out_A[3]),
    .ADR1(DLX_IDinst_reg_out_B[0]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[4]),
    .O(N165601)
  );
  X_BUF \DLX_EXinst_Mshift__n0023_Sh<4>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0023_Sh<4>/F5MUX ),
    .O(\DLX_EXinst_Mshift__n0023_Sh[4] )
  );
  X_MUX2 \DLX_EXinst_Mshift__n0023_Sh<5>281  (
    .IA(N165576),
    .IB(N165578),
    .SEL(DLX_IDinst_reg_out_B[1]),
    .O(\DLX_EXinst_Mshift__n0023_Sh<5>/F5MUX )
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<5>281_G .INIT = 16'hD8D8;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<5>281_G  (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(DLX_IDinst_reg_out_A[2]),
    .ADR2(DLX_IDinst_reg_out_A[3]),
    .ADR3(VCC),
    .O(N165578)
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<5>281_F .INIT = 16'hF3C0;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<5>281_F  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_B[0]),
    .ADR2(DLX_IDinst_reg_out_A[4]),
    .ADR3(DLX_IDinst_reg_out_A[5]),
    .O(N165576)
  );
  X_BUF \DLX_EXinst_Mshift__n0023_Sh<5>/XUSED  (
    .I(\DLX_EXinst_Mshift__n0023_Sh<5>/F5MUX ),
    .O(\DLX_EXinst_Mshift__n0023_Sh[5] )
  );
  X_MUX2 \DLX_EXinst__n0007<24>454_SW01  (
    .IA(N165821),
    .IB(N165823),
    .SEL(DLX_IDinst_IR_opcode_field[0]),
    .O(\N163716/F5MUX )
  );
  defparam \DLX_EXinst__n0007<24>454_SW01_G .INIT = 16'h8C80;
  X_LUT4 \DLX_EXinst__n0007<24>454_SW01_G  (
    .ADR0(\DLX_IDinst_Imm[8] ),
    .ADR1(DLX_EXinst_N76011),
    .ADR2(DLX_IDinst_IR_opcode_field[1]),
    .ADR3(\DLX_IDinst_Imm[31] ),
    .O(N165823)
  );
  defparam \DLX_EXinst__n0007<24>454_SW01_F .INIT = 16'h2800;
  X_LUT4 \DLX_EXinst__n0007<24>454_SW01_F  (
    .ADR0(DLX_EXinst_N76011),
    .ADR1(DLX_IDinst_reg_out_A[24]),
    .ADR2(DLX_IDinst_IR_opcode_field[1]),
    .ADR3(\DLX_IDinst_Imm[31] ),
    .O(N165821)
  );
  X_BUF \N163716/XUSED  (
    .I(\N163716/F5MUX ),
    .O(N163716)
  );
  X_MUX2 \DLX_EXinst__n0007<26>110_SW01  (
    .IA(N165401),
    .IB(N165403),
    .SEL(DLX_IDinst_IR_opcode_field[0]),
    .O(\N163242/F5MUX )
  );
  defparam \DLX_EXinst__n0007<26>110_SW01_G .INIT = 16'hA088;
  X_LUT4 \DLX_EXinst__n0007<26>110_SW01_G  (
    .ADR0(DLX_EXinst_N76011),
    .ADR1(\DLX_IDinst_Imm[31] ),
    .ADR2(\DLX_IDinst_Imm[10] ),
    .ADR3(DLX_IDinst_IR_opcode_field[1]),
    .O(N165403)
  );
  defparam \DLX_EXinst__n0007<26>110_SW01_F .INIT = 16'h4800;
  X_LUT4 \DLX_EXinst__n0007<26>110_SW01_F  (
    .ADR0(DLX_IDinst_IR_opcode_field[1]),
    .ADR1(\DLX_IDinst_Imm[31] ),
    .ADR2(DLX_IDinst_reg_out_A[26]),
    .ADR3(DLX_EXinst_N76011),
    .O(N165401)
  );
  X_BUF \N163242/XUSED  (
    .I(\N163242/F5MUX ),
    .O(N163242)
  );
  X_MUX2 \DLX_IFinst__n0003<0>1  (
    .IA(N165781),
    .IB(N165783),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[0])
  );
  defparam \DLX_IFinst__n0003<0>1_G .INIT = 16'hDD88;
  X_LUT4 \DLX_IFinst__n0003<0>1_G  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(IR[0]),
    .ADR2(VCC),
    .ADR3(DLX_IFinst_IR_previous[0]),
    .O(N165783)
  );
  defparam \DLX_IFinst__n0003<0>1_F .INIT = 16'hF4B0;
  X_LUT4 \DLX_IFinst__n0003<0>1_F  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(DLX_IFinst_stalled),
    .ADR2(IR[0]),
    .ADR3(DLX_IFinst_IR_curr[0]),
    .O(N165781)
  );
  X_MUX2 \DLX_IFinst__n0003<1>1  (
    .IA(N165766),
    .IB(N165768),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[1])
  );
  defparam \DLX_IFinst__n0003<1>1_G .INIT = 16'hBB88;
  X_LUT4 \DLX_IFinst__n0003<1>1_G  (
    .ADR0(IR[1]),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(VCC),
    .ADR3(DLX_IFinst_IR_previous[1]),
    .O(N165768)
  );
  defparam \DLX_IFinst__n0003<1>1_F .INIT = 16'hF0D8;
  X_LUT4 \DLX_IFinst__n0003<1>1_F  (
    .ADR0(DLX_IFinst_stalled),
    .ADR1(DLX_IFinst_IR_curr[1]),
    .ADR2(IR[1]),
    .ADR3(DLX_IDinst_branch_sig),
    .O(N165766)
  );
  X_MUX2 \DLX_IFinst__n0003<2>1  (
    .IA(N165746),
    .IB(N165748),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[2])
  );
  defparam \DLX_IFinst__n0003<2>1_G .INIT = 16'hCCAA;
  X_LUT4 \DLX_IFinst__n0003<2>1_G  (
    .ADR0(DLX_IFinst_IR_previous[2]),
    .ADR1(IR[2]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_branch_sig),
    .O(N165748)
  );
  defparam \DLX_IFinst__n0003<2>1_F .INIT = 16'hAEA2;
  X_LUT4 \DLX_IFinst__n0003<2>1_F  (
    .ADR0(IR[2]),
    .ADR1(DLX_IFinst_stalled),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(DLX_IFinst_IR_curr[2]),
    .O(N165746)
  );
  X_MUX2 \DLX_IFinst__n0003<3>1  (
    .IA(N165726),
    .IB(N165728),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[3])
  );
  defparam \DLX_IFinst__n0003<3>1_G .INIT = 16'hAACC;
  X_LUT4 \DLX_IFinst__n0003<3>1_G  (
    .ADR0(IR[3]),
    .ADR1(DLX_IFinst_IR_previous[3]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_branch_sig),
    .O(N165728)
  );
  defparam \DLX_IFinst__n0003<3>1_F .INIT = 16'hDC8C;
  X_LUT4 \DLX_IFinst__n0003<3>1_F  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(IR[3]),
    .ADR2(DLX_IFinst_stalled),
    .ADR3(DLX_IFinst_IR_curr[3]),
    .O(N165726)
  );
  X_MUX2 \DLX_IFinst__n0003<4>1  (
    .IA(N165721),
    .IB(N165723),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[4])
  );
  defparam \DLX_IFinst__n0003<4>1_G .INIT = 16'hD8D8;
  X_LUT4 \DLX_IFinst__n0003<4>1_G  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(IR[4]),
    .ADR2(DLX_IFinst_IR_previous[4]),
    .ADR3(VCC),
    .O(N165723)
  );
  defparam \DLX_IFinst__n0003<4>1_F .INIT = 16'hDC8C;
  X_LUT4 \DLX_IFinst__n0003<4>1_F  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(IR[4]),
    .ADR2(DLX_IFinst_stalled),
    .ADR3(DLX_IFinst_IR_curr[4]),
    .O(N165721)
  );
  X_MUX2 \DLX_IFinst__n0003<5>1  (
    .IA(N165691),
    .IB(N165693),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[5])
  );
  defparam \DLX_IFinst__n0003<5>1_G .INIT = 16'hCCAA;
  X_LUT4 \DLX_IFinst__n0003<5>1_G  (
    .ADR0(DLX_IFinst_IR_previous[5]),
    .ADR1(IR[5]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_branch_sig),
    .O(N165693)
  );
  defparam \DLX_IFinst__n0003<5>1_F .INIT = 16'hACAA;
  X_LUT4 \DLX_IFinst__n0003<5>1_F  (
    .ADR0(IR[5]),
    .ADR1(DLX_IFinst_IR_curr[5]),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(DLX_IFinst_stalled),
    .O(N165691)
  );
  X_MUX2 \DLX_IFinst__n0003<6>1  (
    .IA(N165701),
    .IB(N165703),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[6])
  );
  defparam \DLX_IFinst__n0003<6>1_G .INIT = 16'hAAF0;
  X_LUT4 \DLX_IFinst__n0003<6>1_G  (
    .ADR0(IR[6]),
    .ADR1(VCC),
    .ADR2(DLX_IFinst_IR_previous[6]),
    .ADR3(DLX_IDinst_branch_sig),
    .O(N165703)
  );
  defparam \DLX_IFinst__n0003<6>1_F .INIT = 16'hAEA2;
  X_LUT4 \DLX_IFinst__n0003<6>1_F  (
    .ADR0(IR[6]),
    .ADR1(DLX_IFinst_stalled),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(DLX_IFinst_IR_curr[6]),
    .O(N165701)
  );
  X_MUX2 \DLX_IFinst__n0003<7>1  (
    .IA(N165796),
    .IB(N165798),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[7])
  );
  defparam \DLX_IFinst__n0003<7>1_G .INIT = 16'hEE44;
  X_LUT4 \DLX_IFinst__n0003<7>1_G  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(DLX_IFinst_IR_previous[7]),
    .ADR2(VCC),
    .ADR3(IR[7]),
    .O(N165798)
  );
  defparam \DLX_IFinst__n0003<7>1_F .INIT = 16'hF4B0;
  X_LUT4 \DLX_IFinst__n0003<7>1_F  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(DLX_IFinst_stalled),
    .ADR2(IR[7]),
    .ADR3(DLX_IFinst_IR_curr[7]),
    .O(N165796)
  );
  X_MUX2 \DLX_IFinst__n0003<8>1  (
    .IA(N165736),
    .IB(N165738),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[8])
  );
  defparam \DLX_IFinst__n0003<8>1_G .INIT = 16'hAFA0;
  X_LUT4 \DLX_IFinst__n0003<8>1_G  (
    .ADR0(IR[8]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(DLX_IFinst_IR_previous[8]),
    .O(N165738)
  );
  defparam \DLX_IFinst__n0003<8>1_F .INIT = 16'hAACA;
  X_LUT4 \DLX_IFinst__n0003<8>1_F  (
    .ADR0(IR[8]),
    .ADR1(DLX_IFinst_IR_curr[8]),
    .ADR2(DLX_IFinst_stalled),
    .ADR3(DLX_IDinst_branch_sig),
    .O(N165736)
  );
  X_MUX2 \DLX_IFinst__n0003<9>1  (
    .IA(N165741),
    .IB(N165743),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[9])
  );
  defparam \DLX_IFinst__n0003<9>1_G .INIT = 16'hEE44;
  X_LUT4 \DLX_IFinst__n0003<9>1_G  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(DLX_IFinst_IR_previous[9]),
    .ADR2(VCC),
    .ADR3(IR[9]),
    .O(N165743)
  );
  defparam \DLX_IFinst__n0003<9>1_F .INIT = 16'hFB40;
  X_LUT4 \DLX_IFinst__n0003<9>1_F  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(DLX_IFinst_stalled),
    .ADR2(DLX_IFinst_IR_curr[9]),
    .ADR3(IR[9]),
    .O(N165741)
  );
  X_MUX2 DLX_IDinst__n0428581 (
    .IA(N165466),
    .IB(N165468),
    .SEL(DLX_IDinst_IR_latched[26]),
    .O(\CHOICE1987/F5MUX )
  );
  defparam DLX_IDinst__n0428581_G.INIT = 16'h31F0;
  X_LUT4 DLX_IDinst__n0428581_G (
    .ADR0(DLX_IDinst_IR_latched[30]),
    .ADR1(DLX_IDinst_IR_latched[27]),
    .ADR2(DLX_IDinst_IR_latched[29]),
    .ADR3(DLX_IDinst_IR_latched[28]),
    .O(N165468)
  );
  defparam DLX_IDinst__n0428581_F.INIT = 16'h7F05;
  X_LUT4 DLX_IDinst__n0428581_F (
    .ADR0(DLX_IDinst_IR_latched[30]),
    .ADR1(DLX_IDinst_IR_latched[28]),
    .ADR2(DLX_IDinst_IR_latched[27]),
    .ADR3(DLX_IDinst_IR_latched[29]),
    .O(N165466)
  );
  X_BUF \CHOICE1987/XUSED  (
    .I(\CHOICE1987/F5MUX ),
    .O(CHOICE1987)
  );
  X_MUX2 DLX_IDinst_Ker1074031 (
    .IA(N165546),
    .IB(N165548),
    .SEL(DLX_IDinst__n0166),
    .O(\DLX_IDinst_N107405/F5MUX )
  );
  defparam DLX_IDinst_Ker1074031_G.INIT = 16'h0313;
  X_LUT4 DLX_IDinst_Ker1074031_G (
    .ADR0(CHOICE1994),
    .ADR1(N135079),
    .ADR2(DLX_IDinst_N108238),
    .ADR3(CHOICE1989),
    .O(N165548)
  );
  defparam DLX_IDinst_Ker1074031_F.INIT = 16'h330A;
  X_LUT4 DLX_IDinst_Ker1074031_F (
    .ADR0(DLX_IDinst__n0434),
    .ADR1(DLX_IDinst__n0433),
    .ADR2(DLX_IDinst__n0436),
    .ADR3(DLX_IDinst__n0167),
    .O(N165546)
  );
  X_BUF \DLX_IDinst_N107405/XUSED  (
    .I(\DLX_IDinst_N107405/F5MUX ),
    .O(DLX_IDinst_N107405)
  );
  X_MUX2 \DLX_EXinst__n0007<19>149_SW01  (
    .IA(N165891),
    .IB(N165893),
    .SEL(DLX_IDinst_IR_opcode_field[0]),
    .O(\N163338/F5MUX )
  );
  defparam \DLX_EXinst__n0007<19>149_SW01_G .INIT = 16'hB080;
  X_LUT4 \DLX_EXinst__n0007<19>149_SW01_G  (
    .ADR0(\DLX_IDinst_Imm[3] ),
    .ADR1(DLX_IDinst_IR_opcode_field[1]),
    .ADR2(DLX_EXinst_N76011),
    .ADR3(\DLX_IDinst_Imm[31] ),
    .O(N165893)
  );
  defparam \DLX_EXinst__n0007<19>149_SW01_F .INIT = 16'h2800;
  X_LUT4 \DLX_EXinst__n0007<19>149_SW01_F  (
    .ADR0(DLX_EXinst_N76011),
    .ADR1(DLX_IDinst_IR_opcode_field[1]),
    .ADR2(DLX_IDinst_reg_out_A[19]),
    .ADR3(\DLX_IDinst_Imm[31] ),
    .O(N165891)
  );
  X_BUF \N163338/XUSED  (
    .I(\N163338/F5MUX ),
    .O(N163338)
  );
  X_MUX2 \DLX_EXinst__n0007<10>2341  (
    .IA(N165706),
    .IB(N165708),
    .SEL(DLX_EXinst__n0036),
    .O(\CHOICE4498/F5MUX )
  );
  defparam \DLX_EXinst__n0007<10>2341_G .INIT = 16'hFEFE;
  X_LUT4 \DLX_EXinst__n0007<10>2341_G  (
    .ADR0(CHOICE4450),
    .ADR1(CHOICE4467),
    .ADR2(CHOICE4445),
    .ADR3(VCC),
    .O(N165708)
  );
  defparam \DLX_EXinst__n0007<10>2341_F .INIT = 16'hFDFC;
  X_LUT4 \DLX_EXinst__n0007<10>2341_F  (
    .ADR0(N146478),
    .ADR1(CHOICE4479),
    .ADR2(CHOICE4495),
    .ADR3(CHOICE4474),
    .O(N165706)
  );
  X_BUF \CHOICE4498/XUSED  (
    .I(\CHOICE4498/F5MUX ),
    .O(CHOICE4498)
  );
  defparam DLX_IDinst_RegFile_28_18_1609.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_28_18_1609 (
    .I(DLX_IDinst_WB_data_eff[18]),
    .CE(DLX_IDinst__n0606),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_28_18)
  );
  X_MUX2 \DLX_EXinst__n0007<11>2341  (
    .IA(N165351),
    .IB(N165353),
    .SEL(DLX_EXinst__n0036),
    .O(\CHOICE4438/F5MUX )
  );
  defparam \DLX_EXinst__n0007<11>2341_G .INIT = 16'hFFEE;
  X_LUT4 \DLX_EXinst__n0007<11>2341_G  (
    .ADR0(CHOICE4385),
    .ADR1(CHOICE4390),
    .ADR2(VCC),
    .ADR3(CHOICE4407),
    .O(N165353)
  );
  defparam \DLX_EXinst__n0007<11>2341_F .INIT = 16'hFCFE;
  X_LUT4 \DLX_EXinst__n0007<11>2341_F  (
    .ADR0(CHOICE4414),
    .ADR1(CHOICE4419),
    .ADR2(CHOICE4435),
    .ADR3(N146478),
    .O(N165351)
  );
  X_BUF \CHOICE4438/XUSED  (
    .I(\CHOICE4438/F5MUX ),
    .O(CHOICE4438)
  );
  X_MUX2 \DLX_EXinst__n0007<12>2261  (
    .IA(N165346),
    .IB(N165348),
    .SEL(DLX_EXinst__n0036),
    .O(\CHOICE3813/F5MUX )
  );
  defparam \DLX_EXinst__n0007<12>2261_G .INIT = 16'hFEEE;
  X_LUT4 \DLX_EXinst__n0007<12>2261_G  (
    .ADR0(CHOICE3766),
    .ADR1(CHOICE3785),
    .ADR2(N134683),
    .ADR3(DLX_IDinst_reg_out_B[4]),
    .O(N165348)
  );
  defparam \DLX_EXinst__n0007<12>2261_F .INIT = 16'hFFEC;
  X_LUT4 \DLX_EXinst__n0007<12>2261_F  (
    .ADR0(CHOICE3793),
    .ADR1(CHOICE3810),
    .ADR2(\DLX_IDinst_Imm[12] ),
    .ADR3(CHOICE3795),
    .O(N165346)
  );
  X_BUF \CHOICE3813/XUSED  (
    .I(\CHOICE3813/F5MUX ),
    .O(CHOICE3813)
  );
  defparam DLX_IDinst_RegFile_29_10_1610.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_29_10_1610 (
    .I(DLX_IDinst_WB_data_eff[10]),
    .CE(DLX_IDinst__n0608),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_29_10)
  );
  X_MUX2 \DLX_EXinst__n0007<13>2261  (
    .IA(N165731),
    .IB(N165733),
    .SEL(DLX_EXinst__n0036),
    .O(\CHOICE3758/F5MUX )
  );
  defparam \DLX_EXinst__n0007<13>2261_G .INIT = 16'hFFF8;
  X_LUT4 \DLX_EXinst__n0007<13>2261_G  (
    .ADR0(N139189),
    .ADR1(DLX_IDinst_reg_out_B[4]),
    .ADR2(CHOICE3711),
    .ADR3(CHOICE3730),
    .O(N165733)
  );
  defparam \DLX_EXinst__n0007<13>2261_F .INIT = 16'hFFEC;
  X_LUT4 \DLX_EXinst__n0007<13>2261_F  (
    .ADR0(CHOICE3738),
    .ADR1(CHOICE3740),
    .ADR2(\DLX_IDinst_Imm[13] ),
    .ADR3(CHOICE3755),
    .O(N165731)
  );
  X_BUF \CHOICE3758/XUSED  (
    .I(\CHOICE3758/F5MUX ),
    .O(CHOICE3758)
  );
  X_MUX2 \DLX_EXinst__n0007<21>1771  (
    .IA(N165561),
    .IB(N165563),
    .SEL(DLX_IDinst_reg_out_B[2]),
    .O(\DLX_IDinst_RegFile_3_12/F5MUX )
  );
  defparam \DLX_EXinst__n0007<21>1771_G .INIT = 16'h44F0;
  X_LUT4 \DLX_EXinst__n0007<21>1771_G  (
    .ADR0(DLX_IDinst_reg_out_B[3]),
    .ADR1(\DLX_EXinst_Mshift__n0023_Sh[1] ),
    .ADR2(DLX_EXinst_N73848),
    .ADR3(DLX_IDinst_reg_out_B[4]),
    .O(N165563)
  );
  defparam \DLX_EXinst__n0007<21>1771_F .INIT = 16'h0ACA;
  X_LUT4 \DLX_EXinst__n0007<21>1771_F  (
    .ADR0(DLX_EXinst_N74024),
    .ADR1(\DLX_EXinst_Mshift__n0023_Sh[5] ),
    .ADR2(DLX_IDinst_reg_out_B[4]),
    .ADR3(DLX_IDinst_reg_out_B[3]),
    .O(N165561)
  );
  X_BUF \DLX_IDinst_RegFile_3_12/XUSED  (
    .I(\DLX_IDinst_RegFile_3_12/F5MUX ),
    .O(CHOICE4167)
  );
  X_MUX2 \DLX_EXinst__n0007<30>2211  (
    .IA(N165441),
    .IB(N165443),
    .SEL(DLX_IDinst_reg_out_B[4]),
    .O(\CHOICE4754/F5MUX )
  );
  defparam \DLX_EXinst__n0007<30>2211_G .INIT = 16'h80A2;
  X_LUT4 \DLX_EXinst__n0007<30>2211_G  (
    .ADR0(DLX_EXinst_N76338),
    .ADR1(DLX_IDinst_reg_out_B[3]),
    .ADR2(DLX_EXinst_N72908),
    .ADR3(N130105),
    .O(N165443)
  );
  defparam \DLX_EXinst__n0007<30>2211_F .INIT = 16'h88C0;
  X_LUT4 \DLX_EXinst__n0007<30>2211_F  (
    .ADR0(N133120),
    .ADR1(DLX_EXinst_N76338),
    .ADR2(CHOICE4748),
    .ADR3(DLX_IDinst_reg_out_B[2]),
    .O(N165441)
  );
  X_BUF \CHOICE4754/XUSED  (
    .I(\CHOICE4754/F5MUX ),
    .O(CHOICE4754)
  );
  X_MUX2 \DLX_EXinst__n0007<14>2261  (
    .IA(N165696),
    .IB(N165698),
    .SEL(DLX_EXinst__n0036),
    .O(\CHOICE3703/F5MUX )
  );
  defparam \DLX_EXinst__n0007<14>2261_G .INIT = 16'hFFF8;
  X_LUT4 \DLX_EXinst__n0007<14>2261_G  (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(N139297),
    .ADR2(CHOICE3656),
    .ADR3(CHOICE3675),
    .O(N165698)
  );
  defparam \DLX_EXinst__n0007<14>2261_F .INIT = 16'hFEFA;
  X_LUT4 \DLX_EXinst__n0007<14>2261_F  (
    .ADR0(CHOICE3685),
    .ADR1(\DLX_IDinst_Imm[14] ),
    .ADR2(CHOICE3700),
    .ADR3(CHOICE3683),
    .O(N165696)
  );
  X_BUF \CHOICE3703/XUSED  (
    .I(\CHOICE3703/F5MUX ),
    .O(CHOICE3703)
  );
  X_MUX2 \DLX_EXinst__n0007<22>1771  (
    .IA(N165391),
    .IB(N165393),
    .SEL(DLX_IDinst_reg_out_B[2]),
    .O(\CHOICE4102/F5MUX )
  );
  defparam \DLX_EXinst__n0007<22>1771_G .INIT = 16'h7430;
  X_LUT4 \DLX_EXinst__n0007<22>1771_G  (
    .ADR0(DLX_IDinst_reg_out_B[3]),
    .ADR1(DLX_IDinst_reg_out_B[4]),
    .ADR2(DLX_EXinst_N73853),
    .ADR3(\DLX_EXinst_Mshift__n0023_Sh[2] ),
    .O(N165393)
  );
  defparam \DLX_EXinst__n0007<22>1771_F .INIT = 16'h50CC;
  X_LUT4 \DLX_EXinst__n0007<22>1771_F  (
    .ADR0(DLX_IDinst_reg_out_B[3]),
    .ADR1(DLX_EXinst_N74029),
    .ADR2(\DLX_EXinst_Mshift__n0023_Sh[6] ),
    .ADR3(DLX_IDinst_reg_out_B[4]),
    .O(N165391)
  );
  X_BUF \CHOICE4102/XUSED  (
    .I(\CHOICE4102/F5MUX ),
    .O(CHOICE4102)
  );
  X_MUX2 \DLX_EXinst__n0007<31>4111  (
    .IA(N165816),
    .IB(N165818),
    .SEL(\DLX_IDinst_Imm[4] ),
    .O(\CHOICE5838/F5MUX )
  );
  defparam \DLX_EXinst__n0007<31>4111_G .INIT = 16'hC480;
  X_LUT4 \DLX_EXinst__n0007<31>4111_G  (
    .ADR0(\DLX_IDinst_Imm[3] ),
    .ADR1(DLX_EXinst__n0055),
    .ADR2(DLX_EXinst_N72998),
    .ADR3(N130415),
    .O(N165818)
  );
  defparam \DLX_EXinst__n0007<31>4111_F .INIT = 16'hC088;
  X_LUT4 \DLX_EXinst__n0007<31>4111_F  (
    .ADR0(N163186),
    .ADR1(DLX_EXinst__n0055),
    .ADR2(N137282),
    .ADR3(\DLX_IDinst_Imm[2] ),
    .O(N165816)
  );
  X_BUF \CHOICE5838/XUSED  (
    .I(\CHOICE5838/F5MUX ),
    .O(CHOICE5838)
  );
  X_MUX2 \DLX_EXinst__n0007<23>1771  (
    .IA(N165461),
    .IB(N165463),
    .SEL(DLX_IDinst_reg_out_B[2]),
    .O(\CHOICE4037/F5MUX )
  );
  defparam \DLX_EXinst__n0007<23>1771_G .INIT = 16'h7520;
  X_LUT4 \DLX_EXinst__n0007<23>1771_G  (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(DLX_IDinst_reg_out_B[3]),
    .ADR2(\DLX_EXinst_Mshift__n0023_Sh[3] ),
    .ADR3(DLX_EXinst_N73858),
    .O(N165463)
  );
  defparam \DLX_EXinst__n0007<23>1771_F .INIT = 16'h7520;
  X_LUT4 \DLX_EXinst__n0007<23>1771_F  (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(DLX_IDinst_reg_out_B[3]),
    .ADR2(\DLX_EXinst_Mshift__n0023_Sh[7] ),
    .ADR3(DLX_EXinst_N74034),
    .O(N165461)
  );
  X_BUF \CHOICE4037/XUSED  (
    .I(\CHOICE4037/F5MUX ),
    .O(CHOICE4037)
  );
  X_MUX2 \DLX_EXinst__n0007<31>5251  (
    .IA(N165711),
    .IB(N165713),
    .SEL(DLX_IDinst_reg_out_A[31]),
    .O(\CHOICE5864/F5MUX )
  );
  defparam \DLX_EXinst__n0007<31>5251_G .INIT = 16'hFEEE;
  X_LUT4 \DLX_EXinst__n0007<31>5251_G  (
    .ADR0(CHOICE5861),
    .ADR1(DLX_EXinst__n0053),
    .ADR2(\DLX_IDinst_Imm[31] ),
    .ADR3(DLX_EXinst__n0052),
    .O(N165713)
  );
  defparam \DLX_EXinst__n0007<31>5251_F .INIT = 16'h6000;
  X_LUT4 \DLX_EXinst__n0007<31>5251_F  (
    .ADR0(DLX_IDinst_IR_opcode_field[0]),
    .ADR1(DLX_IDinst_IR_opcode_field[1]),
    .ADR2(DLX_EXinst_N76011),
    .ADR3(\DLX_IDinst_Imm[31] ),
    .O(N165711)
  );
  X_BUF \CHOICE5864/XUSED  (
    .I(\CHOICE5864/F5MUX ),
    .O(CHOICE5864)
  );
  X_MUX2 \DLX_EXinst__n0007<16>2141  (
    .IA(N165666),
    .IB(N165668),
    .SEL(\DLX_IDinst_Imm[2] ),
    .O(\CHOICE4608/F5MUX )
  );
  defparam \DLX_EXinst__n0007<16>2141_G .INIT = 16'h3210;
  X_LUT4 \DLX_EXinst__n0007<16>2141_G  (
    .ADR0(\DLX_IDinst_Imm[3] ),
    .ADR1(\DLX_IDinst_Imm[4] ),
    .ADR2(\DLX_EXinst_Mshift__n0021_Sh[12] ),
    .ADR3(\DLX_EXinst_Mshift__n0021_Sh[4] ),
    .O(N165668)
  );
  defparam \DLX_EXinst__n0007<16>2141_F .INIT = 16'h00E4;
  X_LUT4 \DLX_EXinst__n0007<16>2141_F  (
    .ADR0(\DLX_IDinst_Imm[3] ),
    .ADR1(\DLX_EXinst_Mshift__n0021_Sh[16] ),
    .ADR2(\DLX_EXinst_Mshift__n0021_Sh[8] ),
    .ADR3(\DLX_IDinst_Imm[4] ),
    .O(N165666)
  );
  X_BUF \CHOICE4608/XUSED  (
    .I(\CHOICE4608/F5MUX ),
    .O(CHOICE4608)
  );
  X_MUX2 \DLX_EXinst__n0007<16>2941  (
    .IA(N165756),
    .IB(N165758),
    .SEL(DLX_IDinst_IR_opcode_field[0]),
    .O(\DLX_IDinst_RegFile_2_31/F5MUX )
  );
  defparam \DLX_EXinst__n0007<16>2941_G .INIT = 16'hD800;
  X_LUT4 \DLX_EXinst__n0007<16>2941_G  (
    .ADR0(DLX_IDinst_IR_opcode_field[1]),
    .ADR1(\DLX_IDinst_Imm[0] ),
    .ADR2(\DLX_IDinst_Imm[31] ),
    .ADR3(DLX_EXinst_N76011),
    .O(N165758)
  );
  defparam \DLX_EXinst__n0007<16>2941_F .INIT = 16'h4080;
  X_LUT4 \DLX_EXinst__n0007<16>2941_F  (
    .ADR0(DLX_IDinst_reg_out_A[16]),
    .ADR1(\DLX_IDinst_Imm[31] ),
    .ADR2(DLX_EXinst_N76011),
    .ADR3(DLX_IDinst_IR_opcode_field[1]),
    .O(N165756)
  );
  X_BUF \DLX_IDinst_RegFile_2_31/XUSED  (
    .I(\DLX_IDinst_RegFile_2_31/F5MUX ),
    .O(CHOICE4624)
  );
  X_MUX2 \DLX_EXinst__n0007<24>2951  (
    .IA(N165826),
    .IB(N165828),
    .SEL(\DLX_IDinst_Imm[5] ),
    .O(\CHOICE5648/F5MUX )
  );
  defparam \DLX_EXinst__n0007<24>2951_G .INIT = 16'h0020;
  X_LUT4 \DLX_EXinst__n0007<24>2951_G  (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(\DLX_IDinst_Imm[4] ),
    .ADR2(N147520),
    .ADR3(\DLX_IDinst_Imm[3] ),
    .O(N165828)
  );
  defparam \DLX_EXinst__n0007<24>2951_F .INIT = 16'hC808;
  X_LUT4 \DLX_EXinst__n0007<24>2951_F  (
    .ADR0(\DLX_EXinst_Mshift__n0020_Sh[88] ),
    .ADR1(N147520),
    .ADR2(\DLX_IDinst_Imm[4] ),
    .ADR3(DLX_IDinst_reg_out_A[31]),
    .O(N165826)
  );
  X_BUF \CHOICE5648/XUSED  (
    .I(\CHOICE5648/F5MUX ),
    .O(CHOICE5648)
  );
  X_MUX2 \DLX_EXinst__n0007<17>2631  (
    .IA(N165536),
    .IB(N165538),
    .SEL(DLX_IDinst_reg_out_B[3]),
    .O(\DLX_IFinst_IR_previous<21>/F5MUX )
  );
  defparam \DLX_EXinst__n0007<17>2631_G .INIT = 16'hB080;
  X_LUT4 \DLX_EXinst__n0007<17>2631_G  (
    .ADR0(\DLX_EXinst_Mshift__n0023_Sh[5] ),
    .ADR1(DLX_IDinst_reg_out_B[2]),
    .ADR2(DLX_EXinst__n0080),
    .ADR3(\DLX_EXinst_Mshift__n0023_Sh[9] ),
    .O(N165538)
  );
  defparam \DLX_EXinst__n0007<17>2631_F .INIT = 16'hC840;
  X_LUT4 \DLX_EXinst__n0007<17>2631_F  (
    .ADR0(DLX_IDinst_reg_out_B[2]),
    .ADR1(DLX_EXinst__n0080),
    .ADR2(N129951),
    .ADR3(\DLX_EXinst_Mshift__n0023_Sh[13] ),
    .O(N165536)
  );
  X_BUF \DLX_IFinst_IR_previous<21>/XUSED  (
    .I(\DLX_IFinst_IR_previous<21>/F5MUX ),
    .O(CHOICE5416)
  );
  defparam DLX_IDinst_RegFile_28_27_1611.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_28_27_1611 (
    .I(DLX_IDinst_WB_data_eff[27]),
    .CE(DLX_IDinst__n0606),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_28_27)
  );
  X_MUX2 \DLX_EXinst__n0007<18>2631  (
    .IA(N165566),
    .IB(N165568),
    .SEL(DLX_IDinst_reg_out_B[3]),
    .O(\CHOICE5258/F5MUX )
  );
  defparam \DLX_EXinst__n0007<18>2631_G .INIT = 16'h8C80;
  X_LUT4 \DLX_EXinst__n0007<18>2631_G  (
    .ADR0(\DLX_EXinst_Mshift__n0023_Sh[6] ),
    .ADR1(DLX_EXinst__n0080),
    .ADR2(DLX_IDinst_reg_out_B[2]),
    .ADR3(\DLX_EXinst_Mshift__n0023_Sh[10] ),
    .O(N165568)
  );
  defparam \DLX_EXinst__n0007<18>2631_F .INIT = 16'hC480;
  X_LUT4 \DLX_EXinst__n0007<18>2631_F  (
    .ADR0(DLX_IDinst_reg_out_B[2]),
    .ADR1(DLX_EXinst__n0080),
    .ADR2(\DLX_EXinst_Mshift__n0023_Sh[14] ),
    .ADR3(N130001),
    .O(N165566)
  );
  X_BUF \CHOICE5258/XUSED  (
    .I(\CHOICE5258/F5MUX ),
    .O(CHOICE5258)
  );
  X_MUX2 \DLX_EXinst__n0007<19>2631  (
    .IA(N165596),
    .IB(N165598),
    .SEL(DLX_IDinst_reg_out_B[3]),
    .O(\DLX_IDinst_RegFile_1_4/F5MUX )
  );
  defparam \DLX_EXinst__n0007<19>2631_G .INIT = 16'hC480;
  X_LUT4 \DLX_EXinst__n0007<19>2631_G  (
    .ADR0(DLX_IDinst_reg_out_B[2]),
    .ADR1(DLX_EXinst__n0080),
    .ADR2(\DLX_EXinst_Mshift__n0023_Sh[7] ),
    .ADR3(\DLX_EXinst_Mshift__n0023_Sh[11] ),
    .O(N165598)
  );
  defparam \DLX_EXinst__n0007<19>2631_F .INIT = 16'hC840;
  X_LUT4 \DLX_EXinst__n0007<19>2631_F  (
    .ADR0(DLX_IDinst_reg_out_B[2]),
    .ADR1(DLX_EXinst__n0080),
    .ADR2(\DLX_EXinst_Mshift__n0023_Sh[19] ),
    .ADR3(\DLX_EXinst_Mshift__n0023_Sh[15] ),
    .O(N165596)
  );
  X_BUF \DLX_IDinst_RegFile_1_4/XUSED  (
    .I(\DLX_IDinst_RegFile_1_4/F5MUX ),
    .O(CHOICE5337)
  );
  X_MUX2 \DLX_EXinst__n0007<28>1191  (
    .IA(N165861),
    .IB(N165863),
    .SEL(DLX_IDinst_IR_opcode_field[0]),
    .O(\CHOICE4874/F5MUX )
  );
  defparam \DLX_EXinst__n0007<28>1191_G .INIT = 16'hC840;
  X_LUT4 \DLX_EXinst__n0007<28>1191_G  (
    .ADR0(DLX_IDinst_IR_opcode_field[1]),
    .ADR1(DLX_EXinst_N76011),
    .ADR2(\DLX_IDinst_Imm[31] ),
    .ADR3(\DLX_IDinst_Imm[12] ),
    .O(N165863)
  );
  defparam \DLX_EXinst__n0007<28>1191_F .INIT = 16'h2800;
  X_LUT4 \DLX_EXinst__n0007<28>1191_F  (
    .ADR0(DLX_EXinst_N76011),
    .ADR1(DLX_IDinst_reg_out_A[28]),
    .ADR2(DLX_IDinst_IR_opcode_field[1]),
    .ADR3(\DLX_IDinst_Imm[31] ),
    .O(N165861)
  );
  X_BUF \CHOICE4874/XUSED  (
    .I(\CHOICE4874/F5MUX ),
    .O(CHOICE4874)
  );
  X_MUX2 \DLX_EXinst__n0007<28>2691  (
    .IA(N165581),
    .IB(N165583),
    .SEL(DLX_IDinst_reg_out_B[4]),
    .O(\DLX_IDinst_RegFile_10_0/F5MUX )
  );
  defparam \DLX_EXinst__n0007<28>2691_G .INIT = 16'hAC00;
  X_LUT4 \DLX_EXinst__n0007<28>2691_G  (
    .ADR0(DLX_EXinst_N72898),
    .ADR1(DLX_EXinst_N74051),
    .ADR2(DLX_IDinst_reg_out_B[3]),
    .ADR3(DLX_EXinst_N76338),
    .O(N165583)
  );
  defparam \DLX_EXinst__n0007<28>2691_F .INIT = 16'h8C80;
  X_LUT4 \DLX_EXinst__n0007<28>2691_F  (
    .ADR0(DLX_EXinst_N75006),
    .ADR1(DLX_EXinst_N76338),
    .ADR2(DLX_IDinst_reg_out_B[3]),
    .ADR3(CHOICE4896),
    .O(N165581)
  );
  X_BUF \DLX_IDinst_RegFile_10_0/XUSED  (
    .I(\DLX_IDinst_RegFile_10_0/F5MUX ),
    .O(CHOICE4902)
  );
  X_MUX2 \DLX_EXinst__n0007<29>2211  (
    .IA(N165481),
    .IB(N165483),
    .SEL(DLX_IDinst_reg_out_B[4]),
    .O(\CHOICE4825/F5MUX )
  );
  defparam \DLX_EXinst__n0007<29>2211_G .INIT = 16'h8D00;
  X_LUT4 \DLX_EXinst__n0007<29>2211_G  (
    .ADR0(DLX_IDinst_reg_out_B[3]),
    .ADR1(DLX_EXinst_N72903),
    .ADR2(N130051),
    .ADR3(DLX_EXinst_N76338),
    .O(N165483)
  );
  defparam \DLX_EXinst__n0007<29>2211_F .INIT = 16'hE400;
  X_LUT4 \DLX_EXinst__n0007<29>2211_F  (
    .ADR0(DLX_IDinst_reg_out_B[2]),
    .ADR1(CHOICE4819),
    .ADR2(N133048),
    .ADR3(DLX_EXinst_N76338),
    .O(N165481)
  );
  X_BUF \CHOICE4825/XUSED  (
    .I(\CHOICE4825/F5MUX ),
    .O(CHOICE4825)
  );
  X_MUX2 \DLX_EXinst__n0007<5>25511  (
    .IA(N165876),
    .IB(N165878),
    .SEL(DLX_EXinst__n0036),
    .O(\DLX_EXinst_ALU_result_5_1/F5MUX )
  );
  defparam \DLX_EXinst__n0007<5>25511_G .INIT = 16'hFAF0;
  X_LUT4 \DLX_EXinst__n0007<5>25511_G  (
    .ADR0(DLX_EXinst__n0012[5]),
    .ADR1(VCC),
    .ADR2(N163182),
    .ADR3(DLX_EXinst__n0127),
    .O(N165878)
  );
  defparam \DLX_EXinst__n0007<5>25511_F .INIT = 16'hFFF8;
  X_LUT4 \DLX_EXinst__n0007<5>25511_F  (
    .ADR0(DLX_EXinst__n0109),
    .ADR1(DLX_EXinst__n0012[5]),
    .ADR2(CHOICE3971),
    .ADR3(CHOICE3987),
    .O(N165876)
  );
  X_BUF \DLX_EXinst_ALU_result_5_1/XUSED  (
    .I(\DLX_EXinst_ALU_result_5_1/F5MUX ),
    .O(N162863)
  );
  X_MUX2 \DLX_EXinst__n0007<6>25511  (
    .IA(N165841),
    .IB(N165843),
    .SEL(DLX_EXinst__n0036),
    .O(\DLX_EXinst_ALU_result_6_1/F5MUX )
  );
  defparam \DLX_EXinst__n0007<6>25511_G .INIT = 16'hFFA0;
  X_LUT4 \DLX_EXinst__n0007<6>25511_G  (
    .ADR0(DLX_EXinst__n0012[6]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst__n0127),
    .ADR3(N163198),
    .O(N165843)
  );
  defparam \DLX_EXinst__n0007<6>25511_F .INIT = 16'hFFEC;
  X_LUT4 \DLX_EXinst__n0007<6>25511_F  (
    .ADR0(DLX_EXinst__n0012[6]),
    .ADR1(CHOICE3912),
    .ADR2(DLX_EXinst__n0109),
    .ADR3(CHOICE3928),
    .O(N165841)
  );
  X_BUF \DLX_EXinst_ALU_result_6_1/XUSED  (
    .I(\DLX_EXinst_ALU_result_6_1/F5MUX ),
    .O(N162801)
  );
  X_MUX2 \DLX_EXinst__n0007<7>25511  (
    .IA(N165801),
    .IB(N165803),
    .SEL(DLX_EXinst__n0036),
    .O(\DLX_EXinst_ALU_result_7_1/F5MUX )
  );
  defparam \DLX_EXinst__n0007<7>25511_G .INIT = 16'hEECC;
  X_LUT4 \DLX_EXinst__n0007<7>25511_G  (
    .ADR0(DLX_EXinst__n0012[7]),
    .ADR1(N163226),
    .ADR2(VCC),
    .ADR3(DLX_EXinst__n0127),
    .O(N165803)
  );
  defparam \DLX_EXinst__n0007<7>25511_F .INIT = 16'hFFF8;
  X_LUT4 \DLX_EXinst__n0007<7>25511_F  (
    .ADR0(DLX_EXinst__n0012[7]),
    .ADR1(DLX_EXinst__n0109),
    .ADR2(CHOICE3869),
    .ADR3(CHOICE3853),
    .O(N165801)
  );
  X_BUF \DLX_EXinst_ALU_result_7_1/XUSED  (
    .I(\DLX_EXinst_ALU_result_7_1/F5MUX ),
    .O(N162807)
  );
  X_MUX2 DLX_EXinst_Ker74226291 (
    .IA(N165436),
    .IB(N165438),
    .SEL(DLX_IDinst_reg_out_B[1]),
    .O(\CHOICE1765/F5MUX )
  );
  defparam DLX_EXinst_Ker74226291_G.INIT = 16'h3202;
  X_LUT4 DLX_EXinst_Ker74226291_G (
    .ADR0(DLX_IDinst_reg_out_A[25]),
    .ADR1(DLX_IDinst_reg_out_B[3]),
    .ADR2(DLX_IDinst_reg_out_B[0]),
    .ADR3(DLX_IDinst_reg_out_A[24]),
    .O(N165438)
  );
  defparam DLX_EXinst_Ker74226291_F.INIT = 16'h4540;
  X_LUT4 DLX_EXinst_Ker74226291_F (
    .ADR0(DLX_IDinst_reg_out_B[3]),
    .ADR1(DLX_IDinst_reg_out_A[26]),
    .ADR2(DLX_IDinst_reg_out_B[0]),
    .ADR3(DLX_IDinst_reg_out_A[27]),
    .O(N165436)
  );
  X_BUF \CHOICE1765/XUSED  (
    .I(\CHOICE1765/F5MUX ),
    .O(CHOICE1765)
  );
  X_MUX2 DLX_EXinst_Ker75142361 (
    .IA(N165626),
    .IB(N165628),
    .SEL(DLX_IDinst_reg_out_B[5]),
    .O(\DLX_IDinst_RegFile_30_10/F5MUX )
  );
  defparam DLX_EXinst_Ker75142361_G.INIT = 16'h2AAA;
  X_LUT4 DLX_EXinst_Ker75142361_G (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(DLX_IDinst_reg_out_B_2_1),
    .ADR2(DLX_IDinst_reg_out_B_3_1),
    .ADR3(DLX_IDinst_reg_out_B[1]),
    .O(N165628)
  );
  defparam DLX_EXinst_Ker75142361_F.INIT = 16'hF5A0;
  X_LUT4 DLX_EXinst_Ker75142361_F (
    .ADR0(DLX_IDinst_reg_out_B_2_1),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N73088),
    .ADR3(DLX_EXinst_N74731),
    .O(N165626)
  );
  X_BUF \DLX_IDinst_RegFile_30_10/XUSED  (
    .I(\DLX_IDinst_RegFile_30_10/F5MUX ),
    .O(N137372)
  );
  X_MUX2 DLX_EXinst_Ker74454481 (
    .IA(N165486),
    .IB(N165488),
    .SEL(DLX_IDinst_reg_out_B[5]),
    .O(\N137952/F5MUX )
  );
  defparam DLX_EXinst_Ker74454481_G.INIT = 16'h00EC;
  X_LUT4 DLX_EXinst_Ker74454481_G (
    .ADR0(\DLX_EXinst_Mshift__n0024_Sh[31] ),
    .ADR1(CHOICE1830),
    .ADR2(DLX_IDinst_reg_out_B_2_1),
    .ADR3(DLX_IDinst_reg_out_B_3_1),
    .O(N165488)
  );
  defparam DLX_EXinst_Ker74454481_F.INIT = 16'hFE22;
  X_LUT4 DLX_EXinst_Ker74454481_F (
    .ADR0(CHOICE1830),
    .ADR1(DLX_IDinst_reg_out_B_3_1),
    .ADR2(DLX_IDinst_reg_out_B_2_1),
    .ADR3(DLX_IDinst_reg_out_A[31]),
    .O(N165486)
  );
  X_BUF \N137952/XUSED  (
    .I(\N137952/F5MUX ),
    .O(N137952)
  );
  X_MUX2 DLX_EXinst_Ker75335361 (
    .IA(N165476),
    .IB(N165478),
    .SEL(\DLX_IDinst_Imm[5] ),
    .O(\DLX_IFinst_IR_previous<24>/F5MUX )
  );
  defparam DLX_EXinst_Ker75335361_G.INIT = 16'h7F00;
  X_LUT4 DLX_EXinst_Ker75335361_G (
    .ADR0(DLX_IDinst_Imm_3_1),
    .ADR1(DLX_IDinst_Imm_1_1),
    .ADR2(DLX_IDinst_Imm_2_1),
    .ADR3(DLX_IDinst_reg_out_A[31]),
    .O(N165478)
  );
  defparam DLX_EXinst_Ker75335361_F.INIT = 16'hD8D8;
  X_LUT4 DLX_EXinst_Ker75335361_F (
    .ADR0(DLX_IDinst_Imm_2_1),
    .ADR1(DLX_EXinst_N73018),
    .ADR2(DLX_EXinst_N74986),
    .ADR3(VCC),
    .O(N165476)
  );
  X_BUF \DLX_IFinst_IR_previous<24>/XUSED  (
    .I(\DLX_IFinst_IR_previous<24>/F5MUX ),
    .O(N137608)
  );
  X_MUX2 DLX_EXinst_Ker75503281 (
    .IA(N165376),
    .IB(N165378),
    .SEL(DLX_IDinst_Imm_3_1),
    .O(\N134488/F5MUX )
  );
  defparam DLX_EXinst_Ker75503281_G.INIT = 16'hCCAA;
  X_LUT4 DLX_EXinst_Ker75503281_G (
    .ADR0(DLX_EXinst_N73128),
    .ADR1(DLX_EXinst_N73524),
    .ADR2(VCC),
    .ADR3(\DLX_IDinst_Imm[0] ),
    .O(N165378)
  );
  defparam DLX_EXinst_Ker75503281_F.INIT = 16'hAACC;
  X_LUT4 DLX_EXinst_Ker75503281_F (
    .ADR0(DLX_EXinst_N73549),
    .ADR1(DLX_EXinst_N73108),
    .ADR2(VCC),
    .ADR3(\DLX_IDinst_Imm[0] ),
    .O(N165376)
  );
  X_BUF \N134488/XUSED  (
    .I(\N134488/F5MUX ),
    .O(N134488)
  );
  X_MUX2 DLX_EXinst_Ker74367531 (
    .IA(N165931),
    .IB(N165933),
    .SEL(DLX_IDinst_reg_out_B[5]),
    .O(\DLX_IDinst_RegFile_2_20/F5MUX )
  );
  defparam DLX_EXinst_Ker74367531_G.INIT = 16'h5C0C;
  X_LUT4 DLX_EXinst_Ker74367531_G (
    .ADR0(DLX_IDinst_reg_out_B[2]),
    .ADR1(DLX_IDinst_reg_out_A[31]),
    .ADR2(DLX_IDinst_reg_out_B[3]),
    .ADR3(\DLX_EXinst_Mshift__n0019_Sh[61] ),
    .O(N165933)
  );
  defparam DLX_EXinst_Ker74367531_F.INIT = 16'hDDCC;
  X_LUT4 DLX_EXinst_Ker74367531_F (
    .ADR0(DLX_IDinst_reg_out_B[2]),
    .ADR1(CHOICE3026),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N73083),
    .O(N165931)
  );
  X_BUF \DLX_IDinst_RegFile_2_20/XUSED  (
    .I(\DLX_IDinst_RegFile_2_20/F5MUX ),
    .O(CHOICE3036)
  );
  X_MUX2 DLX_EXinst_Ker75167391 (
    .IA(N165556),
    .IB(N165558),
    .SEL(DLX_IDinst_reg_out_B[5]),
    .O(\N137859/F5MUX )
  );
  defparam DLX_EXinst_Ker75167391_G.INIT = 16'hDF80;
  X_LUT4 DLX_EXinst_Ker75167391_G (
    .ADR0(DLX_IDinst_reg_out_B_3_1),
    .ADR1(\DLX_EXinst_Mshift__n0019_Sh[61] ),
    .ADR2(DLX_IDinst_reg_out_B_2_1),
    .ADR3(DLX_IDinst_reg_out_A[31]),
    .O(N165558)
  );
  defparam DLX_EXinst_Ker75167391_F.INIT = 16'hCFC0;
  X_LUT4 DLX_EXinst_Ker75167391_F (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N73083),
    .ADR2(DLX_IDinst_reg_out_B_2_1),
    .ADR3(DLX_EXinst_N74726),
    .O(N165556)
  );
  X_BUF \N137859/XUSED  (
    .I(\N137859/F5MUX ),
    .O(N137859)
  );
  X_MUX2 DLX_EXinst_Ker75360281 (
    .IA(N165501),
    .IB(N165503),
    .SEL(DLX_IDinst_reg_out_B[0]),
    .O(\DLX_IDinst_RegFile_26_0/F5MUX )
  );
  defparam DLX_EXinst_Ker75360281_G.INIT = 16'hBB88;
  X_LUT4 DLX_EXinst_Ker75360281_G (
    .ADR0(DLX_EXinst_N73048),
    .ADR1(DLX_IDinst_reg_out_B_3_1),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N73028),
    .O(N165503)
  );
  defparam DLX_EXinst_Ker75360281_F.INIT = 16'hACAC;
  X_LUT4 DLX_EXinst_Ker75360281_F (
    .ADR0(DLX_EXinst_N73394),
    .ADR1(DLX_EXinst_N73424),
    .ADR2(DLX_IDinst_reg_out_B_3_1),
    .ADR3(VCC),
    .O(N165501)
  );
  X_BUF \DLX_IDinst_RegFile_26_0/XUSED  (
    .I(\DLX_IDinst_RegFile_26_0/F5MUX ),
    .O(N133408)
  );
  X_MUX2 DLX_EXinst_Ker75345391 (
    .IA(N165656),
    .IB(N165658),
    .SEL(\DLX_IDinst_Imm[5] ),
    .O(\N138037/F5MUX )
  );
  defparam DLX_EXinst_Ker75345391_G.INIT = 16'hEC4C;
  X_LUT4 DLX_EXinst_Ker75345391_G (
    .ADR0(DLX_IDinst_Imm_3_1),
    .ADR1(DLX_IDinst_reg_out_A[31]),
    .ADR2(DLX_IDinst_Imm_2_1),
    .ADR3(\DLX_EXinst_Mshift__n0020_Sh[61] ),
    .O(N165658)
  );
  defparam DLX_EXinst_Ker75345391_F.INIT = 16'hFC0C;
  X_LUT4 DLX_EXinst_Ker75345391_F (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N74981),
    .ADR2(DLX_IDinst_Imm_2_1),
    .ADR3(DLX_EXinst_N73013),
    .O(N165656)
  );
  X_BUF \N138037/XUSED  (
    .I(\N138037/F5MUX ),
    .O(N138037)
  );
  X_MUX2 DLX_EXinst_Ker75370281 (
    .IA(N165506),
    .IB(N165508),
    .SEL(DLX_IDinst_Imm_3_1),
    .O(\DLX_IDinst_RegFile_17_7/F5MUX )
  );
  defparam DLX_EXinst_Ker75370281_G.INIT = 16'hEE22;
  X_LUT4 DLX_EXinst_Ker75370281_G (
    .ADR0(DLX_EXinst_N72958),
    .ADR1(\DLX_IDinst_Imm[0] ),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N73479),
    .O(N165508)
  );
  defparam DLX_EXinst_Ker75370281_F.INIT = 16'hF3C0;
  X_LUT4 DLX_EXinst_Ker75370281_F (
    .ADR0(VCC),
    .ADR1(\DLX_IDinst_Imm[0] ),
    .ADR2(DLX_EXinst_N73499),
    .ADR3(DLX_EXinst_N72978),
    .O(N165506)
  );
  X_BUF \DLX_IDinst_RegFile_17_7/XUSED  (
    .I(\DLX_IDinst_RegFile_17_7/F5MUX ),
    .O(N133768)
  );
  X_MUX2 DLX_EXinst_Ker74714461 (
    .IA(N165956),
    .IB(N165958),
    .SEL(\DLX_IDinst_Imm[5] ),
    .O(\N137774/F5MUX )
  );
  defparam DLX_EXinst_Ker74714461_G.INIT = 16'h0222;
  X_LUT4 DLX_EXinst_Ker74714461_G (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(DLX_IDinst_Imm_3_1),
    .ADR2(DLX_IDinst_Imm_2_1),
    .ADR3(DLX_EXinst_N73211),
    .O(N165958)
  );
  defparam DLX_EXinst_Ker74714461_F.INIT = 16'hAAB8;
  X_LUT4 DLX_EXinst_Ker74714461_F (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(DLX_IDinst_Imm_3_1),
    .ADR2(\DLX_EXinst_Mshift__n0020_Sh[27] ),
    .ADR3(DLX_IDinst_Imm_2_1),
    .O(N165956)
  );
  X_BUF \N137774/XUSED  (
    .I(\N137774/F5MUX ),
    .O(N137774)
  );
  X_MUX2 DLX_EXinst_Ker75355281 (
    .IA(N165541),
    .IB(N165543),
    .SEL(DLX_IDinst_reg_out_B[0]),
    .O(\DLX_IDinst_RegFile_10_3/F5MUX )
  );
  defparam DLX_EXinst_Ker75355281_G.INIT = 16'hB8B8;
  X_LUT4 DLX_EXinst_Ker75355281_G (
    .ADR0(DLX_EXinst_N73394),
    .ADR1(DLX_IDinst_reg_out_B_3_1),
    .ADR2(DLX_EXinst_N73424),
    .ADR3(VCC),
    .O(N165543)
  );
  defparam DLX_EXinst_Ker75355281_F.INIT = 16'hF5A0;
  X_LUT4 DLX_EXinst_Ker75355281_F (
    .ADR0(DLX_IDinst_reg_out_B_3_1),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N73043),
    .ADR3(DLX_EXinst_N73023),
    .O(N165541)
  );
  X_BUF \DLX_IDinst_RegFile_10_3/XUSED  (
    .I(\DLX_IDinst_RegFile_10_3/F5MUX ),
    .O(N133480)
  );
  X_MUX2 DLX_EXinst_Ker74459291 (
    .IA(N165406),
    .IB(N165408),
    .SEL(DLX_IDinst_Imm_1_1),
    .O(\CHOICE1727/F5MUX )
  );
  defparam DLX_EXinst_Ker74459291_G.INIT = 16'h5410;
  X_LUT4 DLX_EXinst_Ker74459291_G (
    .ADR0(\DLX_IDinst_Imm[3] ),
    .ADR1(\DLX_IDinst_Imm[0] ),
    .ADR2(DLX_IDinst_reg_out_A[25]),
    .ADR3(DLX_IDinst_reg_out_A[24]),
    .O(N165408)
  );
  defparam DLX_EXinst_Ker74459291_F.INIT = 16'h00CA;
  X_LUT4 DLX_EXinst_Ker74459291_F (
    .ADR0(DLX_IDinst_reg_out_A[27]),
    .ADR1(DLX_IDinst_reg_out_A[26]),
    .ADR2(\DLX_IDinst_Imm[0] ),
    .ADR3(\DLX_IDinst_Imm[3] ),
    .O(N165406)
  );
  X_BUF \CHOICE1727/XUSED  (
    .I(\CHOICE1727/F5MUX ),
    .O(CHOICE1727)
  );
  X_MUX2 DLX_EXinst_Ker74629141 (
    .IA(N165671),
    .IB(N165673),
    .SEL(DLX_EXinst__n0036),
    .O(\DLX_IDinst_RegFile_2_28/F5MUX )
  );
  defparam DLX_EXinst_Ker74629141_G.INIT = 16'h0088;
  X_LUT4 DLX_EXinst_Ker74629141_G (
    .ADR0(N148609),
    .ADR1(DLX_IDinst_reg_out_B[4]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[5]),
    .O(N165673)
  );
  defparam DLX_EXinst_Ker74629141_F.INIT = 16'h2020;
  X_LUT4 DLX_EXinst_Ker74629141_F (
    .ADR0(\DLX_IDinst_Imm[4] ),
    .ADR1(\DLX_IDinst_Imm[5] ),
    .ADR2(N147520),
    .ADR3(VCC),
    .O(N165671)
  );
  X_BUF \DLX_IDinst_RegFile_2_28/XUSED  (
    .I(\DLX_IDinst_RegFile_2_28/F5MUX ),
    .O(CHOICE929)
  );
  X_MUX2 DLX_EXinst_Ker75380281 (
    .IA(N165661),
    .IB(N165663),
    .SEL(DLX_IDinst_Imm_3_1),
    .O(\N134128/F5MUX )
  );
  defparam DLX_EXinst_Ker75380281_G.INIT = 16'hAAF0;
  X_LUT4 DLX_EXinst_Ker75380281_G (
    .ADR0(DLX_EXinst_N72958),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N73484),
    .ADR3(\DLX_IDinst_Imm[0] ),
    .O(N165663)
  );
  defparam DLX_EXinst_Ker75380281_F.INIT = 16'hAFA0;
  X_LUT4 DLX_EXinst_Ker75380281_F (
    .ADR0(DLX_EXinst_N72978),
    .ADR1(VCC),
    .ADR2(\DLX_IDinst_Imm[0] ),
    .ADR3(DLX_EXinst_N73374),
    .O(N165661)
  );
  X_BUF \N134128/XUSED  (
    .I(\N134128/F5MUX ),
    .O(N134128)
  );
  X_MUX2 DLX_EXinst_Ker73773171 (
    .IA(N165426),
    .IB(N165428),
    .SEL(DLX_EXinst__n0036),
    .O(\DLX_IFinst_IR_previous<1>/F5MUX )
  );
  defparam DLX_EXinst_Ker73773171_G.INIT = 16'h0C00;
  X_LUT4 DLX_EXinst_Ker73773171_G (
    .ADR0(VCC),
    .ADR1(N148609),
    .ADR2(DLX_IDinst_reg_out_B[4]),
    .ADR3(DLX_IDinst_reg_out_B[5]),
    .O(N165428)
  );
  defparam DLX_EXinst_Ker73773171_F.INIT = 16'h0088;
  X_LUT4 DLX_EXinst_Ker73773171_F (
    .ADR0(N147520),
    .ADR1(\DLX_IDinst_Imm[5] ),
    .ADR2(VCC),
    .ADR3(\DLX_IDinst_Imm[4] ),
    .O(N165426)
  );
  X_BUF \DLX_IFinst_IR_previous<1>/XUSED  (
    .I(\DLX_IFinst_IR_previous<1>/F5MUX ),
    .O(CHOICE1661)
  );
  X_MUX2 DLX_EXinst_Ker75365281 (
    .IA(N165381),
    .IB(N165383),
    .SEL(DLX_IDinst_reg_out_B[0]),
    .O(\N133552/F5MUX )
  );
  defparam DLX_EXinst_Ker75365281_G.INIT = 16'hCCAA;
  X_LUT4 DLX_EXinst_Ker75365281_G (
    .ADR0(DLX_EXinst_N73429),
    .ADR1(DLX_EXinst_N73399),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B_3_1),
    .O(N165383)
  );
  defparam DLX_EXinst_Ker75365281_F.INIT = 16'hF0CC;
  X_LUT4 DLX_EXinst_Ker75365281_F (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N73028),
    .ADR2(DLX_EXinst_N73048),
    .ADR3(DLX_IDinst_reg_out_B_3_1),
    .O(N165381)
  );
  X_BUF \N133552/XUSED  (
    .I(\N133552/F5MUX ),
    .O(N133552)
  );
  X_MUX2 DLX_EXinst_Ker74652581 (
    .IA(N165896),
    .IB(N165898),
    .SEL(\DLX_IDinst_Imm[5] ),
    .O(\DLX_IDinst_RegFile_14_21/F5MUX )
  );
  defparam DLX_EXinst_Ker74652581_G.INIT = 16'h1F00;
  X_LUT4 DLX_EXinst_Ker74652581_G (
    .ADR0(DLX_IDinst_Imm_1_1),
    .ADR1(DLX_IDinst_Imm_2_1),
    .ADR2(DLX_IDinst_Imm_3_1),
    .ADR3(DLX_IDinst_reg_out_A[31]),
    .O(N165898)
  );
  defparam DLX_EXinst_Ker74652581_F.INIT = 16'hFF22;
  X_LUT4 DLX_EXinst_Ker74652581_F (
    .ADR0(DLX_EXinst_N73018),
    .ADR1(DLX_IDinst_Imm_2_1),
    .ADR2(VCC),
    .ADR3(CHOICE2926),
    .O(N165896)
  );
  X_BUF \DLX_IDinst_RegFile_14_21/XUSED  (
    .I(\DLX_IDinst_RegFile_14_21/F5MUX ),
    .O(CHOICE2938)
  );
  X_MUX2 DLX_EXinst_Ker74647601 (
    .IA(N165866),
    .IB(N165868),
    .SEL(\DLX_IDinst_Imm[5] ),
    .O(\CHOICE2965/F5MUX )
  );
  defparam DLX_EXinst_Ker74647601_G.INIT = 16'h2F20;
  X_LUT4 DLX_EXinst_Ker74647601_G (
    .ADR0(\DLX_EXinst_Mshift__n0020_Sh[61] ),
    .ADR1(DLX_IDinst_Imm_2_1),
    .ADR2(DLX_IDinst_Imm_3_1),
    .ADR3(DLX_IDinst_reg_out_A[31]),
    .O(N165868)
  );
  defparam DLX_EXinst_Ker74647601_F.INIT = 16'hFF22;
  X_LUT4 DLX_EXinst_Ker74647601_F (
    .ADR0(DLX_EXinst_N73013),
    .ADR1(DLX_IDinst_Imm_2_1),
    .ADR2(VCC),
    .ADR3(CHOICE2953),
    .O(N165866)
  );
  X_BUF \CHOICE2965/XUSED  (
    .I(\CHOICE2965/F5MUX ),
    .O(CHOICE2965)
  );
  X_MUX2 DLX_EXinst_Ker74674291 (
    .IA(N165386),
    .IB(N165388),
    .SEL(DLX_IDinst_Imm_1_1),
    .O(\DLX_IFinst_IR_previous<4>/F5MUX )
  );
  defparam DLX_EXinst_Ker74674291_G.INIT = 16'h5410;
  X_LUT4 DLX_EXinst_Ker74674291_G (
    .ADR0(DLX_IDinst_Imm_3_1),
    .ADR1(\DLX_IDinst_Imm[0] ),
    .ADR2(DLX_IDinst_reg_out_A[6]),
    .ADR3(DLX_IDinst_reg_out_A[7]),
    .O(N165388)
  );
  defparam DLX_EXinst_Ker74674291_F.INIT = 16'h0C0A;
  X_LUT4 DLX_EXinst_Ker74674291_F (
    .ADR0(DLX_IDinst_reg_out_A[4]),
    .ADR1(DLX_IDinst_reg_out_A[5]),
    .ADR2(DLX_IDinst_Imm_3_1),
    .ADR3(\DLX_IDinst_Imm[0] ),
    .O(N165386)
  );
  X_BUF \DLX_IFinst_IR_previous<4>/XUSED  (
    .I(\DLX_IFinst_IR_previous<4>/F5MUX ),
    .O(CHOICE1791)
  );
  X_MUX2 DLX_EXinst_Ker75493281 (
    .IA(N165356),
    .IB(N165358),
    .SEL(DLX_IDinst_Imm_3_1),
    .O(\N133984/F5MUX )
  );
  defparam DLX_EXinst_Ker75493281_G.INIT = 16'hACAC;
  X_LUT4 DLX_EXinst_Ker75493281_G (
    .ADR0(DLX_EXinst_N73529),
    .ADR1(DLX_EXinst_N73133),
    .ADR2(\DLX_IDinst_Imm[0] ),
    .ADR3(VCC),
    .O(N165358)
  );
  defparam DLX_EXinst_Ker75493281_F.INIT = 16'hCFC0;
  X_LUT4 DLX_EXinst_Ker75493281_F (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N73554),
    .ADR2(\DLX_IDinst_Imm[0] ),
    .ADR3(DLX_EXinst_N73113),
    .O(N165356)
  );
  X_BUF \N133984/XUSED  (
    .I(\N133984/F5MUX ),
    .O(N133984)
  );
  X_MUX2 DLX_EXinst_Ker75498281 (
    .IA(N165456),
    .IB(N165458),
    .SEL(DLX_IDinst_Imm_3_1),
    .O(\DLX_IDinst_RegFile_14_10/F5MUX )
  );
  defparam DLX_EXinst_Ker75498281_G.INIT = 16'hF5A0;
  X_LUT4 DLX_EXinst_Ker75498281_G (
    .ADR0(\DLX_IDinst_Imm[0] ),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N73133),
    .ADR3(DLX_EXinst_N73524),
    .O(N165458)
  );
  defparam DLX_EXinst_Ker75498281_F.INIT = 16'hEE22;
  X_LUT4 DLX_EXinst_Ker75498281_F (
    .ADR0(DLX_EXinst_N73549),
    .ADR1(\DLX_IDinst_Imm[0] ),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N73113),
    .O(N165456)
  );
  X_BUF \DLX_IDinst_RegFile_14_10/XUSED  (
    .I(\DLX_IDinst_RegFile_14_10/F5MUX ),
    .O(N134056)
  );
  X_MUX2 DLX_EXinst_Ker74994281 (
    .IA(N165641),
    .IB(N165643),
    .SEL(DLX_IDinst_reg_out_B[0]),
    .O(\N133048/F5MUX )
  );
  defparam DLX_EXinst_Ker74994281_G.INIT = 16'hD8D8;
  X_LUT4 DLX_EXinst_Ker74994281_G (
    .ADR0(DLX_IDinst_reg_out_B_3_1),
    .ADR1(DLX_EXinst_N73574),
    .ADR2(DLX_EXinst_N73594),
    .ADR3(VCC),
    .O(N165643)
  );
  defparam DLX_EXinst_Ker74994281_F.INIT = 16'hD8D8;
  X_LUT4 DLX_EXinst_Ker74994281_F (
    .ADR0(DLX_IDinst_reg_out_B_3_1),
    .ADR1(DLX_EXinst_N72873),
    .ADR2(DLX_EXinst_N72893),
    .ADR3(VCC),
    .O(N165641)
  );
  X_BUF \N133048/XUSED  (
    .I(\N133048/F5MUX ),
    .O(N133048)
  );
  X_MUX2 DLX_IDinst__n06151 (
    .IA(N165651),
    .IB(N165653),
    .SEL(DLX_IDinst__n0387),
    .O(\DLX_IDinst_RegFile_11_0/F5MUX )
  );
  defparam DLX_IDinst__n06151_G.INIT = 16'h00A0;
  X_LUT4 DLX_IDinst__n06151_G (
    .ADR0(DLX_IDinst_slot_num_FFd3),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_delay_slot),
    .ADR3(DLX_IDinst_slot_num_FFd1),
    .O(N165653)
  );
  defparam DLX_IDinst__n06151_F.INIT = 16'hFFFD;
  X_LUT4 DLX_IDinst__n06151_F (
    .ADR0(DLX_IDinst_stall),
    .ADR1(FREEZE_IBUF),
    .ADR2(DLX_IDinst_N108100),
    .ADR3(DLX_IDinst_delay_slot),
    .O(N165651)
  );
  X_BUF \DLX_IDinst_RegFile_11_0/XUSED  (
    .I(\DLX_IDinst_RegFile_11_0/F5MUX ),
    .O(DLX_IDinst__n0615)
  );
  X_MUX2 DLX_EXinst_Ker74999281 (
    .IA(N165611),
    .IB(N165613),
    .SEL(DLX_IDinst_reg_out_B[0]),
    .O(\N133120/F5MUX )
  );
  defparam DLX_EXinst_Ker74999281_G.INIT = 16'hBB88;
  X_LUT4 DLX_EXinst_Ker74999281_G (
    .ADR0(DLX_EXinst_N72873),
    .ADR1(DLX_IDinst_reg_out_B_3_1),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N72893),
    .O(N165613)
  );
  defparam DLX_EXinst_Ker74999281_F.INIT = 16'hDD88;
  X_LUT4 DLX_EXinst_Ker74999281_F (
    .ADR0(DLX_IDinst_reg_out_B_3_1),
    .ADR1(DLX_EXinst_N73579),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N73354),
    .O(N165611)
  );
  X_BUF \N133120/XUSED  (
    .I(\N133120/F5MUX ),
    .O(N133120)
  );
  X_MUX2 \DLX_EXinst__n0007<8>951  (
    .IA(N165946),
    .IB(N165948),
    .SEL(DLX_IDinst_reg_out_B[4]),
    .O(\DLX_IDinst_RegFile_14_22/F5MUX )
  );
  defparam \DLX_EXinst__n0007<8>951_G .INIT = 16'h0200;
  X_LUT4 \DLX_EXinst__n0007<8>951_G  (
    .ADR0(DLX_EXinst_N73369),
    .ADR1(N148323),
    .ADR2(DLX_IDinst_reg_out_B[3]),
    .ADR3(DLX_EXinst__n0081),
    .O(N165948)
  );
  defparam \DLX_EXinst__n0007<8>951_F .INIT = 16'h3000;
  X_LUT4 \DLX_EXinst__n0007<8>951_F  (
    .ADR0(VCC),
    .ADR1(N148323),
    .ADR2(\DLX_EXinst_Mshift__n0023_Sh[40] ),
    .ADR3(DLX_EXinst__n0080),
    .O(N165946)
  );
  X_BUF \DLX_IDinst_RegFile_14_22/XUSED  (
    .I(\DLX_IDinst_RegFile_14_22/F5MUX ),
    .O(CHOICE5154)
  );
  X_MUX2 \DM_read_data<0>11  (
    .IA(N165686),
    .IB(N165688),
    .SEL(DLX_EXinst_ALU_result[12]),
    .O(\DM_read_data<0>/F5MUX )
  );
  defparam \DM_read_data<0>11_G .INIT = 16'hFAF8;
  X_LUT4 \DM_read_data<0>11_G  (
    .ADR0(DLX_EXinst_ALU_result[13]),
    .ADR1(vram_out_cpu[2]),
    .ADR2(CHOICE246),
    .ADR3(DLX_EXinst_ALU_result[14]),
    .O(N165688)
  );
  defparam \DM_read_data<0>11_F .INIT = 16'hFAF8;
  X_LUT4 \DM_read_data<0>11_F  (
    .ADR0(DLX_EXinst_ALU_result[13]),
    .ADR1(DLX_EXinst_ALU_result[14]),
    .ADR2(CHOICE254),
    .ADR3(vram_out_cpu[1]),
    .O(N165686)
  );
  X_BUF \DM_read_data<0>/XUSED  (
    .I(\DM_read_data<0>/F5MUX ),
    .O(DM_read_data[0])
  );
  X_ONE \vram_out_vga_eff/LOGIC_ONE_1612  (
    .O(\vram_out_vga_eff/LOGIC_ONE )
  );
  X_MUX2 \Mmux__COND_2_inst_mux_f6_0.F51_1613  (
    .IA(\NLW_Mmux__COND_2_inst_mux_f6_0.F51_IA_UNCONNECTED ),
    .IB(\vram_out_vga<4>_rt ),
    .SEL(\vram_out_vga_eff/LOGIC_ONE ),
    .O(\Mmux__COND_2_inst_mux_f6_0.F51 )
  );
  defparam \vram_out_vga<4>_rt_1614 .INIT = 16'hFF00;
  X_LUT4 \vram_out_vga<4>_rt_1614  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vram_out_vga[4]),
    .O(\vram_out_vga<4>_rt )
  );
  X_BUF \vram_out_vga_eff/YUSED  (
    .I(\vram_out_vga_eff/F6MUX ),
    .O(vram_out_vga_eff)
  );
  X_MUX2 Mmux__COND_2_inst_mux_f6_0 (
    .IA(Mmux__COND_2__net2),
    .IB(\Mmux__COND_2_inst_mux_f6_0.F51 ),
    .SEL(vga_address[14]),
    .O(\vram_out_vga_eff/F6MUX )
  );
  X_MUX2 \DLX_EXinst__n0007<15>26211  (
    .IA(N165646),
    .IB(N165648),
    .SEL(DLX_EXinst__n0036),
    .O(N162847)
  );
  defparam \DLX_EXinst__n0007<15>26211_G .INIT = 16'hFCCC;
  X_LUT4 \DLX_EXinst__n0007<15>26211_G  (
    .ADR0(VCC),
    .ADR1(CHOICE4316),
    .ADR2(DLX_EXinst__n0012[15]),
    .ADR3(DLX_EXinst__n0127),
    .O(N165648)
  );
  defparam \DLX_EXinst__n0007<15>26211_F .INIT = 16'hFFEC;
  X_LUT4 \DLX_EXinst__n0007<15>26211_F  (
    .ADR0(DLX_EXinst__n0109),
    .ADR1(CHOICE4316),
    .ADR2(DLX_EXinst__n0012[15]),
    .ADR3(CHOICE4314),
    .O(N165646)
  );
  defparam DLX_IDinst_RegFile_28_19_1615.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_28_19_1615 (
    .I(DLX_IDinst_WB_data_eff[19]),
    .CE(DLX_IDinst__n0606),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_28_19)
  );
  X_MUX2 Mmux__COND_2_inst_mux_f5_0 (
    .IA(Mmux__COND_2__net0),
    .IB(Mmux__COND_2__net1),
    .SEL(vga_address[13]),
    .O(\Mmux__COND_2__net2/F5MUX )
  );
  defparam Mmux__COND_2_inst_lut3_11.INIT = 16'hCCAA;
  X_LUT4 Mmux__COND_2_inst_lut3_11 (
    .ADR0(vram_out_vga[2]),
    .ADR1(vram_out_vga[3]),
    .ADR2(VCC),
    .ADR3(vga_address[12]),
    .O(Mmux__COND_2__net1)
  );
  defparam Mmux__COND_2_inst_lut3_01.INIT = 16'hEE22;
  X_LUT4 Mmux__COND_2_inst_lut3_01 (
    .ADR0(vram_out_vga[0]),
    .ADR1(vga_address[12]),
    .ADR2(VCC),
    .ADR3(vram_out_vga[1]),
    .O(Mmux__COND_2__net0)
  );
  X_BUF \Mmux__COND_2__net2/F5USED  (
    .I(\Mmux__COND_2__net2/F5MUX ),
    .O(Mmux__COND_2__net2)
  );
  X_MUX2 DLX_IDinst_Ker108226201 (
    .IA(N165951),
    .IB(N165953),
    .SEL(DLX_IDinst_IR_latched[26]),
    .O(\DLX_MEMinst_opcode_of_WB<3>/F5MUX )
  );
  defparam DLX_IDinst_Ker108226201_G.INIT = 16'hFFFB;
  X_LUT4 DLX_IDinst_Ker108226201_G (
    .ADR0(DLX_IDinst_IR_latched[31]),
    .ADR1(DLX_IDinst_N108221),
    .ADR2(DLX_IDinst_zflag),
    .ADR3(DLX_IDinst_IR_latched[29]),
    .O(N165953)
  );
  defparam DLX_IDinst_Ker108226201_F.INIT = 16'h77FF;
  X_LUT4 DLX_IDinst_Ker108226201_F (
    .ADR0(DLX_IDinst_IR_latched[30]),
    .ADR1(DLX_IDinst_N108165),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_IR_latched[27]),
    .O(N165951)
  );
  X_BUF \DLX_MEMinst_opcode_of_WB<3>/XUSED  (
    .I(\DLX_MEMinst_opcode_of_WB<3>/F5MUX ),
    .O(CHOICE3373)
  );
  X_MUX2 \DLX_IFinst__n0003<10>1  (
    .IA(N165926),
    .IB(N165928),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[10])
  );
  defparam \DLX_IFinst__n0003<10>1_G .INIT = 16'hFC30;
  X_LUT4 \DLX_IFinst__n0003<10>1_G  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(DLX_IFinst_IR_previous[10]),
    .ADR3(IR[10]),
    .O(N165928)
  );
  defparam \DLX_IFinst__n0003<10>1_F .INIT = 16'hD8CC;
  X_LUT4 \DLX_IFinst__n0003<10>1_F  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(IR[10]),
    .ADR2(DLX_IFinst_IR_curr[10]),
    .ADR3(DLX_IFinst_stalled),
    .O(N165926)
  );
  X_MUX2 \DLX_IFinst__n0003<11>1  (
    .IA(N165791),
    .IB(N165793),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[11])
  );
  defparam \DLX_IFinst__n0003<11>1_G .INIT = 16'hAAF0;
  X_LUT4 \DLX_IFinst__n0003<11>1_G  (
    .ADR0(IR[11]),
    .ADR1(VCC),
    .ADR2(DLX_IFinst_IR_previous[11]),
    .ADR3(DLX_IDinst_branch_sig),
    .O(N165793)
  );
  defparam \DLX_IFinst__n0003<11>1_F .INIT = 16'hF0B8;
  X_LUT4 \DLX_IFinst__n0003<11>1_F  (
    .ADR0(DLX_IFinst_IR_curr[11]),
    .ADR1(DLX_IFinst_stalled),
    .ADR2(IR[11]),
    .ADR3(DLX_IDinst_branch_sig),
    .O(N165791)
  );
  X_MUX2 \DLX_IFinst__n0003<20>1  (
    .IA(N165921),
    .IB(N165923),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[20])
  );
  defparam \DLX_IFinst__n0003<20>1_G .INIT = 16'hE4E4;
  X_LUT4 \DLX_IFinst__n0003<20>1_G  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(DLX_IFinst_IR_previous[20]),
    .ADR2(IR[20]),
    .ADR3(VCC),
    .O(N165923)
  );
  defparam \DLX_IFinst__n0003<20>1_F .INIT = 16'hCCE4;
  X_LUT4 \DLX_IFinst__n0003<20>1_F  (
    .ADR0(DLX_IFinst_stalled),
    .ADR1(IR[20]),
    .ADR2(DLX_IFinst_IR_curr[20]),
    .ADR3(DLX_IDinst_branch_sig),
    .O(N165921)
  );
  X_MUX2 \DLX_IFinst__n0003<12>1  (
    .IA(N165806),
    .IB(N165808),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[12])
  );
  defparam \DLX_IFinst__n0003<12>1_G .INIT = 16'hF3C0;
  X_LUT4 \DLX_IFinst__n0003<12>1_G  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(IR[12]),
    .ADR3(DLX_IFinst_IR_previous[12]),
    .O(N165808)
  );
  defparam \DLX_IFinst__n0003<12>1_F .INIT = 16'hFD20;
  X_LUT4 \DLX_IFinst__n0003<12>1_F  (
    .ADR0(DLX_IFinst_stalled),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(DLX_IFinst_IR_curr[12]),
    .ADR3(IR[12]),
    .O(N165806)
  );
  defparam DLX_IDinst_RegFile_29_11_1616.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_29_11_1616 (
    .I(DLX_IDinst_WB_data_eff[11]),
    .CE(DLX_IDinst__n0608),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_29_11)
  );
  X_MUX2 \DLX_IFinst__n0003<13>1  (
    .IA(N165886),
    .IB(N165888),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[13])
  );
  defparam \DLX_IFinst__n0003<13>1_G .INIT = 16'hEE44;
  X_LUT4 \DLX_IFinst__n0003<13>1_G  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(DLX_IFinst_IR_previous[13]),
    .ADR2(VCC),
    .ADR3(IR[13]),
    .O(N165888)
  );
  defparam \DLX_IFinst__n0003<13>1_F .INIT = 16'hFB40;
  X_LUT4 \DLX_IFinst__n0003<13>1_F  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(DLX_IFinst_stalled),
    .ADR2(DLX_IFinst_IR_curr[13]),
    .ADR3(IR[13]),
    .O(N165886)
  );
  X_MUX2 \DLX_IFinst__n0003<21>1  (
    .IA(N165751),
    .IB(N165753),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[21])
  );
  defparam \DLX_IFinst__n0003<21>1_G .INIT = 16'hFC0C;
  X_LUT4 \DLX_IFinst__n0003<21>1_G  (
    .ADR0(VCC),
    .ADR1(DLX_IFinst_IR_previous[21]),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(IR[21]),
    .O(N165753)
  );
  defparam \DLX_IFinst__n0003<21>1_F .INIT = 16'hF2D0;
  X_LUT4 \DLX_IFinst__n0003<21>1_F  (
    .ADR0(DLX_IFinst_stalled),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(IR[21]),
    .ADR3(DLX_IFinst_IR_curr[21]),
    .O(N165751)
  );
  X_MUX2 \DLX_IFinst__n0003<30>1  (
    .IA(N165911),
    .IB(N165913),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[30])
  );
  defparam \DLX_IFinst__n0003<30>1_G .INIT = 16'hCCF0;
  X_LUT4 \DLX_IFinst__n0003<30>1_G  (
    .ADR0(VCC),
    .ADR1(IR_MSB_6_OBUF),
    .ADR2(DLX_IFinst_IR_previous[30]),
    .ADR3(DLX_IDinst_branch_sig),
    .O(N165913)
  );
  defparam \DLX_IFinst__n0003<30>1_F .INIT = 16'hF2D0;
  X_LUT4 \DLX_IFinst__n0003<30>1_F  (
    .ADR0(DLX_IFinst_stalled),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(IR_MSB_6_OBUF),
    .ADR3(DLX_IFinst_IR_curr[30]),
    .O(N165911)
  );
  X_MUX2 \DLX_IFinst__n0003<14>1  (
    .IA(N165776),
    .IB(N165778),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[14])
  );
  defparam \DLX_IFinst__n0003<14>1_G .INIT = 16'hE4E4;
  X_LUT4 \DLX_IFinst__n0003<14>1_G  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(DLX_IFinst_IR_previous[14]),
    .ADR2(IR[14]),
    .ADR3(VCC),
    .O(N165778)
  );
  defparam \DLX_IFinst__n0003<14>1_F .INIT = 16'hF0D8;
  X_LUT4 \DLX_IFinst__n0003<14>1_F  (
    .ADR0(DLX_IFinst_stalled),
    .ADR1(DLX_IFinst_IR_curr[14]),
    .ADR2(IR[14]),
    .ADR3(DLX_IDinst_branch_sig),
    .O(N165776)
  );
  X_MUX2 \DLX_IFinst__n0003<22>1  (
    .IA(N165396),
    .IB(N165398),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[22])
  );
  defparam \DLX_IFinst__n0003<22>1_G .INIT = 16'hFC30;
  X_LUT4 \DLX_IFinst__n0003<22>1_G  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(DLX_IFinst_IR_previous[22]),
    .ADR3(IR[22]),
    .O(N165398)
  );
  defparam \DLX_IFinst__n0003<22>1_F .INIT = 16'hE4F0;
  X_LUT4 \DLX_IFinst__n0003<22>1_F  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(DLX_IFinst_IR_curr[22]),
    .ADR2(IR[22]),
    .ADR3(DLX_IFinst_stalled),
    .O(N165396)
  );
  X_MUX2 \DLX_IFinst__n0003<23>1  (
    .IA(N165871),
    .IB(N165873),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[23])
  );
  defparam \DLX_IFinst__n0003<23>1_G .INIT = 16'hFC30;
  X_LUT4 \DLX_IFinst__n0003<23>1_G  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(DLX_IFinst_IR_previous[23]),
    .ADR3(IR[23]),
    .O(N165873)
  );
  defparam \DLX_IFinst__n0003<23>1_F .INIT = 16'hE2F0;
  X_LUT4 \DLX_IFinst__n0003<23>1_F  (
    .ADR0(DLX_IFinst_IR_curr[23]),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(IR[23]),
    .ADR3(DLX_IFinst_stalled),
    .O(N165871)
  );
  X_MUX2 \DLX_IFinst__n0003<15>1  (
    .IA(N165836),
    .IB(N165838),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[15])
  );
  defparam \DLX_IFinst__n0003<15>1_G .INIT = 16'hCCF0;
  X_LUT4 \DLX_IFinst__n0003<15>1_G  (
    .ADR0(VCC),
    .ADR1(IR[15]),
    .ADR2(DLX_IFinst_IR_previous[15]),
    .ADR3(DLX_IDinst_branch_sig),
    .O(N165838)
  );
  defparam \DLX_IFinst__n0003<15>1_F .INIT = 16'hFB08;
  X_LUT4 \DLX_IFinst__n0003<15>1_F  (
    .ADR0(DLX_IFinst_IR_curr[15]),
    .ADR1(DLX_IFinst_stalled),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(IR[15]),
    .O(N165836)
  );
  X_MUX2 \DLX_IFinst__n0003<31>1  (
    .IA(N165676),
    .IB(N165678),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[31])
  );
  defparam \DLX_IFinst__n0003<31>1_G .INIT = 16'hF0AA;
  X_LUT4 \DLX_IFinst__n0003<31>1_G  (
    .ADR0(DLX_IFinst_IR_previous[31]),
    .ADR1(VCC),
    .ADR2(IR_MSB_7_OBUF),
    .ADR3(DLX_IDinst_branch_sig),
    .O(N165678)
  );
  defparam \DLX_IFinst__n0003<31>1_F .INIT = 16'hFB40;
  X_LUT4 \DLX_IFinst__n0003<31>1_F  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(DLX_IFinst_stalled),
    .ADR2(DLX_IFinst_IR_curr[31]),
    .ADR3(IR_MSB_7_OBUF),
    .O(N165676)
  );
  X_MUX2 \DLX_IFinst__n0003<24>1  (
    .IA(N165881),
    .IB(N165883),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[24])
  );
  defparam \DLX_IFinst__n0003<24>1_G .INIT = 16'hFC0C;
  X_LUT4 \DLX_IFinst__n0003<24>1_G  (
    .ADR0(VCC),
    .ADR1(DLX_IFinst_IR_previous[24]),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(IR_MSB_0_OBUF),
    .O(N165883)
  );
  defparam \DLX_IFinst__n0003<24>1_F .INIT = 16'hFD08;
  X_LUT4 \DLX_IFinst__n0003<24>1_F  (
    .ADR0(DLX_IFinst_stalled),
    .ADR1(DLX_IFinst_IR_curr[24]),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(IR_MSB_0_OBUF),
    .O(N165881)
  );
  X_MUX2 \DLX_IFinst__n0003<16>1  (
    .IA(N165856),
    .IB(N165858),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[16])
  );
  defparam \DLX_IFinst__n0003<16>1_G .INIT = 16'hBB88;
  X_LUT4 \DLX_IFinst__n0003<16>1_G  (
    .ADR0(IR[16]),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(VCC),
    .ADR3(DLX_IFinst_IR_previous[16]),
    .O(N165858)
  );
  defparam \DLX_IFinst__n0003<16>1_F .INIT = 16'hFD20;
  X_LUT4 \DLX_IFinst__n0003<16>1_F  (
    .ADR0(DLX_IFinst_stalled),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(DLX_IFinst_IR_curr[16]),
    .ADR3(IR[16]),
    .O(N165856)
  );
  X_MUX2 \DLX_IFinst__n0003<17>1  (
    .IA(N165851),
    .IB(N165853),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[17])
  );
  defparam \DLX_IFinst__n0003<17>1_G .INIT = 16'hAACC;
  X_LUT4 \DLX_IFinst__n0003<17>1_G  (
    .ADR0(IR[17]),
    .ADR1(DLX_IFinst_IR_previous[17]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_branch_sig),
    .O(N165853)
  );
  defparam \DLX_IFinst__n0003<17>1_F .INIT = 16'hCCE4;
  X_LUT4 \DLX_IFinst__n0003<17>1_F  (
    .ADR0(DLX_IFinst_stalled),
    .ADR1(IR[17]),
    .ADR2(DLX_IFinst_IR_curr[17]),
    .ADR3(DLX_IDinst_branch_sig),
    .O(N165851)
  );
  X_MUX2 \DLX_IFinst__n0003<25>1  (
    .IA(N165811),
    .IB(N165813),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[25])
  );
  defparam \DLX_IFinst__n0003<25>1_G .INIT = 16'hE2E2;
  X_LUT4 \DLX_IFinst__n0003<25>1_G  (
    .ADR0(DLX_IFinst_IR_previous[25]),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(IR_MSB_1_OBUF),
    .ADR3(VCC),
    .O(N165813)
  );
  defparam \DLX_IFinst__n0003<25>1_F .INIT = 16'hEF20;
  X_LUT4 \DLX_IFinst__n0003<25>1_F  (
    .ADR0(DLX_IFinst_IR_curr[25]),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(DLX_IFinst_stalled),
    .ADR3(IR_MSB_1_OBUF),
    .O(N165811)
  );
  X_MUX2 \DLX_IFinst__n0003<18>1  (
    .IA(N165901),
    .IB(N165903),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[18])
  );
  defparam \DLX_IFinst__n0003<18>1_G .INIT = 16'hFC30;
  X_LUT4 \DLX_IFinst__n0003<18>1_G  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(DLX_IFinst_IR_previous[18]),
    .ADR3(IR[18]),
    .O(N165903)
  );
  defparam \DLX_IFinst__n0003<18>1_F .INIT = 16'hFD08;
  X_LUT4 \DLX_IFinst__n0003<18>1_F  (
    .ADR0(DLX_IFinst_stalled),
    .ADR1(DLX_IFinst_IR_curr[18]),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(IR[18]),
    .O(N165901)
  );
  X_MUX2 \DLX_IFinst__n0003<26>1  (
    .IA(N165716),
    .IB(N165718),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[26])
  );
  defparam \DLX_IFinst__n0003<26>1_G .INIT = 16'hF3C0;
  X_LUT4 \DLX_IFinst__n0003<26>1_G  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(IR_MSB_2_OBUF),
    .ADR3(DLX_IFinst_IR_previous[26]),
    .O(N165718)
  );
  defparam \DLX_IFinst__n0003<26>1_F .INIT = 16'hF2D0;
  X_LUT4 \DLX_IFinst__n0003<26>1_F  (
    .ADR0(DLX_IFinst_stalled),
    .ADR1(DLX_IDinst_branch_sig),
    .ADR2(IR_MSB_2_OBUF),
    .ADR3(DLX_IFinst_IR_curr[26]),
    .O(N165716)
  );
  X_MUX2 \DLX_IFinst__n0003<19>1  (
    .IA(N165906),
    .IB(N165908),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[19])
  );
  defparam \DLX_IFinst__n0003<19>1_G .INIT = 16'hE4E4;
  X_LUT4 \DLX_IFinst__n0003<19>1_G  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(DLX_IFinst_IR_previous[19]),
    .ADR2(IR[19]),
    .ADR3(VCC),
    .O(N165908)
  );
  defparam \DLX_IFinst__n0003<19>1_F .INIT = 16'hF4B0;
  X_LUT4 \DLX_IFinst__n0003<19>1_F  (
    .ADR0(DLX_IDinst_branch_sig),
    .ADR1(DLX_IFinst_stalled),
    .ADR2(IR[19]),
    .ADR3(DLX_IFinst_IR_curr[19]),
    .O(N165906)
  );
  X_MUX2 \DLX_IFinst__n0003<27>1  (
    .IA(N165761),
    .IB(N165763),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[27])
  );
  defparam \DLX_IFinst__n0003<27>1_G .INIT = 16'hCFC0;
  X_LUT4 \DLX_IFinst__n0003<27>1_G  (
    .ADR0(VCC),
    .ADR1(IR_MSB_3_OBUF),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(DLX_IFinst_IR_previous[27]),
    .O(N165763)
  );
  defparam \DLX_IFinst__n0003<27>1_F .INIT = 16'hCACC;
  X_LUT4 \DLX_IFinst__n0003<27>1_F  (
    .ADR0(DLX_IFinst_IR_curr[27]),
    .ADR1(IR_MSB_3_OBUF),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(DLX_IFinst_stalled),
    .O(N165761)
  );
  X_MUX2 \DLX_IFinst__n0003<28>1  (
    .IA(N165936),
    .IB(N165938),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[28])
  );
  defparam \DLX_IFinst__n0003<28>1_G .INIT = 16'hAAF0;
  X_LUT4 \DLX_IFinst__n0003<28>1_G  (
    .ADR0(IR_MSB_4_OBUF),
    .ADR1(VCC),
    .ADR2(DLX_IFinst_IR_previous[28]),
    .ADR3(DLX_IDinst_branch_sig),
    .O(N165938)
  );
  defparam \DLX_IFinst__n0003<28>1_F .INIT = 16'hCACC;
  X_LUT4 \DLX_IFinst__n0003<28>1_F  (
    .ADR0(DLX_IFinst_IR_curr[28]),
    .ADR1(IR_MSB_4_OBUF),
    .ADR2(DLX_IDinst_branch_sig),
    .ADR3(DLX_IFinst_stalled),
    .O(N165936)
  );
  X_MUX2 \DLX_IFinst__n0003<29>1  (
    .IA(N165831),
    .IB(N165833),
    .SEL(DLX_IFinst__n0000),
    .O(DLX_IFinst__n0003[29])
  );
  defparam \DLX_IFinst__n0003<29>1_G .INIT = 16'hF0CC;
  X_LUT4 \DLX_IFinst__n0003<29>1_G  (
    .ADR0(VCC),
    .ADR1(DLX_IFinst_IR_previous[29]),
    .ADR2(IR_MSB_5_OBUF),
    .ADR3(DLX_IDinst_branch_sig),
    .O(N165833)
  );
  defparam \DLX_IFinst__n0003<29>1_F .INIT = 16'hAAE2;
  X_LUT4 \DLX_IFinst__n0003<29>1_F  (
    .ADR0(IR_MSB_5_OBUF),
    .ADR1(DLX_IFinst_stalled),
    .ADR2(DLX_IFinst_IR_curr[29]),
    .ADR3(DLX_IDinst_branch_sig),
    .O(N165831)
  );
  X_MUX2 DLX_EXinst_Ker751521 (
    .IA(N165551),
    .IB(N165553),
    .SEL(DLX_IDinst_Imm_2_1),
    .O(\DLX_EXinst_N75154/F5MUX )
  );
  defparam DLX_EXinst_Ker751521_G.INIT = 16'h2B28;
  X_LUT4 DLX_EXinst_Ker751521_G (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(DLX_IDinst_Imm_3_1),
    .ADR2(\DLX_IDinst_Imm[5] ),
    .ADR3(\DLX_EXinst_Mshift__n0022_Sh[24] ),
    .O(N165553)
  );
  defparam DLX_EXinst_Ker751521_F.INIT = 16'hF0CC;
  X_LUT4 DLX_EXinst_Ker751521_F (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N72797),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(\DLX_IDinst_Imm[5] ),
    .O(N165551)
  );
  X_BUF \DLX_EXinst_N75154/XUSED  (
    .I(\DLX_EXinst_N75154/F5MUX ),
    .O(DLX_EXinst_N75154)
  );
  X_MUX2 DLX_EXinst_Ker749641 (
    .IA(N165431),
    .IB(N165433),
    .SEL(DLX_IDinst_reg_out_B_2_1),
    .O(\DLX_IDinst_RegFile_22_14/F5MUX )
  );
  defparam DLX_EXinst_Ker749641_G.INIT = 16'h7610;
  X_LUT4 DLX_EXinst_Ker749641_G (
    .ADR0(DLX_IDinst_reg_out_B_3_1),
    .ADR1(DLX_IDinst_reg_out_B[5]),
    .ADR2(\DLX_EXinst_Mshift__n0019_Sh[24] ),
    .ADR3(DLX_IDinst_reg_out_A[31]),
    .O(N165433)
  );
  defparam DLX_EXinst_Ker749641_F.INIT = 16'hF3C0;
  X_LUT4 DLX_EXinst_Ker749641_F (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_B[5]),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(DLX_EXinst_N72809),
    .O(N165431)
  );
  X_BUF \DLX_IDinst_RegFile_22_14/XUSED  (
    .I(\DLX_IDinst_RegFile_22_14/F5MUX ),
    .O(DLX_EXinst_N74966)
  );
  X_ZERO \vga_top_vga1_vcounter<0>/LOGIC_ZERO_1617  (
    .O(\vga_top_vga1_vcounter<0>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_vcounter_Madd__n0000_inst_cy_9_1618 (
    .IA(GLOBAL_LOGIC1),
    .IB(\vga_top_vga1_vcounter<0>/LOGIC_ZERO ),
    .SEL(vga_top_vga1_vcounter_Madd__n0000_inst_lut2_9),
    .O(vga_top_vga1_vcounter_Madd__n0000_inst_cy_9)
  );
  defparam vga_top_vga1_vcounter_Madd__n0000_inst_lut2_91.INIT = 16'h3333;
  X_LUT4 vga_top_vga1_vcounter_Madd__n0000_inst_lut2_91 (
    .ADR0(GLOBAL_LOGIC1),
    .ADR1(vga_top_vga1_vcounter[0]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(vga_top_vga1_vcounter_Madd__n0000_inst_lut2_9)
  );
  defparam \vga_top_vga1_vcounter<0>/G .INIT = 16'hFF00;
  X_LUT4 \vga_top_vga1_vcounter<0>/G  (
    .ADR0(GLOBAL_LOGIC0),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_vcounter[1]),
    .O(\vga_top_vga1_vcounter<0>/GROM )
  );
  X_BUF \vga_top_vga1_vcounter<0>/COUTUSED  (
    .I(\vga_top_vga1_vcounter<0>/CYMUXG ),
    .O(vga_top_vga1_vcounter_Madd__n0000_inst_cy_10)
  );
  X_MUX2 vga_top_vga1_vcounter_Madd__n0000_inst_cy_10_1619 (
    .IA(GLOBAL_LOGIC0),
    .IB(vga_top_vga1_vcounter_Madd__n0000_inst_cy_9),
    .SEL(\vga_top_vga1_vcounter<0>/GROM ),
    .O(\vga_top_vga1_vcounter<0>/CYMUXG )
  );
  X_XOR2 vga_top_vga1_vcounter_Madd__n0000_inst_sum_10 (
    .I0(vga_top_vga1_vcounter_Madd__n0000_inst_cy_9),
    .I1(\vga_top_vga1_vcounter<0>/GROM ),
    .O(vga_top_vga1_vcounter__n0000[1])
  );
  X_ZERO \vga_top_vga1_vcounter<2>/LOGIC_ZERO_1620  (
    .O(\vga_top_vga1_vcounter<2>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_vcounter_Madd__n0000_inst_cy_11_1621 (
    .IA(\vga_top_vga1_vcounter<2>/LOGIC_ZERO ),
    .IB(\vga_top_vga1_vcounter<2>/CYINIT ),
    .SEL(\vga_top_vga1_vcounter<2>/FROM ),
    .O(vga_top_vga1_vcounter_Madd__n0000_inst_cy_11)
  );
  X_XOR2 vga_top_vga1_vcounter_Madd__n0000_inst_sum_11 (
    .I0(\vga_top_vga1_vcounter<2>/CYINIT ),
    .I1(\vga_top_vga1_vcounter<2>/FROM ),
    .O(vga_top_vga1_vcounter__n0000[2])
  );
  defparam \vga_top_vga1_vcounter<2>/F .INIT = 16'hFF00;
  X_LUT4 \vga_top_vga1_vcounter<2>/F  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_vcounter[2]),
    .O(\vga_top_vga1_vcounter<2>/FROM )
  );
  defparam \vga_top_vga1_vcounter<2>/G .INIT = 16'hCCCC;
  X_LUT4 \vga_top_vga1_vcounter<2>/G  (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_vcounter[3]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\vga_top_vga1_vcounter<2>/GROM )
  );
  X_BUF \vga_top_vga1_vcounter<2>/COUTUSED  (
    .I(\vga_top_vga1_vcounter<2>/CYMUXG ),
    .O(vga_top_vga1_vcounter_Madd__n0000_inst_cy_12)
  );
  X_MUX2 vga_top_vga1_vcounter_Madd__n0000_inst_cy_12_1622 (
    .IA(\vga_top_vga1_vcounter<2>/LOGIC_ZERO ),
    .IB(vga_top_vga1_vcounter_Madd__n0000_inst_cy_11),
    .SEL(\vga_top_vga1_vcounter<2>/GROM ),
    .O(\vga_top_vga1_vcounter<2>/CYMUXG )
  );
  X_XOR2 vga_top_vga1_vcounter_Madd__n0000_inst_sum_12 (
    .I0(vga_top_vga1_vcounter_Madd__n0000_inst_cy_11),
    .I1(\vga_top_vga1_vcounter<2>/GROM ),
    .O(vga_top_vga1_vcounter__n0000[3])
  );
  X_BUF \vga_top_vga1_vcounter<2>/CYINIT_1623  (
    .I(vga_top_vga1_vcounter_Madd__n0000_inst_cy_10),
    .O(\vga_top_vga1_vcounter<2>/CYINIT )
  );
  X_ZERO \vga_top_vga1_vcounter<4>/LOGIC_ZERO_1624  (
    .O(\vga_top_vga1_vcounter<4>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_vcounter_Madd__n0000_inst_cy_13_1625 (
    .IA(\vga_top_vga1_vcounter<4>/LOGIC_ZERO ),
    .IB(\vga_top_vga1_vcounter<4>/CYINIT ),
    .SEL(\vga_top_vga1_vcounter<4>/FROM ),
    .O(vga_top_vga1_vcounter_Madd__n0000_inst_cy_13)
  );
  X_XOR2 vga_top_vga1_vcounter_Madd__n0000_inst_sum_13 (
    .I0(\vga_top_vga1_vcounter<4>/CYINIT ),
    .I1(\vga_top_vga1_vcounter<4>/FROM ),
    .O(vga_top_vga1_vcounter__n0000[4])
  );
  defparam \vga_top_vga1_vcounter<4>/F .INIT = 16'hAAAA;
  X_LUT4 \vga_top_vga1_vcounter<4>/F  (
    .ADR0(vga_top_vga1_vcounter[4]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\vga_top_vga1_vcounter<4>/FROM )
  );
  defparam \vga_top_vga1_vcounter<4>/G .INIT = 16'hF0F0;
  X_LUT4 \vga_top_vga1_vcounter<4>/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_vcounter[5]),
    .ADR3(VCC),
    .O(\vga_top_vga1_vcounter<4>/GROM )
  );
  X_BUF \vga_top_vga1_vcounter<4>/COUTUSED  (
    .I(\vga_top_vga1_vcounter<4>/CYMUXG ),
    .O(vga_top_vga1_vcounter_Madd__n0000_inst_cy_14)
  );
  X_MUX2 vga_top_vga1_vcounter_Madd__n0000_inst_cy_14_1626 (
    .IA(\vga_top_vga1_vcounter<4>/LOGIC_ZERO ),
    .IB(vga_top_vga1_vcounter_Madd__n0000_inst_cy_13),
    .SEL(\vga_top_vga1_vcounter<4>/GROM ),
    .O(\vga_top_vga1_vcounter<4>/CYMUXG )
  );
  X_XOR2 vga_top_vga1_vcounter_Madd__n0000_inst_sum_14 (
    .I0(vga_top_vga1_vcounter_Madd__n0000_inst_cy_13),
    .I1(\vga_top_vga1_vcounter<4>/GROM ),
    .O(vga_top_vga1_vcounter__n0000[5])
  );
  X_BUF \vga_top_vga1_vcounter<4>/CYINIT_1627  (
    .I(vga_top_vga1_vcounter_Madd__n0000_inst_cy_12),
    .O(\vga_top_vga1_vcounter<4>/CYINIT )
  );
  X_ZERO \vga_top_vga1_vcounter<6>/LOGIC_ZERO_1628  (
    .O(\vga_top_vga1_vcounter<6>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_vcounter_Madd__n0000_inst_cy_15_1629 (
    .IA(\vga_top_vga1_vcounter<6>/LOGIC_ZERO ),
    .IB(\vga_top_vga1_vcounter<6>/CYINIT ),
    .SEL(\vga_top_vga1_vcounter<6>/FROM ),
    .O(vga_top_vga1_vcounter_Madd__n0000_inst_cy_15)
  );
  X_XOR2 vga_top_vga1_vcounter_Madd__n0000_inst_sum_15 (
    .I0(\vga_top_vga1_vcounter<6>/CYINIT ),
    .I1(\vga_top_vga1_vcounter<6>/FROM ),
    .O(vga_top_vga1_vcounter__n0000[6])
  );
  defparam \vga_top_vga1_vcounter<6>/F .INIT = 16'hCCCC;
  X_LUT4 \vga_top_vga1_vcounter<6>/F  (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_vcounter[6]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\vga_top_vga1_vcounter<6>/FROM )
  );
  defparam \vga_top_vga1_vcounter<6>/G .INIT = 16'hF0F0;
  X_LUT4 \vga_top_vga1_vcounter<6>/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_vcounter[7]),
    .ADR3(VCC),
    .O(\vga_top_vga1_vcounter<6>/GROM )
  );
  X_BUF \vga_top_vga1_vcounter<6>/COUTUSED  (
    .I(\vga_top_vga1_vcounter<6>/CYMUXG ),
    .O(vga_top_vga1_vcounter_Madd__n0000_inst_cy_16)
  );
  X_MUX2 vga_top_vga1_vcounter_Madd__n0000_inst_cy_16_1630 (
    .IA(\vga_top_vga1_vcounter<6>/LOGIC_ZERO ),
    .IB(vga_top_vga1_vcounter_Madd__n0000_inst_cy_15),
    .SEL(\vga_top_vga1_vcounter<6>/GROM ),
    .O(\vga_top_vga1_vcounter<6>/CYMUXG )
  );
  X_XOR2 vga_top_vga1_vcounter_Madd__n0000_inst_sum_16 (
    .I0(vga_top_vga1_vcounter_Madd__n0000_inst_cy_15),
    .I1(\vga_top_vga1_vcounter<6>/GROM ),
    .O(vga_top_vga1_vcounter__n0000[7])
  );
  X_BUF \vga_top_vga1_vcounter<6>/CYINIT_1631  (
    .I(vga_top_vga1_vcounter_Madd__n0000_inst_cy_14),
    .O(\vga_top_vga1_vcounter<6>/CYINIT )
  );
  X_ZERO \vga_top_vga1_vcounter<8>/LOGIC_ZERO_1632  (
    .O(\vga_top_vga1_vcounter<8>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_vcounter_Madd__n0000_inst_cy_17_1633 (
    .IA(\vga_top_vga1_vcounter<8>/LOGIC_ZERO ),
    .IB(\vga_top_vga1_vcounter<8>/CYINIT ),
    .SEL(\vga_top_vga1_vcounter<8>/FROM ),
    .O(vga_top_vga1_vcounter_Madd__n0000_inst_cy_17)
  );
  X_XOR2 vga_top_vga1_vcounter_Madd__n0000_inst_sum_17 (
    .I0(\vga_top_vga1_vcounter<8>/CYINIT ),
    .I1(\vga_top_vga1_vcounter<8>/FROM ),
    .O(vga_top_vga1_vcounter__n0000[8])
  );
  defparam \vga_top_vga1_vcounter<8>/F .INIT = 16'hCCCC;
  X_LUT4 \vga_top_vga1_vcounter<8>/F  (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_vcounter[8]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\vga_top_vga1_vcounter<8>/FROM )
  );
  defparam \vga_top_vga1_vcounter<9>_rt_1634 .INIT = 16'hCCCC;
  X_LUT4 \vga_top_vga1_vcounter<9>_rt_1634  (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_vcounter[9]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\vga_top_vga1_vcounter<9>_rt )
  );
  X_XOR2 vga_top_vga1_vcounter_Madd__n0000_inst_sum_18 (
    .I0(vga_top_vga1_vcounter_Madd__n0000_inst_cy_17),
    .I1(\vga_top_vga1_vcounter<9>_rt ),
    .O(vga_top_vga1_vcounter__n0000[9])
  );
  X_BUF \vga_top_vga1_vcounter<8>/CYINIT_1635  (
    .I(vga_top_vga1_vcounter_Madd__n0000_inst_cy_16),
    .O(\vga_top_vga1_vcounter<8>/CYINIT )
  );
  X_ONE \DLX_EXinst_Mcompar__n0059_inst_cy_103/LOGIC_ONE_1636  (
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_103/LOGIC_ONE )
  );
  X_ZERO \DLX_EXinst_Mcompar__n0059_inst_cy_103/LOGIC_ZERO_1637  (
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_103/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0059_inst_cy_102_1638 (
    .IA(\DLX_EXinst_Mcompar__n0059_inst_cy_103/LOGIC_ZERO ),
    .IB(\DLX_EXinst_Mcompar__n0059_inst_cy_103/LOGIC_ONE ),
    .SEL(DLX_EXinst_Mcompar__n0059_inst_lut4_0),
    .O(DLX_EXinst_Mcompar__n0059_inst_cy_102)
  );
  defparam DLX_EXinst_Mcompar__n0059_inst_lut4_01.INIT = 16'h9009;
  X_LUT4 DLX_EXinst_Mcompar__n0059_inst_lut4_01 (
    .ADR0(DLX_IDinst_reg_out_A[0]),
    .ADR1(\DLX_IDinst_Imm[0] ),
    .ADR2(DLX_IDinst_reg_out_A[1]),
    .ADR3(DLX_IDinst_Imm_1_1),
    .O(DLX_EXinst_Mcompar__n0059_inst_lut4_0)
  );
  defparam DLX_EXinst_Mcompar__n0059_inst_lut4_16.INIT = 16'h9009;
  X_LUT4 DLX_EXinst_Mcompar__n0059_inst_lut4_16 (
    .ADR0(DLX_IDinst_reg_out_A[3]),
    .ADR1(DLX_IDinst_Imm_3_1),
    .ADR2(DLX_IDinst_Imm_2_1),
    .ADR3(DLX_IDinst_reg_out_A[2]),
    .O(DLX_EXinst_Mcompar__n0059_inst_lut4_1)
  );
  X_BUF \DLX_EXinst_Mcompar__n0059_inst_cy_103/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0059_inst_cy_103/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0059_inst_cy_103)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0059_inst_cy_103_1639 (
    .IA(\DLX_EXinst_Mcompar__n0059_inst_cy_103/LOGIC_ZERO ),
    .IB(DLX_EXinst_Mcompar__n0059_inst_cy_102),
    .SEL(DLX_EXinst_Mcompar__n0059_inst_lut4_1),
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_103/CYMUXG )
  );
  X_ZERO \DLX_EXinst_Mcompar__n0059_inst_cy_105/LOGIC_ZERO_1640  (
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_105/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0059_inst_cy_104_1641 (
    .IA(\DLX_EXinst_Mcompar__n0059_inst_cy_105/LOGIC_ZERO ),
    .IB(\DLX_EXinst_Mcompar__n0059_inst_cy_105/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0059_inst_lut4_2),
    .O(DLX_EXinst_Mcompar__n0059_inst_cy_104)
  );
  defparam DLX_EXinst_Mcompar__n0059_inst_lut4_21.INIT = 16'h8421;
  X_LUT4 DLX_EXinst_Mcompar__n0059_inst_lut4_21 (
    .ADR0(\DLX_IDinst_Imm[5] ),
    .ADR1(DLX_IDinst_reg_out_A[4]),
    .ADR2(DLX_IDinst_reg_out_A[5]),
    .ADR3(\DLX_IDinst_Imm[4] ),
    .O(DLX_EXinst_Mcompar__n0059_inst_lut4_2)
  );
  defparam DLX_EXinst_Mcompar__n0059_inst_lut4_31.INIT = 16'h8421;
  X_LUT4 DLX_EXinst_Mcompar__n0059_inst_lut4_31 (
    .ADR0(\DLX_IDinst_Imm[7] ),
    .ADR1(DLX_IDinst_reg_out_A[6]),
    .ADR2(DLX_IDinst_reg_out_A[7]),
    .ADR3(\DLX_IDinst_Imm[6] ),
    .O(DLX_EXinst_Mcompar__n0059_inst_lut4_3)
  );
  X_BUF \DLX_EXinst_Mcompar__n0059_inst_cy_105/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0059_inst_cy_105/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0059_inst_cy_105)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0059_inst_cy_105_1642 (
    .IA(\DLX_EXinst_Mcompar__n0059_inst_cy_105/LOGIC_ZERO ),
    .IB(DLX_EXinst_Mcompar__n0059_inst_cy_104),
    .SEL(DLX_EXinst_Mcompar__n0059_inst_lut4_3),
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_105/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0059_inst_cy_105/CYINIT_1643  (
    .I(DLX_EXinst_Mcompar__n0059_inst_cy_103),
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_105/CYINIT )
  );
  X_ZERO \DLX_EXinst_Mcompar__n0059_inst_cy_107/LOGIC_ZERO_1644  (
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_107/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0059_inst_cy_106_1645 (
    .IA(\DLX_EXinst_Mcompar__n0059_inst_cy_107/LOGIC_ZERO ),
    .IB(\DLX_EXinst_Mcompar__n0059_inst_cy_107/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0059_inst_lut4_4),
    .O(DLX_EXinst_Mcompar__n0059_inst_cy_106)
  );
  defparam DLX_EXinst_Mcompar__n0059_inst_lut4_41.INIT = 16'h8421;
  X_LUT4 DLX_EXinst_Mcompar__n0059_inst_lut4_41 (
    .ADR0(DLX_IDinst_reg_out_A[9]),
    .ADR1(\DLX_IDinst_Imm[8] ),
    .ADR2(\DLX_IDinst_Imm[9] ),
    .ADR3(DLX_IDinst_reg_out_A[8]),
    .O(DLX_EXinst_Mcompar__n0059_inst_lut4_4)
  );
  defparam DLX_EXinst_Mcompar__n0059_inst_lut4_51.INIT = 16'h8421;
  X_LUT4 DLX_EXinst_Mcompar__n0059_inst_lut4_51 (
    .ADR0(DLX_IDinst_reg_out_A[11]),
    .ADR1(DLX_IDinst_reg_out_A[10]),
    .ADR2(\DLX_IDinst_Imm[11] ),
    .ADR3(\DLX_IDinst_Imm[10] ),
    .O(DLX_EXinst_Mcompar__n0059_inst_lut4_5)
  );
  X_BUF \DLX_EXinst_Mcompar__n0059_inst_cy_107/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0059_inst_cy_107/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0059_inst_cy_107)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0059_inst_cy_107_1646 (
    .IA(\DLX_EXinst_Mcompar__n0059_inst_cy_107/LOGIC_ZERO ),
    .IB(DLX_EXinst_Mcompar__n0059_inst_cy_106),
    .SEL(DLX_EXinst_Mcompar__n0059_inst_lut4_5),
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_107/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0059_inst_cy_107/CYINIT_1647  (
    .I(DLX_EXinst_Mcompar__n0059_inst_cy_105),
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_107/CYINIT )
  );
  defparam DLX_IDinst_RegFile_28_28_1648.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_28_28_1648 (
    .I(DLX_IDinst_WB_data_eff[28]),
    .CE(DLX_IDinst__n0606),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_28_28)
  );
  X_ZERO \DLX_EXinst_Mcompar__n0059_inst_cy_109/LOGIC_ZERO_1649  (
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_109/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0059_inst_cy_108_1650 (
    .IA(\DLX_EXinst_Mcompar__n0059_inst_cy_109/LOGIC_ZERO ),
    .IB(\DLX_EXinst_Mcompar__n0059_inst_cy_109/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0059_inst_lut4_6),
    .O(DLX_EXinst_Mcompar__n0059_inst_cy_108)
  );
  defparam DLX_EXinst_Mcompar__n0059_inst_lut4_61.INIT = 16'h8421;
  X_LUT4 DLX_EXinst_Mcompar__n0059_inst_lut4_61 (
    .ADR0(DLX_IDinst_reg_out_A[12]),
    .ADR1(\DLX_IDinst_Imm[13] ),
    .ADR2(\DLX_IDinst_Imm[12] ),
    .ADR3(DLX_IDinst_reg_out_A[13]),
    .O(DLX_EXinst_Mcompar__n0059_inst_lut4_6)
  );
  defparam DLX_EXinst_Mcompar__n0059_inst_lut4_71.INIT = 16'h8241;
  X_LUT4 DLX_EXinst_Mcompar__n0059_inst_lut4_71 (
    .ADR0(\DLX_IDinst_Imm[15] ),
    .ADR1(\DLX_IDinst_Imm[14] ),
    .ADR2(DLX_IDinst_reg_out_A[14]),
    .ADR3(DLX_IDinst_reg_out_A[15]),
    .O(DLX_EXinst_Mcompar__n0059_inst_lut4_7)
  );
  X_BUF \DLX_EXinst_Mcompar__n0059_inst_cy_109/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0059_inst_cy_109/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0059_inst_cy_109)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0059_inst_cy_109_1651 (
    .IA(\DLX_EXinst_Mcompar__n0059_inst_cy_109/LOGIC_ZERO ),
    .IB(DLX_EXinst_Mcompar__n0059_inst_cy_108),
    .SEL(DLX_EXinst_Mcompar__n0059_inst_lut4_7),
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_109/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0059_inst_cy_109/CYINIT_1652  (
    .I(DLX_EXinst_Mcompar__n0059_inst_cy_107),
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_109/CYINIT )
  );
  X_ZERO \DLX_EXinst_Mcompar__n0059_inst_cy_111/LOGIC_ZERO_1653  (
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_111/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0059_inst_cy_110_1654 (
    .IA(\DLX_EXinst_Mcompar__n0059_inst_cy_111/LOGIC_ZERO ),
    .IB(\DLX_EXinst_Mcompar__n0059_inst_cy_111/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0059_inst_lut4_8),
    .O(DLX_EXinst_Mcompar__n0059_inst_cy_110)
  );
  defparam DLX_EXinst_Mcompar__n0059_inst_lut4_81.INIT = 16'hA005;
  X_LUT4 DLX_EXinst_Mcompar__n0059_inst_lut4_81 (
    .ADR0(DLX_IDinst_reg_out_A[17]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[16]),
    .ADR3(\DLX_IDinst_Imm[31] ),
    .O(DLX_EXinst_Mcompar__n0059_inst_lut4_8)
  );
  defparam DLX_EXinst_Mcompar__n0059_inst_lut4_91.INIT = 16'hA005;
  X_LUT4 DLX_EXinst_Mcompar__n0059_inst_lut4_91 (
    .ADR0(DLX_IDinst_reg_out_A[19]),
    .ADR1(VCC),
    .ADR2(\DLX_IDinst_Imm[31] ),
    .ADR3(DLX_IDinst_reg_out_A[18]),
    .O(DLX_EXinst_Mcompar__n0059_inst_lut4_9)
  );
  X_BUF \DLX_EXinst_Mcompar__n0059_inst_cy_111/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0059_inst_cy_111/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0059_inst_cy_111)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0059_inst_cy_111_1655 (
    .IA(\DLX_EXinst_Mcompar__n0059_inst_cy_111/LOGIC_ZERO ),
    .IB(DLX_EXinst_Mcompar__n0059_inst_cy_110),
    .SEL(DLX_EXinst_Mcompar__n0059_inst_lut4_9),
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_111/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0059_inst_cy_111/CYINIT_1656  (
    .I(DLX_EXinst_Mcompar__n0059_inst_cy_109),
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_111/CYINIT )
  );
  defparam DLX_IDinst_RegFile_29_12_1657.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_29_12_1657 (
    .I(DLX_IDinst_WB_data_eff[12]),
    .CE(DLX_IDinst__n0608),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_29_12)
  );
  X_ZERO \DLX_IDinst_RegFile_14_12/LOGIC_ZERO_1658  (
    .O(\DLX_IDinst_RegFile_14_12/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0059_inst_cy_112_1659 (
    .IA(\DLX_IDinst_RegFile_14_12/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_14_12/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0059_inst_lut4_10),
    .O(DLX_EXinst_Mcompar__n0059_inst_cy_112)
  );
  defparam DLX_EXinst_Mcompar__n0059_inst_lut4_101.INIT = 16'h8181;
  X_LUT4 DLX_EXinst_Mcompar__n0059_inst_lut4_101 (
    .ADR0(DLX_IDinst_reg_out_A[20]),
    .ADR1(\DLX_IDinst_Imm[31] ),
    .ADR2(DLX_IDinst_reg_out_A[21]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0059_inst_lut4_10)
  );
  defparam DLX_EXinst_Mcompar__n0059_inst_lut4_111.INIT = 16'hC003;
  X_LUT4 DLX_EXinst_Mcompar__n0059_inst_lut4_111 (
    .ADR0(VCC),
    .ADR1(\DLX_IDinst_Imm[31] ),
    .ADR2(DLX_IDinst_reg_out_A[23]),
    .ADR3(DLX_IDinst_reg_out_A[22]),
    .O(DLX_EXinst_Mcompar__n0059_inst_lut4_11)
  );
  X_BUF \DLX_IDinst_RegFile_14_12/COUTUSED  (
    .I(\DLX_IDinst_RegFile_14_12/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0059_inst_cy_113)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0059_inst_cy_113_1660 (
    .IA(\DLX_IDinst_RegFile_14_12/LOGIC_ZERO ),
    .IB(DLX_EXinst_Mcompar__n0059_inst_cy_112),
    .SEL(DLX_EXinst_Mcompar__n0059_inst_lut4_11),
    .O(\DLX_IDinst_RegFile_14_12/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_14_12/CYINIT_1661  (
    .I(DLX_EXinst_Mcompar__n0059_inst_cy_111),
    .O(\DLX_IDinst_RegFile_14_12/CYINIT )
  );
  X_ZERO \DLX_EXinst_Mcompar__n0059_inst_cy_115/LOGIC_ZERO_1662  (
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_115/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0059_inst_cy_114_1663 (
    .IA(\DLX_EXinst_Mcompar__n0059_inst_cy_115/LOGIC_ZERO ),
    .IB(\DLX_EXinst_Mcompar__n0059_inst_cy_115/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0059_inst_lut4_12),
    .O(DLX_EXinst_Mcompar__n0059_inst_cy_114)
  );
  defparam DLX_EXinst_Mcompar__n0059_inst_lut4_121.INIT = 16'hA005;
  X_LUT4 DLX_EXinst_Mcompar__n0059_inst_lut4_121 (
    .ADR0(DLX_IDinst_reg_out_A[25]),
    .ADR1(VCC),
    .ADR2(\DLX_IDinst_Imm[31] ),
    .ADR3(DLX_IDinst_reg_out_A[24]),
    .O(DLX_EXinst_Mcompar__n0059_inst_lut4_12)
  );
  defparam DLX_EXinst_Mcompar__n0059_inst_lut4_131.INIT = 16'hA005;
  X_LUT4 DLX_EXinst_Mcompar__n0059_inst_lut4_131 (
    .ADR0(DLX_IDinst_reg_out_A[27]),
    .ADR1(VCC),
    .ADR2(\DLX_IDinst_Imm[31] ),
    .ADR3(DLX_IDinst_reg_out_A[26]),
    .O(DLX_EXinst_Mcompar__n0059_inst_lut4_13)
  );
  X_BUF \DLX_EXinst_Mcompar__n0059_inst_cy_115/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0059_inst_cy_115/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0059_inst_cy_115)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0059_inst_cy_115_1664 (
    .IA(\DLX_EXinst_Mcompar__n0059_inst_cy_115/LOGIC_ZERO ),
    .IB(DLX_EXinst_Mcompar__n0059_inst_cy_114),
    .SEL(DLX_EXinst_Mcompar__n0059_inst_lut4_13),
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_115/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0059_inst_cy_115/CYINIT_1665  (
    .I(DLX_EXinst_Mcompar__n0059_inst_cy_113),
    .O(\DLX_EXinst_Mcompar__n0059_inst_cy_115/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_30_17/LOGIC_ZERO_1666  (
    .O(\DLX_IDinst_RegFile_30_17/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0059_inst_cy_116_1667 (
    .IA(\DLX_IDinst_RegFile_30_17/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_30_17/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0059_inst_lut4_14),
    .O(DLX_EXinst_Mcompar__n0059_inst_cy_116)
  );
  defparam DLX_EXinst_Mcompar__n0059_inst_lut4_141.INIT = 16'h8811;
  X_LUT4 DLX_EXinst_Mcompar__n0059_inst_lut4_141 (
    .ADR0(DLX_IDinst_reg_out_A[28]),
    .ADR1(\DLX_IDinst_Imm[31] ),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[29]),
    .O(DLX_EXinst_Mcompar__n0059_inst_lut4_14)
  );
  defparam DLX_EXinst_Mcompar__n0059_inst_lut4_151.INIT = 16'h8181;
  X_LUT4 DLX_EXinst_Mcompar__n0059_inst_lut4_151 (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(\DLX_IDinst_Imm[31] ),
    .ADR2(DLX_IDinst_reg_out_A[30]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0059_inst_lut4_15)
  );
  X_BUF \DLX_IDinst_RegFile_30_17/COUTUSED  (
    .I(\DLX_IDinst_RegFile_30_17/CYMUXG ),
    .O(DLX_EXinst__n0059)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0059_inst_cy_117 (
    .IA(\DLX_IDinst_RegFile_30_17/LOGIC_ZERO ),
    .IB(DLX_EXinst_Mcompar__n0059_inst_cy_116),
    .SEL(DLX_EXinst_Mcompar__n0059_inst_lut4_15),
    .O(\DLX_IDinst_RegFile_30_17/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_30_17/CYINIT_1668  (
    .I(DLX_EXinst_Mcompar__n0059_inst_cy_115),
    .O(\DLX_IDinst_RegFile_30_17/CYINIT )
  );
  X_ZERO \DLX_EXinst_Mcompar__n0067_inst_cy_199/LOGIC_ZERO_1669  (
    .O(\DLX_EXinst_Mcompar__n0067_inst_cy_199/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0067_inst_cy_198_1670 (
    .IA(DLX_IDinst_reg_out_A[0]),
    .IB(\DLX_EXinst_Mcompar__n0067_inst_cy_199/LOGIC_ZERO ),
    .SEL(DLX_EXinst_Mcompar__n0067_inst_lut2_134),
    .O(DLX_EXinst_Mcompar__n0067_inst_cy_198)
  );
  defparam DLX_EXinst_Mcompar__n0067_inst_lut2_1341.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0067_inst_lut2_1341 (
    .ADR0(DLX_IDinst_reg_out_A[0]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(\DLX_IDinst_Imm[0] ),
    .O(DLX_EXinst_Mcompar__n0067_inst_lut2_134)
  );
  defparam DLX_EXinst_Mcompar__n0067_inst_lut2_1351.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0067_inst_lut2_1351 (
    .ADR0(DLX_IDinst_reg_out_A[1]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_Imm_1_1),
    .O(DLX_EXinst_Mcompar__n0067_inst_lut2_135)
  );
  X_BUF \DLX_EXinst_Mcompar__n0067_inst_cy_199/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0067_inst_cy_199/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0067_inst_cy_199)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0067_inst_cy_199_1671 (
    .IA(DLX_IDinst_reg_out_A[1]),
    .IB(DLX_EXinst_Mcompar__n0067_inst_cy_198),
    .SEL(DLX_EXinst_Mcompar__n0067_inst_lut2_135),
    .O(\DLX_EXinst_Mcompar__n0067_inst_cy_199/CYMUXG )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0067_inst_cy_200_1672 (
    .IA(DLX_IDinst_reg_out_A[2]),
    .IB(\DLX_IDinst_RegFile_11_3/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0067_inst_lut2_136),
    .O(DLX_EXinst_Mcompar__n0067_inst_cy_200)
  );
  defparam DLX_EXinst_Mcompar__n0067_inst_lut2_1361.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0067_inst_lut2_1361 (
    .ADR0(DLX_IDinst_reg_out_A[2]),
    .ADR1(DLX_IDinst_Imm_2_1),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0067_inst_lut2_136)
  );
  defparam DLX_EXinst_Mcompar__n0067_inst_lut2_1371.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0067_inst_lut2_1371 (
    .ADR0(DLX_IDinst_reg_out_A[3]),
    .ADR1(DLX_IDinst_Imm_3_1),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0067_inst_lut2_137)
  );
  X_BUF \DLX_IDinst_RegFile_11_3/COUTUSED  (
    .I(\DLX_IDinst_RegFile_11_3/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0067_inst_cy_201)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0067_inst_cy_201_1673 (
    .IA(DLX_IDinst_reg_out_A[3]),
    .IB(DLX_EXinst_Mcompar__n0067_inst_cy_200),
    .SEL(DLX_EXinst_Mcompar__n0067_inst_lut2_137),
    .O(\DLX_IDinst_RegFile_11_3/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_11_3/CYINIT_1674  (
    .I(DLX_EXinst_Mcompar__n0067_inst_cy_199),
    .O(\DLX_IDinst_RegFile_11_3/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0067_inst_cy_202_1675 (
    .IA(DLX_IDinst_reg_out_A[4]),
    .IB(\DLX_EXinst_Mcompar__n0067_inst_cy_203/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0067_inst_lut2_138),
    .O(DLX_EXinst_Mcompar__n0067_inst_cy_202)
  );
  defparam DLX_EXinst_Mcompar__n0067_inst_lut2_1381.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0067_inst_lut2_1381 (
    .ADR0(DLX_IDinst_reg_out_A[4]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(\DLX_IDinst_Imm[4] ),
    .O(DLX_EXinst_Mcompar__n0067_inst_lut2_138)
  );
  defparam DLX_EXinst_Mcompar__n0067_inst_lut2_1391.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0067_inst_lut2_1391 (
    .ADR0(DLX_IDinst_reg_out_A[5]),
    .ADR1(\DLX_IDinst_Imm[5] ),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0067_inst_lut2_139)
  );
  X_BUF \DLX_EXinst_Mcompar__n0067_inst_cy_203/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0067_inst_cy_203/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0067_inst_cy_203)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0067_inst_cy_203_1676 (
    .IA(DLX_IDinst_reg_out_A[5]),
    .IB(DLX_EXinst_Mcompar__n0067_inst_cy_202),
    .SEL(DLX_EXinst_Mcompar__n0067_inst_lut2_139),
    .O(\DLX_EXinst_Mcompar__n0067_inst_cy_203/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0067_inst_cy_203/CYINIT_1677  (
    .I(DLX_EXinst_Mcompar__n0067_inst_cy_201),
    .O(\DLX_EXinst_Mcompar__n0067_inst_cy_203/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0067_inst_cy_204_1678 (
    .IA(DLX_IDinst_reg_out_A[6]),
    .IB(\DLX_IDinst_RegFile_14_17/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0067_inst_lut2_140),
    .O(DLX_EXinst_Mcompar__n0067_inst_cy_204)
  );
  defparam DLX_EXinst_Mcompar__n0067_inst_lut2_1401.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0067_inst_lut2_1401 (
    .ADR0(DLX_IDinst_reg_out_A[6]),
    .ADR1(VCC),
    .ADR2(\DLX_IDinst_Imm[6] ),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0067_inst_lut2_140)
  );
  defparam DLX_EXinst_Mcompar__n0067_inst_lut2_1411.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0067_inst_lut2_1411 (
    .ADR0(DLX_IDinst_reg_out_A[7]),
    .ADR1(VCC),
    .ADR2(\DLX_IDinst_Imm[7] ),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0067_inst_lut2_141)
  );
  X_BUF \DLX_IDinst_RegFile_14_17/COUTUSED  (
    .I(\DLX_IDinst_RegFile_14_17/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0067_inst_cy_205)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0067_inst_cy_205_1679 (
    .IA(DLX_IDinst_reg_out_A[7]),
    .IB(DLX_EXinst_Mcompar__n0067_inst_cy_204),
    .SEL(DLX_EXinst_Mcompar__n0067_inst_lut2_141),
    .O(\DLX_IDinst_RegFile_14_17/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_14_17/CYINIT_1680  (
    .I(DLX_EXinst_Mcompar__n0067_inst_cy_203),
    .O(\DLX_IDinst_RegFile_14_17/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0067_inst_cy_206_1681 (
    .IA(DLX_IDinst_reg_out_A[8]),
    .IB(\DLX_EXinst_Mcompar__n0067_inst_cy_207/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0067_inst_lut2_142),
    .O(DLX_EXinst_Mcompar__n0067_inst_cy_206)
  );
  defparam DLX_EXinst_Mcompar__n0067_inst_lut2_1421.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0067_inst_lut2_1421 (
    .ADR0(DLX_IDinst_reg_out_A[8]),
    .ADR1(\DLX_IDinst_Imm[8] ),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0067_inst_lut2_142)
  );
  defparam DLX_EXinst_Mcompar__n0067_inst_lut2_1431.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0067_inst_lut2_1431 (
    .ADR0(DLX_IDinst_reg_out_A[9]),
    .ADR1(VCC),
    .ADR2(\DLX_IDinst_Imm[9] ),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0067_inst_lut2_143)
  );
  X_BUF \DLX_EXinst_Mcompar__n0067_inst_cy_207/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0067_inst_cy_207/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0067_inst_cy_207)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0067_inst_cy_207_1682 (
    .IA(DLX_IDinst_reg_out_A[9]),
    .IB(DLX_EXinst_Mcompar__n0067_inst_cy_206),
    .SEL(DLX_EXinst_Mcompar__n0067_inst_lut2_143),
    .O(\DLX_EXinst_Mcompar__n0067_inst_cy_207/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0067_inst_cy_207/CYINIT_1683  (
    .I(DLX_EXinst_Mcompar__n0067_inst_cy_205),
    .O(\DLX_EXinst_Mcompar__n0067_inst_cy_207/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0067_inst_cy_208_1684 (
    .IA(DLX_IDinst_reg_out_A[10]),
    .IB(\DLX_IDinst_RegFile_30_20/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0067_inst_lut2_144),
    .O(DLX_EXinst_Mcompar__n0067_inst_cy_208)
  );
  defparam DLX_EXinst_Mcompar__n0067_inst_lut2_1441.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0067_inst_lut2_1441 (
    .ADR0(DLX_IDinst_reg_out_A[10]),
    .ADR1(\DLX_IDinst_Imm[10] ),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0067_inst_lut2_144)
  );
  defparam DLX_EXinst_Mcompar__n0067_inst_lut2_1451.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0067_inst_lut2_1451 (
    .ADR0(DLX_IDinst_reg_out_A[11]),
    .ADR1(\DLX_IDinst_Imm[11] ),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0067_inst_lut2_145)
  );
  X_BUF \DLX_IDinst_RegFile_30_20/COUTUSED  (
    .I(\DLX_IDinst_RegFile_30_20/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0067_inst_cy_209)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0067_inst_cy_209_1685 (
    .IA(DLX_IDinst_reg_out_A[11]),
    .IB(DLX_EXinst_Mcompar__n0067_inst_cy_208),
    .SEL(DLX_EXinst_Mcompar__n0067_inst_lut2_145),
    .O(\DLX_IDinst_RegFile_30_20/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_30_20/CYINIT_1686  (
    .I(DLX_EXinst_Mcompar__n0067_inst_cy_207),
    .O(\DLX_IDinst_RegFile_30_20/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0067_inst_cy_210_1687 (
    .IA(DLX_IDinst_reg_out_A[12]),
    .IB(\DLX_EXinst_Mcompar__n0067_inst_cy_211/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0067_inst_lut2_146),
    .O(DLX_EXinst_Mcompar__n0067_inst_cy_210)
  );
  defparam DLX_EXinst_Mcompar__n0067_inst_lut2_1461.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0067_inst_lut2_1461 (
    .ADR0(DLX_IDinst_reg_out_A[12]),
    .ADR1(\DLX_IDinst_Imm[12] ),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0067_inst_lut2_146)
  );
  defparam DLX_EXinst_Mcompar__n0067_inst_lut2_1471.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0067_inst_lut2_1471 (
    .ADR0(DLX_IDinst_reg_out_A[13]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(\DLX_IDinst_Imm[13] ),
    .O(DLX_EXinst_Mcompar__n0067_inst_lut2_147)
  );
  X_BUF \DLX_EXinst_Mcompar__n0067_inst_cy_211/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0067_inst_cy_211/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0067_inst_cy_211)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0067_inst_cy_211_1688 (
    .IA(DLX_IDinst_reg_out_A[13]),
    .IB(DLX_EXinst_Mcompar__n0067_inst_cy_210),
    .SEL(DLX_EXinst_Mcompar__n0067_inst_lut2_147),
    .O(\DLX_EXinst_Mcompar__n0067_inst_cy_211/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0067_inst_cy_211/CYINIT_1689  (
    .I(DLX_EXinst_Mcompar__n0067_inst_cy_209),
    .O(\DLX_EXinst_Mcompar__n0067_inst_cy_211/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0067_inst_cy_212_1690 (
    .IA(DLX_IDinst_reg_out_A[14]),
    .IB(\DLX_IDinst_RegFile_11_27/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0067_inst_lut2_148),
    .O(DLX_EXinst_Mcompar__n0067_inst_cy_212)
  );
  defparam DLX_EXinst_Mcompar__n0067_inst_lut2_1481.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0067_inst_lut2_1481 (
    .ADR0(DLX_IDinst_reg_out_A[14]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(\DLX_IDinst_Imm[14] ),
    .O(DLX_EXinst_Mcompar__n0067_inst_lut2_148)
  );
  defparam DLX_EXinst_Mcompar__n0067_inst_lut2_1491.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0067_inst_lut2_1491 (
    .ADR0(DLX_IDinst_reg_out_A[15]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(\DLX_IDinst_Imm[15] ),
    .O(DLX_EXinst_Mcompar__n0067_inst_lut2_149)
  );
  X_BUF \DLX_IDinst_RegFile_11_27/COUTUSED  (
    .I(\DLX_IDinst_RegFile_11_27/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0067_inst_cy_213)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0067_inst_cy_213_1691 (
    .IA(DLX_IDinst_reg_out_A[15]),
    .IB(DLX_EXinst_Mcompar__n0067_inst_cy_212),
    .SEL(DLX_EXinst_Mcompar__n0067_inst_lut2_149),
    .O(\DLX_IDinst_RegFile_11_27/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_11_27/CYINIT_1692  (
    .I(DLX_EXinst_Mcompar__n0067_inst_cy_211),
    .O(\DLX_IDinst_RegFile_11_27/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0067_inst_cy_214_1693 (
    .IA(DLX_IDinst_reg_out_A[16]),
    .IB(\DLX_EXinst_Mcompar__n0067_inst_cy_215/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0067_inst_lut2_150),
    .O(DLX_EXinst_Mcompar__n0067_inst_cy_214)
  );
  defparam DLX_EXinst_Mcompar__n0067_inst_lut2_1501.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0067_inst_lut2_1501 (
    .ADR0(DLX_IDinst_reg_out_A[16]),
    .ADR1(DLX_IDinst_Imm_31_1),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0067_inst_lut2_150)
  );
  defparam DLX_EXinst_Mcompar__n0067_inst_lut2_1511.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0067_inst_lut2_1511 (
    .ADR0(DLX_IDinst_reg_out_A[17]),
    .ADR1(DLX_IDinst_Imm_31_1),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0067_inst_lut2_151)
  );
  X_BUF \DLX_EXinst_Mcompar__n0067_inst_cy_215/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0067_inst_cy_215/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0067_inst_cy_215)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0067_inst_cy_215_1694 (
    .IA(DLX_IDinst_reg_out_A[17]),
    .IB(DLX_EXinst_Mcompar__n0067_inst_cy_214),
    .SEL(DLX_EXinst_Mcompar__n0067_inst_lut2_151),
    .O(\DLX_EXinst_Mcompar__n0067_inst_cy_215/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0067_inst_cy_215/CYINIT_1695  (
    .I(DLX_EXinst_Mcompar__n0067_inst_cy_213),
    .O(\DLX_EXinst_Mcompar__n0067_inst_cy_215/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0067_inst_cy_216_1696 (
    .IA(DLX_IDinst_reg_out_A[18]),
    .IB(\DLX_IDinst_RegFile_18_3/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0067_inst_lut2_152),
    .O(DLX_EXinst_Mcompar__n0067_inst_cy_216)
  );
  defparam DLX_EXinst_Mcompar__n0067_inst_lut2_1521.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0067_inst_lut2_1521 (
    .ADR0(DLX_IDinst_reg_out_A[18]),
    .ADR1(DLX_IDinst_Imm_31_1),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0067_inst_lut2_152)
  );
  defparam DLX_EXinst_Mcompar__n0067_inst_lut2_1531.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0067_inst_lut2_1531 (
    .ADR0(DLX_IDinst_reg_out_A[19]),
    .ADR1(DLX_IDinst_Imm_31_1),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0067_inst_lut2_153)
  );
  X_BUF \DLX_IDinst_RegFile_18_3/COUTUSED  (
    .I(\DLX_IDinst_RegFile_18_3/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0067_inst_cy_217)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0067_inst_cy_217_1697 (
    .IA(DLX_IDinst_reg_out_A[19]),
    .IB(DLX_EXinst_Mcompar__n0067_inst_cy_216),
    .SEL(DLX_EXinst_Mcompar__n0067_inst_lut2_153),
    .O(\DLX_IDinst_RegFile_18_3/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_18_3/CYINIT_1698  (
    .I(DLX_EXinst_Mcompar__n0067_inst_cy_215),
    .O(\DLX_IDinst_RegFile_18_3/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0067_inst_cy_218_1699 (
    .IA(DLX_IDinst_reg_out_A[20]),
    .IB(\DLX_EXinst_Mcompar__n0067_inst_cy_219/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0067_inst_lut2_154),
    .O(DLX_EXinst_Mcompar__n0067_inst_cy_218)
  );
  defparam DLX_EXinst_Mcompar__n0067_inst_lut2_1541.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0067_inst_lut2_1541 (
    .ADR0(DLX_IDinst_reg_out_A[20]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_Imm_31_1),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0067_inst_lut2_154)
  );
  defparam DLX_EXinst_Mcompar__n0067_inst_lut2_1551.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0067_inst_lut2_1551 (
    .ADR0(DLX_IDinst_reg_out_A[21]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_Imm_31_1),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0067_inst_lut2_155)
  );
  X_BUF \DLX_EXinst_Mcompar__n0067_inst_cy_219/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0067_inst_cy_219/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0067_inst_cy_219)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0067_inst_cy_219_1700 (
    .IA(DLX_IDinst_reg_out_A[21]),
    .IB(DLX_EXinst_Mcompar__n0067_inst_cy_218),
    .SEL(DLX_EXinst_Mcompar__n0067_inst_lut2_155),
    .O(\DLX_EXinst_Mcompar__n0067_inst_cy_219/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0067_inst_cy_219/CYINIT_1701  (
    .I(DLX_EXinst_Mcompar__n0067_inst_cy_217),
    .O(\DLX_EXinst_Mcompar__n0067_inst_cy_219/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0067_inst_cy_220_1702 (
    .IA(DLX_IDinst_reg_out_A[22]),
    .IB(\DLX_IDinst_RegFile_22_26/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0067_inst_lut2_156),
    .O(DLX_EXinst_Mcompar__n0067_inst_cy_220)
  );
  defparam DLX_EXinst_Mcompar__n0067_inst_lut2_1561.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0067_inst_lut2_1561 (
    .ADR0(DLX_IDinst_reg_out_A[22]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_Imm_31_1),
    .O(DLX_EXinst_Mcompar__n0067_inst_lut2_156)
  );
  defparam DLX_EXinst_Mcompar__n0067_inst_lut2_1571.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0067_inst_lut2_1571 (
    .ADR0(DLX_IDinst_reg_out_A[23]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_Imm_31_1),
    .O(DLX_EXinst_Mcompar__n0067_inst_lut2_157)
  );
  X_BUF \DLX_IDinst_RegFile_22_26/COUTUSED  (
    .I(\DLX_IDinst_RegFile_22_26/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0067_inst_cy_221)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0067_inst_cy_221_1703 (
    .IA(DLX_IDinst_reg_out_A[23]),
    .IB(DLX_EXinst_Mcompar__n0067_inst_cy_220),
    .SEL(DLX_EXinst_Mcompar__n0067_inst_lut2_157),
    .O(\DLX_IDinst_RegFile_22_26/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_22_26/CYINIT_1704  (
    .I(DLX_EXinst_Mcompar__n0067_inst_cy_219),
    .O(\DLX_IDinst_RegFile_22_26/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0067_inst_cy_222_1705 (
    .IA(DLX_IDinst_reg_out_A[24]),
    .IB(\DLX_EXinst_Mcompar__n0067_inst_cy_223/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0067_inst_lut2_158),
    .O(DLX_EXinst_Mcompar__n0067_inst_cy_222)
  );
  defparam DLX_EXinst_Mcompar__n0067_inst_lut2_1581.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0067_inst_lut2_1581 (
    .ADR0(DLX_IDinst_reg_out_A[24]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_Imm_31_1),
    .O(DLX_EXinst_Mcompar__n0067_inst_lut2_158)
  );
  defparam DLX_EXinst_Mcompar__n0067_inst_lut2_1591.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0067_inst_lut2_1591 (
    .ADR0(DLX_IDinst_reg_out_A[25]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_Imm_31_1),
    .O(DLX_EXinst_Mcompar__n0067_inst_lut2_159)
  );
  X_BUF \DLX_EXinst_Mcompar__n0067_inst_cy_223/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0067_inst_cy_223/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0067_inst_cy_223)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0067_inst_cy_223_1706 (
    .IA(DLX_IDinst_reg_out_A[25]),
    .IB(DLX_EXinst_Mcompar__n0067_inst_cy_222),
    .SEL(DLX_EXinst_Mcompar__n0067_inst_lut2_159),
    .O(\DLX_EXinst_Mcompar__n0067_inst_cy_223/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0067_inst_cy_223/CYINIT_1707  (
    .I(DLX_EXinst_Mcompar__n0067_inst_cy_221),
    .O(\DLX_EXinst_Mcompar__n0067_inst_cy_223/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0067_inst_cy_224_1708 (
    .IA(DLX_IDinst_reg_out_A[26]),
    .IB(\DLX_IDinst_RegFile_30_13/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0067_inst_lut2_160),
    .O(DLX_EXinst_Mcompar__n0067_inst_cy_224)
  );
  defparam DLX_EXinst_Mcompar__n0067_inst_lut2_1601.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0067_inst_lut2_1601 (
    .ADR0(DLX_IDinst_reg_out_A[26]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_Imm_31_1),
    .O(DLX_EXinst_Mcompar__n0067_inst_lut2_160)
  );
  defparam DLX_EXinst_Mcompar__n0067_inst_lut2_1611.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0067_inst_lut2_1611 (
    .ADR0(DLX_IDinst_reg_out_A[27]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_Imm_31_1),
    .O(DLX_EXinst_Mcompar__n0067_inst_lut2_161)
  );
  X_BUF \DLX_IDinst_RegFile_30_13/COUTUSED  (
    .I(\DLX_IDinst_RegFile_30_13/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0067_inst_cy_225)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0067_inst_cy_225_1709 (
    .IA(DLX_IDinst_reg_out_A[27]),
    .IB(DLX_EXinst_Mcompar__n0067_inst_cy_224),
    .SEL(DLX_EXinst_Mcompar__n0067_inst_lut2_161),
    .O(\DLX_IDinst_RegFile_30_13/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_30_13/CYINIT_1710  (
    .I(DLX_EXinst_Mcompar__n0067_inst_cy_223),
    .O(\DLX_IDinst_RegFile_30_13/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0067_inst_cy_226_1711 (
    .IA(DLX_IDinst_reg_out_A[28]),
    .IB(\DLX_EXinst_Mcompar__n0067_inst_cy_227/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0067_inst_lut2_162),
    .O(DLX_EXinst_Mcompar__n0067_inst_cy_226)
  );
  defparam DLX_EXinst_Mcompar__n0067_inst_lut2_1621.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0067_inst_lut2_1621 (
    .ADR0(DLX_IDinst_reg_out_A[28]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_Imm_31_1),
    .O(DLX_EXinst_Mcompar__n0067_inst_lut2_162)
  );
  defparam DLX_EXinst_Mcompar__n0067_inst_lut2_1631.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0067_inst_lut2_1631 (
    .ADR0(DLX_IDinst_reg_out_A[29]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_Imm_31_1),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0067_inst_lut2_163)
  );
  X_BUF \DLX_EXinst_Mcompar__n0067_inst_cy_227/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0067_inst_cy_227/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0067_inst_cy_227)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0067_inst_cy_227_1712 (
    .IA(DLX_IDinst_reg_out_A[29]),
    .IB(DLX_EXinst_Mcompar__n0067_inst_cy_226),
    .SEL(DLX_EXinst_Mcompar__n0067_inst_lut2_163),
    .O(\DLX_EXinst_Mcompar__n0067_inst_cy_227/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0067_inst_cy_227/CYINIT_1713  (
    .I(DLX_EXinst_Mcompar__n0067_inst_cy_225),
    .O(\DLX_EXinst_Mcompar__n0067_inst_cy_227/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0067_inst_cy_228_1714 (
    .IA(DLX_IDinst_reg_out_A[30]),
    .IB(\DLX_EXinst_Mcompar__n0067_inst_cy_228/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0067_inst_lut2_164),
    .O(\DLX_EXinst_Mcompar__n0067_inst_cy_228/CYMUXF )
  );
  defparam DLX_EXinst_Mcompar__n0067_inst_lut2_1641.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0067_inst_lut2_1641 (
    .ADR0(DLX_IDinst_reg_out_A[30]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_Imm_31_1),
    .O(DLX_EXinst_Mcompar__n0067_inst_lut2_164)
  );
  X_BUF \DLX_EXinst_Mcompar__n0067_inst_cy_228/XBUSED  (
    .I(\DLX_EXinst_Mcompar__n0067_inst_cy_228/CYMUXF ),
    .O(DLX_EXinst_Mcompar__n0067_inst_cy_228)
  );
  X_BUF \DLX_EXinst_Mcompar__n0067_inst_cy_228/CYINIT_1715  (
    .I(DLX_EXinst_Mcompar__n0067_inst_cy_227),
    .O(\DLX_EXinst_Mcompar__n0067_inst_cy_228/CYINIT )
  );
  X_ZERO \vga_top_vga1_gridvcounter<0>/LOGIC_ZERO_1716  (
    .O(\vga_top_vga1_gridvcounter<0>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_0_1717 (
    .IA(GLOBAL_LOGIC1),
    .IB(\vga_top_vga1_gridvcounter<0>/LOGIC_ZERO ),
    .SEL(vga_top_vga1_gridvcounter_Madd__n0000_inst_lut2_0),
    .O(vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_0)
  );
  defparam vga_top_vga1_gridvcounter_Madd__n0000_inst_lut2_01.INIT = 16'h3333;
  X_LUT4 vga_top_vga1_gridvcounter_Madd__n0000_inst_lut2_01 (
    .ADR0(GLOBAL_LOGIC1),
    .ADR1(vga_top_vga1_gridvcounter[0]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(vga_top_vga1_gridvcounter_Madd__n0000_inst_lut2_0)
  );
  defparam \vga_top_vga1_gridvcounter<0>/G .INIT = 16'hF0F0;
  X_LUT4 \vga_top_vga1_gridvcounter<0>/G  (
    .ADR0(GLOBAL_LOGIC0),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_gridvcounter[1]),
    .ADR3(VCC),
    .O(\vga_top_vga1_gridvcounter<0>/GROM )
  );
  X_BUF \vga_top_vga1_gridvcounter<0>/COUTUSED  (
    .I(\vga_top_vga1_gridvcounter<0>/CYMUXG ),
    .O(vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_1)
  );
  X_MUX2 vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_1_1718 (
    .IA(GLOBAL_LOGIC0),
    .IB(vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_0),
    .SEL(\vga_top_vga1_gridvcounter<0>/GROM ),
    .O(\vga_top_vga1_gridvcounter<0>/CYMUXG )
  );
  X_XOR2 vga_top_vga1_gridvcounter_Madd__n0000_inst_sum_1 (
    .I0(vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_0),
    .I1(\vga_top_vga1_gridvcounter<0>/GROM ),
    .O(vga_top_vga1_gridvcounter__n0000[1])
  );
  X_ZERO \vga_top_vga1_gridvcounter<2>/LOGIC_ZERO_1719  (
    .O(\vga_top_vga1_gridvcounter<2>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_2_1720 (
    .IA(\vga_top_vga1_gridvcounter<2>/LOGIC_ZERO ),
    .IB(\vga_top_vga1_gridvcounter<2>/CYINIT ),
    .SEL(\vga_top_vga1_gridvcounter<2>/FROM ),
    .O(vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_2)
  );
  X_XOR2 vga_top_vga1_gridvcounter_Madd__n0000_inst_sum_2 (
    .I0(\vga_top_vga1_gridvcounter<2>/CYINIT ),
    .I1(\vga_top_vga1_gridvcounter<2>/FROM ),
    .O(vga_top_vga1_gridvcounter__n0000[2])
  );
  defparam \vga_top_vga1_gridvcounter<2>/F .INIT = 16'hCCCC;
  X_LUT4 \vga_top_vga1_gridvcounter<2>/F  (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_gridvcounter[2]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\vga_top_vga1_gridvcounter<2>/FROM )
  );
  defparam \vga_top_vga1_gridvcounter<2>/G .INIT = 16'hF0F0;
  X_LUT4 \vga_top_vga1_gridvcounter<2>/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_gridvcounter[3]),
    .ADR3(VCC),
    .O(\vga_top_vga1_gridvcounter<2>/GROM )
  );
  X_BUF \vga_top_vga1_gridvcounter<2>/COUTUSED  (
    .I(\vga_top_vga1_gridvcounter<2>/CYMUXG ),
    .O(vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_3)
  );
  X_MUX2 vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_3_1721 (
    .IA(\vga_top_vga1_gridvcounter<2>/LOGIC_ZERO ),
    .IB(vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_2),
    .SEL(\vga_top_vga1_gridvcounter<2>/GROM ),
    .O(\vga_top_vga1_gridvcounter<2>/CYMUXG )
  );
  X_XOR2 vga_top_vga1_gridvcounter_Madd__n0000_inst_sum_3 (
    .I0(vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_2),
    .I1(\vga_top_vga1_gridvcounter<2>/GROM ),
    .O(vga_top_vga1_gridvcounter__n0000[3])
  );
  X_BUF \vga_top_vga1_gridvcounter<2>/CYINIT_1722  (
    .I(vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_1),
    .O(\vga_top_vga1_gridvcounter<2>/CYINIT )
  );
  X_ZERO \vga_top_vga1_gridvcounter<4>/LOGIC_ZERO_1723  (
    .O(\vga_top_vga1_gridvcounter<4>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_4_1724 (
    .IA(\vga_top_vga1_gridvcounter<4>/LOGIC_ZERO ),
    .IB(\vga_top_vga1_gridvcounter<4>/CYINIT ),
    .SEL(\vga_top_vga1_gridvcounter<4>/FROM ),
    .O(vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_4)
  );
  X_XOR2 vga_top_vga1_gridvcounter_Madd__n0000_inst_sum_4 (
    .I0(\vga_top_vga1_gridvcounter<4>/CYINIT ),
    .I1(\vga_top_vga1_gridvcounter<4>/FROM ),
    .O(vga_top_vga1_gridvcounter__n0000[4])
  );
  defparam \vga_top_vga1_gridvcounter<4>/F .INIT = 16'hCCCC;
  X_LUT4 \vga_top_vga1_gridvcounter<4>/F  (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_gridvcounter[4]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\vga_top_vga1_gridvcounter<4>/FROM )
  );
  defparam \vga_top_vga1_gridvcounter<4>/G .INIT = 16'hAAAA;
  X_LUT4 \vga_top_vga1_gridvcounter<4>/G  (
    .ADR0(vga_top_vga1_gridvcounter[5]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\vga_top_vga1_gridvcounter<4>/GROM )
  );
  X_BUF \vga_top_vga1_gridvcounter<4>/COUTUSED  (
    .I(\vga_top_vga1_gridvcounter<4>/CYMUXG ),
    .O(vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_5)
  );
  X_MUX2 vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_5_1725 (
    .IA(\vga_top_vga1_gridvcounter<4>/LOGIC_ZERO ),
    .IB(vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_4),
    .SEL(\vga_top_vga1_gridvcounter<4>/GROM ),
    .O(\vga_top_vga1_gridvcounter<4>/CYMUXG )
  );
  X_XOR2 vga_top_vga1_gridvcounter_Madd__n0000_inst_sum_5 (
    .I0(vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_4),
    .I1(\vga_top_vga1_gridvcounter<4>/GROM ),
    .O(vga_top_vga1_gridvcounter__n0000[5])
  );
  X_BUF \vga_top_vga1_gridvcounter<4>/CYINIT_1726  (
    .I(vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_3),
    .O(\vga_top_vga1_gridvcounter<4>/CYINIT )
  );
  X_ZERO \vga_top_vga1_gridvcounter<6>/LOGIC_ZERO_1727  (
    .O(\vga_top_vga1_gridvcounter<6>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_6_1728 (
    .IA(\vga_top_vga1_gridvcounter<6>/LOGIC_ZERO ),
    .IB(\vga_top_vga1_gridvcounter<6>/CYINIT ),
    .SEL(\vga_top_vga1_gridvcounter<6>/FROM ),
    .O(vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_6)
  );
  X_XOR2 vga_top_vga1_gridvcounter_Madd__n0000_inst_sum_6 (
    .I0(\vga_top_vga1_gridvcounter<6>/CYINIT ),
    .I1(\vga_top_vga1_gridvcounter<6>/FROM ),
    .O(vga_top_vga1_gridvcounter__n0000[6])
  );
  defparam \vga_top_vga1_gridvcounter<6>/F .INIT = 16'hAAAA;
  X_LUT4 \vga_top_vga1_gridvcounter<6>/F  (
    .ADR0(vga_top_vga1_gridvcounter[6]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\vga_top_vga1_gridvcounter<6>/FROM )
  );
  defparam \vga_top_vga1_gridvcounter<6>/G .INIT = 16'hF0F0;
  X_LUT4 \vga_top_vga1_gridvcounter<6>/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_gridvcounter[7]),
    .ADR3(VCC),
    .O(\vga_top_vga1_gridvcounter<6>/GROM )
  );
  X_BUF \vga_top_vga1_gridvcounter<6>/COUTUSED  (
    .I(\vga_top_vga1_gridvcounter<6>/CYMUXG ),
    .O(vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_7)
  );
  X_MUX2 vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_7_1729 (
    .IA(\vga_top_vga1_gridvcounter<6>/LOGIC_ZERO ),
    .IB(vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_6),
    .SEL(\vga_top_vga1_gridvcounter<6>/GROM ),
    .O(\vga_top_vga1_gridvcounter<6>/CYMUXG )
  );
  X_XOR2 vga_top_vga1_gridvcounter_Madd__n0000_inst_sum_7 (
    .I0(vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_6),
    .I1(\vga_top_vga1_gridvcounter<6>/GROM ),
    .O(vga_top_vga1_gridvcounter__n0000[7])
  );
  X_BUF \vga_top_vga1_gridvcounter<6>/CYINIT_1730  (
    .I(vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_5),
    .O(\vga_top_vga1_gridvcounter<6>/CYINIT )
  );
  X_XOR2 vga_top_vga1_gridvcounter_Madd__n0000_inst_sum_8 (
    .I0(\vga_top_vga1_gridvcounter<8>/CYINIT ),
    .I1(\vga_top_vga1_gridvcounter<8>_rt ),
    .O(vga_top_vga1_gridvcounter__n0000[8])
  );
  defparam \vga_top_vga1_gridvcounter<8>_rt_1731 .INIT = 16'hCCCC;
  X_LUT4 \vga_top_vga1_gridvcounter<8>_rt_1731  (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_gridvcounter[8]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\vga_top_vga1_gridvcounter<8>_rt )
  );
  X_BUF \vga_top_vga1_gridvcounter<8>/CYINIT_1732  (
    .I(vga_top_vga1_gridvcounter_Madd__n0000_inst_cy_7),
    .O(\vga_top_vga1_gridvcounter<8>/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_30_27/LOGIC_ZERO_1733  (
    .O(\DLX_IDinst_RegFile_30_27/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_166_1734 (
    .IA(DLX_IDinst_reg_out_A[0]),
    .IB(\DLX_IDinst_RegFile_30_27/LOGIC_ZERO ),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_102),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_166)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1021.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1021 (
    .ADR0(DLX_IDinst_reg_out_A[0]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[0]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_102)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1031.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1031 (
    .ADR0(DLX_IDinst_reg_out_A[1]),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_103)
  );
  X_BUF \DLX_IDinst_RegFile_30_27/COUTUSED  (
    .I(\DLX_IDinst_RegFile_30_27/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_167)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_167_1735 (
    .IA(DLX_IDinst_reg_out_A[1]),
    .IB(DLX_EXinst_Mcompar__n0091_inst_cy_166),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_103),
    .O(\DLX_IDinst_RegFile_30_27/CYMUXG )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_168_1736 (
    .IA(DLX_IDinst_reg_out_A[2]),
    .IB(\DLX_EXinst_Mcompar__n0091_inst_cy_169/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_104),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_168)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1041.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1041 (
    .ADR0(DLX_IDinst_reg_out_A[2]),
    .ADR1(DLX_IDinst_reg_out_B_2_1),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_104)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1051.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1051 (
    .ADR0(DLX_IDinst_reg_out_A[3]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B_3_1),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_105)
  );
  X_BUF \DLX_EXinst_Mcompar__n0091_inst_cy_169/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0091_inst_cy_169/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_169)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_169_1737 (
    .IA(DLX_IDinst_reg_out_A[3]),
    .IB(DLX_EXinst_Mcompar__n0091_inst_cy_168),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_105),
    .O(\DLX_EXinst_Mcompar__n0091_inst_cy_169/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0091_inst_cy_169/CYINIT_1738  (
    .I(DLX_EXinst_Mcompar__n0091_inst_cy_167),
    .O(\DLX_EXinst_Mcompar__n0091_inst_cy_169/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_170_1739 (
    .IA(DLX_IDinst_reg_out_A[4]),
    .IB(\DLX_IDinst_RegFile_22_30/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_106),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_170)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1061.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1061 (
    .ADR0(DLX_IDinst_reg_out_A[4]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[4]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_106)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1071.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1071 (
    .ADR0(DLX_IDinst_reg_out_A[5]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[5]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_107)
  );
  X_BUF \DLX_IDinst_RegFile_22_30/COUTUSED  (
    .I(\DLX_IDinst_RegFile_22_30/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_171)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_171_1740 (
    .IA(DLX_IDinst_reg_out_A[5]),
    .IB(DLX_EXinst_Mcompar__n0091_inst_cy_170),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_107),
    .O(\DLX_IDinst_RegFile_22_30/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_22_30/CYINIT_1741  (
    .I(DLX_EXinst_Mcompar__n0091_inst_cy_169),
    .O(\DLX_IDinst_RegFile_22_30/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_172_1742 (
    .IA(DLX_IDinst_reg_out_A[6]),
    .IB(\DLX_EXinst_Mcompar__n0091_inst_cy_173/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_108),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_172)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1081.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1081 (
    .ADR0(DLX_IDinst_reg_out_A[6]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[6]),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_108)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1091.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1091 (
    .ADR0(DLX_IDinst_reg_out_A[7]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[7]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_109)
  );
  X_BUF \DLX_EXinst_Mcompar__n0091_inst_cy_173/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0091_inst_cy_173/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_173)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_173_1743 (
    .IA(DLX_IDinst_reg_out_A[7]),
    .IB(DLX_EXinst_Mcompar__n0091_inst_cy_172),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_109),
    .O(\DLX_EXinst_Mcompar__n0091_inst_cy_173/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0091_inst_cy_173/CYINIT_1744  (
    .I(DLX_EXinst_Mcompar__n0091_inst_cy_171),
    .O(\DLX_EXinst_Mcompar__n0091_inst_cy_173/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_174_1745 (
    .IA(DLX_IDinst_reg_out_A[8]),
    .IB(\DLX_IDinst_RegFile_1_6/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_110),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_174)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1101.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1101 (
    .ADR0(DLX_IDinst_reg_out_A[8]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[8]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_110)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1111.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1111 (
    .ADR0(DLX_IDinst_reg_out_A[9]),
    .ADR1(DLX_IDinst_reg_out_B[9]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_111)
  );
  X_BUF \DLX_IDinst_RegFile_1_6/COUTUSED  (
    .I(\DLX_IDinst_RegFile_1_6/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_175)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_175_1746 (
    .IA(DLX_IDinst_reg_out_A[9]),
    .IB(DLX_EXinst_Mcompar__n0091_inst_cy_174),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_111),
    .O(\DLX_IDinst_RegFile_1_6/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_1_6/CYINIT_1747  (
    .I(DLX_EXinst_Mcompar__n0091_inst_cy_173),
    .O(\DLX_IDinst_RegFile_1_6/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_176_1748 (
    .IA(DLX_IDinst_reg_out_A[10]),
    .IB(\DLX_EXinst_Mcompar__n0091_inst_cy_177/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_112),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_176)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1121.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1121 (
    .ADR0(DLX_IDinst_reg_out_A[10]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[10]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_112)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1131.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1131 (
    .ADR0(DLX_IDinst_reg_out_A[11]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[11]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_113)
  );
  X_BUF \DLX_EXinst_Mcompar__n0091_inst_cy_177/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0091_inst_cy_177/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_177)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_177_1749 (
    .IA(DLX_IDinst_reg_out_A[11]),
    .IB(DLX_EXinst_Mcompar__n0091_inst_cy_176),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_113),
    .O(\DLX_EXinst_Mcompar__n0091_inst_cy_177/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0091_inst_cy_177/CYINIT_1750  (
    .I(DLX_EXinst_Mcompar__n0091_inst_cy_175),
    .O(\DLX_EXinst_Mcompar__n0091_inst_cy_177/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_178_1751 (
    .IA(DLX_IDinst_reg_out_A[12]),
    .IB(\DLX_IDinst_RegFile_30_22/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_114),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_178)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1141.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1141 (
    .ADR0(DLX_IDinst_reg_out_A[12]),
    .ADR1(DLX_IDinst_reg_out_B[12]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_114)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1151.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1151 (
    .ADR0(DLX_IDinst_reg_out_A[13]),
    .ADR1(DLX_IDinst_reg_out_B[13]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_115)
  );
  X_BUF \DLX_IDinst_RegFile_30_22/COUTUSED  (
    .I(\DLX_IDinst_RegFile_30_22/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_179)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_179_1752 (
    .IA(DLX_IDinst_reg_out_A[13]),
    .IB(DLX_EXinst_Mcompar__n0091_inst_cy_178),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_115),
    .O(\DLX_IDinst_RegFile_30_22/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_30_22/CYINIT_1753  (
    .I(DLX_EXinst_Mcompar__n0091_inst_cy_177),
    .O(\DLX_IDinst_RegFile_30_22/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_180_1754 (
    .IA(DLX_IDinst_reg_out_A[14]),
    .IB(\DLX_EXinst_Mcompar__n0091_inst_cy_181/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_116),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_180)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1161.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1161 (
    .ADR0(DLX_IDinst_reg_out_A[14]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[14]),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_116)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1171.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1171 (
    .ADR0(DLX_IDinst_reg_out_A[15]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[15]),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_117)
  );
  X_BUF \DLX_EXinst_Mcompar__n0091_inst_cy_181/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0091_inst_cy_181/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_181)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_181_1755 (
    .IA(DLX_IDinst_reg_out_A[15]),
    .IB(DLX_EXinst_Mcompar__n0091_inst_cy_180),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_117),
    .O(\DLX_EXinst_Mcompar__n0091_inst_cy_181/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0091_inst_cy_181/CYINIT_1756  (
    .I(DLX_EXinst_Mcompar__n0091_inst_cy_179),
    .O(\DLX_EXinst_Mcompar__n0091_inst_cy_181/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_182_1757 (
    .IA(DLX_IDinst_reg_out_A[16]),
    .IB(\DLX_IDinst_RegFile_30_18/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_118),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_182)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1181.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1181 (
    .ADR0(DLX_IDinst_reg_out_A[16]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[16]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_118)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1191.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1191 (
    .ADR0(DLX_IDinst_reg_out_A[17]),
    .ADR1(DLX_IDinst_reg_out_B[17]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_119)
  );
  X_BUF \DLX_IDinst_RegFile_30_18/COUTUSED  (
    .I(\DLX_IDinst_RegFile_30_18/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_183)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_183_1758 (
    .IA(DLX_IDinst_reg_out_A[17]),
    .IB(DLX_EXinst_Mcompar__n0091_inst_cy_182),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_119),
    .O(\DLX_IDinst_RegFile_30_18/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_30_18/CYINIT_1759  (
    .I(DLX_EXinst_Mcompar__n0091_inst_cy_181),
    .O(\DLX_IDinst_RegFile_30_18/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_184_1760 (
    .IA(DLX_IDinst_reg_out_A[18]),
    .IB(\DLX_EXinst_Mcompar__n0091_inst_cy_185/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_120),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_184)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1201.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1201 (
    .ADR0(DLX_IDinst_reg_out_A[18]),
    .ADR1(DLX_IDinst_reg_out_B[18]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_120)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1211.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1211 (
    .ADR0(DLX_IDinst_reg_out_A[19]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[19]),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_121)
  );
  X_BUF \DLX_EXinst_Mcompar__n0091_inst_cy_185/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0091_inst_cy_185/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_185)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_185_1761 (
    .IA(DLX_IDinst_reg_out_A[19]),
    .IB(DLX_EXinst_Mcompar__n0091_inst_cy_184),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_121),
    .O(\DLX_EXinst_Mcompar__n0091_inst_cy_185/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0091_inst_cy_185/CYINIT_1762  (
    .I(DLX_EXinst_Mcompar__n0091_inst_cy_183),
    .O(\DLX_EXinst_Mcompar__n0091_inst_cy_185/CYINIT )
  );
  defparam DLX_IDinst_RegFile_29_20_1763.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_29_20_1763 (
    .I(DLX_IDinst_WB_data_eff[20]),
    .CE(DLX_IDinst__n0608),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_29_20)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_186_1764 (
    .IA(DLX_IDinst_reg_out_A[20]),
    .IB(\DLX_IDinst_RegFile_22_23/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_122),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_186)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1221.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1221 (
    .ADR0(DLX_IDinst_reg_out_A[20]),
    .ADR1(DLX_IDinst_reg_out_B[20]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_122)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1231.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1231 (
    .ADR0(DLX_IDinst_reg_out_A[21]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[21]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_123)
  );
  X_BUF \DLX_IDinst_RegFile_22_23/COUTUSED  (
    .I(\DLX_IDinst_RegFile_22_23/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_187)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_187_1765 (
    .IA(DLX_IDinst_reg_out_A[21]),
    .IB(DLX_EXinst_Mcompar__n0091_inst_cy_186),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_123),
    .O(\DLX_IDinst_RegFile_22_23/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_22_23/CYINIT_1766  (
    .I(DLX_EXinst_Mcompar__n0091_inst_cy_185),
    .O(\DLX_IDinst_RegFile_22_23/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_188_1767 (
    .IA(DLX_IDinst_reg_out_A[22]),
    .IB(\DLX_EXinst_Mcompar__n0091_inst_cy_189/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_124),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_188)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1241.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1241 (
    .ADR0(DLX_IDinst_reg_out_A[22]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[22]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_124)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1251.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1251 (
    .ADR0(DLX_IDinst_reg_out_A[23]),
    .ADR1(DLX_IDinst_reg_out_B[23]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_125)
  );
  X_BUF \DLX_EXinst_Mcompar__n0091_inst_cy_189/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0091_inst_cy_189/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_189)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_189_1768 (
    .IA(DLX_IDinst_reg_out_A[23]),
    .IB(DLX_EXinst_Mcompar__n0091_inst_cy_188),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_125),
    .O(\DLX_EXinst_Mcompar__n0091_inst_cy_189/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0091_inst_cy_189/CYINIT_1769  (
    .I(DLX_EXinst_Mcompar__n0091_inst_cy_187),
    .O(\DLX_EXinst_Mcompar__n0091_inst_cy_189/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_190_1770 (
    .IA(DLX_IDinst_reg_out_A[24]),
    .IB(\DLX_IDinst_RegFile_15_11/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_126),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_190)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1261.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1261 (
    .ADR0(DLX_IDinst_reg_out_A[24]),
    .ADR1(DLX_IDinst_reg_out_B[24]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_126)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1271.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1271 (
    .ADR0(DLX_IDinst_reg_out_A[25]),
    .ADR1(DLX_IDinst_reg_out_B[25]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_127)
  );
  X_BUF \DLX_IDinst_RegFile_15_11/COUTUSED  (
    .I(\DLX_IDinst_RegFile_15_11/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_191)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_191_1771 (
    .IA(DLX_IDinst_reg_out_A[25]),
    .IB(DLX_EXinst_Mcompar__n0091_inst_cy_190),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_127),
    .O(\DLX_IDinst_RegFile_15_11/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_15_11/CYINIT_1772  (
    .I(DLX_EXinst_Mcompar__n0091_inst_cy_189),
    .O(\DLX_IDinst_RegFile_15_11/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_192_1773 (
    .IA(DLX_IDinst_reg_out_A[26]),
    .IB(\DLX_EXinst_Mcompar__n0091_inst_cy_193/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_128),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_192)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1281.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1281 (
    .ADR0(DLX_IDinst_reg_out_A[26]),
    .ADR1(DLX_IDinst_reg_out_B[26]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_128)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1291.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1291 (
    .ADR0(DLX_IDinst_reg_out_A[27]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[27]),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_129)
  );
  X_BUF \DLX_EXinst_Mcompar__n0091_inst_cy_193/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0091_inst_cy_193/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_193)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_193_1774 (
    .IA(DLX_IDinst_reg_out_A[27]),
    .IB(DLX_EXinst_Mcompar__n0091_inst_cy_192),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_129),
    .O(\DLX_EXinst_Mcompar__n0091_inst_cy_193/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0091_inst_cy_193/CYINIT_1775  (
    .I(DLX_EXinst_Mcompar__n0091_inst_cy_191),
    .O(\DLX_EXinst_Mcompar__n0091_inst_cy_193/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_194_1776 (
    .IA(DLX_IDinst_reg_out_A[28]),
    .IB(\DLX_IDinst_RegFile_3_6/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_130),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_194)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1301.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1301 (
    .ADR0(DLX_IDinst_reg_out_A[28]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[28]),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_130)
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1311.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1311 (
    .ADR0(DLX_IDinst_reg_out_A[29]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[29]),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_131)
  );
  X_BUF \DLX_IDinst_RegFile_3_6/COUTUSED  (
    .I(\DLX_IDinst_RegFile_3_6/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_195)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_195_1777 (
    .IA(DLX_IDinst_reg_out_A[29]),
    .IB(DLX_EXinst_Mcompar__n0091_inst_cy_194),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_131),
    .O(\DLX_IDinst_RegFile_3_6/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_3_6/CYINIT_1778  (
    .I(DLX_EXinst_Mcompar__n0091_inst_cy_193),
    .O(\DLX_IDinst_RegFile_3_6/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0091_inst_cy_196_1779 (
    .IA(DLX_IDinst_reg_out_A[30]),
    .IB(\DLX_EXinst_mem_to_reg_EX/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0091_inst_lut2_132),
    .O(\DLX_EXinst_mem_to_reg_EX/CYMUXF )
  );
  defparam DLX_EXinst_Mcompar__n0091_inst_lut2_1321.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0091_inst_lut2_1321 (
    .ADR0(DLX_IDinst_reg_out_A[30]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[30]),
    .O(DLX_EXinst_Mcompar__n0091_inst_lut2_132)
  );
  defparam \DLX_EXinst__n0008<30>1 .INIT = 16'h8888;
  X_LUT4 \DLX_EXinst__n0008<30>1  (
    .ADR0(DLX_IDinst_reg_out_B[30]),
    .ADR1(DLX_EXinst_N72746),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst__n0008[30])
  );
  X_BUF \DLX_EXinst_mem_to_reg_EX/XBUSED  (
    .I(\DLX_EXinst_mem_to_reg_EX/CYMUXF ),
    .O(DLX_EXinst_Mcompar__n0091_inst_cy_196)
  );
  X_BUF \DLX_EXinst_mem_to_reg_EX/CYINIT_1780  (
    .I(DLX_EXinst_Mcompar__n0091_inst_cy_195),
    .O(\DLX_EXinst_mem_to_reg_EX/CYINIT )
  );
  X_ONE \DLX_IDinst_RegFile_23_21/LOGIC_ONE_1781  (
    .O(\DLX_IDinst_RegFile_23_21/LOGIC_ONE )
  );
  X_MUX2 DLX_IDinst_Msub__n0157_inst_cy_265_1782 (
    .IA(DLX_IDinst_Madd__n0158_inst_lut2_230),
    .IB(\DLX_IDinst_RegFile_23_21/CYINIT ),
    .SEL(DLX_IDinst_Msub__n0157_inst_lut2_198),
    .O(DLX_IDinst_Msub__n0157_inst_cy_265)
  );
  X_XOR2 DLX_IDinst_Msub__n0157_inst_sum_102 (
    .I0(\DLX_IDinst_RegFile_23_21/CYINIT ),
    .I1(DLX_IDinst_Msub__n0157_inst_lut2_198),
    .O(\DLX_IDinst_RegFile_23_21/XORF )
  );
  defparam DLX_IDinst_Msub__n0157_inst_lut2_1981.INIT = 16'hC3C3;
  X_LUT4 DLX_IDinst_Msub__n0157_inst_lut2_1981 (
    .ADR0(DLX_IDinst_Madd__n0158_inst_lut2_230),
    .ADR1(DLX_IDinst_jtarget[0]),
    .ADR2(DLX_IFinst_NPC[0]),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0157_inst_lut2_198)
  );
  defparam DLX_IDinst_Msub__n0157_inst_lut2_1991.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0157_inst_lut2_1991 (
    .ADR0(DLX_IDinst__n0158[1]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0157_inst_lut2_199)
  );
  X_BUF \DLX_IDinst_RegFile_23_21/COUTUSED  (
    .I(\DLX_IDinst_RegFile_23_21/CYMUXG ),
    .O(DLX_IDinst_Msub__n0157_inst_cy_266)
  );
  X_BUF \DLX_IDinst_RegFile_23_21/XUSED  (
    .I(\DLX_IDinst_RegFile_23_21/XORF ),
    .O(DLX_IDinst__n0157[0])
  );
  X_BUF \DLX_IDinst_RegFile_23_21/YUSED  (
    .I(\DLX_IDinst_RegFile_23_21/XORG ),
    .O(DLX_IDinst__n0157[1])
  );
  X_MUX2 DLX_IDinst_Msub__n0157_inst_cy_266_1783 (
    .IA(DLX_IDinst__n0158[1]),
    .IB(DLX_IDinst_Msub__n0157_inst_cy_265),
    .SEL(DLX_IDinst_Msub__n0157_inst_lut2_199),
    .O(\DLX_IDinst_RegFile_23_21/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Msub__n0157_inst_sum_103 (
    .I0(DLX_IDinst_Msub__n0157_inst_cy_265),
    .I1(DLX_IDinst_Msub__n0157_inst_lut2_199),
    .O(\DLX_IDinst_RegFile_23_21/XORG )
  );
  X_BUF \DLX_IDinst_RegFile_23_21/CYINIT_1784  (
    .I(\DLX_IDinst_RegFile_23_21/LOGIC_ONE ),
    .O(\DLX_IDinst_RegFile_23_21/CYINIT )
  );
  X_MUX2 DLX_IDinst_Msub__n0157_inst_cy_267_1785 (
    .IA(GLOBAL_LOGIC0),
    .IB(\DLX_IDinst__n0157<2>/CYINIT ),
    .SEL(\DLX_IDinst__n0157<2>/FROM ),
    .O(DLX_IDinst_Msub__n0157_inst_cy_267)
  );
  X_XOR2 DLX_IDinst_Msub__n0157_inst_sum_104 (
    .I0(\DLX_IDinst__n0157<2>/CYINIT ),
    .I1(\DLX_IDinst__n0157<2>/FROM ),
    .O(\DLX_IDinst__n0157<2>/XORF )
  );
  defparam \DLX_IDinst__n0157<2>/F .INIT = 16'hCCCC;
  X_LUT4 \DLX_IDinst__n0157<2>/F  (
    .ADR0(GLOBAL_LOGIC0),
    .ADR1(DLX_IDinst__n0158[2]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IDinst__n0157<2>/FROM )
  );
  defparam DLX_IDinst_Msub__n0157_inst_lut2_2011.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0157_inst_lut2_2011 (
    .ADR0(DLX_IDinst__n0158[3]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0157_inst_lut2_201)
  );
  X_BUF \DLX_IDinst__n0157<2>/COUTUSED  (
    .I(\DLX_IDinst__n0157<2>/CYMUXG ),
    .O(DLX_IDinst_Msub__n0157_inst_cy_268)
  );
  X_BUF \DLX_IDinst__n0157<2>/XUSED  (
    .I(\DLX_IDinst__n0157<2>/XORF ),
    .O(DLX_IDinst__n0157[2])
  );
  X_BUF \DLX_IDinst__n0157<2>/YUSED  (
    .I(\DLX_IDinst__n0157<2>/XORG ),
    .O(DLX_IDinst__n0157[3])
  );
  X_MUX2 DLX_IDinst_Msub__n0157_inst_cy_268_1786 (
    .IA(DLX_IDinst__n0158[3]),
    .IB(DLX_IDinst_Msub__n0157_inst_cy_267),
    .SEL(DLX_IDinst_Msub__n0157_inst_lut2_201),
    .O(\DLX_IDinst__n0157<2>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Msub__n0157_inst_sum_105 (
    .I0(DLX_IDinst_Msub__n0157_inst_cy_267),
    .I1(DLX_IDinst_Msub__n0157_inst_lut2_201),
    .O(\DLX_IDinst__n0157<2>/XORG )
  );
  X_BUF \DLX_IDinst__n0157<2>/CYINIT_1787  (
    .I(DLX_IDinst_Msub__n0157_inst_cy_266),
    .O(\DLX_IDinst__n0157<2>/CYINIT )
  );
  X_MUX2 DLX_IDinst_Msub__n0157_inst_cy_269_1788 (
    .IA(DLX_IDinst__n0158[4]),
    .IB(\DLX_IDinst__n0157<4>/CYINIT ),
    .SEL(DLX_IDinst_Msub__n0157_inst_lut2_202),
    .O(DLX_IDinst_Msub__n0157_inst_cy_269)
  );
  X_XOR2 DLX_IDinst_Msub__n0157_inst_sum_106 (
    .I0(\DLX_IDinst__n0157<4>/CYINIT ),
    .I1(DLX_IDinst_Msub__n0157_inst_lut2_202),
    .O(\DLX_IDinst__n0157<4>/XORF )
  );
  defparam DLX_IDinst_Msub__n0157_inst_lut2_2021.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0157_inst_lut2_2021 (
    .ADR0(DLX_IDinst__n0158[4]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0157_inst_lut2_202)
  );
  defparam DLX_IDinst_Msub__n0157_inst_lut2_2031.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0157_inst_lut2_2031 (
    .ADR0(DLX_IDinst__n0158[5]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0157_inst_lut2_203)
  );
  X_BUF \DLX_IDinst__n0157<4>/COUTUSED  (
    .I(\DLX_IDinst__n0157<4>/CYMUXG ),
    .O(DLX_IDinst_Msub__n0157_inst_cy_270)
  );
  X_BUF \DLX_IDinst__n0157<4>/XUSED  (
    .I(\DLX_IDinst__n0157<4>/XORF ),
    .O(DLX_IDinst__n0157[4])
  );
  X_BUF \DLX_IDinst__n0157<4>/YUSED  (
    .I(\DLX_IDinst__n0157<4>/XORG ),
    .O(DLX_IDinst__n0157[5])
  );
  X_MUX2 DLX_IDinst_Msub__n0157_inst_cy_270_1789 (
    .IA(DLX_IDinst__n0158[5]),
    .IB(DLX_IDinst_Msub__n0157_inst_cy_269),
    .SEL(DLX_IDinst_Msub__n0157_inst_lut2_203),
    .O(\DLX_IDinst__n0157<4>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Msub__n0157_inst_sum_107 (
    .I0(DLX_IDinst_Msub__n0157_inst_cy_269),
    .I1(DLX_IDinst_Msub__n0157_inst_lut2_203),
    .O(\DLX_IDinst__n0157<4>/XORG )
  );
  X_BUF \DLX_IDinst__n0157<4>/CYINIT_1790  (
    .I(DLX_IDinst_Msub__n0157_inst_cy_268),
    .O(\DLX_IDinst__n0157<4>/CYINIT )
  );
  X_MUX2 DLX_IDinst_Msub__n0157_inst_cy_271_1791 (
    .IA(DLX_IDinst__n0158[6]),
    .IB(\DLX_IDinst_RegFile_6_20/CYINIT ),
    .SEL(DLX_IDinst_Msub__n0157_inst_lut2_204),
    .O(DLX_IDinst_Msub__n0157_inst_cy_271)
  );
  X_XOR2 DLX_IDinst_Msub__n0157_inst_sum_108 (
    .I0(\DLX_IDinst_RegFile_6_20/CYINIT ),
    .I1(DLX_IDinst_Msub__n0157_inst_lut2_204),
    .O(\DLX_IDinst_RegFile_6_20/XORF )
  );
  defparam DLX_IDinst_Msub__n0157_inst_lut2_2041.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0157_inst_lut2_2041 (
    .ADR0(DLX_IDinst__n0158[6]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0157_inst_lut2_204)
  );
  defparam DLX_IDinst_Msub__n0157_inst_lut2_2051.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0157_inst_lut2_2051 (
    .ADR0(DLX_IDinst__n0158[7]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0157_inst_lut2_205)
  );
  X_BUF \DLX_IDinst_RegFile_6_20/COUTUSED  (
    .I(\DLX_IDinst_RegFile_6_20/CYMUXG ),
    .O(DLX_IDinst_Msub__n0157_inst_cy_272)
  );
  X_BUF \DLX_IDinst_RegFile_6_20/XUSED  (
    .I(\DLX_IDinst_RegFile_6_20/XORF ),
    .O(DLX_IDinst__n0157[6])
  );
  X_BUF \DLX_IDinst_RegFile_6_20/YUSED  (
    .I(\DLX_IDinst_RegFile_6_20/XORG ),
    .O(DLX_IDinst__n0157[7])
  );
  X_MUX2 DLX_IDinst_Msub__n0157_inst_cy_272_1792 (
    .IA(DLX_IDinst__n0158[7]),
    .IB(DLX_IDinst_Msub__n0157_inst_cy_271),
    .SEL(DLX_IDinst_Msub__n0157_inst_lut2_205),
    .O(\DLX_IDinst_RegFile_6_20/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Msub__n0157_inst_sum_109 (
    .I0(DLX_IDinst_Msub__n0157_inst_cy_271),
    .I1(DLX_IDinst_Msub__n0157_inst_lut2_205),
    .O(\DLX_IDinst_RegFile_6_20/XORG )
  );
  X_BUF \DLX_IDinst_RegFile_6_20/CYINIT_1793  (
    .I(DLX_IDinst_Msub__n0157_inst_cy_270),
    .O(\DLX_IDinst_RegFile_6_20/CYINIT )
  );
  X_MUX2 DLX_IDinst_Msub__n0157_inst_cy_273_1794 (
    .IA(DLX_IDinst__n0158[8]),
    .IB(\DLX_IDinst__n0157<8>/CYINIT ),
    .SEL(DLX_IDinst_Msub__n0157_inst_lut2_206),
    .O(DLX_IDinst_Msub__n0157_inst_cy_273)
  );
  X_XOR2 DLX_IDinst_Msub__n0157_inst_sum_110 (
    .I0(\DLX_IDinst__n0157<8>/CYINIT ),
    .I1(DLX_IDinst_Msub__n0157_inst_lut2_206),
    .O(\DLX_IDinst__n0157<8>/XORF )
  );
  defparam DLX_IDinst_Msub__n0157_inst_lut2_2061.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0157_inst_lut2_2061 (
    .ADR0(DLX_IDinst__n0158[8]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0157_inst_lut2_206)
  );
  defparam DLX_IDinst_Msub__n0157_inst_lut2_2071.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0157_inst_lut2_2071 (
    .ADR0(DLX_IDinst__n0158[9]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0157_inst_lut2_207)
  );
  X_BUF \DLX_IDinst__n0157<8>/COUTUSED  (
    .I(\DLX_IDinst__n0157<8>/CYMUXG ),
    .O(DLX_IDinst_Msub__n0157_inst_cy_274)
  );
  X_BUF \DLX_IDinst__n0157<8>/XUSED  (
    .I(\DLX_IDinst__n0157<8>/XORF ),
    .O(DLX_IDinst__n0157[8])
  );
  X_BUF \DLX_IDinst__n0157<8>/YUSED  (
    .I(\DLX_IDinst__n0157<8>/XORG ),
    .O(DLX_IDinst__n0157[9])
  );
  X_MUX2 DLX_IDinst_Msub__n0157_inst_cy_274_1795 (
    .IA(DLX_IDinst__n0158[9]),
    .IB(DLX_IDinst_Msub__n0157_inst_cy_273),
    .SEL(DLX_IDinst_Msub__n0157_inst_lut2_207),
    .O(\DLX_IDinst__n0157<8>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Msub__n0157_inst_sum_111 (
    .I0(DLX_IDinst_Msub__n0157_inst_cy_273),
    .I1(DLX_IDinst_Msub__n0157_inst_lut2_207),
    .O(\DLX_IDinst__n0157<8>/XORG )
  );
  X_BUF \DLX_IDinst__n0157<8>/CYINIT_1796  (
    .I(DLX_IDinst_Msub__n0157_inst_cy_272),
    .O(\DLX_IDinst__n0157<8>/CYINIT )
  );
  X_MUX2 DLX_IDinst_Msub__n0157_inst_cy_275_1797 (
    .IA(DLX_IDinst__n0158[10]),
    .IB(\DLX_IDinst_RegFile_15_20/CYINIT ),
    .SEL(DLX_IDinst_Msub__n0157_inst_lut2_208),
    .O(DLX_IDinst_Msub__n0157_inst_cy_275)
  );
  X_XOR2 DLX_IDinst_Msub__n0157_inst_sum_112 (
    .I0(\DLX_IDinst_RegFile_15_20/CYINIT ),
    .I1(DLX_IDinst_Msub__n0157_inst_lut2_208),
    .O(\DLX_IDinst_RegFile_15_20/XORF )
  );
  defparam DLX_IDinst_Msub__n0157_inst_lut2_2081.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0157_inst_lut2_2081 (
    .ADR0(DLX_IDinst__n0158[10]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0157_inst_lut2_208)
  );
  defparam DLX_IDinst_Msub__n0157_inst_lut2_2091.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0157_inst_lut2_2091 (
    .ADR0(DLX_IDinst__n0158[11]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0157_inst_lut2_209)
  );
  X_BUF \DLX_IDinst_RegFile_15_20/COUTUSED  (
    .I(\DLX_IDinst_RegFile_15_20/CYMUXG ),
    .O(DLX_IDinst_Msub__n0157_inst_cy_276)
  );
  X_BUF \DLX_IDinst_RegFile_15_20/XUSED  (
    .I(\DLX_IDinst_RegFile_15_20/XORF ),
    .O(DLX_IDinst__n0157[10])
  );
  X_BUF \DLX_IDinst_RegFile_15_20/YUSED  (
    .I(\DLX_IDinst_RegFile_15_20/XORG ),
    .O(DLX_IDinst__n0157[11])
  );
  X_MUX2 DLX_IDinst_Msub__n0157_inst_cy_276_1798 (
    .IA(DLX_IDinst__n0158[11]),
    .IB(DLX_IDinst_Msub__n0157_inst_cy_275),
    .SEL(DLX_IDinst_Msub__n0157_inst_lut2_209),
    .O(\DLX_IDinst_RegFile_15_20/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Msub__n0157_inst_sum_113 (
    .I0(DLX_IDinst_Msub__n0157_inst_cy_275),
    .I1(DLX_IDinst_Msub__n0157_inst_lut2_209),
    .O(\DLX_IDinst_RegFile_15_20/XORG )
  );
  X_BUF \DLX_IDinst_RegFile_15_20/CYINIT_1799  (
    .I(DLX_IDinst_Msub__n0157_inst_cy_274),
    .O(\DLX_IDinst_RegFile_15_20/CYINIT )
  );
  X_MUX2 DLX_IDinst_Msub__n0157_inst_cy_277_1800 (
    .IA(DLX_IDinst__n0158[12]),
    .IB(\DLX_IDinst__n0157<12>/CYINIT ),
    .SEL(DLX_IDinst_Msub__n0157_inst_lut2_210),
    .O(DLX_IDinst_Msub__n0157_inst_cy_277)
  );
  X_XOR2 DLX_IDinst_Msub__n0157_inst_sum_114 (
    .I0(\DLX_IDinst__n0157<12>/CYINIT ),
    .I1(DLX_IDinst_Msub__n0157_inst_lut2_210),
    .O(\DLX_IDinst__n0157<12>/XORF )
  );
  defparam DLX_IDinst_Msub__n0157_inst_lut2_2101.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0157_inst_lut2_2101 (
    .ADR0(DLX_IDinst__n0158[12]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0157_inst_lut2_210)
  );
  defparam DLX_IDinst_Msub__n0157_inst_lut2_2111.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0157_inst_lut2_2111 (
    .ADR0(DLX_IDinst__n0158[13]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0157_inst_lut2_211)
  );
  X_BUF \DLX_IDinst__n0157<12>/COUTUSED  (
    .I(\DLX_IDinst__n0157<12>/CYMUXG ),
    .O(DLX_IDinst_Msub__n0157_inst_cy_278)
  );
  X_BUF \DLX_IDinst__n0157<12>/XUSED  (
    .I(\DLX_IDinst__n0157<12>/XORF ),
    .O(DLX_IDinst__n0157[12])
  );
  X_BUF \DLX_IDinst__n0157<12>/YUSED  (
    .I(\DLX_IDinst__n0157<12>/XORG ),
    .O(DLX_IDinst__n0157[13])
  );
  X_MUX2 DLX_IDinst_Msub__n0157_inst_cy_278_1801 (
    .IA(DLX_IDinst__n0158[13]),
    .IB(DLX_IDinst_Msub__n0157_inst_cy_277),
    .SEL(DLX_IDinst_Msub__n0157_inst_lut2_211),
    .O(\DLX_IDinst__n0157<12>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Msub__n0157_inst_sum_115 (
    .I0(DLX_IDinst_Msub__n0157_inst_cy_277),
    .I1(DLX_IDinst_Msub__n0157_inst_lut2_211),
    .O(\DLX_IDinst__n0157<12>/XORG )
  );
  X_BUF \DLX_IDinst__n0157<12>/CYINIT_1802  (
    .I(DLX_IDinst_Msub__n0157_inst_cy_276),
    .O(\DLX_IDinst__n0157<12>/CYINIT )
  );
  X_MUX2 DLX_IDinst_Msub__n0157_inst_cy_279_1803 (
    .IA(DLX_IDinst__n0158[14]),
    .IB(\DLX_IDinst_RegFile_14_16/CYINIT ),
    .SEL(DLX_IDinst_Msub__n0157_inst_lut2_212),
    .O(DLX_IDinst_Msub__n0157_inst_cy_279)
  );
  X_XOR2 DLX_IDinst_Msub__n0157_inst_sum_116 (
    .I0(\DLX_IDinst_RegFile_14_16/CYINIT ),
    .I1(DLX_IDinst_Msub__n0157_inst_lut2_212),
    .O(\DLX_IDinst_RegFile_14_16/XORF )
  );
  defparam DLX_IDinst_Msub__n0157_inst_lut2_2121.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0157_inst_lut2_2121 (
    .ADR0(DLX_IDinst__n0158[14]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0157_inst_lut2_212)
  );
  defparam DLX_IDinst_Msub__n0157_inst_lut2_2131.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0157_inst_lut2_2131 (
    .ADR0(DLX_IDinst__n0158[15]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0157_inst_lut2_213)
  );
  X_BUF \DLX_IDinst_RegFile_14_16/COUTUSED  (
    .I(\DLX_IDinst_RegFile_14_16/CYMUXG ),
    .O(DLX_IDinst_Msub__n0157_inst_cy_280)
  );
  X_BUF \DLX_IDinst_RegFile_14_16/XUSED  (
    .I(\DLX_IDinst_RegFile_14_16/XORF ),
    .O(DLX_IDinst__n0157[14])
  );
  X_BUF \DLX_IDinst_RegFile_14_16/YUSED  (
    .I(\DLX_IDinst_RegFile_14_16/XORG ),
    .O(DLX_IDinst__n0157[15])
  );
  X_MUX2 DLX_IDinst_Msub__n0157_inst_cy_280_1804 (
    .IA(DLX_IDinst__n0158[15]),
    .IB(DLX_IDinst_Msub__n0157_inst_cy_279),
    .SEL(DLX_IDinst_Msub__n0157_inst_lut2_213),
    .O(\DLX_IDinst_RegFile_14_16/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Msub__n0157_inst_sum_117 (
    .I0(DLX_IDinst_Msub__n0157_inst_cy_279),
    .I1(DLX_IDinst_Msub__n0157_inst_lut2_213),
    .O(\DLX_IDinst_RegFile_14_16/XORG )
  );
  X_BUF \DLX_IDinst_RegFile_14_16/CYINIT_1805  (
    .I(DLX_IDinst_Msub__n0157_inst_cy_278),
    .O(\DLX_IDinst_RegFile_14_16/CYINIT )
  );
  X_MUX2 DLX_IDinst_Msub__n0157_inst_cy_281_1806 (
    .IA(DLX_IDinst__n0158[16]),
    .IB(\DLX_IDinst__n0157<16>/CYINIT ),
    .SEL(DLX_IDinst_Msub__n0157_inst_lut2_214),
    .O(DLX_IDinst_Msub__n0157_inst_cy_281)
  );
  X_XOR2 DLX_IDinst_Msub__n0157_inst_sum_118 (
    .I0(\DLX_IDinst__n0157<16>/CYINIT ),
    .I1(DLX_IDinst_Msub__n0157_inst_lut2_214),
    .O(\DLX_IDinst__n0157<16>/XORF )
  );
  defparam DLX_IDinst_Msub__n0157_inst_lut2_2141.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0157_inst_lut2_2141 (
    .ADR0(DLX_IDinst__n0158[16]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0157_inst_lut2_214)
  );
  defparam DLX_IDinst_Msub__n0157_inst_lut2_2151.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0157_inst_lut2_2151 (
    .ADR0(DLX_IDinst__n0158[17]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0157_inst_lut2_215)
  );
  X_BUF \DLX_IDinst__n0157<16>/COUTUSED  (
    .I(\DLX_IDinst__n0157<16>/CYMUXG ),
    .O(DLX_IDinst_Msub__n0157_inst_cy_282)
  );
  X_BUF \DLX_IDinst__n0157<16>/XUSED  (
    .I(\DLX_IDinst__n0157<16>/XORF ),
    .O(DLX_IDinst__n0157[16])
  );
  X_BUF \DLX_IDinst__n0157<16>/YUSED  (
    .I(\DLX_IDinst__n0157<16>/XORG ),
    .O(DLX_IDinst__n0157[17])
  );
  X_MUX2 DLX_IDinst_Msub__n0157_inst_cy_282_1807 (
    .IA(DLX_IDinst__n0158[17]),
    .IB(DLX_IDinst_Msub__n0157_inst_cy_281),
    .SEL(DLX_IDinst_Msub__n0157_inst_lut2_215),
    .O(\DLX_IDinst__n0157<16>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Msub__n0157_inst_sum_119 (
    .I0(DLX_IDinst_Msub__n0157_inst_cy_281),
    .I1(DLX_IDinst_Msub__n0157_inst_lut2_215),
    .O(\DLX_IDinst__n0157<16>/XORG )
  );
  X_BUF \DLX_IDinst__n0157<16>/CYINIT_1808  (
    .I(DLX_IDinst_Msub__n0157_inst_cy_280),
    .O(\DLX_IDinst__n0157<16>/CYINIT )
  );
  X_MUX2 DLX_IDinst_Msub__n0157_inst_cy_283_1809 (
    .IA(DLX_IDinst__n0158[18]),
    .IB(\DLX_IDinst_RegFile_23_12/CYINIT ),
    .SEL(DLX_IDinst_Msub__n0157_inst_lut2_216),
    .O(DLX_IDinst_Msub__n0157_inst_cy_283)
  );
  X_XOR2 DLX_IDinst_Msub__n0157_inst_sum_120 (
    .I0(\DLX_IDinst_RegFile_23_12/CYINIT ),
    .I1(DLX_IDinst_Msub__n0157_inst_lut2_216),
    .O(\DLX_IDinst_RegFile_23_12/XORF )
  );
  defparam DLX_IDinst_Msub__n0157_inst_lut2_2161.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0157_inst_lut2_2161 (
    .ADR0(DLX_IDinst__n0158[18]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0157_inst_lut2_216)
  );
  defparam DLX_IDinst_Msub__n0157_inst_lut2_2171.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0157_inst_lut2_2171 (
    .ADR0(DLX_IDinst__n0158[19]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0157_inst_lut2_217)
  );
  X_BUF \DLX_IDinst_RegFile_23_12/COUTUSED  (
    .I(\DLX_IDinst_RegFile_23_12/CYMUXG ),
    .O(DLX_IDinst_Msub__n0157_inst_cy_284)
  );
  X_BUF \DLX_IDinst_RegFile_23_12/XUSED  (
    .I(\DLX_IDinst_RegFile_23_12/XORF ),
    .O(DLX_IDinst__n0157[18])
  );
  X_BUF \DLX_IDinst_RegFile_23_12/YUSED  (
    .I(\DLX_IDinst_RegFile_23_12/XORG ),
    .O(DLX_IDinst__n0157[19])
  );
  X_MUX2 DLX_IDinst_Msub__n0157_inst_cy_284_1810 (
    .IA(DLX_IDinst__n0158[19]),
    .IB(DLX_IDinst_Msub__n0157_inst_cy_283),
    .SEL(DLX_IDinst_Msub__n0157_inst_lut2_217),
    .O(\DLX_IDinst_RegFile_23_12/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Msub__n0157_inst_sum_121 (
    .I0(DLX_IDinst_Msub__n0157_inst_cy_283),
    .I1(DLX_IDinst_Msub__n0157_inst_lut2_217),
    .O(\DLX_IDinst_RegFile_23_12/XORG )
  );
  X_BUF \DLX_IDinst_RegFile_23_12/CYINIT_1811  (
    .I(DLX_IDinst_Msub__n0157_inst_cy_282),
    .O(\DLX_IDinst_RegFile_23_12/CYINIT )
  );
  X_MUX2 DLX_IDinst_Msub__n0157_inst_cy_285_1812 (
    .IA(DLX_IDinst__n0158[20]),
    .IB(\DLX_IDinst__n0157<20>/CYINIT ),
    .SEL(DLX_IDinst_Msub__n0157_inst_lut2_218),
    .O(DLX_IDinst_Msub__n0157_inst_cy_285)
  );
  X_XOR2 DLX_IDinst_Msub__n0157_inst_sum_122 (
    .I0(\DLX_IDinst__n0157<20>/CYINIT ),
    .I1(DLX_IDinst_Msub__n0157_inst_lut2_218),
    .O(\DLX_IDinst__n0157<20>/XORF )
  );
  defparam DLX_IDinst_Msub__n0157_inst_lut2_2181.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0157_inst_lut2_2181 (
    .ADR0(DLX_IDinst__n0158[20]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0157_inst_lut2_218)
  );
  defparam DLX_IDinst_Msub__n0157_inst_lut2_2191.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0157_inst_lut2_2191 (
    .ADR0(DLX_IDinst__n0158[21]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0157_inst_lut2_219)
  );
  X_BUF \DLX_IDinst__n0157<20>/COUTUSED  (
    .I(\DLX_IDinst__n0157<20>/CYMUXG ),
    .O(DLX_IDinst_Msub__n0157_inst_cy_286)
  );
  X_BUF \DLX_IDinst__n0157<20>/XUSED  (
    .I(\DLX_IDinst__n0157<20>/XORF ),
    .O(DLX_IDinst__n0157[20])
  );
  X_BUF \DLX_IDinst__n0157<20>/YUSED  (
    .I(\DLX_IDinst__n0157<20>/XORG ),
    .O(DLX_IDinst__n0157[21])
  );
  X_MUX2 DLX_IDinst_Msub__n0157_inst_cy_286_1813 (
    .IA(DLX_IDinst__n0158[21]),
    .IB(DLX_IDinst_Msub__n0157_inst_cy_285),
    .SEL(DLX_IDinst_Msub__n0157_inst_lut2_219),
    .O(\DLX_IDinst__n0157<20>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Msub__n0157_inst_sum_123 (
    .I0(DLX_IDinst_Msub__n0157_inst_cy_285),
    .I1(DLX_IDinst_Msub__n0157_inst_lut2_219),
    .O(\DLX_IDinst__n0157<20>/XORG )
  );
  X_BUF \DLX_IDinst__n0157<20>/CYINIT_1814  (
    .I(DLX_IDinst_Msub__n0157_inst_cy_284),
    .O(\DLX_IDinst__n0157<20>/CYINIT )
  );
  defparam DLX_IDinst_RegFile_28_29_1815.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_28_29_1815 (
    .I(DLX_IDinst_WB_data_eff[29]),
    .CE(DLX_IDinst__n0606),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_28_29)
  );
  X_MUX2 DLX_IDinst_Msub__n0157_inst_cy_287_1816 (
    .IA(DLX_IDinst__n0158[22]),
    .IB(\DLX_IDinst_RegFile_6_12/CYINIT ),
    .SEL(DLX_IDinst_Msub__n0157_inst_lut2_220),
    .O(DLX_IDinst_Msub__n0157_inst_cy_287)
  );
  X_XOR2 DLX_IDinst_Msub__n0157_inst_sum_124 (
    .I0(\DLX_IDinst_RegFile_6_12/CYINIT ),
    .I1(DLX_IDinst_Msub__n0157_inst_lut2_220),
    .O(\DLX_IDinst_RegFile_6_12/XORF )
  );
  defparam DLX_IDinst_Msub__n0157_inst_lut2_2201.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0157_inst_lut2_2201 (
    .ADR0(DLX_IDinst__n0158[22]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0157_inst_lut2_220)
  );
  defparam DLX_IDinst_Msub__n0157_inst_lut2_2211.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0157_inst_lut2_2211 (
    .ADR0(DLX_IDinst__n0158[23]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0157_inst_lut2_221)
  );
  X_BUF \DLX_IDinst_RegFile_6_12/COUTUSED  (
    .I(\DLX_IDinst_RegFile_6_12/CYMUXG ),
    .O(DLX_IDinst_Msub__n0157_inst_cy_288)
  );
  X_BUF \DLX_IDinst_RegFile_6_12/XUSED  (
    .I(\DLX_IDinst_RegFile_6_12/XORF ),
    .O(DLX_IDinst__n0157[22])
  );
  X_BUF \DLX_IDinst_RegFile_6_12/YUSED  (
    .I(\DLX_IDinst_RegFile_6_12/XORG ),
    .O(DLX_IDinst__n0157[23])
  );
  X_MUX2 DLX_IDinst_Msub__n0157_inst_cy_288_1817 (
    .IA(DLX_IDinst__n0158[23]),
    .IB(DLX_IDinst_Msub__n0157_inst_cy_287),
    .SEL(DLX_IDinst_Msub__n0157_inst_lut2_221),
    .O(\DLX_IDinst_RegFile_6_12/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Msub__n0157_inst_sum_125 (
    .I0(DLX_IDinst_Msub__n0157_inst_cy_287),
    .I1(DLX_IDinst_Msub__n0157_inst_lut2_221),
    .O(\DLX_IDinst_RegFile_6_12/XORG )
  );
  X_BUF \DLX_IDinst_RegFile_6_12/CYINIT_1818  (
    .I(DLX_IDinst_Msub__n0157_inst_cy_286),
    .O(\DLX_IDinst_RegFile_6_12/CYINIT )
  );
  X_MUX2 DLX_IDinst_Msub__n0157_inst_cy_289_1819 (
    .IA(DLX_IDinst__n0158[24]),
    .IB(\DLX_IDinst__n0157<24>/CYINIT ),
    .SEL(DLX_IDinst_Msub__n0157_inst_lut2_222),
    .O(DLX_IDinst_Msub__n0157_inst_cy_289)
  );
  X_XOR2 DLX_IDinst_Msub__n0157_inst_sum_126 (
    .I0(\DLX_IDinst__n0157<24>/CYINIT ),
    .I1(DLX_IDinst_Msub__n0157_inst_lut2_222),
    .O(\DLX_IDinst__n0157<24>/XORF )
  );
  defparam DLX_IDinst_Msub__n0157_inst_lut2_2221.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0157_inst_lut2_2221 (
    .ADR0(DLX_IDinst__n0158[24]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0157_inst_lut2_222)
  );
  defparam DLX_IDinst_Msub__n0157_inst_lut2_2231.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0157_inst_lut2_2231 (
    .ADR0(DLX_IDinst__n0158[25]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0157_inst_lut2_223)
  );
  X_BUF \DLX_IDinst__n0157<24>/COUTUSED  (
    .I(\DLX_IDinst__n0157<24>/CYMUXG ),
    .O(DLX_IDinst_Msub__n0157_inst_cy_290)
  );
  X_BUF \DLX_IDinst__n0157<24>/XUSED  (
    .I(\DLX_IDinst__n0157<24>/XORF ),
    .O(DLX_IDinst__n0157[24])
  );
  X_BUF \DLX_IDinst__n0157<24>/YUSED  (
    .I(\DLX_IDinst__n0157<24>/XORG ),
    .O(DLX_IDinst__n0157[25])
  );
  X_MUX2 DLX_IDinst_Msub__n0157_inst_cy_290_1820 (
    .IA(DLX_IDinst__n0158[25]),
    .IB(DLX_IDinst_Msub__n0157_inst_cy_289),
    .SEL(DLX_IDinst_Msub__n0157_inst_lut2_223),
    .O(\DLX_IDinst__n0157<24>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Msub__n0157_inst_sum_127 (
    .I0(DLX_IDinst_Msub__n0157_inst_cy_289),
    .I1(DLX_IDinst_Msub__n0157_inst_lut2_223),
    .O(\DLX_IDinst__n0157<24>/XORG )
  );
  X_BUF \DLX_IDinst__n0157<24>/CYINIT_1821  (
    .I(DLX_IDinst_Msub__n0157_inst_cy_288),
    .O(\DLX_IDinst__n0157<24>/CYINIT )
  );
  X_MUX2 DLX_IDinst_Msub__n0157_inst_cy_291_1822 (
    .IA(DLX_IDinst__n0158[26]),
    .IB(\DLX_IDinst_RegFile_1_7/CYINIT ),
    .SEL(DLX_IDinst_Msub__n0157_inst_lut2_224),
    .O(DLX_IDinst_Msub__n0157_inst_cy_291)
  );
  X_XOR2 DLX_IDinst_Msub__n0157_inst_sum_128 (
    .I0(\DLX_IDinst_RegFile_1_7/CYINIT ),
    .I1(DLX_IDinst_Msub__n0157_inst_lut2_224),
    .O(\DLX_IDinst_RegFile_1_7/XORF )
  );
  defparam DLX_IDinst_Msub__n0157_inst_lut2_2241.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0157_inst_lut2_2241 (
    .ADR0(DLX_IDinst__n0158[26]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0157_inst_lut2_224)
  );
  defparam DLX_IDinst_Msub__n0157_inst_lut2_2251.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0157_inst_lut2_2251 (
    .ADR0(DLX_IDinst__n0158[27]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0157_inst_lut2_225)
  );
  X_BUF \DLX_IDinst_RegFile_1_7/COUTUSED  (
    .I(\DLX_IDinst_RegFile_1_7/CYMUXG ),
    .O(DLX_IDinst_Msub__n0157_inst_cy_292)
  );
  X_BUF \DLX_IDinst_RegFile_1_7/XUSED  (
    .I(\DLX_IDinst_RegFile_1_7/XORF ),
    .O(DLX_IDinst__n0157[26])
  );
  X_BUF \DLX_IDinst_RegFile_1_7/YUSED  (
    .I(\DLX_IDinst_RegFile_1_7/XORG ),
    .O(DLX_IDinst__n0157[27])
  );
  X_MUX2 DLX_IDinst_Msub__n0157_inst_cy_292_1823 (
    .IA(DLX_IDinst__n0158[27]),
    .IB(DLX_IDinst_Msub__n0157_inst_cy_291),
    .SEL(DLX_IDinst_Msub__n0157_inst_lut2_225),
    .O(\DLX_IDinst_RegFile_1_7/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Msub__n0157_inst_sum_129 (
    .I0(DLX_IDinst_Msub__n0157_inst_cy_291),
    .I1(DLX_IDinst_Msub__n0157_inst_lut2_225),
    .O(\DLX_IDinst_RegFile_1_7/XORG )
  );
  X_BUF \DLX_IDinst_RegFile_1_7/CYINIT_1824  (
    .I(DLX_IDinst_Msub__n0157_inst_cy_290),
    .O(\DLX_IDinst_RegFile_1_7/CYINIT )
  );
  X_MUX2 DLX_IDinst_Msub__n0157_inst_cy_293_1825 (
    .IA(DLX_IDinst__n0158[28]),
    .IB(\DLX_IDinst__n0157<28>/CYINIT ),
    .SEL(DLX_IDinst_Msub__n0157_inst_lut2_226),
    .O(DLX_IDinst_Msub__n0157_inst_cy_293)
  );
  X_XOR2 DLX_IDinst_Msub__n0157_inst_sum_130 (
    .I0(\DLX_IDinst__n0157<28>/CYINIT ),
    .I1(DLX_IDinst_Msub__n0157_inst_lut2_226),
    .O(\DLX_IDinst__n0157<28>/XORF )
  );
  defparam DLX_IDinst_Msub__n0157_inst_lut2_2261.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0157_inst_lut2_2261 (
    .ADR0(DLX_IDinst__n0158[28]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0157_inst_lut2_226)
  );
  defparam DLX_IDinst_Msub__n0157_inst_lut2_2271.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0157_inst_lut2_2271 (
    .ADR0(DLX_IDinst__n0158[29]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0157_inst_lut2_227)
  );
  X_BUF \DLX_IDinst__n0157<28>/COUTUSED  (
    .I(\DLX_IDinst__n0157<28>/CYMUXG ),
    .O(DLX_IDinst_Msub__n0157_inst_cy_294)
  );
  X_BUF \DLX_IDinst__n0157<28>/XUSED  (
    .I(\DLX_IDinst__n0157<28>/XORF ),
    .O(DLX_IDinst__n0157[28])
  );
  X_BUF \DLX_IDinst__n0157<28>/YUSED  (
    .I(\DLX_IDinst__n0157<28>/XORG ),
    .O(DLX_IDinst__n0157[29])
  );
  X_MUX2 DLX_IDinst_Msub__n0157_inst_cy_294_1826 (
    .IA(DLX_IDinst__n0158[29]),
    .IB(DLX_IDinst_Msub__n0157_inst_cy_293),
    .SEL(DLX_IDinst_Msub__n0157_inst_lut2_227),
    .O(\DLX_IDinst__n0157<28>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Msub__n0157_inst_sum_131 (
    .I0(DLX_IDinst_Msub__n0157_inst_cy_293),
    .I1(DLX_IDinst_Msub__n0157_inst_lut2_227),
    .O(\DLX_IDinst__n0157<28>/XORG )
  );
  X_BUF \DLX_IDinst__n0157<28>/CYINIT_1827  (
    .I(DLX_IDinst_Msub__n0157_inst_cy_292),
    .O(\DLX_IDinst__n0157<28>/CYINIT )
  );
  X_MUX2 DLX_IDinst_Msub__n0157_inst_cy_295_1828 (
    .IA(DLX_IDinst__n0158[30]),
    .IB(\DLX_IDinst_RegFile_10_9/CYINIT ),
    .SEL(DLX_IDinst_Msub__n0157_inst_lut2_228),
    .O(DLX_IDinst_Msub__n0157_inst_cy_295)
  );
  X_XOR2 DLX_IDinst_Msub__n0157_inst_sum_132 (
    .I0(\DLX_IDinst_RegFile_10_9/CYINIT ),
    .I1(DLX_IDinst_Msub__n0157_inst_lut2_228),
    .O(\DLX_IDinst_RegFile_10_9/XORF )
  );
  defparam DLX_IDinst_Msub__n0157_inst_lut2_2281.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0157_inst_lut2_2281 (
    .ADR0(DLX_IDinst__n0158[30]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0157_inst_lut2_228)
  );
  defparam DLX_IDinst_Msub__n0157_inst_lut2_2291.INIT = 16'h5555;
  X_LUT4 DLX_IDinst_Msub__n0157_inst_lut2_2291 (
    .ADR0(DLX_IDinst__n0158[31]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_IDinst_Msub__n0157_inst_lut2_229)
  );
  X_BUF \DLX_IDinst_RegFile_10_9/XUSED  (
    .I(\DLX_IDinst_RegFile_10_9/XORF ),
    .O(DLX_IDinst__n0157[30])
  );
  X_BUF \DLX_IDinst_RegFile_10_9/YUSED  (
    .I(\DLX_IDinst_RegFile_10_9/XORG ),
    .O(DLX_IDinst__n0157[31])
  );
  X_XOR2 DLX_IDinst_Msub__n0157_inst_sum_133 (
    .I0(DLX_IDinst_Msub__n0157_inst_cy_295),
    .I1(DLX_IDinst_Msub__n0157_inst_lut2_229),
    .O(\DLX_IDinst_RegFile_10_9/XORG )
  );
  X_BUF \DLX_IDinst_RegFile_10_9/CYINIT_1829  (
    .I(DLX_IDinst_Msub__n0157_inst_cy_294),
    .O(\DLX_IDinst_RegFile_10_9/CYINIT )
  );
  X_ZERO \vga_top_vga1_gridhcounter<0>/LOGIC_ZERO_1830  (
    .O(\vga_top_vga1_gridhcounter<0>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_0_1831 (
    .IA(GLOBAL_LOGIC1),
    .IB(\vga_top_vga1_gridhcounter<0>/LOGIC_ZERO ),
    .SEL(vga_top_vga1_gridhcounter_Madd__n0000_inst_lut2_0),
    .O(vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_0)
  );
  defparam vga_top_vga1_gridhcounter_Madd__n0000_inst_lut2_01.INIT = 16'h3333;
  X_LUT4 vga_top_vga1_gridhcounter_Madd__n0000_inst_lut2_01 (
    .ADR0(GLOBAL_LOGIC1),
    .ADR1(vga_top_vga1_gridhcounter[0]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(vga_top_vga1_gridhcounter_Madd__n0000_inst_lut2_0)
  );
  defparam \vga_top_vga1_gridhcounter<0>/G .INIT = 16'hFF00;
  X_LUT4 \vga_top_vga1_gridhcounter<0>/G  (
    .ADR0(GLOBAL_LOGIC0),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_gridhcounter[1]),
    .O(\vga_top_vga1_gridhcounter<0>/GROM )
  );
  X_BUF \vga_top_vga1_gridhcounter<0>/COUTUSED  (
    .I(\vga_top_vga1_gridhcounter<0>/CYMUXG ),
    .O(vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_1)
  );
  X_MUX2 vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_1_1832 (
    .IA(GLOBAL_LOGIC0),
    .IB(vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_0),
    .SEL(\vga_top_vga1_gridhcounter<0>/GROM ),
    .O(\vga_top_vga1_gridhcounter<0>/CYMUXG )
  );
  X_XOR2 vga_top_vga1_gridhcounter_Madd__n0000_inst_sum_1 (
    .I0(vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_0),
    .I1(\vga_top_vga1_gridhcounter<0>/GROM ),
    .O(vga_top_vga1_gridhcounter__n0000[1])
  );
  X_ZERO \vga_top_vga1_gridhcounter<2>/LOGIC_ZERO_1833  (
    .O(\vga_top_vga1_gridhcounter<2>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_2_1834 (
    .IA(\vga_top_vga1_gridhcounter<2>/LOGIC_ZERO ),
    .IB(\vga_top_vga1_gridhcounter<2>/CYINIT ),
    .SEL(\vga_top_vga1_gridhcounter<2>/FROM ),
    .O(vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_2)
  );
  X_XOR2 vga_top_vga1_gridhcounter_Madd__n0000_inst_sum_2 (
    .I0(\vga_top_vga1_gridhcounter<2>/CYINIT ),
    .I1(\vga_top_vga1_gridhcounter<2>/FROM ),
    .O(vga_top_vga1_gridhcounter__n0000[2])
  );
  defparam \vga_top_vga1_gridhcounter<2>/F .INIT = 16'hCCCC;
  X_LUT4 \vga_top_vga1_gridhcounter<2>/F  (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_gridhcounter[2]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\vga_top_vga1_gridhcounter<2>/FROM )
  );
  defparam \vga_top_vga1_gridhcounter<2>/G .INIT = 16'hF0F0;
  X_LUT4 \vga_top_vga1_gridhcounter<2>/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_gridhcounter[3]),
    .ADR3(VCC),
    .O(\vga_top_vga1_gridhcounter<2>/GROM )
  );
  X_BUF \vga_top_vga1_gridhcounter<2>/COUTUSED  (
    .I(\vga_top_vga1_gridhcounter<2>/CYMUXG ),
    .O(vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_3)
  );
  X_MUX2 vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_3_1835 (
    .IA(\vga_top_vga1_gridhcounter<2>/LOGIC_ZERO ),
    .IB(vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_2),
    .SEL(\vga_top_vga1_gridhcounter<2>/GROM ),
    .O(\vga_top_vga1_gridhcounter<2>/CYMUXG )
  );
  X_XOR2 vga_top_vga1_gridhcounter_Madd__n0000_inst_sum_3 (
    .I0(vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_2),
    .I1(\vga_top_vga1_gridhcounter<2>/GROM ),
    .O(vga_top_vga1_gridhcounter__n0000[3])
  );
  X_BUF \vga_top_vga1_gridhcounter<2>/CYINIT_1836  (
    .I(vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_1),
    .O(\vga_top_vga1_gridhcounter<2>/CYINIT )
  );
  X_ZERO \vga_top_vga1_gridhcounter<4>/LOGIC_ZERO_1837  (
    .O(\vga_top_vga1_gridhcounter<4>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_4_1838 (
    .IA(\vga_top_vga1_gridhcounter<4>/LOGIC_ZERO ),
    .IB(\vga_top_vga1_gridhcounter<4>/CYINIT ),
    .SEL(\vga_top_vga1_gridhcounter<4>/FROM ),
    .O(vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_4)
  );
  X_XOR2 vga_top_vga1_gridhcounter_Madd__n0000_inst_sum_4 (
    .I0(\vga_top_vga1_gridhcounter<4>/CYINIT ),
    .I1(\vga_top_vga1_gridhcounter<4>/FROM ),
    .O(vga_top_vga1_gridhcounter__n0000[4])
  );
  defparam \vga_top_vga1_gridhcounter<4>/F .INIT = 16'hCCCC;
  X_LUT4 \vga_top_vga1_gridhcounter<4>/F  (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_gridhcounter[4]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\vga_top_vga1_gridhcounter<4>/FROM )
  );
  defparam \vga_top_vga1_gridhcounter<4>/G .INIT = 16'hF0F0;
  X_LUT4 \vga_top_vga1_gridhcounter<4>/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_gridhcounter[5]),
    .ADR3(VCC),
    .O(\vga_top_vga1_gridhcounter<4>/GROM )
  );
  X_BUF \vga_top_vga1_gridhcounter<4>/COUTUSED  (
    .I(\vga_top_vga1_gridhcounter<4>/CYMUXG ),
    .O(vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_5)
  );
  X_MUX2 vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_5_1839 (
    .IA(\vga_top_vga1_gridhcounter<4>/LOGIC_ZERO ),
    .IB(vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_4),
    .SEL(\vga_top_vga1_gridhcounter<4>/GROM ),
    .O(\vga_top_vga1_gridhcounter<4>/CYMUXG )
  );
  X_XOR2 vga_top_vga1_gridhcounter_Madd__n0000_inst_sum_5 (
    .I0(vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_4),
    .I1(\vga_top_vga1_gridhcounter<4>/GROM ),
    .O(vga_top_vga1_gridhcounter__n0000[5])
  );
  X_BUF \vga_top_vga1_gridhcounter<4>/CYINIT_1840  (
    .I(vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_3),
    .O(\vga_top_vga1_gridhcounter<4>/CYINIT )
  );
  X_ZERO \vga_top_vga1_gridhcounter<6>/LOGIC_ZERO_1841  (
    .O(\vga_top_vga1_gridhcounter<6>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_6_1842 (
    .IA(\vga_top_vga1_gridhcounter<6>/LOGIC_ZERO ),
    .IB(\vga_top_vga1_gridhcounter<6>/CYINIT ),
    .SEL(\vga_top_vga1_gridhcounter<6>/FROM ),
    .O(vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_6)
  );
  X_XOR2 vga_top_vga1_gridhcounter_Madd__n0000_inst_sum_6 (
    .I0(\vga_top_vga1_gridhcounter<6>/CYINIT ),
    .I1(\vga_top_vga1_gridhcounter<6>/FROM ),
    .O(vga_top_vga1_gridhcounter__n0000[6])
  );
  defparam \vga_top_vga1_gridhcounter<6>/F .INIT = 16'hCCCC;
  X_LUT4 \vga_top_vga1_gridhcounter<6>/F  (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_gridhcounter[6]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\vga_top_vga1_gridhcounter<6>/FROM )
  );
  defparam \vga_top_vga1_gridhcounter<6>/G .INIT = 16'hF0F0;
  X_LUT4 \vga_top_vga1_gridhcounter<6>/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_gridhcounter[7]),
    .ADR3(VCC),
    .O(\vga_top_vga1_gridhcounter<6>/GROM )
  );
  X_BUF \vga_top_vga1_gridhcounter<6>/COUTUSED  (
    .I(\vga_top_vga1_gridhcounter<6>/CYMUXG ),
    .O(vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_7)
  );
  X_MUX2 vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_7_1843 (
    .IA(\vga_top_vga1_gridhcounter<6>/LOGIC_ZERO ),
    .IB(vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_6),
    .SEL(\vga_top_vga1_gridhcounter<6>/GROM ),
    .O(\vga_top_vga1_gridhcounter<6>/CYMUXG )
  );
  X_XOR2 vga_top_vga1_gridhcounter_Madd__n0000_inst_sum_7 (
    .I0(vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_6),
    .I1(\vga_top_vga1_gridhcounter<6>/GROM ),
    .O(vga_top_vga1_gridhcounter__n0000[7])
  );
  X_BUF \vga_top_vga1_gridhcounter<6>/CYINIT_1844  (
    .I(vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_5),
    .O(\vga_top_vga1_gridhcounter<6>/CYINIT )
  );
  X_XOR2 vga_top_vga1_gridhcounter_Madd__n0000_inst_sum_8 (
    .I0(\vga_top_vga1_gridhcounter<8>/CYINIT ),
    .I1(\vga_top_vga1_gridhcounter<8>_rt ),
    .O(vga_top_vga1_gridhcounter__n0000[8])
  );
  defparam \vga_top_vga1_gridhcounter<8>_rt_1845 .INIT = 16'hCCCC;
  X_LUT4 \vga_top_vga1_gridhcounter<8>_rt_1845  (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_gridhcounter[8]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\vga_top_vga1_gridhcounter<8>_rt )
  );
  X_BUF \vga_top_vga1_gridhcounter<8>/CYINIT_1846  (
    .I(vga_top_vga1_gridhcounter_Madd__n0000_inst_cy_7),
    .O(\vga_top_vga1_gridhcounter<8>/CYINIT )
  );
  X_ZERO \vga_top_vga1_hcounter<0>/LOGIC_ZERO_1847  (
    .O(\vga_top_vga1_hcounter<0>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_hcounter_Madd__n0000_inst_cy_19_1848 (
    .IA(GLOBAL_LOGIC1),
    .IB(\vga_top_vga1_hcounter<0>/LOGIC_ZERO ),
    .SEL(vga_top_vga1_hcounter_Madd__n0000_inst_lut2_19),
    .O(vga_top_vga1_hcounter_Madd__n0000_inst_cy_19)
  );
  defparam vga_top_vga1_hcounter_Madd__n0000_inst_lut2_191.INIT = 16'h3333;
  X_LUT4 vga_top_vga1_hcounter_Madd__n0000_inst_lut2_191 (
    .ADR0(GLOBAL_LOGIC1),
    .ADR1(vga_top_vga1_hcounter[0]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(vga_top_vga1_hcounter_Madd__n0000_inst_lut2_19)
  );
  defparam \vga_top_vga1_hcounter<0>/G .INIT = 16'hF0F0;
  X_LUT4 \vga_top_vga1_hcounter<0>/G  (
    .ADR0(GLOBAL_LOGIC0),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_hcounter[1]),
    .ADR3(VCC),
    .O(\vga_top_vga1_hcounter<0>/GROM )
  );
  X_BUF \vga_top_vga1_hcounter<0>/COUTUSED  (
    .I(\vga_top_vga1_hcounter<0>/CYMUXG ),
    .O(vga_top_vga1_hcounter_Madd__n0000_inst_cy_20)
  );
  X_MUX2 vga_top_vga1_hcounter_Madd__n0000_inst_cy_20_1849 (
    .IA(GLOBAL_LOGIC0),
    .IB(vga_top_vga1_hcounter_Madd__n0000_inst_cy_19),
    .SEL(\vga_top_vga1_hcounter<0>/GROM ),
    .O(\vga_top_vga1_hcounter<0>/CYMUXG )
  );
  X_XOR2 vga_top_vga1_hcounter_Madd__n0000_inst_sum_20 (
    .I0(vga_top_vga1_hcounter_Madd__n0000_inst_cy_19),
    .I1(\vga_top_vga1_hcounter<0>/GROM ),
    .O(vga_top_vga1_hcounter__n0000[1])
  );
  X_ZERO \vga_top_vga1_hcounter<2>/LOGIC_ZERO_1850  (
    .O(\vga_top_vga1_hcounter<2>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_hcounter_Madd__n0000_inst_cy_21_1851 (
    .IA(\vga_top_vga1_hcounter<2>/LOGIC_ZERO ),
    .IB(\vga_top_vga1_hcounter<2>/CYINIT ),
    .SEL(\vga_top_vga1_hcounter<2>/FROM ),
    .O(vga_top_vga1_hcounter_Madd__n0000_inst_cy_21)
  );
  X_XOR2 vga_top_vga1_hcounter_Madd__n0000_inst_sum_21 (
    .I0(\vga_top_vga1_hcounter<2>/CYINIT ),
    .I1(\vga_top_vga1_hcounter<2>/FROM ),
    .O(vga_top_vga1_hcounter__n0000[2])
  );
  defparam \vga_top_vga1_hcounter<2>/F .INIT = 16'hFF00;
  X_LUT4 \vga_top_vga1_hcounter<2>/F  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[2]),
    .O(\vga_top_vga1_hcounter<2>/FROM )
  );
  defparam \vga_top_vga1_hcounter<2>/G .INIT = 16'hF0F0;
  X_LUT4 \vga_top_vga1_hcounter<2>/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_hcounter[3]),
    .ADR3(VCC),
    .O(\vga_top_vga1_hcounter<2>/GROM )
  );
  X_BUF \vga_top_vga1_hcounter<2>/COUTUSED  (
    .I(\vga_top_vga1_hcounter<2>/CYMUXG ),
    .O(vga_top_vga1_hcounter_Madd__n0000_inst_cy_22)
  );
  X_MUX2 vga_top_vga1_hcounter_Madd__n0000_inst_cy_22_1852 (
    .IA(\vga_top_vga1_hcounter<2>/LOGIC_ZERO ),
    .IB(vga_top_vga1_hcounter_Madd__n0000_inst_cy_21),
    .SEL(\vga_top_vga1_hcounter<2>/GROM ),
    .O(\vga_top_vga1_hcounter<2>/CYMUXG )
  );
  X_XOR2 vga_top_vga1_hcounter_Madd__n0000_inst_sum_22 (
    .I0(vga_top_vga1_hcounter_Madd__n0000_inst_cy_21),
    .I1(\vga_top_vga1_hcounter<2>/GROM ),
    .O(vga_top_vga1_hcounter__n0000[3])
  );
  X_BUF \vga_top_vga1_hcounter<2>/CYINIT_1853  (
    .I(vga_top_vga1_hcounter_Madd__n0000_inst_cy_20),
    .O(\vga_top_vga1_hcounter<2>/CYINIT )
  );
  defparam DLX_IDinst_RegFile_29_13_1854.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_29_13_1854 (
    .I(DLX_IDinst_WB_data_eff[13]),
    .CE(DLX_IDinst__n0608),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_29_13)
  );
  X_ZERO \vga_top_vga1_hcounter<4>/LOGIC_ZERO_1855  (
    .O(\vga_top_vga1_hcounter<4>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_hcounter_Madd__n0000_inst_cy_23_1856 (
    .IA(\vga_top_vga1_hcounter<4>/LOGIC_ZERO ),
    .IB(\vga_top_vga1_hcounter<4>/CYINIT ),
    .SEL(\vga_top_vga1_hcounter<4>/FROM ),
    .O(vga_top_vga1_hcounter_Madd__n0000_inst_cy_23)
  );
  X_XOR2 vga_top_vga1_hcounter_Madd__n0000_inst_sum_23 (
    .I0(\vga_top_vga1_hcounter<4>/CYINIT ),
    .I1(\vga_top_vga1_hcounter<4>/FROM ),
    .O(vga_top_vga1_hcounter__n0000[4])
  );
  defparam \vga_top_vga1_hcounter<4>/F .INIT = 16'hFF00;
  X_LUT4 \vga_top_vga1_hcounter<4>/F  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[4]),
    .O(\vga_top_vga1_hcounter<4>/FROM )
  );
  defparam \vga_top_vga1_hcounter<4>/G .INIT = 16'hF0F0;
  X_LUT4 \vga_top_vga1_hcounter<4>/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_hcounter[5]),
    .ADR3(VCC),
    .O(\vga_top_vga1_hcounter<4>/GROM )
  );
  X_BUF \vga_top_vga1_hcounter<4>/COUTUSED  (
    .I(\vga_top_vga1_hcounter<4>/CYMUXG ),
    .O(vga_top_vga1_hcounter_Madd__n0000_inst_cy_24)
  );
  X_MUX2 vga_top_vga1_hcounter_Madd__n0000_inst_cy_24_1857 (
    .IA(\vga_top_vga1_hcounter<4>/LOGIC_ZERO ),
    .IB(vga_top_vga1_hcounter_Madd__n0000_inst_cy_23),
    .SEL(\vga_top_vga1_hcounter<4>/GROM ),
    .O(\vga_top_vga1_hcounter<4>/CYMUXG )
  );
  X_XOR2 vga_top_vga1_hcounter_Madd__n0000_inst_sum_24 (
    .I0(vga_top_vga1_hcounter_Madd__n0000_inst_cy_23),
    .I1(\vga_top_vga1_hcounter<4>/GROM ),
    .O(vga_top_vga1_hcounter__n0000[5])
  );
  X_BUF \vga_top_vga1_hcounter<4>/CYINIT_1858  (
    .I(vga_top_vga1_hcounter_Madd__n0000_inst_cy_22),
    .O(\vga_top_vga1_hcounter<4>/CYINIT )
  );
  X_ZERO \vga_top_vga1_hcounter<6>/LOGIC_ZERO_1859  (
    .O(\vga_top_vga1_hcounter<6>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_hcounter_Madd__n0000_inst_cy_25_1860 (
    .IA(\vga_top_vga1_hcounter<6>/LOGIC_ZERO ),
    .IB(\vga_top_vga1_hcounter<6>/CYINIT ),
    .SEL(\vga_top_vga1_hcounter<6>/FROM ),
    .O(vga_top_vga1_hcounter_Madd__n0000_inst_cy_25)
  );
  X_XOR2 vga_top_vga1_hcounter_Madd__n0000_inst_sum_25 (
    .I0(\vga_top_vga1_hcounter<6>/CYINIT ),
    .I1(\vga_top_vga1_hcounter<6>/FROM ),
    .O(vga_top_vga1_hcounter__n0000[6])
  );
  defparam \vga_top_vga1_hcounter<6>/F .INIT = 16'hCCCC;
  X_LUT4 \vga_top_vga1_hcounter<6>/F  (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_hcounter[6]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\vga_top_vga1_hcounter<6>/FROM )
  );
  defparam \vga_top_vga1_hcounter<6>/G .INIT = 16'hF0F0;
  X_LUT4 \vga_top_vga1_hcounter<6>/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_hcounter[7]),
    .ADR3(VCC),
    .O(\vga_top_vga1_hcounter<6>/GROM )
  );
  X_BUF \vga_top_vga1_hcounter<6>/COUTUSED  (
    .I(\vga_top_vga1_hcounter<6>/CYMUXG ),
    .O(vga_top_vga1_hcounter_Madd__n0000_inst_cy_26)
  );
  X_MUX2 vga_top_vga1_hcounter_Madd__n0000_inst_cy_26_1861 (
    .IA(\vga_top_vga1_hcounter<6>/LOGIC_ZERO ),
    .IB(vga_top_vga1_hcounter_Madd__n0000_inst_cy_25),
    .SEL(\vga_top_vga1_hcounter<6>/GROM ),
    .O(\vga_top_vga1_hcounter<6>/CYMUXG )
  );
  X_XOR2 vga_top_vga1_hcounter_Madd__n0000_inst_sum_26 (
    .I0(vga_top_vga1_hcounter_Madd__n0000_inst_cy_25),
    .I1(\vga_top_vga1_hcounter<6>/GROM ),
    .O(vga_top_vga1_hcounter__n0000[7])
  );
  X_BUF \vga_top_vga1_hcounter<6>/CYINIT_1862  (
    .I(vga_top_vga1_hcounter_Madd__n0000_inst_cy_24),
    .O(\vga_top_vga1_hcounter<6>/CYINIT )
  );
  X_ZERO \vga_top_vga1_hcounter<8>/LOGIC_ZERO_1863  (
    .O(\vga_top_vga1_hcounter<8>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_hcounter_Madd__n0000_inst_cy_27_1864 (
    .IA(\vga_top_vga1_hcounter<8>/LOGIC_ZERO ),
    .IB(\vga_top_vga1_hcounter<8>/CYINIT ),
    .SEL(\vga_top_vga1_hcounter<8>/FROM ),
    .O(vga_top_vga1_hcounter_Madd__n0000_inst_cy_27)
  );
  X_XOR2 vga_top_vga1_hcounter_Madd__n0000_inst_sum_27 (
    .I0(\vga_top_vga1_hcounter<8>/CYINIT ),
    .I1(\vga_top_vga1_hcounter<8>/FROM ),
    .O(vga_top_vga1_hcounter__n0000[8])
  );
  defparam \vga_top_vga1_hcounter<8>/F .INIT = 16'hCCCC;
  X_LUT4 \vga_top_vga1_hcounter<8>/F  (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_hcounter[8]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\vga_top_vga1_hcounter<8>/FROM )
  );
  defparam \vga_top_vga1_hcounter<8>/G .INIT = 16'hFF00;
  X_LUT4 \vga_top_vga1_hcounter<8>/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[9]),
    .O(\vga_top_vga1_hcounter<8>/GROM )
  );
  X_BUF \vga_top_vga1_hcounter<8>/COUTUSED  (
    .I(\vga_top_vga1_hcounter<8>/CYMUXG ),
    .O(vga_top_vga1_hcounter_Madd__n0000_inst_cy_28)
  );
  X_MUX2 vga_top_vga1_hcounter_Madd__n0000_inst_cy_28_1865 (
    .IA(\vga_top_vga1_hcounter<8>/LOGIC_ZERO ),
    .IB(vga_top_vga1_hcounter_Madd__n0000_inst_cy_27),
    .SEL(\vga_top_vga1_hcounter<8>/GROM ),
    .O(\vga_top_vga1_hcounter<8>/CYMUXG )
  );
  X_XOR2 vga_top_vga1_hcounter_Madd__n0000_inst_sum_28 (
    .I0(vga_top_vga1_hcounter_Madd__n0000_inst_cy_27),
    .I1(\vga_top_vga1_hcounter<8>/GROM ),
    .O(vga_top_vga1_hcounter__n0000[9])
  );
  X_BUF \vga_top_vga1_hcounter<8>/CYINIT_1866  (
    .I(vga_top_vga1_hcounter_Madd__n0000_inst_cy_26),
    .O(\vga_top_vga1_hcounter<8>/CYINIT )
  );
  X_ZERO \vga_top_vga1_hcounter<10>/LOGIC_ZERO_1867  (
    .O(\vga_top_vga1_hcounter<10>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_hcounter_Madd__n0000_inst_cy_29_1868 (
    .IA(\vga_top_vga1_hcounter<10>/LOGIC_ZERO ),
    .IB(\vga_top_vga1_hcounter<10>/CYINIT ),
    .SEL(\vga_top_vga1_hcounter<10>/FROM ),
    .O(vga_top_vga1_hcounter_Madd__n0000_inst_cy_29)
  );
  X_XOR2 vga_top_vga1_hcounter_Madd__n0000_inst_sum_29 (
    .I0(\vga_top_vga1_hcounter<10>/CYINIT ),
    .I1(\vga_top_vga1_hcounter<10>/FROM ),
    .O(vga_top_vga1_hcounter__n0000[10])
  );
  defparam \vga_top_vga1_hcounter<10>/F .INIT = 16'hCCCC;
  X_LUT4 \vga_top_vga1_hcounter<10>/F  (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_hcounter[10]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\vga_top_vga1_hcounter<10>/FROM )
  );
  defparam \vga_top_vga1_hcounter<10>/G .INIT = 16'hF0F0;
  X_LUT4 \vga_top_vga1_hcounter<10>/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_hcounter[11]),
    .ADR3(VCC),
    .O(\vga_top_vga1_hcounter<10>/GROM )
  );
  X_BUF \vga_top_vga1_hcounter<10>/COUTUSED  (
    .I(\vga_top_vga1_hcounter<10>/CYMUXG ),
    .O(vga_top_vga1_hcounter_Madd__n0000_inst_cy_30)
  );
  X_MUX2 vga_top_vga1_hcounter_Madd__n0000_inst_cy_30_1869 (
    .IA(\vga_top_vga1_hcounter<10>/LOGIC_ZERO ),
    .IB(vga_top_vga1_hcounter_Madd__n0000_inst_cy_29),
    .SEL(\vga_top_vga1_hcounter<10>/GROM ),
    .O(\vga_top_vga1_hcounter<10>/CYMUXG )
  );
  X_XOR2 vga_top_vga1_hcounter_Madd__n0000_inst_sum_30 (
    .I0(vga_top_vga1_hcounter_Madd__n0000_inst_cy_29),
    .I1(\vga_top_vga1_hcounter<10>/GROM ),
    .O(vga_top_vga1_hcounter__n0000[11])
  );
  X_BUF \vga_top_vga1_hcounter<10>/CYINIT_1870  (
    .I(vga_top_vga1_hcounter_Madd__n0000_inst_cy_28),
    .O(\vga_top_vga1_hcounter<10>/CYINIT )
  );
  X_ZERO \vga_top_vga1_hcounter<12>/LOGIC_ZERO_1871  (
    .O(\vga_top_vga1_hcounter<12>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_hcounter_Madd__n0000_inst_cy_31_1872 (
    .IA(\vga_top_vga1_hcounter<12>/LOGIC_ZERO ),
    .IB(\vga_top_vga1_hcounter<12>/CYINIT ),
    .SEL(\vga_top_vga1_hcounter<12>/FROM ),
    .O(vga_top_vga1_hcounter_Madd__n0000_inst_cy_31)
  );
  X_XOR2 vga_top_vga1_hcounter_Madd__n0000_inst_sum_31 (
    .I0(\vga_top_vga1_hcounter<12>/CYINIT ),
    .I1(\vga_top_vga1_hcounter<12>/FROM ),
    .O(vga_top_vga1_hcounter__n0000[12])
  );
  defparam \vga_top_vga1_hcounter<12>/F .INIT = 16'hCCCC;
  X_LUT4 \vga_top_vga1_hcounter<12>/F  (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_hcounter[12]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\vga_top_vga1_hcounter<12>/FROM )
  );
  defparam \vga_top_vga1_hcounter<12>/G .INIT = 16'hF0F0;
  X_LUT4 \vga_top_vga1_hcounter<12>/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_hcounter[13]),
    .ADR3(VCC),
    .O(\vga_top_vga1_hcounter<12>/GROM )
  );
  X_BUF \vga_top_vga1_hcounter<12>/COUTUSED  (
    .I(\vga_top_vga1_hcounter<12>/CYMUXG ),
    .O(vga_top_vga1_hcounter_Madd__n0000_inst_cy_32)
  );
  X_MUX2 vga_top_vga1_hcounter_Madd__n0000_inst_cy_32_1873 (
    .IA(\vga_top_vga1_hcounter<12>/LOGIC_ZERO ),
    .IB(vga_top_vga1_hcounter_Madd__n0000_inst_cy_31),
    .SEL(\vga_top_vga1_hcounter<12>/GROM ),
    .O(\vga_top_vga1_hcounter<12>/CYMUXG )
  );
  X_XOR2 vga_top_vga1_hcounter_Madd__n0000_inst_sum_32 (
    .I0(vga_top_vga1_hcounter_Madd__n0000_inst_cy_31),
    .I1(\vga_top_vga1_hcounter<12>/GROM ),
    .O(vga_top_vga1_hcounter__n0000[13])
  );
  X_BUF \vga_top_vga1_hcounter<12>/CYINIT_1874  (
    .I(vga_top_vga1_hcounter_Madd__n0000_inst_cy_30),
    .O(\vga_top_vga1_hcounter<12>/CYINIT )
  );
  X_ZERO \vga_top_vga1_hcounter<14>/LOGIC_ZERO_1875  (
    .O(\vga_top_vga1_hcounter<14>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_hcounter_Madd__n0000_inst_cy_33_1876 (
    .IA(\vga_top_vga1_hcounter<14>/LOGIC_ZERO ),
    .IB(\vga_top_vga1_hcounter<14>/CYINIT ),
    .SEL(\vga_top_vga1_hcounter<14>/FROM ),
    .O(vga_top_vga1_hcounter_Madd__n0000_inst_cy_33)
  );
  X_XOR2 vga_top_vga1_hcounter_Madd__n0000_inst_sum_33 (
    .I0(\vga_top_vga1_hcounter<14>/CYINIT ),
    .I1(\vga_top_vga1_hcounter<14>/FROM ),
    .O(vga_top_vga1_hcounter__n0000[14])
  );
  defparam \vga_top_vga1_hcounter<14>/F .INIT = 16'hF0F0;
  X_LUT4 \vga_top_vga1_hcounter<14>/F  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_hcounter[14]),
    .ADR3(VCC),
    .O(\vga_top_vga1_hcounter<14>/FROM )
  );
  defparam \vga_top_vga1_hcounter<15>_rt_1877 .INIT = 16'hAAAA;
  X_LUT4 \vga_top_vga1_hcounter<15>_rt_1877  (
    .ADR0(vga_top_vga1_hcounter[15]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\vga_top_vga1_hcounter<15>_rt )
  );
  X_XOR2 vga_top_vga1_hcounter_Madd__n0000_inst_sum_34 (
    .I0(vga_top_vga1_hcounter_Madd__n0000_inst_cy_33),
    .I1(\vga_top_vga1_hcounter<15>_rt ),
    .O(vga_top_vga1_hcounter__n0000[15])
  );
  X_BUF \vga_top_vga1_hcounter<14>/CYINIT_1878  (
    .I(vga_top_vga1_hcounter_Madd__n0000_inst_cy_32),
    .O(\vga_top_vga1_hcounter<14>/CYINIT )
  );
  X_ZERO \vga_top_vga1_Mmult__n0043_inst_lut2_317/LOGIC_ZERO_1879  (
    .O(\vga_top_vga1_Mmult__n0043_inst_lut2_317/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_Mmult__n0043_inst_cy_436_1880 (
    .IA(vga_top_vga1_gridvcounter[2]),
    .IB(\vga_top_vga1_Mmult__n0043_inst_lut2_317/LOGIC_ZERO ),
    .SEL(vga_top_vga1_Mmult__n0043_inst_lut2_303),
    .O(vga_top_vga1_Mmult__n0043_inst_cy_436)
  );
  defparam vga_top_vga1_Mmult__n0043_inst_lut2_3031.INIT = 16'h55AA;
  X_LUT4 vga_top_vga1_Mmult__n0043_inst_lut2_3031 (
    .ADR0(vga_top_vga1_gridvcounter[2]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_gridvcounter[0]),
    .O(vga_top_vga1_Mmult__n0043_inst_lut2_303)
  );
  defparam vga_top_vga1_Mmult__n0043_inst_lut2_3041.INIT = 16'h55AA;
  X_LUT4 vga_top_vga1_Mmult__n0043_inst_lut2_3041 (
    .ADR0(vga_top_vga1_gridvcounter[3]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_gridvcounter[1]),
    .O(vga_top_vga1_Mmult__n0043_inst_lut2_304)
  );
  X_BUF \vga_top_vga1_Mmult__n0043_inst_lut2_317/COUTUSED  (
    .I(\vga_top_vga1_Mmult__n0043_inst_lut2_317/CYMUXG ),
    .O(vga_top_vga1_Mmult__n0043_inst_cy_437)
  );
  X_BUF \vga_top_vga1_Mmult__n0043_inst_lut2_317/YUSED  (
    .I(\vga_top_vga1_Mmult__n0043_inst_lut2_317/XORG ),
    .O(vga_top_vga1_Mmult__n0043_inst_lut2_317)
  );
  X_MUX2 vga_top_vga1_Mmult__n0043_inst_cy_437_1881 (
    .IA(vga_top_vga1_gridvcounter[3]),
    .IB(vga_top_vga1_Mmult__n0043_inst_cy_436),
    .SEL(vga_top_vga1_Mmult__n0043_inst_lut2_304),
    .O(\vga_top_vga1_Mmult__n0043_inst_lut2_317/CYMUXG )
  );
  X_XOR2 vga_top_vga1_Mmult__n0043_inst_sum_226 (
    .I0(vga_top_vga1_Mmult__n0043_inst_cy_436),
    .I1(vga_top_vga1_Mmult__n0043_inst_lut2_304),
    .O(\vga_top_vga1_Mmult__n0043_inst_lut2_317/XORG )
  );
  X_MUX2 vga_top_vga1_Mmult__n0043_inst_cy_438_1882 (
    .IA(vga_top_vga1_gridvcounter[4]),
    .IB(\DLX_IDinst_RegFile_3_14/CYINIT ),
    .SEL(vga_top_vga1_Mmult__n0043_inst_lut2_305),
    .O(vga_top_vga1_Mmult__n0043_inst_cy_438)
  );
  X_XOR2 vga_top_vga1_Mmult__n0043_inst_sum_227 (
    .I0(\DLX_IDinst_RegFile_3_14/CYINIT ),
    .I1(vga_top_vga1_Mmult__n0043_inst_lut2_305),
    .O(\DLX_IDinst_RegFile_3_14/XORF )
  );
  defparam vga_top_vga1_Mmult__n0043_inst_lut2_3051.INIT = 16'h6666;
  X_LUT4 vga_top_vga1_Mmult__n0043_inst_lut2_3051 (
    .ADR0(vga_top_vga1_gridvcounter[4]),
    .ADR1(vga_top_vga1_gridvcounter[2]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(vga_top_vga1_Mmult__n0043_inst_lut2_305)
  );
  defparam vga_top_vga1_Mmult__n0043_inst_lut2_3061.INIT = 16'h5A5A;
  X_LUT4 vga_top_vga1_Mmult__n0043_inst_lut2_3061 (
    .ADR0(vga_top_vga1_gridvcounter[5]),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_gridvcounter[3]),
    .ADR3(VCC),
    .O(vga_top_vga1_Mmult__n0043_inst_lut2_306)
  );
  X_BUF \DLX_IDinst_RegFile_3_14/COUTUSED  (
    .I(\DLX_IDinst_RegFile_3_14/CYMUXG ),
    .O(vga_top_vga1_Mmult__n0043_inst_cy_439)
  );
  X_BUF \DLX_IDinst_RegFile_3_14/XUSED  (
    .I(\DLX_IDinst_RegFile_3_14/XORF ),
    .O(vga_top_vga1_Mmult__n0043_inst_lut2_318)
  );
  X_BUF \DLX_IDinst_RegFile_3_14/YUSED  (
    .I(\DLX_IDinst_RegFile_3_14/XORG ),
    .O(vga_top_vga1_Mmult__n0043_inst_lut2_319)
  );
  X_MUX2 vga_top_vga1_Mmult__n0043_inst_cy_439_1883 (
    .IA(vga_top_vga1_gridvcounter[5]),
    .IB(vga_top_vga1_Mmult__n0043_inst_cy_438),
    .SEL(vga_top_vga1_Mmult__n0043_inst_lut2_306),
    .O(\DLX_IDinst_RegFile_3_14/CYMUXG )
  );
  X_XOR2 vga_top_vga1_Mmult__n0043_inst_sum_228 (
    .I0(vga_top_vga1_Mmult__n0043_inst_cy_438),
    .I1(vga_top_vga1_Mmult__n0043_inst_lut2_306),
    .O(\DLX_IDinst_RegFile_3_14/XORG )
  );
  X_BUF \DLX_IDinst_RegFile_3_14/CYINIT_1884  (
    .I(vga_top_vga1_Mmult__n0043_inst_cy_437),
    .O(\DLX_IDinst_RegFile_3_14/CYINIT )
  );
  X_MUX2 vga_top_vga1_Mmult__n0043_inst_cy_440_1885 (
    .IA(vga_top_vga1_gridvcounter[6]),
    .IB(\vga_top_vga1_Mmult__n0043_inst_lut2_320/CYINIT ),
    .SEL(vga_top_vga1_Mmult__n0043_inst_lut2_307),
    .O(vga_top_vga1_Mmult__n0043_inst_cy_440)
  );
  X_XOR2 vga_top_vga1_Mmult__n0043_inst_sum_229 (
    .I0(\vga_top_vga1_Mmult__n0043_inst_lut2_320/CYINIT ),
    .I1(vga_top_vga1_Mmult__n0043_inst_lut2_307),
    .O(\vga_top_vga1_Mmult__n0043_inst_lut2_320/XORF )
  );
  defparam vga_top_vga1_Mmult__n0043_inst_lut2_3071.INIT = 16'h55AA;
  X_LUT4 vga_top_vga1_Mmult__n0043_inst_lut2_3071 (
    .ADR0(vga_top_vga1_gridvcounter[6]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_gridvcounter[4]),
    .O(vga_top_vga1_Mmult__n0043_inst_lut2_307)
  );
  defparam vga_top_vga1_Mmult__n0043_inst_lut2_3081.INIT = 16'h6666;
  X_LUT4 vga_top_vga1_Mmult__n0043_inst_lut2_3081 (
    .ADR0(vga_top_vga1_gridvcounter[7]),
    .ADR1(vga_top_vga1_gridvcounter[5]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(vga_top_vga1_Mmult__n0043_inst_lut2_308)
  );
  X_BUF \vga_top_vga1_Mmult__n0043_inst_lut2_320/COUTUSED  (
    .I(\vga_top_vga1_Mmult__n0043_inst_lut2_320/CYMUXG ),
    .O(vga_top_vga1_Mmult__n0043_inst_cy_441)
  );
  X_BUF \vga_top_vga1_Mmult__n0043_inst_lut2_320/XUSED  (
    .I(\vga_top_vga1_Mmult__n0043_inst_lut2_320/XORF ),
    .O(vga_top_vga1_Mmult__n0043_inst_lut2_320)
  );
  X_BUF \vga_top_vga1_Mmult__n0043_inst_lut2_320/YUSED  (
    .I(\vga_top_vga1_Mmult__n0043_inst_lut2_320/XORG ),
    .O(vga_top_vga1_Mmult__n0043_inst_lut2_321)
  );
  X_MUX2 vga_top_vga1_Mmult__n0043_inst_cy_441_1886 (
    .IA(vga_top_vga1_gridvcounter[7]),
    .IB(vga_top_vga1_Mmult__n0043_inst_cy_440),
    .SEL(vga_top_vga1_Mmult__n0043_inst_lut2_308),
    .O(\vga_top_vga1_Mmult__n0043_inst_lut2_320/CYMUXG )
  );
  X_XOR2 vga_top_vga1_Mmult__n0043_inst_sum_230 (
    .I0(vga_top_vga1_Mmult__n0043_inst_cy_440),
    .I1(vga_top_vga1_Mmult__n0043_inst_lut2_308),
    .O(\vga_top_vga1_Mmult__n0043_inst_lut2_320/XORG )
  );
  X_BUF \vga_top_vga1_Mmult__n0043_inst_lut2_320/CYINIT_1887  (
    .I(vga_top_vga1_Mmult__n0043_inst_cy_439),
    .O(\vga_top_vga1_Mmult__n0043_inst_lut2_320/CYINIT )
  );
  defparam DLX_IDinst_RegFile_29_21_1888.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_29_21_1888 (
    .I(DLX_IDinst_WB_data_eff[21]),
    .CE(DLX_IDinst__n0608),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_29_21)
  );
  X_MUX2 vga_top_vga1_Mmult__n0043_inst_cy_442_1889 (
    .IA(vga_top_vga1_gridvcounter[8]),
    .IB(\vga_top_vga1_Mmult__n0043_inst_lut2_322/CYINIT ),
    .SEL(vga_top_vga1_Mmult__n0043_inst_lut2_309),
    .O(vga_top_vga1_Mmult__n0043_inst_cy_442)
  );
  X_XOR2 vga_top_vga1_Mmult__n0043_inst_sum_231 (
    .I0(\vga_top_vga1_Mmult__n0043_inst_lut2_322/CYINIT ),
    .I1(vga_top_vga1_Mmult__n0043_inst_lut2_309),
    .O(\vga_top_vga1_Mmult__n0043_inst_lut2_322/XORF )
  );
  defparam vga_top_vga1_Mmult__n0043_inst_lut2_3091.INIT = 16'h55AA;
  X_LUT4 vga_top_vga1_Mmult__n0043_inst_lut2_3091 (
    .ADR0(vga_top_vga1_gridvcounter[8]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_gridvcounter[6]),
    .O(vga_top_vga1_Mmult__n0043_inst_lut2_309)
  );
  defparam \$BEL_0 .INIT = 16'hAAAA;
  X_LUT4 \$BEL_0  (
    .ADR0(vga_top_vga1_gridvcounter[7]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\$SIG_0 )
  );
  X_BUF \vga_top_vga1_Mmult__n0043_inst_lut2_322/XUSED  (
    .I(\vga_top_vga1_Mmult__n0043_inst_lut2_322/XORF ),
    .O(vga_top_vga1_Mmult__n0043_inst_lut2_322)
  );
  X_BUF \vga_top_vga1_Mmult__n0043_inst_lut2_322/YUSED  (
    .I(\vga_top_vga1_Mmult__n0043_inst_lut2_322/XORG ),
    .O(vga_top_vga1_Mmult__n0043_inst_lut2_323)
  );
  X_XOR2 vga_top_vga1_Mmult__n0043_inst_sum_232 (
    .I0(vga_top_vga1_Mmult__n0043_inst_cy_442),
    .I1(\$SIG_0 ),
    .O(\vga_top_vga1_Mmult__n0043_inst_lut2_322/XORG )
  );
  X_BUF \vga_top_vga1_Mmult__n0043_inst_lut2_322/CYINIT_1890  (
    .I(vga_top_vga1_Mmult__n0043_inst_cy_441),
    .O(\vga_top_vga1_Mmult__n0043_inst_lut2_322/CYINIT )
  );
  X_ONE \vga_top_vga1_Mcompar__n0034_inst_cy_329/LOGIC_ONE_1891  (
    .O(\vga_top_vga1_Mcompar__n0034_inst_cy_329/LOGIC_ONE )
  );
  X_ZERO \vga_top_vga1_Mcompar__n0034_inst_cy_329/LOGIC_ZERO_1892  (
    .O(\vga_top_vga1_Mcompar__n0034_inst_cy_329/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0034_inst_cy_328_1893 (
    .IA(\vga_top_vga1_Mcompar__n0034_inst_cy_329/LOGIC_ZERO ),
    .IB(\vga_top_vga1_Mcompar__n0034_inst_cy_329/LOGIC_ONE ),
    .SEL(\$SIG_1 ),
    .O(vga_top_vga1_Mcompar__n0034_inst_cy_328)
  );
  defparam \$BEL_1 .INIT = 16'hFF00;
  X_LUT4 \$BEL_1  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[2]),
    .O(\$SIG_1 )
  );
  defparam \$BEL_2 .INIT = 16'hFF00;
  X_LUT4 \$BEL_2  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[2]),
    .O(\$SIG_2 )
  );
  X_BUF \vga_top_vga1_Mcompar__n0034_inst_cy_329/COUTUSED  (
    .I(\vga_top_vga1_Mcompar__n0034_inst_cy_329/CYMUXG ),
    .O(vga_top_vga1_Mcompar__n0034_inst_cy_329)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0034_inst_cy_329_1894 (
    .IA(\vga_top_vga1_Mcompar__n0034_inst_cy_329/LOGIC_ZERO ),
    .IB(vga_top_vga1_Mcompar__n0034_inst_cy_328),
    .SEL(\$SIG_2 ),
    .O(\vga_top_vga1_Mcompar__n0034_inst_cy_329/CYMUXG )
  );
  X_ONE \DLX_IDinst_RegFile_6_13/LOGIC_ONE_1895  (
    .O(\DLX_IDinst_RegFile_6_13/LOGIC_ONE )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0034_inst_cy_330_1896 (
    .IA(\DLX_IDinst_RegFile_6_13/LOGIC_ONE ),
    .IB(\DLX_IDinst_RegFile_6_13/CYINIT ),
    .SEL(vga_top_vga1_Mcompar__n0034_inst_lut2_262),
    .O(vga_top_vga1_Mcompar__n0034_inst_cy_330)
  );
  defparam vga_top_vga1_Mcompar__n0034_inst_lut2_2621.INIT = 16'h0055;
  X_LUT4 vga_top_vga1_Mcompar__n0034_inst_lut2_2621 (
    .ADR0(vga_top_vga1_hcounter[3]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[4]),
    .O(vga_top_vga1_Mcompar__n0034_inst_lut2_262)
  );
  defparam vga_top_vga1_Mcompar__n0034_inst_lut2_2631.INIT = 16'h000F;
  X_LUT4 vga_top_vga1_Mcompar__n0034_inst_lut2_2631 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_hcounter[3]),
    .ADR3(vga_top_vga1_hcounter[4]),
    .O(vga_top_vga1_Mcompar__n0034_inst_lut2_263)
  );
  X_BUF \DLX_IDinst_RegFile_6_13/COUTUSED  (
    .I(\DLX_IDinst_RegFile_6_13/CYMUXG ),
    .O(vga_top_vga1_Mcompar__n0034_inst_cy_331)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0034_inst_cy_331_1897 (
    .IA(\DLX_IDinst_RegFile_6_13/LOGIC_ONE ),
    .IB(vga_top_vga1_Mcompar__n0034_inst_cy_330),
    .SEL(vga_top_vga1_Mcompar__n0034_inst_lut2_263),
    .O(\DLX_IDinst_RegFile_6_13/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_6_13/CYINIT_1898  (
    .I(vga_top_vga1_Mcompar__n0034_inst_cy_329),
    .O(\DLX_IDinst_RegFile_6_13/CYINIT )
  );
  X_ZERO \vga_top_vga1_Mcompar__n0034_inst_cy_333/LOGIC_ZERO_1899  (
    .O(\vga_top_vga1_Mcompar__n0034_inst_cy_333/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0034_inst_cy_332_1900 (
    .IA(\vga_top_vga1_Mcompar__n0034_inst_cy_333/LOGIC_ZERO ),
    .IB(\vga_top_vga1_Mcompar__n0034_inst_cy_333/CYINIT ),
    .SEL(\$SIG_3 ),
    .O(vga_top_vga1_Mcompar__n0034_inst_cy_332)
  );
  defparam \$BEL_3 .INIT = 16'hAAAA;
  X_LUT4 \$BEL_3  (
    .ADR0(vga_top_vga1_hcounter[5]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\$SIG_3 )
  );
  defparam \$BEL_4 .INIT = 16'hFF00;
  X_LUT4 \$BEL_4  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[5]),
    .O(\$SIG_4 )
  );
  X_BUF \vga_top_vga1_Mcompar__n0034_inst_cy_333/COUTUSED  (
    .I(\vga_top_vga1_Mcompar__n0034_inst_cy_333/CYMUXG ),
    .O(vga_top_vga1_Mcompar__n0034_inst_cy_333)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0034_inst_cy_333_1901 (
    .IA(\vga_top_vga1_Mcompar__n0034_inst_cy_333/LOGIC_ZERO ),
    .IB(vga_top_vga1_Mcompar__n0034_inst_cy_332),
    .SEL(\$SIG_4 ),
    .O(\vga_top_vga1_Mcompar__n0034_inst_cy_333/CYMUXG )
  );
  X_BUF \vga_top_vga1_Mcompar__n0034_inst_cy_333/CYINIT_1902  (
    .I(vga_top_vga1_Mcompar__n0034_inst_cy_331),
    .O(\vga_top_vga1_Mcompar__n0034_inst_cy_333/CYINIT )
  );
  X_ONE \vga_top_vga1_Mcompar__n0034_inst_cy_335/LOGIC_ONE_1903  (
    .O(\vga_top_vga1_Mcompar__n0034_inst_cy_335/LOGIC_ONE )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0034_inst_cy_334_1904 (
    .IA(\vga_top_vga1_Mcompar__n0034_inst_cy_335/LOGIC_ONE ),
    .IB(\vga_top_vga1_Mcompar__n0034_inst_cy_335/CYINIT ),
    .SEL(vga_top_vga1_Mcompar__n0034_inst_lut2_264),
    .O(vga_top_vga1_Mcompar__n0034_inst_cy_334)
  );
  defparam vga_top_vga1_Mcompar__n0034_inst_lut2_2641.INIT = 16'h0055;
  X_LUT4 vga_top_vga1_Mcompar__n0034_inst_lut2_2641 (
    .ADR0(vga_top_vga1_hcounter[7]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[6]),
    .O(vga_top_vga1_Mcompar__n0034_inst_lut2_264)
  );
  defparam vga_top_vga1_Mcompar__n0034_inst_lut2_2651.INIT = 16'h0033;
  X_LUT4 vga_top_vga1_Mcompar__n0034_inst_lut2_2651 (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_hcounter[6]),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[7]),
    .O(vga_top_vga1_Mcompar__n0034_inst_lut2_265)
  );
  X_BUF \vga_top_vga1_Mcompar__n0034_inst_cy_335/COUTUSED  (
    .I(\vga_top_vga1_Mcompar__n0034_inst_cy_335/CYMUXG ),
    .O(vga_top_vga1_Mcompar__n0034_inst_cy_335)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0034_inst_cy_335_1905 (
    .IA(\vga_top_vga1_Mcompar__n0034_inst_cy_335/LOGIC_ONE ),
    .IB(vga_top_vga1_Mcompar__n0034_inst_cy_334),
    .SEL(vga_top_vga1_Mcompar__n0034_inst_lut2_265),
    .O(\vga_top_vga1_Mcompar__n0034_inst_cy_335/CYMUXG )
  );
  X_BUF \vga_top_vga1_Mcompar__n0034_inst_cy_335/CYINIT_1906  (
    .I(vga_top_vga1_Mcompar__n0034_inst_cy_333),
    .O(\vga_top_vga1_Mcompar__n0034_inst_cy_335/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_14_29/LOGIC_ZERO_1907  (
    .O(\DLX_IDinst_RegFile_14_29/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0034_inst_cy_336_1908 (
    .IA(\DLX_IDinst_RegFile_14_29/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_14_29/CYINIT ),
    .SEL(vga_top_vga1_Mcompar__n0034_inst_lut2_266),
    .O(vga_top_vga1_Mcompar__n0034_inst_cy_336)
  );
  defparam vga_top_vga1_Mcompar__n0034_inst_lut2_2661.INIT = 16'h8888;
  X_LUT4 vga_top_vga1_Mcompar__n0034_inst_lut2_2661 (
    .ADR0(vga_top_vga1_hcounter[9]),
    .ADR1(vga_top_vga1_hcounter[8]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(vga_top_vga1_Mcompar__n0034_inst_lut2_266)
  );
  defparam vga_top_vga1_Mcompar__n0034_inst_lut2_2671.INIT = 16'hF000;
  X_LUT4 vga_top_vga1_Mcompar__n0034_inst_lut2_2671 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_hcounter[9]),
    .ADR3(vga_top_vga1_hcounter[8]),
    .O(vga_top_vga1_Mcompar__n0034_inst_lut2_267)
  );
  X_BUF \DLX_IDinst_RegFile_14_29/COUTUSED  (
    .I(\DLX_IDinst_RegFile_14_29/CYMUXG ),
    .O(vga_top_vga1_Mcompar__n0034_inst_cy_337)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0034_inst_cy_337_1909 (
    .IA(\DLX_IDinst_RegFile_14_29/LOGIC_ZERO ),
    .IB(vga_top_vga1_Mcompar__n0034_inst_cy_336),
    .SEL(vga_top_vga1_Mcompar__n0034_inst_lut2_267),
    .O(\DLX_IDinst_RegFile_14_29/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_14_29/CYINIT_1910  (
    .I(vga_top_vga1_Mcompar__n0034_inst_cy_335),
    .O(\DLX_IDinst_RegFile_14_29/CYINIT )
  );
  X_ONE \vga_top_vga1__n0034/LOGIC_ONE_1911  (
    .O(\vga_top_vga1__n0034/LOGIC_ONE )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0034_inst_cy_338_1912 (
    .IA(\vga_top_vga1__n0034/LOGIC_ONE ),
    .IB(\vga_top_vga1__n0034/CYINIT ),
    .SEL(vga_top_vga1_Mcompar__n0034_inst_lut4_1099),
    .O(vga_top_vga1_Mcompar__n0034_inst_cy_338)
  );
  defparam vga_top_vga1_Mcompar__n0034_inst_lut4_10991.INIT = 16'h0001;
  X_LUT4 vga_top_vga1_Mcompar__n0034_inst_lut4_10991 (
    .ADR0(vga_top_vga1_hcounter[10]),
    .ADR1(vga_top_vga1_hcounter[11]),
    .ADR2(vga_top_vga1_hcounter[12]),
    .ADR3(vga_top_vga1_hcounter[13]),
    .O(vga_top_vga1_Mcompar__n0034_inst_lut4_1099)
  );
  defparam vga_top_vga1_Mcompar__n0034_inst_lut2_2681.INIT = 16'h000F;
  X_LUT4 vga_top_vga1_Mcompar__n0034_inst_lut2_2681 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_hcounter[15]),
    .ADR3(vga_top_vga1_hcounter[14]),
    .O(vga_top_vga1_Mcompar__n0034_inst_lut2_268)
  );
  X_BUF \vga_top_vga1__n0034/COUTUSED  (
    .I(\vga_top_vga1__n0034/CYMUXG ),
    .O(vga_top_vga1__n0034)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0034_inst_cy_339 (
    .IA(\vga_top_vga1__n0034/LOGIC_ONE ),
    .IB(vga_top_vga1_Mcompar__n0034_inst_cy_338),
    .SEL(vga_top_vga1_Mcompar__n0034_inst_lut2_268),
    .O(\vga_top_vga1__n0034/CYMUXG )
  );
  X_BUF \vga_top_vga1__n0034/CYINIT_1913  (
    .I(vga_top_vga1_Mcompar__n0034_inst_cy_337),
    .O(\vga_top_vga1__n0034/CYINIT )
  );
  X_ONE \DLX_IDinst_Mmux__COND_4_inst_cy_97/LOGIC_ONE_1914  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_97/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_4_inst_cy_97/LOGIC_ZERO_1915  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_97/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_96_1916 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_97/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_4_inst_cy_97/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_155),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_96)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1551.INIT = 16'hFB3B;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1551 (
    .ADR0(DLX_IDinst_RegFile_0_6),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_43),
    .ADR2(DLX_IDinst_jtarget[16]),
    .ADR3(DLX_IDinst_RegFile_1_6),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_155)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1561.INIT = 16'hACFF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1561 (
    .ADR0(DLX_IDinst_RegFile_3_6),
    .ADR1(DLX_IDinst_RegFile_2_6),
    .ADR2(DLX_IDinst_jtarget[16]),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_44),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_156)
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_cy_97/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_4_inst_cy_97/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_97)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_97_1917 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_97/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_96),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_156),
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_97/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mmux__COND_4_inst_cy_193/LOGIC_ONE_1918  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_193/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_4_inst_cy_193/LOGIC_ZERO_1919  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_193/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_192_1920 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_193/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_4_inst_cy_193/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_251),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_192)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2511.INIT = 16'hF7B3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2511 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_43),
    .ADR2(DLX_IDinst_RegFile_1_12),
    .ADR3(DLX_IDinst_RegFile_0_12),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_251)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2521.INIT = 16'hF7B3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2521 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_44),
    .ADR2(DLX_IDinst_RegFile_3_12),
    .ADR3(DLX_IDinst_RegFile_2_12),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_252)
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_cy_193/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_4_inst_cy_193/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_193)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_193_1921 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_193/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_192),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_252),
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_193/CYMUXG )
  );
  X_ONE \DLX_EXinst_reg_write_EX/LOGIC_ONE_1922  (
    .O(\DLX_EXinst_reg_write_EX/LOGIC_ONE )
  );
  X_ZERO \DLX_EXinst_reg_write_EX/LOGIC_ZERO_1923  (
    .O(\DLX_EXinst_reg_write_EX/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_112_1924 (
    .IA(\DLX_EXinst_reg_write_EX/LOGIC_ZERO ),
    .IB(\DLX_EXinst_reg_write_EX/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_171),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_112)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1711.INIT = 16'hE2FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1711 (
    .ADR0(DLX_IDinst_RegFile_0_7),
    .ADR1(DLX_IDinst_jtarget[16]),
    .ADR2(DLX_IDinst_RegFile_1_7),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_43),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_171)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1721.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1721 (
    .ADR0(DLX_IDinst_RegFile_2_7),
    .ADR1(DLX_IDinst_jtarget[16]),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_44),
    .ADR3(DLX_IDinst_RegFile_3_7),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_172)
  );
  X_BUF \DLX_EXinst_reg_write_EX/COUTUSED  (
    .I(\DLX_EXinst_reg_write_EX/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_113)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_113_1925 (
    .IA(\DLX_EXinst_reg_write_EX/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_112),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_172),
    .O(\DLX_EXinst_reg_write_EX/CYMUXG )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_4_inst_cy_121/LOGIC_ZERO_1926  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_121/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_120_1927 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_121/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_4_inst_cy_121/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_179),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_120)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1791.INIT = 16'hBF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1791 (
    .ADR0(DLX_IDinst_RegFile_17_7),
    .ADR1(DLX_IDinst_jtarget[16]),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_51),
    .ADR3(DLX_IDinst_RegFile_16_7),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_179)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1801.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1801 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_52),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR2(DLX_IDinst_RegFile_18_7),
    .ADR3(DLX_IDinst_RegFile_19_7),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_180)
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_cy_121/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_4_inst_cy_121/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_121)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_121_1928 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_121/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_120),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_180),
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_121/CYMUXG )
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_cy_121/CYINIT_1929  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_119),
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_121/CYINIT )
  );
  X_ONE \DLX_IDinst_Mmux__COND_4_inst_cy_209/LOGIC_ONE_1930  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_209/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_4_inst_cy_209/LOGIC_ZERO_1931  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_209/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_208_1932 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_209/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_4_inst_cy_209/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_267),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_208)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2671.INIT = 16'hBF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2671 (
    .ADR0(DLX_IDinst_RegFile_1_13),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_43),
    .ADR3(DLX_IDinst_RegFile_0_13),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_267)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2681.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2681 (
    .ADR0(DLX_IDinst_RegFile_3_13),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_44),
    .ADR2(DLX_IDinst_RegFile_2_13),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_268)
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_cy_209/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_4_inst_cy_209/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_209)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_209_1933 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_209/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_208),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_268),
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_209/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mmux__COND_4_inst_cy_129/LOGIC_ONE_1934  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_129/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_4_inst_cy_129/LOGIC_ZERO_1935  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_129/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_128_1936 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_129/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_4_inst_cy_129/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_187),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_128)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1871.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1871 (
    .ADR0(DLX_IDinst_RegFile_0_8),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_43),
    .ADR2(DLX_IDinst_RegFile_1_8),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_187)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1881.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1881 (
    .ADR0(DLX_IDinst_RegFile_3_8),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_44),
    .ADR2(DLX_IDinst_RegFile_2_8),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_188)
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_cy_129/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_4_inst_cy_129/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_129)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_129_1937 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_129/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_128),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_188),
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_129/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mmux__COND_4_inst_cy_289/LOGIC_ONE_1938  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_289/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_4_inst_cy_289/LOGIC_ZERO_1939  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_289/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_288_1940 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_289/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_4_inst_cy_289/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_347),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_288)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3471.INIT = 16'hDFD5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3471 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_43),
    .ADR1(DLX_IDinst_RegFile_1_18),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR3(DLX_IDinst_RegFile_0_18),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_347)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3481.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3481 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR1(DLX_IDinst_RegFile_2_18),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_44),
    .ADR3(DLX_IDinst_RegFile_3_18),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_348)
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_cy_289/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_4_inst_cy_289/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_289)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_289_1941 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_289/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_288),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_348),
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_289/CYMUXG )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_4_inst_cy_295/LOGIC_ZERO_1942  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_295/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_294_1943 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_295/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_4_inst_cy_295/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_353),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_294)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3531.INIT = 16'hB8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3531 (
    .ADR0(DLX_IDinst_RegFile_13_18),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR2(DLX_IDinst_RegFile_12_18),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_49),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_353)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3541.INIT = 16'hBFB3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3541 (
    .ADR0(DLX_IDinst_RegFile_15_18),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_50),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR3(DLX_IDinst_RegFile_14_18),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_354)
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_cy_295/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_4_inst_cy_295/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_295)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_295_1944 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_295/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_294),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_354),
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_295/CYMUXG )
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_cy_295/CYINIT_1945  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_293),
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_295/CYINIT )
  );
  X_ONE \DLX_IDinst_Mmux__COND_4_inst_cy_305/LOGIC_ONE_1946  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_305/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_4_inst_cy_305/LOGIC_ZERO_1947  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_305/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_304_1948 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_305/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_4_inst_cy_305/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_363),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_304)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3631.INIT = 16'hE2FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3631 (
    .ADR0(DLX_IDinst_RegFile_0_19),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR2(DLX_IDinst_RegFile_1_19),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_43),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_363)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3641.INIT = 16'hCFAF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3641 (
    .ADR0(DLX_IDinst_RegFile_2_19),
    .ADR1(DLX_IDinst_RegFile_3_19),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_44),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_364)
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_cy_305/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_4_inst_cy_305/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_305)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_305_1949 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_305/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_304),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_364),
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_305/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mmux__COND_4_inst_cy_225/LOGIC_ONE_1950  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_225/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_4_inst_cy_225/LOGIC_ZERO_1951  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_225/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_224_1952 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_225/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_4_inst_cy_225/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_283),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_224)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2831.INIT = 16'hBFB3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2831 (
    .ADR0(DLX_IDinst_RegFile_1_14),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_43),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR3(DLX_IDinst_RegFile_0_14),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_283)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2841.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2841 (
    .ADR0(DLX_IDinst_RegFile_2_14),
    .ADR1(DLX_IDinst_RegFile_3_14),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_44),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_284)
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_cy_225/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_4_inst_cy_225/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_225)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_225_1953 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_225/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_224),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_284),
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_225/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mmux__COND_4_inst_cy_145/LOGIC_ONE_1954  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_145/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_4_inst_cy_145/LOGIC_ZERO_1955  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_145/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_144_1956 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_145/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_4_inst_cy_145/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_203),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_144)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2031.INIT = 16'hE4FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2031 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR1(DLX_IDinst_RegFile_0_9),
    .ADR2(DLX_IDinst_RegFile_1_9),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_43),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_203)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2041.INIT = 16'hD8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2041 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR1(DLX_IDinst_RegFile_3_9),
    .ADR2(DLX_IDinst_RegFile_2_9),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_44),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_204)
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_cy_145/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_4_inst_cy_145/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_145)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_145_1957 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_145/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_144),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_204),
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_145/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mmux__COND_4_inst_cy_401/LOGIC_ONE_1958  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_401/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_4_inst_cy_401/LOGIC_ZERO_1959  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_401/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_400_1960 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_401/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_4_inst_cy_401/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_459),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_400)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4591.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4591 (
    .ADR0(DLX_IDinst_RegFile_0_25),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_43),
    .ADR2(DLX_IDinst_RegFile_1_25),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_459)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4601.INIT = 16'hDDF5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4601 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_44),
    .ADR1(DLX_IDinst_RegFile_3_25),
    .ADR2(DLX_IDinst_RegFile_2_25),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_460)
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_cy_401/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_4_inst_cy_401/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_401)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_401_1961 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_401/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_400),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_460),
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_401/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mmux__COND_4_inst_cy_321/LOGIC_ONE_1962  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_321/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_4_inst_cy_321/LOGIC_ZERO_1963  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_321/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_320_1964 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_321/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_4_inst_cy_321/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_379),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_320)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3791.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3791 (
    .ADR0(DLX_IDinst_RegFile_1_20),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_43),
    .ADR2(DLX_IDinst_RegFile_0_20),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_379)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3801.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3801 (
    .ADR0(DLX_IDinst_RegFile_2_20),
    .ADR1(DLX_IDinst_RegFile_3_20),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_44),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_380)
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_cy_321/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_4_inst_cy_321/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_321)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_321_1965 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_321/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_320),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_380),
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_321/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mmux__COND_4_inst_cy_241/LOGIC_ONE_1966  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_241/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_4_inst_cy_241/LOGIC_ZERO_1967  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_241/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_240_1968 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_241/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_4_inst_cy_241/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_299),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_240)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2991.INIT = 16'hBFB3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2991 (
    .ADR0(DLX_IDinst_RegFile_1_15),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_43),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR3(DLX_IDinst_RegFile_0_15),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_299)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3001.INIT = 16'hACFF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3001 (
    .ADR0(DLX_IDinst_RegFile_3_15),
    .ADR1(DLX_IDinst_RegFile_2_15),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_44),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_300)
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_cy_241/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_4_inst_cy_241/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_241)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_241_1969 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_241/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_240),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_300),
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_241/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mmux__COND_4_inst_cy_161/LOGIC_ONE_1970  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_161/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_4_inst_cy_161/LOGIC_ZERO_1971  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_161/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_160_1972 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_161/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_4_inst_cy_161/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_219),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_160)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2191.INIT = 16'hFB3B;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2191 (
    .ADR0(DLX_IDinst_RegFile_0_10),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_43),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR3(DLX_IDinst_RegFile_1_10),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_219)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2201.INIT = 16'hF7B3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2201 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_44),
    .ADR2(DLX_IDinst_RegFile_3_10),
    .ADR3(DLX_IDinst_RegFile_2_10),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_220)
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_cy_161/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_4_inst_cy_161/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_161)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_161_1973 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_161/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_160),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_220),
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_161/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mmux__COND_4_inst_cy_497/LOGIC_ONE_1974  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_497/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_4_inst_cy_497/LOGIC_ZERO_1975  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_497/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_496_1976 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_497/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_4_inst_cy_497/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_555),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_496)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5551.INIT = 16'hB8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5551 (
    .ADR0(DLX_IDinst_RegFile_1_31),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR2(DLX_IDinst_RegFile_0_31),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_43),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_555)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5561.INIT = 16'hE4FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5561 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR1(DLX_IDinst_RegFile_2_31),
    .ADR2(DLX_IDinst_RegFile_3_31),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_44),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_556)
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_cy_497/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_4_inst_cy_497/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_497)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_497_1977 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_497/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_496),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_556),
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_497/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mmux__COND_4_inst_cy_417/LOGIC_ONE_1978  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_417/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_4_inst_cy_417/LOGIC_ZERO_1979  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_417/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_416_1980 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_417/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_4_inst_cy_417/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_475),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_416)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4751.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4751 (
    .ADR0(DLX_IDinst_RegFile_0_26),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_43),
    .ADR3(DLX_IDinst_RegFile_1_26),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_475)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4761.INIT = 16'hE4FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4761 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR1(DLX_IDinst_RegFile_2_26),
    .ADR2(DLX_IDinst_RegFile_3_26),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_44),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_476)
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_cy_417/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_4_inst_cy_417/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_417)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_417_1981 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_417/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_416),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_476),
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_417/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mmux__COND_4_inst_cy_337/LOGIC_ONE_1982  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_337/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_4_inst_cy_337/LOGIC_ZERO_1983  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_337/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_336_1984 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_337/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_4_inst_cy_337/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_395),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_336)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3951.INIT = 16'hE4FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3951 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR1(DLX_IDinst_RegFile_0_21),
    .ADR2(DLX_IDinst_RegFile_1_21),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_43),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_395)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3961.INIT = 16'hFB73;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3961 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_44),
    .ADR2(DLX_IDinst_RegFile_2_21),
    .ADR3(DLX_IDinst_RegFile_3_21),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_396)
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_cy_337/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_4_inst_cy_337/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_337)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_337_1985 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_337/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_336),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_396),
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_337/CYMUXG )
  );
  X_ONE \DLX_EXinst_reg_out_B_EX<3>/LOGIC_ONE_1986  (
    .O(\DLX_EXinst_reg_out_B_EX<3>/LOGIC_ONE )
  );
  X_ZERO \DLX_EXinst_reg_out_B_EX<3>/LOGIC_ZERO_1987  (
    .O(\DLX_EXinst_reg_out_B_EX<3>/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_256_1988 (
    .IA(\DLX_EXinst_reg_out_B_EX<3>/LOGIC_ZERO ),
    .IB(\DLX_EXinst_reg_out_B_EX<3>/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_315),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_256)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3151.INIT = 16'hE2FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3151 (
    .ADR0(DLX_IDinst_RegFile_0_16),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR2(DLX_IDinst_RegFile_1_16),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_43),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_315)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3161.INIT = 16'hF7B3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3161 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_44),
    .ADR2(DLX_IDinst_RegFile_3_16),
    .ADR3(DLX_IDinst_RegFile_2_16),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_316)
  );
  X_BUF \DLX_EXinst_reg_out_B_EX<3>/COUTUSED  (
    .I(\DLX_EXinst_reg_out_B_EX<3>/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_257)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_257_1989 (
    .IA(\DLX_EXinst_reg_out_B_EX<3>/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_256),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_316),
    .O(\DLX_EXinst_reg_out_B_EX<3>/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mmux__COND_4_inst_cy_177/LOGIC_ONE_1990  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_177/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_4_inst_cy_177/LOGIC_ZERO_1991  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_177/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_176_1992 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_177/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_4_inst_cy_177/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_235),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_176)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2351.INIT = 16'hAFCF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2351 (
    .ADR0(DLX_IDinst_RegFile_1_11),
    .ADR1(DLX_IDinst_RegFile_0_11),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_43),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_235)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2361.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2361 (
    .ADR0(DLX_IDinst_RegFile_3_11),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_44),
    .ADR2(DLX_IDinst_RegFile_2_11),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_236)
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_cy_177/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_4_inst_cy_177/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_177)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_177_1993 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_177/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_176),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_236),
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_177/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mmux__COND_4_inst_cy_433/LOGIC_ONE_1994  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_433/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_4_inst_cy_433/LOGIC_ZERO_1995  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_433/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_432_1996 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_433/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_4_inst_cy_433/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_491),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_432)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4911.INIT = 16'hDFD5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4911 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_43),
    .ADR1(DLX_IDinst_RegFile_1_27),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR3(DLX_IDinst_RegFile_0_27),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_491)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4921.INIT = 16'hDF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4921 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR1(DLX_IDinst_RegFile_3_27),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_44),
    .ADR3(DLX_IDinst_RegFile_2_27),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_492)
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_cy_433/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_4_inst_cy_433/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_433)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_433_1997 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_433/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_432),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_492),
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_433/CYMUXG )
  );
  defparam DLX_IDinst_RegFile_29_30_1998.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_29_30_1998 (
    .I(DLX_IDinst_WB_data_eff[30]),
    .CE(DLX_IDinst__n0608),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_29_30)
  );
  X_ONE \DLX_IDinst_Mmux__COND_4_inst_cy_353/LOGIC_ONE_1999  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_353/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_4_inst_cy_353/LOGIC_ZERO_2000  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_353/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_352_2001 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_353/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_4_inst_cy_353/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_411),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_352)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4111.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4111 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR1(DLX_IDinst_RegFile_0_22),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_43),
    .ADR3(DLX_IDinst_RegFile_1_22),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_411)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4121.INIT = 16'hDF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4121 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR1(DLX_IDinst_RegFile_3_22),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_44),
    .ADR3(DLX_IDinst_RegFile_2_22),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_412)
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_cy_353/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_4_inst_cy_353/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_353)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_353_2002 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_353/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_352),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_412),
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_353/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mmux__COND_4_inst_cy_273/LOGIC_ONE_2003  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_273/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_4_inst_cy_273/LOGIC_ZERO_2004  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_273/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_272_2005 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_273/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_4_inst_cy_273/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_331),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_272)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3311.INIT = 16'hAFCF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3311 (
    .ADR0(DLX_IDinst_RegFile_1_17),
    .ADR1(DLX_IDinst_RegFile_0_17),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_43),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_331)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3321.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3321 (
    .ADR0(DLX_IDinst_RegFile_2_17),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_44),
    .ADR3(DLX_IDinst_RegFile_3_17),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_332)
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_cy_273/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_4_inst_cy_273/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_273)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_273_2006 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_273/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_272),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_332),
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_273/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mmux__COND_4_inst_cy_449/LOGIC_ONE_2007  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_449/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_4_inst_cy_449/LOGIC_ZERO_2008  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_449/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_448_2009 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_449/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_4_inst_cy_449/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_507),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_448)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5071.INIT = 16'hF7B3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5071 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_43),
    .ADR2(DLX_IDinst_RegFile_1_28),
    .ADR3(DLX_IDinst_RegFile_0_28),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_507)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5081.INIT = 16'hFB3B;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5081 (
    .ADR0(DLX_IDinst_RegFile_2_28),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_44),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR3(DLX_IDinst_RegFile_3_28),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_508)
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_cy_449/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_4_inst_cy_449/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_449)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_449_2010 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_449/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_448),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_508),
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_449/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mmux__COND_4_inst_cy_369/LOGIC_ONE_2011  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_369/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_4_inst_cy_369/LOGIC_ZERO_2012  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_369/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_368_2013 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_369/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_4_inst_cy_369/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_427),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_368)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4271.INIT = 16'hDFD5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4271 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_43),
    .ADR1(DLX_IDinst_RegFile_1_23),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR3(DLX_IDinst_RegFile_0_23),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_427)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4281.INIT = 16'hBF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4281 (
    .ADR0(DLX_IDinst_RegFile_3_23),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_44),
    .ADR3(DLX_IDinst_RegFile_2_23),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_428)
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_cy_369/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_4_inst_cy_369/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_369)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_369_2014 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_369/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_368),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_428),
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_369/CYMUXG )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_4_inst_cy_381/LOGIC_ZERO_2015  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_381/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_380_2016 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_381/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_4_inst_cy_381/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_439),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_380)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4391.INIT = 16'hACFF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4391 (
    .ADR0(DLX_IDinst_RegFile_25_23),
    .ADR1(DLX_IDinst_RegFile_24_23),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_55),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_439)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4401.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4401 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_56),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR2(DLX_IDinst_RegFile_26_23),
    .ADR3(DLX_IDinst_RegFile_27_23),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_440)
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_cy_381/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_4_inst_cy_381/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_381)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_381_2017 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_381/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_380),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_440),
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_381/CYMUXG )
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_cy_381/CYINIT_2018  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_379),
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_381/CYINIT )
  );
  X_ONE \DLX_IDinst_Mmux__COND_4_inst_cy_465/LOGIC_ONE_2019  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_465/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_4_inst_cy_465/LOGIC_ZERO_2020  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_465/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_464_2021 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_465/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_4_inst_cy_465/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_523),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_464)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5231.INIT = 16'hAFCF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5231 (
    .ADR0(DLX_IDinst_RegFile_1_29),
    .ADR1(DLX_IDinst_RegFile_0_29),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_43),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_523)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5241.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5241 (
    .ADR0(DLX_IDinst_RegFile_2_29),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_44),
    .ADR2(DLX_IDinst_RegFile_3_29),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_524)
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_cy_465/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_4_inst_cy_465/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_465)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_465_2022 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_465/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_464),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_524),
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_465/CYMUXG )
  );
  defparam DLX_IDinst_RegFile_29_14_2023.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_29_14_2023 (
    .I(DLX_IDinst_WB_data_eff[14]),
    .CE(DLX_IDinst__n0608),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_29_14)
  );
  X_ZERO \DLX_IDinst_Mmux__COND_4_inst_cy_467/LOGIC_ZERO_2024  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_467/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_466_2025 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_467/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_4_inst_cy_467/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_525),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_466)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5251.INIT = 16'hAFCF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5251 (
    .ADR0(DLX_IDinst_RegFile_5_29),
    .ADR1(DLX_IDinst_RegFile_4_29),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_45),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_525)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5261.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5261 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_46),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR2(DLX_IDinst_RegFile_6_29),
    .ADR3(DLX_IDinst_RegFile_7_29),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_526)
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_cy_467/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_4_inst_cy_467/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_467)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_467_2026 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_467/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_466),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_526),
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_467/CYMUXG )
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_cy_467/CYINIT_2027  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_465),
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_467/CYINIT )
  );
  X_ONE \DLX_IDinst_Mmux__COND_4_inst_cy_385/LOGIC_ONE_2028  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_385/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_4_inst_cy_385/LOGIC_ZERO_2029  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_385/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_384_2030 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_385/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_4_inst_cy_385/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_443),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_384)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4431.INIT = 16'hFB3B;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4431 (
    .ADR0(DLX_IDinst_RegFile_0_24),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_43),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR3(DLX_IDinst_RegFile_1_24),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_443)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4441.INIT = 16'hFB73;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4441 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_44),
    .ADR2(DLX_IDinst_RegFile_2_24),
    .ADR3(DLX_IDinst_RegFile_3_24),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_444)
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_cy_385/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_4_inst_cy_385/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_385)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_385_2031 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_385/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_384),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_444),
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_385/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mmux__COND_4_inst_cy_481/LOGIC_ONE_2032  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_481/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_4_inst_cy_481/LOGIC_ZERO_2033  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_481/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_480_2034 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_481/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_4_inst_cy_481/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_539),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_480)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5391.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5391 (
    .ADR0(DLX_IDinst_RegFile_0_30),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_43),
    .ADR2(DLX_IDinst_RegFile_1_30),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_539)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5401.INIT = 16'hE4FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5401 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR1(DLX_IDinst_RegFile_2_30),
    .ADR2(DLX_IDinst_RegFile_3_30),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_44),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_540)
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_cy_481/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_4_inst_cy_481/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_481)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_481_2035 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_481/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_480),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_540),
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_481/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mmux__COND_4_inst_cy_1/LOGIC_ONE_2036  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_1/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_4_inst_cy_1/LOGIC_ZERO_2037  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_1/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_0_2038 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_1/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_4_inst_cy_1/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_59),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_0)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_591.INIT = 16'hBF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_591 (
    .ADR0(DLX_IDinst_RegFile_1_0),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_43),
    .ADR3(DLX_IDinst_RegFile_0_0),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_59)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_601.INIT = 16'hF5DD;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_601 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_44),
    .ADR1(DLX_IDinst_RegFile_2_0),
    .ADR2(DLX_IDinst_RegFile_3_0),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_60)
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_cy_1/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_4_inst_cy_1/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_1)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_1_2039 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_1/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_0),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_60),
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_1/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mmux__COND_4_inst_cy_17/LOGIC_ONE_2040  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_17/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_4_inst_cy_17/LOGIC_ZERO_2041  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_17/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_16_2042 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_17/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_4_inst_cy_17/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_75),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_16)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_751.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_751 (
    .ADR0(DLX_IDinst_RegFile_0_1),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_43),
    .ADR3(DLX_IDinst_RegFile_1_1),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_75)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_761.INIT = 16'hF7D5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_761 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_44),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR2(DLX_IDinst_RegFile_3_1),
    .ADR3(DLX_IDinst_RegFile_2_1),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_76)
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_cy_17/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_4_inst_cy_17/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_17)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_17_2043 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_17/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_16),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_76),
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_17/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mmux__COND_4_inst_cy_33/LOGIC_ONE_2044  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_33/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_4_inst_cy_33/LOGIC_ZERO_2045  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_33/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_32_2046 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_33/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_4_inst_cy_33/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_91),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_32)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_911.INIT = 16'hE2FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_911 (
    .ADR0(DLX_IDinst_RegFile_0_2),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR2(DLX_IDinst_RegFile_1_2),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_43),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_91)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_921.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_921 (
    .ADR0(DLX_IDinst_RegFile_2_2),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_44),
    .ADR2(DLX_IDinst_RegFile_3_2),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_92)
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_cy_33/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_4_inst_cy_33/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_33)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_33_2047 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_33/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_32),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_92),
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_33/CYMUXG )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_4_inst_cy_41/LOGIC_ZERO_2048  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_41/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_40_2049 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_41/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_4_inst_cy_41/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_99),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_40)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_991.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_991 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_51),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR2(DLX_IDinst_RegFile_16_2),
    .ADR3(DLX_IDinst_RegFile_17_2),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_99)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1001.INIT = 16'hF5DD;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1001 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_52),
    .ADR1(DLX_IDinst_RegFile_18_2),
    .ADR2(DLX_IDinst_RegFile_19_2),
    .ADR3(DLX_IDinst_jtarget[16]),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_100)
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_cy_41/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_4_inst_cy_41/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_41)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_41_2050 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_41/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_40),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_100),
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_41/CYMUXG )
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_cy_41/CYINIT_2051  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_39),
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_41/CYINIT )
  );
  X_ONE \DLX_IDinst_Cause_Reg<6>/LOGIC_ONE_2052  (
    .O(\DLX_IDinst_Cause_Reg<6>/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Cause_Reg<6>/LOGIC_ZERO_2053  (
    .O(\DLX_IDinst_Cause_Reg<6>/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_48_2054 (
    .IA(\DLX_IDinst_Cause_Reg<6>/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Cause_Reg<6>/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_107),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_48)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1071.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1071 (
    .ADR0(DLX_IDinst_RegFile_0_3),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_43),
    .ADR2(DLX_IDinst_RegFile_1_3),
    .ADR3(DLX_IDinst_jtarget[16]),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_107)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1081.INIT = 16'hDDF5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1081 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_44),
    .ADR1(DLX_IDinst_RegFile_3_3),
    .ADR2(DLX_IDinst_RegFile_2_3),
    .ADR3(DLX_IDinst_jtarget[16]),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_108)
  );
  X_BUF \DLX_IDinst_Cause_Reg<6>/COUTUSED  (
    .I(\DLX_IDinst_Cause_Reg<6>/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_49)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_49_2055 (
    .IA(\DLX_IDinst_Cause_Reg<6>/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_48),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_108),
    .O(\DLX_IDinst_Cause_Reg<6>/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mmux__COND_4_inst_cy_65/LOGIC_ONE_2056  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_65/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_4_inst_cy_65/LOGIC_ZERO_2057  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_65/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_64_2058 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_65/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_4_inst_cy_65/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_123),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_64)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1231.INIT = 16'hAFCF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1231 (
    .ADR0(DLX_IDinst_RegFile_1_4),
    .ADR1(DLX_IDinst_RegFile_0_4),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_43),
    .ADR3(DLX_IDinst_jtarget[16]),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_123)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1241.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1241 (
    .ADR0(DLX_IDinst_RegFile_2_4),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_44),
    .ADR2(DLX_IDinst_RegFile_3_4),
    .ADR3(DLX_IDinst_jtarget[16]),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_124)
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_cy_65/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_4_inst_cy_65/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_65)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_65_2059 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_65/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_64),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_124),
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_65/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mmux__COND_4_inst_cy_81/LOGIC_ONE_2060  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_81/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_4_inst_cy_81/LOGIC_ZERO_2061  (
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_81/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_80_2062 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_81/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_4_inst_cy_81/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_139),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_80)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1391.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1391 (
    .ADR0(DLX_IDinst_RegFile_1_5),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_43),
    .ADR2(DLX_IDinst_RegFile_0_5),
    .ADR3(DLX_IDinst_jtarget[16]),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_139)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_1401.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_1401 (
    .ADR0(DLX_IDinst_RegFile_3_5),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_44),
    .ADR2(DLX_IDinst_RegFile_2_5),
    .ADR3(DLX_IDinst_jtarget[16]),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_140)
  );
  X_BUF \DLX_IDinst_Mmux__COND_4_inst_cy_81/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_4_inst_cy_81/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_81)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_81_2063 (
    .IA(\DLX_IDinst_Mmux__COND_4_inst_cy_81/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_80),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_140),
    .O(\DLX_IDinst_Mmux__COND_4_inst_cy_81/CYMUXG )
  );
  X_ZERO \DLX_EXinst_Mcompar__n0065_inst_cy_167/LOGIC_ZERO_2064  (
    .O(\DLX_EXinst_Mcompar__n0065_inst_cy_167/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0065_inst_cy_166_2065 (
    .IA(DLX_IDinst_reg_out_A[0]),
    .IB(\DLX_EXinst_Mcompar__n0065_inst_cy_167/LOGIC_ZERO ),
    .SEL(DLX_EXinst_Mcompar__n0065_inst_lut2_102),
    .O(DLX_EXinst_Mcompar__n0065_inst_cy_166)
  );
  defparam DLX_EXinst_Mcompar__n0065_inst_lut2_1021.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0065_inst_lut2_1021 (
    .ADR0(DLX_IDinst_reg_out_A[0]),
    .ADR1(VCC),
    .ADR2(\DLX_IDinst_Imm[0] ),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0065_inst_lut2_102)
  );
  defparam DLX_EXinst_Mcompar__n0065_inst_lut2_1031.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0065_inst_lut2_1031 (
    .ADR0(DLX_IDinst_reg_out_A[1]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_Imm_1_1),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0065_inst_lut2_103)
  );
  X_BUF \DLX_EXinst_Mcompar__n0065_inst_cy_167/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0065_inst_cy_167/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0065_inst_cy_167)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0065_inst_cy_167_2066 (
    .IA(DLX_IDinst_reg_out_A[1]),
    .IB(DLX_EXinst_Mcompar__n0065_inst_cy_166),
    .SEL(DLX_EXinst_Mcompar__n0065_inst_lut2_103),
    .O(\DLX_EXinst_Mcompar__n0065_inst_cy_167/CYMUXG )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0065_inst_cy_168_2067 (
    .IA(DLX_IDinst_reg_out_A[2]),
    .IB(\DLX_IDinst_RegFile_3_0/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0065_inst_lut2_104),
    .O(DLX_EXinst_Mcompar__n0065_inst_cy_168)
  );
  defparam DLX_EXinst_Mcompar__n0065_inst_lut2_1041.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0065_inst_lut2_1041 (
    .ADR0(DLX_IDinst_reg_out_A[2]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_Imm_2_1),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0065_inst_lut2_104)
  );
  defparam DLX_EXinst_Mcompar__n0065_inst_lut2_1051.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0065_inst_lut2_1051 (
    .ADR0(DLX_IDinst_reg_out_A[3]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_Imm_3_1),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0065_inst_lut2_105)
  );
  X_BUF \DLX_IDinst_RegFile_3_0/COUTUSED  (
    .I(\DLX_IDinst_RegFile_3_0/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0065_inst_cy_169)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0065_inst_cy_169_2068 (
    .IA(DLX_IDinst_reg_out_A[3]),
    .IB(DLX_EXinst_Mcompar__n0065_inst_cy_168),
    .SEL(DLX_EXinst_Mcompar__n0065_inst_lut2_105),
    .O(\DLX_IDinst_RegFile_3_0/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_3_0/CYINIT_2069  (
    .I(DLX_EXinst_Mcompar__n0065_inst_cy_167),
    .O(\DLX_IDinst_RegFile_3_0/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0065_inst_cy_170_2070 (
    .IA(DLX_IDinst_reg_out_A[4]),
    .IB(\DLX_EXinst_Mcompar__n0065_inst_cy_171/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0065_inst_lut2_106),
    .O(DLX_EXinst_Mcompar__n0065_inst_cy_170)
  );
  defparam DLX_EXinst_Mcompar__n0065_inst_lut2_1061.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0065_inst_lut2_1061 (
    .ADR0(DLX_IDinst_reg_out_A[4]),
    .ADR1(VCC),
    .ADR2(\DLX_IDinst_Imm[4] ),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0065_inst_lut2_106)
  );
  defparam DLX_EXinst_Mcompar__n0065_inst_lut2_1071.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0065_inst_lut2_1071 (
    .ADR0(DLX_IDinst_reg_out_A[5]),
    .ADR1(\DLX_IDinst_Imm[5] ),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0065_inst_lut2_107)
  );
  X_BUF \DLX_EXinst_Mcompar__n0065_inst_cy_171/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0065_inst_cy_171/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0065_inst_cy_171)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0065_inst_cy_171_2071 (
    .IA(DLX_IDinst_reg_out_A[5]),
    .IB(DLX_EXinst_Mcompar__n0065_inst_cy_170),
    .SEL(DLX_EXinst_Mcompar__n0065_inst_lut2_107),
    .O(\DLX_EXinst_Mcompar__n0065_inst_cy_171/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0065_inst_cy_171/CYINIT_2072  (
    .I(DLX_EXinst_Mcompar__n0065_inst_cy_169),
    .O(\DLX_EXinst_Mcompar__n0065_inst_cy_171/CYINIT )
  );
  defparam DLX_IDinst_RegFile_29_22_2073.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_29_22_2073 (
    .I(DLX_IDinst_WB_data_eff[22]),
    .CE(DLX_IDinst__n0608),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_29_22)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0065_inst_cy_172_2074 (
    .IA(DLX_IDinst_reg_out_A[6]),
    .IB(\DLX_IDinst_RegFile_31_11/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0065_inst_lut2_108),
    .O(DLX_EXinst_Mcompar__n0065_inst_cy_172)
  );
  defparam DLX_EXinst_Mcompar__n0065_inst_lut2_1081.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0065_inst_lut2_1081 (
    .ADR0(DLX_IDinst_reg_out_A[6]),
    .ADR1(VCC),
    .ADR2(\DLX_IDinst_Imm[6] ),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0065_inst_lut2_108)
  );
  defparam DLX_EXinst_Mcompar__n0065_inst_lut2_1091.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0065_inst_lut2_1091 (
    .ADR0(DLX_IDinst_reg_out_A[7]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(\DLX_IDinst_Imm[7] ),
    .O(DLX_EXinst_Mcompar__n0065_inst_lut2_109)
  );
  X_BUF \DLX_IDinst_RegFile_31_11/COUTUSED  (
    .I(\DLX_IDinst_RegFile_31_11/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0065_inst_cy_173)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0065_inst_cy_173_2075 (
    .IA(DLX_IDinst_reg_out_A[7]),
    .IB(DLX_EXinst_Mcompar__n0065_inst_cy_172),
    .SEL(DLX_EXinst_Mcompar__n0065_inst_lut2_109),
    .O(\DLX_IDinst_RegFile_31_11/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_31_11/CYINIT_2076  (
    .I(DLX_EXinst_Mcompar__n0065_inst_cy_171),
    .O(\DLX_IDinst_RegFile_31_11/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0065_inst_cy_174_2077 (
    .IA(DLX_IDinst_reg_out_A[8]),
    .IB(\DLX_EXinst_Mcompar__n0065_inst_cy_175/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0065_inst_lut2_110),
    .O(DLX_EXinst_Mcompar__n0065_inst_cy_174)
  );
  defparam DLX_EXinst_Mcompar__n0065_inst_lut2_1101.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0065_inst_lut2_1101 (
    .ADR0(DLX_IDinst_reg_out_A[8]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(\DLX_IDinst_Imm[8] ),
    .O(DLX_EXinst_Mcompar__n0065_inst_lut2_110)
  );
  defparam DLX_EXinst_Mcompar__n0065_inst_lut2_1111.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0065_inst_lut2_1111 (
    .ADR0(DLX_IDinst_reg_out_A[9]),
    .ADR1(\DLX_IDinst_Imm[9] ),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0065_inst_lut2_111)
  );
  X_BUF \DLX_EXinst_Mcompar__n0065_inst_cy_175/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0065_inst_cy_175/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0065_inst_cy_175)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0065_inst_cy_175_2078 (
    .IA(DLX_IDinst_reg_out_A[9]),
    .IB(DLX_EXinst_Mcompar__n0065_inst_cy_174),
    .SEL(DLX_EXinst_Mcompar__n0065_inst_lut2_111),
    .O(\DLX_EXinst_Mcompar__n0065_inst_cy_175/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0065_inst_cy_175/CYINIT_2079  (
    .I(DLX_EXinst_Mcompar__n0065_inst_cy_173),
    .O(\DLX_EXinst_Mcompar__n0065_inst_cy_175/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0065_inst_cy_176_2080 (
    .IA(DLX_IDinst_reg_out_A[10]),
    .IB(\DLX_IDinst_RegFile_3_30/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0065_inst_lut2_112),
    .O(DLX_EXinst_Mcompar__n0065_inst_cy_176)
  );
  defparam DLX_EXinst_Mcompar__n0065_inst_lut2_1121.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0065_inst_lut2_1121 (
    .ADR0(DLX_IDinst_reg_out_A[10]),
    .ADR1(VCC),
    .ADR2(\DLX_IDinst_Imm[10] ),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0065_inst_lut2_112)
  );
  defparam DLX_EXinst_Mcompar__n0065_inst_lut2_1131.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0065_inst_lut2_1131 (
    .ADR0(DLX_IDinst_reg_out_A[11]),
    .ADR1(\DLX_IDinst_Imm[11] ),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0065_inst_lut2_113)
  );
  X_BUF \DLX_IDinst_RegFile_3_30/COUTUSED  (
    .I(\DLX_IDinst_RegFile_3_30/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0065_inst_cy_177)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0065_inst_cy_177_2081 (
    .IA(DLX_IDinst_reg_out_A[11]),
    .IB(DLX_EXinst_Mcompar__n0065_inst_cy_176),
    .SEL(DLX_EXinst_Mcompar__n0065_inst_lut2_113),
    .O(\DLX_IDinst_RegFile_3_30/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_3_30/CYINIT_2082  (
    .I(DLX_EXinst_Mcompar__n0065_inst_cy_175),
    .O(\DLX_IDinst_RegFile_3_30/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0065_inst_cy_178_2083 (
    .IA(DLX_IDinst_reg_out_A[12]),
    .IB(\DLX_EXinst_Mcompar__n0065_inst_cy_179/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0065_inst_lut2_114),
    .O(DLX_EXinst_Mcompar__n0065_inst_cy_178)
  );
  defparam DLX_EXinst_Mcompar__n0065_inst_lut2_1141.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0065_inst_lut2_1141 (
    .ADR0(DLX_IDinst_reg_out_A[12]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(\DLX_IDinst_Imm[12] ),
    .O(DLX_EXinst_Mcompar__n0065_inst_lut2_114)
  );
  defparam DLX_EXinst_Mcompar__n0065_inst_lut2_1151.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0065_inst_lut2_1151 (
    .ADR0(DLX_IDinst_reg_out_A[13]),
    .ADR1(VCC),
    .ADR2(\DLX_IDinst_Imm[13] ),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0065_inst_lut2_115)
  );
  X_BUF \DLX_EXinst_Mcompar__n0065_inst_cy_179/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0065_inst_cy_179/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0065_inst_cy_179)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0065_inst_cy_179_2084 (
    .IA(DLX_IDinst_reg_out_A[13]),
    .IB(DLX_EXinst_Mcompar__n0065_inst_cy_178),
    .SEL(DLX_EXinst_Mcompar__n0065_inst_lut2_115),
    .O(\DLX_EXinst_Mcompar__n0065_inst_cy_179/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0065_inst_cy_179/CYINIT_2085  (
    .I(DLX_EXinst_Mcompar__n0065_inst_cy_177),
    .O(\DLX_EXinst_Mcompar__n0065_inst_cy_179/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0065_inst_cy_180_2086 (
    .IA(DLX_IDinst_reg_out_A[14]),
    .IB(\DLX_IDinst_RegFile_22_28/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0065_inst_lut2_116),
    .O(DLX_EXinst_Mcompar__n0065_inst_cy_180)
  );
  defparam DLX_EXinst_Mcompar__n0065_inst_lut2_1161.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0065_inst_lut2_1161 (
    .ADR0(DLX_IDinst_reg_out_A[14]),
    .ADR1(\DLX_IDinst_Imm[14] ),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0065_inst_lut2_116)
  );
  defparam DLX_EXinst_Mcompar__n0065_inst_lut2_1171.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0065_inst_lut2_1171 (
    .ADR0(DLX_IDinst_reg_out_A[15]),
    .ADR1(VCC),
    .ADR2(\DLX_IDinst_Imm[15] ),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0065_inst_lut2_117)
  );
  X_BUF \DLX_IDinst_RegFile_22_28/COUTUSED  (
    .I(\DLX_IDinst_RegFile_22_28/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0065_inst_cy_181)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0065_inst_cy_181_2087 (
    .IA(DLX_IDinst_reg_out_A[15]),
    .IB(DLX_EXinst_Mcompar__n0065_inst_cy_180),
    .SEL(DLX_EXinst_Mcompar__n0065_inst_lut2_117),
    .O(\DLX_IDinst_RegFile_22_28/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_22_28/CYINIT_2088  (
    .I(DLX_EXinst_Mcompar__n0065_inst_cy_179),
    .O(\DLX_IDinst_RegFile_22_28/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0065_inst_cy_182_2089 (
    .IA(DLX_IDinst_reg_out_A[16]),
    .IB(\DLX_EXinst_Mcompar__n0065_inst_cy_183/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0065_inst_lut2_118),
    .O(DLX_EXinst_Mcompar__n0065_inst_cy_182)
  );
  defparam DLX_EXinst_Mcompar__n0065_inst_lut2_1181.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0065_inst_lut2_1181 (
    .ADR0(DLX_IDinst_reg_out_A[16]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_Imm_31_1),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0065_inst_lut2_118)
  );
  defparam DLX_EXinst_Mcompar__n0065_inst_lut2_1191.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0065_inst_lut2_1191 (
    .ADR0(DLX_IDinst_reg_out_A[17]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_Imm_31_1),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0065_inst_lut2_119)
  );
  X_BUF \DLX_EXinst_Mcompar__n0065_inst_cy_183/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0065_inst_cy_183/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0065_inst_cy_183)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0065_inst_cy_183_2090 (
    .IA(DLX_IDinst_reg_out_A[17]),
    .IB(DLX_EXinst_Mcompar__n0065_inst_cy_182),
    .SEL(DLX_EXinst_Mcompar__n0065_inst_lut2_119),
    .O(\DLX_EXinst_Mcompar__n0065_inst_cy_183/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0065_inst_cy_183/CYINIT_2091  (
    .I(DLX_EXinst_Mcompar__n0065_inst_cy_181),
    .O(\DLX_EXinst_Mcompar__n0065_inst_cy_183/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0065_inst_cy_184_2092 (
    .IA(DLX_IDinst_reg_out_A[18]),
    .IB(\DLX_IDinst_RegFile_1_8/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0065_inst_lut2_120),
    .O(DLX_EXinst_Mcompar__n0065_inst_cy_184)
  );
  defparam DLX_EXinst_Mcompar__n0065_inst_lut2_1201.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0065_inst_lut2_1201 (
    .ADR0(DLX_IDinst_reg_out_A[18]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_Imm_31_1),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0065_inst_lut2_120)
  );
  defparam DLX_EXinst_Mcompar__n0065_inst_lut2_1211.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0065_inst_lut2_1211 (
    .ADR0(DLX_IDinst_reg_out_A[19]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_Imm_31_1),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0065_inst_lut2_121)
  );
  X_BUF \DLX_IDinst_RegFile_1_8/COUTUSED  (
    .I(\DLX_IDinst_RegFile_1_8/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0065_inst_cy_185)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0065_inst_cy_185_2093 (
    .IA(DLX_IDinst_reg_out_A[19]),
    .IB(DLX_EXinst_Mcompar__n0065_inst_cy_184),
    .SEL(DLX_EXinst_Mcompar__n0065_inst_lut2_121),
    .O(\DLX_IDinst_RegFile_1_8/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_1_8/CYINIT_2094  (
    .I(DLX_EXinst_Mcompar__n0065_inst_cy_183),
    .O(\DLX_IDinst_RegFile_1_8/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0065_inst_cy_186_2095 (
    .IA(DLX_IDinst_reg_out_A[20]),
    .IB(\DLX_EXinst_Mcompar__n0065_inst_cy_187/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0065_inst_lut2_122),
    .O(DLX_EXinst_Mcompar__n0065_inst_cy_186)
  );
  defparam DLX_EXinst_Mcompar__n0065_inst_lut2_1221.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0065_inst_lut2_1221 (
    .ADR0(DLX_IDinst_reg_out_A[20]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_Imm_31_1),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0065_inst_lut2_122)
  );
  defparam DLX_EXinst_Mcompar__n0065_inst_lut2_1231.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0065_inst_lut2_1231 (
    .ADR0(DLX_IDinst_reg_out_A[21]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_Imm_31_1),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0065_inst_lut2_123)
  );
  X_BUF \DLX_EXinst_Mcompar__n0065_inst_cy_187/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0065_inst_cy_187/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0065_inst_cy_187)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0065_inst_cy_187_2096 (
    .IA(DLX_IDinst_reg_out_A[21]),
    .IB(DLX_EXinst_Mcompar__n0065_inst_cy_186),
    .SEL(DLX_EXinst_Mcompar__n0065_inst_lut2_123),
    .O(\DLX_EXinst_Mcompar__n0065_inst_cy_187/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0065_inst_cy_187/CYINIT_2097  (
    .I(DLX_EXinst_Mcompar__n0065_inst_cy_185),
    .O(\DLX_EXinst_Mcompar__n0065_inst_cy_187/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0065_inst_cy_188_2098 (
    .IA(DLX_IDinst_reg_out_A[22]),
    .IB(\DLX_IDinst_RegFile_31_20/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0065_inst_lut2_124),
    .O(DLX_EXinst_Mcompar__n0065_inst_cy_188)
  );
  defparam DLX_EXinst_Mcompar__n0065_inst_lut2_1241.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0065_inst_lut2_1241 (
    .ADR0(DLX_IDinst_reg_out_A[22]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_Imm_31_1),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0065_inst_lut2_124)
  );
  defparam DLX_EXinst_Mcompar__n0065_inst_lut2_1251.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0065_inst_lut2_1251 (
    .ADR0(DLX_IDinst_reg_out_A[23]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_Imm_31_1),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0065_inst_lut2_125)
  );
  X_BUF \DLX_IDinst_RegFile_31_20/COUTUSED  (
    .I(\DLX_IDinst_RegFile_31_20/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0065_inst_cy_189)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0065_inst_cy_189_2099 (
    .IA(DLX_IDinst_reg_out_A[23]),
    .IB(DLX_EXinst_Mcompar__n0065_inst_cy_188),
    .SEL(DLX_EXinst_Mcompar__n0065_inst_lut2_125),
    .O(\DLX_IDinst_RegFile_31_20/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_31_20/CYINIT_2100  (
    .I(DLX_EXinst_Mcompar__n0065_inst_cy_187),
    .O(\DLX_IDinst_RegFile_31_20/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0065_inst_cy_190_2101 (
    .IA(DLX_IDinst_reg_out_A[24]),
    .IB(\DLX_EXinst_Mcompar__n0065_inst_cy_191/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0065_inst_lut2_126),
    .O(DLX_EXinst_Mcompar__n0065_inst_cy_190)
  );
  defparam DLX_EXinst_Mcompar__n0065_inst_lut2_1261.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0065_inst_lut2_1261 (
    .ADR0(DLX_IDinst_reg_out_A[24]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_Imm_31_1),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0065_inst_lut2_126)
  );
  defparam DLX_EXinst_Mcompar__n0065_inst_lut2_1271.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0065_inst_lut2_1271 (
    .ADR0(DLX_IDinst_reg_out_A[25]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_Imm_31_1),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0065_inst_lut2_127)
  );
  X_BUF \DLX_EXinst_Mcompar__n0065_inst_cy_191/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0065_inst_cy_191/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0065_inst_cy_191)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0065_inst_cy_191_2102 (
    .IA(DLX_IDinst_reg_out_A[25]),
    .IB(DLX_EXinst_Mcompar__n0065_inst_cy_190),
    .SEL(DLX_EXinst_Mcompar__n0065_inst_lut2_127),
    .O(\DLX_EXinst_Mcompar__n0065_inst_cy_191/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0065_inst_cy_191/CYINIT_2103  (
    .I(DLX_EXinst_Mcompar__n0065_inst_cy_189),
    .O(\DLX_EXinst_Mcompar__n0065_inst_cy_191/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0065_inst_cy_192_2104 (
    .IA(DLX_IDinst_reg_out_A[26]),
    .IB(\DLX_IDinst_RegFile_24_12/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0065_inst_lut2_128),
    .O(DLX_EXinst_Mcompar__n0065_inst_cy_192)
  );
  defparam DLX_EXinst_Mcompar__n0065_inst_lut2_1281.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0065_inst_lut2_1281 (
    .ADR0(DLX_IDinst_reg_out_A[26]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_Imm_31_1),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0065_inst_lut2_128)
  );
  defparam DLX_EXinst_Mcompar__n0065_inst_lut2_1291.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0065_inst_lut2_1291 (
    .ADR0(DLX_IDinst_reg_out_A[27]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_Imm_31_1),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0065_inst_lut2_129)
  );
  X_BUF \DLX_IDinst_RegFile_24_12/COUTUSED  (
    .I(\DLX_IDinst_RegFile_24_12/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0065_inst_cy_193)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0065_inst_cy_193_2105 (
    .IA(DLX_IDinst_reg_out_A[27]),
    .IB(DLX_EXinst_Mcompar__n0065_inst_cy_192),
    .SEL(DLX_EXinst_Mcompar__n0065_inst_lut2_129),
    .O(\DLX_IDinst_RegFile_24_12/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_24_12/CYINIT_2106  (
    .I(DLX_EXinst_Mcompar__n0065_inst_cy_191),
    .O(\DLX_IDinst_RegFile_24_12/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0065_inst_cy_194_2107 (
    .IA(DLX_IDinst_reg_out_A[28]),
    .IB(\DLX_EXinst_Mcompar__n0065_inst_cy_195/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0065_inst_lut2_130),
    .O(DLX_EXinst_Mcompar__n0065_inst_cy_194)
  );
  defparam DLX_EXinst_Mcompar__n0065_inst_lut2_1301.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0065_inst_lut2_1301 (
    .ADR0(DLX_IDinst_reg_out_A[28]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_Imm_31_1),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0065_inst_lut2_130)
  );
  defparam DLX_EXinst_Mcompar__n0065_inst_lut2_1311.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0065_inst_lut2_1311 (
    .ADR0(DLX_IDinst_reg_out_A[29]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_Imm_31_1),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0065_inst_lut2_131)
  );
  X_BUF \DLX_EXinst_Mcompar__n0065_inst_cy_195/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0065_inst_cy_195/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0065_inst_cy_195)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0065_inst_cy_195_2108 (
    .IA(DLX_IDinst_reg_out_A[29]),
    .IB(DLX_EXinst_Mcompar__n0065_inst_cy_194),
    .SEL(DLX_EXinst_Mcompar__n0065_inst_lut2_131),
    .O(\DLX_EXinst_Mcompar__n0065_inst_cy_195/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0065_inst_cy_195/CYINIT_2109  (
    .I(DLX_EXinst_Mcompar__n0065_inst_cy_193),
    .O(\DLX_EXinst_Mcompar__n0065_inst_cy_195/CYINIT )
  );
  defparam DLX_IDinst_RegFile_29_15_2110.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_29_15_2110 (
    .I(DLX_IDinst_WB_data_eff[15]),
    .CE(DLX_IDinst__n0608),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_29_15)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0065_inst_cy_196_2111 (
    .IA(DLX_IDinst_reg_out_A[30]),
    .IB(\DLX_EXinst_Mcompar__n0065_inst_cy_196/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0065_inst_lut2_132),
    .O(\DLX_EXinst_Mcompar__n0065_inst_cy_196/CYMUXF )
  );
  defparam DLX_EXinst_Mcompar__n0065_inst_lut2_1321.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0065_inst_lut2_1321 (
    .ADR0(DLX_IDinst_reg_out_A[30]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_Imm_31_1),
    .O(DLX_EXinst_Mcompar__n0065_inst_lut2_132)
  );
  X_BUF \DLX_EXinst_Mcompar__n0065_inst_cy_196/XBUSED  (
    .I(\DLX_EXinst_Mcompar__n0065_inst_cy_196/CYMUXF ),
    .O(DLX_EXinst_Mcompar__n0065_inst_cy_196)
  );
  X_BUF \DLX_EXinst_Mcompar__n0065_inst_cy_196/CYINIT_2112  (
    .I(DLX_EXinst_Mcompar__n0065_inst_cy_195),
    .O(\DLX_EXinst_Mcompar__n0065_inst_cy_196/CYINIT )
  );
  X_ONE \DLX_IDinst_RegFile_15_13/LOGIC_ONE_2113  (
    .O(\DLX_IDinst_RegFile_15_13/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_RegFile_15_13/LOGIC_ZERO_2114  (
    .O(\DLX_IDinst_RegFile_15_13/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0029_inst_cy_370_2115 (
    .IA(\DLX_IDinst_RegFile_15_13/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_15_13/LOGIC_ONE ),
    .SEL(vga_top_vga1_Mcompar__n0029_inst_lut1_22),
    .O(vga_top_vga1_Mcompar__n0029_inst_cy_370)
  );
  defparam vga_top_vga1_Mcompar__n0029_inst_lut1_221.INIT = 16'h00FF;
  X_LUT4 vga_top_vga1_Mcompar__n0029_inst_lut1_221 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[4]),
    .O(vga_top_vga1_Mcompar__n0029_inst_lut1_22)
  );
  defparam vga_top_vga1_Mcompar__n0029_inst_lut1_231.INIT = 16'h00FF;
  X_LUT4 vga_top_vga1_Mcompar__n0029_inst_lut1_231 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[4]),
    .O(vga_top_vga1_Mcompar__n0029_inst_lut1_23)
  );
  X_BUF \DLX_IDinst_RegFile_15_13/COUTUSED  (
    .I(\DLX_IDinst_RegFile_15_13/CYMUXG ),
    .O(vga_top_vga1_Mcompar__n0029_inst_cy_371)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0029_inst_cy_371_2116 (
    .IA(\DLX_IDinst_RegFile_15_13/LOGIC_ZERO ),
    .IB(vga_top_vga1_Mcompar__n0029_inst_cy_370),
    .SEL(vga_top_vga1_Mcompar__n0029_inst_lut1_23),
    .O(\DLX_IDinst_RegFile_15_13/CYMUXG )
  );
  X_ONE \vga_top_vga1_Mcompar__n0029_inst_cy_373/LOGIC_ONE_2117  (
    .O(\vga_top_vga1_Mcompar__n0029_inst_cy_373/LOGIC_ONE )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0029_inst_cy_372_2118 (
    .IA(\vga_top_vga1_Mcompar__n0029_inst_cy_373/LOGIC_ONE ),
    .IB(\vga_top_vga1_Mcompar__n0029_inst_cy_373/CYINIT ),
    .SEL(\$SIG_5 ),
    .O(vga_top_vga1_Mcompar__n0029_inst_cy_372)
  );
  defparam \$BEL_5 .INIT = 16'hF0F0;
  X_LUT4 \$BEL_5  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_hcounter[5]),
    .ADR3(VCC),
    .O(\$SIG_5 )
  );
  defparam \$BEL_6 .INIT = 16'hF0F0;
  X_LUT4 \$BEL_6  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_hcounter[5]),
    .ADR3(VCC),
    .O(\$SIG_6 )
  );
  X_BUF \vga_top_vga1_Mcompar__n0029_inst_cy_373/COUTUSED  (
    .I(\vga_top_vga1_Mcompar__n0029_inst_cy_373/CYMUXG ),
    .O(vga_top_vga1_Mcompar__n0029_inst_cy_373)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0029_inst_cy_373_2119 (
    .IA(\vga_top_vga1_Mcompar__n0029_inst_cy_373/LOGIC_ONE ),
    .IB(vga_top_vga1_Mcompar__n0029_inst_cy_372),
    .SEL(\$SIG_6 ),
    .O(\vga_top_vga1_Mcompar__n0029_inst_cy_373/CYMUXG )
  );
  X_BUF \vga_top_vga1_Mcompar__n0029_inst_cy_373/CYINIT_2120  (
    .I(vga_top_vga1_Mcompar__n0029_inst_cy_371),
    .O(\vga_top_vga1_Mcompar__n0029_inst_cy_373/CYINIT )
  );
  X_ZERO \vga_top_vga1_Mcompar__n0029_inst_cy_375/LOGIC_ZERO_2121  (
    .O(\vga_top_vga1_Mcompar__n0029_inst_cy_375/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0029_inst_cy_374_2122 (
    .IA(\vga_top_vga1_Mcompar__n0029_inst_cy_375/LOGIC_ZERO ),
    .IB(\vga_top_vga1_Mcompar__n0029_inst_cy_375/CYINIT ),
    .SEL(vga_top_vga1_Mcompar__n0029_inst_lut4_1104),
    .O(vga_top_vga1_Mcompar__n0029_inst_cy_374)
  );
  defparam vga_top_vga1_Mcompar__n0029_inst_lut4_11041.INIT = 16'h0001;
  X_LUT4 vga_top_vga1_Mcompar__n0029_inst_lut4_11041 (
    .ADR0(vga_top_vga1_hcounter[6]),
    .ADR1(vga_top_vga1_hcounter[8]),
    .ADR2(vga_top_vga1_hcounter[7]),
    .ADR3(vga_top_vga1_hcounter[9]),
    .O(vga_top_vga1_Mcompar__n0029_inst_lut4_1104)
  );
  defparam vga_top_vga1_Mcompar__n0029_inst_lut4_11051.INIT = 16'h0001;
  X_LUT4 vga_top_vga1_Mcompar__n0029_inst_lut4_11051 (
    .ADR0(vga_top_vga1_hcounter[8]),
    .ADR1(vga_top_vga1_hcounter[9]),
    .ADR2(vga_top_vga1_hcounter[6]),
    .ADR3(vga_top_vga1_hcounter[7]),
    .O(vga_top_vga1_Mcompar__n0029_inst_lut4_1105)
  );
  X_BUF \vga_top_vga1_Mcompar__n0029_inst_cy_375/COUTUSED  (
    .I(\vga_top_vga1_Mcompar__n0029_inst_cy_375/CYMUXG ),
    .O(vga_top_vga1_Mcompar__n0029_inst_cy_375)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0029_inst_cy_375_2123 (
    .IA(\vga_top_vga1_Mcompar__n0029_inst_cy_375/LOGIC_ZERO ),
    .IB(vga_top_vga1_Mcompar__n0029_inst_cy_374),
    .SEL(vga_top_vga1_Mcompar__n0029_inst_lut4_1105),
    .O(\vga_top_vga1_Mcompar__n0029_inst_cy_375/CYMUXG )
  );
  X_BUF \vga_top_vga1_Mcompar__n0029_inst_cy_375/CYINIT_2124  (
    .I(vga_top_vga1_Mcompar__n0029_inst_cy_373),
    .O(\vga_top_vga1_Mcompar__n0029_inst_cy_375/CYINIT )
  );
  X_ZERO \DLX_IFinst_IR_curr<10>/LOGIC_ZERO_2125  (
    .O(\DLX_IFinst_IR_curr<10>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0029_inst_cy_376_2126 (
    .IA(\DLX_IFinst_IR_curr<10>/LOGIC_ZERO ),
    .IB(\DLX_IFinst_IR_curr<10>/CYINIT ),
    .SEL(vga_top_vga1_Mcompar__n0029_inst_lut4_1106),
    .O(vga_top_vga1_Mcompar__n0029_inst_cy_376)
  );
  defparam vga_top_vga1_Mcompar__n0029_inst_lut4_11061.INIT = 16'h0001;
  X_LUT4 vga_top_vga1_Mcompar__n0029_inst_lut4_11061 (
    .ADR0(vga_top_vga1_hcounter[10]),
    .ADR1(vga_top_vga1_hcounter[12]),
    .ADR2(vga_top_vga1_hcounter[11]),
    .ADR3(vga_top_vga1_hcounter[13]),
    .O(vga_top_vga1_Mcompar__n0029_inst_lut4_1106)
  );
  defparam vga_top_vga1_Mcompar__n0029_inst_lut2_2751.INIT = 16'h0505;
  X_LUT4 vga_top_vga1_Mcompar__n0029_inst_lut2_2751 (
    .ADR0(vga_top_vga1_hcounter[14]),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_hcounter[15]),
    .ADR3(VCC),
    .O(vga_top_vga1_Mcompar__n0029_inst_lut2_275)
  );
  X_BUF \DLX_IFinst_IR_curr<10>/COUTUSED  (
    .I(\DLX_IFinst_IR_curr<10>/CYMUXG ),
    .O(vga_top_vga1__n0029)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0029_inst_cy_377 (
    .IA(\DLX_IFinst_IR_curr<10>/LOGIC_ZERO ),
    .IB(vga_top_vga1_Mcompar__n0029_inst_cy_376),
    .SEL(vga_top_vga1_Mcompar__n0029_inst_lut2_275),
    .O(\DLX_IFinst_IR_curr<10>/CYMUXG )
  );
  X_BUF \DLX_IFinst_IR_curr<10>/CYINIT_2127  (
    .I(vga_top_vga1_Mcompar__n0029_inst_cy_375),
    .O(\DLX_IFinst_IR_curr<10>/CYINIT )
  );
  X_ONE \vga_top_vga1_Mcompar__n0037_inst_cy_472/LOGIC_ONE_2128  (
    .O(\vga_top_vga1_Mcompar__n0037_inst_cy_472/LOGIC_ONE )
  );
  X_ZERO \vga_top_vga1_Mcompar__n0037_inst_cy_472/LOGIC_ZERO_2129  (
    .O(\vga_top_vga1_Mcompar__n0037_inst_cy_472/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0037_inst_cy_471_2130 (
    .IA(\vga_top_vga1_Mcompar__n0037_inst_cy_472/LOGIC_ZERO ),
    .IB(\vga_top_vga1_Mcompar__n0037_inst_cy_472/LOGIC_ONE ),
    .SEL(vga_top_vga1_Mcompar__n0037_inst_lut2_341),
    .O(vga_top_vga1_Mcompar__n0037_inst_cy_471)
  );
  defparam vga_top_vga1_Mcompar__n0037_inst_lut2_3411.INIT = 16'h8888;
  X_LUT4 vga_top_vga1_Mcompar__n0037_inst_lut2_3411 (
    .ADR0(vga_top_vga1_hcounter[4]),
    .ADR1(vga_top_vga1_hcounter[5]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(vga_top_vga1_Mcompar__n0037_inst_lut2_341)
  );
  defparam vga_top_vga1_Mcompar__n0037_inst_lut2_3421.INIT = 16'hAA00;
  X_LUT4 vga_top_vga1_Mcompar__n0037_inst_lut2_3421 (
    .ADR0(vga_top_vga1_hcounter[5]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[4]),
    .O(vga_top_vga1_Mcompar__n0037_inst_lut2_342)
  );
  X_BUF \vga_top_vga1_Mcompar__n0037_inst_cy_472/COUTUSED  (
    .I(\vga_top_vga1_Mcompar__n0037_inst_cy_472/CYMUXG ),
    .O(vga_top_vga1_Mcompar__n0037_inst_cy_472)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0037_inst_cy_472_2131 (
    .IA(\vga_top_vga1_Mcompar__n0037_inst_cy_472/LOGIC_ZERO ),
    .IB(vga_top_vga1_Mcompar__n0037_inst_cy_471),
    .SEL(vga_top_vga1_Mcompar__n0037_inst_lut2_342),
    .O(\vga_top_vga1_Mcompar__n0037_inst_cy_472/CYMUXG )
  );
  X_ONE \DLX_IDinst_RegFile_30_29/LOGIC_ONE_2132  (
    .O(\DLX_IDinst_RegFile_30_29/LOGIC_ONE )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0037_inst_cy_473_2133 (
    .IA(\DLX_IDinst_RegFile_30_29/LOGIC_ONE ),
    .IB(\DLX_IDinst_RegFile_30_29/CYINIT ),
    .SEL(vga_top_vga1_Mcompar__n0037_inst_lut4_1139),
    .O(vga_top_vga1_Mcompar__n0037_inst_cy_473)
  );
  defparam vga_top_vga1_Mcompar__n0037_inst_lut4_11391.INIT = 16'h0001;
  X_LUT4 vga_top_vga1_Mcompar__n0037_inst_lut4_11391 (
    .ADR0(vga_top_vga1_hcounter[8]),
    .ADR1(vga_top_vga1_hcounter[6]),
    .ADR2(vga_top_vga1_hcounter[7]),
    .ADR3(vga_top_vga1_hcounter[9]),
    .O(vga_top_vga1_Mcompar__n0037_inst_lut4_1139)
  );
  defparam vga_top_vga1_Mcompar__n0037_inst_lut4_11401.INIT = 16'h0001;
  X_LUT4 vga_top_vga1_Mcompar__n0037_inst_lut4_11401 (
    .ADR0(vga_top_vga1_hcounter[8]),
    .ADR1(vga_top_vga1_hcounter[6]),
    .ADR2(vga_top_vga1_hcounter[9]),
    .ADR3(vga_top_vga1_hcounter[7]),
    .O(vga_top_vga1_Mcompar__n0037_inst_lut4_1140)
  );
  X_BUF \DLX_IDinst_RegFile_30_29/COUTUSED  (
    .I(\DLX_IDinst_RegFile_30_29/CYMUXG ),
    .O(vga_top_vga1_Mcompar__n0037_inst_cy_474)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0037_inst_cy_474_2134 (
    .IA(\DLX_IDinst_RegFile_30_29/LOGIC_ONE ),
    .IB(vga_top_vga1_Mcompar__n0037_inst_cy_473),
    .SEL(vga_top_vga1_Mcompar__n0037_inst_lut4_1140),
    .O(\DLX_IDinst_RegFile_30_29/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_30_29/CYINIT_2135  (
    .I(vga_top_vga1_Mcompar__n0037_inst_cy_472),
    .O(\DLX_IDinst_RegFile_30_29/CYINIT )
  );
  X_ONE \vga_top_vga1__n0037/LOGIC_ONE_2136  (
    .O(\vga_top_vga1__n0037/LOGIC_ONE )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0037_inst_cy_475_2137 (
    .IA(\vga_top_vga1__n0037/LOGIC_ONE ),
    .IB(\vga_top_vga1__n0037/CYINIT ),
    .SEL(vga_top_vga1_Mcompar__n0037_inst_lut4_1141),
    .O(vga_top_vga1_Mcompar__n0037_inst_cy_475)
  );
  defparam vga_top_vga1_Mcompar__n0037_inst_lut4_11411.INIT = 16'h0001;
  X_LUT4 vga_top_vga1_Mcompar__n0037_inst_lut4_11411 (
    .ADR0(vga_top_vga1_hcounter[11]),
    .ADR1(vga_top_vga1_hcounter[12]),
    .ADR2(vga_top_vga1_hcounter[13]),
    .ADR3(vga_top_vga1_hcounter[10]),
    .O(vga_top_vga1_Mcompar__n0037_inst_lut4_1141)
  );
  defparam vga_top_vga1_Mcompar__n0037_inst_lut2_3431.INIT = 16'h0033;
  X_LUT4 vga_top_vga1_Mcompar__n0037_inst_lut2_3431 (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_hcounter[15]),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[14]),
    .O(vga_top_vga1_Mcompar__n0037_inst_lut2_343)
  );
  X_BUF \vga_top_vga1__n0037/COUTUSED  (
    .I(\vga_top_vga1__n0037/CYMUXG ),
    .O(vga_top_vga1__n0037)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0037_inst_cy_476 (
    .IA(\vga_top_vga1__n0037/LOGIC_ONE ),
    .IB(vga_top_vga1_Mcompar__n0037_inst_cy_475),
    .SEL(vga_top_vga1_Mcompar__n0037_inst_lut2_343),
    .O(\vga_top_vga1__n0037/CYMUXG )
  );
  X_BUF \vga_top_vga1__n0037/CYINIT_2138  (
    .I(vga_top_vga1_Mcompar__n0037_inst_cy_474),
    .O(\vga_top_vga1__n0037/CYINIT )
  );
  X_ONE \DLX_IDinst_Mcompar__n0368_inst_cy_263/LOGIC_ONE_2139  (
    .O(\DLX_IDinst_Mcompar__n0368_inst_cy_263/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mcompar__n0368_inst_cy_263/LOGIC_ZERO_2140  (
    .O(\DLX_IDinst_Mcompar__n0368_inst_cy_263/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mcompar__n0368_inst_cy_262_2141 (
    .IA(\DLX_IDinst_Mcompar__n0368_inst_cy_263/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mcompar__n0368_inst_cy_263/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mcompar__n0368_inst_lut4_40),
    .O(DLX_IDinst_Mcompar__n0368_inst_cy_262)
  );
  defparam DLX_IDinst_Mcompar__n0368_inst_lut4_401.INIT = 16'h9009;
  X_LUT4 DLX_IDinst_Mcompar__n0368_inst_lut4_401 (
    .ADR0(DLX_MEMinst_reg_dst_out[0]),
    .ADR1(DLX_IDinst_jtarget[16]),
    .ADR2(DLX_MEMinst_reg_dst_out[1]),
    .ADR3(DLX_IDinst_jtarget[17]),
    .O(DLX_IDinst_Mcompar__n0368_inst_lut4_40)
  );
  defparam DLX_IDinst_Mcompar__n0368_inst_lut4_411.INIT = 16'h8241;
  X_LUT4 DLX_IDinst_Mcompar__n0368_inst_lut4_411 (
    .ADR0(DLX_IDinst_jtarget[19]),
    .ADR1(DLX_IDinst_jtarget[18]),
    .ADR2(DLX_MEMinst_reg_dst_out[2]),
    .ADR3(DLX_MEMinst_reg_dst_out[3]),
    .O(DLX_IDinst_Mcompar__n0368_inst_lut4_41)
  );
  X_BUF \DLX_IDinst_Mcompar__n0368_inst_cy_263/COUTUSED  (
    .I(\DLX_IDinst_Mcompar__n0368_inst_cy_263/CYMUXG ),
    .O(DLX_IDinst_Mcompar__n0368_inst_cy_263)
  );
  X_MUX2 DLX_IDinst_Mcompar__n0368_inst_cy_263_2142 (
    .IA(\DLX_IDinst_Mcompar__n0368_inst_cy_263/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mcompar__n0368_inst_cy_262),
    .SEL(DLX_IDinst_Mcompar__n0368_inst_lut4_41),
    .O(\DLX_IDinst_Mcompar__n0368_inst_cy_263/CYMUXG )
  );
  X_ZERO \DLX_EXinst_Mcompar__n0063_inst_cy_135/LOGIC_ZERO_2143  (
    .O(\DLX_EXinst_Mcompar__n0063_inst_cy_135/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_134_2144 (
    .IA(\DLX_IDinst_Imm[0] ),
    .IB(\DLX_EXinst_Mcompar__n0063_inst_cy_135/LOGIC_ZERO ),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_70),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_134)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_701.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_701 (
    .ADR0(\DLX_IDinst_Imm[0] ),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[0]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_70)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_711.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_711 (
    .ADR0(DLX_IDinst_Imm_1_1),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[1]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_71)
  );
  X_BUF \DLX_EXinst_Mcompar__n0063_inst_cy_135/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0063_inst_cy_135/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_135)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_135_2145 (
    .IA(DLX_IDinst_Imm_1_1),
    .IB(DLX_EXinst_Mcompar__n0063_inst_cy_134),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_71),
    .O(\DLX_EXinst_Mcompar__n0063_inst_cy_135/CYMUXG )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_136_2146 (
    .IA(DLX_IDinst_Imm_2_1),
    .IB(\DLX_IDinst_RegFile_15_22/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_72),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_136)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_721.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_721 (
    .ADR0(DLX_IDinst_Imm_2_1),
    .ADR1(DLX_IDinst_reg_out_A[2]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_72)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_731.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_731 (
    .ADR0(DLX_IDinst_Imm_3_1),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[3]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_73)
  );
  X_BUF \DLX_IDinst_RegFile_15_22/COUTUSED  (
    .I(\DLX_IDinst_RegFile_15_22/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_137)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_137_2147 (
    .IA(DLX_IDinst_Imm_3_1),
    .IB(DLX_EXinst_Mcompar__n0063_inst_cy_136),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_73),
    .O(\DLX_IDinst_RegFile_15_22/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_15_22/CYINIT_2148  (
    .I(DLX_EXinst_Mcompar__n0063_inst_cy_135),
    .O(\DLX_IDinst_RegFile_15_22/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_138_2149 (
    .IA(\DLX_IDinst_Imm[4] ),
    .IB(\DLX_EXinst_Mcompar__n0063_inst_cy_139/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_74),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_138)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_741.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_741 (
    .ADR0(\DLX_IDinst_Imm[4] ),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[4]),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_74)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_751.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_751 (
    .ADR0(\DLX_IDinst_Imm[5] ),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[5]),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_75)
  );
  X_BUF \DLX_EXinst_Mcompar__n0063_inst_cy_139/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0063_inst_cy_139/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_139)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_139_2150 (
    .IA(\DLX_IDinst_Imm[5] ),
    .IB(DLX_EXinst_Mcompar__n0063_inst_cy_138),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_75),
    .O(\DLX_EXinst_Mcompar__n0063_inst_cy_139/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0063_inst_cy_139/CYINIT_2151  (
    .I(DLX_EXinst_Mcompar__n0063_inst_cy_137),
    .O(\DLX_EXinst_Mcompar__n0063_inst_cy_139/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_140_2152 (
    .IA(\DLX_IDinst_Imm[6] ),
    .IB(\DLX_IFinst_IR_curr<11>/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_76),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_140)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_761.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_761 (
    .ADR0(\DLX_IDinst_Imm[6] ),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[6]),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_76)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_771.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_771 (
    .ADR0(\DLX_IDinst_Imm[7] ),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[7]),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_77)
  );
  X_BUF \DLX_IFinst_IR_curr<11>/COUTUSED  (
    .I(\DLX_IFinst_IR_curr<11>/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_141)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_141_2153 (
    .IA(\DLX_IDinst_Imm[7] ),
    .IB(DLX_EXinst_Mcompar__n0063_inst_cy_140),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_77),
    .O(\DLX_IFinst_IR_curr<11>/CYMUXG )
  );
  X_BUF \DLX_IFinst_IR_curr<11>/CYINIT_2154  (
    .I(DLX_EXinst_Mcompar__n0063_inst_cy_139),
    .O(\DLX_IFinst_IR_curr<11>/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_142_2155 (
    .IA(\DLX_IDinst_Imm[8] ),
    .IB(\DLX_EXinst_Mcompar__n0063_inst_cy_143/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_78),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_142)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_781.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_781 (
    .ADR0(\DLX_IDinst_Imm[8] ),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[8]),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_78)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_791.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_791 (
    .ADR0(\DLX_IDinst_Imm[9] ),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[9]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_79)
  );
  X_BUF \DLX_EXinst_Mcompar__n0063_inst_cy_143/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0063_inst_cy_143/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_143)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_143_2156 (
    .IA(\DLX_IDinst_Imm[9] ),
    .IB(DLX_EXinst_Mcompar__n0063_inst_cy_142),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_79),
    .O(\DLX_EXinst_Mcompar__n0063_inst_cy_143/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0063_inst_cy_143/CYINIT_2157  (
    .I(DLX_EXinst_Mcompar__n0063_inst_cy_141),
    .O(\DLX_EXinst_Mcompar__n0063_inst_cy_143/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_144_2158 (
    .IA(\DLX_IDinst_Imm[10] ),
    .IB(\DLX_IDinst_RegFile_23_14/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_80),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_144)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_801.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_801 (
    .ADR0(\DLX_IDinst_Imm[10] ),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[10]),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_80)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_811.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_811 (
    .ADR0(\DLX_IDinst_Imm[11] ),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[11]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_81)
  );
  X_BUF \DLX_IDinst_RegFile_23_14/COUTUSED  (
    .I(\DLX_IDinst_RegFile_23_14/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_145)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_145_2159 (
    .IA(\DLX_IDinst_Imm[11] ),
    .IB(DLX_EXinst_Mcompar__n0063_inst_cy_144),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_81),
    .O(\DLX_IDinst_RegFile_23_14/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_23_14/CYINIT_2160  (
    .I(DLX_EXinst_Mcompar__n0063_inst_cy_143),
    .O(\DLX_IDinst_RegFile_23_14/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_146_2161 (
    .IA(\DLX_IDinst_Imm[12] ),
    .IB(\DLX_EXinst_Mcompar__n0063_inst_cy_147/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_82),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_146)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_821.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_821 (
    .ADR0(\DLX_IDinst_Imm[12] ),
    .ADR1(DLX_IDinst_reg_out_A[12]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_82)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_831.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_831 (
    .ADR0(\DLX_IDinst_Imm[13] ),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[13]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_83)
  );
  X_BUF \DLX_EXinst_Mcompar__n0063_inst_cy_147/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0063_inst_cy_147/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_147)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_147_2162 (
    .IA(\DLX_IDinst_Imm[13] ),
    .IB(DLX_EXinst_Mcompar__n0063_inst_cy_146),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_83),
    .O(\DLX_EXinst_Mcompar__n0063_inst_cy_147/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0063_inst_cy_147/CYINIT_2163  (
    .I(DLX_EXinst_Mcompar__n0063_inst_cy_145),
    .O(\DLX_EXinst_Mcompar__n0063_inst_cy_147/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_148_2164 (
    .IA(\DLX_IDinst_Imm[14] ),
    .IB(\DLX_IDinst_RegFile_26_3/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_84),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_148)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_841.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_841 (
    .ADR0(\DLX_IDinst_Imm[14] ),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[14]),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_84)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_851.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_851 (
    .ADR0(\DLX_IDinst_Imm[15] ),
    .ADR1(DLX_IDinst_reg_out_A[15]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_85)
  );
  X_BUF \DLX_IDinst_RegFile_26_3/COUTUSED  (
    .I(\DLX_IDinst_RegFile_26_3/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_149)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_149_2165 (
    .IA(\DLX_IDinst_Imm[15] ),
    .IB(DLX_EXinst_Mcompar__n0063_inst_cy_148),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_85),
    .O(\DLX_IDinst_RegFile_26_3/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_26_3/CYINIT_2166  (
    .I(DLX_EXinst_Mcompar__n0063_inst_cy_147),
    .O(\DLX_IDinst_RegFile_26_3/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_150_2167 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(\DLX_EXinst_Mcompar__n0063_inst_cy_151/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_86),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_150)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_861.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_861 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[16]),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_86)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_871.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_871 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(DLX_IDinst_reg_out_A[17]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_87)
  );
  X_BUF \DLX_EXinst_Mcompar__n0063_inst_cy_151/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0063_inst_cy_151/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_151)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_151_2168 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(DLX_EXinst_Mcompar__n0063_inst_cy_150),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_87),
    .O(\DLX_EXinst_Mcompar__n0063_inst_cy_151/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0063_inst_cy_151/CYINIT_2169  (
    .I(DLX_EXinst_Mcompar__n0063_inst_cy_149),
    .O(\DLX_EXinst_Mcompar__n0063_inst_cy_151/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_152_2170 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(\DLX_IDinst_RegFile_15_23/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_88),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_152)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_881.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_881 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[18]),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_88)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_891.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_891 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[19]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_89)
  );
  X_BUF \DLX_IDinst_RegFile_15_23/COUTUSED  (
    .I(\DLX_IDinst_RegFile_15_23/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_153)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_153_2171 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(DLX_EXinst_Mcompar__n0063_inst_cy_152),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_89),
    .O(\DLX_IDinst_RegFile_15_23/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_15_23/CYINIT_2172  (
    .I(DLX_EXinst_Mcompar__n0063_inst_cy_151),
    .O(\DLX_IDinst_RegFile_15_23/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_154_2173 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(\DLX_EXinst_Mcompar__n0063_inst_cy_155/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_90),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_154)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_901.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_901 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(DLX_IDinst_reg_out_A[20]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_90)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_911.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_911 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[21]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_91)
  );
  X_BUF \DLX_EXinst_Mcompar__n0063_inst_cy_155/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0063_inst_cy_155/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_155)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_155_2174 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(DLX_EXinst_Mcompar__n0063_inst_cy_154),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_91),
    .O(\DLX_EXinst_Mcompar__n0063_inst_cy_155/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0063_inst_cy_155/CYINIT_2175  (
    .I(DLX_EXinst_Mcompar__n0063_inst_cy_153),
    .O(\DLX_EXinst_Mcompar__n0063_inst_cy_155/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_156_2176 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(\DLX_IFinst_IR_curr<20>/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_92),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_156)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_921.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_921 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[22]),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_92)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_931.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_931 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[23]),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_93)
  );
  X_BUF \DLX_IFinst_IR_curr<20>/COUTUSED  (
    .I(\DLX_IFinst_IR_curr<20>/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_157)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_157_2177 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(DLX_EXinst_Mcompar__n0063_inst_cy_156),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_93),
    .O(\DLX_IFinst_IR_curr<20>/CYMUXG )
  );
  X_BUF \DLX_IFinst_IR_curr<20>/CYINIT_2178  (
    .I(DLX_EXinst_Mcompar__n0063_inst_cy_155),
    .O(\DLX_IFinst_IR_curr<20>/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_158_2179 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(\DLX_EXinst_Mcompar__n0063_inst_cy_159/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_94),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_158)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_941.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_941 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(DLX_IDinst_reg_out_A[24]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_94)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_951.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_951 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(DLX_IDinst_reg_out_A[25]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_95)
  );
  X_BUF \DLX_EXinst_Mcompar__n0063_inst_cy_159/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0063_inst_cy_159/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_159)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_159_2180 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(DLX_EXinst_Mcompar__n0063_inst_cy_158),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_95),
    .O(\DLX_EXinst_Mcompar__n0063_inst_cy_159/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0063_inst_cy_159/CYINIT_2181  (
    .I(DLX_EXinst_Mcompar__n0063_inst_cy_157),
    .O(\DLX_EXinst_Mcompar__n0063_inst_cy_159/CYINIT )
  );
  defparam DLX_IDinst_RegFile_29_23_2182.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_29_23_2182 (
    .I(DLX_IDinst_WB_data_eff[23]),
    .CE(DLX_IDinst__n0608),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_29_23)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_160_2183 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(\DLX_IDinst_RegFile_31_23/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_96),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_160)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_961.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_961 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[26]),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_96)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_971.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_971 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[27]),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_97)
  );
  X_BUF \DLX_IDinst_RegFile_31_23/COUTUSED  (
    .I(\DLX_IDinst_RegFile_31_23/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_161)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_161_2184 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(DLX_EXinst_Mcompar__n0063_inst_cy_160),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_97),
    .O(\DLX_IDinst_RegFile_31_23/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_31_23/CYINIT_2185  (
    .I(DLX_EXinst_Mcompar__n0063_inst_cy_159),
    .O(\DLX_IDinst_RegFile_31_23/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_162_2186 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(\DLX_EXinst_Mcompar__n0063_inst_cy_163/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_98),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_162)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_981.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_981 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(DLX_IDinst_reg_out_A[28]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_98)
  );
  defparam DLX_EXinst_Mcompar__n0063_inst_lut2_991.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0063_inst_lut2_991 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(DLX_IDinst_reg_out_A[29]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0063_inst_lut2_99)
  );
  X_BUF \DLX_EXinst_Mcompar__n0063_inst_cy_163/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0063_inst_cy_163/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0063_inst_cy_163)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0063_inst_cy_163_2187 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(DLX_EXinst_Mcompar__n0063_inst_cy_162),
    .SEL(DLX_EXinst_Mcompar__n0063_inst_lut2_99),
    .O(\DLX_EXinst_Mcompar__n0063_inst_cy_163/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0063_inst_cy_163/CYINIT_2188  (
    .I(DLX_EXinst_Mcompar__n0063_inst_cy_161),
    .O(\DLX_EXinst_Mcompar__n0063_inst_cy_163/CYINIT )
  );
  X_ONE \DLX_IDinst_RegFile_31_29/LOGIC_ONE_2189  (
    .O(\DLX_IDinst_RegFile_31_29/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_RegFile_31_29/LOGIC_ZERO_2190  (
    .O(\DLX_IDinst_RegFile_31_29/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0030_inst_cy_354_2191 (
    .IA(\DLX_IDinst_RegFile_31_29/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_31_29/LOGIC_ONE ),
    .SEL(vga_top_vga1_Mcompar__n0030_inst_lut4_1101),
    .O(vga_top_vga1_Mcompar__n0030_inst_cy_354)
  );
  defparam vga_top_vga1_Mcompar__n0030_inst_lut4_11011.INIT = 16'h8000;
  X_LUT4 vga_top_vga1_Mcompar__n0030_inst_lut4_11011 (
    .ADR0(vga_top_vga1_hcounter[1]),
    .ADR1(vga_top_vga1_hcounter[3]),
    .ADR2(vga_top_vga1_hcounter[0]),
    .ADR3(vga_top_vga1_hcounter[2]),
    .O(vga_top_vga1_Mcompar__n0030_inst_lut4_1101)
  );
  defparam vga_top_vga1_Mcompar__n0030_inst_lut4_11021.INIT = 16'h8000;
  X_LUT4 vga_top_vga1_Mcompar__n0030_inst_lut4_11021 (
    .ADR0(vga_top_vga1_hcounter[2]),
    .ADR1(vga_top_vga1_hcounter[3]),
    .ADR2(vga_top_vga1_hcounter[1]),
    .ADR3(vga_top_vga1_hcounter[0]),
    .O(vga_top_vga1_Mcompar__n0030_inst_lut4_1102)
  );
  X_BUF \DLX_IDinst_RegFile_31_29/COUTUSED  (
    .I(\DLX_IDinst_RegFile_31_29/CYMUXG ),
    .O(vga_top_vga1_Mcompar__n0030_inst_cy_355)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0030_inst_cy_355_2192 (
    .IA(\DLX_IDinst_RegFile_31_29/LOGIC_ZERO ),
    .IB(vga_top_vga1_Mcompar__n0030_inst_cy_354),
    .SEL(vga_top_vga1_Mcompar__n0030_inst_lut4_1102),
    .O(\DLX_IDinst_RegFile_31_29/CYMUXG )
  );
  X_ONE \vga_top_vga1_Mcompar__n0030_inst_cy_357/LOGIC_ONE_2193  (
    .O(\vga_top_vga1_Mcompar__n0030_inst_cy_357/LOGIC_ONE )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0030_inst_cy_356_2194 (
    .IA(\vga_top_vga1_Mcompar__n0030_inst_cy_357/LOGIC_ONE ),
    .IB(\vga_top_vga1_Mcompar__n0030_inst_cy_357/CYINIT ),
    .SEL(vga_top_vga1_Mcompar__n0030_inst_lut1_10),
    .O(vga_top_vga1_Mcompar__n0030_inst_cy_356)
  );
  defparam vga_top_vga1_Mcompar__n0030_inst_lut1_101.INIT = 16'h0F0F;
  X_LUT4 vga_top_vga1_Mcompar__n0030_inst_lut1_101 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_hcounter[4]),
    .ADR3(VCC),
    .O(vga_top_vga1_Mcompar__n0030_inst_lut1_10)
  );
  defparam vga_top_vga1_Mcompar__n0030_inst_lut1_111.INIT = 16'h5555;
  X_LUT4 vga_top_vga1_Mcompar__n0030_inst_lut1_111 (
    .ADR0(vga_top_vga1_hcounter[4]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(vga_top_vga1_Mcompar__n0030_inst_lut1_11)
  );
  X_BUF \vga_top_vga1_Mcompar__n0030_inst_cy_357/COUTUSED  (
    .I(\vga_top_vga1_Mcompar__n0030_inst_cy_357/CYMUXG ),
    .O(vga_top_vga1_Mcompar__n0030_inst_cy_357)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0030_inst_cy_357_2195 (
    .IA(\vga_top_vga1_Mcompar__n0030_inst_cy_357/LOGIC_ONE ),
    .IB(vga_top_vga1_Mcompar__n0030_inst_cy_356),
    .SEL(vga_top_vga1_Mcompar__n0030_inst_lut1_11),
    .O(\vga_top_vga1_Mcompar__n0030_inst_cy_357/CYMUXG )
  );
  X_BUF \vga_top_vga1_Mcompar__n0030_inst_cy_357/CYINIT_2196  (
    .I(vga_top_vga1_Mcompar__n0030_inst_cy_355),
    .O(\vga_top_vga1_Mcompar__n0030_inst_cy_357/CYINIT )
  );
  X_ZERO \vga_top_vga1_Mcompar__n0030_inst_cy_359/LOGIC_ZERO_2197  (
    .O(\vga_top_vga1_Mcompar__n0030_inst_cy_359/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0030_inst_cy_358_2198 (
    .IA(\vga_top_vga1_Mcompar__n0030_inst_cy_359/LOGIC_ZERO ),
    .IB(\vga_top_vga1_Mcompar__n0030_inst_cy_359/CYINIT ),
    .SEL(\$SIG_7 ),
    .O(vga_top_vga1_Mcompar__n0030_inst_cy_358)
  );
  defparam \$BEL_7 .INIT = 16'hFF00;
  X_LUT4 \$BEL_7  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[5]),
    .O(\$SIG_7 )
  );
  defparam \$BEL_8 .INIT = 16'hCCCC;
  X_LUT4 \$BEL_8  (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_hcounter[5]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\$SIG_8 )
  );
  X_BUF \vga_top_vga1_Mcompar__n0030_inst_cy_359/COUTUSED  (
    .I(\vga_top_vga1_Mcompar__n0030_inst_cy_359/CYMUXG ),
    .O(vga_top_vga1_Mcompar__n0030_inst_cy_359)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0030_inst_cy_359_2199 (
    .IA(\vga_top_vga1_Mcompar__n0030_inst_cy_359/LOGIC_ZERO ),
    .IB(vga_top_vga1_Mcompar__n0030_inst_cy_358),
    .SEL(\$SIG_8 ),
    .O(\vga_top_vga1_Mcompar__n0030_inst_cy_359/CYMUXG )
  );
  X_BUF \vga_top_vga1_Mcompar__n0030_inst_cy_359/CYINIT_2200  (
    .I(vga_top_vga1_Mcompar__n0030_inst_cy_357),
    .O(\vga_top_vga1_Mcompar__n0030_inst_cy_359/CYINIT )
  );
  X_ONE \DLX_IDinst_RegFile_31_31/LOGIC_ONE_2201  (
    .O(\DLX_IDinst_RegFile_31_31/LOGIC_ONE )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0030_inst_cy_360_2202 (
    .IA(\DLX_IDinst_RegFile_31_31/LOGIC_ONE ),
    .IB(\DLX_IDinst_RegFile_31_31/CYINIT ),
    .SEL(vga_top_vga1_Mcompar__n0030_inst_lut1_14),
    .O(vga_top_vga1_Mcompar__n0030_inst_cy_360)
  );
  defparam vga_top_vga1_Mcompar__n0030_inst_lut1_141.INIT = 16'h0F0F;
  X_LUT4 vga_top_vga1_Mcompar__n0030_inst_lut1_141 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_hcounter[6]),
    .ADR3(VCC),
    .O(vga_top_vga1_Mcompar__n0030_inst_lut1_14)
  );
  defparam vga_top_vga1_Mcompar__n0030_inst_lut1_151.INIT = 16'h00FF;
  X_LUT4 vga_top_vga1_Mcompar__n0030_inst_lut1_151 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[6]),
    .O(vga_top_vga1_Mcompar__n0030_inst_lut1_15)
  );
  X_BUF \DLX_IDinst_RegFile_31_31/COUTUSED  (
    .I(\DLX_IDinst_RegFile_31_31/CYMUXG ),
    .O(vga_top_vga1_Mcompar__n0030_inst_cy_361)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0030_inst_cy_361_2203 (
    .IA(\DLX_IDinst_RegFile_31_31/LOGIC_ONE ),
    .IB(vga_top_vga1_Mcompar__n0030_inst_cy_360),
    .SEL(vga_top_vga1_Mcompar__n0030_inst_lut1_15),
    .O(\DLX_IDinst_RegFile_31_31/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_31_31/CYINIT_2204  (
    .I(vga_top_vga1_Mcompar__n0030_inst_cy_359),
    .O(\DLX_IDinst_RegFile_31_31/CYINIT )
  );
  X_ZERO \vga_top_vga1_Mcompar__n0030_inst_cy_363/LOGIC_ZERO_2205  (
    .O(\vga_top_vga1_Mcompar__n0030_inst_cy_363/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0030_inst_cy_362_2206 (
    .IA(\vga_top_vga1_Mcompar__n0030_inst_cy_363/LOGIC_ZERO ),
    .IB(\vga_top_vga1_Mcompar__n0030_inst_cy_363/CYINIT ),
    .SEL(\$SIG_9 ),
    .O(vga_top_vga1_Mcompar__n0030_inst_cy_362)
  );
  defparam \$BEL_9 .INIT = 16'hF0F0;
  X_LUT4 \$BEL_9  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_hcounter[7]),
    .ADR3(VCC),
    .O(\$SIG_9 )
  );
  defparam \$BEL_10 .INIT = 16'hCCCC;
  X_LUT4 \$BEL_10  (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_hcounter[7]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\$SIG_10 )
  );
  X_BUF \vga_top_vga1_Mcompar__n0030_inst_cy_363/COUTUSED  (
    .I(\vga_top_vga1_Mcompar__n0030_inst_cy_363/CYMUXG ),
    .O(vga_top_vga1_Mcompar__n0030_inst_cy_363)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0030_inst_cy_363_2207 (
    .IA(\vga_top_vga1_Mcompar__n0030_inst_cy_363/LOGIC_ZERO ),
    .IB(vga_top_vga1_Mcompar__n0030_inst_cy_362),
    .SEL(\$SIG_10 ),
    .O(\vga_top_vga1_Mcompar__n0030_inst_cy_363/CYMUXG )
  );
  X_BUF \vga_top_vga1_Mcompar__n0030_inst_cy_363/CYINIT_2208  (
    .I(vga_top_vga1_Mcompar__n0030_inst_cy_361),
    .O(\vga_top_vga1_Mcompar__n0030_inst_cy_363/CYINIT )
  );
  X_ONE \vga_top_vga1_Mcompar__n0030_inst_cy_365/LOGIC_ONE_2209  (
    .O(\vga_top_vga1_Mcompar__n0030_inst_cy_365/LOGIC_ONE )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0030_inst_cy_364_2210 (
    .IA(\vga_top_vga1_Mcompar__n0030_inst_cy_365/LOGIC_ONE ),
    .IB(\vga_top_vga1_Mcompar__n0030_inst_cy_365/CYINIT ),
    .SEL(vga_top_vga1_Mcompar__n0030_inst_lut1_18),
    .O(vga_top_vga1_Mcompar__n0030_inst_cy_364)
  );
  defparam vga_top_vga1_Mcompar__n0030_inst_lut1_181.INIT = 16'h00FF;
  X_LUT4 vga_top_vga1_Mcompar__n0030_inst_lut1_181 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[8]),
    .O(vga_top_vga1_Mcompar__n0030_inst_lut1_18)
  );
  defparam vga_top_vga1_Mcompar__n0030_inst_lut1_191.INIT = 16'h00FF;
  X_LUT4 vga_top_vga1_Mcompar__n0030_inst_lut1_191 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[8]),
    .O(vga_top_vga1_Mcompar__n0030_inst_lut1_19)
  );
  X_BUF \vga_top_vga1_Mcompar__n0030_inst_cy_365/COUTUSED  (
    .I(\vga_top_vga1_Mcompar__n0030_inst_cy_365/CYMUXG ),
    .O(vga_top_vga1_Mcompar__n0030_inst_cy_365)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0030_inst_cy_365_2211 (
    .IA(\vga_top_vga1_Mcompar__n0030_inst_cy_365/LOGIC_ONE ),
    .IB(vga_top_vga1_Mcompar__n0030_inst_cy_364),
    .SEL(vga_top_vga1_Mcompar__n0030_inst_lut1_19),
    .O(\vga_top_vga1_Mcompar__n0030_inst_cy_365/CYMUXG )
  );
  X_BUF \vga_top_vga1_Mcompar__n0030_inst_cy_365/CYINIT_2212  (
    .I(vga_top_vga1_Mcompar__n0030_inst_cy_363),
    .O(\vga_top_vga1_Mcompar__n0030_inst_cy_365/CYINIT )
  );
  X_ZERO \vga_top_vga1_Mcompar__n0030_inst_cy_367/LOGIC_ZERO_2213  (
    .O(\vga_top_vga1_Mcompar__n0030_inst_cy_367/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0030_inst_cy_366_2214 (
    .IA(\vga_top_vga1_Mcompar__n0030_inst_cy_367/LOGIC_ZERO ),
    .IB(\vga_top_vga1_Mcompar__n0030_inst_cy_367/CYINIT ),
    .SEL(\$SIG_11 ),
    .O(vga_top_vga1_Mcompar__n0030_inst_cy_366)
  );
  defparam \$BEL_11 .INIT = 16'hFF00;
  X_LUT4 \$BEL_11  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[9]),
    .O(\$SIG_11 )
  );
  defparam \$BEL_12 .INIT = 16'hCCCC;
  X_LUT4 \$BEL_12  (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_hcounter[9]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\$SIG_12 )
  );
  X_BUF \vga_top_vga1_Mcompar__n0030_inst_cy_367/COUTUSED  (
    .I(\vga_top_vga1_Mcompar__n0030_inst_cy_367/CYMUXG ),
    .O(vga_top_vga1_Mcompar__n0030_inst_cy_367)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0030_inst_cy_367_2215 (
    .IA(\vga_top_vga1_Mcompar__n0030_inst_cy_367/LOGIC_ZERO ),
    .IB(vga_top_vga1_Mcompar__n0030_inst_cy_366),
    .SEL(\$SIG_12 ),
    .O(\vga_top_vga1_Mcompar__n0030_inst_cy_367/CYMUXG )
  );
  X_BUF \vga_top_vga1_Mcompar__n0030_inst_cy_367/CYINIT_2216  (
    .I(vga_top_vga1_Mcompar__n0030_inst_cy_365),
    .O(\vga_top_vga1_Mcompar__n0030_inst_cy_367/CYINIT )
  );
  X_ONE \DLX_IFinst_IR_curr<12>/LOGIC_ONE_2217  (
    .O(\DLX_IFinst_IR_curr<12>/LOGIC_ONE )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0030_inst_cy_368_2218 (
    .IA(\DLX_IFinst_IR_curr<12>/LOGIC_ONE ),
    .IB(\DLX_IFinst_IR_curr<12>/CYINIT ),
    .SEL(vga_top_vga1_Mcompar__n0030_inst_lut4_1103),
    .O(vga_top_vga1_Mcompar__n0030_inst_cy_368)
  );
  defparam vga_top_vga1_Mcompar__n0030_inst_lut4_11031.INIT = 16'h0001;
  X_LUT4 vga_top_vga1_Mcompar__n0030_inst_lut4_11031 (
    .ADR0(vga_top_vga1_hcounter[10]),
    .ADR1(vga_top_vga1_hcounter[13]),
    .ADR2(vga_top_vga1_hcounter[12]),
    .ADR3(vga_top_vga1_hcounter[11]),
    .O(vga_top_vga1_Mcompar__n0030_inst_lut4_1103)
  );
  defparam vga_top_vga1_Mcompar__n0030_inst_lut2_2741.INIT = 16'h0505;
  X_LUT4 vga_top_vga1_Mcompar__n0030_inst_lut2_2741 (
    .ADR0(vga_top_vga1_hcounter[14]),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_hcounter[15]),
    .ADR3(VCC),
    .O(vga_top_vga1_Mcompar__n0030_inst_lut2_274)
  );
  X_BUF \DLX_IFinst_IR_curr<12>/COUTUSED  (
    .I(\DLX_IFinst_IR_curr<12>/CYMUXG ),
    .O(vga_top_vga1__n0030)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0030_inst_cy_369 (
    .IA(\DLX_IFinst_IR_curr<12>/LOGIC_ONE ),
    .IB(vga_top_vga1_Mcompar__n0030_inst_cy_368),
    .SEL(vga_top_vga1_Mcompar__n0030_inst_lut2_274),
    .O(\DLX_IFinst_IR_curr<12>/CYMUXG )
  );
  X_BUF \DLX_IFinst_IR_curr<12>/CYINIT_2219  (
    .I(vga_top_vga1_Mcompar__n0030_inst_cy_367),
    .O(\DLX_IFinst_IR_curr<12>/CYINIT )
  );
  X_ZERO \DLX_EXinst_Mcompar__n0089_inst_cy_135/LOGIC_ZERO_2220  (
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_135/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_134_2221 (
    .IA(DLX_IDinst_reg_out_B[0]),
    .IB(\DLX_EXinst_Mcompar__n0089_inst_cy_135/LOGIC_ZERO ),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_70),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_134)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_701.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_701 (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(DLX_IDinst_reg_out_A[0]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_70)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_711.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_711 (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[1]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_71)
  );
  X_BUF \DLX_EXinst_Mcompar__n0089_inst_cy_135/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0089_inst_cy_135/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_135)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_135_2222 (
    .IA(DLX_IDinst_reg_out_B[1]),
    .IB(DLX_EXinst_Mcompar__n0089_inst_cy_134),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_71),
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_135/CYMUXG )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_136_2223 (
    .IA(DLX_IDinst_reg_out_B_2_1),
    .IB(\DLX_IDinst_RegFile_23_16/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_72),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_136)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_721.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_721 (
    .ADR0(DLX_IDinst_reg_out_B_2_1),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[2]),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_72)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_731.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_731 (
    .ADR0(DLX_IDinst_reg_out_B_3_1),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[3]),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_73)
  );
  X_BUF \DLX_IDinst_RegFile_23_16/COUTUSED  (
    .I(\DLX_IDinst_RegFile_23_16/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_137)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_137_2224 (
    .IA(DLX_IDinst_reg_out_B_3_1),
    .IB(DLX_EXinst_Mcompar__n0089_inst_cy_136),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_73),
    .O(\DLX_IDinst_RegFile_23_16/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_23_16/CYINIT_2225  (
    .I(DLX_EXinst_Mcompar__n0089_inst_cy_135),
    .O(\DLX_IDinst_RegFile_23_16/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_138_2226 (
    .IA(DLX_IDinst_reg_out_B[4]),
    .IB(\DLX_EXinst_Mcompar__n0089_inst_cy_139/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_74),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_138)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_741.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_741 (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(DLX_IDinst_reg_out_A[4]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_74)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_751.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_751 (
    .ADR0(DLX_IDinst_reg_out_B[5]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[5]),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_75)
  );
  X_BUF \DLX_EXinst_Mcompar__n0089_inst_cy_139/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0089_inst_cy_139/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_139)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_139_2227 (
    .IA(DLX_IDinst_reg_out_B[5]),
    .IB(DLX_EXinst_Mcompar__n0089_inst_cy_138),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_75),
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_139/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0089_inst_cy_139/CYINIT_2228  (
    .I(DLX_EXinst_Mcompar__n0089_inst_cy_137),
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_139/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_140_2229 (
    .IA(DLX_IDinst_reg_out_B[6]),
    .IB(\vga_top_vga1_clockcounter_FFd2/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_76),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_140)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_761.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_761 (
    .ADR0(DLX_IDinst_reg_out_B[6]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[6]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_76)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_771.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_771 (
    .ADR0(DLX_IDinst_reg_out_B[7]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[7]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_77)
  );
  X_BUF \vga_top_vga1_clockcounter_FFd2/COUTUSED  (
    .I(\vga_top_vga1_clockcounter_FFd2/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_141)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_141_2230 (
    .IA(DLX_IDinst_reg_out_B[7]),
    .IB(DLX_EXinst_Mcompar__n0089_inst_cy_140),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_77),
    .O(\vga_top_vga1_clockcounter_FFd2/CYMUXG )
  );
  X_BUF \vga_top_vga1_clockcounter_FFd2/CYINIT_2231  (
    .I(DLX_EXinst_Mcompar__n0089_inst_cy_139),
    .O(\vga_top_vga1_clockcounter_FFd2/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_142_2232 (
    .IA(DLX_IDinst_reg_out_B[8]),
    .IB(\DLX_EXinst_Mcompar__n0089_inst_cy_143/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_78),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_142)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_781.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_781 (
    .ADR0(DLX_IDinst_reg_out_B[8]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[8]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_78)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_791.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_791 (
    .ADR0(DLX_IDinst_reg_out_B[9]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[9]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_79)
  );
  X_BUF \DLX_EXinst_Mcompar__n0089_inst_cy_143/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0089_inst_cy_143/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_143)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_143_2233 (
    .IA(DLX_IDinst_reg_out_B[9]),
    .IB(DLX_EXinst_Mcompar__n0089_inst_cy_142),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_79),
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_143/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0089_inst_cy_143/CYINIT_2234  (
    .I(DLX_EXinst_Mcompar__n0089_inst_cy_141),
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_143/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_144_2235 (
    .IA(DLX_IDinst_reg_out_B[10]),
    .IB(\DLX_IDinst_RegFile_6_26/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_80),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_144)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_801.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_801 (
    .ADR0(DLX_IDinst_reg_out_B[10]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[10]),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_80)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_811.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_811 (
    .ADR0(DLX_IDinst_reg_out_B[11]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[11]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_81)
  );
  X_BUF \DLX_IDinst_RegFile_6_26/COUTUSED  (
    .I(\DLX_IDinst_RegFile_6_26/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_145)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_145_2236 (
    .IA(DLX_IDinst_reg_out_B[11]),
    .IB(DLX_EXinst_Mcompar__n0089_inst_cy_144),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_81),
    .O(\DLX_IDinst_RegFile_6_26/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_6_26/CYINIT_2237  (
    .I(DLX_EXinst_Mcompar__n0089_inst_cy_143),
    .O(\DLX_IDinst_RegFile_6_26/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_146_2238 (
    .IA(DLX_IDinst_reg_out_B[12]),
    .IB(\DLX_EXinst_Mcompar__n0089_inst_cy_147/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_82),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_146)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_821.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_821 (
    .ADR0(DLX_IDinst_reg_out_B[12]),
    .ADR1(DLX_IDinst_reg_out_A[12]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_82)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_831.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_831 (
    .ADR0(DLX_IDinst_reg_out_B[13]),
    .ADR1(DLX_IDinst_reg_out_A[13]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_83)
  );
  X_BUF \DLX_EXinst_Mcompar__n0089_inst_cy_147/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0089_inst_cy_147/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_147)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_147_2239 (
    .IA(DLX_IDinst_reg_out_B[13]),
    .IB(DLX_EXinst_Mcompar__n0089_inst_cy_146),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_83),
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_147/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0089_inst_cy_147/CYINIT_2240  (
    .I(DLX_EXinst_Mcompar__n0089_inst_cy_145),
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_147/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_148_2241 (
    .IA(DLX_IDinst_reg_out_B[14]),
    .IB(\DLX_IFinst_IR_curr<21>/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_84),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_148)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_841.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_841 (
    .ADR0(DLX_IDinst_reg_out_B[14]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[14]),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_84)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_851.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_851 (
    .ADR0(DLX_IDinst_reg_out_B[15]),
    .ADR1(DLX_IDinst_reg_out_A[15]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_85)
  );
  X_BUF \DLX_IFinst_IR_curr<21>/COUTUSED  (
    .I(\DLX_IFinst_IR_curr<21>/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_149)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_149_2242 (
    .IA(DLX_IDinst_reg_out_B[15]),
    .IB(DLX_EXinst_Mcompar__n0089_inst_cy_148),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_85),
    .O(\DLX_IFinst_IR_curr<21>/CYMUXG )
  );
  X_BUF \DLX_IFinst_IR_curr<21>/CYINIT_2243  (
    .I(DLX_EXinst_Mcompar__n0089_inst_cy_147),
    .O(\DLX_IFinst_IR_curr<21>/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_150_2244 (
    .IA(DLX_IDinst_reg_out_B[16]),
    .IB(\DLX_EXinst_Mcompar__n0089_inst_cy_151/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_86),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_150)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_861.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_861 (
    .ADR0(DLX_IDinst_reg_out_B[16]),
    .ADR1(DLX_IDinst_reg_out_A[16]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_86)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_871.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_871 (
    .ADR0(DLX_IDinst_reg_out_B[17]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[17]),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_87)
  );
  X_BUF \DLX_EXinst_Mcompar__n0089_inst_cy_151/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0089_inst_cy_151/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_151)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_151_2245 (
    .IA(DLX_IDinst_reg_out_B[17]),
    .IB(DLX_EXinst_Mcompar__n0089_inst_cy_150),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_87),
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_151/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0089_inst_cy_151/CYINIT_2246  (
    .I(DLX_EXinst_Mcompar__n0089_inst_cy_149),
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_151/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_152_2247 (
    .IA(DLX_IDinst_reg_out_B[18]),
    .IB(\DLX_IDinst_RegFile_7_11/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_88),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_152)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_881.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_881 (
    .ADR0(DLX_IDinst_reg_out_B[18]),
    .ADR1(DLX_IDinst_reg_out_A[18]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_88)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_891.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_891 (
    .ADR0(DLX_IDinst_reg_out_B[19]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[19]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_89)
  );
  X_BUF \DLX_IDinst_RegFile_7_11/COUTUSED  (
    .I(\DLX_IDinst_RegFile_7_11/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_153)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_153_2248 (
    .IA(DLX_IDinst_reg_out_B[19]),
    .IB(DLX_EXinst_Mcompar__n0089_inst_cy_152),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_89),
    .O(\DLX_IDinst_RegFile_7_11/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_7_11/CYINIT_2249  (
    .I(DLX_EXinst_Mcompar__n0089_inst_cy_151),
    .O(\DLX_IDinst_RegFile_7_11/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_154_2250 (
    .IA(DLX_IDinst_reg_out_B[20]),
    .IB(\DLX_EXinst_Mcompar__n0089_inst_cy_155/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_90),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_154)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_901.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_901 (
    .ADR0(DLX_IDinst_reg_out_B[20]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[20]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_90)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_911.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_911 (
    .ADR0(DLX_IDinst_reg_out_B[21]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[21]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_91)
  );
  X_BUF \DLX_EXinst_Mcompar__n0089_inst_cy_155/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0089_inst_cy_155/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_155)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_155_2251 (
    .IA(DLX_IDinst_reg_out_B[21]),
    .IB(DLX_EXinst_Mcompar__n0089_inst_cy_154),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_91),
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_155/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0089_inst_cy_155/CYINIT_2252  (
    .I(DLX_EXinst_Mcompar__n0089_inst_cy_153),
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_155/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_156_2253 (
    .IA(DLX_IDinst_reg_out_B[22]),
    .IB(\DLX_IDinst_RegFile_3_23/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_92),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_156)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_921.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_921 (
    .ADR0(DLX_IDinst_reg_out_B[22]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[22]),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_92)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_931.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_931 (
    .ADR0(DLX_IDinst_reg_out_B[23]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[23]),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_93)
  );
  X_BUF \DLX_IDinst_RegFile_3_23/COUTUSED  (
    .I(\DLX_IDinst_RegFile_3_23/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_157)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_157_2254 (
    .IA(DLX_IDinst_reg_out_B[23]),
    .IB(DLX_EXinst_Mcompar__n0089_inst_cy_156),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_93),
    .O(\DLX_IDinst_RegFile_3_23/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_3_23/CYINIT_2255  (
    .I(DLX_EXinst_Mcompar__n0089_inst_cy_155),
    .O(\DLX_IDinst_RegFile_3_23/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_158_2256 (
    .IA(DLX_IDinst_reg_out_B[24]),
    .IB(\DLX_EXinst_Mcompar__n0089_inst_cy_159/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_94),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_158)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_941.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_941 (
    .ADR0(DLX_IDinst_reg_out_B[24]),
    .ADR1(DLX_IDinst_reg_out_A[24]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_94)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_951.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_951 (
    .ADR0(DLX_IDinst_reg_out_B[25]),
    .ADR1(DLX_IDinst_reg_out_A[25]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_95)
  );
  X_BUF \DLX_EXinst_Mcompar__n0089_inst_cy_159/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0089_inst_cy_159/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_159)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_159_2257 (
    .IA(DLX_IDinst_reg_out_B[25]),
    .IB(DLX_EXinst_Mcompar__n0089_inst_cy_158),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_95),
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_159/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0089_inst_cy_159/CYINIT_2258  (
    .I(DLX_EXinst_Mcompar__n0089_inst_cy_157),
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_159/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_160_2259 (
    .IA(DLX_IDinst_reg_out_B[26]),
    .IB(\DLX_IDinst_RegFile_31_17/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_96),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_160)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_961.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_961 (
    .ADR0(DLX_IDinst_reg_out_B[26]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[26]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_96)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_971.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_971 (
    .ADR0(DLX_IDinst_reg_out_B[27]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[27]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_97)
  );
  X_BUF \DLX_IDinst_RegFile_31_17/COUTUSED  (
    .I(\DLX_IDinst_RegFile_31_17/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_161)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_161_2260 (
    .IA(DLX_IDinst_reg_out_B[27]),
    .IB(DLX_EXinst_Mcompar__n0089_inst_cy_160),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_97),
    .O(\DLX_IDinst_RegFile_31_17/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_31_17/CYINIT_2261  (
    .I(DLX_EXinst_Mcompar__n0089_inst_cy_159),
    .O(\DLX_IDinst_RegFile_31_17/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_162_2262 (
    .IA(DLX_IDinst_reg_out_B[28]),
    .IB(\DLX_EXinst_Mcompar__n0089_inst_cy_163/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_98),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_162)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_981.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_981 (
    .ADR0(DLX_IDinst_reg_out_B[28]),
    .ADR1(DLX_IDinst_reg_out_A[28]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_98)
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_991.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_991 (
    .ADR0(DLX_IDinst_reg_out_B[29]),
    .ADR1(DLX_IDinst_reg_out_A[29]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_99)
  );
  X_BUF \DLX_EXinst_Mcompar__n0089_inst_cy_163/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0089_inst_cy_163/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_163)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_163_2263 (
    .IA(DLX_IDinst_reg_out_B[29]),
    .IB(DLX_EXinst_Mcompar__n0089_inst_cy_162),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_99),
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_163/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0089_inst_cy_163/CYINIT_2264  (
    .I(DLX_EXinst_Mcompar__n0089_inst_cy_161),
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_163/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0089_inst_cy_164_2265 (
    .IA(DLX_IDinst_reg_out_B[30]),
    .IB(\DLX_EXinst_Mcompar__n0089_inst_cy_164/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0089_inst_lut2_100),
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_164/CYMUXF )
  );
  defparam DLX_EXinst_Mcompar__n0089_inst_lut2_1001.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0089_inst_lut2_1001 (
    .ADR0(DLX_IDinst_reg_out_B[30]),
    .ADR1(DLX_IDinst_reg_out_A[30]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0089_inst_lut2_100)
  );
  X_BUF \DLX_EXinst_Mcompar__n0089_inst_cy_164/XBUSED  (
    .I(\DLX_EXinst_Mcompar__n0089_inst_cy_164/CYMUXF ),
    .O(DLX_EXinst_Mcompar__n0089_inst_cy_164)
  );
  X_BUF \DLX_EXinst_Mcompar__n0089_inst_cy_164/CYINIT_2266  (
    .I(DLX_EXinst_Mcompar__n0089_inst_cy_163),
    .O(\DLX_EXinst_Mcompar__n0089_inst_cy_164/CYINIT )
  );
  X_ONE \DLX_IDinst_Mcompar__n0104_inst_cy_263/LOGIC_ONE_2267  (
    .O(\DLX_IDinst_Mcompar__n0104_inst_cy_263/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mcompar__n0104_inst_cy_263/LOGIC_ZERO_2268  (
    .O(\DLX_IDinst_Mcompar__n0104_inst_cy_263/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mcompar__n0104_inst_cy_262_2269 (
    .IA(\DLX_IDinst_Mcompar__n0104_inst_cy_263/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mcompar__n0104_inst_cy_263/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mcompar__n0104_inst_lut4_40),
    .O(DLX_IDinst_Mcompar__n0104_inst_cy_262)
  );
  defparam DLX_IDinst_Mcompar__n0104_inst_lut4_401.INIT = 16'h9009;
  X_LUT4 DLX_IDinst_Mcompar__n0104_inst_lut4_401 (
    .ADR0(DLX_EXinst_reg_dst_out[1]),
    .ADR1(DLX_IDinst_jtarget[22]),
    .ADR2(DLX_EXinst_reg_dst_out[0]),
    .ADR3(DLX_IDinst_jtarget[21]),
    .O(DLX_IDinst_Mcompar__n0104_inst_lut4_40)
  );
  defparam DLX_IDinst_Mcompar__n0104_inst_lut4_411.INIT = 16'h9009;
  X_LUT4 DLX_IDinst_Mcompar__n0104_inst_lut4_411 (
    .ADR0(DLX_IDinst_jtarget[23]),
    .ADR1(DLX_EXinst_reg_dst_out[2]),
    .ADR2(DLX_IDinst_jtarget[24]),
    .ADR3(DLX_EXinst_reg_dst_out[3]),
    .O(DLX_IDinst_Mcompar__n0104_inst_lut4_41)
  );
  X_BUF \DLX_IDinst_Mcompar__n0104_inst_cy_263/COUTUSED  (
    .I(\DLX_IDinst_Mcompar__n0104_inst_cy_263/CYMUXG ),
    .O(DLX_IDinst_Mcompar__n0104_inst_cy_263)
  );
  X_MUX2 DLX_IDinst_Mcompar__n0104_inst_cy_263_2270 (
    .IA(\DLX_IDinst_Mcompar__n0104_inst_cy_263/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mcompar__n0104_inst_cy_262),
    .SEL(DLX_IDinst_Mcompar__n0104_inst_lut4_41),
    .O(\DLX_IDinst_Mcompar__n0104_inst_cy_263/CYMUXG )
  );
  X_ZERO \DLX_IDinst__n0104/LOGIC_ZERO_2271  (
    .O(\DLX_IDinst__n0104/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mcompar__n0104_inst_cy_264 (
    .IA(\DLX_IDinst__n0104/LOGIC_ZERO ),
    .IB(\DLX_IDinst__n0104/CYINIT ),
    .SEL(DLX_IDinst_Mcompar__n0104_inst_lut4_42),
    .O(\DLX_IDinst__n0104/CYMUXF )
  );
  defparam DLX_IDinst_Mcompar__n0104_inst_lut4_421.INIT = 16'h99A5;
  X_LUT4 DLX_IDinst_Mcompar__n0104_inst_lut4_421 (
    .ADR0(DLX_EXinst_reg_dst_out[4]),
    .ADR1(DLX_IFinst_IR_latched[25]),
    .ADR2(DLX_IDinst_current_IR[25]),
    .ADR3(DLX_EXinst__n0144),
    .O(DLX_IDinst_Mcompar__n0104_inst_lut4_42)
  );
  X_BUF \DLX_IDinst__n0104/XBUSED  (
    .I(\DLX_IDinst__n0104/CYMUXF ),
    .O(DLX_IDinst__n0104)
  );
  X_BUF \DLX_IDinst__n0104/CYINIT_2272  (
    .I(DLX_IDinst_Mcompar__n0104_inst_cy_263),
    .O(\DLX_IDinst__n0104/CYINIT )
  );
  X_ZERO \DLX_EXinst_Mcompar__n0061_inst_cy_119/LOGIC_ZERO_2273  (
    .O(\DLX_EXinst_Mcompar__n0061_inst_cy_119/LOGIC_ZERO )
  );
  X_ONE \DLX_EXinst_Mcompar__n0061_inst_cy_119/LOGIC_ONE_2274  (
    .O(\DLX_EXinst_Mcompar__n0061_inst_cy_119/LOGIC_ONE )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0061_inst_cy_118_2275 (
    .IA(\DLX_EXinst_Mcompar__n0061_inst_cy_119/LOGIC_ONE ),
    .IB(\DLX_EXinst_Mcompar__n0061_inst_cy_119/LOGIC_ZERO ),
    .SEL(DLX_EXinst_Mcompar__n0061_inst_lut4_16),
    .O(DLX_EXinst_Mcompar__n0061_inst_cy_118)
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_lut4_161.INIT = 16'h8421;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_lut4_161 (
    .ADR0(DLX_IDinst_reg_out_A[1]),
    .ADR1(\DLX_IDinst_Imm[0] ),
    .ADR2(DLX_IDinst_Imm_1_1),
    .ADR3(DLX_IDinst_reg_out_A[0]),
    .O(DLX_EXinst_Mcompar__n0061_inst_lut4_16)
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_lut4_171.INIT = 16'h9009;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_lut4_171 (
    .ADR0(DLX_IDinst_Imm_3_1),
    .ADR1(DLX_IDinst_reg_out_A[3]),
    .ADR2(DLX_IDinst_Imm_2_1),
    .ADR3(DLX_IDinst_reg_out_A[2]),
    .O(DLX_EXinst_Mcompar__n0061_inst_lut4_17)
  );
  X_BUF \DLX_EXinst_Mcompar__n0061_inst_cy_119/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0061_inst_cy_119/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0061_inst_cy_119)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0061_inst_cy_119_2276 (
    .IA(\DLX_EXinst_Mcompar__n0061_inst_cy_119/LOGIC_ONE ),
    .IB(DLX_EXinst_Mcompar__n0061_inst_cy_118),
    .SEL(DLX_EXinst_Mcompar__n0061_inst_lut4_17),
    .O(\DLX_EXinst_Mcompar__n0061_inst_cy_119/CYMUXG )
  );
  X_ONE \DLX_EXinst_Mcompar__n0061_inst_cy_121/LOGIC_ONE_2277  (
    .O(\DLX_EXinst_Mcompar__n0061_inst_cy_121/LOGIC_ONE )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0061_inst_cy_120_2278 (
    .IA(\DLX_EXinst_Mcompar__n0061_inst_cy_121/LOGIC_ONE ),
    .IB(\DLX_EXinst_Mcompar__n0061_inst_cy_121/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0061_inst_lut4_18),
    .O(DLX_EXinst_Mcompar__n0061_inst_cy_120)
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_lut4_181.INIT = 16'h8241;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_lut4_181 (
    .ADR0(DLX_IDinst_reg_out_A[5]),
    .ADR1(\DLX_IDinst_Imm[4] ),
    .ADR2(DLX_IDinst_reg_out_A[4]),
    .ADR3(\DLX_IDinst_Imm[5] ),
    .O(DLX_EXinst_Mcompar__n0061_inst_lut4_18)
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_lut4_191.INIT = 16'h8421;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_lut4_191 (
    .ADR0(DLX_IDinst_reg_out_A[7]),
    .ADR1(\DLX_IDinst_Imm[6] ),
    .ADR2(\DLX_IDinst_Imm[7] ),
    .ADR3(DLX_IDinst_reg_out_A[6]),
    .O(DLX_EXinst_Mcompar__n0061_inst_lut4_19)
  );
  X_BUF \DLX_EXinst_Mcompar__n0061_inst_cy_121/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0061_inst_cy_121/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0061_inst_cy_121)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0061_inst_cy_121_2279 (
    .IA(\DLX_EXinst_Mcompar__n0061_inst_cy_121/LOGIC_ONE ),
    .IB(DLX_EXinst_Mcompar__n0061_inst_cy_120),
    .SEL(DLX_EXinst_Mcompar__n0061_inst_lut4_19),
    .O(\DLX_EXinst_Mcompar__n0061_inst_cy_121/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0061_inst_cy_121/CYINIT_2280  (
    .I(DLX_EXinst_Mcompar__n0061_inst_cy_119),
    .O(\DLX_EXinst_Mcompar__n0061_inst_cy_121/CYINIT )
  );
  X_ONE \DLX_EXinst_Mcompar__n0061_inst_cy_123/LOGIC_ONE_2281  (
    .O(\DLX_EXinst_Mcompar__n0061_inst_cy_123/LOGIC_ONE )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0061_inst_cy_122_2282 (
    .IA(\DLX_EXinst_Mcompar__n0061_inst_cy_123/LOGIC_ONE ),
    .IB(\DLX_EXinst_Mcompar__n0061_inst_cy_123/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0061_inst_lut4_20),
    .O(DLX_EXinst_Mcompar__n0061_inst_cy_122)
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_lut4_201.INIT = 16'h8241;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_lut4_201 (
    .ADR0(DLX_IDinst_reg_out_A[9]),
    .ADR1(DLX_IDinst_reg_out_A[8]),
    .ADR2(\DLX_IDinst_Imm[8] ),
    .ADR3(\DLX_IDinst_Imm[9] ),
    .O(DLX_EXinst_Mcompar__n0061_inst_lut4_20)
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_lut4_211.INIT = 16'h9009;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_lut4_211 (
    .ADR0(\DLX_IDinst_Imm[10] ),
    .ADR1(DLX_IDinst_reg_out_A[10]),
    .ADR2(DLX_IDinst_reg_out_A[11]),
    .ADR3(\DLX_IDinst_Imm[11] ),
    .O(DLX_EXinst_Mcompar__n0061_inst_lut4_21)
  );
  X_BUF \DLX_EXinst_Mcompar__n0061_inst_cy_123/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0061_inst_cy_123/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0061_inst_cy_123)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0061_inst_cy_123_2283 (
    .IA(\DLX_EXinst_Mcompar__n0061_inst_cy_123/LOGIC_ONE ),
    .IB(DLX_EXinst_Mcompar__n0061_inst_cy_122),
    .SEL(DLX_EXinst_Mcompar__n0061_inst_lut4_21),
    .O(\DLX_EXinst_Mcompar__n0061_inst_cy_123/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0061_inst_cy_123/CYINIT_2284  (
    .I(DLX_EXinst_Mcompar__n0061_inst_cy_121),
    .O(\DLX_EXinst_Mcompar__n0061_inst_cy_123/CYINIT )
  );
  X_ONE \DLX_MEMinst_opcode_of_WB<0>/LOGIC_ONE_2285  (
    .O(\DLX_MEMinst_opcode_of_WB<0>/LOGIC_ONE )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0061_inst_cy_124_2286 (
    .IA(\DLX_MEMinst_opcode_of_WB<0>/LOGIC_ONE ),
    .IB(\DLX_MEMinst_opcode_of_WB<0>/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0061_inst_lut4_22),
    .O(DLX_EXinst_Mcompar__n0061_inst_cy_124)
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_lut4_221.INIT = 16'h9009;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_lut4_221 (
    .ADR0(DLX_IDinst_reg_out_A[13]),
    .ADR1(\DLX_IDinst_Imm[13] ),
    .ADR2(\DLX_IDinst_Imm[12] ),
    .ADR3(DLX_IDinst_reg_out_A[12]),
    .O(DLX_EXinst_Mcompar__n0061_inst_lut4_22)
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_lut4_231.INIT = 16'h9009;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_lut4_231 (
    .ADR0(\DLX_IDinst_Imm[15] ),
    .ADR1(DLX_IDinst_reg_out_A[15]),
    .ADR2(\DLX_IDinst_Imm[14] ),
    .ADR3(DLX_IDinst_reg_out_A[14]),
    .O(DLX_EXinst_Mcompar__n0061_inst_lut4_23)
  );
  X_BUF \DLX_MEMinst_opcode_of_WB<0>/COUTUSED  (
    .I(\DLX_MEMinst_opcode_of_WB<0>/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0061_inst_cy_125)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0061_inst_cy_125_2287 (
    .IA(\DLX_MEMinst_opcode_of_WB<0>/LOGIC_ONE ),
    .IB(DLX_EXinst_Mcompar__n0061_inst_cy_124),
    .SEL(DLX_EXinst_Mcompar__n0061_inst_lut4_23),
    .O(\DLX_MEMinst_opcode_of_WB<0>/CYMUXG )
  );
  X_BUF \DLX_MEMinst_opcode_of_WB<0>/CYINIT_2288  (
    .I(DLX_EXinst_Mcompar__n0061_inst_cy_123),
    .O(\DLX_MEMinst_opcode_of_WB<0>/CYINIT )
  );
  defparam DLX_IDinst_RegFile_29_31_2289.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_29_31_2289 (
    .I(DLX_IDinst_WB_data_eff[31]),
    .CE(DLX_IDinst__n0608),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_29_31)
  );
  X_ONE \DLX_EXinst_Mcompar__n0061_inst_cy_127/LOGIC_ONE_2290  (
    .O(\DLX_EXinst_Mcompar__n0061_inst_cy_127/LOGIC_ONE )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0061_inst_cy_126_2291 (
    .IA(\DLX_EXinst_Mcompar__n0061_inst_cy_127/LOGIC_ONE ),
    .IB(\DLX_EXinst_Mcompar__n0061_inst_cy_127/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0061_inst_lut4_24),
    .O(DLX_EXinst_Mcompar__n0061_inst_cy_126)
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_lut4_241.INIT = 16'h8421;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_lut4_241 (
    .ADR0(\DLX_IDinst_Imm[31] ),
    .ADR1(DLX_IDinst_reg_out_A[16]),
    .ADR2(DLX_IDinst_reg_out_A[17]),
    .ADR3(DLX_IDinst_Imm_31_1),
    .O(DLX_EXinst_Mcompar__n0061_inst_lut4_24)
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_lut4_251.INIT = 16'h8811;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_lut4_251 (
    .ADR0(DLX_IDinst_reg_out_A[18]),
    .ADR1(DLX_IDinst_reg_out_A[19]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_Imm_31_1),
    .O(DLX_EXinst_Mcompar__n0061_inst_lut4_25)
  );
  X_BUF \DLX_EXinst_Mcompar__n0061_inst_cy_127/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0061_inst_cy_127/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0061_inst_cy_127)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0061_inst_cy_127_2292 (
    .IA(\DLX_EXinst_Mcompar__n0061_inst_cy_127/LOGIC_ONE ),
    .IB(DLX_EXinst_Mcompar__n0061_inst_cy_126),
    .SEL(DLX_EXinst_Mcompar__n0061_inst_lut4_25),
    .O(\DLX_EXinst_Mcompar__n0061_inst_cy_127/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0061_inst_cy_127/CYINIT_2293  (
    .I(DLX_EXinst_Mcompar__n0061_inst_cy_125),
    .O(\DLX_EXinst_Mcompar__n0061_inst_cy_127/CYINIT )
  );
  X_ONE \DLX_IDinst_RegFile_23_26/LOGIC_ONE_2294  (
    .O(\DLX_IDinst_RegFile_23_26/LOGIC_ONE )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0061_inst_cy_128_2295 (
    .IA(\DLX_IDinst_RegFile_23_26/LOGIC_ONE ),
    .IB(\DLX_IDinst_RegFile_23_26/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0061_inst_lut4_26),
    .O(DLX_EXinst_Mcompar__n0061_inst_cy_128)
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_lut4_261.INIT = 16'h8811;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_lut4_261 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(DLX_IDinst_reg_out_A[21]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[20]),
    .O(DLX_EXinst_Mcompar__n0061_inst_lut4_26)
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_lut4_271.INIT = 16'h8811;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_lut4_271 (
    .ADR0(DLX_IDinst_reg_out_A[22]),
    .ADR1(DLX_IDinst_Imm_31_1),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[23]),
    .O(DLX_EXinst_Mcompar__n0061_inst_lut4_27)
  );
  X_BUF \DLX_IDinst_RegFile_23_26/COUTUSED  (
    .I(\DLX_IDinst_RegFile_23_26/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0061_inst_cy_129)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0061_inst_cy_129_2296 (
    .IA(\DLX_IDinst_RegFile_23_26/LOGIC_ONE ),
    .IB(DLX_EXinst_Mcompar__n0061_inst_cy_128),
    .SEL(DLX_EXinst_Mcompar__n0061_inst_lut4_27),
    .O(\DLX_IDinst_RegFile_23_26/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_23_26/CYINIT_2297  (
    .I(DLX_EXinst_Mcompar__n0061_inst_cy_127),
    .O(\DLX_IDinst_RegFile_23_26/CYINIT )
  );
  X_ONE \DLX_EXinst_Mcompar__n0061_inst_cy_131/LOGIC_ONE_2298  (
    .O(\DLX_EXinst_Mcompar__n0061_inst_cy_131/LOGIC_ONE )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0061_inst_cy_130_2299 (
    .IA(\DLX_EXinst_Mcompar__n0061_inst_cy_131/LOGIC_ONE ),
    .IB(\DLX_EXinst_Mcompar__n0061_inst_cy_131/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0061_inst_lut4_28),
    .O(DLX_EXinst_Mcompar__n0061_inst_cy_130)
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_lut4_281.INIT = 16'hC003;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_lut4_281 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_reg_out_A[24]),
    .ADR2(DLX_IDinst_Imm_31_1),
    .ADR3(DLX_IDinst_reg_out_A[25]),
    .O(DLX_EXinst_Mcompar__n0061_inst_lut4_28)
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_lut4_291.INIT = 16'h8181;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_lut4_291 (
    .ADR0(DLX_IDinst_reg_out_A[27]),
    .ADR1(DLX_IDinst_reg_out_A[26]),
    .ADR2(DLX_IDinst_Imm_31_1),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0061_inst_lut4_29)
  );
  X_BUF \DLX_EXinst_Mcompar__n0061_inst_cy_131/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0061_inst_cy_131/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0061_inst_cy_131)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0061_inst_cy_131_2300 (
    .IA(\DLX_EXinst_Mcompar__n0061_inst_cy_131/LOGIC_ONE ),
    .IB(DLX_EXinst_Mcompar__n0061_inst_cy_130),
    .SEL(DLX_EXinst_Mcompar__n0061_inst_lut4_29),
    .O(\DLX_EXinst_Mcompar__n0061_inst_cy_131/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0061_inst_cy_131/CYINIT_2301  (
    .I(DLX_EXinst_Mcompar__n0061_inst_cy_129),
    .O(\DLX_EXinst_Mcompar__n0061_inst_cy_131/CYINIT )
  );
  X_ONE \DLX_IDinst_RegFile_16_13/LOGIC_ONE_2302  (
    .O(\DLX_IDinst_RegFile_16_13/LOGIC_ONE )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0061_inst_cy_132_2303 (
    .IA(\DLX_IDinst_RegFile_16_13/LOGIC_ONE ),
    .IB(\DLX_IDinst_RegFile_16_13/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0061_inst_lut4_30),
    .O(DLX_EXinst_Mcompar__n0061_inst_cy_132)
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_lut4_301.INIT = 16'hA005;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_lut4_301 (
    .ADR0(DLX_IDinst_reg_out_A[29]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_Imm_31_1),
    .ADR3(DLX_IDinst_reg_out_A[28]),
    .O(DLX_EXinst_Mcompar__n0061_inst_lut4_30)
  );
  defparam DLX_EXinst_Mcompar__n0061_inst_lut4_311.INIT = 16'hA005;
  X_LUT4 DLX_EXinst_Mcompar__n0061_inst_lut4_311 (
    .ADR0(DLX_IDinst_reg_out_A[30]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_Imm_31_1),
    .ADR3(DLX_IDinst_reg_out_A[31]),
    .O(DLX_EXinst_Mcompar__n0061_inst_lut4_31)
  );
  X_BUF \DLX_IDinst_RegFile_16_13/COUTUSED  (
    .I(\DLX_IDinst_RegFile_16_13/CYMUXG ),
    .O(DLX_EXinst__n0061)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0061_inst_cy_133 (
    .IA(\DLX_IDinst_RegFile_16_13/LOGIC_ONE ),
    .IB(DLX_EXinst_Mcompar__n0061_inst_cy_132),
    .SEL(DLX_EXinst_Mcompar__n0061_inst_lut4_31),
    .O(\DLX_IDinst_RegFile_16_13/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_16_13/CYINIT_2304  (
    .I(DLX_EXinst_Mcompar__n0061_inst_cy_131),
    .O(\DLX_IDinst_RegFile_16_13/CYINIT )
  );
  X_ONE \DLX_IDinst_Mmux__COND_5_inst_cy_593/LOGIC_ONE_2305  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_593/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_5_inst_cy_593/LOGIC_ZERO_2306  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_593/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_592_2307 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_593/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_5_inst_cy_593/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_667),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_592)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6671.INIT = 16'hFB3B;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6671 (
    .ADR0(DLX_IDinst_RegFile_0_5),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_571),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR3(DLX_IDinst_RegFile_1_5),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_667)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6681.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6681 (
    .ADR0(DLX_IDinst_RegFile_2_5),
    .ADR1(DLX_IDinst_RegFile_3_5),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_572),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_668)
  );
  X_BUF \DLX_IDinst_Mmux__COND_5_inst_cy_593/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_5_inst_cy_593/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_593)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_593_2308 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_593/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_592),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_668),
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_593/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mmux__COND_5_inst_cy_513/LOGIC_ONE_2309  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_513/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_5_inst_cy_513/LOGIC_ZERO_2310  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_513/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_512_2311 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_513/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_5_inst_cy_513/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_587),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_512)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_5871.INIT = 16'hAFCF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_5871 (
    .ADR0(DLX_IDinst_RegFile_1_0),
    .ADR1(DLX_IDinst_RegFile_0_0),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_571),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_587)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_5881.INIT = 16'hFB73;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_5881 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_572),
    .ADR2(DLX_IDinst_RegFile_2_0),
    .ADR3(DLX_IDinst_RegFile_3_0),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_588)
  );
  X_BUF \DLX_IDinst_Mmux__COND_5_inst_cy_513/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_5_inst_cy_513/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_513)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_513_2312 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_513/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_512),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_588),
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_513/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mmux__COND_5_inst_cy_609/LOGIC_ONE_2313  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_609/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_5_inst_cy_609/LOGIC_ZERO_2314  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_609/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_608_2315 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_609/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_5_inst_cy_609/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_683),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_608)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6831.INIT = 16'hFB73;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6831 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_571),
    .ADR2(DLX_IDinst_RegFile_0_6),
    .ADR3(DLX_IDinst_RegFile_1_6),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_683)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6841.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6841 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_572),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR2(DLX_IDinst_RegFile_2_6),
    .ADR3(DLX_IDinst_RegFile_3_6),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_684)
  );
  X_BUF \DLX_IDinst_Mmux__COND_5_inst_cy_609/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_5_inst_cy_609/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_609)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_609_2316 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_609/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_608),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_684),
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_609/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mmux__COND_5_inst_cy_529/LOGIC_ONE_2317  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_529/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_5_inst_cy_529/LOGIC_ZERO_2318  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_529/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_528_2319 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_529/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_5_inst_cy_529/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_603),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_528)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6031.INIT = 16'hF7D5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6031 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_571),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR2(DLX_IDinst_RegFile_1_1),
    .ADR3(DLX_IDinst_RegFile_0_1),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_603)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6041.INIT = 16'hCFAF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6041 (
    .ADR0(DLX_IDinst_RegFile_2_1),
    .ADR1(DLX_IDinst_RegFile_3_1),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_572),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_604)
  );
  X_BUF \DLX_IDinst_Mmux__COND_5_inst_cy_529/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_5_inst_cy_529/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_529)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_529_2320 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_529/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_528),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_604),
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_529/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mmux__COND_5_inst_cy_689/LOGIC_ONE_2321  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_689/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_5_inst_cy_689/LOGIC_ZERO_2322  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_689/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_688_2323 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_689/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_5_inst_cy_689/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_763),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_688)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7631.INIT = 16'hF7D5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7631 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_571),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR2(DLX_IDinst_RegFile_1_11),
    .ADR3(DLX_IDinst_RegFile_0_11),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_763)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7641.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7641 (
    .ADR0(DLX_IDinst_RegFile_2_11),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_572),
    .ADR3(DLX_IDinst_RegFile_3_11),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_764)
  );
  X_BUF \DLX_IDinst_Mmux__COND_5_inst_cy_689/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_5_inst_cy_689/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_689)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_689_2324 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_689/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_688),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_764),
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_689/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mmux__COND_5_inst_cy_705/LOGIC_ONE_2325  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_705/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_5_inst_cy_705/LOGIC_ZERO_2326  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_705/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_704_2327 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_705/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_5_inst_cy_705/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_779),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_704)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7791.INIT = 16'hE2FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7791 (
    .ADR0(DLX_IDinst_RegFile_0_12),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR2(DLX_IDinst_RegFile_1_12),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_571),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_779)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7801.INIT = 16'hFD5D;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7801 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_572),
    .ADR1(DLX_IDinst_RegFile_2_12),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR3(DLX_IDinst_RegFile_3_12),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_780)
  );
  X_BUF \DLX_IDinst_Mmux__COND_5_inst_cy_705/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_5_inst_cy_705/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_705)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_705_2328 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_705/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_704),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_780),
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_705/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mmux__COND_5_inst_cy_625/LOGIC_ONE_2329  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_625/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_5_inst_cy_625/LOGIC_ZERO_2330  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_625/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_624_2331 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_625/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_5_inst_cy_625/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_699),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_624)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6991.INIT = 16'hD8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6991 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR1(DLX_IDinst_RegFile_1_7),
    .ADR2(DLX_IDinst_RegFile_0_7),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_571),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_699)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7001.INIT = 16'hBF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7001 (
    .ADR0(DLX_IDinst_RegFile_3_7),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_572),
    .ADR3(DLX_IDinst_RegFile_2_7),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_700)
  );
  X_BUF \DLX_IDinst_Mmux__COND_5_inst_cy_625/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_5_inst_cy_625/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_625)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_625_2332 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_625/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_624),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_700),
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_625/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mmux__COND_5_inst_cy_545/LOGIC_ONE_2333  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_545/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_5_inst_cy_545/LOGIC_ZERO_2334  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_545/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_544_2335 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_545/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_5_inst_cy_545/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_619),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_544)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6191.INIT = 16'hACFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6191 (
    .ADR0(DLX_IDinst_RegFile_1_2),
    .ADR1(DLX_IDinst_RegFile_0_2),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_571),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_619)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6201.INIT = 16'hF7B3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6201 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_572),
    .ADR2(DLX_IDinst_RegFile_3_2),
    .ADR3(DLX_IDinst_RegFile_2_2),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_620)
  );
  X_BUF \DLX_IDinst_Mmux__COND_5_inst_cy_545/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_5_inst_cy_545/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_545)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_545_2336 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_545/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_544),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_620),
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_545/CYMUXG )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_5_inst_cy_557/LOGIC_ZERO_2337  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_557/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_556_2338 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_557/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_5_inst_cy_557/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_631),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_556)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6311.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6311 (
    .ADR0(DLX_IDinst_RegFile_24_2),
    .ADR1(DLX_IDinst_RegFile_25_2),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_583),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_631)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6321.INIT = 16'hE4FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6321 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR1(DLX_IDinst_RegFile_26_2),
    .ADR2(DLX_IDinst_RegFile_27_2),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_584),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_632)
  );
  X_BUF \DLX_IDinst_Mmux__COND_5_inst_cy_557/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_5_inst_cy_557/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_557)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_557_2339 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_557/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_556),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_632),
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_557/CYMUXG )
  );
  X_BUF \DLX_IDinst_Mmux__COND_5_inst_cy_557/CYINIT_2340  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_555),
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_557/CYINIT )
  );
  X_ONE \DLX_IDinst_Mmux__COND_5_inst_cy_801/LOGIC_ONE_2341  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_801/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_5_inst_cy_801/LOGIC_ZERO_2342  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_801/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_800_2343 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_801/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_5_inst_cy_801/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_875),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_800)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8751.INIT = 16'hDFD5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8751 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_571),
    .ADR1(DLX_IDinst_RegFile_1_18),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR3(DLX_IDinst_RegFile_0_18),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_875)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8761.INIT = 16'hDF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8761 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR1(DLX_IDinst_RegFile_3_18),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_572),
    .ADR3(DLX_IDinst_RegFile_2_18),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_876)
  );
  X_BUF \DLX_IDinst_Mmux__COND_5_inst_cy_801/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_5_inst_cy_801/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_801)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_801_2344 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_801/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_800),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_876),
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_801/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mmux__COND_5_inst_cy_721/LOGIC_ONE_2345  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_721/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_5_inst_cy_721/LOGIC_ZERO_2346  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_721/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_720_2347 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_721/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_5_inst_cy_721/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_795),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_720)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7951.INIT = 16'hE4FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7951 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR1(DLX_IDinst_RegFile_0_13),
    .ADR2(DLX_IDinst_RegFile_1_13),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_571),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_795)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7961.INIT = 16'hB8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7961 (
    .ADR0(DLX_IDinst_RegFile_3_13),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR2(DLX_IDinst_RegFile_2_13),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_572),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_796)
  );
  X_BUF \DLX_IDinst_Mmux__COND_5_inst_cy_721/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_5_inst_cy_721/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_721)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_721_2348 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_721/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_720),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_796),
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_721/CYMUXG )
  );
  X_ONE \DLX_EXinst_reg_out_B_EX<5>/LOGIC_ONE_2349  (
    .O(\DLX_EXinst_reg_out_B_EX<5>/LOGIC_ONE )
  );
  X_ZERO \DLX_EXinst_reg_out_B_EX<5>/LOGIC_ZERO_2350  (
    .O(\DLX_EXinst_reg_out_B_EX<5>/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_640_2351 (
    .IA(\DLX_EXinst_reg_out_B_EX<5>/LOGIC_ZERO ),
    .IB(\DLX_EXinst_reg_out_B_EX<5>/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_715),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_640)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7151.INIT = 16'hE4FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7151 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR1(DLX_IDinst_RegFile_0_8),
    .ADR2(DLX_IDinst_RegFile_1_8),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_571),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_715)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7161.INIT = 16'hFB73;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7161 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_572),
    .ADR2(DLX_IDinst_RegFile_2_8),
    .ADR3(DLX_IDinst_RegFile_3_8),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_716)
  );
  X_BUF \DLX_EXinst_reg_out_B_EX<5>/COUTUSED  (
    .I(\DLX_EXinst_reg_out_B_EX<5>/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_641)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_641_2352 (
    .IA(\DLX_EXinst_reg_out_B_EX<5>/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_640),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_716),
    .O(\DLX_EXinst_reg_out_B_EX<5>/CYMUXG )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_5_inst_cy_649/LOGIC_ZERO_2353  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_649/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_648_2354 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_649/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_5_inst_cy_649/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_723),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_648)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7231.INIT = 16'hF7B3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7231 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_579),
    .ADR2(DLX_IDinst_RegFile_17_8),
    .ADR3(DLX_IDinst_RegFile_16_8),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_723)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7241.INIT = 16'hBF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7241 (
    .ADR0(DLX_IDinst_RegFile_19_8),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_580),
    .ADR3(DLX_IDinst_RegFile_18_8),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_724)
  );
  X_BUF \DLX_IDinst_Mmux__COND_5_inst_cy_649/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_5_inst_cy_649/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_649)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_649_2355 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_649/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_648),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_724),
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_649/CYMUXG )
  );
  X_BUF \DLX_IDinst_Mmux__COND_5_inst_cy_649/CYINIT_2356  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_647),
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_649/CYINIT )
  );
  X_ONE \DLX_IDinst_Mmux__COND_5_inst_cy_561/LOGIC_ONE_2357  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_561/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_5_inst_cy_561/LOGIC_ZERO_2358  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_561/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_560_2359 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_561/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_5_inst_cy_561/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_635),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_560)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6351.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6351 (
    .ADR0(DLX_IDinst_RegFile_0_3),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_571),
    .ADR3(DLX_IDinst_RegFile_1_3),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_635)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6361.INIT = 16'hBF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6361 (
    .ADR0(DLX_IDinst_RegFile_3_3),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_572),
    .ADR3(DLX_IDinst_RegFile_2_3),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_636)
  );
  X_BUF \DLX_IDinst_Mmux__COND_5_inst_cy_561/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_5_inst_cy_561/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_561)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_561_2360 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_561/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_560),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_636),
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_561/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mmux__COND_5_inst_cy_897/LOGIC_ONE_2361  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_897/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_5_inst_cy_897/LOGIC_ZERO_2362  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_897/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_896_2363 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_897/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_5_inst_cy_897/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_971),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_896)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9711.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9711 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR1(DLX_IDinst_RegFile_0_24),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_571),
    .ADR3(DLX_IDinst_RegFile_1_24),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_971)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9721.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9721 (
    .ADR0(DLX_IDinst_RegFile_3_24),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_572),
    .ADR2(DLX_IDinst_RegFile_2_24),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_972)
  );
  X_BUF \DLX_IDinst_Mmux__COND_5_inst_cy_897/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_5_inst_cy_897/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_897)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_897_2364 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_897/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_896),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_972),
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_897/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mmux__COND_5_inst_cy_817/LOGIC_ONE_2365  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_817/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_5_inst_cy_817/LOGIC_ZERO_2366  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_817/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_816_2367 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_817/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_5_inst_cy_817/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_891),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_816)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8911.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8911 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR1(DLX_IDinst_RegFile_0_19),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_571),
    .ADR3(DLX_IDinst_RegFile_1_19),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_891)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8921.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8921 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_572),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR2(DLX_IDinst_RegFile_2_19),
    .ADR3(DLX_IDinst_RegFile_3_19),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_892)
  );
  X_BUF \DLX_IDinst_Mmux__COND_5_inst_cy_817/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_5_inst_cy_817/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_817)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_817_2368 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_817/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_816),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_892),
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_817/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mmux__COND_5_inst_cy_737/LOGIC_ONE_2369  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_737/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_5_inst_cy_737/LOGIC_ZERO_2370  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_737/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_736_2371 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_737/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_5_inst_cy_737/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_811),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_736)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8111.INIT = 16'hDDF5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8111 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_571),
    .ADR1(DLX_IDinst_RegFile_1_14),
    .ADR2(DLX_IDinst_RegFile_0_14),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_811)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8121.INIT = 16'hAFCF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8121 (
    .ADR0(DLX_IDinst_RegFile_3_14),
    .ADR1(DLX_IDinst_RegFile_2_14),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_572),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_812)
  );
  X_BUF \DLX_IDinst_Mmux__COND_5_inst_cy_737/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_5_inst_cy_737/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_737)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_737_2372 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_737/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_736),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_812),
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_737/CYMUXG )
  );
  defparam DLX_IDinst_RegFile_29_16_2373.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_29_16_2373 (
    .I(DLX_IDinst_WB_data_eff[16]),
    .CE(DLX_IDinst__n0608),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_29_16)
  );
  X_ZERO \DLX_IDinst_Mmux__COND_5_inst_cy_741/LOGIC_ZERO_2374  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_741/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_740_2375 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_741/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_5_inst_cy_741/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_815),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_740)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8151.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8151 (
    .ADR0(DLX_IDinst_RegFile_8_14),
    .ADR1(DLX_IDinst_RegFile_9_14),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_575),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_815)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8161.INIT = 16'hF7D5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8161 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_576),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR2(DLX_IDinst_RegFile_11_14),
    .ADR3(DLX_IDinst_RegFile_10_14),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_816)
  );
  X_BUF \DLX_IDinst_Mmux__COND_5_inst_cy_741/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_5_inst_cy_741/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_741)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_741_2376 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_741/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_740),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_816),
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_741/CYMUXG )
  );
  X_BUF \DLX_IDinst_Mmux__COND_5_inst_cy_741/CYINIT_2377  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_739),
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_741/CYINIT )
  );
  X_ONE \DLX_IDinst_Mmux__COND_5_inst_cy_657/LOGIC_ONE_2378  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_657/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_5_inst_cy_657/LOGIC_ZERO_2379  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_657/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_656_2380 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_657/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_5_inst_cy_657/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_731),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_656)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7311.INIT = 16'hAFCF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7311 (
    .ADR0(DLX_IDinst_RegFile_1_9),
    .ADR1(DLX_IDinst_RegFile_0_9),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_571),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_731)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7321.INIT = 16'hDF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7321 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR1(DLX_IDinst_RegFile_3_9),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_572),
    .ADR3(DLX_IDinst_RegFile_2_9),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_732)
  );
  X_BUF \DLX_IDinst_Mmux__COND_5_inst_cy_657/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_5_inst_cy_657/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_657)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_657_2381 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_657/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_656),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_732),
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_657/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mmux__COND_5_inst_cy_577/LOGIC_ONE_2382  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_577/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_5_inst_cy_577/LOGIC_ZERO_2383  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_577/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_576_2384 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_577/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_5_inst_cy_577/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_651),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_576)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6511.INIT = 16'hDF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6511 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR1(DLX_IDinst_RegFile_1_4),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_571),
    .ADR3(DLX_IDinst_RegFile_0_4),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_651)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_6521.INIT = 16'hB8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_6521 (
    .ADR0(DLX_IDinst_RegFile_3_4),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_4 ),
    .ADR2(DLX_IDinst_RegFile_2_4),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_572),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_652)
  );
  X_BUF \DLX_IDinst_Mmux__COND_5_inst_cy_577/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_5_inst_cy_577/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_577)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_577_2385 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_577/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_576),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_652),
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_577/CYMUXG )
  );
  defparam DLX_IDinst_RegFile_29_24_2386.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_29_24_2386 (
    .I(DLX_IDinst_WB_data_eff[24]),
    .CE(DLX_IDinst__n0608),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_29_24)
  );
  X_ONE \DLX_IDinst_Mmux__COND_5_inst_cy_913/LOGIC_ONE_2387  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_913/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_5_inst_cy_913/LOGIC_ZERO_2388  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_913/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_912_2389 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_913/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_5_inst_cy_913/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_987),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_912)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9871.INIT = 16'hACFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9871 (
    .ADR0(DLX_IDinst_RegFile_1_25),
    .ADR1(DLX_IDinst_RegFile_0_25),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_571),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_987)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9881.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9881 (
    .ADR0(DLX_IDinst_RegFile_2_25),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_572),
    .ADR3(DLX_IDinst_RegFile_3_25),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_988)
  );
  X_BUF \DLX_IDinst_Mmux__COND_5_inst_cy_913/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_5_inst_cy_913/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_913)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_913_2390 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_913/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_912),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_988),
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_913/CYMUXG )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_5_inst_cy_925/LOGIC_ZERO_2391  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_925/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_924_2392 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_925/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_5_inst_cy_925/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_999),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_924)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9991.INIT = 16'hBF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9991 (
    .ADR0(DLX_IDinst_RegFile_25_25),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_583),
    .ADR3(DLX_IDinst_RegFile_24_25),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_999)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10001.INIT = 16'hE4FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10001 (
    .ADR0(DLX_IDinst_jtarget[21]),
    .ADR1(DLX_IDinst_RegFile_26_25),
    .ADR2(DLX_IDinst_RegFile_27_25),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_584),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1000)
  );
  X_BUF \DLX_IDinst_Mmux__COND_5_inst_cy_925/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_5_inst_cy_925/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_925)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_925_2393 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_925/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_924),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1000),
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_925/CYMUXG )
  );
  X_BUF \DLX_IDinst_Mmux__COND_5_inst_cy_925/CYINIT_2394  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_923),
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_925/CYINIT )
  );
  X_ONE \DLX_IDinst_Mmux__COND_5_inst_cy_833/LOGIC_ONE_2395  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_833/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_5_inst_cy_833/LOGIC_ZERO_2396  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_833/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_832_2397 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_833/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_5_inst_cy_833/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_907),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_832)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9071.INIT = 16'hF5DD;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9071 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_571),
    .ADR1(DLX_IDinst_RegFile_0_20),
    .ADR2(DLX_IDinst_RegFile_1_20),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_907)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9081.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9081 (
    .ADR0(DLX_IDinst_RegFile_2_20),
    .ADR1(DLX_IDinst_RegFile_3_20),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_572),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_908)
  );
  X_BUF \DLX_IDinst_Mmux__COND_5_inst_cy_833/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_5_inst_cy_833/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_833)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_833_2398 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_833/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_832),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_908),
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_833/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mmux__COND_5_inst_cy_753/LOGIC_ONE_2399  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_753/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_5_inst_cy_753/LOGIC_ZERO_2400  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_753/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_752_2401 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_753/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_5_inst_cy_753/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_827),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_752)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8271.INIT = 16'hD8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8271 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR1(DLX_IDinst_RegFile_1_15),
    .ADR2(DLX_IDinst_RegFile_0_15),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_571),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_827)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8281.INIT = 16'hF7D5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8281 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_572),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR2(DLX_IDinst_RegFile_3_15),
    .ADR3(DLX_IDinst_RegFile_2_15),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_828)
  );
  X_BUF \DLX_IDinst_Mmux__COND_5_inst_cy_753/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_5_inst_cy_753/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_753)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_753_2402 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_753/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_752),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_828),
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_753/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mmux__COND_5_inst_cy_673/LOGIC_ONE_2403  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_673/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_5_inst_cy_673/LOGIC_ZERO_2404  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_673/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_672_2405 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_673/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_5_inst_cy_673/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_747),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_672)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7471.INIT = 16'hDF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7471 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR1(DLX_IDinst_RegFile_1_10),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_571),
    .ADR3(DLX_IDinst_RegFile_0_10),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_747)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7481.INIT = 16'hCFAF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7481 (
    .ADR0(DLX_IDinst_RegFile_2_10),
    .ADR1(DLX_IDinst_RegFile_3_10),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_572),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_748)
  );
  X_BUF \DLX_IDinst_Mmux__COND_5_inst_cy_673/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_5_inst_cy_673/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_673)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_673_2406 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_673/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_672),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_748),
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_673/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mmux__COND_5_inst_cy_929/LOGIC_ONE_2407  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_929/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_5_inst_cy_929/LOGIC_ZERO_2408  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_929/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_928_2409 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_929/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_5_inst_cy_929/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1003),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_928)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10031.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10031 (
    .ADR0(DLX_IDinst_RegFile_0_26),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_571),
    .ADR2(DLX_IDinst_RegFile_1_26),
    .ADR3(DLX_IDinst_jtarget[21]),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1003)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10041.INIT = 16'hFD5D;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10041 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_572),
    .ADR1(DLX_IDinst_RegFile_2_26),
    .ADR2(DLX_IDinst_jtarget[21]),
    .ADR3(DLX_IDinst_RegFile_3_26),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1004)
  );
  X_BUF \DLX_IDinst_Mmux__COND_5_inst_cy_929/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_5_inst_cy_929/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_929)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_929_2410 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_929/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_928),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1004),
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_929/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mmux__COND_5_inst_cy_849/LOGIC_ONE_2411  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_849/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_5_inst_cy_849/LOGIC_ZERO_2412  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_849/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_848_2413 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_849/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_5_inst_cy_849/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_923),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_848)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9231.INIT = 16'hCFAF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9231 (
    .ADR0(DLX_IDinst_RegFile_0_21),
    .ADR1(DLX_IDinst_RegFile_1_21),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_571),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_923)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9241.INIT = 16'hF5DD;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9241 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_572),
    .ADR1(DLX_IDinst_RegFile_2_21),
    .ADR2(DLX_IDinst_RegFile_3_21),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_924)
  );
  X_BUF \DLX_IDinst_Mmux__COND_5_inst_cy_849/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_5_inst_cy_849/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_849)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_849_2414 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_849/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_848),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_924),
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_849/CYMUXG )
  );
  X_ONE \DLX_MEMinst_opcode_of_WB<4>/LOGIC_ONE_2415  (
    .O(\DLX_MEMinst_opcode_of_WB<4>/LOGIC_ONE )
  );
  X_ZERO \DLX_MEMinst_opcode_of_WB<4>/LOGIC_ZERO_2416  (
    .O(\DLX_MEMinst_opcode_of_WB<4>/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_768_2417 (
    .IA(\DLX_MEMinst_opcode_of_WB<4>/LOGIC_ZERO ),
    .IB(\DLX_MEMinst_opcode_of_WB<4>/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_843),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_768)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8431.INIT = 16'hDFD5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8431 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_571),
    .ADR1(DLX_IDinst_RegFile_1_16),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR3(DLX_IDinst_RegFile_0_16),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_843)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8441.INIT = 16'hACFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8441 (
    .ADR0(DLX_IDinst_RegFile_3_16),
    .ADR1(DLX_IDinst_RegFile_2_16),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_572),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_844)
  );
  X_BUF \DLX_MEMinst_opcode_of_WB<4>/COUTUSED  (
    .I(\DLX_MEMinst_opcode_of_WB<4>/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_769)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_769_2418 (
    .IA(\DLX_MEMinst_opcode_of_WB<4>/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_768),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_844),
    .O(\DLX_MEMinst_opcode_of_WB<4>/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mmux__COND_5_inst_cy_865/LOGIC_ONE_2419  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_865/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_5_inst_cy_865/LOGIC_ZERO_2420  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_865/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_864_2421 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_865/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_5_inst_cy_865/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_939),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_864)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9391.INIT = 16'hBFB3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9391 (
    .ADR0(DLX_IDinst_RegFile_1_22),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_571),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR3(DLX_IDinst_RegFile_0_22),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_939)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9401.INIT = 16'hF7D5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9401 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_572),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR2(DLX_IDinst_RegFile_3_22),
    .ADR3(DLX_IDinst_RegFile_2_22),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_940)
  );
  X_BUF \DLX_IDinst_Mmux__COND_5_inst_cy_865/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_5_inst_cy_865/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_865)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_865_2422 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_865/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_864),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_940),
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_865/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mmux__COND_5_inst_cy_785/LOGIC_ONE_2423  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_785/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_5_inst_cy_785/LOGIC_ZERO_2424  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_785/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_784_2425 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_785/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_5_inst_cy_785/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_859),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_784)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8591.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8591 (
    .ADR0(DLX_IDinst_RegFile_0_17),
    .ADR1(DLX_IDinst_RegFile_1_17),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_571),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_859)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8601.INIT = 16'hCFAF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8601 (
    .ADR0(DLX_IDinst_RegFile_2_17),
    .ADR1(DLX_IDinst_RegFile_3_17),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_572),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_860)
  );
  X_BUF \DLX_IDinst_Mmux__COND_5_inst_cy_785/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_5_inst_cy_785/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_785)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_785_2426 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_785/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_784),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_860),
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_785/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mmux__COND_5_inst_cy_945/LOGIC_ONE_2427  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_945/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_5_inst_cy_945/LOGIC_ZERO_2428  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_945/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_944_2429 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_945/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_5_inst_cy_945/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1019),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_944)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10191.INIT = 16'hF5DD;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10191 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_571),
    .ADR1(DLX_IDinst_RegFile_0_27),
    .ADR2(DLX_IDinst_RegFile_1_27),
    .ADR3(DLX_IDinst_jtarget[21]),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1019)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10201.INIT = 16'hDF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10201 (
    .ADR0(DLX_IDinst_jtarget[21]),
    .ADR1(DLX_IDinst_RegFile_3_27),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_572),
    .ADR3(DLX_IDinst_RegFile_2_27),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1020)
  );
  X_BUF \DLX_IDinst_Mmux__COND_5_inst_cy_945/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_5_inst_cy_945/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_945)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_945_2430 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_945/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_944),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1020),
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_945/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mmux__COND_5_inst_cy_881/LOGIC_ONE_2431  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_881/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_5_inst_cy_881/LOGIC_ZERO_2432  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_881/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_880_2433 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_881/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_5_inst_cy_881/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_955),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_880)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9551.INIT = 16'hE2FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9551 (
    .ADR0(DLX_IDinst_RegFile_0_23),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR2(DLX_IDinst_RegFile_1_23),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_571),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_955)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9561.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9561 (
    .ADR0(DLX_IDinst_RegFile_2_23),
    .ADR1(DLX_IDinst_RegFile_3_23),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_572),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_956)
  );
  X_BUF \DLX_IDinst_Mmux__COND_5_inst_cy_881/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_5_inst_cy_881/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_881)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_881_2434 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_881/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_880),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_956),
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_881/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mmux__COND_5_inst_cy_961/LOGIC_ONE_2435  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_961/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_5_inst_cy_961/LOGIC_ZERO_2436  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_961/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_960_2437 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_961/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_5_inst_cy_961/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1035),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_960)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10351.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10351 (
    .ADR0(DLX_IDinst_RegFile_1_28),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_571),
    .ADR2(DLX_IDinst_RegFile_0_28),
    .ADR3(DLX_IDinst_jtarget[21]),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1035)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10361.INIT = 16'hD8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10361 (
    .ADR0(DLX_IDinst_jtarget[21]),
    .ADR1(DLX_IDinst_RegFile_3_28),
    .ADR2(DLX_IDinst_RegFile_2_28),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_572),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1036)
  );
  X_BUF \DLX_IDinst_Mmux__COND_5_inst_cy_961/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_5_inst_cy_961/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_961)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_961_2438 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_961/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_960),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1036),
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_961/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mmux__COND_5_inst_cy_977/LOGIC_ONE_2439  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_977/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_5_inst_cy_977/LOGIC_ZERO_2440  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_977/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_976_2441 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_977/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_5_inst_cy_977/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1051),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_976)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10511.INIT = 16'hBF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10511 (
    .ADR0(DLX_IDinst_RegFile_1_29),
    .ADR1(DLX_IDinst_jtarget[21]),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_571),
    .ADR3(DLX_IDinst_RegFile_0_29),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1051)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10521.INIT = 16'hAFCF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10521 (
    .ADR0(DLX_IDinst_RegFile_3_29),
    .ADR1(DLX_IDinst_RegFile_2_29),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_572),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1052)
  );
  X_BUF \DLX_IDinst_Mmux__COND_5_inst_cy_977/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_5_inst_cy_977/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_977)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_977_2442 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_977/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_976),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1052),
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_977/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mmux__COND_5_inst_cy_993/LOGIC_ONE_2443  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_993/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_5_inst_cy_993/LOGIC_ZERO_2444  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_993/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_992_2445 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_993/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_5_inst_cy_993/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1067),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_992)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10671.INIT = 16'hFB3B;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10671 (
    .ADR0(DLX_IDinst_RegFile_0_30),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_571),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR3(DLX_IDinst_RegFile_1_30),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1067)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10681.INIT = 16'hDF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10681 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR1(DLX_IDinst_RegFile_3_30),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_572),
    .ADR3(DLX_IDinst_RegFile_2_30),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1068)
  );
  X_BUF \DLX_IDinst_Mmux__COND_5_inst_cy_993/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_5_inst_cy_993/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_993)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_993_2446 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_993/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_992),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1068),
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_993/CYMUXG )
  );
  X_MUX2 DLX_EXinst_Maddsub__n0012_inst_cy_70_2447 (
    .IA(DLX_IDinst_reg_out_A[0]),
    .IB(\DLX_IDinst_RegFile_3_16/CYINIT ),
    .SEL(DLX_EXinst_Maddsub__n0012_inst_lut3_2),
    .O(DLX_EXinst_Maddsub__n0012_inst_cy_70)
  );
  X_XOR2 DLX_EXinst_Maddsub__n0012_inst_sum_70 (
    .I0(\DLX_IDinst_RegFile_3_16/CYINIT ),
    .I1(DLX_EXinst_Maddsub__n0012_inst_lut3_2),
    .O(\DLX_IDinst_RegFile_3_16/XORF )
  );
  defparam DLX_EXinst_Maddsub__n0012_inst_lut3_210.INIT = 16'h9696;
  X_LUT4 DLX_EXinst_Maddsub__n0012_inst_lut3_210 (
    .ADR0(DLX_IDinst_reg_out_A[0]),
    .ADR1(DLX_EXinst__n0013[0]),
    .ADR2(N144912),
    .ADR3(VCC),
    .O(DLX_EXinst_Maddsub__n0012_inst_lut3_2)
  );
  defparam DLX_EXinst_Maddsub__n0012_inst_lut3_34.INIT = 16'h9696;
  X_LUT4 DLX_EXinst_Maddsub__n0012_inst_lut3_34 (
    .ADR0(DLX_IDinst_reg_out_A[1]),
    .ADR1(DLX_EXinst__n0013[1]),
    .ADR2(N144912),
    .ADR3(VCC),
    .O(DLX_EXinst_Maddsub__n0012_inst_lut3_3)
  );
  X_BUF \DLX_IDinst_RegFile_3_16/COUTUSED  (
    .I(\DLX_IDinst_RegFile_3_16/CYMUXG ),
    .O(DLX_EXinst_Maddsub__n0012_inst_cy_71)
  );
  X_BUF \DLX_IDinst_RegFile_3_16/XUSED  (
    .I(\DLX_IDinst_RegFile_3_16/XORF ),
    .O(DLX_EXinst__n0012[0])
  );
  X_BUF \DLX_IDinst_RegFile_3_16/YUSED  (
    .I(\DLX_IDinst_RegFile_3_16/XORG ),
    .O(DLX_EXinst__n0012[1])
  );
  X_MUX2 DLX_EXinst_Maddsub__n0012_inst_cy_71_2448 (
    .IA(DLX_IDinst_reg_out_A[1]),
    .IB(DLX_EXinst_Maddsub__n0012_inst_cy_70),
    .SEL(DLX_EXinst_Maddsub__n0012_inst_lut3_3),
    .O(\DLX_IDinst_RegFile_3_16/CYMUXG )
  );
  X_XOR2 DLX_EXinst_Maddsub__n0012_inst_sum_71 (
    .I0(DLX_EXinst_Maddsub__n0012_inst_cy_70),
    .I1(DLX_EXinst_Maddsub__n0012_inst_lut3_3),
    .O(\DLX_IDinst_RegFile_3_16/XORG )
  );
  X_BUF \DLX_IDinst_RegFile_3_16/CYINIT_2449  (
    .I(N144912),
    .O(\DLX_IDinst_RegFile_3_16/CYINIT )
  );
  X_MUX2 DLX_EXinst_Maddsub__n0012_inst_cy_72_2450 (
    .IA(DLX_IDinst_reg_out_A[2]),
    .IB(\DLX_EXinst__n0012<2>/CYINIT ),
    .SEL(DLX_EXinst_Maddsub__n0012_inst_lut3_4),
    .O(DLX_EXinst_Maddsub__n0012_inst_cy_72)
  );
  X_XOR2 DLX_EXinst_Maddsub__n0012_inst_sum_72 (
    .I0(\DLX_EXinst__n0012<2>/CYINIT ),
    .I1(DLX_EXinst_Maddsub__n0012_inst_lut3_4),
    .O(\DLX_EXinst__n0012<2>/XORF )
  );
  defparam DLX_EXinst_Maddsub__n0012_inst_lut3_41.INIT = 16'hA55A;
  X_LUT4 DLX_EXinst_Maddsub__n0012_inst_lut3_41 (
    .ADR0(DLX_IDinst_reg_out_A[2]),
    .ADR1(VCC),
    .ADR2(N144912),
    .ADR3(DLX_EXinst__n0013[2]),
    .O(DLX_EXinst_Maddsub__n0012_inst_lut3_4)
  );
  defparam DLX_EXinst_Maddsub__n0012_inst_lut3_51.INIT = 16'hA55A;
  X_LUT4 DLX_EXinst_Maddsub__n0012_inst_lut3_51 (
    .ADR0(DLX_IDinst_reg_out_A[3]),
    .ADR1(VCC),
    .ADR2(N144912),
    .ADR3(DLX_EXinst__n0013[3]),
    .O(DLX_EXinst_Maddsub__n0012_inst_lut3_5)
  );
  X_BUF \DLX_EXinst__n0012<2>/COUTUSED  (
    .I(\DLX_EXinst__n0012<2>/CYMUXG ),
    .O(DLX_EXinst_Maddsub__n0012_inst_cy_73)
  );
  X_BUF \DLX_EXinst__n0012<2>/XUSED  (
    .I(\DLX_EXinst__n0012<2>/XORF ),
    .O(DLX_EXinst__n0012[2])
  );
  X_BUF \DLX_EXinst__n0012<2>/YUSED  (
    .I(\DLX_EXinst__n0012<2>/XORG ),
    .O(DLX_EXinst__n0012[3])
  );
  X_MUX2 DLX_EXinst_Maddsub__n0012_inst_cy_73_2451 (
    .IA(DLX_IDinst_reg_out_A[3]),
    .IB(DLX_EXinst_Maddsub__n0012_inst_cy_72),
    .SEL(DLX_EXinst_Maddsub__n0012_inst_lut3_5),
    .O(\DLX_EXinst__n0012<2>/CYMUXG )
  );
  X_XOR2 DLX_EXinst_Maddsub__n0012_inst_sum_73 (
    .I0(DLX_EXinst_Maddsub__n0012_inst_cy_72),
    .I1(DLX_EXinst_Maddsub__n0012_inst_lut3_5),
    .O(\DLX_EXinst__n0012<2>/XORG )
  );
  X_BUF \DLX_EXinst__n0012<2>/CYINIT_2452  (
    .I(DLX_EXinst_Maddsub__n0012_inst_cy_71),
    .O(\DLX_EXinst__n0012<2>/CYINIT )
  );
  X_MUX2 DLX_EXinst_Maddsub__n0012_inst_cy_74_2453 (
    .IA(DLX_IDinst_reg_out_A[4]),
    .IB(\DLX_EXinst__n0012<4>/CYINIT ),
    .SEL(DLX_EXinst_Maddsub__n0012_inst_lut3_6),
    .O(DLX_EXinst_Maddsub__n0012_inst_cy_74)
  );
  X_XOR2 DLX_EXinst_Maddsub__n0012_inst_sum_74 (
    .I0(\DLX_EXinst__n0012<4>/CYINIT ),
    .I1(DLX_EXinst_Maddsub__n0012_inst_lut3_6),
    .O(\DLX_EXinst__n0012<4>/XORF )
  );
  defparam DLX_EXinst_Maddsub__n0012_inst_lut3_61.INIT = 16'hA55A;
  X_LUT4 DLX_EXinst_Maddsub__n0012_inst_lut3_61 (
    .ADR0(DLX_IDinst_reg_out_A[4]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst__n0013[4]),
    .ADR3(N144912),
    .O(DLX_EXinst_Maddsub__n0012_inst_lut3_6)
  );
  defparam DLX_EXinst_Maddsub__n0012_inst_lut3_71.INIT = 16'hA55A;
  X_LUT4 DLX_EXinst_Maddsub__n0012_inst_lut3_71 (
    .ADR0(DLX_IDinst_reg_out_A[5]),
    .ADR1(VCC),
    .ADR2(N144912),
    .ADR3(DLX_EXinst__n0013[5]),
    .O(DLX_EXinst_Maddsub__n0012_inst_lut3_7)
  );
  X_BUF \DLX_EXinst__n0012<4>/COUTUSED  (
    .I(\DLX_EXinst__n0012<4>/CYMUXG ),
    .O(DLX_EXinst_Maddsub__n0012_inst_cy_75)
  );
  X_BUF \DLX_EXinst__n0012<4>/XUSED  (
    .I(\DLX_EXinst__n0012<4>/XORF ),
    .O(DLX_EXinst__n0012[4])
  );
  X_BUF \DLX_EXinst__n0012<4>/YUSED  (
    .I(\DLX_EXinst__n0012<4>/XORG ),
    .O(DLX_EXinst__n0012[5])
  );
  X_MUX2 DLX_EXinst_Maddsub__n0012_inst_cy_75_2454 (
    .IA(DLX_IDinst_reg_out_A[5]),
    .IB(DLX_EXinst_Maddsub__n0012_inst_cy_74),
    .SEL(DLX_EXinst_Maddsub__n0012_inst_lut3_7),
    .O(\DLX_EXinst__n0012<4>/CYMUXG )
  );
  X_XOR2 DLX_EXinst_Maddsub__n0012_inst_sum_75 (
    .I0(DLX_EXinst_Maddsub__n0012_inst_cy_74),
    .I1(DLX_EXinst_Maddsub__n0012_inst_lut3_7),
    .O(\DLX_EXinst__n0012<4>/XORG )
  );
  X_BUF \DLX_EXinst__n0012<4>/CYINIT_2455  (
    .I(DLX_EXinst_Maddsub__n0012_inst_cy_73),
    .O(\DLX_EXinst__n0012<4>/CYINIT )
  );
  X_MUX2 DLX_EXinst_Maddsub__n0012_inst_cy_76_2456 (
    .IA(DLX_IDinst_reg_out_A[6]),
    .IB(\DLX_EXinst__n0012<6>/CYINIT ),
    .SEL(DLX_EXinst_Maddsub__n0012_inst_lut3_8),
    .O(DLX_EXinst_Maddsub__n0012_inst_cy_76)
  );
  X_XOR2 DLX_EXinst_Maddsub__n0012_inst_sum_76 (
    .I0(\DLX_EXinst__n0012<6>/CYINIT ),
    .I1(DLX_EXinst_Maddsub__n0012_inst_lut3_8),
    .O(\DLX_EXinst__n0012<6>/XORF )
  );
  defparam DLX_EXinst_Maddsub__n0012_inst_lut3_81.INIT = 16'hA55A;
  X_LUT4 DLX_EXinst_Maddsub__n0012_inst_lut3_81 (
    .ADR0(DLX_IDinst_reg_out_A[6]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst__n0013[6]),
    .ADR3(N144912),
    .O(DLX_EXinst_Maddsub__n0012_inst_lut3_8)
  );
  defparam DLX_EXinst_Maddsub__n0012_inst_lut3_91.INIT = 16'h9966;
  X_LUT4 DLX_EXinst_Maddsub__n0012_inst_lut3_91 (
    .ADR0(DLX_IDinst_reg_out_A[7]),
    .ADR1(N144912),
    .ADR2(VCC),
    .ADR3(DLX_EXinst__n0013[7]),
    .O(DLX_EXinst_Maddsub__n0012_inst_lut3_9)
  );
  X_BUF \DLX_EXinst__n0012<6>/COUTUSED  (
    .I(\DLX_EXinst__n0012<6>/CYMUXG ),
    .O(DLX_EXinst_Maddsub__n0012_inst_cy_77)
  );
  X_BUF \DLX_EXinst__n0012<6>/XUSED  (
    .I(\DLX_EXinst__n0012<6>/XORF ),
    .O(DLX_EXinst__n0012[6])
  );
  X_BUF \DLX_EXinst__n0012<6>/YUSED  (
    .I(\DLX_EXinst__n0012<6>/XORG ),
    .O(DLX_EXinst__n0012[7])
  );
  X_MUX2 DLX_EXinst_Maddsub__n0012_inst_cy_77_2457 (
    .IA(DLX_IDinst_reg_out_A[7]),
    .IB(DLX_EXinst_Maddsub__n0012_inst_cy_76),
    .SEL(DLX_EXinst_Maddsub__n0012_inst_lut3_9),
    .O(\DLX_EXinst__n0012<6>/CYMUXG )
  );
  X_XOR2 DLX_EXinst_Maddsub__n0012_inst_sum_77 (
    .I0(DLX_EXinst_Maddsub__n0012_inst_cy_76),
    .I1(DLX_EXinst_Maddsub__n0012_inst_lut3_9),
    .O(\DLX_EXinst__n0012<6>/XORG )
  );
  X_BUF \DLX_EXinst__n0012<6>/CYINIT_2458  (
    .I(DLX_EXinst_Maddsub__n0012_inst_cy_75),
    .O(\DLX_EXinst__n0012<6>/CYINIT )
  );
  X_MUX2 DLX_EXinst_Maddsub__n0012_inst_cy_78_2459 (
    .IA(DLX_IDinst_reg_out_A[8]),
    .IB(\DLX_IDinst_RegFile_26_10/CYINIT ),
    .SEL(DLX_EXinst_Maddsub__n0012_inst_lut3_10),
    .O(DLX_EXinst_Maddsub__n0012_inst_cy_78)
  );
  X_XOR2 DLX_EXinst_Maddsub__n0012_inst_sum_78 (
    .I0(\DLX_IDinst_RegFile_26_10/CYINIT ),
    .I1(DLX_EXinst_Maddsub__n0012_inst_lut3_10),
    .O(\DLX_IDinst_RegFile_26_10/XORF )
  );
  defparam DLX_EXinst_Maddsub__n0012_inst_lut3_101.INIT = 16'h9966;
  X_LUT4 DLX_EXinst_Maddsub__n0012_inst_lut3_101 (
    .ADR0(DLX_IDinst_reg_out_A[8]),
    .ADR1(DLX_EXinst__n0013[8]),
    .ADR2(VCC),
    .ADR3(N144912),
    .O(DLX_EXinst_Maddsub__n0012_inst_lut3_10)
  );
  defparam DLX_EXinst_Maddsub__n0012_inst_lut3_111.INIT = 16'hA55A;
  X_LUT4 DLX_EXinst_Maddsub__n0012_inst_lut3_111 (
    .ADR0(DLX_IDinst_reg_out_A[9]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst__n0013[9]),
    .ADR3(N144912),
    .O(DLX_EXinst_Maddsub__n0012_inst_lut3_11)
  );
  X_BUF \DLX_IDinst_RegFile_26_10/COUTUSED  (
    .I(\DLX_IDinst_RegFile_26_10/CYMUXG ),
    .O(DLX_EXinst_Maddsub__n0012_inst_cy_79)
  );
  X_BUF \DLX_IDinst_RegFile_26_10/XUSED  (
    .I(\DLX_IDinst_RegFile_26_10/XORF ),
    .O(DLX_EXinst__n0012[8])
  );
  X_BUF \DLX_IDinst_RegFile_26_10/YUSED  (
    .I(\DLX_IDinst_RegFile_26_10/XORG ),
    .O(DLX_EXinst__n0012[9])
  );
  X_MUX2 DLX_EXinst_Maddsub__n0012_inst_cy_79_2460 (
    .IA(DLX_IDinst_reg_out_A[9]),
    .IB(DLX_EXinst_Maddsub__n0012_inst_cy_78),
    .SEL(DLX_EXinst_Maddsub__n0012_inst_lut3_11),
    .O(\DLX_IDinst_RegFile_26_10/CYMUXG )
  );
  X_XOR2 DLX_EXinst_Maddsub__n0012_inst_sum_79 (
    .I0(DLX_EXinst_Maddsub__n0012_inst_cy_78),
    .I1(DLX_EXinst_Maddsub__n0012_inst_lut3_11),
    .O(\DLX_IDinst_RegFile_26_10/XORG )
  );
  X_BUF \DLX_IDinst_RegFile_26_10/CYINIT_2461  (
    .I(DLX_EXinst_Maddsub__n0012_inst_cy_77),
    .O(\DLX_IDinst_RegFile_26_10/CYINIT )
  );
  X_MUX2 DLX_EXinst_Maddsub__n0012_inst_cy_80_2462 (
    .IA(DLX_IDinst_reg_out_A[10]),
    .IB(\DLX_EXinst__n0012<10>/CYINIT ),
    .SEL(DLX_EXinst_Maddsub__n0012_inst_lut3_12),
    .O(DLX_EXinst_Maddsub__n0012_inst_cy_80)
  );
  X_XOR2 DLX_EXinst_Maddsub__n0012_inst_sum_80 (
    .I0(\DLX_EXinst__n0012<10>/CYINIT ),
    .I1(DLX_EXinst_Maddsub__n0012_inst_lut3_12),
    .O(\DLX_EXinst__n0012<10>/XORF )
  );
  defparam DLX_EXinst_Maddsub__n0012_inst_lut3_121.INIT = 16'hA55A;
  X_LUT4 DLX_EXinst_Maddsub__n0012_inst_lut3_121 (
    .ADR0(DLX_IDinst_reg_out_A[10]),
    .ADR1(VCC),
    .ADR2(N144912),
    .ADR3(DLX_EXinst__n0013[10]),
    .O(DLX_EXinst_Maddsub__n0012_inst_lut3_12)
  );
  defparam DLX_EXinst_Maddsub__n0012_inst_lut3_131.INIT = 16'h9696;
  X_LUT4 DLX_EXinst_Maddsub__n0012_inst_lut3_131 (
    .ADR0(DLX_IDinst_reg_out_A[11]),
    .ADR1(DLX_EXinst__n0013[11]),
    .ADR2(N144912),
    .ADR3(VCC),
    .O(DLX_EXinst_Maddsub__n0012_inst_lut3_13)
  );
  X_BUF \DLX_EXinst__n0012<10>/COUTUSED  (
    .I(\DLX_EXinst__n0012<10>/CYMUXG ),
    .O(DLX_EXinst_Maddsub__n0012_inst_cy_81)
  );
  X_BUF \DLX_EXinst__n0012<10>/XUSED  (
    .I(\DLX_EXinst__n0012<10>/XORF ),
    .O(DLX_EXinst__n0012[10])
  );
  X_BUF \DLX_EXinst__n0012<10>/YUSED  (
    .I(\DLX_EXinst__n0012<10>/XORG ),
    .O(DLX_EXinst__n0012[11])
  );
  X_MUX2 DLX_EXinst_Maddsub__n0012_inst_cy_81_2463 (
    .IA(DLX_IDinst_reg_out_A[11]),
    .IB(DLX_EXinst_Maddsub__n0012_inst_cy_80),
    .SEL(DLX_EXinst_Maddsub__n0012_inst_lut3_13),
    .O(\DLX_EXinst__n0012<10>/CYMUXG )
  );
  X_XOR2 DLX_EXinst_Maddsub__n0012_inst_sum_81 (
    .I0(DLX_EXinst_Maddsub__n0012_inst_cy_80),
    .I1(DLX_EXinst_Maddsub__n0012_inst_lut3_13),
    .O(\DLX_EXinst__n0012<10>/XORG )
  );
  X_BUF \DLX_EXinst__n0012<10>/CYINIT_2464  (
    .I(DLX_EXinst_Maddsub__n0012_inst_cy_79),
    .O(\DLX_EXinst__n0012<10>/CYINIT )
  );
  X_MUX2 DLX_EXinst_Maddsub__n0012_inst_cy_82_2465 (
    .IA(DLX_IDinst_reg_out_A[12]),
    .IB(\DLX_EXinst__n0012<12>/CYINIT ),
    .SEL(DLX_EXinst_Maddsub__n0012_inst_lut3_14),
    .O(DLX_EXinst_Maddsub__n0012_inst_cy_82)
  );
  X_XOR2 DLX_EXinst_Maddsub__n0012_inst_sum_82 (
    .I0(\DLX_EXinst__n0012<12>/CYINIT ),
    .I1(DLX_EXinst_Maddsub__n0012_inst_lut3_14),
    .O(\DLX_EXinst__n0012<12>/XORF )
  );
  defparam DLX_EXinst_Maddsub__n0012_inst_lut3_141.INIT = 16'h9966;
  X_LUT4 DLX_EXinst_Maddsub__n0012_inst_lut3_141 (
    .ADR0(DLX_IDinst_reg_out_A[12]),
    .ADR1(N144912),
    .ADR2(VCC),
    .ADR3(DLX_EXinst__n0013[12]),
    .O(DLX_EXinst_Maddsub__n0012_inst_lut3_14)
  );
  defparam DLX_EXinst_Maddsub__n0012_inst_lut3_151.INIT = 16'h9696;
  X_LUT4 DLX_EXinst_Maddsub__n0012_inst_lut3_151 (
    .ADR0(DLX_IDinst_reg_out_A[13]),
    .ADR1(N144912),
    .ADR2(DLX_EXinst__n0013[13]),
    .ADR3(VCC),
    .O(DLX_EXinst_Maddsub__n0012_inst_lut3_15)
  );
  X_BUF \DLX_EXinst__n0012<12>/COUTUSED  (
    .I(\DLX_EXinst__n0012<12>/CYMUXG ),
    .O(DLX_EXinst_Maddsub__n0012_inst_cy_83)
  );
  X_BUF \DLX_EXinst__n0012<12>/XUSED  (
    .I(\DLX_EXinst__n0012<12>/XORF ),
    .O(DLX_EXinst__n0012[12])
  );
  X_BUF \DLX_EXinst__n0012<12>/YUSED  (
    .I(\DLX_EXinst__n0012<12>/XORG ),
    .O(DLX_EXinst__n0012[13])
  );
  X_MUX2 DLX_EXinst_Maddsub__n0012_inst_cy_83_2466 (
    .IA(DLX_IDinst_reg_out_A[13]),
    .IB(DLX_EXinst_Maddsub__n0012_inst_cy_82),
    .SEL(DLX_EXinst_Maddsub__n0012_inst_lut3_15),
    .O(\DLX_EXinst__n0012<12>/CYMUXG )
  );
  X_XOR2 DLX_EXinst_Maddsub__n0012_inst_sum_83 (
    .I0(DLX_EXinst_Maddsub__n0012_inst_cy_82),
    .I1(DLX_EXinst_Maddsub__n0012_inst_lut3_15),
    .O(\DLX_EXinst__n0012<12>/XORG )
  );
  X_BUF \DLX_EXinst__n0012<12>/CYINIT_2467  (
    .I(DLX_EXinst_Maddsub__n0012_inst_cy_81),
    .O(\DLX_EXinst__n0012<12>/CYINIT )
  );
  X_MUX2 DLX_EXinst_Maddsub__n0012_inst_cy_84_2468 (
    .IA(DLX_IDinst_reg_out_A[14]),
    .IB(\DLX_EXinst__n0012<14>/CYINIT ),
    .SEL(DLX_EXinst_Maddsub__n0012_inst_lut3_16),
    .O(DLX_EXinst_Maddsub__n0012_inst_cy_84)
  );
  X_XOR2 DLX_EXinst_Maddsub__n0012_inst_sum_84 (
    .I0(\DLX_EXinst__n0012<14>/CYINIT ),
    .I1(DLX_EXinst_Maddsub__n0012_inst_lut3_16),
    .O(\DLX_EXinst__n0012<14>/XORF )
  );
  defparam DLX_EXinst_Maddsub__n0012_inst_lut3_161.INIT = 16'h9696;
  X_LUT4 DLX_EXinst_Maddsub__n0012_inst_lut3_161 (
    .ADR0(DLX_IDinst_reg_out_A[14]),
    .ADR1(DLX_EXinst__n0013[14]),
    .ADR2(N144912),
    .ADR3(VCC),
    .O(DLX_EXinst_Maddsub__n0012_inst_lut3_16)
  );
  defparam DLX_EXinst_Maddsub__n0012_inst_lut3_171.INIT = 16'h9696;
  X_LUT4 DLX_EXinst_Maddsub__n0012_inst_lut3_171 (
    .ADR0(DLX_IDinst_reg_out_A[15]),
    .ADR1(N144912),
    .ADR2(DLX_EXinst__n0013[15]),
    .ADR3(VCC),
    .O(DLX_EXinst_Maddsub__n0012_inst_lut3_17)
  );
  X_BUF \DLX_EXinst__n0012<14>/COUTUSED  (
    .I(\DLX_EXinst__n0012<14>/CYMUXG ),
    .O(DLX_EXinst_Maddsub__n0012_inst_cy_85)
  );
  X_BUF \DLX_EXinst__n0012<14>/XUSED  (
    .I(\DLX_EXinst__n0012<14>/XORF ),
    .O(DLX_EXinst__n0012[14])
  );
  X_BUF \DLX_EXinst__n0012<14>/YUSED  (
    .I(\DLX_EXinst__n0012<14>/XORG ),
    .O(DLX_EXinst__n0012[15])
  );
  X_MUX2 DLX_EXinst_Maddsub__n0012_inst_cy_85_2469 (
    .IA(DLX_IDinst_reg_out_A[15]),
    .IB(DLX_EXinst_Maddsub__n0012_inst_cy_84),
    .SEL(DLX_EXinst_Maddsub__n0012_inst_lut3_17),
    .O(\DLX_EXinst__n0012<14>/CYMUXG )
  );
  X_XOR2 DLX_EXinst_Maddsub__n0012_inst_sum_85 (
    .I0(DLX_EXinst_Maddsub__n0012_inst_cy_84),
    .I1(DLX_EXinst_Maddsub__n0012_inst_lut3_17),
    .O(\DLX_EXinst__n0012<14>/XORG )
  );
  X_BUF \DLX_EXinst__n0012<14>/CYINIT_2470  (
    .I(DLX_EXinst_Maddsub__n0012_inst_cy_83),
    .O(\DLX_EXinst__n0012<14>/CYINIT )
  );
  X_MUX2 DLX_EXinst_Maddsub__n0012_inst_cy_86_2471 (
    .IA(DLX_IDinst_reg_out_A[16]),
    .IB(\DLX_IDinst_RegFile_18_5/CYINIT ),
    .SEL(DLX_EXinst_Maddsub__n0012_inst_lut3_18),
    .O(DLX_EXinst_Maddsub__n0012_inst_cy_86)
  );
  X_XOR2 DLX_EXinst_Maddsub__n0012_inst_sum_86 (
    .I0(\DLX_IDinst_RegFile_18_5/CYINIT ),
    .I1(DLX_EXinst_Maddsub__n0012_inst_lut3_18),
    .O(\DLX_IDinst_RegFile_18_5/XORF )
  );
  defparam DLX_EXinst_Maddsub__n0012_inst_lut3_181.INIT = 16'hA55A;
  X_LUT4 DLX_EXinst_Maddsub__n0012_inst_lut3_181 (
    .ADR0(DLX_IDinst_reg_out_A[16]),
    .ADR1(VCC),
    .ADR2(N144912),
    .ADR3(DLX_EXinst__n0013[16]),
    .O(DLX_EXinst_Maddsub__n0012_inst_lut3_18)
  );
  defparam DLX_EXinst_Maddsub__n0012_inst_lut3_191.INIT = 16'hA55A;
  X_LUT4 DLX_EXinst_Maddsub__n0012_inst_lut3_191 (
    .ADR0(DLX_IDinst_reg_out_A[17]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst__n0013[17]),
    .ADR3(N144912),
    .O(DLX_EXinst_Maddsub__n0012_inst_lut3_19)
  );
  X_BUF \DLX_IDinst_RegFile_18_5/COUTUSED  (
    .I(\DLX_IDinst_RegFile_18_5/CYMUXG ),
    .O(DLX_EXinst_Maddsub__n0012_inst_cy_87)
  );
  X_BUF \DLX_IDinst_RegFile_18_5/XUSED  (
    .I(\DLX_IDinst_RegFile_18_5/XORF ),
    .O(DLX_EXinst__n0012[16])
  );
  X_BUF \DLX_IDinst_RegFile_18_5/YUSED  (
    .I(\DLX_IDinst_RegFile_18_5/XORG ),
    .O(DLX_EXinst__n0012[17])
  );
  X_MUX2 DLX_EXinst_Maddsub__n0012_inst_cy_87_2472 (
    .IA(DLX_IDinst_reg_out_A[17]),
    .IB(DLX_EXinst_Maddsub__n0012_inst_cy_86),
    .SEL(DLX_EXinst_Maddsub__n0012_inst_lut3_19),
    .O(\DLX_IDinst_RegFile_18_5/CYMUXG )
  );
  X_XOR2 DLX_EXinst_Maddsub__n0012_inst_sum_87 (
    .I0(DLX_EXinst_Maddsub__n0012_inst_cy_86),
    .I1(DLX_EXinst_Maddsub__n0012_inst_lut3_19),
    .O(\DLX_IDinst_RegFile_18_5/XORG )
  );
  X_BUF \DLX_IDinst_RegFile_18_5/CYINIT_2473  (
    .I(DLX_EXinst_Maddsub__n0012_inst_cy_85),
    .O(\DLX_IDinst_RegFile_18_5/CYINIT )
  );
  X_MUX2 DLX_EXinst_Maddsub__n0012_inst_cy_88_2474 (
    .IA(DLX_IDinst_reg_out_A[18]),
    .IB(\DLX_EXinst__n0012<18>/CYINIT ),
    .SEL(DLX_EXinst_Maddsub__n0012_inst_lut3_20),
    .O(DLX_EXinst_Maddsub__n0012_inst_cy_88)
  );
  X_XOR2 DLX_EXinst_Maddsub__n0012_inst_sum_88 (
    .I0(\DLX_EXinst__n0012<18>/CYINIT ),
    .I1(DLX_EXinst_Maddsub__n0012_inst_lut3_20),
    .O(\DLX_EXinst__n0012<18>/XORF )
  );
  defparam DLX_EXinst_Maddsub__n0012_inst_lut3_201.INIT = 16'h9696;
  X_LUT4 DLX_EXinst_Maddsub__n0012_inst_lut3_201 (
    .ADR0(DLX_IDinst_reg_out_A[18]),
    .ADR1(DLX_EXinst__n0013[18]),
    .ADR2(N144912),
    .ADR3(VCC),
    .O(DLX_EXinst_Maddsub__n0012_inst_lut3_20)
  );
  defparam DLX_EXinst_Maddsub__n0012_inst_lut3_211.INIT = 16'hA55A;
  X_LUT4 DLX_EXinst_Maddsub__n0012_inst_lut3_211 (
    .ADR0(DLX_IDinst_reg_out_A[19]),
    .ADR1(VCC),
    .ADR2(N144912),
    .ADR3(DLX_EXinst__n0013[19]),
    .O(DLX_EXinst_Maddsub__n0012_inst_lut3_21)
  );
  X_BUF \DLX_EXinst__n0012<18>/COUTUSED  (
    .I(\DLX_EXinst__n0012<18>/CYMUXG ),
    .O(DLX_EXinst_Maddsub__n0012_inst_cy_89)
  );
  X_BUF \DLX_EXinst__n0012<18>/XUSED  (
    .I(\DLX_EXinst__n0012<18>/XORF ),
    .O(DLX_EXinst__n0012[18])
  );
  X_BUF \DLX_EXinst__n0012<18>/YUSED  (
    .I(\DLX_EXinst__n0012<18>/XORG ),
    .O(DLX_EXinst__n0012[19])
  );
  X_MUX2 DLX_EXinst_Maddsub__n0012_inst_cy_89_2475 (
    .IA(DLX_IDinst_reg_out_A[19]),
    .IB(DLX_EXinst_Maddsub__n0012_inst_cy_88),
    .SEL(DLX_EXinst_Maddsub__n0012_inst_lut3_21),
    .O(\DLX_EXinst__n0012<18>/CYMUXG )
  );
  X_XOR2 DLX_EXinst_Maddsub__n0012_inst_sum_89 (
    .I0(DLX_EXinst_Maddsub__n0012_inst_cy_88),
    .I1(DLX_EXinst_Maddsub__n0012_inst_lut3_21),
    .O(\DLX_EXinst__n0012<18>/XORG )
  );
  X_BUF \DLX_EXinst__n0012<18>/CYINIT_2476  (
    .I(DLX_EXinst_Maddsub__n0012_inst_cy_87),
    .O(\DLX_EXinst__n0012<18>/CYINIT )
  );
  X_MUX2 DLX_EXinst_Maddsub__n0012_inst_cy_90_2477 (
    .IA(DLX_IDinst_reg_out_A[20]),
    .IB(\DLX_EXinst__n0012<20>/CYINIT ),
    .SEL(DLX_EXinst_Maddsub__n0012_inst_lut3_22),
    .O(DLX_EXinst_Maddsub__n0012_inst_cy_90)
  );
  X_XOR2 DLX_EXinst_Maddsub__n0012_inst_sum_90 (
    .I0(\DLX_EXinst__n0012<20>/CYINIT ),
    .I1(DLX_EXinst_Maddsub__n0012_inst_lut3_22),
    .O(\DLX_EXinst__n0012<20>/XORF )
  );
  defparam DLX_EXinst_Maddsub__n0012_inst_lut3_221.INIT = 16'h9696;
  X_LUT4 DLX_EXinst_Maddsub__n0012_inst_lut3_221 (
    .ADR0(DLX_IDinst_reg_out_A[20]),
    .ADR1(DLX_EXinst__n0013[20]),
    .ADR2(N144912),
    .ADR3(VCC),
    .O(DLX_EXinst_Maddsub__n0012_inst_lut3_22)
  );
  defparam DLX_EXinst_Maddsub__n0012_inst_lut3_231.INIT = 16'hA55A;
  X_LUT4 DLX_EXinst_Maddsub__n0012_inst_lut3_231 (
    .ADR0(DLX_IDinst_reg_out_A[21]),
    .ADR1(VCC),
    .ADR2(N144912),
    .ADR3(DLX_EXinst__n0013[21]),
    .O(DLX_EXinst_Maddsub__n0012_inst_lut3_23)
  );
  X_BUF \DLX_EXinst__n0012<20>/COUTUSED  (
    .I(\DLX_EXinst__n0012<20>/CYMUXG ),
    .O(DLX_EXinst_Maddsub__n0012_inst_cy_91)
  );
  X_BUF \DLX_EXinst__n0012<20>/XUSED  (
    .I(\DLX_EXinst__n0012<20>/XORF ),
    .O(DLX_EXinst__n0012[20])
  );
  X_BUF \DLX_EXinst__n0012<20>/YUSED  (
    .I(\DLX_EXinst__n0012<20>/XORG ),
    .O(DLX_EXinst__n0012[21])
  );
  X_MUX2 DLX_EXinst_Maddsub__n0012_inst_cy_91_2478 (
    .IA(DLX_IDinst_reg_out_A[21]),
    .IB(DLX_EXinst_Maddsub__n0012_inst_cy_90),
    .SEL(DLX_EXinst_Maddsub__n0012_inst_lut3_23),
    .O(\DLX_EXinst__n0012<20>/CYMUXG )
  );
  X_XOR2 DLX_EXinst_Maddsub__n0012_inst_sum_91 (
    .I0(DLX_EXinst_Maddsub__n0012_inst_cy_90),
    .I1(DLX_EXinst_Maddsub__n0012_inst_lut3_23),
    .O(\DLX_EXinst__n0012<20>/XORG )
  );
  X_BUF \DLX_EXinst__n0012<20>/CYINIT_2479  (
    .I(DLX_EXinst_Maddsub__n0012_inst_cy_89),
    .O(\DLX_EXinst__n0012<20>/CYINIT )
  );
  X_MUX2 DLX_EXinst_Maddsub__n0012_inst_cy_92_2480 (
    .IA(DLX_IDinst_reg_out_A[22]),
    .IB(\DLX_EXinst__n0012<22>/CYINIT ),
    .SEL(DLX_EXinst_Maddsub__n0012_inst_lut3_24),
    .O(DLX_EXinst_Maddsub__n0012_inst_cy_92)
  );
  X_XOR2 DLX_EXinst_Maddsub__n0012_inst_sum_92 (
    .I0(\DLX_EXinst__n0012<22>/CYINIT ),
    .I1(DLX_EXinst_Maddsub__n0012_inst_lut3_24),
    .O(\DLX_EXinst__n0012<22>/XORF )
  );
  defparam DLX_EXinst_Maddsub__n0012_inst_lut3_241.INIT = 16'h9966;
  X_LUT4 DLX_EXinst_Maddsub__n0012_inst_lut3_241 (
    .ADR0(DLX_IDinst_reg_out_A[22]),
    .ADR1(DLX_EXinst__n0013[22]),
    .ADR2(VCC),
    .ADR3(N144912),
    .O(DLX_EXinst_Maddsub__n0012_inst_lut3_24)
  );
  defparam DLX_EXinst_Maddsub__n0012_inst_lut3_251.INIT = 16'h9966;
  X_LUT4 DLX_EXinst_Maddsub__n0012_inst_lut3_251 (
    .ADR0(DLX_IDinst_reg_out_A[23]),
    .ADR1(DLX_EXinst__n0013[23]),
    .ADR2(VCC),
    .ADR3(N144912),
    .O(DLX_EXinst_Maddsub__n0012_inst_lut3_25)
  );
  X_BUF \DLX_EXinst__n0012<22>/COUTUSED  (
    .I(\DLX_EXinst__n0012<22>/CYMUXG ),
    .O(DLX_EXinst_Maddsub__n0012_inst_cy_93)
  );
  X_BUF \DLX_EXinst__n0012<22>/XUSED  (
    .I(\DLX_EXinst__n0012<22>/XORF ),
    .O(DLX_EXinst__n0012[22])
  );
  X_BUF \DLX_EXinst__n0012<22>/YUSED  (
    .I(\DLX_EXinst__n0012<22>/XORG ),
    .O(DLX_EXinst__n0012[23])
  );
  X_MUX2 DLX_EXinst_Maddsub__n0012_inst_cy_93_2481 (
    .IA(DLX_IDinst_reg_out_A[23]),
    .IB(DLX_EXinst_Maddsub__n0012_inst_cy_92),
    .SEL(DLX_EXinst_Maddsub__n0012_inst_lut3_25),
    .O(\DLX_EXinst__n0012<22>/CYMUXG )
  );
  X_XOR2 DLX_EXinst_Maddsub__n0012_inst_sum_93 (
    .I0(DLX_EXinst_Maddsub__n0012_inst_cy_92),
    .I1(DLX_EXinst_Maddsub__n0012_inst_lut3_25),
    .O(\DLX_EXinst__n0012<22>/XORG )
  );
  X_BUF \DLX_EXinst__n0012<22>/CYINIT_2482  (
    .I(DLX_EXinst_Maddsub__n0012_inst_cy_91),
    .O(\DLX_EXinst__n0012<22>/CYINIT )
  );
  defparam DLX_IDinst_RegFile_29_25_2483.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_29_25_2483 (
    .I(DLX_IDinst_WB_data_eff[25]),
    .CE(DLX_IDinst__n0608),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_29_25)
  );
  X_MUX2 DLX_EXinst_Maddsub__n0012_inst_cy_94_2484 (
    .IA(DLX_IDinst_reg_out_A[24]),
    .IB(\DLX_IDinst_EPC<29>/CYINIT ),
    .SEL(DLX_EXinst_Maddsub__n0012_inst_lut3_26),
    .O(DLX_EXinst_Maddsub__n0012_inst_cy_94)
  );
  X_XOR2 DLX_EXinst_Maddsub__n0012_inst_sum_94 (
    .I0(\DLX_IDinst_EPC<29>/CYINIT ),
    .I1(DLX_EXinst_Maddsub__n0012_inst_lut3_26),
    .O(\DLX_IDinst_EPC<29>/XORF )
  );
  defparam DLX_EXinst_Maddsub__n0012_inst_lut3_261.INIT = 16'h9696;
  X_LUT4 DLX_EXinst_Maddsub__n0012_inst_lut3_261 (
    .ADR0(DLX_IDinst_reg_out_A[24]),
    .ADR1(N144912),
    .ADR2(DLX_EXinst__n0013[24]),
    .ADR3(VCC),
    .O(DLX_EXinst_Maddsub__n0012_inst_lut3_26)
  );
  defparam DLX_EXinst_Maddsub__n0012_inst_lut3_271.INIT = 16'hA55A;
  X_LUT4 DLX_EXinst_Maddsub__n0012_inst_lut3_271 (
    .ADR0(DLX_IDinst_reg_out_A[25]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst__n0013[25]),
    .ADR3(N144912),
    .O(DLX_EXinst_Maddsub__n0012_inst_lut3_27)
  );
  X_BUF \DLX_IDinst_EPC<29>/COUTUSED  (
    .I(\DLX_IDinst_EPC<29>/CYMUXG ),
    .O(DLX_EXinst_Maddsub__n0012_inst_cy_95)
  );
  X_BUF \DLX_IDinst_EPC<29>/XUSED  (
    .I(\DLX_IDinst_EPC<29>/XORF ),
    .O(DLX_EXinst__n0012[24])
  );
  X_BUF \DLX_IDinst_EPC<29>/YUSED  (
    .I(\DLX_IDinst_EPC<29>/XORG ),
    .O(DLX_EXinst__n0012[25])
  );
  X_MUX2 DLX_EXinst_Maddsub__n0012_inst_cy_95_2485 (
    .IA(DLX_IDinst_reg_out_A[25]),
    .IB(DLX_EXinst_Maddsub__n0012_inst_cy_94),
    .SEL(DLX_EXinst_Maddsub__n0012_inst_lut3_27),
    .O(\DLX_IDinst_EPC<29>/CYMUXG )
  );
  X_XOR2 DLX_EXinst_Maddsub__n0012_inst_sum_95 (
    .I0(DLX_EXinst_Maddsub__n0012_inst_cy_94),
    .I1(DLX_EXinst_Maddsub__n0012_inst_lut3_27),
    .O(\DLX_IDinst_EPC<29>/XORG )
  );
  X_BUF \DLX_IDinst_EPC<29>/CYINIT_2486  (
    .I(DLX_EXinst_Maddsub__n0012_inst_cy_93),
    .O(\DLX_IDinst_EPC<29>/CYINIT )
  );
  X_MUX2 DLX_EXinst_Maddsub__n0012_inst_cy_96_2487 (
    .IA(DLX_IDinst_reg_out_A[26]),
    .IB(\DLX_EXinst__n0012<26>/CYINIT ),
    .SEL(DLX_EXinst_Maddsub__n0012_inst_lut3_28),
    .O(DLX_EXinst_Maddsub__n0012_inst_cy_96)
  );
  X_XOR2 DLX_EXinst_Maddsub__n0012_inst_sum_96 (
    .I0(\DLX_EXinst__n0012<26>/CYINIT ),
    .I1(DLX_EXinst_Maddsub__n0012_inst_lut3_28),
    .O(\DLX_EXinst__n0012<26>/XORF )
  );
  defparam DLX_EXinst_Maddsub__n0012_inst_lut3_281.INIT = 16'h9966;
  X_LUT4 DLX_EXinst_Maddsub__n0012_inst_lut3_281 (
    .ADR0(DLX_IDinst_reg_out_A[26]),
    .ADR1(DLX_EXinst__n0013[26]),
    .ADR2(VCC),
    .ADR3(N144912),
    .O(DLX_EXinst_Maddsub__n0012_inst_lut3_28)
  );
  defparam DLX_EXinst_Maddsub__n0012_inst_lut3_291.INIT = 16'h9696;
  X_LUT4 DLX_EXinst_Maddsub__n0012_inst_lut3_291 (
    .ADR0(DLX_IDinst_reg_out_A[27]),
    .ADR1(N144912),
    .ADR2(DLX_EXinst__n0013[27]),
    .ADR3(VCC),
    .O(DLX_EXinst_Maddsub__n0012_inst_lut3_29)
  );
  X_BUF \DLX_EXinst__n0012<26>/COUTUSED  (
    .I(\DLX_EXinst__n0012<26>/CYMUXG ),
    .O(DLX_EXinst_Maddsub__n0012_inst_cy_97)
  );
  X_BUF \DLX_EXinst__n0012<26>/XUSED  (
    .I(\DLX_EXinst__n0012<26>/XORF ),
    .O(DLX_EXinst__n0012[26])
  );
  X_BUF \DLX_EXinst__n0012<26>/YUSED  (
    .I(\DLX_EXinst__n0012<26>/XORG ),
    .O(DLX_EXinst__n0012[27])
  );
  X_MUX2 DLX_EXinst_Maddsub__n0012_inst_cy_97_2488 (
    .IA(DLX_IDinst_reg_out_A[27]),
    .IB(DLX_EXinst_Maddsub__n0012_inst_cy_96),
    .SEL(DLX_EXinst_Maddsub__n0012_inst_lut3_29),
    .O(\DLX_EXinst__n0012<26>/CYMUXG )
  );
  X_XOR2 DLX_EXinst_Maddsub__n0012_inst_sum_97 (
    .I0(DLX_EXinst_Maddsub__n0012_inst_cy_96),
    .I1(DLX_EXinst_Maddsub__n0012_inst_lut3_29),
    .O(\DLX_EXinst__n0012<26>/XORG )
  );
  X_BUF \DLX_EXinst__n0012<26>/CYINIT_2489  (
    .I(DLX_EXinst_Maddsub__n0012_inst_cy_95),
    .O(\DLX_EXinst__n0012<26>/CYINIT )
  );
  X_MUX2 DLX_EXinst_Maddsub__n0012_inst_cy_98_2490 (
    .IA(DLX_IDinst_reg_out_A[28]),
    .IB(\DLX_EXinst__n0012<28>/CYINIT ),
    .SEL(DLX_EXinst_Maddsub__n0012_inst_lut3_30),
    .O(DLX_EXinst_Maddsub__n0012_inst_cy_98)
  );
  X_XOR2 DLX_EXinst_Maddsub__n0012_inst_sum_98 (
    .I0(\DLX_EXinst__n0012<28>/CYINIT ),
    .I1(DLX_EXinst_Maddsub__n0012_inst_lut3_30),
    .O(\DLX_EXinst__n0012<28>/XORF )
  );
  defparam DLX_EXinst_Maddsub__n0012_inst_lut3_301.INIT = 16'hA55A;
  X_LUT4 DLX_EXinst_Maddsub__n0012_inst_lut3_301 (
    .ADR0(DLX_IDinst_reg_out_A[28]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst__n0013[28]),
    .ADR3(N144912),
    .O(DLX_EXinst_Maddsub__n0012_inst_lut3_30)
  );
  defparam DLX_EXinst_Maddsub__n0012_inst_lut3_311.INIT = 16'hA55A;
  X_LUT4 DLX_EXinst_Maddsub__n0012_inst_lut3_311 (
    .ADR0(DLX_IDinst_reg_out_A[29]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst__n0013[29]),
    .ADR3(N144912),
    .O(DLX_EXinst_Maddsub__n0012_inst_lut3_31)
  );
  X_BUF \DLX_EXinst__n0012<28>/COUTUSED  (
    .I(\DLX_EXinst__n0012<28>/CYMUXG ),
    .O(DLX_EXinst_Maddsub__n0012_inst_cy_99)
  );
  X_BUF \DLX_EXinst__n0012<28>/XUSED  (
    .I(\DLX_EXinst__n0012<28>/XORF ),
    .O(DLX_EXinst__n0012[28])
  );
  X_BUF \DLX_EXinst__n0012<28>/YUSED  (
    .I(\DLX_EXinst__n0012<28>/XORG ),
    .O(DLX_EXinst__n0012[29])
  );
  X_MUX2 DLX_EXinst_Maddsub__n0012_inst_cy_99_2491 (
    .IA(DLX_IDinst_reg_out_A[29]),
    .IB(DLX_EXinst_Maddsub__n0012_inst_cy_98),
    .SEL(DLX_EXinst_Maddsub__n0012_inst_lut3_31),
    .O(\DLX_EXinst__n0012<28>/CYMUXG )
  );
  X_XOR2 DLX_EXinst_Maddsub__n0012_inst_sum_99 (
    .I0(DLX_EXinst_Maddsub__n0012_inst_cy_98),
    .I1(DLX_EXinst_Maddsub__n0012_inst_lut3_31),
    .O(\DLX_EXinst__n0012<28>/XORG )
  );
  X_BUF \DLX_EXinst__n0012<28>/CYINIT_2492  (
    .I(DLX_EXinst_Maddsub__n0012_inst_cy_97),
    .O(\DLX_EXinst__n0012<28>/CYINIT )
  );
  X_MUX2 DLX_EXinst_Maddsub__n0012_inst_cy_100_2493 (
    .IA(DLX_IDinst_reg_out_A[30]),
    .IB(\DLX_EXinst__n0012<30>/CYINIT ),
    .SEL(DLX_EXinst_Maddsub__n0012_inst_lut3_32),
    .O(DLX_EXinst_Maddsub__n0012_inst_cy_100)
  );
  X_XOR2 DLX_EXinst_Maddsub__n0012_inst_sum_100 (
    .I0(\DLX_EXinst__n0012<30>/CYINIT ),
    .I1(DLX_EXinst_Maddsub__n0012_inst_lut3_32),
    .O(\DLX_EXinst__n0012<30>/XORF )
  );
  defparam DLX_EXinst_Maddsub__n0012_inst_lut3_321.INIT = 16'h9966;
  X_LUT4 DLX_EXinst_Maddsub__n0012_inst_lut3_321 (
    .ADR0(DLX_IDinst_reg_out_A[30]),
    .ADR1(N144912),
    .ADR2(VCC),
    .ADR3(DLX_EXinst__n0013[30]),
    .O(DLX_EXinst_Maddsub__n0012_inst_lut3_32)
  );
  defparam DLX_EXinst_Maddsub__n0012_inst_lut3_331.INIT = 16'h9966;
  X_LUT4 DLX_EXinst_Maddsub__n0012_inst_lut3_331 (
    .ADR0(DLX_IDinst_reg_out_A[31]),
    .ADR1(DLX_EXinst__n0013[31]),
    .ADR2(VCC),
    .ADR3(N144912),
    .O(DLX_EXinst_Maddsub__n0012_inst_lut3_33)
  );
  X_BUF \DLX_EXinst__n0012<30>/XUSED  (
    .I(\DLX_EXinst__n0012<30>/XORF ),
    .O(DLX_EXinst__n0012[30])
  );
  X_BUF \DLX_EXinst__n0012<30>/YUSED  (
    .I(\DLX_EXinst__n0012<30>/XORG ),
    .O(DLX_EXinst__n0012[31])
  );
  X_XOR2 DLX_EXinst_Maddsub__n0012_inst_sum_101 (
    .I0(DLX_EXinst_Maddsub__n0012_inst_cy_100),
    .I1(DLX_EXinst_Maddsub__n0012_inst_lut3_33),
    .O(\DLX_EXinst__n0012<30>/XORG )
  );
  X_BUF \DLX_EXinst__n0012<30>/CYINIT_2494  (
    .I(DLX_EXinst_Maddsub__n0012_inst_cy_99),
    .O(\DLX_EXinst__n0012<30>/CYINIT )
  );
  X_ZERO \DLX_EXinst_Mcompar__n0087_inst_cy_119/LOGIC_ZERO_2495  (
    .O(\DLX_EXinst_Mcompar__n0087_inst_cy_119/LOGIC_ZERO )
  );
  X_ONE \DLX_EXinst_Mcompar__n0087_inst_cy_119/LOGIC_ONE_2496  (
    .O(\DLX_EXinst_Mcompar__n0087_inst_cy_119/LOGIC_ONE )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0087_inst_cy_118_2497 (
    .IA(\DLX_EXinst_Mcompar__n0087_inst_cy_119/LOGIC_ONE ),
    .IB(\DLX_EXinst_Mcompar__n0087_inst_cy_119/LOGIC_ZERO ),
    .SEL(DLX_EXinst_Mcompar__n0087_inst_lut4_16),
    .O(DLX_EXinst_Mcompar__n0087_inst_cy_118)
  );
  defparam DLX_EXinst_Mcompar__n0087_inst_lut4_161.INIT = 16'h8421;
  X_LUT4 DLX_EXinst_Mcompar__n0087_inst_lut4_161 (
    .ADR0(DLX_IDinst_reg_out_A[1]),
    .ADR1(DLX_IDinst_reg_out_B[0]),
    .ADR2(DLX_IDinst_reg_out_B[1]),
    .ADR3(DLX_IDinst_reg_out_A[0]),
    .O(DLX_EXinst_Mcompar__n0087_inst_lut4_16)
  );
  defparam DLX_EXinst_Mcompar__n0087_inst_lut4_171.INIT = 16'h9009;
  X_LUT4 DLX_EXinst_Mcompar__n0087_inst_lut4_171 (
    .ADR0(DLX_IDinst_reg_out_B_3_1),
    .ADR1(DLX_IDinst_reg_out_A[3]),
    .ADR2(DLX_IDinst_reg_out_B_2_1),
    .ADR3(DLX_IDinst_reg_out_A[2]),
    .O(DLX_EXinst_Mcompar__n0087_inst_lut4_17)
  );
  X_BUF \DLX_EXinst_Mcompar__n0087_inst_cy_119/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0087_inst_cy_119/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0087_inst_cy_119)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0087_inst_cy_119_2498 (
    .IA(\DLX_EXinst_Mcompar__n0087_inst_cy_119/LOGIC_ONE ),
    .IB(DLX_EXinst_Mcompar__n0087_inst_cy_118),
    .SEL(DLX_EXinst_Mcompar__n0087_inst_lut4_17),
    .O(\DLX_EXinst_Mcompar__n0087_inst_cy_119/CYMUXG )
  );
  X_ONE \DLX_EXinst_Mcompar__n0087_inst_cy_121/LOGIC_ONE_2499  (
    .O(\DLX_EXinst_Mcompar__n0087_inst_cy_121/LOGIC_ONE )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0087_inst_cy_120_2500 (
    .IA(\DLX_EXinst_Mcompar__n0087_inst_cy_121/LOGIC_ONE ),
    .IB(\DLX_EXinst_Mcompar__n0087_inst_cy_121/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0087_inst_lut4_18),
    .O(DLX_EXinst_Mcompar__n0087_inst_cy_120)
  );
  defparam DLX_EXinst_Mcompar__n0087_inst_lut4_181.INIT = 16'h8421;
  X_LUT4 DLX_EXinst_Mcompar__n0087_inst_lut4_181 (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(DLX_IDinst_reg_out_B[5]),
    .ADR2(DLX_IDinst_reg_out_A[4]),
    .ADR3(DLX_IDinst_reg_out_A[5]),
    .O(DLX_EXinst_Mcompar__n0087_inst_lut4_18)
  );
  defparam DLX_EXinst_Mcompar__n0087_inst_lut4_191.INIT = 16'h8241;
  X_LUT4 DLX_EXinst_Mcompar__n0087_inst_lut4_191 (
    .ADR0(DLX_IDinst_reg_out_A[7]),
    .ADR1(DLX_IDinst_reg_out_B[6]),
    .ADR2(DLX_IDinst_reg_out_A[6]),
    .ADR3(DLX_IDinst_reg_out_B[7]),
    .O(DLX_EXinst_Mcompar__n0087_inst_lut4_19)
  );
  X_BUF \DLX_EXinst_Mcompar__n0087_inst_cy_121/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0087_inst_cy_121/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0087_inst_cy_121)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0087_inst_cy_121_2501 (
    .IA(\DLX_EXinst_Mcompar__n0087_inst_cy_121/LOGIC_ONE ),
    .IB(DLX_EXinst_Mcompar__n0087_inst_cy_120),
    .SEL(DLX_EXinst_Mcompar__n0087_inst_lut4_19),
    .O(\DLX_EXinst_Mcompar__n0087_inst_cy_121/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0087_inst_cy_121/CYINIT_2502  (
    .I(DLX_EXinst_Mcompar__n0087_inst_cy_119),
    .O(\DLX_EXinst_Mcompar__n0087_inst_cy_121/CYINIT )
  );
  defparam DLX_IDinst_RegFile_29_17_2503.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_29_17_2503 (
    .I(DLX_IDinst_WB_data_eff[17]),
    .CE(DLX_IDinst__n0608),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_29_17)
  );
  X_ONE \DLX_EXinst_Mcompar__n0087_inst_cy_123/LOGIC_ONE_2504  (
    .O(\DLX_EXinst_Mcompar__n0087_inst_cy_123/LOGIC_ONE )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0087_inst_cy_122_2505 (
    .IA(\DLX_EXinst_Mcompar__n0087_inst_cy_123/LOGIC_ONE ),
    .IB(\DLX_EXinst_Mcompar__n0087_inst_cy_123/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0087_inst_lut4_20),
    .O(DLX_EXinst_Mcompar__n0087_inst_cy_122)
  );
  defparam DLX_EXinst_Mcompar__n0087_inst_lut4_201.INIT = 16'h9009;
  X_LUT4 DLX_EXinst_Mcompar__n0087_inst_lut4_201 (
    .ADR0(DLX_IDinst_reg_out_B[8]),
    .ADR1(DLX_IDinst_reg_out_A[8]),
    .ADR2(DLX_IDinst_reg_out_B[9]),
    .ADR3(DLX_IDinst_reg_out_A[9]),
    .O(DLX_EXinst_Mcompar__n0087_inst_lut4_20)
  );
  defparam DLX_EXinst_Mcompar__n0087_inst_lut4_211.INIT = 16'h9009;
  X_LUT4 DLX_EXinst_Mcompar__n0087_inst_lut4_211 (
    .ADR0(DLX_IDinst_reg_out_A[11]),
    .ADR1(DLX_IDinst_reg_out_B[11]),
    .ADR2(DLX_IDinst_reg_out_A[10]),
    .ADR3(DLX_IDinst_reg_out_B[10]),
    .O(DLX_EXinst_Mcompar__n0087_inst_lut4_21)
  );
  X_BUF \DLX_EXinst_Mcompar__n0087_inst_cy_123/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0087_inst_cy_123/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0087_inst_cy_123)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0087_inst_cy_123_2506 (
    .IA(\DLX_EXinst_Mcompar__n0087_inst_cy_123/LOGIC_ONE ),
    .IB(DLX_EXinst_Mcompar__n0087_inst_cy_122),
    .SEL(DLX_EXinst_Mcompar__n0087_inst_lut4_21),
    .O(\DLX_EXinst_Mcompar__n0087_inst_cy_123/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0087_inst_cy_123/CYINIT_2507  (
    .I(DLX_EXinst_Mcompar__n0087_inst_cy_121),
    .O(\DLX_EXinst_Mcompar__n0087_inst_cy_123/CYINIT )
  );
  X_ONE \DLX_EXinst_Mcompar__n0087_inst_cy_125/LOGIC_ONE_2508  (
    .O(\DLX_EXinst_Mcompar__n0087_inst_cy_125/LOGIC_ONE )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0087_inst_cy_124_2509 (
    .IA(\DLX_EXinst_Mcompar__n0087_inst_cy_125/LOGIC_ONE ),
    .IB(\DLX_EXinst_Mcompar__n0087_inst_cy_125/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0087_inst_lut4_22),
    .O(DLX_EXinst_Mcompar__n0087_inst_cy_124)
  );
  defparam DLX_EXinst_Mcompar__n0087_inst_lut4_221.INIT = 16'h8241;
  X_LUT4 DLX_EXinst_Mcompar__n0087_inst_lut4_221 (
    .ADR0(DLX_IDinst_reg_out_A[13]),
    .ADR1(DLX_IDinst_reg_out_B[12]),
    .ADR2(DLX_IDinst_reg_out_A[12]),
    .ADR3(DLX_IDinst_reg_out_B[13]),
    .O(DLX_EXinst_Mcompar__n0087_inst_lut4_22)
  );
  defparam DLX_EXinst_Mcompar__n0087_inst_lut4_231.INIT = 16'h8241;
  X_LUT4 DLX_EXinst_Mcompar__n0087_inst_lut4_231 (
    .ADR0(DLX_IDinst_reg_out_A[14]),
    .ADR1(DLX_IDinst_reg_out_A[15]),
    .ADR2(DLX_IDinst_reg_out_B[15]),
    .ADR3(DLX_IDinst_reg_out_B[14]),
    .O(DLX_EXinst_Mcompar__n0087_inst_lut4_23)
  );
  X_BUF \DLX_EXinst_Mcompar__n0087_inst_cy_125/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0087_inst_cy_125/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0087_inst_cy_125)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0087_inst_cy_125_2510 (
    .IA(\DLX_EXinst_Mcompar__n0087_inst_cy_125/LOGIC_ONE ),
    .IB(DLX_EXinst_Mcompar__n0087_inst_cy_124),
    .SEL(DLX_EXinst_Mcompar__n0087_inst_lut4_23),
    .O(\DLX_EXinst_Mcompar__n0087_inst_cy_125/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0087_inst_cy_125/CYINIT_2511  (
    .I(DLX_EXinst_Mcompar__n0087_inst_cy_123),
    .O(\DLX_EXinst_Mcompar__n0087_inst_cy_125/CYINIT )
  );
  X_ONE \DLX_EXinst_Mcompar__n0087_inst_cy_127/LOGIC_ONE_2512  (
    .O(\DLX_EXinst_Mcompar__n0087_inst_cy_127/LOGIC_ONE )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0087_inst_cy_126_2513 (
    .IA(\DLX_EXinst_Mcompar__n0087_inst_cy_127/LOGIC_ONE ),
    .IB(\DLX_EXinst_Mcompar__n0087_inst_cy_127/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0087_inst_lut4_24),
    .O(DLX_EXinst_Mcompar__n0087_inst_cy_126)
  );
  defparam DLX_EXinst_Mcompar__n0087_inst_lut4_241.INIT = 16'h9009;
  X_LUT4 DLX_EXinst_Mcompar__n0087_inst_lut4_241 (
    .ADR0(DLX_IDinst_reg_out_A[16]),
    .ADR1(DLX_IDinst_reg_out_B[16]),
    .ADR2(DLX_IDinst_reg_out_B[17]),
    .ADR3(DLX_IDinst_reg_out_A[17]),
    .O(DLX_EXinst_Mcompar__n0087_inst_lut4_24)
  );
  defparam DLX_EXinst_Mcompar__n0087_inst_lut4_251.INIT = 16'h8241;
  X_LUT4 DLX_EXinst_Mcompar__n0087_inst_lut4_251 (
    .ADR0(DLX_IDinst_reg_out_A[18]),
    .ADR1(DLX_IDinst_reg_out_B[19]),
    .ADR2(DLX_IDinst_reg_out_A[19]),
    .ADR3(DLX_IDinst_reg_out_B[18]),
    .O(DLX_EXinst_Mcompar__n0087_inst_lut4_25)
  );
  X_BUF \DLX_EXinst_Mcompar__n0087_inst_cy_127/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0087_inst_cy_127/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0087_inst_cy_127)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0087_inst_cy_127_2514 (
    .IA(\DLX_EXinst_Mcompar__n0087_inst_cy_127/LOGIC_ONE ),
    .IB(DLX_EXinst_Mcompar__n0087_inst_cy_126),
    .SEL(DLX_EXinst_Mcompar__n0087_inst_lut4_25),
    .O(\DLX_EXinst_Mcompar__n0087_inst_cy_127/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0087_inst_cy_127/CYINIT_2515  (
    .I(DLX_EXinst_Mcompar__n0087_inst_cy_125),
    .O(\DLX_EXinst_Mcompar__n0087_inst_cy_127/CYINIT )
  );
  X_ONE \DLX_EXinst_Mcompar__n0087_inst_cy_129/LOGIC_ONE_2516  (
    .O(\DLX_EXinst_Mcompar__n0087_inst_cy_129/LOGIC_ONE )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0087_inst_cy_128_2517 (
    .IA(\DLX_EXinst_Mcompar__n0087_inst_cy_129/LOGIC_ONE ),
    .IB(\DLX_EXinst_Mcompar__n0087_inst_cy_129/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0087_inst_lut4_26),
    .O(DLX_EXinst_Mcompar__n0087_inst_cy_128)
  );
  defparam DLX_EXinst_Mcompar__n0087_inst_lut4_261.INIT = 16'h8241;
  X_LUT4 DLX_EXinst_Mcompar__n0087_inst_lut4_261 (
    .ADR0(DLX_IDinst_reg_out_B[20]),
    .ADR1(DLX_IDinst_reg_out_B[21]),
    .ADR2(DLX_IDinst_reg_out_A[21]),
    .ADR3(DLX_IDinst_reg_out_A[20]),
    .O(DLX_EXinst_Mcompar__n0087_inst_lut4_26)
  );
  defparam DLX_EXinst_Mcompar__n0087_inst_lut4_271.INIT = 16'h8421;
  X_LUT4 DLX_EXinst_Mcompar__n0087_inst_lut4_271 (
    .ADR0(DLX_IDinst_reg_out_A[23]),
    .ADR1(DLX_IDinst_reg_out_A[22]),
    .ADR2(DLX_IDinst_reg_out_B[23]),
    .ADR3(DLX_IDinst_reg_out_B[22]),
    .O(DLX_EXinst_Mcompar__n0087_inst_lut4_27)
  );
  X_BUF \DLX_EXinst_Mcompar__n0087_inst_cy_129/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0087_inst_cy_129/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0087_inst_cy_129)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0087_inst_cy_129_2518 (
    .IA(\DLX_EXinst_Mcompar__n0087_inst_cy_129/LOGIC_ONE ),
    .IB(DLX_EXinst_Mcompar__n0087_inst_cy_128),
    .SEL(DLX_EXinst_Mcompar__n0087_inst_lut4_27),
    .O(\DLX_EXinst_Mcompar__n0087_inst_cy_129/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0087_inst_cy_129/CYINIT_2519  (
    .I(DLX_EXinst_Mcompar__n0087_inst_cy_127),
    .O(\DLX_EXinst_Mcompar__n0087_inst_cy_129/CYINIT )
  );
  X_ONE \DLX_EXinst_Mcompar__n0087_inst_cy_131/LOGIC_ONE_2520  (
    .O(\DLX_EXinst_Mcompar__n0087_inst_cy_131/LOGIC_ONE )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0087_inst_cy_130_2521 (
    .IA(\DLX_EXinst_Mcompar__n0087_inst_cy_131/LOGIC_ONE ),
    .IB(\DLX_EXinst_Mcompar__n0087_inst_cy_131/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0087_inst_lut4_28),
    .O(DLX_EXinst_Mcompar__n0087_inst_cy_130)
  );
  defparam DLX_EXinst_Mcompar__n0087_inst_lut4_281.INIT = 16'h8241;
  X_LUT4 DLX_EXinst_Mcompar__n0087_inst_lut4_281 (
    .ADR0(DLX_IDinst_reg_out_A[25]),
    .ADR1(DLX_IDinst_reg_out_A[24]),
    .ADR2(DLX_IDinst_reg_out_B[24]),
    .ADR3(DLX_IDinst_reg_out_B[25]),
    .O(DLX_EXinst_Mcompar__n0087_inst_lut4_28)
  );
  defparam DLX_EXinst_Mcompar__n0087_inst_lut4_291.INIT = 16'h8421;
  X_LUT4 DLX_EXinst_Mcompar__n0087_inst_lut4_291 (
    .ADR0(DLX_IDinst_reg_out_B[27]),
    .ADR1(DLX_IDinst_reg_out_B[26]),
    .ADR2(DLX_IDinst_reg_out_A[27]),
    .ADR3(DLX_IDinst_reg_out_A[26]),
    .O(DLX_EXinst_Mcompar__n0087_inst_lut4_29)
  );
  X_BUF \DLX_EXinst_Mcompar__n0087_inst_cy_131/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0087_inst_cy_131/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0087_inst_cy_131)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0087_inst_cy_131_2522 (
    .IA(\DLX_EXinst_Mcompar__n0087_inst_cy_131/LOGIC_ONE ),
    .IB(DLX_EXinst_Mcompar__n0087_inst_cy_130),
    .SEL(DLX_EXinst_Mcompar__n0087_inst_lut4_29),
    .O(\DLX_EXinst_Mcompar__n0087_inst_cy_131/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0087_inst_cy_131/CYINIT_2523  (
    .I(DLX_EXinst_Mcompar__n0087_inst_cy_129),
    .O(\DLX_EXinst_Mcompar__n0087_inst_cy_131/CYINIT )
  );
  X_ONE \DLX_EXinst__n0087/LOGIC_ONE_2524  (
    .O(\DLX_EXinst__n0087/LOGIC_ONE )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0087_inst_cy_132_2525 (
    .IA(\DLX_EXinst__n0087/LOGIC_ONE ),
    .IB(\DLX_EXinst__n0087/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0087_inst_lut4_30),
    .O(DLX_EXinst_Mcompar__n0087_inst_cy_132)
  );
  defparam DLX_EXinst_Mcompar__n0087_inst_lut4_301.INIT = 16'h9009;
  X_LUT4 DLX_EXinst_Mcompar__n0087_inst_lut4_301 (
    .ADR0(DLX_IDinst_reg_out_B[28]),
    .ADR1(DLX_IDinst_reg_out_A[28]),
    .ADR2(DLX_IDinst_reg_out_A[29]),
    .ADR3(DLX_IDinst_reg_out_B[29]),
    .O(DLX_EXinst_Mcompar__n0087_inst_lut4_30)
  );
  defparam DLX_EXinst_Mcompar__n0087_inst_lut4_311.INIT = 16'h8421;
  X_LUT4 DLX_EXinst_Mcompar__n0087_inst_lut4_311 (
    .ADR0(DLX_IDinst_reg_out_B[31]),
    .ADR1(DLX_IDinst_reg_out_A[30]),
    .ADR2(DLX_IDinst_reg_out_A[31]),
    .ADR3(DLX_IDinst_reg_out_B[30]),
    .O(DLX_EXinst_Mcompar__n0087_inst_lut4_31)
  );
  X_BUF \DLX_EXinst__n0087/COUTUSED  (
    .I(\DLX_EXinst__n0087/CYMUXG ),
    .O(DLX_EXinst__n0087)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0087_inst_cy_133 (
    .IA(\DLX_EXinst__n0087/LOGIC_ONE ),
    .IB(DLX_EXinst_Mcompar__n0087_inst_cy_132),
    .SEL(DLX_EXinst_Mcompar__n0087_inst_lut4_31),
    .O(\DLX_EXinst__n0087/CYMUXG )
  );
  X_BUF \DLX_EXinst__n0087/CYINIT_2526  (
    .I(DLX_EXinst_Mcompar__n0087_inst_cy_131),
    .O(\DLX_EXinst__n0087/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_2_25/LOGIC_ZERO_2527  (
    .O(\DLX_IDinst_RegFile_2_25/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_230_2528 (
    .IA(DLX_IDinst_reg_out_B[0]),
    .IB(\DLX_IDinst_RegFile_2_25/LOGIC_ZERO ),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_166),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_230)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1661.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1661 (
    .ADR0(DLX_IDinst_reg_out_B[0]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[0]),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_166)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1671.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1671 (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[1]),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_167)
  );
  X_BUF \DLX_IDinst_RegFile_2_25/COUTUSED  (
    .I(\DLX_IDinst_RegFile_2_25/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_231)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_231_2529 (
    .IA(DLX_IDinst_reg_out_B[1]),
    .IB(DLX_EXinst_Mcompar__n0095_inst_cy_230),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_167),
    .O(\DLX_IDinst_RegFile_2_25/CYMUXG )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_232_2530 (
    .IA(DLX_IDinst_reg_out_B_2_1),
    .IB(\DLX_EXinst_Mcompar__n0095_inst_cy_233/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_168),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_232)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1681.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1681 (
    .ADR0(DLX_IDinst_reg_out_B_2_1),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[2]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_168)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1691.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1691 (
    .ADR0(DLX_IDinst_reg_out_B_3_1),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[3]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_169)
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_233/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0095_inst_cy_233/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_233)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_233_2531 (
    .IA(DLX_IDinst_reg_out_B_3_1),
    .IB(DLX_EXinst_Mcompar__n0095_inst_cy_232),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_169),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_233/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_233/CYINIT_2532  (
    .I(DLX_EXinst_Mcompar__n0095_inst_cy_231),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_233/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_234_2533 (
    .IA(DLX_IDinst_reg_out_B[4]),
    .IB(\DLX_EXinst_Mcompar__n0095_inst_cy_235/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_170),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_234)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1701.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1701 (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[4]),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_170)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1711.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1711 (
    .ADR0(DLX_IDinst_reg_out_B[5]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[5]),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_171)
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_235/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0095_inst_cy_235/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_235)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_235_2534 (
    .IA(DLX_IDinst_reg_out_B[5]),
    .IB(DLX_EXinst_Mcompar__n0095_inst_cy_234),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_171),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_235/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_235/CYINIT_2535  (
    .I(DLX_EXinst_Mcompar__n0095_inst_cy_233),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_235/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_236_2536 (
    .IA(DLX_IDinst_reg_out_B[6]),
    .IB(\DLX_EXinst_Mcompar__n0095_inst_cy_237/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_172),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_236)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1721.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1721 (
    .ADR0(DLX_IDinst_reg_out_B[6]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[6]),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_172)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1731.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1731 (
    .ADR0(DLX_IDinst_reg_out_B[7]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[7]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_173)
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_237/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0095_inst_cy_237/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_237)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_237_2537 (
    .IA(DLX_IDinst_reg_out_B[7]),
    .IB(DLX_EXinst_Mcompar__n0095_inst_cy_236),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_173),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_237/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_237/CYINIT_2538  (
    .I(DLX_EXinst_Mcompar__n0095_inst_cy_235),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_237/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_238_2539 (
    .IA(DLX_IDinst_reg_out_B[8]),
    .IB(\DLX_IFinst_IR_curr<15>/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_174),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_238)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1741.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1741 (
    .ADR0(DLX_IDinst_reg_out_B[8]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[8]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_174)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1751.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1751 (
    .ADR0(DLX_IDinst_reg_out_B[9]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[9]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_175)
  );
  X_BUF \DLX_IFinst_IR_curr<15>/COUTUSED  (
    .I(\DLX_IFinst_IR_curr<15>/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_239)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_239_2540 (
    .IA(DLX_IDinst_reg_out_B[9]),
    .IB(DLX_EXinst_Mcompar__n0095_inst_cy_238),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_175),
    .O(\DLX_IFinst_IR_curr<15>/CYMUXG )
  );
  X_BUF \DLX_IFinst_IR_curr<15>/CYINIT_2541  (
    .I(DLX_EXinst_Mcompar__n0095_inst_cy_237),
    .O(\DLX_IFinst_IR_curr<15>/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_240_2542 (
    .IA(DLX_IDinst_reg_out_B[10]),
    .IB(\DLX_EXinst_Mcompar__n0095_inst_cy_241/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_176),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_240)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1761.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1761 (
    .ADR0(DLX_IDinst_reg_out_B[10]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[10]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_176)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1771.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1771 (
    .ADR0(DLX_IDinst_reg_out_B[11]),
    .ADR1(DLX_IDinst_reg_out_A[11]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_177)
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_241/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0095_inst_cy_241/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_241)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_241_2543 (
    .IA(DLX_IDinst_reg_out_B[11]),
    .IB(DLX_EXinst_Mcompar__n0095_inst_cy_240),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_177),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_241/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_241/CYINIT_2544  (
    .I(DLX_EXinst_Mcompar__n0095_inst_cy_239),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_241/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_242_2545 (
    .IA(DLX_IDinst_reg_out_B[12]),
    .IB(\DLX_EXinst_Mcompar__n0095_inst_cy_243/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_178),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_242)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1781.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1781 (
    .ADR0(DLX_IDinst_reg_out_B[12]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[12]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_178)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1791.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1791 (
    .ADR0(DLX_IDinst_reg_out_B[13]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[13]),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_179)
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_243/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0095_inst_cy_243/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_243)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_243_2546 (
    .IA(DLX_IDinst_reg_out_B[13]),
    .IB(DLX_EXinst_Mcompar__n0095_inst_cy_242),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_179),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_243/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_243/CYINIT_2547  (
    .I(DLX_EXinst_Mcompar__n0095_inst_cy_241),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_243/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_244_2548 (
    .IA(DLX_IDinst_reg_out_B[14]),
    .IB(\DLX_EXinst_Mcompar__n0095_inst_cy_245/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_180),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_244)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1801.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1801 (
    .ADR0(DLX_IDinst_reg_out_B[14]),
    .ADR1(DLX_IDinst_reg_out_A[14]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_180)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1811.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1811 (
    .ADR0(DLX_IDinst_reg_out_B[15]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[15]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_181)
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_245/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0095_inst_cy_245/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_245)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_245_2549 (
    .IA(DLX_IDinst_reg_out_B[15]),
    .IB(DLX_EXinst_Mcompar__n0095_inst_cy_244),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_181),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_245/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_245/CYINIT_2550  (
    .I(DLX_EXinst_Mcompar__n0095_inst_cy_243),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_245/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_246_2551 (
    .IA(DLX_IDinst_reg_out_B[16]),
    .IB(\DLX_IFinst_IR_curr<4>/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_182),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_246)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1821.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1821 (
    .ADR0(DLX_IDinst_reg_out_B[16]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[16]),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_182)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1831.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1831 (
    .ADR0(DLX_IDinst_reg_out_B[17]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[17]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_183)
  );
  X_BUF \DLX_IFinst_IR_curr<4>/COUTUSED  (
    .I(\DLX_IFinst_IR_curr<4>/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_247)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_247_2552 (
    .IA(DLX_IDinst_reg_out_B[17]),
    .IB(DLX_EXinst_Mcompar__n0095_inst_cy_246),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_183),
    .O(\DLX_IFinst_IR_curr<4>/CYMUXG )
  );
  X_BUF \DLX_IFinst_IR_curr<4>/CYINIT_2553  (
    .I(DLX_EXinst_Mcompar__n0095_inst_cy_245),
    .O(\DLX_IFinst_IR_curr<4>/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_248_2554 (
    .IA(DLX_IDinst_reg_out_B[18]),
    .IB(\DLX_EXinst_Mcompar__n0095_inst_cy_249/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_184),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_248)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1841.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1841 (
    .ADR0(DLX_IDinst_reg_out_B[18]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[18]),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_184)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1851.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1851 (
    .ADR0(DLX_IDinst_reg_out_B[19]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[19]),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_185)
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_249/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0095_inst_cy_249/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_249)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_249_2555 (
    .IA(DLX_IDinst_reg_out_B[19]),
    .IB(DLX_EXinst_Mcompar__n0095_inst_cy_248),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_185),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_249/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_249/CYINIT_2556  (
    .I(DLX_EXinst_Mcompar__n0095_inst_cy_247),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_249/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_250_2557 (
    .IA(DLX_IDinst_reg_out_B[20]),
    .IB(\DLX_EXinst_Mcompar__n0095_inst_cy_251/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_186),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_250)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1861.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1861 (
    .ADR0(DLX_IDinst_reg_out_B[20]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[20]),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_186)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1871.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1871 (
    .ADR0(DLX_IDinst_reg_out_B[21]),
    .ADR1(DLX_IDinst_reg_out_A[21]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_187)
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_251/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0095_inst_cy_251/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_251)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_251_2558 (
    .IA(DLX_IDinst_reg_out_B[21]),
    .IB(DLX_EXinst_Mcompar__n0095_inst_cy_250),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_187),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_251/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_251/CYINIT_2559  (
    .I(DLX_EXinst_Mcompar__n0095_inst_cy_249),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_251/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_252_2560 (
    .IA(DLX_IDinst_reg_out_B[22]),
    .IB(\DLX_EXinst_Mcompar__n0095_inst_cy_253/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_188),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_252)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1881.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1881 (
    .ADR0(DLX_IDinst_reg_out_B[22]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[22]),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_188)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1891.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1891 (
    .ADR0(DLX_IDinst_reg_out_B[23]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[23]),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_189)
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_253/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0095_inst_cy_253/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_253)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_253_2561 (
    .IA(DLX_IDinst_reg_out_B[23]),
    .IB(DLX_EXinst_Mcompar__n0095_inst_cy_252),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_189),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_253/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_253/CYINIT_2562  (
    .I(DLX_EXinst_Mcompar__n0095_inst_cy_251),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_253/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_254_2563 (
    .IA(DLX_IDinst_reg_out_B[24]),
    .IB(\DLX_IFinst_IR_curr<31>/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_190),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_254)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1901.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1901 (
    .ADR0(DLX_IDinst_reg_out_B[24]),
    .ADR1(DLX_IDinst_reg_out_A[24]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_190)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1911.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1911 (
    .ADR0(DLX_IDinst_reg_out_B[25]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[25]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_191)
  );
  X_BUF \DLX_IFinst_IR_curr<31>/COUTUSED  (
    .I(\DLX_IFinst_IR_curr<31>/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_255)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_255_2564 (
    .IA(DLX_IDinst_reg_out_B[25]),
    .IB(DLX_EXinst_Mcompar__n0095_inst_cy_254),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_191),
    .O(\DLX_IFinst_IR_curr<31>/CYMUXG )
  );
  X_BUF \DLX_IFinst_IR_curr<31>/CYINIT_2565  (
    .I(DLX_EXinst_Mcompar__n0095_inst_cy_253),
    .O(\DLX_IFinst_IR_curr<31>/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_256_2566 (
    .IA(DLX_IDinst_reg_out_B[26]),
    .IB(\DLX_EXinst_Mcompar__n0095_inst_cy_257/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_192),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_256)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1921.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1921 (
    .ADR0(DLX_IDinst_reg_out_B[26]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[26]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_192)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1931.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1931 (
    .ADR0(DLX_IDinst_reg_out_B[27]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[27]),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_193)
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_257/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0095_inst_cy_257/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_257)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_257_2567 (
    .IA(DLX_IDinst_reg_out_B[27]),
    .IB(DLX_EXinst_Mcompar__n0095_inst_cy_256),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_193),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_257/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_257/CYINIT_2568  (
    .I(DLX_EXinst_Mcompar__n0095_inst_cy_255),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_257/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_258_2569 (
    .IA(DLX_IDinst_reg_out_B[28]),
    .IB(\DLX_EXinst_Mcompar__n0095_inst_cy_259/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_194),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_258)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1941.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1941 (
    .ADR0(DLX_IDinst_reg_out_B[28]),
    .ADR1(DLX_IDinst_reg_out_A[28]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_194)
  );
  defparam DLX_EXinst_Mcompar__n0095_inst_lut2_1951.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0095_inst_lut2_1951 (
    .ADR0(DLX_IDinst_reg_out_B[29]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[29]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0095_inst_lut2_195)
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_259/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0095_inst_cy_259/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0095_inst_cy_259)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0095_inst_cy_259_2570 (
    .IA(DLX_IDinst_reg_out_B[29]),
    .IB(DLX_EXinst_Mcompar__n0095_inst_cy_258),
    .SEL(DLX_EXinst_Mcompar__n0095_inst_lut2_195),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_259/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0095_inst_cy_259/CYINIT_2571  (
    .I(DLX_EXinst_Mcompar__n0095_inst_cy_257),
    .O(\DLX_EXinst_Mcompar__n0095_inst_cy_259/CYINIT )
  );
  X_ZERO \DLX_IDinst_Madd__n0158_inst_lut2_230/LOGIC_ZERO_2572  (
    .O(\DLX_IDinst_Madd__n0158_inst_lut2_230/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Madd__n0158_inst_cy_297_2573 (
    .IA(DLX_IFinst_NPC[0]),
    .IB(\DLX_IDinst_Madd__n0158_inst_lut2_230/LOGIC_ZERO ),
    .SEL(\DLX_IDinst_Madd__n0158_inst_lut2_230/FROM ),
    .O(DLX_IDinst_Madd__n0158_inst_cy_297)
  );
  defparam DLX_IDinst_Madd__n0158_inst_lut2_2301.INIT = 16'h5A5A;
  X_LUT4 DLX_IDinst_Madd__n0158_inst_lut2_2301 (
    .ADR0(DLX_IFinst_NPC[0]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_jtarget[0]),
    .ADR3(VCC),
    .O(\DLX_IDinst_Madd__n0158_inst_lut2_230/FROM )
  );
  defparam DLX_IDinst_Madd__n0158_inst_lut2_2311.INIT = 16'h656A;
  X_LUT4 DLX_IDinst_Madd__n0158_inst_lut2_2311 (
    .ADR0(DLX_IFinst_NPC[1]),
    .ADR1(DLX_IFinst_IR_latched[1]),
    .ADR2(DLX_EXinst__n0144),
    .ADR3(DLX_IDinst_current_IR[1]),
    .O(DLX_IDinst_Madd__n0158_inst_lut2_231)
  );
  X_BUF \DLX_IDinst_Madd__n0158_inst_lut2_230/COUTUSED  (
    .I(\DLX_IDinst_Madd__n0158_inst_lut2_230/CYMUXG ),
    .O(DLX_IDinst_Madd__n0158_inst_cy_298)
  );
  X_BUF \DLX_IDinst_Madd__n0158_inst_lut2_230/XUSED  (
    .I(\DLX_IDinst_Madd__n0158_inst_lut2_230/FROM ),
    .O(DLX_IDinst_Madd__n0158_inst_lut2_230)
  );
  X_BUF \DLX_IDinst_Madd__n0158_inst_lut2_230/YUSED  (
    .I(\DLX_IDinst_Madd__n0158_inst_lut2_230/XORG ),
    .O(DLX_IDinst__n0158[1])
  );
  X_MUX2 DLX_IDinst_Madd__n0158_inst_cy_298_2574 (
    .IA(DLX_IFinst_NPC[1]),
    .IB(DLX_IDinst_Madd__n0158_inst_cy_297),
    .SEL(DLX_IDinst_Madd__n0158_inst_lut2_231),
    .O(\DLX_IDinst_Madd__n0158_inst_lut2_230/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Madd__n0158_inst_sum_135 (
    .I0(DLX_IDinst_Madd__n0158_inst_cy_297),
    .I1(DLX_IDinst_Madd__n0158_inst_lut2_231),
    .O(\DLX_IDinst_Madd__n0158_inst_lut2_230/XORG )
  );
  X_MUX2 DLX_IDinst_Madd__n0158_inst_cy_299_2575 (
    .IA(DLX_IFinst_NPC[2]),
    .IB(\DLX_IDinst_RegFile_2_30/CYINIT ),
    .SEL(DLX_IDinst_Madd__n0158_inst_lut2_232),
    .O(DLX_IDinst_Madd__n0158_inst_cy_299)
  );
  X_XOR2 DLX_IDinst_Madd__n0158_inst_sum_136 (
    .I0(\DLX_IDinst_RegFile_2_30/CYINIT ),
    .I1(DLX_IDinst_Madd__n0158_inst_lut2_232),
    .O(\DLX_IDinst_RegFile_2_30/XORF )
  );
  defparam DLX_IDinst_Madd__n0158_inst_lut2_2321.INIT = 16'h56A6;
  X_LUT4 DLX_IDinst_Madd__n0158_inst_lut2_2321 (
    .ADR0(DLX_IFinst_NPC[2]),
    .ADR1(DLX_IDinst_current_IR[2]),
    .ADR2(DLX_EXinst__n0144),
    .ADR3(DLX_IFinst_IR_latched[2]),
    .O(DLX_IDinst_Madd__n0158_inst_lut2_232)
  );
  defparam DLX_IDinst_Madd__n0158_inst_lut2_2331.INIT = 16'h5A66;
  X_LUT4 DLX_IDinst_Madd__n0158_inst_lut2_2331 (
    .ADR0(DLX_IFinst_NPC[3]),
    .ADR1(DLX_IDinst_current_IR[3]),
    .ADR2(DLX_IFinst_IR_latched[3]),
    .ADR3(DLX_EXinst__n0144),
    .O(DLX_IDinst_Madd__n0158_inst_lut2_233)
  );
  X_BUF \DLX_IDinst_RegFile_2_30/COUTUSED  (
    .I(\DLX_IDinst_RegFile_2_30/CYMUXG ),
    .O(DLX_IDinst_Madd__n0158_inst_cy_300)
  );
  X_BUF \DLX_IDinst_RegFile_2_30/XUSED  (
    .I(\DLX_IDinst_RegFile_2_30/XORF ),
    .O(DLX_IDinst__n0158[2])
  );
  X_BUF \DLX_IDinst_RegFile_2_30/YUSED  (
    .I(\DLX_IDinst_RegFile_2_30/XORG ),
    .O(DLX_IDinst__n0158[3])
  );
  X_MUX2 DLX_IDinst_Madd__n0158_inst_cy_300_2576 (
    .IA(DLX_IFinst_NPC[3]),
    .IB(DLX_IDinst_Madd__n0158_inst_cy_299),
    .SEL(DLX_IDinst_Madd__n0158_inst_lut2_233),
    .O(\DLX_IDinst_RegFile_2_30/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Madd__n0158_inst_sum_137 (
    .I0(DLX_IDinst_Madd__n0158_inst_cy_299),
    .I1(DLX_IDinst_Madd__n0158_inst_lut2_233),
    .O(\DLX_IDinst_RegFile_2_30/XORG )
  );
  X_BUF \DLX_IDinst_RegFile_2_30/CYINIT_2577  (
    .I(DLX_IDinst_Madd__n0158_inst_cy_298),
    .O(\DLX_IDinst_RegFile_2_30/CYINIT )
  );
  X_MUX2 DLX_IDinst_Madd__n0158_inst_cy_301_2578 (
    .IA(DLX_IFinst_NPC[4]),
    .IB(\DLX_IDinst__n0158<4>/CYINIT ),
    .SEL(DLX_IDinst_Madd__n0158_inst_lut2_234),
    .O(DLX_IDinst_Madd__n0158_inst_cy_301)
  );
  X_XOR2 DLX_IDinst_Madd__n0158_inst_sum_138 (
    .I0(\DLX_IDinst__n0158<4>/CYINIT ),
    .I1(DLX_IDinst_Madd__n0158_inst_lut2_234),
    .O(\DLX_IDinst__n0158<4>/XORF )
  );
  defparam DLX_IDinst_Madd__n0158_inst_lut2_2341.INIT = 16'h5A66;
  X_LUT4 DLX_IDinst_Madd__n0158_inst_lut2_2341 (
    .ADR0(DLX_IFinst_NPC[4]),
    .ADR1(DLX_IDinst_current_IR[4]),
    .ADR2(DLX_IFinst_IR_latched[4]),
    .ADR3(DLX_EXinst__n0144),
    .O(DLX_IDinst_Madd__n0158_inst_lut2_234)
  );
  defparam DLX_IDinst_Madd__n0158_inst_lut2_2351.INIT = 16'h5A66;
  X_LUT4 DLX_IDinst_Madd__n0158_inst_lut2_2351 (
    .ADR0(DLX_IFinst_NPC[5]),
    .ADR1(DLX_IDinst_current_IR[5]),
    .ADR2(DLX_IFinst_IR_latched[5]),
    .ADR3(DLX_EXinst__n0144),
    .O(DLX_IDinst_Madd__n0158_inst_lut2_235)
  );
  X_BUF \DLX_IDinst__n0158<4>/COUTUSED  (
    .I(\DLX_IDinst__n0158<4>/CYMUXG ),
    .O(DLX_IDinst_Madd__n0158_inst_cy_302)
  );
  X_BUF \DLX_IDinst__n0158<4>/XUSED  (
    .I(\DLX_IDinst__n0158<4>/XORF ),
    .O(DLX_IDinst__n0158[4])
  );
  X_BUF \DLX_IDinst__n0158<4>/YUSED  (
    .I(\DLX_IDinst__n0158<4>/XORG ),
    .O(DLX_IDinst__n0158[5])
  );
  X_MUX2 DLX_IDinst_Madd__n0158_inst_cy_302_2579 (
    .IA(DLX_IFinst_NPC[5]),
    .IB(DLX_IDinst_Madd__n0158_inst_cy_301),
    .SEL(DLX_IDinst_Madd__n0158_inst_lut2_235),
    .O(\DLX_IDinst__n0158<4>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Madd__n0158_inst_sum_139 (
    .I0(DLX_IDinst_Madd__n0158_inst_cy_301),
    .I1(DLX_IDinst_Madd__n0158_inst_lut2_235),
    .O(\DLX_IDinst__n0158<4>/XORG )
  );
  X_BUF \DLX_IDinst__n0158<4>/CYINIT_2580  (
    .I(DLX_IDinst_Madd__n0158_inst_cy_300),
    .O(\DLX_IDinst__n0158<4>/CYINIT )
  );
  X_MUX2 DLX_IDinst_Madd__n0158_inst_cy_303_2581 (
    .IA(DLX_IFinst_NPC[6]),
    .IB(\DLX_IDinst__n0158<6>/CYINIT ),
    .SEL(DLX_IDinst_Madd__n0158_inst_lut2_236),
    .O(DLX_IDinst_Madd__n0158_inst_cy_303)
  );
  X_XOR2 DLX_IDinst_Madd__n0158_inst_sum_140 (
    .I0(\DLX_IDinst__n0158<6>/CYINIT ),
    .I1(DLX_IDinst_Madd__n0158_inst_lut2_236),
    .O(\DLX_IDinst__n0158<6>/XORF )
  );
  defparam DLX_IDinst_Madd__n0158_inst_lut2_2361.INIT = 16'h665A;
  X_LUT4 DLX_IDinst_Madd__n0158_inst_lut2_2361 (
    .ADR0(DLX_IFinst_NPC[6]),
    .ADR1(DLX_IFinst_IR_latched[6]),
    .ADR2(DLX_IDinst_current_IR[6]),
    .ADR3(DLX_EXinst__n0144),
    .O(DLX_IDinst_Madd__n0158_inst_lut2_236)
  );
  defparam DLX_IDinst_Madd__n0158_inst_lut2_2371.INIT = 16'h596A;
  X_LUT4 DLX_IDinst_Madd__n0158_inst_lut2_2371 (
    .ADR0(DLX_IFinst_NPC[7]),
    .ADR1(DLX_EXinst__n0144),
    .ADR2(DLX_IFinst_IR_latched[7]),
    .ADR3(DLX_IDinst_current_IR[7]),
    .O(DLX_IDinst_Madd__n0158_inst_lut2_237)
  );
  X_BUF \DLX_IDinst__n0158<6>/COUTUSED  (
    .I(\DLX_IDinst__n0158<6>/CYMUXG ),
    .O(DLX_IDinst_Madd__n0158_inst_cy_304)
  );
  X_BUF \DLX_IDinst__n0158<6>/XUSED  (
    .I(\DLX_IDinst__n0158<6>/XORF ),
    .O(DLX_IDinst__n0158[6])
  );
  X_BUF \DLX_IDinst__n0158<6>/YUSED  (
    .I(\DLX_IDinst__n0158<6>/XORG ),
    .O(DLX_IDinst__n0158[7])
  );
  X_MUX2 DLX_IDinst_Madd__n0158_inst_cy_304_2582 (
    .IA(DLX_IFinst_NPC[7]),
    .IB(DLX_IDinst_Madd__n0158_inst_cy_303),
    .SEL(DLX_IDinst_Madd__n0158_inst_lut2_237),
    .O(\DLX_IDinst__n0158<6>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Madd__n0158_inst_sum_141 (
    .I0(DLX_IDinst_Madd__n0158_inst_cy_303),
    .I1(DLX_IDinst_Madd__n0158_inst_lut2_237),
    .O(\DLX_IDinst__n0158<6>/XORG )
  );
  X_BUF \DLX_IDinst__n0158<6>/CYINIT_2583  (
    .I(DLX_IDinst_Madd__n0158_inst_cy_302),
    .O(\DLX_IDinst__n0158<6>/CYINIT )
  );
  X_MUX2 DLX_IDinst_Madd__n0158_inst_cy_305_2584 (
    .IA(DLX_IFinst_NPC[8]),
    .IB(\DLX_IDinst__n0158<8>/CYINIT ),
    .SEL(DLX_IDinst_Madd__n0158_inst_lut2_238),
    .O(DLX_IDinst_Madd__n0158_inst_cy_305)
  );
  X_XOR2 DLX_IDinst_Madd__n0158_inst_sum_142 (
    .I0(\DLX_IDinst__n0158<8>/CYINIT ),
    .I1(DLX_IDinst_Madd__n0158_inst_lut2_238),
    .O(\DLX_IDinst__n0158<8>/XORF )
  );
  defparam DLX_IDinst_Madd__n0158_inst_lut2_2381.INIT = 16'h569A;
  X_LUT4 DLX_IDinst_Madd__n0158_inst_lut2_2381 (
    .ADR0(DLX_IFinst_NPC[8]),
    .ADR1(DLX_EXinst__n0144),
    .ADR2(DLX_IDinst_current_IR[8]),
    .ADR3(DLX_IFinst_IR_latched[8]),
    .O(DLX_IDinst_Madd__n0158_inst_lut2_238)
  );
  defparam DLX_IDinst_Madd__n0158_inst_lut2_2391.INIT = 16'h665A;
  X_LUT4 DLX_IDinst_Madd__n0158_inst_lut2_2391 (
    .ADR0(DLX_IFinst_NPC[9]),
    .ADR1(DLX_IFinst_IR_latched[9]),
    .ADR2(DLX_IDinst_current_IR[9]),
    .ADR3(DLX_EXinst__n0144),
    .O(DLX_IDinst_Madd__n0158_inst_lut2_239)
  );
  X_BUF \DLX_IDinst__n0158<8>/COUTUSED  (
    .I(\DLX_IDinst__n0158<8>/CYMUXG ),
    .O(DLX_IDinst_Madd__n0158_inst_cy_306)
  );
  X_BUF \DLX_IDinst__n0158<8>/XUSED  (
    .I(\DLX_IDinst__n0158<8>/XORF ),
    .O(DLX_IDinst__n0158[8])
  );
  X_BUF \DLX_IDinst__n0158<8>/YUSED  (
    .I(\DLX_IDinst__n0158<8>/XORG ),
    .O(DLX_IDinst__n0158[9])
  );
  X_MUX2 DLX_IDinst_Madd__n0158_inst_cy_306_2585 (
    .IA(DLX_IFinst_NPC[9]),
    .IB(DLX_IDinst_Madd__n0158_inst_cy_305),
    .SEL(DLX_IDinst_Madd__n0158_inst_lut2_239),
    .O(\DLX_IDinst__n0158<8>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Madd__n0158_inst_sum_143 (
    .I0(DLX_IDinst_Madd__n0158_inst_cy_305),
    .I1(DLX_IDinst_Madd__n0158_inst_lut2_239),
    .O(\DLX_IDinst__n0158<8>/XORG )
  );
  X_BUF \DLX_IDinst__n0158<8>/CYINIT_2586  (
    .I(DLX_IDinst_Madd__n0158_inst_cy_304),
    .O(\DLX_IDinst__n0158<8>/CYINIT )
  );
  X_MUX2 DLX_IDinst_Madd__n0158_inst_cy_307_2587 (
    .IA(DLX_IFinst_NPC[10]),
    .IB(\DLX_IFinst_IR_curr<24>/CYINIT ),
    .SEL(DLX_IDinst_Madd__n0158_inst_lut2_240),
    .O(DLX_IDinst_Madd__n0158_inst_cy_307)
  );
  X_XOR2 DLX_IDinst_Madd__n0158_inst_sum_144 (
    .I0(\DLX_IFinst_IR_curr<24>/CYINIT ),
    .I1(DLX_IDinst_Madd__n0158_inst_lut2_240),
    .O(\DLX_IFinst_IR_curr<24>/XORF )
  );
  defparam DLX_IDinst_Madd__n0158_inst_lut2_2401.INIT = 16'h665A;
  X_LUT4 DLX_IDinst_Madd__n0158_inst_lut2_2401 (
    .ADR0(DLX_IFinst_NPC[10]),
    .ADR1(DLX_IFinst_IR_latched[10]),
    .ADR2(DLX_IDinst_current_IR[10]),
    .ADR3(DLX_EXinst__n0144),
    .O(DLX_IDinst_Madd__n0158_inst_lut2_240)
  );
  defparam DLX_IDinst_Madd__n0158_inst_lut2_2411.INIT = 16'h5A66;
  X_LUT4 DLX_IDinst_Madd__n0158_inst_lut2_2411 (
    .ADR0(DLX_IFinst_NPC[11]),
    .ADR1(DLX_IDinst_current_IR[11]),
    .ADR2(DLX_IFinst_IR_latched[11]),
    .ADR3(DLX_EXinst__n0144),
    .O(DLX_IDinst_Madd__n0158_inst_lut2_241)
  );
  X_BUF \DLX_IFinst_IR_curr<24>/COUTUSED  (
    .I(\DLX_IFinst_IR_curr<24>/CYMUXG ),
    .O(DLX_IDinst_Madd__n0158_inst_cy_308)
  );
  X_BUF \DLX_IFinst_IR_curr<24>/XUSED  (
    .I(\DLX_IFinst_IR_curr<24>/XORF ),
    .O(DLX_IDinst__n0158[10])
  );
  X_BUF \DLX_IFinst_IR_curr<24>/YUSED  (
    .I(\DLX_IFinst_IR_curr<24>/XORG ),
    .O(DLX_IDinst__n0158[11])
  );
  X_MUX2 DLX_IDinst_Madd__n0158_inst_cy_308_2588 (
    .IA(DLX_IFinst_NPC[11]),
    .IB(DLX_IDinst_Madd__n0158_inst_cy_307),
    .SEL(DLX_IDinst_Madd__n0158_inst_lut2_241),
    .O(\DLX_IFinst_IR_curr<24>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Madd__n0158_inst_sum_145 (
    .I0(DLX_IDinst_Madd__n0158_inst_cy_307),
    .I1(DLX_IDinst_Madd__n0158_inst_lut2_241),
    .O(\DLX_IFinst_IR_curr<24>/XORG )
  );
  X_BUF \DLX_IFinst_IR_curr<24>/CYINIT_2589  (
    .I(DLX_IDinst_Madd__n0158_inst_cy_306),
    .O(\DLX_IFinst_IR_curr<24>/CYINIT )
  );
  defparam DLX_IDinst_RegFile_29_26_2590.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_29_26_2590 (
    .I(DLX_IDinst_WB_data_eff[26]),
    .CE(DLX_IDinst__n0608),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_29_26)
  );
  X_MUX2 DLX_IDinst_Madd__n0158_inst_cy_309_2591 (
    .IA(DLX_IFinst_NPC[12]),
    .IB(\DLX_IDinst__n0158<12>/CYINIT ),
    .SEL(DLX_IDinst_Madd__n0158_inst_lut2_242),
    .O(DLX_IDinst_Madd__n0158_inst_cy_309)
  );
  X_XOR2 DLX_IDinst_Madd__n0158_inst_sum_146 (
    .I0(\DLX_IDinst__n0158<12>/CYINIT ),
    .I1(DLX_IDinst_Madd__n0158_inst_lut2_242),
    .O(\DLX_IDinst__n0158<12>/XORF )
  );
  defparam DLX_IDinst_Madd__n0158_inst_lut2_2421.INIT = 16'h5A66;
  X_LUT4 DLX_IDinst_Madd__n0158_inst_lut2_2421 (
    .ADR0(DLX_IFinst_NPC[12]),
    .ADR1(DLX_IDinst_current_IR[12]),
    .ADR2(DLX_IFinst_IR_latched[12]),
    .ADR3(DLX_EXinst__n0144),
    .O(DLX_IDinst_Madd__n0158_inst_lut2_242)
  );
  defparam DLX_IDinst_Madd__n0158_inst_lut2_2431.INIT = 16'h656A;
  X_LUT4 DLX_IDinst_Madd__n0158_inst_lut2_2431 (
    .ADR0(DLX_IFinst_NPC[13]),
    .ADR1(DLX_IFinst_IR_latched[13]),
    .ADR2(DLX_EXinst__n0144),
    .ADR3(DLX_IDinst_current_IR[13]),
    .O(DLX_IDinst_Madd__n0158_inst_lut2_243)
  );
  X_BUF \DLX_IDinst__n0158<12>/COUTUSED  (
    .I(\DLX_IDinst__n0158<12>/CYMUXG ),
    .O(DLX_IDinst_Madd__n0158_inst_cy_310)
  );
  X_BUF \DLX_IDinst__n0158<12>/XUSED  (
    .I(\DLX_IDinst__n0158<12>/XORF ),
    .O(DLX_IDinst__n0158[12])
  );
  X_BUF \DLX_IDinst__n0158<12>/YUSED  (
    .I(\DLX_IDinst__n0158<12>/XORG ),
    .O(DLX_IDinst__n0158[13])
  );
  X_MUX2 DLX_IDinst_Madd__n0158_inst_cy_310_2592 (
    .IA(DLX_IFinst_NPC[13]),
    .IB(DLX_IDinst_Madd__n0158_inst_cy_309),
    .SEL(DLX_IDinst_Madd__n0158_inst_lut2_243),
    .O(\DLX_IDinst__n0158<12>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Madd__n0158_inst_sum_147 (
    .I0(DLX_IDinst_Madd__n0158_inst_cy_309),
    .I1(DLX_IDinst_Madd__n0158_inst_lut2_243),
    .O(\DLX_IDinst__n0158<12>/XORG )
  );
  X_BUF \DLX_IDinst__n0158<12>/CYINIT_2593  (
    .I(DLX_IDinst_Madd__n0158_inst_cy_308),
    .O(\DLX_IDinst__n0158<12>/CYINIT )
  );
  X_MUX2 DLX_IDinst_Madd__n0158_inst_cy_311_2594 (
    .IA(DLX_IFinst_NPC[14]),
    .IB(\DLX_IDinst__n0158<14>/CYINIT ),
    .SEL(DLX_IDinst_Madd__n0158_inst_lut2_244),
    .O(DLX_IDinst_Madd__n0158_inst_cy_311)
  );
  X_XOR2 DLX_IDinst_Madd__n0158_inst_sum_148 (
    .I0(\DLX_IDinst__n0158<14>/CYINIT ),
    .I1(DLX_IDinst_Madd__n0158_inst_lut2_244),
    .O(\DLX_IDinst__n0158<14>/XORF )
  );
  defparam DLX_IDinst_Madd__n0158_inst_lut2_2441.INIT = 16'h569A;
  X_LUT4 DLX_IDinst_Madd__n0158_inst_lut2_2441 (
    .ADR0(DLX_IFinst_NPC[14]),
    .ADR1(DLX_EXinst__n0144),
    .ADR2(DLX_IDinst_current_IR[14]),
    .ADR3(DLX_IFinst_IR_latched[14]),
    .O(DLX_IDinst_Madd__n0158_inst_lut2_244)
  );
  defparam DLX_IDinst_Madd__n0158_inst_lut2_2451.INIT = 16'h656A;
  X_LUT4 DLX_IDinst_Madd__n0158_inst_lut2_2451 (
    .ADR0(DLX_IFinst_NPC[15]),
    .ADR1(DLX_IFinst_IR_latched[15]),
    .ADR2(DLX_EXinst__n0144),
    .ADR3(DLX_IDinst_current_IR[15]),
    .O(DLX_IDinst_Madd__n0158_inst_lut2_245)
  );
  X_BUF \DLX_IDinst__n0158<14>/COUTUSED  (
    .I(\DLX_IDinst__n0158<14>/CYMUXG ),
    .O(DLX_IDinst_Madd__n0158_inst_cy_312)
  );
  X_BUF \DLX_IDinst__n0158<14>/XUSED  (
    .I(\DLX_IDinst__n0158<14>/XORF ),
    .O(DLX_IDinst__n0158[14])
  );
  X_BUF \DLX_IDinst__n0158<14>/YUSED  (
    .I(\DLX_IDinst__n0158<14>/XORG ),
    .O(DLX_IDinst__n0158[15])
  );
  X_MUX2 DLX_IDinst_Madd__n0158_inst_cy_312_2595 (
    .IA(DLX_IFinst_NPC[15]),
    .IB(DLX_IDinst_Madd__n0158_inst_cy_311),
    .SEL(DLX_IDinst_Madd__n0158_inst_lut2_245),
    .O(\DLX_IDinst__n0158<14>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Madd__n0158_inst_sum_149 (
    .I0(DLX_IDinst_Madd__n0158_inst_cy_311),
    .I1(DLX_IDinst_Madd__n0158_inst_lut2_245),
    .O(\DLX_IDinst__n0158<14>/XORG )
  );
  X_BUF \DLX_IDinst__n0158<14>/CYINIT_2596  (
    .I(DLX_IDinst_Madd__n0158_inst_cy_310),
    .O(\DLX_IDinst__n0158<14>/CYINIT )
  );
  X_MUX2 DLX_IDinst_Madd__n0158_inst_cy_313_2597 (
    .IA(DLX_IFinst_NPC[16]),
    .IB(\DLX_IDinst__n0158<16>/CYINIT ),
    .SEL(DLX_IDinst_Madd__n0158_inst_lut2_246),
    .O(DLX_IDinst_Madd__n0158_inst_cy_313)
  );
  X_XOR2 DLX_IDinst_Madd__n0158_inst_sum_150 (
    .I0(\DLX_IDinst__n0158<16>/CYINIT ),
    .I1(DLX_IDinst_Madd__n0158_inst_lut2_246),
    .O(\DLX_IDinst__n0158<16>/XORF )
  );
  defparam DLX_IDinst_Madd__n0158_inst_lut2_2461.INIT = 16'h569A;
  X_LUT4 DLX_IDinst_Madd__n0158_inst_lut2_2461 (
    .ADR0(DLX_IFinst_NPC[16]),
    .ADR1(DLX_IDinst__n0635),
    .ADR2(DLX_IDinst_jtarget[15]),
    .ADR3(DLX_IDinst_jtarget[16]),
    .O(DLX_IDinst_Madd__n0158_inst_lut2_246)
  );
  defparam DLX_IDinst_Madd__n0158_inst_lut2_2471.INIT = 16'h596A;
  X_LUT4 DLX_IDinst_Madd__n0158_inst_lut2_2471 (
    .ADR0(DLX_IFinst_NPC[17]),
    .ADR1(DLX_IDinst__n0635),
    .ADR2(DLX_IDinst_jtarget[17]),
    .ADR3(DLX_IDinst_jtarget[15]),
    .O(DLX_IDinst_Madd__n0158_inst_lut2_247)
  );
  X_BUF \DLX_IDinst__n0158<16>/COUTUSED  (
    .I(\DLX_IDinst__n0158<16>/CYMUXG ),
    .O(DLX_IDinst_Madd__n0158_inst_cy_314)
  );
  X_BUF \DLX_IDinst__n0158<16>/XUSED  (
    .I(\DLX_IDinst__n0158<16>/XORF ),
    .O(DLX_IDinst__n0158[16])
  );
  X_BUF \DLX_IDinst__n0158<16>/YUSED  (
    .I(\DLX_IDinst__n0158<16>/XORG ),
    .O(DLX_IDinst__n0158[17])
  );
  X_MUX2 DLX_IDinst_Madd__n0158_inst_cy_314_2598 (
    .IA(DLX_IFinst_NPC[17]),
    .IB(DLX_IDinst_Madd__n0158_inst_cy_313),
    .SEL(DLX_IDinst_Madd__n0158_inst_lut2_247),
    .O(\DLX_IDinst__n0158<16>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Madd__n0158_inst_sum_151 (
    .I0(DLX_IDinst_Madd__n0158_inst_cy_313),
    .I1(DLX_IDinst_Madd__n0158_inst_lut2_247),
    .O(\DLX_IDinst__n0158<16>/XORG )
  );
  X_BUF \DLX_IDinst__n0158<16>/CYINIT_2599  (
    .I(DLX_IDinst_Madd__n0158_inst_cy_312),
    .O(\DLX_IDinst__n0158<16>/CYINIT )
  );
  X_MUX2 DLX_IDinst_Madd__n0158_inst_cy_315_2600 (
    .IA(DLX_IFinst_NPC[18]),
    .IB(\DLX_IDinst_RegFile_0_6/CYINIT ),
    .SEL(DLX_IDinst_Madd__n0158_inst_lut2_248),
    .O(DLX_IDinst_Madd__n0158_inst_cy_315)
  );
  X_XOR2 DLX_IDinst_Madd__n0158_inst_sum_152 (
    .I0(\DLX_IDinst_RegFile_0_6/CYINIT ),
    .I1(DLX_IDinst_Madd__n0158_inst_lut2_248),
    .O(\DLX_IDinst_RegFile_0_6/XORF )
  );
  defparam DLX_IDinst_Madd__n0158_inst_lut2_2481.INIT = 16'h656A;
  X_LUT4 DLX_IDinst_Madd__n0158_inst_lut2_2481 (
    .ADR0(DLX_IFinst_NPC[18]),
    .ADR1(DLX_IDinst_jtarget[18]),
    .ADR2(DLX_IDinst__n0635),
    .ADR3(DLX_IDinst_jtarget[15]),
    .O(DLX_IDinst_Madd__n0158_inst_lut2_248)
  );
  defparam DLX_IDinst_Madd__n0158_inst_lut2_2491.INIT = 16'h656A;
  X_LUT4 DLX_IDinst_Madd__n0158_inst_lut2_2491 (
    .ADR0(DLX_IFinst_NPC[19]),
    .ADR1(DLX_IDinst_jtarget[19]),
    .ADR2(DLX_IDinst__n0635),
    .ADR3(DLX_IDinst_jtarget[15]),
    .O(DLX_IDinst_Madd__n0158_inst_lut2_249)
  );
  X_BUF \DLX_IDinst_RegFile_0_6/COUTUSED  (
    .I(\DLX_IDinst_RegFile_0_6/CYMUXG ),
    .O(DLX_IDinst_Madd__n0158_inst_cy_316)
  );
  X_BUF \DLX_IDinst_RegFile_0_6/XUSED  (
    .I(\DLX_IDinst_RegFile_0_6/XORF ),
    .O(DLX_IDinst__n0158[18])
  );
  X_BUF \DLX_IDinst_RegFile_0_6/YUSED  (
    .I(\DLX_IDinst_RegFile_0_6/XORG ),
    .O(DLX_IDinst__n0158[19])
  );
  X_MUX2 DLX_IDinst_Madd__n0158_inst_cy_316_2601 (
    .IA(DLX_IFinst_NPC[19]),
    .IB(DLX_IDinst_Madd__n0158_inst_cy_315),
    .SEL(DLX_IDinst_Madd__n0158_inst_lut2_249),
    .O(\DLX_IDinst_RegFile_0_6/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Madd__n0158_inst_sum_153 (
    .I0(DLX_IDinst_Madd__n0158_inst_cy_315),
    .I1(DLX_IDinst_Madd__n0158_inst_lut2_249),
    .O(\DLX_IDinst_RegFile_0_6/XORG )
  );
  X_BUF \DLX_IDinst_RegFile_0_6/CYINIT_2602  (
    .I(DLX_IDinst_Madd__n0158_inst_cy_314),
    .O(\DLX_IDinst_RegFile_0_6/CYINIT )
  );
  X_MUX2 DLX_IDinst_Madd__n0158_inst_cy_317_2603 (
    .IA(DLX_IFinst_NPC[20]),
    .IB(\DLX_IDinst__n0158<20>/CYINIT ),
    .SEL(DLX_IDinst_Madd__n0158_inst_lut2_250),
    .O(DLX_IDinst_Madd__n0158_inst_cy_317)
  );
  X_XOR2 DLX_IDinst_Madd__n0158_inst_sum_154 (
    .I0(\DLX_IDinst__n0158<20>/CYINIT ),
    .I1(DLX_IDinst_Madd__n0158_inst_lut2_250),
    .O(\DLX_IDinst__n0158<20>/XORF )
  );
  defparam DLX_IDinst_Madd__n0158_inst_lut2_2501.INIT = 16'h596A;
  X_LUT4 DLX_IDinst_Madd__n0158_inst_lut2_2501 (
    .ADR0(DLX_IFinst_NPC[20]),
    .ADR1(DLX_IDinst__n0635),
    .ADR2(DLX_IDinst_jtarget[20]),
    .ADR3(DLX_IDinst_jtarget[15]),
    .O(DLX_IDinst_Madd__n0158_inst_lut2_250)
  );
  defparam DLX_IDinst_Madd__n0158_inst_lut2_2511.INIT = 16'h569A;
  X_LUT4 DLX_IDinst_Madd__n0158_inst_lut2_2511 (
    .ADR0(DLX_IFinst_NPC[21]),
    .ADR1(DLX_IDinst__n0635),
    .ADR2(DLX_IDinst_jtarget[15]),
    .ADR3(DLX_IDinst_jtarget[21]),
    .O(DLX_IDinst_Madd__n0158_inst_lut2_251)
  );
  X_BUF \DLX_IDinst__n0158<20>/COUTUSED  (
    .I(\DLX_IDinst__n0158<20>/CYMUXG ),
    .O(DLX_IDinst_Madd__n0158_inst_cy_318)
  );
  X_BUF \DLX_IDinst__n0158<20>/XUSED  (
    .I(\DLX_IDinst__n0158<20>/XORF ),
    .O(DLX_IDinst__n0158[20])
  );
  X_BUF \DLX_IDinst__n0158<20>/YUSED  (
    .I(\DLX_IDinst__n0158<20>/XORG ),
    .O(DLX_IDinst__n0158[21])
  );
  X_MUX2 DLX_IDinst_Madd__n0158_inst_cy_318_2604 (
    .IA(DLX_IFinst_NPC[21]),
    .IB(DLX_IDinst_Madd__n0158_inst_cy_317),
    .SEL(DLX_IDinst_Madd__n0158_inst_lut2_251),
    .O(\DLX_IDinst__n0158<20>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Madd__n0158_inst_sum_155 (
    .I0(DLX_IDinst_Madd__n0158_inst_cy_317),
    .I1(DLX_IDinst_Madd__n0158_inst_lut2_251),
    .O(\DLX_IDinst__n0158<20>/XORG )
  );
  X_BUF \DLX_IDinst__n0158<20>/CYINIT_2605  (
    .I(DLX_IDinst_Madd__n0158_inst_cy_316),
    .O(\DLX_IDinst__n0158<20>/CYINIT )
  );
  X_MUX2 DLX_IDinst_Madd__n0158_inst_cy_319_2606 (
    .IA(DLX_IFinst_NPC[22]),
    .IB(\DLX_IDinst__n0158<22>/CYINIT ),
    .SEL(DLX_IDinst_Madd__n0158_inst_lut2_252),
    .O(DLX_IDinst_Madd__n0158_inst_cy_319)
  );
  X_XOR2 DLX_IDinst_Madd__n0158_inst_sum_156 (
    .I0(\DLX_IDinst__n0158<22>/CYINIT ),
    .I1(DLX_IDinst_Madd__n0158_inst_lut2_252),
    .O(\DLX_IDinst__n0158<22>/XORF )
  );
  defparam DLX_IDinst_Madd__n0158_inst_lut2_2521.INIT = 16'h569A;
  X_LUT4 DLX_IDinst_Madd__n0158_inst_lut2_2521 (
    .ADR0(DLX_IFinst_NPC[22]),
    .ADR1(DLX_IDinst__n0635),
    .ADR2(DLX_IDinst_jtarget[15]),
    .ADR3(DLX_IDinst_jtarget[22]),
    .O(DLX_IDinst_Madd__n0158_inst_lut2_252)
  );
  defparam DLX_IDinst_Madd__n0158_inst_lut2_2531.INIT = 16'h596A;
  X_LUT4 DLX_IDinst_Madd__n0158_inst_lut2_2531 (
    .ADR0(DLX_IFinst_NPC[23]),
    .ADR1(DLX_IDinst__n0635),
    .ADR2(DLX_IDinst_jtarget[23]),
    .ADR3(DLX_IDinst_jtarget[15]),
    .O(DLX_IDinst_Madd__n0158_inst_lut2_253)
  );
  X_BUF \DLX_IDinst__n0158<22>/COUTUSED  (
    .I(\DLX_IDinst__n0158<22>/CYMUXG ),
    .O(DLX_IDinst_Madd__n0158_inst_cy_320)
  );
  X_BUF \DLX_IDinst__n0158<22>/XUSED  (
    .I(\DLX_IDinst__n0158<22>/XORF ),
    .O(DLX_IDinst__n0158[22])
  );
  X_BUF \DLX_IDinst__n0158<22>/YUSED  (
    .I(\DLX_IDinst__n0158<22>/XORG ),
    .O(DLX_IDinst__n0158[23])
  );
  X_MUX2 DLX_IDinst_Madd__n0158_inst_cy_320_2607 (
    .IA(DLX_IFinst_NPC[23]),
    .IB(DLX_IDinst_Madd__n0158_inst_cy_319),
    .SEL(DLX_IDinst_Madd__n0158_inst_lut2_253),
    .O(\DLX_IDinst__n0158<22>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Madd__n0158_inst_sum_157 (
    .I0(DLX_IDinst_Madd__n0158_inst_cy_319),
    .I1(DLX_IDinst_Madd__n0158_inst_lut2_253),
    .O(\DLX_IDinst__n0158<22>/XORG )
  );
  X_BUF \DLX_IDinst__n0158<22>/CYINIT_2608  (
    .I(DLX_IDinst_Madd__n0158_inst_cy_318),
    .O(\DLX_IDinst__n0158<22>/CYINIT )
  );
  X_MUX2 DLX_IDinst_Madd__n0158_inst_cy_321_2609 (
    .IA(DLX_IFinst_NPC[24]),
    .IB(\DLX_IDinst__n0158<24>/CYINIT ),
    .SEL(DLX_IDinst_Madd__n0158_inst_lut2_254),
    .O(DLX_IDinst_Madd__n0158_inst_cy_321)
  );
  X_XOR2 DLX_IDinst_Madd__n0158_inst_sum_158 (
    .I0(\DLX_IDinst__n0158<24>/CYINIT ),
    .I1(DLX_IDinst_Madd__n0158_inst_lut2_254),
    .O(\DLX_IDinst__n0158<24>/XORF )
  );
  defparam DLX_IDinst_Madd__n0158_inst_lut2_2541.INIT = 16'h596A;
  X_LUT4 DLX_IDinst_Madd__n0158_inst_lut2_2541 (
    .ADR0(DLX_IFinst_NPC[24]),
    .ADR1(DLX_IDinst__n0635),
    .ADR2(DLX_IDinst_jtarget[24]),
    .ADR3(DLX_IDinst_jtarget[15]),
    .O(DLX_IDinst_Madd__n0158_inst_lut2_254)
  );
  defparam DLX_IDinst_Madd__n0158_inst_lut2_2551.INIT = 16'h656A;
  X_LUT4 DLX_IDinst_Madd__n0158_inst_lut2_2551 (
    .ADR0(DLX_IFinst_NPC[25]),
    .ADR1(DLX_IDinst_jtarget[25]),
    .ADR2(DLX_IDinst__n0635),
    .ADR3(DLX_IDinst_jtarget[15]),
    .O(DLX_IDinst_Madd__n0158_inst_lut2_255)
  );
  X_BUF \DLX_IDinst__n0158<24>/COUTUSED  (
    .I(\DLX_IDinst__n0158<24>/CYMUXG ),
    .O(DLX_IDinst_Madd__n0158_inst_cy_322)
  );
  X_BUF \DLX_IDinst__n0158<24>/XUSED  (
    .I(\DLX_IDinst__n0158<24>/XORF ),
    .O(DLX_IDinst__n0158[24])
  );
  X_BUF \DLX_IDinst__n0158<24>/YUSED  (
    .I(\DLX_IDinst__n0158<24>/XORG ),
    .O(DLX_IDinst__n0158[25])
  );
  X_MUX2 DLX_IDinst_Madd__n0158_inst_cy_322_2610 (
    .IA(DLX_IFinst_NPC[25]),
    .IB(DLX_IDinst_Madd__n0158_inst_cy_321),
    .SEL(DLX_IDinst_Madd__n0158_inst_lut2_255),
    .O(\DLX_IDinst__n0158<24>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Madd__n0158_inst_sum_159 (
    .I0(DLX_IDinst_Madd__n0158_inst_cy_321),
    .I1(DLX_IDinst_Madd__n0158_inst_lut2_255),
    .O(\DLX_IDinst__n0158<24>/XORG )
  );
  X_BUF \DLX_IDinst__n0158<24>/CYINIT_2611  (
    .I(DLX_IDinst_Madd__n0158_inst_cy_320),
    .O(\DLX_IDinst__n0158<24>/CYINIT )
  );
  X_MUX2 DLX_IDinst_Madd__n0158_inst_cy_323_2612 (
    .IA(DLX_IFinst_NPC[26]),
    .IB(\DLX_IFinst_IR_curr<16>/CYINIT ),
    .SEL(DLX_IDinst_Madd__n0158_inst_lut2_256),
    .O(DLX_IDinst_Madd__n0158_inst_cy_323)
  );
  X_XOR2 DLX_IDinst_Madd__n0158_inst_sum_160 (
    .I0(\DLX_IFinst_IR_curr<16>/CYINIT ),
    .I1(DLX_IDinst_Madd__n0158_inst_lut2_256),
    .O(\DLX_IFinst_IR_curr<16>/XORF )
  );
  defparam DLX_IDinst_Madd__n0158_inst_lut2_2561.INIT = 16'h656A;
  X_LUT4 DLX_IDinst_Madd__n0158_inst_lut2_2561 (
    .ADR0(DLX_IFinst_NPC[26]),
    .ADR1(DLX_IDinst_jtarget[25]),
    .ADR2(DLX_IDinst__n0635),
    .ADR3(DLX_IDinst_jtarget[15]),
    .O(DLX_IDinst_Madd__n0158_inst_lut2_256)
  );
  defparam DLX_IDinst_Madd__n0158_inst_lut2_2571.INIT = 16'h656A;
  X_LUT4 DLX_IDinst_Madd__n0158_inst_lut2_2571 (
    .ADR0(DLX_IFinst_NPC[27]),
    .ADR1(DLX_IDinst_jtarget[25]),
    .ADR2(DLX_IDinst__n0635),
    .ADR3(DLX_IDinst_jtarget[15]),
    .O(DLX_IDinst_Madd__n0158_inst_lut2_257)
  );
  X_BUF \DLX_IFinst_IR_curr<16>/COUTUSED  (
    .I(\DLX_IFinst_IR_curr<16>/CYMUXG ),
    .O(DLX_IDinst_Madd__n0158_inst_cy_324)
  );
  X_BUF \DLX_IFinst_IR_curr<16>/XUSED  (
    .I(\DLX_IFinst_IR_curr<16>/XORF ),
    .O(DLX_IDinst__n0158[26])
  );
  X_BUF \DLX_IFinst_IR_curr<16>/YUSED  (
    .I(\DLX_IFinst_IR_curr<16>/XORG ),
    .O(DLX_IDinst__n0158[27])
  );
  X_MUX2 DLX_IDinst_Madd__n0158_inst_cy_324_2613 (
    .IA(DLX_IFinst_NPC[27]),
    .IB(DLX_IDinst_Madd__n0158_inst_cy_323),
    .SEL(DLX_IDinst_Madd__n0158_inst_lut2_257),
    .O(\DLX_IFinst_IR_curr<16>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Madd__n0158_inst_sum_161 (
    .I0(DLX_IDinst_Madd__n0158_inst_cy_323),
    .I1(DLX_IDinst_Madd__n0158_inst_lut2_257),
    .O(\DLX_IFinst_IR_curr<16>/XORG )
  );
  X_BUF \DLX_IFinst_IR_curr<16>/CYINIT_2614  (
    .I(DLX_IDinst_Madd__n0158_inst_cy_322),
    .O(\DLX_IFinst_IR_curr<16>/CYINIT )
  );
  X_MUX2 DLX_IDinst_Madd__n0158_inst_cy_325_2615 (
    .IA(DLX_IFinst_NPC[28]),
    .IB(\DLX_IDinst__n0158<28>/CYINIT ),
    .SEL(DLX_IDinst_Madd__n0158_inst_lut2_258),
    .O(DLX_IDinst_Madd__n0158_inst_cy_325)
  );
  X_XOR2 DLX_IDinst_Madd__n0158_inst_sum_162 (
    .I0(\DLX_IDinst__n0158<28>/CYINIT ),
    .I1(DLX_IDinst_Madd__n0158_inst_lut2_258),
    .O(\DLX_IDinst__n0158<28>/XORF )
  );
  defparam DLX_IDinst_Madd__n0158_inst_lut2_2581.INIT = 16'h596A;
  X_LUT4 DLX_IDinst_Madd__n0158_inst_lut2_2581 (
    .ADR0(DLX_IFinst_NPC[28]),
    .ADR1(DLX_IDinst__n0635),
    .ADR2(DLX_IDinst_jtarget[25]),
    .ADR3(DLX_IDinst_jtarget[15]),
    .O(DLX_IDinst_Madd__n0158_inst_lut2_258)
  );
  defparam DLX_IDinst_Madd__n0158_inst_lut2_2591.INIT = 16'h596A;
  X_LUT4 DLX_IDinst_Madd__n0158_inst_lut2_2591 (
    .ADR0(DLX_IFinst_NPC[29]),
    .ADR1(DLX_IDinst__n0635),
    .ADR2(DLX_IDinst_jtarget[25]),
    .ADR3(DLX_IDinst_jtarget[15]),
    .O(DLX_IDinst_Madd__n0158_inst_lut2_259)
  );
  X_BUF \DLX_IDinst__n0158<28>/COUTUSED  (
    .I(\DLX_IDinst__n0158<28>/CYMUXG ),
    .O(DLX_IDinst_Madd__n0158_inst_cy_326)
  );
  X_BUF \DLX_IDinst__n0158<28>/XUSED  (
    .I(\DLX_IDinst__n0158<28>/XORF ),
    .O(DLX_IDinst__n0158[28])
  );
  X_BUF \DLX_IDinst__n0158<28>/YUSED  (
    .I(\DLX_IDinst__n0158<28>/XORG ),
    .O(DLX_IDinst__n0158[29])
  );
  X_MUX2 DLX_IDinst_Madd__n0158_inst_cy_326_2616 (
    .IA(DLX_IFinst_NPC[29]),
    .IB(DLX_IDinst_Madd__n0158_inst_cy_325),
    .SEL(DLX_IDinst_Madd__n0158_inst_lut2_259),
    .O(\DLX_IDinst__n0158<28>/CYMUXG )
  );
  X_XOR2 DLX_IDinst_Madd__n0158_inst_sum_163 (
    .I0(DLX_IDinst_Madd__n0158_inst_cy_325),
    .I1(DLX_IDinst_Madd__n0158_inst_lut2_259),
    .O(\DLX_IDinst__n0158<28>/XORG )
  );
  X_BUF \DLX_IDinst__n0158<28>/CYINIT_2617  (
    .I(DLX_IDinst_Madd__n0158_inst_cy_324),
    .O(\DLX_IDinst__n0158<28>/CYINIT )
  );
  X_MUX2 DLX_IDinst_Madd__n0158_inst_cy_327_2618 (
    .IA(DLX_IFinst_NPC[30]),
    .IB(\DLX_IDinst__n0158<30>/CYINIT ),
    .SEL(DLX_IDinst_Madd__n0158_inst_lut2_260),
    .O(DLX_IDinst_Madd__n0158_inst_cy_327)
  );
  X_XOR2 DLX_IDinst_Madd__n0158_inst_sum_164 (
    .I0(\DLX_IDinst__n0158<30>/CYINIT ),
    .I1(DLX_IDinst_Madd__n0158_inst_lut2_260),
    .O(\DLX_IDinst__n0158<30>/XORF )
  );
  defparam DLX_IDinst_Madd__n0158_inst_lut2_2601.INIT = 16'h656A;
  X_LUT4 DLX_IDinst_Madd__n0158_inst_lut2_2601 (
    .ADR0(DLX_IFinst_NPC[30]),
    .ADR1(DLX_IDinst_jtarget[25]),
    .ADR2(DLX_IDinst__n0635),
    .ADR3(DLX_IDinst_jtarget[15]),
    .O(DLX_IDinst_Madd__n0158_inst_lut2_260)
  );
  defparam DLX_IDinst_Madd__n0158_inst_lut2_2611.INIT = 16'h596A;
  X_LUT4 DLX_IDinst_Madd__n0158_inst_lut2_2611 (
    .ADR0(DLX_IFinst_NPC[31]),
    .ADR1(DLX_IDinst__n0635),
    .ADR2(DLX_IDinst_jtarget[25]),
    .ADR3(DLX_IDinst_jtarget[15]),
    .O(DLX_IDinst_Madd__n0158_inst_lut2_261)
  );
  X_BUF \DLX_IDinst__n0158<30>/XUSED  (
    .I(\DLX_IDinst__n0158<30>/XORF ),
    .O(DLX_IDinst__n0158[30])
  );
  X_BUF \DLX_IDinst__n0158<30>/YUSED  (
    .I(\DLX_IDinst__n0158<30>/XORG ),
    .O(DLX_IDinst__n0158[31])
  );
  X_XOR2 DLX_IDinst_Madd__n0158_inst_sum_165 (
    .I0(DLX_IDinst_Madd__n0158_inst_cy_327),
    .I1(DLX_IDinst_Madd__n0158_inst_lut2_261),
    .O(\DLX_IDinst__n0158<30>/XORG )
  );
  X_BUF \DLX_IDinst__n0158<30>/CYINIT_2619  (
    .I(DLX_IDinst_Madd__n0158_inst_cy_326),
    .O(\DLX_IDinst__n0158<30>/CYINIT )
  );
  X_ONE \DLX_IDinst_Mcompar__n0102_inst_cy_263/LOGIC_ONE_2620  (
    .O(\DLX_IDinst_Mcompar__n0102_inst_cy_263/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mcompar__n0102_inst_cy_263/LOGIC_ZERO_2621  (
    .O(\DLX_IDinst_Mcompar__n0102_inst_cy_263/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mcompar__n0102_inst_cy_262_2622 (
    .IA(\DLX_IDinst_Mcompar__n0102_inst_cy_263/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mcompar__n0102_inst_cy_263/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mcompar__n0102_inst_lut4_40),
    .O(DLX_IDinst_Mcompar__n0102_inst_cy_262)
  );
  defparam DLX_IDinst_Mcompar__n0102_inst_lut4_401.INIT = 16'h8241;
  X_LUT4 DLX_IDinst_Mcompar__n0102_inst_lut4_401 (
    .ADR0(DLX_reg_dst_of_EX[0]),
    .ADR1(DLX_reg_dst_of_EX[1]),
    .ADR2(DLX_IDinst_jtarget[17]),
    .ADR3(DLX_IDinst_jtarget[16]),
    .O(DLX_IDinst_Mcompar__n0102_inst_lut4_40)
  );
  defparam DLX_IDinst_Mcompar__n0102_inst_lut4_411.INIT = 16'h8241;
  X_LUT4 DLX_IDinst_Mcompar__n0102_inst_lut4_411 (
    .ADR0(DLX_reg_dst_of_EX[2]),
    .ADR1(DLX_reg_dst_of_EX[3]),
    .ADR2(DLX_IDinst_jtarget[19]),
    .ADR3(DLX_IDinst_jtarget[18]),
    .O(DLX_IDinst_Mcompar__n0102_inst_lut4_41)
  );
  X_BUF \DLX_IDinst_Mcompar__n0102_inst_cy_263/COUTUSED  (
    .I(\DLX_IDinst_Mcompar__n0102_inst_cy_263/CYMUXG ),
    .O(DLX_IDinst_Mcompar__n0102_inst_cy_263)
  );
  X_MUX2 DLX_IDinst_Mcompar__n0102_inst_cy_263_2623 (
    .IA(\DLX_IDinst_Mcompar__n0102_inst_cy_263/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mcompar__n0102_inst_cy_262),
    .SEL(DLX_IDinst_Mcompar__n0102_inst_lut4_41),
    .O(\DLX_IDinst_Mcompar__n0102_inst_cy_263/CYMUXG )
  );
  X_ZERO \DLX_IDinst__n0102/LOGIC_ZERO_2624  (
    .O(\DLX_IDinst__n0102/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mcompar__n0102_inst_cy_264 (
    .IA(\DLX_IDinst__n0102/LOGIC_ZERO ),
    .IB(\DLX_IDinst__n0102/CYINIT ),
    .SEL(DLX_IDinst_Mcompar__n0102_inst_lut4_42),
    .O(\DLX_IDinst__n0102/CYMUXF )
  );
  defparam DLX_IDinst_Mcompar__n0102_inst_lut4_421.INIT = 16'hE14B;
  X_LUT4 DLX_IDinst_Mcompar__n0102_inst_lut4_421 (
    .ADR0(DLX_EXinst__n0144),
    .ADR1(DLX_IDinst_current_IR[20]),
    .ADR2(DLX_reg_dst_of_EX[4]),
    .ADR3(DLX_IFinst_IR_latched[20]),
    .O(DLX_IDinst_Mcompar__n0102_inst_lut4_42)
  );
  X_BUF \DLX_IDinst__n0102/XBUSED  (
    .I(\DLX_IDinst__n0102/CYMUXF ),
    .O(DLX_IDinst__n0102)
  );
  X_BUF \DLX_IDinst__n0102/CYINIT_2625  (
    .I(DLX_IDinst_Mcompar__n0102_inst_cy_263),
    .O(\DLX_IDinst__n0102/CYINIT )
  );
  X_ONE \DLX_IDinst_RegFile_2_18/LOGIC_ONE_2626  (
    .O(\DLX_IDinst_RegFile_2_18/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_RegFile_2_18/LOGIC_ZERO_2627  (
    .O(\DLX_IDinst_RegFile_2_18/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0033_inst_cy_340_2628 (
    .IA(\DLX_IDinst_RegFile_2_18/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_2_18/LOGIC_ONE ),
    .SEL(vga_top_vga1_Mcompar__n0033_inst_lut1_4),
    .O(vga_top_vga1_Mcompar__n0033_inst_cy_340)
  );
  defparam vga_top_vga1_Mcompar__n0033_inst_lut1_41.INIT = 16'h5555;
  X_LUT4 vga_top_vga1_Mcompar__n0033_inst_lut1_41 (
    .ADR0(vga_top_vga1_hcounter[0]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(vga_top_vga1_Mcompar__n0033_inst_lut1_4)
  );
  defparam vga_top_vga1_Mcompar__n0033_inst_lut1_51.INIT = 16'h0F0F;
  X_LUT4 vga_top_vga1_Mcompar__n0033_inst_lut1_51 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_hcounter[0]),
    .ADR3(VCC),
    .O(vga_top_vga1_Mcompar__n0033_inst_lut1_5)
  );
  X_BUF \DLX_IDinst_RegFile_2_18/COUTUSED  (
    .I(\DLX_IDinst_RegFile_2_18/CYMUXG ),
    .O(vga_top_vga1_Mcompar__n0033_inst_cy_341)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0033_inst_cy_341_2629 (
    .IA(\DLX_IDinst_RegFile_2_18/LOGIC_ZERO ),
    .IB(vga_top_vga1_Mcompar__n0033_inst_cy_340),
    .SEL(vga_top_vga1_Mcompar__n0033_inst_lut1_5),
    .O(\DLX_IDinst_RegFile_2_18/CYMUXG )
  );
  X_ONE \vga_top_vga1_Mcompar__n0033_inst_cy_343/LOGIC_ONE_2630  (
    .O(\vga_top_vga1_Mcompar__n0033_inst_cy_343/LOGIC_ONE )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0033_inst_cy_342_2631 (
    .IA(\vga_top_vga1_Mcompar__n0033_inst_cy_343/LOGIC_ONE ),
    .IB(\vga_top_vga1_Mcompar__n0033_inst_cy_343/CYINIT ),
    .SEL(vga_top_vga1_Mcompar__n0033_inst_lut2_269),
    .O(vga_top_vga1_Mcompar__n0033_inst_cy_342)
  );
  defparam vga_top_vga1_Mcompar__n0033_inst_lut2_2691.INIT = 16'hAA00;
  X_LUT4 vga_top_vga1_Mcompar__n0033_inst_lut2_2691 (
    .ADR0(vga_top_vga1_hcounter[1]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[2]),
    .O(vga_top_vga1_Mcompar__n0033_inst_lut2_269)
  );
  defparam vga_top_vga1_Mcompar__n0033_inst_lut2_2701.INIT = 16'hAA00;
  X_LUT4 vga_top_vga1_Mcompar__n0033_inst_lut2_2701 (
    .ADR0(vga_top_vga1_hcounter[1]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[2]),
    .O(vga_top_vga1_Mcompar__n0033_inst_lut2_270)
  );
  X_BUF \vga_top_vga1_Mcompar__n0033_inst_cy_343/COUTUSED  (
    .I(\vga_top_vga1_Mcompar__n0033_inst_cy_343/CYMUXG ),
    .O(vga_top_vga1_Mcompar__n0033_inst_cy_343)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0033_inst_cy_343_2632 (
    .IA(\vga_top_vga1_Mcompar__n0033_inst_cy_343/LOGIC_ONE ),
    .IB(vga_top_vga1_Mcompar__n0033_inst_cy_342),
    .SEL(vga_top_vga1_Mcompar__n0033_inst_lut2_270),
    .O(\vga_top_vga1_Mcompar__n0033_inst_cy_343/CYMUXG )
  );
  X_BUF \vga_top_vga1_Mcompar__n0033_inst_cy_343/CYINIT_2633  (
    .I(vga_top_vga1_Mcompar__n0033_inst_cy_341),
    .O(\vga_top_vga1_Mcompar__n0033_inst_cy_343/CYINIT )
  );
  X_ZERO \vga_top_vga1_Mcompar__n0033_inst_cy_345/LOGIC_ZERO_2634  (
    .O(\vga_top_vga1_Mcompar__n0033_inst_cy_345/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0033_inst_cy_344_2635 (
    .IA(\vga_top_vga1_Mcompar__n0033_inst_cy_345/LOGIC_ZERO ),
    .IB(\vga_top_vga1_Mcompar__n0033_inst_cy_345/CYINIT ),
    .SEL(vga_top_vga1_Mcompar__n0033_inst_lut3_98),
    .O(vga_top_vga1_Mcompar__n0033_inst_cy_344)
  );
  defparam vga_top_vga1_Mcompar__n0033_inst_lut3_981.INIT = 16'h0101;
  X_LUT4 vga_top_vga1_Mcompar__n0033_inst_lut3_981 (
    .ADR0(vga_top_vga1_hcounter[4]),
    .ADR1(vga_top_vga1_hcounter[3]),
    .ADR2(vga_top_vga1_hcounter[5]),
    .ADR3(VCC),
    .O(vga_top_vga1_Mcompar__n0033_inst_lut3_98)
  );
  defparam vga_top_vga1_Mcompar__n0033_inst_lut3_991.INIT = 16'h0101;
  X_LUT4 vga_top_vga1_Mcompar__n0033_inst_lut3_991 (
    .ADR0(vga_top_vga1_hcounter[4]),
    .ADR1(vga_top_vga1_hcounter[3]),
    .ADR2(vga_top_vga1_hcounter[5]),
    .ADR3(VCC),
    .O(vga_top_vga1_Mcompar__n0033_inst_lut3_99)
  );
  X_BUF \vga_top_vga1_Mcompar__n0033_inst_cy_345/COUTUSED  (
    .I(\vga_top_vga1_Mcompar__n0033_inst_cy_345/CYMUXG ),
    .O(vga_top_vga1_Mcompar__n0033_inst_cy_345)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0033_inst_cy_345_2636 (
    .IA(\vga_top_vga1_Mcompar__n0033_inst_cy_345/LOGIC_ZERO ),
    .IB(vga_top_vga1_Mcompar__n0033_inst_cy_344),
    .SEL(vga_top_vga1_Mcompar__n0033_inst_lut3_99),
    .O(\vga_top_vga1_Mcompar__n0033_inst_cy_345/CYMUXG )
  );
  X_BUF \vga_top_vga1_Mcompar__n0033_inst_cy_345/CYINIT_2637  (
    .I(vga_top_vga1_Mcompar__n0033_inst_cy_343),
    .O(\vga_top_vga1_Mcompar__n0033_inst_cy_345/CYINIT )
  );
  X_ONE \vga_top_vga1_Mcompar__n0033_inst_cy_347/LOGIC_ONE_2638  (
    .O(\vga_top_vga1_Mcompar__n0033_inst_cy_347/LOGIC_ONE )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0033_inst_cy_346_2639 (
    .IA(\vga_top_vga1_Mcompar__n0033_inst_cy_347/LOGIC_ONE ),
    .IB(\vga_top_vga1_Mcompar__n0033_inst_cy_347/CYINIT ),
    .SEL(vga_top_vga1_Mcompar__n0033_inst_lut2_271),
    .O(vga_top_vga1_Mcompar__n0033_inst_cy_346)
  );
  defparam vga_top_vga1_Mcompar__n0033_inst_lut2_2711.INIT = 16'hAA00;
  X_LUT4 vga_top_vga1_Mcompar__n0033_inst_lut2_2711 (
    .ADR0(vga_top_vga1_hcounter[6]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[7]),
    .O(vga_top_vga1_Mcompar__n0033_inst_lut2_271)
  );
  defparam vga_top_vga1_Mcompar__n0033_inst_lut2_2721.INIT = 16'hA0A0;
  X_LUT4 vga_top_vga1_Mcompar__n0033_inst_lut2_2721 (
    .ADR0(vga_top_vga1_hcounter[6]),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_hcounter[7]),
    .ADR3(VCC),
    .O(vga_top_vga1_Mcompar__n0033_inst_lut2_272)
  );
  X_BUF \vga_top_vga1_Mcompar__n0033_inst_cy_347/COUTUSED  (
    .I(\vga_top_vga1_Mcompar__n0033_inst_cy_347/CYMUXG ),
    .O(vga_top_vga1_Mcompar__n0033_inst_cy_347)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0033_inst_cy_347_2640 (
    .IA(\vga_top_vga1_Mcompar__n0033_inst_cy_347/LOGIC_ONE ),
    .IB(vga_top_vga1_Mcompar__n0033_inst_cy_346),
    .SEL(vga_top_vga1_Mcompar__n0033_inst_lut2_272),
    .O(\vga_top_vga1_Mcompar__n0033_inst_cy_347/CYMUXG )
  );
  X_BUF \vga_top_vga1_Mcompar__n0033_inst_cy_347/CYINIT_2641  (
    .I(vga_top_vga1_Mcompar__n0033_inst_cy_345),
    .O(\vga_top_vga1_Mcompar__n0033_inst_cy_347/CYINIT )
  );
  X_ZERO \DLX_IFinst_IR_curr<25>/LOGIC_ZERO_2642  (
    .O(\DLX_IFinst_IR_curr<25>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0033_inst_cy_348_2643 (
    .IA(\DLX_IFinst_IR_curr<25>/LOGIC_ZERO ),
    .IB(\DLX_IFinst_IR_curr<25>/CYINIT ),
    .SEL(vga_top_vga1_Mcompar__n0033_inst_lut1_6),
    .O(vga_top_vga1_Mcompar__n0033_inst_cy_348)
  );
  defparam vga_top_vga1_Mcompar__n0033_inst_lut1_61.INIT = 16'h00FF;
  X_LUT4 vga_top_vga1_Mcompar__n0033_inst_lut1_61 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[8]),
    .O(vga_top_vga1_Mcompar__n0033_inst_lut1_6)
  );
  defparam vga_top_vga1_Mcompar__n0033_inst_lut1_71.INIT = 16'h00FF;
  X_LUT4 vga_top_vga1_Mcompar__n0033_inst_lut1_71 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(vga_top_vga1_hcounter[8]),
    .O(vga_top_vga1_Mcompar__n0033_inst_lut1_7)
  );
  X_BUF \DLX_IFinst_IR_curr<25>/COUTUSED  (
    .I(\DLX_IFinst_IR_curr<25>/CYMUXG ),
    .O(vga_top_vga1_Mcompar__n0033_inst_cy_349)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0033_inst_cy_349_2644 (
    .IA(\DLX_IFinst_IR_curr<25>/LOGIC_ZERO ),
    .IB(vga_top_vga1_Mcompar__n0033_inst_cy_348),
    .SEL(vga_top_vga1_Mcompar__n0033_inst_lut1_7),
    .O(\DLX_IFinst_IR_curr<25>/CYMUXG )
  );
  X_BUF \DLX_IFinst_IR_curr<25>/CYINIT_2645  (
    .I(vga_top_vga1_Mcompar__n0033_inst_cy_347),
    .O(\DLX_IFinst_IR_curr<25>/CYINIT )
  );
  X_ONE \vga_top_vga1_Mcompar__n0033_inst_cy_351/LOGIC_ONE_2646  (
    .O(\vga_top_vga1_Mcompar__n0033_inst_cy_351/LOGIC_ONE )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0033_inst_cy_350_2647 (
    .IA(\vga_top_vga1_Mcompar__n0033_inst_cy_351/LOGIC_ONE ),
    .IB(\vga_top_vga1_Mcompar__n0033_inst_cy_351/CYINIT ),
    .SEL(\$SIG_13 ),
    .O(vga_top_vga1_Mcompar__n0033_inst_cy_350)
  );
  defparam \$BEL_13 .INIT = 16'hCCCC;
  X_LUT4 \$BEL_13  (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_hcounter[9]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\$SIG_13 )
  );
  defparam \$BEL_14 .INIT = 16'hCCCC;
  X_LUT4 \$BEL_14  (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_hcounter[9]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\$SIG_14 )
  );
  X_BUF \vga_top_vga1_Mcompar__n0033_inst_cy_351/COUTUSED  (
    .I(\vga_top_vga1_Mcompar__n0033_inst_cy_351/CYMUXG ),
    .O(vga_top_vga1_Mcompar__n0033_inst_cy_351)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0033_inst_cy_351_2648 (
    .IA(\vga_top_vga1_Mcompar__n0033_inst_cy_351/LOGIC_ONE ),
    .IB(vga_top_vga1_Mcompar__n0033_inst_cy_350),
    .SEL(\$SIG_14 ),
    .O(\vga_top_vga1_Mcompar__n0033_inst_cy_351/CYMUXG )
  );
  X_BUF \vga_top_vga1_Mcompar__n0033_inst_cy_351/CYINIT_2649  (
    .I(vga_top_vga1_Mcompar__n0033_inst_cy_349),
    .O(\vga_top_vga1_Mcompar__n0033_inst_cy_351/CYINIT )
  );
  X_ZERO \vga_top_vga1__n0033/LOGIC_ZERO_2650  (
    .O(\vga_top_vga1__n0033/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_Mcompar__n0033_inst_cy_352_2651 (
    .IA(\vga_top_vga1__n0033/LOGIC_ZERO ),
    .IB(\vga_top_vga1__n0033/CYINIT ),
    .SEL(vga_top_vga1_Mcompar__n0033_inst_lut4_1100),
    .O(vga_top_vga1_Mcompar__n0033_inst_cy_352)
  );
  defparam vga_top_vga1_Mcompar__n0033_inst_lut4_11001.INIT = 16'h0001;
  X_LUT4 vga_top_vga1_Mcompar__n0033_inst_lut4_11001 (
    .ADR0(vga_top_vga1_hcounter[10]),
    .ADR1(vga_top_vga1_hcounter[11]),
    .ADR2(vga_top_vga1_hcounter[12]),
    .ADR3(vga_top_vga1_hcounter[13]),
    .O(vga_top_vga1_Mcompar__n0033_inst_lut4_1100)
  );
  defparam vga_top_vga1_Mcompar__n0033_inst_lut2_2731.INIT = 16'h1111;
  X_LUT4 vga_top_vga1_Mcompar__n0033_inst_lut2_2731 (
    .ADR0(vga_top_vga1_hcounter[14]),
    .ADR1(vga_top_vga1_hcounter[15]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(vga_top_vga1_Mcompar__n0033_inst_lut2_273)
  );
  X_BUF \vga_top_vga1__n0033/COUTUSED  (
    .I(\vga_top_vga1__n0033/CYMUXG ),
    .O(vga_top_vga1__n0033)
  );
  X_MUX2 vga_top_vga1_Mcompar__n0033_inst_cy_353 (
    .IA(\vga_top_vga1__n0033/LOGIC_ZERO ),
    .IB(vga_top_vga1_Mcompar__n0033_inst_cy_352),
    .SEL(vga_top_vga1_Mcompar__n0033_inst_lut2_273),
    .O(\vga_top_vga1__n0033/CYMUXG )
  );
  X_BUF \vga_top_vga1__n0033/CYINIT_2652  (
    .I(vga_top_vga1_Mcompar__n0033_inst_cy_351),
    .O(\vga_top_vga1__n0033/CYINIT )
  );
  X_ZERO \vga_top_vga1_Madd_addressout_inst_lut2_331/LOGIC_ZERO_2653  (
    .O(\vga_top_vga1_Madd_addressout_inst_lut2_331/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_Madd_addressout_inst_cy_462_2654 (
    .IA(vga_top_vga1_gridhcounter[5]),
    .IB(\vga_top_vga1_Madd_addressout_inst_lut2_331/LOGIC_ZERO ),
    .SEL(\vga_top_vga1_Madd_addressout_inst_lut2_331/FROM ),
    .O(vga_top_vga1_Madd_addressout_inst_cy_462)
  );
  defparam vga_top_vga1_Madd_addressout_inst_lut2_3311.INIT = 16'h5A5A;
  X_LUT4 vga_top_vga1_Madd_addressout_inst_lut2_3311 (
    .ADR0(vga_top_vga1_gridhcounter[5]),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_gridvcounter[0]),
    .ADR3(VCC),
    .O(\vga_top_vga1_Madd_addressout_inst_lut2_331/FROM )
  );
  defparam vga_top_vga1_Madd_addressout_inst_lut2_3321.INIT = 16'h5A5A;
  X_LUT4 vga_top_vga1_Madd_addressout_inst_lut2_3321 (
    .ADR0(vga_top_vga1_gridhcounter[6]),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_gridvcounter[1]),
    .ADR3(VCC),
    .O(vga_top_vga1_Madd_addressout_inst_lut2_332)
  );
  X_BUF \vga_top_vga1_Madd_addressout_inst_lut2_331/COUTUSED  (
    .I(\vga_top_vga1_Madd_addressout_inst_lut2_331/CYMUXG ),
    .O(vga_top_vga1_Madd_addressout_inst_cy_463)
  );
  X_BUF \vga_top_vga1_Madd_addressout_inst_lut2_331/XUSED  (
    .I(\vga_top_vga1_Madd_addressout_inst_lut2_331/FROM ),
    .O(vga_top_vga1_Madd_addressout_inst_lut2_331)
  );
  X_BUF \vga_top_vga1_Madd_addressout_inst_lut2_331/YUSED  (
    .I(\vga_top_vga1_Madd_addressout_inst_lut2_331/XORG ),
    .O(vga_address[6])
  );
  X_MUX2 vga_top_vga1_Madd_addressout_inst_cy_463_2655 (
    .IA(vga_top_vga1_gridhcounter[6]),
    .IB(vga_top_vga1_Madd_addressout_inst_cy_462),
    .SEL(vga_top_vga1_Madd_addressout_inst_lut2_332),
    .O(\vga_top_vga1_Madd_addressout_inst_lut2_331/CYMUXG )
  );
  X_XOR2 vga_top_vga1_Madd_addressout_inst_sum_254 (
    .I0(vga_top_vga1_Madd_addressout_inst_cy_462),
    .I1(vga_top_vga1_Madd_addressout_inst_lut2_332),
    .O(\vga_top_vga1_Madd_addressout_inst_lut2_331/XORG )
  );
  defparam DLX_IDinst_RegFile_29_18_2656.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_29_18_2656 (
    .I(DLX_IDinst_WB_data_eff[18]),
    .CE(DLX_IDinst__n0608),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_29_18)
  );
  X_MUX2 vga_top_vga1_Madd_addressout_inst_cy_464_2657 (
    .IA(vga_top_vga1_gridhcounter[7]),
    .IB(\vga_address<7>/CYINIT ),
    .SEL(vga_top_vga1_Madd_addressout_inst_lut2_333),
    .O(vga_top_vga1_Madd_addressout_inst_cy_464)
  );
  X_XOR2 vga_top_vga1_Madd_addressout_inst_sum_255 (
    .I0(\vga_address<7>/CYINIT ),
    .I1(vga_top_vga1_Madd_addressout_inst_lut2_333),
    .O(\vga_address<7>/XORF )
  );
  defparam vga_top_vga1_Madd_addressout_inst_lut2_3331.INIT = 16'h9696;
  X_LUT4 vga_top_vga1_Madd_addressout_inst_lut2_3331 (
    .ADR0(vga_top_vga1_gridhcounter[7]),
    .ADR1(vga_top_vga1_gridvcounter[0]),
    .ADR2(vga_top_vga1_gridvcounter[2]),
    .ADR3(VCC),
    .O(vga_top_vga1_Madd_addressout_inst_lut2_333)
  );
  defparam vga_top_vga1_Madd_addressout_inst_lut2_3341.INIT = 16'h5A5A;
  X_LUT4 vga_top_vga1_Madd_addressout_inst_lut2_3341 (
    .ADR0(vga_top_vga1_gridhcounter[8]),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_Mmult__n0043_inst_lut2_317),
    .ADR3(VCC),
    .O(vga_top_vga1_Madd_addressout_inst_lut2_334)
  );
  X_BUF \vga_address<7>/COUTUSED  (
    .I(\vga_address<7>/CYMUXG ),
    .O(vga_top_vga1_Madd_addressout_inst_cy_465)
  );
  X_BUF \vga_address<7>/XUSED  (
    .I(\vga_address<7>/XORF ),
    .O(vga_address[7])
  );
  X_BUF \vga_address<7>/YUSED  (
    .I(\vga_address<7>/XORG ),
    .O(vga_address[8])
  );
  X_MUX2 vga_top_vga1_Madd_addressout_inst_cy_465_2658 (
    .IA(vga_top_vga1_gridhcounter[8]),
    .IB(vga_top_vga1_Madd_addressout_inst_cy_464),
    .SEL(vga_top_vga1_Madd_addressout_inst_lut2_334),
    .O(\vga_address<7>/CYMUXG )
  );
  X_XOR2 vga_top_vga1_Madd_addressout_inst_sum_256 (
    .I0(vga_top_vga1_Madd_addressout_inst_cy_464),
    .I1(vga_top_vga1_Madd_addressout_inst_lut2_334),
    .O(\vga_address<7>/XORG )
  );
  X_BUF \vga_address<7>/CYINIT_2659  (
    .I(vga_top_vga1_Madd_addressout_inst_cy_463),
    .O(\vga_address<7>/CYINIT )
  );
  X_ZERO \vga_address<9>/LOGIC_ZERO_2660  (
    .O(\vga_address<9>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_Madd_addressout_inst_cy_466_2661 (
    .IA(\vga_address<9>/LOGIC_ZERO ),
    .IB(\vga_address<9>/CYINIT ),
    .SEL(\vga_address<9>/FROM ),
    .O(vga_top_vga1_Madd_addressout_inst_cy_466)
  );
  X_XOR2 vga_top_vga1_Madd_addressout_inst_sum_257 (
    .I0(\vga_address<9>/CYINIT ),
    .I1(\vga_address<9>/FROM ),
    .O(\vga_address<9>/XORF )
  );
  defparam \vga_address<9>/F .INIT = 16'hF0F0;
  X_LUT4 \vga_address<9>/F  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_Mmult__n0043_inst_lut2_318),
    .ADR3(VCC),
    .O(\vga_address<9>/FROM )
  );
  defparam \vga_address<9>/G .INIT = 16'hF0F0;
  X_LUT4 \vga_address<9>/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_Mmult__n0043_inst_lut2_319),
    .ADR3(VCC),
    .O(\vga_address<9>/GROM )
  );
  X_BUF \vga_address<9>/COUTUSED  (
    .I(\vga_address<9>/CYMUXG ),
    .O(vga_top_vga1_Madd_addressout_inst_cy_467)
  );
  X_BUF \vga_address<9>/XUSED  (
    .I(\vga_address<9>/XORF ),
    .O(vga_address[9])
  );
  X_BUF \vga_address<9>/YUSED  (
    .I(\vga_address<9>/XORG ),
    .O(vga_address[10])
  );
  X_MUX2 vga_top_vga1_Madd_addressout_inst_cy_467_2662 (
    .IA(\vga_address<9>/LOGIC_ZERO ),
    .IB(vga_top_vga1_Madd_addressout_inst_cy_466),
    .SEL(\vga_address<9>/GROM ),
    .O(\vga_address<9>/CYMUXG )
  );
  X_XOR2 vga_top_vga1_Madd_addressout_inst_sum_258 (
    .I0(vga_top_vga1_Madd_addressout_inst_cy_466),
    .I1(\vga_address<9>/GROM ),
    .O(\vga_address<9>/XORG )
  );
  X_BUF \vga_address<9>/CYINIT_2663  (
    .I(vga_top_vga1_Madd_addressout_inst_cy_465),
    .O(\vga_address<9>/CYINIT )
  );
  X_ZERO \vga_address<11>/LOGIC_ZERO_2664  (
    .O(\vga_address<11>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_Madd_addressout_inst_cy_468_2665 (
    .IA(\vga_address<11>/LOGIC_ZERO ),
    .IB(\vga_address<11>/CYINIT ),
    .SEL(\vga_address<11>/FROM ),
    .O(vga_top_vga1_Madd_addressout_inst_cy_468)
  );
  X_XOR2 vga_top_vga1_Madd_addressout_inst_sum_259 (
    .I0(\vga_address<11>/CYINIT ),
    .I1(\vga_address<11>/FROM ),
    .O(\vga_address<11>/XORF )
  );
  defparam \vga_address<11>/F .INIT = 16'hF0F0;
  X_LUT4 \vga_address<11>/F  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_Mmult__n0043_inst_lut2_320),
    .ADR3(VCC),
    .O(\vga_address<11>/FROM )
  );
  defparam \vga_address<11>/G .INIT = 16'hCCCC;
  X_LUT4 \vga_address<11>/G  (
    .ADR0(VCC),
    .ADR1(vga_top_vga1_Mmult__n0043_inst_lut2_321),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\vga_address<11>/GROM )
  );
  X_BUF \vga_address<11>/COUTUSED  (
    .I(\vga_address<11>/CYMUXG ),
    .O(vga_top_vga1_Madd_addressout_inst_cy_469)
  );
  X_BUF \vga_address<11>/XUSED  (
    .I(\vga_address<11>/XORF ),
    .O(vga_address[11])
  );
  X_BUF \vga_address<11>/YUSED  (
    .I(\vga_address<11>/XORG ),
    .O(vga_address[12])
  );
  X_MUX2 vga_top_vga1_Madd_addressout_inst_cy_469_2666 (
    .IA(\vga_address<11>/LOGIC_ZERO ),
    .IB(vga_top_vga1_Madd_addressout_inst_cy_468),
    .SEL(\vga_address<11>/GROM ),
    .O(\vga_address<11>/CYMUXG )
  );
  X_XOR2 vga_top_vga1_Madd_addressout_inst_sum_260 (
    .I0(vga_top_vga1_Madd_addressout_inst_cy_468),
    .I1(\vga_address<11>/GROM ),
    .O(\vga_address<11>/XORG )
  );
  X_BUF \vga_address<11>/CYINIT_2667  (
    .I(vga_top_vga1_Madd_addressout_inst_cy_467),
    .O(\vga_address<11>/CYINIT )
  );
  X_ZERO \vga_address<13>/LOGIC_ZERO_2668  (
    .O(\vga_address<13>/LOGIC_ZERO )
  );
  X_MUX2 vga_top_vga1_Madd_addressout_inst_cy_470_2669 (
    .IA(\vga_address<13>/LOGIC_ZERO ),
    .IB(\vga_address<13>/CYINIT ),
    .SEL(\vga_address<13>/FROM ),
    .O(vga_top_vga1_Madd_addressout_inst_cy_470)
  );
  X_XOR2 vga_top_vga1_Madd_addressout_inst_sum_261 (
    .I0(\vga_address<13>/CYINIT ),
    .I1(\vga_address<13>/FROM ),
    .O(\vga_address<13>/XORF )
  );
  defparam \vga_address<13>/F .INIT = 16'hF0F0;
  X_LUT4 \vga_address<13>/F  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_Mmult__n0043_inst_lut2_322),
    .ADR3(VCC),
    .O(\vga_address<13>/FROM )
  );
  defparam vga_top_vga1_Mmult__n0043_inst_lut2_323_rt_2670.INIT = 16'hF0F0;
  X_LUT4 vga_top_vga1_Mmult__n0043_inst_lut2_323_rt_2670 (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(vga_top_vga1_Mmult__n0043_inst_lut2_323),
    .ADR3(VCC),
    .O(vga_top_vga1_Mmult__n0043_inst_lut2_323_rt)
  );
  X_BUF \vga_address<13>/XUSED  (
    .I(\vga_address<13>/XORF ),
    .O(vga_address[13])
  );
  X_BUF \vga_address<13>/YUSED  (
    .I(\vga_address<13>/XORG ),
    .O(vga_address[14])
  );
  X_XOR2 vga_top_vga1_Madd_addressout_inst_sum_262 (
    .I0(vga_top_vga1_Madd_addressout_inst_cy_470),
    .I1(vga_top_vga1_Mmult__n0043_inst_lut2_323_rt),
    .O(\vga_address<13>/XORG )
  );
  X_BUF \vga_address<13>/CYINIT_2671  (
    .I(vga_top_vga1_Madd_addressout_inst_cy_469),
    .O(\vga_address<13>/CYINIT )
  );
  X_ZERO \DLX_IFinst__n0015<3>/LOGIC_ZERO_2672  (
    .O(\DLX_IFinst__n0015<3>/LOGIC_ZERO )
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_40_2673 (
    .IA(GLOBAL_LOGIC1),
    .IB(\DLX_IFinst__n0015<3>/LOGIC_ZERO ),
    .SEL(DLX_IFinst_Madd__n0005_inst_lut2_40),
    .O(DLX_IFinst_Madd__n0005_inst_cy_40)
  );
  defparam DLX_IFinst_Madd__n0005_inst_lut2_401.INIT = 16'h00FF;
  X_LUT4 DLX_IFinst_Madd__n0005_inst_lut2_401 (
    .ADR0(GLOBAL_LOGIC1),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IFinst_NPC[2]),
    .O(DLX_IFinst_Madd__n0005_inst_lut2_40)
  );
  defparam \DLX_IFinst__n0015<3>/G .INIT = 16'hFF00;
  X_LUT4 \DLX_IFinst__n0015<3>/G  (
    .ADR0(GLOBAL_LOGIC0),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IFinst_NPC[3]),
    .O(\DLX_IFinst__n0015<3>/GROM )
  );
  X_BUF \DLX_IFinst__n0015<3>/COUTUSED  (
    .I(\DLX_IFinst__n0015<3>/CYMUXG ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_41)
  );
  X_BUF \DLX_IFinst__n0015<3>/YUSED  (
    .I(\DLX_IFinst__n0015<3>/XORG ),
    .O(DLX_IFinst__n0015[3])
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_41_2674 (
    .IA(GLOBAL_LOGIC0),
    .IB(DLX_IFinst_Madd__n0005_inst_cy_40),
    .SEL(\DLX_IFinst__n0015<3>/GROM ),
    .O(\DLX_IFinst__n0015<3>/CYMUXG )
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_41 (
    .I0(DLX_IFinst_Madd__n0005_inst_cy_40),
    .I1(\DLX_IFinst__n0015<3>/GROM ),
    .O(\DLX_IFinst__n0015<3>/XORG )
  );
  X_ZERO \DLX_IFinst__n0015<4>/LOGIC_ZERO_2675  (
    .O(\DLX_IFinst__n0015<4>/LOGIC_ZERO )
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_42_2676 (
    .IA(\DLX_IFinst__n0015<4>/LOGIC_ZERO ),
    .IB(\DLX_IFinst__n0015<4>/CYINIT ),
    .SEL(\DLX_IFinst__n0015<4>/FROM ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_42)
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_42 (
    .I0(\DLX_IFinst__n0015<4>/CYINIT ),
    .I1(\DLX_IFinst__n0015<4>/FROM ),
    .O(\DLX_IFinst__n0015<4>/XORF )
  );
  defparam \DLX_IFinst__n0015<4>/F .INIT = 16'hCCCC;
  X_LUT4 \DLX_IFinst__n0015<4>/F  (
    .ADR0(VCC),
    .ADR1(DLX_IFinst_NPC[4]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IFinst__n0015<4>/FROM )
  );
  defparam \DLX_IFinst__n0015<4>/G .INIT = 16'hCCCC;
  X_LUT4 \DLX_IFinst__n0015<4>/G  (
    .ADR0(VCC),
    .ADR1(DLX_IFinst_NPC[5]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IFinst__n0015<4>/GROM )
  );
  X_BUF \DLX_IFinst__n0015<4>/COUTUSED  (
    .I(\DLX_IFinst__n0015<4>/CYMUXG ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_43)
  );
  X_BUF \DLX_IFinst__n0015<4>/XUSED  (
    .I(\DLX_IFinst__n0015<4>/XORF ),
    .O(DLX_IFinst__n0015[4])
  );
  X_BUF \DLX_IFinst__n0015<4>/YUSED  (
    .I(\DLX_IFinst__n0015<4>/XORG ),
    .O(DLX_IFinst__n0015[5])
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_43_2677 (
    .IA(\DLX_IFinst__n0015<4>/LOGIC_ZERO ),
    .IB(DLX_IFinst_Madd__n0005_inst_cy_42),
    .SEL(\DLX_IFinst__n0015<4>/GROM ),
    .O(\DLX_IFinst__n0015<4>/CYMUXG )
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_43 (
    .I0(DLX_IFinst_Madd__n0005_inst_cy_42),
    .I1(\DLX_IFinst__n0015<4>/GROM ),
    .O(\DLX_IFinst__n0015<4>/XORG )
  );
  X_BUF \DLX_IFinst__n0015<4>/CYINIT_2678  (
    .I(DLX_IFinst_Madd__n0005_inst_cy_41),
    .O(\DLX_IFinst__n0015<4>/CYINIT )
  );
  X_ZERO \DLX_IFinst__n0015<6>/LOGIC_ZERO_2679  (
    .O(\DLX_IFinst__n0015<6>/LOGIC_ZERO )
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_44_2680 (
    .IA(\DLX_IFinst__n0015<6>/LOGIC_ZERO ),
    .IB(\DLX_IFinst__n0015<6>/CYINIT ),
    .SEL(\DLX_IFinst__n0015<6>/FROM ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_44)
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_44 (
    .I0(\DLX_IFinst__n0015<6>/CYINIT ),
    .I1(\DLX_IFinst__n0015<6>/FROM ),
    .O(\DLX_IFinst__n0015<6>/XORF )
  );
  defparam \DLX_IFinst__n0015<6>/F .INIT = 16'hAAAA;
  X_LUT4 \DLX_IFinst__n0015<6>/F  (
    .ADR0(DLX_IFinst_NPC[6]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IFinst__n0015<6>/FROM )
  );
  defparam \DLX_IFinst__n0015<6>/G .INIT = 16'hF0F0;
  X_LUT4 \DLX_IFinst__n0015<6>/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IFinst_NPC[7]),
    .ADR3(VCC),
    .O(\DLX_IFinst__n0015<6>/GROM )
  );
  X_BUF \DLX_IFinst__n0015<6>/COUTUSED  (
    .I(\DLX_IFinst__n0015<6>/CYMUXG ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_45)
  );
  X_BUF \DLX_IFinst__n0015<6>/XUSED  (
    .I(\DLX_IFinst__n0015<6>/XORF ),
    .O(DLX_IFinst__n0015[6])
  );
  X_BUF \DLX_IFinst__n0015<6>/YUSED  (
    .I(\DLX_IFinst__n0015<6>/XORG ),
    .O(DLX_IFinst__n0015[7])
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_45_2681 (
    .IA(\DLX_IFinst__n0015<6>/LOGIC_ZERO ),
    .IB(DLX_IFinst_Madd__n0005_inst_cy_44),
    .SEL(\DLX_IFinst__n0015<6>/GROM ),
    .O(\DLX_IFinst__n0015<6>/CYMUXG )
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_45 (
    .I0(DLX_IFinst_Madd__n0005_inst_cy_44),
    .I1(\DLX_IFinst__n0015<6>/GROM ),
    .O(\DLX_IFinst__n0015<6>/XORG )
  );
  X_BUF \DLX_IFinst__n0015<6>/CYINIT_2682  (
    .I(DLX_IFinst_Madd__n0005_inst_cy_43),
    .O(\DLX_IFinst__n0015<6>/CYINIT )
  );
  X_ZERO \DLX_IFinst__n0015<8>/LOGIC_ZERO_2683  (
    .O(\DLX_IFinst__n0015<8>/LOGIC_ZERO )
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_46_2684 (
    .IA(\DLX_IFinst__n0015<8>/LOGIC_ZERO ),
    .IB(\DLX_IFinst__n0015<8>/CYINIT ),
    .SEL(\DLX_IFinst__n0015<8>/FROM ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_46)
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_46 (
    .I0(\DLX_IFinst__n0015<8>/CYINIT ),
    .I1(\DLX_IFinst__n0015<8>/FROM ),
    .O(\DLX_IFinst__n0015<8>/XORF )
  );
  defparam \DLX_IFinst__n0015<8>/F .INIT = 16'hFF00;
  X_LUT4 \DLX_IFinst__n0015<8>/F  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IFinst_NPC[8]),
    .O(\DLX_IFinst__n0015<8>/FROM )
  );
  defparam \DLX_IFinst__n0015<8>/G .INIT = 16'hAAAA;
  X_LUT4 \DLX_IFinst__n0015<8>/G  (
    .ADR0(DLX_IFinst_NPC[9]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IFinst__n0015<8>/GROM )
  );
  X_BUF \DLX_IFinst__n0015<8>/COUTUSED  (
    .I(\DLX_IFinst__n0015<8>/CYMUXG ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_47)
  );
  X_BUF \DLX_IFinst__n0015<8>/XUSED  (
    .I(\DLX_IFinst__n0015<8>/XORF ),
    .O(DLX_IFinst__n0015[8])
  );
  X_BUF \DLX_IFinst__n0015<8>/YUSED  (
    .I(\DLX_IFinst__n0015<8>/XORG ),
    .O(DLX_IFinst__n0015[9])
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_47_2685 (
    .IA(\DLX_IFinst__n0015<8>/LOGIC_ZERO ),
    .IB(DLX_IFinst_Madd__n0005_inst_cy_46),
    .SEL(\DLX_IFinst__n0015<8>/GROM ),
    .O(\DLX_IFinst__n0015<8>/CYMUXG )
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_47 (
    .I0(DLX_IFinst_Madd__n0005_inst_cy_46),
    .I1(\DLX_IFinst__n0015<8>/GROM ),
    .O(\DLX_IFinst__n0015<8>/XORG )
  );
  X_BUF \DLX_IFinst__n0015<8>/CYINIT_2686  (
    .I(DLX_IFinst_Madd__n0005_inst_cy_45),
    .O(\DLX_IFinst__n0015<8>/CYINIT )
  );
  X_ZERO \DLX_IFinst__n0015<10>/LOGIC_ZERO_2687  (
    .O(\DLX_IFinst__n0015<10>/LOGIC_ZERO )
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_48_2688 (
    .IA(\DLX_IFinst__n0015<10>/LOGIC_ZERO ),
    .IB(\DLX_IFinst__n0015<10>/CYINIT ),
    .SEL(\DLX_IFinst__n0015<10>/FROM ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_48)
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_48 (
    .I0(\DLX_IFinst__n0015<10>/CYINIT ),
    .I1(\DLX_IFinst__n0015<10>/FROM ),
    .O(\DLX_IFinst__n0015<10>/XORF )
  );
  defparam \DLX_IFinst__n0015<10>/F .INIT = 16'hFF00;
  X_LUT4 \DLX_IFinst__n0015<10>/F  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IFinst_NPC[10]),
    .O(\DLX_IFinst__n0015<10>/FROM )
  );
  defparam \DLX_IFinst__n0015<10>/G .INIT = 16'hAAAA;
  X_LUT4 \DLX_IFinst__n0015<10>/G  (
    .ADR0(DLX_IFinst_NPC[11]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IFinst__n0015<10>/GROM )
  );
  X_BUF \DLX_IFinst__n0015<10>/COUTUSED  (
    .I(\DLX_IFinst__n0015<10>/CYMUXG ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_49)
  );
  X_BUF \DLX_IFinst__n0015<10>/XUSED  (
    .I(\DLX_IFinst__n0015<10>/XORF ),
    .O(DLX_IFinst__n0015[10])
  );
  X_BUF \DLX_IFinst__n0015<10>/YUSED  (
    .I(\DLX_IFinst__n0015<10>/XORG ),
    .O(DLX_IFinst__n0015[11])
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_49_2689 (
    .IA(\DLX_IFinst__n0015<10>/LOGIC_ZERO ),
    .IB(DLX_IFinst_Madd__n0005_inst_cy_48),
    .SEL(\DLX_IFinst__n0015<10>/GROM ),
    .O(\DLX_IFinst__n0015<10>/CYMUXG )
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_49 (
    .I0(DLX_IFinst_Madd__n0005_inst_cy_48),
    .I1(\DLX_IFinst__n0015<10>/GROM ),
    .O(\DLX_IFinst__n0015<10>/XORG )
  );
  X_BUF \DLX_IFinst__n0015<10>/CYINIT_2690  (
    .I(DLX_IFinst_Madd__n0005_inst_cy_47),
    .O(\DLX_IFinst__n0015<10>/CYINIT )
  );
  X_ZERO \DLX_IFinst__n0015<12>/LOGIC_ZERO_2691  (
    .O(\DLX_IFinst__n0015<12>/LOGIC_ZERO )
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_50_2692 (
    .IA(\DLX_IFinst__n0015<12>/LOGIC_ZERO ),
    .IB(\DLX_IFinst__n0015<12>/CYINIT ),
    .SEL(\DLX_IFinst__n0015<12>/FROM ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_50)
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_50 (
    .I0(\DLX_IFinst__n0015<12>/CYINIT ),
    .I1(\DLX_IFinst__n0015<12>/FROM ),
    .O(\DLX_IFinst__n0015<12>/XORF )
  );
  defparam \DLX_IFinst__n0015<12>/F .INIT = 16'hAAAA;
  X_LUT4 \DLX_IFinst__n0015<12>/F  (
    .ADR0(DLX_IFinst_NPC[12]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IFinst__n0015<12>/FROM )
  );
  defparam \DLX_IFinst__n0015<12>/G .INIT = 16'hF0F0;
  X_LUT4 \DLX_IFinst__n0015<12>/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IFinst_NPC[13]),
    .ADR3(VCC),
    .O(\DLX_IFinst__n0015<12>/GROM )
  );
  X_BUF \DLX_IFinst__n0015<12>/COUTUSED  (
    .I(\DLX_IFinst__n0015<12>/CYMUXG ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_51)
  );
  X_BUF \DLX_IFinst__n0015<12>/XUSED  (
    .I(\DLX_IFinst__n0015<12>/XORF ),
    .O(DLX_IFinst__n0015[12])
  );
  X_BUF \DLX_IFinst__n0015<12>/YUSED  (
    .I(\DLX_IFinst__n0015<12>/XORG ),
    .O(DLX_IFinst__n0015[13])
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_51_2693 (
    .IA(\DLX_IFinst__n0015<12>/LOGIC_ZERO ),
    .IB(DLX_IFinst_Madd__n0005_inst_cy_50),
    .SEL(\DLX_IFinst__n0015<12>/GROM ),
    .O(\DLX_IFinst__n0015<12>/CYMUXG )
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_51 (
    .I0(DLX_IFinst_Madd__n0005_inst_cy_50),
    .I1(\DLX_IFinst__n0015<12>/GROM ),
    .O(\DLX_IFinst__n0015<12>/XORG )
  );
  X_BUF \DLX_IFinst__n0015<12>/CYINIT_2694  (
    .I(DLX_IFinst_Madd__n0005_inst_cy_49),
    .O(\DLX_IFinst__n0015<12>/CYINIT )
  );
  X_ZERO \DLX_IFinst__n0015<14>/LOGIC_ZERO_2695  (
    .O(\DLX_IFinst__n0015<14>/LOGIC_ZERO )
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_52_2696 (
    .IA(\DLX_IFinst__n0015<14>/LOGIC_ZERO ),
    .IB(\DLX_IFinst__n0015<14>/CYINIT ),
    .SEL(\DLX_IFinst__n0015<14>/FROM ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_52)
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_52 (
    .I0(\DLX_IFinst__n0015<14>/CYINIT ),
    .I1(\DLX_IFinst__n0015<14>/FROM ),
    .O(\DLX_IFinst__n0015<14>/XORF )
  );
  defparam \DLX_IFinst__n0015<14>/F .INIT = 16'hAAAA;
  X_LUT4 \DLX_IFinst__n0015<14>/F  (
    .ADR0(DLX_IFinst_NPC[14]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IFinst__n0015<14>/FROM )
  );
  defparam \DLX_IFinst__n0015<14>/G .INIT = 16'hAAAA;
  X_LUT4 \DLX_IFinst__n0015<14>/G  (
    .ADR0(DLX_IFinst_NPC[15]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IFinst__n0015<14>/GROM )
  );
  X_BUF \DLX_IFinst__n0015<14>/COUTUSED  (
    .I(\DLX_IFinst__n0015<14>/CYMUXG ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_53)
  );
  X_BUF \DLX_IFinst__n0015<14>/XUSED  (
    .I(\DLX_IFinst__n0015<14>/XORF ),
    .O(DLX_IFinst__n0015[14])
  );
  X_BUF \DLX_IFinst__n0015<14>/YUSED  (
    .I(\DLX_IFinst__n0015<14>/XORG ),
    .O(DLX_IFinst__n0015[15])
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_53_2697 (
    .IA(\DLX_IFinst__n0015<14>/LOGIC_ZERO ),
    .IB(DLX_IFinst_Madd__n0005_inst_cy_52),
    .SEL(\DLX_IFinst__n0015<14>/GROM ),
    .O(\DLX_IFinst__n0015<14>/CYMUXG )
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_53 (
    .I0(DLX_IFinst_Madd__n0005_inst_cy_52),
    .I1(\DLX_IFinst__n0015<14>/GROM ),
    .O(\DLX_IFinst__n0015<14>/XORG )
  );
  X_BUF \DLX_IFinst__n0015<14>/CYINIT_2698  (
    .I(DLX_IFinst_Madd__n0005_inst_cy_51),
    .O(\DLX_IFinst__n0015<14>/CYINIT )
  );
  X_ZERO \DLX_IFinst__n0015<16>/LOGIC_ZERO_2699  (
    .O(\DLX_IFinst__n0015<16>/LOGIC_ZERO )
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_54_2700 (
    .IA(\DLX_IFinst__n0015<16>/LOGIC_ZERO ),
    .IB(\DLX_IFinst__n0015<16>/CYINIT ),
    .SEL(\DLX_IFinst__n0015<16>/FROM ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_54)
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_54 (
    .I0(\DLX_IFinst__n0015<16>/CYINIT ),
    .I1(\DLX_IFinst__n0015<16>/FROM ),
    .O(\DLX_IFinst__n0015<16>/XORF )
  );
  defparam \DLX_IFinst__n0015<16>/F .INIT = 16'hAAAA;
  X_LUT4 \DLX_IFinst__n0015<16>/F  (
    .ADR0(DLX_IFinst_NPC[16]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IFinst__n0015<16>/FROM )
  );
  defparam \DLX_IFinst__n0015<16>/G .INIT = 16'hCCCC;
  X_LUT4 \DLX_IFinst__n0015<16>/G  (
    .ADR0(VCC),
    .ADR1(DLX_IFinst_NPC[17]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IFinst__n0015<16>/GROM )
  );
  X_BUF \DLX_IFinst__n0015<16>/COUTUSED  (
    .I(\DLX_IFinst__n0015<16>/CYMUXG ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_55)
  );
  X_BUF \DLX_IFinst__n0015<16>/XUSED  (
    .I(\DLX_IFinst__n0015<16>/XORF ),
    .O(DLX_IFinst__n0015[16])
  );
  X_BUF \DLX_IFinst__n0015<16>/YUSED  (
    .I(\DLX_IFinst__n0015<16>/XORG ),
    .O(DLX_IFinst__n0015[17])
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_55_2701 (
    .IA(\DLX_IFinst__n0015<16>/LOGIC_ZERO ),
    .IB(DLX_IFinst_Madd__n0005_inst_cy_54),
    .SEL(\DLX_IFinst__n0015<16>/GROM ),
    .O(\DLX_IFinst__n0015<16>/CYMUXG )
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_55 (
    .I0(DLX_IFinst_Madd__n0005_inst_cy_54),
    .I1(\DLX_IFinst__n0015<16>/GROM ),
    .O(\DLX_IFinst__n0015<16>/XORG )
  );
  X_BUF \DLX_IFinst__n0015<16>/CYINIT_2702  (
    .I(DLX_IFinst_Madd__n0005_inst_cy_53),
    .O(\DLX_IFinst__n0015<16>/CYINIT )
  );
  defparam DLX_IDinst_RegFile_29_27_2703.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_29_27_2703 (
    .I(DLX_IDinst_WB_data_eff[27]),
    .CE(DLX_IDinst__n0608),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_29_27)
  );
  X_ZERO \DLX_IFinst__n0015<18>/LOGIC_ZERO_2704  (
    .O(\DLX_IFinst__n0015<18>/LOGIC_ZERO )
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_56_2705 (
    .IA(\DLX_IFinst__n0015<18>/LOGIC_ZERO ),
    .IB(\DLX_IFinst__n0015<18>/CYINIT ),
    .SEL(\DLX_IFinst__n0015<18>/FROM ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_56)
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_56 (
    .I0(\DLX_IFinst__n0015<18>/CYINIT ),
    .I1(\DLX_IFinst__n0015<18>/FROM ),
    .O(\DLX_IFinst__n0015<18>/XORF )
  );
  defparam \DLX_IFinst__n0015<18>/F .INIT = 16'hF0F0;
  X_LUT4 \DLX_IFinst__n0015<18>/F  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IFinst_NPC[18]),
    .ADR3(VCC),
    .O(\DLX_IFinst__n0015<18>/FROM )
  );
  defparam \DLX_IFinst__n0015<18>/G .INIT = 16'hFF00;
  X_LUT4 \DLX_IFinst__n0015<18>/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IFinst_NPC[19]),
    .O(\DLX_IFinst__n0015<18>/GROM )
  );
  X_BUF \DLX_IFinst__n0015<18>/COUTUSED  (
    .I(\DLX_IFinst__n0015<18>/CYMUXG ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_57)
  );
  X_BUF \DLX_IFinst__n0015<18>/XUSED  (
    .I(\DLX_IFinst__n0015<18>/XORF ),
    .O(DLX_IFinst__n0015[18])
  );
  X_BUF \DLX_IFinst__n0015<18>/YUSED  (
    .I(\DLX_IFinst__n0015<18>/XORG ),
    .O(DLX_IFinst__n0015[19])
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_57_2706 (
    .IA(\DLX_IFinst__n0015<18>/LOGIC_ZERO ),
    .IB(DLX_IFinst_Madd__n0005_inst_cy_56),
    .SEL(\DLX_IFinst__n0015<18>/GROM ),
    .O(\DLX_IFinst__n0015<18>/CYMUXG )
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_57 (
    .I0(DLX_IFinst_Madd__n0005_inst_cy_56),
    .I1(\DLX_IFinst__n0015<18>/GROM ),
    .O(\DLX_IFinst__n0015<18>/XORG )
  );
  X_BUF \DLX_IFinst__n0015<18>/CYINIT_2707  (
    .I(DLX_IFinst_Madd__n0005_inst_cy_55),
    .O(\DLX_IFinst__n0015<18>/CYINIT )
  );
  X_ZERO \DLX_IFinst__n0015<20>/LOGIC_ZERO_2708  (
    .O(\DLX_IFinst__n0015<20>/LOGIC_ZERO )
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_58_2709 (
    .IA(\DLX_IFinst__n0015<20>/LOGIC_ZERO ),
    .IB(\DLX_IFinst__n0015<20>/CYINIT ),
    .SEL(\DLX_IFinst__n0015<20>/FROM ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_58)
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_58 (
    .I0(\DLX_IFinst__n0015<20>/CYINIT ),
    .I1(\DLX_IFinst__n0015<20>/FROM ),
    .O(\DLX_IFinst__n0015<20>/XORF )
  );
  defparam \DLX_IFinst__n0015<20>/F .INIT = 16'hCCCC;
  X_LUT4 \DLX_IFinst__n0015<20>/F  (
    .ADR0(VCC),
    .ADR1(DLX_IFinst_NPC[20]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IFinst__n0015<20>/FROM )
  );
  defparam \DLX_IFinst__n0015<20>/G .INIT = 16'hFF00;
  X_LUT4 \DLX_IFinst__n0015<20>/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IFinst_NPC[21]),
    .O(\DLX_IFinst__n0015<20>/GROM )
  );
  X_BUF \DLX_IFinst__n0015<20>/COUTUSED  (
    .I(\DLX_IFinst__n0015<20>/CYMUXG ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_59)
  );
  X_BUF \DLX_IFinst__n0015<20>/XUSED  (
    .I(\DLX_IFinst__n0015<20>/XORF ),
    .O(DLX_IFinst__n0015[20])
  );
  X_BUF \DLX_IFinst__n0015<20>/YUSED  (
    .I(\DLX_IFinst__n0015<20>/XORG ),
    .O(DLX_IFinst__n0015[21])
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_59_2710 (
    .IA(\DLX_IFinst__n0015<20>/LOGIC_ZERO ),
    .IB(DLX_IFinst_Madd__n0005_inst_cy_58),
    .SEL(\DLX_IFinst__n0015<20>/GROM ),
    .O(\DLX_IFinst__n0015<20>/CYMUXG )
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_59 (
    .I0(DLX_IFinst_Madd__n0005_inst_cy_58),
    .I1(\DLX_IFinst__n0015<20>/GROM ),
    .O(\DLX_IFinst__n0015<20>/XORG )
  );
  X_BUF \DLX_IFinst__n0015<20>/CYINIT_2711  (
    .I(DLX_IFinst_Madd__n0005_inst_cy_57),
    .O(\DLX_IFinst__n0015<20>/CYINIT )
  );
  X_ZERO \DLX_IFinst__n0015<22>/LOGIC_ZERO_2712  (
    .O(\DLX_IFinst__n0015<22>/LOGIC_ZERO )
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_60_2713 (
    .IA(\DLX_IFinst__n0015<22>/LOGIC_ZERO ),
    .IB(\DLX_IFinst__n0015<22>/CYINIT ),
    .SEL(\DLX_IFinst__n0015<22>/FROM ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_60)
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_60 (
    .I0(\DLX_IFinst__n0015<22>/CYINIT ),
    .I1(\DLX_IFinst__n0015<22>/FROM ),
    .O(\DLX_IFinst__n0015<22>/XORF )
  );
  defparam \DLX_IFinst__n0015<22>/F .INIT = 16'hFF00;
  X_LUT4 \DLX_IFinst__n0015<22>/F  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IFinst_NPC[22]),
    .O(\DLX_IFinst__n0015<22>/FROM )
  );
  defparam \DLX_IFinst__n0015<22>/G .INIT = 16'hAAAA;
  X_LUT4 \DLX_IFinst__n0015<22>/G  (
    .ADR0(DLX_IFinst_NPC[23]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IFinst__n0015<22>/GROM )
  );
  X_BUF \DLX_IFinst__n0015<22>/COUTUSED  (
    .I(\DLX_IFinst__n0015<22>/CYMUXG ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_61)
  );
  X_BUF \DLX_IFinst__n0015<22>/XUSED  (
    .I(\DLX_IFinst__n0015<22>/XORF ),
    .O(DLX_IFinst__n0015[22])
  );
  X_BUF \DLX_IFinst__n0015<22>/YUSED  (
    .I(\DLX_IFinst__n0015<22>/XORG ),
    .O(DLX_IFinst__n0015[23])
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_61_2714 (
    .IA(\DLX_IFinst__n0015<22>/LOGIC_ZERO ),
    .IB(DLX_IFinst_Madd__n0005_inst_cy_60),
    .SEL(\DLX_IFinst__n0015<22>/GROM ),
    .O(\DLX_IFinst__n0015<22>/CYMUXG )
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_61 (
    .I0(DLX_IFinst_Madd__n0005_inst_cy_60),
    .I1(\DLX_IFinst__n0015<22>/GROM ),
    .O(\DLX_IFinst__n0015<22>/XORG )
  );
  X_BUF \DLX_IFinst__n0015<22>/CYINIT_2715  (
    .I(DLX_IFinst_Madd__n0005_inst_cy_59),
    .O(\DLX_IFinst__n0015<22>/CYINIT )
  );
  X_ZERO \DLX_IFinst__n0015<24>/LOGIC_ZERO_2716  (
    .O(\DLX_IFinst__n0015<24>/LOGIC_ZERO )
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_62_2717 (
    .IA(\DLX_IFinst__n0015<24>/LOGIC_ZERO ),
    .IB(\DLX_IFinst__n0015<24>/CYINIT ),
    .SEL(\DLX_IFinst__n0015<24>/FROM ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_62)
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_62 (
    .I0(\DLX_IFinst__n0015<24>/CYINIT ),
    .I1(\DLX_IFinst__n0015<24>/FROM ),
    .O(\DLX_IFinst__n0015<24>/XORF )
  );
  defparam \DLX_IFinst__n0015<24>/F .INIT = 16'hFF00;
  X_LUT4 \DLX_IFinst__n0015<24>/F  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IFinst_NPC[24]),
    .O(\DLX_IFinst__n0015<24>/FROM )
  );
  defparam \DLX_IFinst__n0015<24>/G .INIT = 16'hCCCC;
  X_LUT4 \DLX_IFinst__n0015<24>/G  (
    .ADR0(VCC),
    .ADR1(DLX_IFinst_NPC[25]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IFinst__n0015<24>/GROM )
  );
  X_BUF \DLX_IFinst__n0015<24>/COUTUSED  (
    .I(\DLX_IFinst__n0015<24>/CYMUXG ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_63)
  );
  X_BUF \DLX_IFinst__n0015<24>/XUSED  (
    .I(\DLX_IFinst__n0015<24>/XORF ),
    .O(DLX_IFinst__n0015[24])
  );
  X_BUF \DLX_IFinst__n0015<24>/YUSED  (
    .I(\DLX_IFinst__n0015<24>/XORG ),
    .O(DLX_IFinst__n0015[25])
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_63_2718 (
    .IA(\DLX_IFinst__n0015<24>/LOGIC_ZERO ),
    .IB(DLX_IFinst_Madd__n0005_inst_cy_62),
    .SEL(\DLX_IFinst__n0015<24>/GROM ),
    .O(\DLX_IFinst__n0015<24>/CYMUXG )
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_63 (
    .I0(DLX_IFinst_Madd__n0005_inst_cy_62),
    .I1(\DLX_IFinst__n0015<24>/GROM ),
    .O(\DLX_IFinst__n0015<24>/XORG )
  );
  X_BUF \DLX_IFinst__n0015<24>/CYINIT_2719  (
    .I(DLX_IFinst_Madd__n0005_inst_cy_61),
    .O(\DLX_IFinst__n0015<24>/CYINIT )
  );
  X_ZERO \DLX_IFinst__n0015<26>/LOGIC_ZERO_2720  (
    .O(\DLX_IFinst__n0015<26>/LOGIC_ZERO )
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_64_2721 (
    .IA(\DLX_IFinst__n0015<26>/LOGIC_ZERO ),
    .IB(\DLX_IFinst__n0015<26>/CYINIT ),
    .SEL(\DLX_IFinst__n0015<26>/FROM ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_64)
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_64 (
    .I0(\DLX_IFinst__n0015<26>/CYINIT ),
    .I1(\DLX_IFinst__n0015<26>/FROM ),
    .O(\DLX_IFinst__n0015<26>/XORF )
  );
  defparam \DLX_IFinst__n0015<26>/F .INIT = 16'hFF00;
  X_LUT4 \DLX_IFinst__n0015<26>/F  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IFinst_NPC[26]),
    .O(\DLX_IFinst__n0015<26>/FROM )
  );
  defparam \DLX_IFinst__n0015<26>/G .INIT = 16'hF0F0;
  X_LUT4 \DLX_IFinst__n0015<26>/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IFinst_NPC[27]),
    .ADR3(VCC),
    .O(\DLX_IFinst__n0015<26>/GROM )
  );
  X_BUF \DLX_IFinst__n0015<26>/COUTUSED  (
    .I(\DLX_IFinst__n0015<26>/CYMUXG ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_65)
  );
  X_BUF \DLX_IFinst__n0015<26>/XUSED  (
    .I(\DLX_IFinst__n0015<26>/XORF ),
    .O(DLX_IFinst__n0015[26])
  );
  X_BUF \DLX_IFinst__n0015<26>/YUSED  (
    .I(\DLX_IFinst__n0015<26>/XORG ),
    .O(DLX_IFinst__n0015[27])
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_65_2722 (
    .IA(\DLX_IFinst__n0015<26>/LOGIC_ZERO ),
    .IB(DLX_IFinst_Madd__n0005_inst_cy_64),
    .SEL(\DLX_IFinst__n0015<26>/GROM ),
    .O(\DLX_IFinst__n0015<26>/CYMUXG )
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_65 (
    .I0(DLX_IFinst_Madd__n0005_inst_cy_64),
    .I1(\DLX_IFinst__n0015<26>/GROM ),
    .O(\DLX_IFinst__n0015<26>/XORG )
  );
  X_BUF \DLX_IFinst__n0015<26>/CYINIT_2723  (
    .I(DLX_IFinst_Madd__n0005_inst_cy_63),
    .O(\DLX_IFinst__n0015<26>/CYINIT )
  );
  X_ZERO \DLX_IFinst__n0015<28>/LOGIC_ZERO_2724  (
    .O(\DLX_IFinst__n0015<28>/LOGIC_ZERO )
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_66_2725 (
    .IA(\DLX_IFinst__n0015<28>/LOGIC_ZERO ),
    .IB(\DLX_IFinst__n0015<28>/CYINIT ),
    .SEL(\DLX_IFinst__n0015<28>/FROM ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_66)
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_66 (
    .I0(\DLX_IFinst__n0015<28>/CYINIT ),
    .I1(\DLX_IFinst__n0015<28>/FROM ),
    .O(\DLX_IFinst__n0015<28>/XORF )
  );
  defparam \DLX_IFinst__n0015<28>/F .INIT = 16'hFF00;
  X_LUT4 \DLX_IFinst__n0015<28>/F  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IFinst_NPC[28]),
    .O(\DLX_IFinst__n0015<28>/FROM )
  );
  defparam \DLX_IFinst__n0015<28>/G .INIT = 16'hAAAA;
  X_LUT4 \DLX_IFinst__n0015<28>/G  (
    .ADR0(DLX_IFinst_NPC[29]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\DLX_IFinst__n0015<28>/GROM )
  );
  X_BUF \DLX_IFinst__n0015<28>/COUTUSED  (
    .I(\DLX_IFinst__n0015<28>/CYMUXG ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_67)
  );
  X_BUF \DLX_IFinst__n0015<28>/XUSED  (
    .I(\DLX_IFinst__n0015<28>/XORF ),
    .O(DLX_IFinst__n0015[28])
  );
  X_BUF \DLX_IFinst__n0015<28>/YUSED  (
    .I(\DLX_IFinst__n0015<28>/XORG ),
    .O(DLX_IFinst__n0015[29])
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_67_2726 (
    .IA(\DLX_IFinst__n0015<28>/LOGIC_ZERO ),
    .IB(DLX_IFinst_Madd__n0005_inst_cy_66),
    .SEL(\DLX_IFinst__n0015<28>/GROM ),
    .O(\DLX_IFinst__n0015<28>/CYMUXG )
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_67 (
    .I0(DLX_IFinst_Madd__n0005_inst_cy_66),
    .I1(\DLX_IFinst__n0015<28>/GROM ),
    .O(\DLX_IFinst__n0015<28>/XORG )
  );
  X_BUF \DLX_IFinst__n0015<28>/CYINIT_2727  (
    .I(DLX_IFinst_Madd__n0005_inst_cy_65),
    .O(\DLX_IFinst__n0015<28>/CYINIT )
  );
  X_ZERO \DLX_IFinst__n0015<30>/LOGIC_ZERO_2728  (
    .O(\DLX_IFinst__n0015<30>/LOGIC_ZERO )
  );
  X_MUX2 DLX_IFinst_Madd__n0005_inst_cy_68_2729 (
    .IA(\DLX_IFinst__n0015<30>/LOGIC_ZERO ),
    .IB(\DLX_IFinst__n0015<30>/CYINIT ),
    .SEL(\DLX_IFinst__n0015<30>/FROM ),
    .O(DLX_IFinst_Madd__n0005_inst_cy_68)
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_68 (
    .I0(\DLX_IFinst__n0015<30>/CYINIT ),
    .I1(\DLX_IFinst__n0015<30>/FROM ),
    .O(\DLX_IFinst__n0015<30>/XORF )
  );
  defparam \DLX_IFinst__n0015<30>/F .INIT = 16'hFF00;
  X_LUT4 \DLX_IFinst__n0015<30>/F  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IFinst_NPC[30]),
    .O(\DLX_IFinst__n0015<30>/FROM )
  );
  defparam \DLX_IFinst_NPC<31>_rt_2730 .INIT = 16'hFF00;
  X_LUT4 \DLX_IFinst_NPC<31>_rt_2730  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IFinst_NPC[31]),
    .O(\DLX_IFinst_NPC<31>_rt )
  );
  X_BUF \DLX_IFinst__n0015<30>/XUSED  (
    .I(\DLX_IFinst__n0015<30>/XORF ),
    .O(DLX_IFinst__n0015[30])
  );
  X_BUF \DLX_IFinst__n0015<30>/YUSED  (
    .I(\DLX_IFinst__n0015<30>/XORG ),
    .O(DLX_IFinst__n0015[31])
  );
  X_XOR2 DLX_IFinst_Madd__n0005_inst_sum_69 (
    .I0(DLX_IFinst_Madd__n0005_inst_cy_68),
    .I1(\DLX_IFinst_NPC<31>_rt ),
    .O(\DLX_IFinst__n0015<30>/XORG )
  );
  X_BUF \DLX_IFinst__n0015<30>/CYINIT_2731  (
    .I(DLX_IFinst_Madd__n0005_inst_cy_67),
    .O(\DLX_IFinst__n0015<30>/CYINIT )
  );
  X_ONE \DLX_EXinst_Mcompar__n0085_inst_cy_103/LOGIC_ONE_2732  (
    .O(\DLX_EXinst_Mcompar__n0085_inst_cy_103/LOGIC_ONE )
  );
  X_ZERO \DLX_EXinst_Mcompar__n0085_inst_cy_103/LOGIC_ZERO_2733  (
    .O(\DLX_EXinst_Mcompar__n0085_inst_cy_103/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0085_inst_cy_102_2734 (
    .IA(\DLX_EXinst_Mcompar__n0085_inst_cy_103/LOGIC_ZERO ),
    .IB(\DLX_EXinst_Mcompar__n0085_inst_cy_103/LOGIC_ONE ),
    .SEL(DLX_EXinst_Mcompar__n0085_inst_lut4_0),
    .O(DLX_EXinst_Mcompar__n0085_inst_cy_102)
  );
  defparam DLX_EXinst_Mcompar__n0085_inst_lut4_01.INIT = 16'h8241;
  X_LUT4 DLX_EXinst_Mcompar__n0085_inst_lut4_01 (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(DLX_IDinst_reg_out_B[0]),
    .ADR2(DLX_IDinst_reg_out_A[0]),
    .ADR3(DLX_IDinst_reg_out_A[1]),
    .O(DLX_EXinst_Mcompar__n0085_inst_lut4_0)
  );
  defparam DLX_EXinst_Mcompar__n0085_inst_lut4_16.INIT = 16'h9009;
  X_LUT4 DLX_EXinst_Mcompar__n0085_inst_lut4_16 (
    .ADR0(DLX_IDinst_reg_out_B_3_1),
    .ADR1(DLX_IDinst_reg_out_A[3]),
    .ADR2(DLX_IDinst_reg_out_B_2_1),
    .ADR3(DLX_IDinst_reg_out_A[2]),
    .O(DLX_EXinst_Mcompar__n0085_inst_lut4_1)
  );
  X_BUF \DLX_EXinst_Mcompar__n0085_inst_cy_103/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0085_inst_cy_103/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0085_inst_cy_103)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0085_inst_cy_103_2735 (
    .IA(\DLX_EXinst_Mcompar__n0085_inst_cy_103/LOGIC_ZERO ),
    .IB(DLX_EXinst_Mcompar__n0085_inst_cy_102),
    .SEL(DLX_EXinst_Mcompar__n0085_inst_lut4_1),
    .O(\DLX_EXinst_Mcompar__n0085_inst_cy_103/CYMUXG )
  );
  defparam DLX_IDinst_RegFile_29_28_2736.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_29_28_2736 (
    .I(DLX_IDinst_WB_data_eff[28]),
    .CE(DLX_IDinst__n0608),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_29_28)
  );
  X_ZERO \DLX_EXinst_Mcompar__n0085_inst_cy_105/LOGIC_ZERO_2737  (
    .O(\DLX_EXinst_Mcompar__n0085_inst_cy_105/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0085_inst_cy_104_2738 (
    .IA(\DLX_EXinst_Mcompar__n0085_inst_cy_105/LOGIC_ZERO ),
    .IB(\DLX_EXinst_Mcompar__n0085_inst_cy_105/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0085_inst_lut4_2),
    .O(DLX_EXinst_Mcompar__n0085_inst_cy_104)
  );
  defparam DLX_EXinst_Mcompar__n0085_inst_lut4_21.INIT = 16'h8241;
  X_LUT4 DLX_EXinst_Mcompar__n0085_inst_lut4_21 (
    .ADR0(DLX_IDinst_reg_out_B[4]),
    .ADR1(DLX_IDinst_reg_out_A[5]),
    .ADR2(DLX_IDinst_reg_out_B[5]),
    .ADR3(DLX_IDinst_reg_out_A[4]),
    .O(DLX_EXinst_Mcompar__n0085_inst_lut4_2)
  );
  defparam DLX_EXinst_Mcompar__n0085_inst_lut4_31.INIT = 16'h9009;
  X_LUT4 DLX_EXinst_Mcompar__n0085_inst_lut4_31 (
    .ADR0(DLX_IDinst_reg_out_A[6]),
    .ADR1(DLX_IDinst_reg_out_B[6]),
    .ADR2(DLX_IDinst_reg_out_B[7]),
    .ADR3(DLX_IDinst_reg_out_A[7]),
    .O(DLX_EXinst_Mcompar__n0085_inst_lut4_3)
  );
  X_BUF \DLX_EXinst_Mcompar__n0085_inst_cy_105/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0085_inst_cy_105/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0085_inst_cy_105)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0085_inst_cy_105_2739 (
    .IA(\DLX_EXinst_Mcompar__n0085_inst_cy_105/LOGIC_ZERO ),
    .IB(DLX_EXinst_Mcompar__n0085_inst_cy_104),
    .SEL(DLX_EXinst_Mcompar__n0085_inst_lut4_3),
    .O(\DLX_EXinst_Mcompar__n0085_inst_cy_105/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0085_inst_cy_105/CYINIT_2740  (
    .I(DLX_EXinst_Mcompar__n0085_inst_cy_103),
    .O(\DLX_EXinst_Mcompar__n0085_inst_cy_105/CYINIT )
  );
  X_ZERO \DLX_EXinst_Mcompar__n0085_inst_cy_107/LOGIC_ZERO_2741  (
    .O(\DLX_EXinst_Mcompar__n0085_inst_cy_107/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0085_inst_cy_106_2742 (
    .IA(\DLX_EXinst_Mcompar__n0085_inst_cy_107/LOGIC_ZERO ),
    .IB(\DLX_EXinst_Mcompar__n0085_inst_cy_107/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0085_inst_lut4_4),
    .O(DLX_EXinst_Mcompar__n0085_inst_cy_106)
  );
  defparam DLX_EXinst_Mcompar__n0085_inst_lut4_41.INIT = 16'h9009;
  X_LUT4 DLX_EXinst_Mcompar__n0085_inst_lut4_41 (
    .ADR0(DLX_IDinst_reg_out_A[9]),
    .ADR1(DLX_IDinst_reg_out_B[9]),
    .ADR2(DLX_IDinst_reg_out_A[8]),
    .ADR3(DLX_IDinst_reg_out_B[8]),
    .O(DLX_EXinst_Mcompar__n0085_inst_lut4_4)
  );
  defparam DLX_EXinst_Mcompar__n0085_inst_lut4_51.INIT = 16'h8241;
  X_LUT4 DLX_EXinst_Mcompar__n0085_inst_lut4_51 (
    .ADR0(DLX_IDinst_reg_out_B[10]),
    .ADR1(DLX_IDinst_reg_out_B[11]),
    .ADR2(DLX_IDinst_reg_out_A[11]),
    .ADR3(DLX_IDinst_reg_out_A[10]),
    .O(DLX_EXinst_Mcompar__n0085_inst_lut4_5)
  );
  X_BUF \DLX_EXinst_Mcompar__n0085_inst_cy_107/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0085_inst_cy_107/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0085_inst_cy_107)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0085_inst_cy_107_2743 (
    .IA(\DLX_EXinst_Mcompar__n0085_inst_cy_107/LOGIC_ZERO ),
    .IB(DLX_EXinst_Mcompar__n0085_inst_cy_106),
    .SEL(DLX_EXinst_Mcompar__n0085_inst_lut4_5),
    .O(\DLX_EXinst_Mcompar__n0085_inst_cy_107/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0085_inst_cy_107/CYINIT_2744  (
    .I(DLX_EXinst_Mcompar__n0085_inst_cy_105),
    .O(\DLX_EXinst_Mcompar__n0085_inst_cy_107/CYINIT )
  );
  X_ZERO \DLX_EXinst_Mcompar__n0085_inst_cy_109/LOGIC_ZERO_2745  (
    .O(\DLX_EXinst_Mcompar__n0085_inst_cy_109/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0085_inst_cy_108_2746 (
    .IA(\DLX_EXinst_Mcompar__n0085_inst_cy_109/LOGIC_ZERO ),
    .IB(\DLX_EXinst_Mcompar__n0085_inst_cy_109/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0085_inst_lut4_6),
    .O(DLX_EXinst_Mcompar__n0085_inst_cy_108)
  );
  defparam DLX_EXinst_Mcompar__n0085_inst_lut4_61.INIT = 16'h9009;
  X_LUT4 DLX_EXinst_Mcompar__n0085_inst_lut4_61 (
    .ADR0(DLX_IDinst_reg_out_B[12]),
    .ADR1(DLX_IDinst_reg_out_A[12]),
    .ADR2(DLX_IDinst_reg_out_A[13]),
    .ADR3(DLX_IDinst_reg_out_B[13]),
    .O(DLX_EXinst_Mcompar__n0085_inst_lut4_6)
  );
  defparam DLX_EXinst_Mcompar__n0085_inst_lut4_71.INIT = 16'h8241;
  X_LUT4 DLX_EXinst_Mcompar__n0085_inst_lut4_71 (
    .ADR0(DLX_IDinst_reg_out_B[15]),
    .ADR1(DLX_IDinst_reg_out_B[14]),
    .ADR2(DLX_IDinst_reg_out_A[14]),
    .ADR3(DLX_IDinst_reg_out_A[15]),
    .O(DLX_EXinst_Mcompar__n0085_inst_lut4_7)
  );
  X_BUF \DLX_EXinst_Mcompar__n0085_inst_cy_109/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0085_inst_cy_109/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0085_inst_cy_109)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0085_inst_cy_109_2747 (
    .IA(\DLX_EXinst_Mcompar__n0085_inst_cy_109/LOGIC_ZERO ),
    .IB(DLX_EXinst_Mcompar__n0085_inst_cy_108),
    .SEL(DLX_EXinst_Mcompar__n0085_inst_lut4_7),
    .O(\DLX_EXinst_Mcompar__n0085_inst_cy_109/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0085_inst_cy_109/CYINIT_2748  (
    .I(DLX_EXinst_Mcompar__n0085_inst_cy_107),
    .O(\DLX_EXinst_Mcompar__n0085_inst_cy_109/CYINIT )
  );
  X_ZERO \DLX_EXinst_Mcompar__n0085_inst_cy_111/LOGIC_ZERO_2749  (
    .O(\DLX_EXinst_Mcompar__n0085_inst_cy_111/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0085_inst_cy_110_2750 (
    .IA(\DLX_EXinst_Mcompar__n0085_inst_cy_111/LOGIC_ZERO ),
    .IB(\DLX_EXinst_Mcompar__n0085_inst_cy_111/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0085_inst_lut4_8),
    .O(DLX_EXinst_Mcompar__n0085_inst_cy_110)
  );
  defparam DLX_EXinst_Mcompar__n0085_inst_lut4_81.INIT = 16'h9009;
  X_LUT4 DLX_EXinst_Mcompar__n0085_inst_lut4_81 (
    .ADR0(DLX_IDinst_reg_out_A[17]),
    .ADR1(DLX_IDinst_reg_out_B[17]),
    .ADR2(DLX_IDinst_reg_out_B[16]),
    .ADR3(DLX_IDinst_reg_out_A[16]),
    .O(DLX_EXinst_Mcompar__n0085_inst_lut4_8)
  );
  defparam DLX_EXinst_Mcompar__n0085_inst_lut4_91.INIT = 16'h8241;
  X_LUT4 DLX_EXinst_Mcompar__n0085_inst_lut4_91 (
    .ADR0(DLX_IDinst_reg_out_B[19]),
    .ADR1(DLX_IDinst_reg_out_A[18]),
    .ADR2(DLX_IDinst_reg_out_B[18]),
    .ADR3(DLX_IDinst_reg_out_A[19]),
    .O(DLX_EXinst_Mcompar__n0085_inst_lut4_9)
  );
  X_BUF \DLX_EXinst_Mcompar__n0085_inst_cy_111/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0085_inst_cy_111/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0085_inst_cy_111)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0085_inst_cy_111_2751 (
    .IA(\DLX_EXinst_Mcompar__n0085_inst_cy_111/LOGIC_ZERO ),
    .IB(DLX_EXinst_Mcompar__n0085_inst_cy_110),
    .SEL(DLX_EXinst_Mcompar__n0085_inst_lut4_9),
    .O(\DLX_EXinst_Mcompar__n0085_inst_cy_111/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0085_inst_cy_111/CYINIT_2752  (
    .I(DLX_EXinst_Mcompar__n0085_inst_cy_109),
    .O(\DLX_EXinst_Mcompar__n0085_inst_cy_111/CYINIT )
  );
  X_ZERO \DLX_EXinst_Mcompar__n0085_inst_cy_113/LOGIC_ZERO_2753  (
    .O(\DLX_EXinst_Mcompar__n0085_inst_cy_113/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0085_inst_cy_112_2754 (
    .IA(\DLX_EXinst_Mcompar__n0085_inst_cy_113/LOGIC_ZERO ),
    .IB(\DLX_EXinst_Mcompar__n0085_inst_cy_113/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0085_inst_lut4_10),
    .O(DLX_EXinst_Mcompar__n0085_inst_cy_112)
  );
  defparam DLX_EXinst_Mcompar__n0085_inst_lut4_101.INIT = 16'h9009;
  X_LUT4 DLX_EXinst_Mcompar__n0085_inst_lut4_101 (
    .ADR0(DLX_IDinst_reg_out_A[20]),
    .ADR1(DLX_IDinst_reg_out_B[20]),
    .ADR2(DLX_IDinst_reg_out_A[21]),
    .ADR3(DLX_IDinst_reg_out_B[21]),
    .O(DLX_EXinst_Mcompar__n0085_inst_lut4_10)
  );
  defparam DLX_EXinst_Mcompar__n0085_inst_lut4_111.INIT = 16'h9009;
  X_LUT4 DLX_EXinst_Mcompar__n0085_inst_lut4_111 (
    .ADR0(DLX_IDinst_reg_out_A[22]),
    .ADR1(DLX_IDinst_reg_out_B[22]),
    .ADR2(DLX_IDinst_reg_out_B[23]),
    .ADR3(DLX_IDinst_reg_out_A[23]),
    .O(DLX_EXinst_Mcompar__n0085_inst_lut4_11)
  );
  X_BUF \DLX_EXinst_Mcompar__n0085_inst_cy_113/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0085_inst_cy_113/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0085_inst_cy_113)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0085_inst_cy_113_2755 (
    .IA(\DLX_EXinst_Mcompar__n0085_inst_cy_113/LOGIC_ZERO ),
    .IB(DLX_EXinst_Mcompar__n0085_inst_cy_112),
    .SEL(DLX_EXinst_Mcompar__n0085_inst_lut4_11),
    .O(\DLX_EXinst_Mcompar__n0085_inst_cy_113/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0085_inst_cy_113/CYINIT_2756  (
    .I(DLX_EXinst_Mcompar__n0085_inst_cy_111),
    .O(\DLX_EXinst_Mcompar__n0085_inst_cy_113/CYINIT )
  );
  X_ZERO \DLX_EXinst_Mcompar__n0085_inst_cy_115/LOGIC_ZERO_2757  (
    .O(\DLX_EXinst_Mcompar__n0085_inst_cy_115/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0085_inst_cy_114_2758 (
    .IA(\DLX_EXinst_Mcompar__n0085_inst_cy_115/LOGIC_ZERO ),
    .IB(\DLX_EXinst_Mcompar__n0085_inst_cy_115/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0085_inst_lut4_12),
    .O(DLX_EXinst_Mcompar__n0085_inst_cy_114)
  );
  defparam DLX_EXinst_Mcompar__n0085_inst_lut4_121.INIT = 16'h9009;
  X_LUT4 DLX_EXinst_Mcompar__n0085_inst_lut4_121 (
    .ADR0(DLX_IDinst_reg_out_B[24]),
    .ADR1(DLX_IDinst_reg_out_A[24]),
    .ADR2(DLX_IDinst_reg_out_B[25]),
    .ADR3(DLX_IDinst_reg_out_A[25]),
    .O(DLX_EXinst_Mcompar__n0085_inst_lut4_12)
  );
  defparam DLX_EXinst_Mcompar__n0085_inst_lut4_131.INIT = 16'h8421;
  X_LUT4 DLX_EXinst_Mcompar__n0085_inst_lut4_131 (
    .ADR0(DLX_IDinst_reg_out_B[26]),
    .ADR1(DLX_IDinst_reg_out_B[27]),
    .ADR2(DLX_IDinst_reg_out_A[26]),
    .ADR3(DLX_IDinst_reg_out_A[27]),
    .O(DLX_EXinst_Mcompar__n0085_inst_lut4_13)
  );
  X_BUF \DLX_EXinst_Mcompar__n0085_inst_cy_115/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0085_inst_cy_115/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0085_inst_cy_115)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0085_inst_cy_115_2759 (
    .IA(\DLX_EXinst_Mcompar__n0085_inst_cy_115/LOGIC_ZERO ),
    .IB(DLX_EXinst_Mcompar__n0085_inst_cy_114),
    .SEL(DLX_EXinst_Mcompar__n0085_inst_lut4_13),
    .O(\DLX_EXinst_Mcompar__n0085_inst_cy_115/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0085_inst_cy_115/CYINIT_2760  (
    .I(DLX_EXinst_Mcompar__n0085_inst_cy_113),
    .O(\DLX_EXinst_Mcompar__n0085_inst_cy_115/CYINIT )
  );
  X_ZERO \DLX_EXinst__n0085/LOGIC_ZERO_2761  (
    .O(\DLX_EXinst__n0085/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0085_inst_cy_116_2762 (
    .IA(\DLX_EXinst__n0085/LOGIC_ZERO ),
    .IB(\DLX_EXinst__n0085/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0085_inst_lut4_14),
    .O(DLX_EXinst_Mcompar__n0085_inst_cy_116)
  );
  defparam DLX_EXinst_Mcompar__n0085_inst_lut4_141.INIT = 16'h8241;
  X_LUT4 DLX_EXinst_Mcompar__n0085_inst_lut4_141 (
    .ADR0(DLX_IDinst_reg_out_B[28]),
    .ADR1(DLX_IDinst_reg_out_A[29]),
    .ADR2(DLX_IDinst_reg_out_B[29]),
    .ADR3(DLX_IDinst_reg_out_A[28]),
    .O(DLX_EXinst_Mcompar__n0085_inst_lut4_14)
  );
  defparam DLX_EXinst_Mcompar__n0085_inst_lut4_151.INIT = 16'h9009;
  X_LUT4 DLX_EXinst_Mcompar__n0085_inst_lut4_151 (
    .ADR0(DLX_IDinst_reg_out_B[30]),
    .ADR1(DLX_IDinst_reg_out_A[30]),
    .ADR2(DLX_IDinst_reg_out_B[31]),
    .ADR3(DLX_IDinst_reg_out_A[31]),
    .O(DLX_EXinst_Mcompar__n0085_inst_lut4_15)
  );
  X_BUF \DLX_EXinst__n0085/COUTUSED  (
    .I(\DLX_EXinst__n0085/CYMUXG ),
    .O(DLX_EXinst__n0085)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0085_inst_cy_117 (
    .IA(\DLX_EXinst__n0085/LOGIC_ZERO ),
    .IB(DLX_EXinst_Mcompar__n0085_inst_cy_116),
    .SEL(DLX_EXinst_Mcompar__n0085_inst_lut4_15),
    .O(\DLX_EXinst__n0085/CYMUXG )
  );
  X_BUF \DLX_EXinst__n0085/CYINIT_2763  (
    .I(DLX_EXinst_Mcompar__n0085_inst_cy_115),
    .O(\DLX_EXinst__n0085/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_1_19/LOGIC_ZERO_2764  (
    .O(\DLX_IDinst_RegFile_1_19/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_198_2765 (
    .IA(DLX_IDinst_reg_out_A[0]),
    .IB(\DLX_IDinst_RegFile_1_19/LOGIC_ZERO ),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_134),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_198)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1341.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1341 (
    .ADR0(DLX_IDinst_reg_out_A[0]),
    .ADR1(DLX_IDinst_reg_out_B[0]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_134)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1351.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1351 (
    .ADR0(DLX_IDinst_reg_out_A[1]),
    .ADR1(DLX_IDinst_reg_out_B[1]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_135)
  );
  X_BUF \DLX_IDinst_RegFile_1_19/COUTUSED  (
    .I(\DLX_IDinst_RegFile_1_19/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_199)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_199_2766 (
    .IA(DLX_IDinst_reg_out_A[1]),
    .IB(DLX_EXinst_Mcompar__n0093_inst_cy_198),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_135),
    .O(\DLX_IDinst_RegFile_1_19/CYMUXG )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_200_2767 (
    .IA(DLX_IDinst_reg_out_A[2]),
    .IB(\DLX_EXinst_Mcompar__n0093_inst_cy_201/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_136),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_200)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1361.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1361 (
    .ADR0(DLX_IDinst_reg_out_A[2]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B_2_1),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_136)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1371.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1371 (
    .ADR0(DLX_IDinst_reg_out_A[3]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B_3_1),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_137)
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_201/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0093_inst_cy_201/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_201)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_201_2768 (
    .IA(DLX_IDinst_reg_out_A[3]),
    .IB(DLX_EXinst_Mcompar__n0093_inst_cy_200),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_137),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_201/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_201/CYINIT_2769  (
    .I(DLX_EXinst_Mcompar__n0093_inst_cy_199),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_201/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_202_2770 (
    .IA(DLX_IDinst_reg_out_A[4]),
    .IB(\DLX_EXinst_Mcompar__n0093_inst_cy_203/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_138),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_202)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1381.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1381 (
    .ADR0(DLX_IDinst_reg_out_A[4]),
    .ADR1(DLX_IDinst_reg_out_B[4]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_138)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1391.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1391 (
    .ADR0(DLX_IDinst_reg_out_A[5]),
    .ADR1(DLX_IDinst_reg_out_B[5]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_139)
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_203/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0093_inst_cy_203/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_203)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_203_2771 (
    .IA(DLX_IDinst_reg_out_A[5]),
    .IB(DLX_EXinst_Mcompar__n0093_inst_cy_202),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_139),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_203/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_203/CYINIT_2772  (
    .I(DLX_EXinst_Mcompar__n0093_inst_cy_201),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_203/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_204_2773 (
    .IA(DLX_IDinst_reg_out_A[6]),
    .IB(\DLX_EXinst_Mcompar__n0093_inst_cy_205/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_140),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_204)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1401.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1401 (
    .ADR0(DLX_IDinst_reg_out_A[6]),
    .ADR1(DLX_IDinst_reg_out_B[6]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_140)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1411.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1411 (
    .ADR0(DLX_IDinst_reg_out_A[7]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[7]),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_141)
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_205/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0093_inst_cy_205/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_205)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_205_2774 (
    .IA(DLX_IDinst_reg_out_A[7]),
    .IB(DLX_EXinst_Mcompar__n0093_inst_cy_204),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_141),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_205/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_205/CYINIT_2775  (
    .I(DLX_EXinst_Mcompar__n0093_inst_cy_203),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_205/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_206_2776 (
    .IA(DLX_IDinst_reg_out_A[8]),
    .IB(\DLX_IDinst_RegFile_23_2/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_142),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_206)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1421.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1421 (
    .ADR0(DLX_IDinst_reg_out_A[8]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[8]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_142)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1431.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1431 (
    .ADR0(DLX_IDinst_reg_out_A[9]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[9]),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_143)
  );
  X_BUF \DLX_IDinst_RegFile_23_2/COUTUSED  (
    .I(\DLX_IDinst_RegFile_23_2/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_207)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_207_2777 (
    .IA(DLX_IDinst_reg_out_A[9]),
    .IB(DLX_EXinst_Mcompar__n0093_inst_cy_206),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_143),
    .O(\DLX_IDinst_RegFile_23_2/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_23_2/CYINIT_2778  (
    .I(DLX_EXinst_Mcompar__n0093_inst_cy_205),
    .O(\DLX_IDinst_RegFile_23_2/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_208_2779 (
    .IA(DLX_IDinst_reg_out_A[10]),
    .IB(\DLX_EXinst_Mcompar__n0093_inst_cy_209/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_144),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_208)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1441.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1441 (
    .ADR0(DLX_IDinst_reg_out_A[10]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[10]),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_144)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1451.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1451 (
    .ADR0(DLX_IDinst_reg_out_A[11]),
    .ADR1(DLX_IDinst_reg_out_B[11]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_145)
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_209/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0093_inst_cy_209/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_209)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_209_2780 (
    .IA(DLX_IDinst_reg_out_A[11]),
    .IB(DLX_EXinst_Mcompar__n0093_inst_cy_208),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_145),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_209/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_209/CYINIT_2781  (
    .I(DLX_EXinst_Mcompar__n0093_inst_cy_207),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_209/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_210_2782 (
    .IA(DLX_IDinst_reg_out_A[12]),
    .IB(\DLX_EXinst_Mcompar__n0093_inst_cy_211/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_146),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_210)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1461.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1461 (
    .ADR0(DLX_IDinst_reg_out_A[12]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[12]),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_146)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1471.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1471 (
    .ADR0(DLX_IDinst_reg_out_A[13]),
    .ADR1(DLX_IDinst_reg_out_B[13]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_147)
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_211/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0093_inst_cy_211/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_211)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_211_2783 (
    .IA(DLX_IDinst_reg_out_A[13]),
    .IB(DLX_EXinst_Mcompar__n0093_inst_cy_210),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_147),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_211/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_211/CYINIT_2784  (
    .I(DLX_EXinst_Mcompar__n0093_inst_cy_209),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_211/CYINIT )
  );
  defparam DLX_IDinst_RegFile_29_19_2785.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_29_19_2785 (
    .I(DLX_IDinst_WB_data_eff[19]),
    .CE(DLX_IDinst__n0608),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_29_19)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_212_2786 (
    .IA(DLX_IDinst_reg_out_A[14]),
    .IB(\DLX_EXinst_Mcompar__n0093_inst_cy_213/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_148),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_212)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1481.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1481 (
    .ADR0(DLX_IDinst_reg_out_A[14]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[14]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_148)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1491.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1491 (
    .ADR0(DLX_IDinst_reg_out_A[15]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[15]),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_149)
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_213/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0093_inst_cy_213/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_213)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_213_2787 (
    .IA(DLX_IDinst_reg_out_A[15]),
    .IB(DLX_EXinst_Mcompar__n0093_inst_cy_212),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_149),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_213/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_213/CYINIT_2788  (
    .I(DLX_EXinst_Mcompar__n0093_inst_cy_211),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_213/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_214_2789 (
    .IA(DLX_IDinst_reg_out_A[16]),
    .IB(\DLX_IDinst_RegFile_3_18/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_150),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_214)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1501.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1501 (
    .ADR0(DLX_IDinst_reg_out_A[16]),
    .ADR1(DLX_IDinst_reg_out_B[16]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_150)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1511.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1511 (
    .ADR0(DLX_IDinst_reg_out_A[17]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[17]),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_151)
  );
  X_BUF \DLX_IDinst_RegFile_3_18/COUTUSED  (
    .I(\DLX_IDinst_RegFile_3_18/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_215)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_215_2790 (
    .IA(DLX_IDinst_reg_out_A[17]),
    .IB(DLX_EXinst_Mcompar__n0093_inst_cy_214),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_151),
    .O(\DLX_IDinst_RegFile_3_18/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_3_18/CYINIT_2791  (
    .I(DLX_EXinst_Mcompar__n0093_inst_cy_213),
    .O(\DLX_IDinst_RegFile_3_18/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_216_2792 (
    .IA(DLX_IDinst_reg_out_A[18]),
    .IB(\DLX_EXinst_Mcompar__n0093_inst_cy_217/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_152),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_216)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1521.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1521 (
    .ADR0(DLX_IDinst_reg_out_A[18]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[18]),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_152)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1531.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1531 (
    .ADR0(DLX_IDinst_reg_out_A[19]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[19]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_153)
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_217/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0093_inst_cy_217/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_217)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_217_2793 (
    .IA(DLX_IDinst_reg_out_A[19]),
    .IB(DLX_EXinst_Mcompar__n0093_inst_cy_216),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_153),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_217/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_217/CYINIT_2794  (
    .I(DLX_EXinst_Mcompar__n0093_inst_cy_215),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_217/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_218_2795 (
    .IA(DLX_IDinst_reg_out_A[20]),
    .IB(\DLX_EXinst_Mcompar__n0093_inst_cy_219/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_154),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_218)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1541.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1541 (
    .ADR0(DLX_IDinst_reg_out_A[20]),
    .ADR1(DLX_IDinst_reg_out_B[20]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_154)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1551.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1551 (
    .ADR0(DLX_IDinst_reg_out_A[21]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[21]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_155)
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_219/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0093_inst_cy_219/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_219)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_219_2796 (
    .IA(DLX_IDinst_reg_out_A[21]),
    .IB(DLX_EXinst_Mcompar__n0093_inst_cy_218),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_155),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_219/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_219/CYINIT_2797  (
    .I(DLX_EXinst_Mcompar__n0093_inst_cy_217),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_219/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_220_2798 (
    .IA(DLX_IDinst_reg_out_A[22]),
    .IB(\DLX_EXinst_Mcompar__n0093_inst_cy_221/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_156),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_220)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1561.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1561 (
    .ADR0(DLX_IDinst_reg_out_A[22]),
    .ADR1(DLX_IDinst_reg_out_B[22]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_156)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1571.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1571 (
    .ADR0(DLX_IDinst_reg_out_A[23]),
    .ADR1(DLX_IDinst_reg_out_B[23]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_157)
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_221/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0093_inst_cy_221/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_221)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_221_2799 (
    .IA(DLX_IDinst_reg_out_A[23]),
    .IB(DLX_EXinst_Mcompar__n0093_inst_cy_220),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_157),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_221/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_221/CYINIT_2800  (
    .I(DLX_EXinst_Mcompar__n0093_inst_cy_219),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_221/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_222_2801 (
    .IA(DLX_IDinst_reg_out_A[24]),
    .IB(\DLX_IFinst_IR_curr<6>/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_158),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_222)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1581.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1581 (
    .ADR0(DLX_IDinst_reg_out_A[24]),
    .ADR1(DLX_IDinst_reg_out_B[24]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_158)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1591.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1591 (
    .ADR0(DLX_IDinst_reg_out_A[25]),
    .ADR1(DLX_IDinst_reg_out_B[25]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_159)
  );
  X_BUF \DLX_IFinst_IR_curr<6>/COUTUSED  (
    .I(\DLX_IFinst_IR_curr<6>/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_223)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_223_2802 (
    .IA(DLX_IDinst_reg_out_A[25]),
    .IB(DLX_EXinst_Mcompar__n0093_inst_cy_222),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_159),
    .O(\DLX_IFinst_IR_curr<6>/CYMUXG )
  );
  X_BUF \DLX_IFinst_IR_curr<6>/CYINIT_2803  (
    .I(DLX_EXinst_Mcompar__n0093_inst_cy_221),
    .O(\DLX_IFinst_IR_curr<6>/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_224_2804 (
    .IA(DLX_IDinst_reg_out_A[26]),
    .IB(\DLX_EXinst_Mcompar__n0093_inst_cy_225/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_160),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_224)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1601.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1601 (
    .ADR0(DLX_IDinst_reg_out_A[26]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[26]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_160)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1611.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1611 (
    .ADR0(DLX_IDinst_reg_out_A[27]),
    .ADR1(DLX_IDinst_reg_out_B[27]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_161)
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_225/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0093_inst_cy_225/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_225)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_225_2805 (
    .IA(DLX_IDinst_reg_out_A[27]),
    .IB(DLX_EXinst_Mcompar__n0093_inst_cy_224),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_161),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_225/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_225/CYINIT_2806  (
    .I(DLX_EXinst_Mcompar__n0093_inst_cy_223),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_225/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_226_2807 (
    .IA(DLX_IDinst_reg_out_A[28]),
    .IB(\DLX_EXinst_Mcompar__n0093_inst_cy_227/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_162),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_226)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1621.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1621 (
    .ADR0(DLX_IDinst_reg_out_A[28]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[28]),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_162)
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1631.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1631 (
    .ADR0(DLX_IDinst_reg_out_A[29]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[29]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_163)
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_227/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0093_inst_cy_227/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_227)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_227_2808 (
    .IA(DLX_IDinst_reg_out_A[29]),
    .IB(DLX_EXinst_Mcompar__n0093_inst_cy_226),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_163),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_227/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_227/CYINIT_2809  (
    .I(DLX_EXinst_Mcompar__n0093_inst_cy_225),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_227/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0093_inst_cy_228_2810 (
    .IA(DLX_IDinst_reg_out_A[30]),
    .IB(\DLX_EXinst_Mcompar__n0093_inst_cy_228/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0093_inst_lut2_164),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_228/CYMUXF )
  );
  defparam DLX_EXinst_Mcompar__n0093_inst_lut2_1641.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0093_inst_lut2_1641 (
    .ADR0(DLX_IDinst_reg_out_A[30]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[30]),
    .O(DLX_EXinst_Mcompar__n0093_inst_lut2_164)
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_228/XBUSED  (
    .I(\DLX_EXinst_Mcompar__n0093_inst_cy_228/CYMUXF ),
    .O(DLX_EXinst_Mcompar__n0093_inst_cy_228)
  );
  X_BUF \DLX_EXinst_Mcompar__n0093_inst_cy_228/CYINIT_2811  (
    .I(DLX_EXinst_Mcompar__n0093_inst_cy_227),
    .O(\DLX_EXinst_Mcompar__n0093_inst_cy_228/CYINIT )
  );
  X_ZERO \DLX_EXinst_Mcompar__n0069_inst_cy_231/LOGIC_ZERO_2812  (
    .O(\DLX_EXinst_Mcompar__n0069_inst_cy_231/LOGIC_ZERO )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0069_inst_cy_230_2813 (
    .IA(DLX_IDinst_Imm_0_1),
    .IB(\DLX_EXinst_Mcompar__n0069_inst_cy_231/LOGIC_ZERO ),
    .SEL(DLX_EXinst_Mcompar__n0069_inst_lut2_166),
    .O(DLX_EXinst_Mcompar__n0069_inst_cy_230)
  );
  defparam DLX_EXinst_Mcompar__n0069_inst_lut2_1661.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0069_inst_lut2_1661 (
    .ADR0(DLX_IDinst_Imm_0_1),
    .ADR1(DLX_IDinst_reg_out_A[0]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0069_inst_lut2_166)
  );
  defparam DLX_EXinst_Mcompar__n0069_inst_lut2_1671.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0069_inst_lut2_1671 (
    .ADR0(DLX_IDinst_Imm_1_1),
    .ADR1(DLX_IDinst_reg_out_A[1]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0069_inst_lut2_167)
  );
  X_BUF \DLX_EXinst_Mcompar__n0069_inst_cy_231/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0069_inst_cy_231/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0069_inst_cy_231)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0069_inst_cy_231_2814 (
    .IA(DLX_IDinst_Imm_1_1),
    .IB(DLX_EXinst_Mcompar__n0069_inst_cy_230),
    .SEL(DLX_EXinst_Mcompar__n0069_inst_lut2_167),
    .O(\DLX_EXinst_Mcompar__n0069_inst_cy_231/CYMUXG )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0069_inst_cy_232_2815 (
    .IA(DLX_IDinst_Imm_2_1),
    .IB(\DLX_IDinst_RegFile_2_26/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0069_inst_lut2_168),
    .O(DLX_EXinst_Mcompar__n0069_inst_cy_232)
  );
  defparam DLX_EXinst_Mcompar__n0069_inst_lut2_1681.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0069_inst_lut2_1681 (
    .ADR0(DLX_IDinst_Imm_2_1),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[2]),
    .O(DLX_EXinst_Mcompar__n0069_inst_lut2_168)
  );
  defparam DLX_EXinst_Mcompar__n0069_inst_lut2_1691.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0069_inst_lut2_1691 (
    .ADR0(DLX_IDinst_Imm_3_1),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[3]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0069_inst_lut2_169)
  );
  X_BUF \DLX_IDinst_RegFile_2_26/COUTUSED  (
    .I(\DLX_IDinst_RegFile_2_26/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0069_inst_cy_233)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0069_inst_cy_233_2816 (
    .IA(DLX_IDinst_Imm_3_1),
    .IB(DLX_EXinst_Mcompar__n0069_inst_cy_232),
    .SEL(DLX_EXinst_Mcompar__n0069_inst_lut2_169),
    .O(\DLX_IDinst_RegFile_2_26/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_2_26/CYINIT_2817  (
    .I(DLX_EXinst_Mcompar__n0069_inst_cy_231),
    .O(\DLX_IDinst_RegFile_2_26/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0069_inst_cy_234_2818 (
    .IA(\DLX_IDinst_Imm[4] ),
    .IB(\DLX_EXinst_Mcompar__n0069_inst_cy_235/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0069_inst_lut2_170),
    .O(DLX_EXinst_Mcompar__n0069_inst_cy_234)
  );
  defparam DLX_EXinst_Mcompar__n0069_inst_lut2_1701.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0069_inst_lut2_1701 (
    .ADR0(\DLX_IDinst_Imm[4] ),
    .ADR1(DLX_IDinst_reg_out_A[4]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0069_inst_lut2_170)
  );
  defparam DLX_EXinst_Mcompar__n0069_inst_lut2_1711.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0069_inst_lut2_1711 (
    .ADR0(\DLX_IDinst_Imm[5] ),
    .ADR1(DLX_IDinst_reg_out_A[5]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0069_inst_lut2_171)
  );
  X_BUF \DLX_EXinst_Mcompar__n0069_inst_cy_235/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0069_inst_cy_235/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0069_inst_cy_235)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0069_inst_cy_235_2819 (
    .IA(\DLX_IDinst_Imm[5] ),
    .IB(DLX_EXinst_Mcompar__n0069_inst_cy_234),
    .SEL(DLX_EXinst_Mcompar__n0069_inst_lut2_171),
    .O(\DLX_EXinst_Mcompar__n0069_inst_cy_235/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0069_inst_cy_235/CYINIT_2820  (
    .I(DLX_EXinst_Mcompar__n0069_inst_cy_233),
    .O(\DLX_EXinst_Mcompar__n0069_inst_cy_235/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0069_inst_cy_236_2821 (
    .IA(\DLX_IDinst_Imm[6] ),
    .IB(\DLX_EXinst_Mcompar__n0069_inst_cy_237/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0069_inst_lut2_172),
    .O(DLX_EXinst_Mcompar__n0069_inst_cy_236)
  );
  defparam DLX_EXinst_Mcompar__n0069_inst_lut2_1721.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0069_inst_lut2_1721 (
    .ADR0(\DLX_IDinst_Imm[6] ),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[6]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0069_inst_lut2_172)
  );
  defparam DLX_EXinst_Mcompar__n0069_inst_lut2_1731.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0069_inst_lut2_1731 (
    .ADR0(\DLX_IDinst_Imm[7] ),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[7]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0069_inst_lut2_173)
  );
  X_BUF \DLX_EXinst_Mcompar__n0069_inst_cy_237/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0069_inst_cy_237/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0069_inst_cy_237)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0069_inst_cy_237_2822 (
    .IA(\DLX_IDinst_Imm[7] ),
    .IB(DLX_EXinst_Mcompar__n0069_inst_cy_236),
    .SEL(DLX_EXinst_Mcompar__n0069_inst_lut2_173),
    .O(\DLX_EXinst_Mcompar__n0069_inst_cy_237/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0069_inst_cy_237/CYINIT_2823  (
    .I(DLX_EXinst_Mcompar__n0069_inst_cy_235),
    .O(\DLX_EXinst_Mcompar__n0069_inst_cy_237/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0069_inst_cy_238_2824 (
    .IA(\DLX_IDinst_Imm[8] ),
    .IB(\DLX_EXinst_Mcompar__n0069_inst_cy_239/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0069_inst_lut2_174),
    .O(DLX_EXinst_Mcompar__n0069_inst_cy_238)
  );
  defparam DLX_EXinst_Mcompar__n0069_inst_lut2_1741.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0069_inst_lut2_1741 (
    .ADR0(\DLX_IDinst_Imm[8] ),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[8]),
    .O(DLX_EXinst_Mcompar__n0069_inst_lut2_174)
  );
  defparam DLX_EXinst_Mcompar__n0069_inst_lut2_1751.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0069_inst_lut2_1751 (
    .ADR0(\DLX_IDinst_Imm[9] ),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[9]),
    .O(DLX_EXinst_Mcompar__n0069_inst_lut2_175)
  );
  X_BUF \DLX_EXinst_Mcompar__n0069_inst_cy_239/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0069_inst_cy_239/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0069_inst_cy_239)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0069_inst_cy_239_2825 (
    .IA(\DLX_IDinst_Imm[9] ),
    .IB(DLX_EXinst_Mcompar__n0069_inst_cy_238),
    .SEL(DLX_EXinst_Mcompar__n0069_inst_lut2_175),
    .O(\DLX_EXinst_Mcompar__n0069_inst_cy_239/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0069_inst_cy_239/CYINIT_2826  (
    .I(DLX_EXinst_Mcompar__n0069_inst_cy_237),
    .O(\DLX_EXinst_Mcompar__n0069_inst_cy_239/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0069_inst_cy_240_2827 (
    .IA(\DLX_IDinst_Imm[10] ),
    .IB(\DLX_IFinst_IR_curr<27>/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0069_inst_lut2_176),
    .O(DLX_EXinst_Mcompar__n0069_inst_cy_240)
  );
  defparam DLX_EXinst_Mcompar__n0069_inst_lut2_1761.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0069_inst_lut2_1761 (
    .ADR0(\DLX_IDinst_Imm[10] ),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[10]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0069_inst_lut2_176)
  );
  defparam DLX_EXinst_Mcompar__n0069_inst_lut2_1771.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0069_inst_lut2_1771 (
    .ADR0(\DLX_IDinst_Imm[11] ),
    .ADR1(DLX_IDinst_reg_out_A[11]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0069_inst_lut2_177)
  );
  X_BUF \DLX_IFinst_IR_curr<27>/COUTUSED  (
    .I(\DLX_IFinst_IR_curr<27>/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0069_inst_cy_241)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0069_inst_cy_241_2828 (
    .IA(\DLX_IDinst_Imm[11] ),
    .IB(DLX_EXinst_Mcompar__n0069_inst_cy_240),
    .SEL(DLX_EXinst_Mcompar__n0069_inst_lut2_177),
    .O(\DLX_IFinst_IR_curr<27>/CYMUXG )
  );
  X_BUF \DLX_IFinst_IR_curr<27>/CYINIT_2829  (
    .I(DLX_EXinst_Mcompar__n0069_inst_cy_239),
    .O(\DLX_IFinst_IR_curr<27>/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0069_inst_cy_242_2830 (
    .IA(\DLX_IDinst_Imm[12] ),
    .IB(\DLX_EXinst_Mcompar__n0069_inst_cy_243/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0069_inst_lut2_178),
    .O(DLX_EXinst_Mcompar__n0069_inst_cy_242)
  );
  defparam DLX_EXinst_Mcompar__n0069_inst_lut2_1781.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0069_inst_lut2_1781 (
    .ADR0(\DLX_IDinst_Imm[12] ),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[12]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0069_inst_lut2_178)
  );
  defparam DLX_EXinst_Mcompar__n0069_inst_lut2_1791.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0069_inst_lut2_1791 (
    .ADR0(\DLX_IDinst_Imm[13] ),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[13]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0069_inst_lut2_179)
  );
  X_BUF \DLX_EXinst_Mcompar__n0069_inst_cy_243/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0069_inst_cy_243/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0069_inst_cy_243)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0069_inst_cy_243_2831 (
    .IA(\DLX_IDinst_Imm[13] ),
    .IB(DLX_EXinst_Mcompar__n0069_inst_cy_242),
    .SEL(DLX_EXinst_Mcompar__n0069_inst_lut2_179),
    .O(\DLX_EXinst_Mcompar__n0069_inst_cy_243/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0069_inst_cy_243/CYINIT_2832  (
    .I(DLX_EXinst_Mcompar__n0069_inst_cy_241),
    .O(\DLX_EXinst_Mcompar__n0069_inst_cy_243/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0069_inst_cy_244_2833 (
    .IA(\DLX_IDinst_Imm[14] ),
    .IB(\DLX_EXinst_Mcompar__n0069_inst_cy_245/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0069_inst_lut2_180),
    .O(DLX_EXinst_Mcompar__n0069_inst_cy_244)
  );
  defparam DLX_EXinst_Mcompar__n0069_inst_lut2_1801.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0069_inst_lut2_1801 (
    .ADR0(\DLX_IDinst_Imm[14] ),
    .ADR1(DLX_IDinst_reg_out_A[14]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0069_inst_lut2_180)
  );
  defparam DLX_EXinst_Mcompar__n0069_inst_lut2_1811.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0069_inst_lut2_1811 (
    .ADR0(\DLX_IDinst_Imm[15] ),
    .ADR1(DLX_IDinst_reg_out_A[15]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0069_inst_lut2_181)
  );
  X_BUF \DLX_EXinst_Mcompar__n0069_inst_cy_245/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0069_inst_cy_245/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0069_inst_cy_245)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0069_inst_cy_245_2834 (
    .IA(\DLX_IDinst_Imm[15] ),
    .IB(DLX_EXinst_Mcompar__n0069_inst_cy_244),
    .SEL(DLX_EXinst_Mcompar__n0069_inst_lut2_181),
    .O(\DLX_EXinst_Mcompar__n0069_inst_cy_245/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0069_inst_cy_245/CYINIT_2835  (
    .I(DLX_EXinst_Mcompar__n0069_inst_cy_243),
    .O(\DLX_EXinst_Mcompar__n0069_inst_cy_245/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0069_inst_cy_246_2836 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(\DLX_EXinst_Mcompar__n0069_inst_cy_247/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0069_inst_lut2_182),
    .O(DLX_EXinst_Mcompar__n0069_inst_cy_246)
  );
  defparam DLX_EXinst_Mcompar__n0069_inst_lut2_1821.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0069_inst_lut2_1821 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[16]),
    .O(DLX_EXinst_Mcompar__n0069_inst_lut2_182)
  );
  defparam DLX_EXinst_Mcompar__n0069_inst_lut2_1831.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0069_inst_lut2_1831 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[17]),
    .O(DLX_EXinst_Mcompar__n0069_inst_lut2_183)
  );
  X_BUF \DLX_EXinst_Mcompar__n0069_inst_cy_247/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0069_inst_cy_247/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0069_inst_cy_247)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0069_inst_cy_247_2837 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(DLX_EXinst_Mcompar__n0069_inst_cy_246),
    .SEL(DLX_EXinst_Mcompar__n0069_inst_lut2_183),
    .O(\DLX_EXinst_Mcompar__n0069_inst_cy_247/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0069_inst_cy_247/CYINIT_2838  (
    .I(DLX_EXinst_Mcompar__n0069_inst_cy_245),
    .O(\DLX_EXinst_Mcompar__n0069_inst_cy_247/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0069_inst_cy_248_2839 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(\DLX_IDinst_RegFile_3_26/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0069_inst_lut2_184),
    .O(DLX_EXinst_Mcompar__n0069_inst_cy_248)
  );
  defparam DLX_EXinst_Mcompar__n0069_inst_lut2_1841.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0069_inst_lut2_1841 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[18]),
    .O(DLX_EXinst_Mcompar__n0069_inst_lut2_184)
  );
  defparam DLX_EXinst_Mcompar__n0069_inst_lut2_1851.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0069_inst_lut2_1851 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[19]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0069_inst_lut2_185)
  );
  X_BUF \DLX_IDinst_RegFile_3_26/COUTUSED  (
    .I(\DLX_IDinst_RegFile_3_26/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0069_inst_cy_249)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0069_inst_cy_249_2840 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(DLX_EXinst_Mcompar__n0069_inst_cy_248),
    .SEL(DLX_EXinst_Mcompar__n0069_inst_lut2_185),
    .O(\DLX_IDinst_RegFile_3_26/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_3_26/CYINIT_2841  (
    .I(DLX_EXinst_Mcompar__n0069_inst_cy_247),
    .O(\DLX_IDinst_RegFile_3_26/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0069_inst_cy_250_2842 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(\DLX_EXinst_Mcompar__n0069_inst_cy_251/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0069_inst_lut2_186),
    .O(DLX_EXinst_Mcompar__n0069_inst_cy_250)
  );
  defparam DLX_EXinst_Mcompar__n0069_inst_lut2_1861.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0069_inst_lut2_1861 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(DLX_IDinst_reg_out_A[20]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0069_inst_lut2_186)
  );
  defparam DLX_EXinst_Mcompar__n0069_inst_lut2_1871.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0069_inst_lut2_1871 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[21]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0069_inst_lut2_187)
  );
  X_BUF \DLX_EXinst_Mcompar__n0069_inst_cy_251/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0069_inst_cy_251/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0069_inst_cy_251)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0069_inst_cy_251_2843 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(DLX_EXinst_Mcompar__n0069_inst_cy_250),
    .SEL(DLX_EXinst_Mcompar__n0069_inst_lut2_187),
    .O(\DLX_EXinst_Mcompar__n0069_inst_cy_251/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0069_inst_cy_251/CYINIT_2844  (
    .I(DLX_EXinst_Mcompar__n0069_inst_cy_249),
    .O(\DLX_EXinst_Mcompar__n0069_inst_cy_251/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0069_inst_cy_252_2845 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(\DLX_EXinst_Mcompar__n0069_inst_cy_253/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0069_inst_lut2_188),
    .O(DLX_EXinst_Mcompar__n0069_inst_cy_252)
  );
  defparam DLX_EXinst_Mcompar__n0069_inst_lut2_1881.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0069_inst_lut2_1881 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(DLX_IDinst_reg_out_A[22]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0069_inst_lut2_188)
  );
  defparam DLX_EXinst_Mcompar__n0069_inst_lut2_1891.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0069_inst_lut2_1891 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[23]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0069_inst_lut2_189)
  );
  X_BUF \DLX_EXinst_Mcompar__n0069_inst_cy_253/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0069_inst_cy_253/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0069_inst_cy_253)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0069_inst_cy_253_2846 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(DLX_EXinst_Mcompar__n0069_inst_cy_252),
    .SEL(DLX_EXinst_Mcompar__n0069_inst_lut2_189),
    .O(\DLX_EXinst_Mcompar__n0069_inst_cy_253/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0069_inst_cy_253/CYINIT_2847  (
    .I(DLX_EXinst_Mcompar__n0069_inst_cy_251),
    .O(\DLX_EXinst_Mcompar__n0069_inst_cy_253/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0069_inst_cy_254_2848 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(\DLX_EXinst_Mcompar__n0069_inst_cy_255/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0069_inst_lut2_190),
    .O(DLX_EXinst_Mcompar__n0069_inst_cy_254)
  );
  defparam DLX_EXinst_Mcompar__n0069_inst_lut2_1901.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0069_inst_lut2_1901 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[24]),
    .O(DLX_EXinst_Mcompar__n0069_inst_lut2_190)
  );
  defparam DLX_EXinst_Mcompar__n0069_inst_lut2_1911.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0069_inst_lut2_1911 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[25]),
    .O(DLX_EXinst_Mcompar__n0069_inst_lut2_191)
  );
  X_BUF \DLX_EXinst_Mcompar__n0069_inst_cy_255/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0069_inst_cy_255/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0069_inst_cy_255)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0069_inst_cy_255_2849 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(DLX_EXinst_Mcompar__n0069_inst_cy_254),
    .SEL(DLX_EXinst_Mcompar__n0069_inst_lut2_191),
    .O(\DLX_EXinst_Mcompar__n0069_inst_cy_255/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0069_inst_cy_255/CYINIT_2850  (
    .I(DLX_EXinst_Mcompar__n0069_inst_cy_253),
    .O(\DLX_EXinst_Mcompar__n0069_inst_cy_255/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0069_inst_cy_256_2851 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(\DLX_IFinst_IR_curr<19>/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0069_inst_lut2_192),
    .O(DLX_EXinst_Mcompar__n0069_inst_cy_256)
  );
  defparam DLX_EXinst_Mcompar__n0069_inst_lut2_1921.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0069_inst_lut2_1921 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[26]),
    .O(DLX_EXinst_Mcompar__n0069_inst_lut2_192)
  );
  defparam DLX_EXinst_Mcompar__n0069_inst_lut2_1931.INIT = 16'hAA55;
  X_LUT4 DLX_EXinst_Mcompar__n0069_inst_lut2_1931 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_A[27]),
    .O(DLX_EXinst_Mcompar__n0069_inst_lut2_193)
  );
  X_BUF \DLX_IFinst_IR_curr<19>/COUTUSED  (
    .I(\DLX_IFinst_IR_curr<19>/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0069_inst_cy_257)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0069_inst_cy_257_2852 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(DLX_EXinst_Mcompar__n0069_inst_cy_256),
    .SEL(DLX_EXinst_Mcompar__n0069_inst_lut2_193),
    .O(\DLX_IFinst_IR_curr<19>/CYMUXG )
  );
  X_BUF \DLX_IFinst_IR_curr<19>/CYINIT_2853  (
    .I(DLX_EXinst_Mcompar__n0069_inst_cy_255),
    .O(\DLX_IFinst_IR_curr<19>/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0069_inst_cy_258_2854 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(\DLX_EXinst_Mcompar__n0069_inst_cy_259/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0069_inst_lut2_194),
    .O(DLX_EXinst_Mcompar__n0069_inst_cy_258)
  );
  defparam DLX_EXinst_Mcompar__n0069_inst_lut2_1941.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0069_inst_lut2_1941 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(DLX_IDinst_reg_out_A[28]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0069_inst_lut2_194)
  );
  defparam DLX_EXinst_Mcompar__n0069_inst_lut2_1951.INIT = 16'h9999;
  X_LUT4 DLX_EXinst_Mcompar__n0069_inst_lut2_1951 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(DLX_IDinst_reg_out_A[29]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0069_inst_lut2_195)
  );
  X_BUF \DLX_EXinst_Mcompar__n0069_inst_cy_259/COUTUSED  (
    .I(\DLX_EXinst_Mcompar__n0069_inst_cy_259/CYMUXG ),
    .O(DLX_EXinst_Mcompar__n0069_inst_cy_259)
  );
  X_MUX2 DLX_EXinst_Mcompar__n0069_inst_cy_259_2855 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(DLX_EXinst_Mcompar__n0069_inst_cy_258),
    .SEL(DLX_EXinst_Mcompar__n0069_inst_lut2_195),
    .O(\DLX_EXinst_Mcompar__n0069_inst_cy_259/CYMUXG )
  );
  X_BUF \DLX_EXinst_Mcompar__n0069_inst_cy_259/CYINIT_2856  (
    .I(DLX_EXinst_Mcompar__n0069_inst_cy_257),
    .O(\DLX_EXinst_Mcompar__n0069_inst_cy_259/CYINIT )
  );
  X_MUX2 DLX_EXinst_Mcompar__n0069_inst_cy_260_2857 (
    .IA(DLX_IDinst_Imm_31_1),
    .IB(\DLX_EXinst_Mcompar__n0069_inst_cy_260/CYINIT ),
    .SEL(DLX_EXinst_Mcompar__n0069_inst_lut2_196),
    .O(\DLX_EXinst_Mcompar__n0069_inst_cy_260/CYMUXF )
  );
  defparam DLX_EXinst_Mcompar__n0069_inst_lut2_1961.INIT = 16'hA5A5;
  X_LUT4 DLX_EXinst_Mcompar__n0069_inst_lut2_1961 (
    .ADR0(DLX_IDinst_Imm_31_1),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_A[30]),
    .ADR3(VCC),
    .O(DLX_EXinst_Mcompar__n0069_inst_lut2_196)
  );
  X_BUF \DLX_EXinst_Mcompar__n0069_inst_cy_260/XBUSED  (
    .I(\DLX_EXinst_Mcompar__n0069_inst_cy_260/CYMUXF ),
    .O(DLX_EXinst_Mcompar__n0069_inst_cy_260)
  );
  X_BUF \DLX_EXinst_Mcompar__n0069_inst_cy_260/CYINIT_2858  (
    .I(DLX_EXinst_Mcompar__n0069_inst_cy_259),
    .O(\DLX_EXinst_Mcompar__n0069_inst_cy_260/CYINIT )
  );
  X_ONE \DLX_IDinst_Mcompar__n0100_inst_cy_263/LOGIC_ONE_2859  (
    .O(\DLX_IDinst_Mcompar__n0100_inst_cy_263/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mcompar__n0100_inst_cy_263/LOGIC_ZERO_2860  (
    .O(\DLX_IDinst_Mcompar__n0100_inst_cy_263/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mcompar__n0100_inst_cy_262_2861 (
    .IA(\DLX_IDinst_Mcompar__n0100_inst_cy_263/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mcompar__n0100_inst_cy_263/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mcompar__n0100_inst_lut4_40),
    .O(DLX_IDinst_Mcompar__n0100_inst_cy_262)
  );
  defparam DLX_IDinst_Mcompar__n0100_inst_lut4_401.INIT = 16'h8241;
  X_LUT4 DLX_IDinst_Mcompar__n0100_inst_lut4_401 (
    .ADR0(DLX_IDinst_jtarget[22]),
    .ADR1(DLX_reg_dst_of_EX[0]),
    .ADR2(DLX_IDinst_jtarget[21]),
    .ADR3(DLX_reg_dst_of_EX[1]),
    .O(DLX_IDinst_Mcompar__n0100_inst_lut4_40)
  );
  defparam DLX_IDinst_Mcompar__n0100_inst_lut4_411.INIT = 16'h8241;
  X_LUT4 DLX_IDinst_Mcompar__n0100_inst_lut4_411 (
    .ADR0(DLX_reg_dst_of_EX[2]),
    .ADR1(DLX_reg_dst_of_EX[3]),
    .ADR2(DLX_IDinst_jtarget[24]),
    .ADR3(DLX_IDinst_jtarget[23]),
    .O(DLX_IDinst_Mcompar__n0100_inst_lut4_41)
  );
  X_BUF \DLX_IDinst_Mcompar__n0100_inst_cy_263/COUTUSED  (
    .I(\DLX_IDinst_Mcompar__n0100_inst_cy_263/CYMUXG ),
    .O(DLX_IDinst_Mcompar__n0100_inst_cy_263)
  );
  X_MUX2 DLX_IDinst_Mcompar__n0100_inst_cy_263_2862 (
    .IA(\DLX_IDinst_Mcompar__n0100_inst_cy_263/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mcompar__n0100_inst_cy_262),
    .SEL(DLX_IDinst_Mcompar__n0100_inst_lut4_41),
    .O(\DLX_IDinst_Mcompar__n0100_inst_cy_263/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mmux__COND_5_inst_cy_1009/LOGIC_ONE_2863  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_1009/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mmux__COND_5_inst_cy_1009/LOGIC_ZERO_2864  (
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_1009/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_1008_2865 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_1009/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mmux__COND_5_inst_cy_1009/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1083),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_1008)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10831.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10831 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR1(DLX_IDinst_RegFile_0_31),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_571),
    .ADR3(DLX_IDinst_RegFile_1_31),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1083)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10841.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10841 (
    .ADR0(DLX_IDinst_RegFile_2_31),
    .ADR1(DLX_IDinst_RegFile_3_31),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_572),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1084)
  );
  X_BUF \DLX_IDinst_Mmux__COND_5_inst_cy_1009/COUTUSED  (
    .I(\DLX_IDinst_Mmux__COND_5_inst_cy_1009/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_1009)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_1009_2866 (
    .IA(\DLX_IDinst_Mmux__COND_5_inst_cy_1009/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_1008),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1084),
    .O(\DLX_IDinst_Mmux__COND_5_inst_cy_1009/CYMUXG )
  );
  X_ONE \DLX_IDinst_Mcompar__n0105_inst_cy_263/LOGIC_ONE_2867  (
    .O(\DLX_IDinst_Mcompar__n0105_inst_cy_263/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mcompar__n0105_inst_cy_263/LOGIC_ZERO_2868  (
    .O(\DLX_IDinst_Mcompar__n0105_inst_cy_263/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mcompar__n0105_inst_cy_262_2869 (
    .IA(\DLX_IDinst_Mcompar__n0105_inst_cy_263/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mcompar__n0105_inst_cy_263/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mcompar__n0105_inst_lut4_40),
    .O(DLX_IDinst_Mcompar__n0105_inst_cy_262)
  );
  defparam DLX_IDinst_Mcompar__n0105_inst_lut4_401.INIT = 16'h8241;
  X_LUT4 DLX_IDinst_Mcompar__n0105_inst_lut4_401 (
    .ADR0(DLX_IDinst_jtarget[16]),
    .ADR1(DLX_EXinst_reg_dst_out[1]),
    .ADR2(DLX_IDinst_jtarget[17]),
    .ADR3(DLX_EXinst_reg_dst_out[0]),
    .O(DLX_IDinst_Mcompar__n0105_inst_lut4_40)
  );
  defparam DLX_IDinst_Mcompar__n0105_inst_lut4_411.INIT = 16'h8421;
  X_LUT4 DLX_IDinst_Mcompar__n0105_inst_lut4_411 (
    .ADR0(DLX_IDinst_jtarget[18]),
    .ADR1(DLX_IDinst_jtarget[19]),
    .ADR2(DLX_EXinst_reg_dst_out[2]),
    .ADR3(DLX_EXinst_reg_dst_out[3]),
    .O(DLX_IDinst_Mcompar__n0105_inst_lut4_41)
  );
  X_BUF \DLX_IDinst_Mcompar__n0105_inst_cy_263/COUTUSED  (
    .I(\DLX_IDinst_Mcompar__n0105_inst_cy_263/CYMUXG ),
    .O(DLX_IDinst_Mcompar__n0105_inst_cy_263)
  );
  X_MUX2 DLX_IDinst_Mcompar__n0105_inst_cy_263_2870 (
    .IA(\DLX_IDinst_Mcompar__n0105_inst_cy_263/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mcompar__n0105_inst_cy_262),
    .SEL(DLX_IDinst_Mcompar__n0105_inst_lut4_41),
    .O(\DLX_IDinst_Mcompar__n0105_inst_cy_263/CYMUXG )
  );
  X_ZERO \DLX_IDinst__n0105/LOGIC_ZERO_2871  (
    .O(\DLX_IDinst__n0105/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mcompar__n0105_inst_cy_264 (
    .IA(\DLX_IDinst__n0105/LOGIC_ZERO ),
    .IB(\DLX_IDinst__n0105/CYINIT ),
    .SEL(DLX_IDinst_Mcompar__n0105_inst_lut4_42),
    .O(\DLX_IDinst__n0105/CYMUXF )
  );
  defparam DLX_IDinst_Mcompar__n0105_inst_lut4_421.INIT = 16'h9A95;
  X_LUT4 DLX_IDinst_Mcompar__n0105_inst_lut4_421 (
    .ADR0(DLX_EXinst_reg_dst_out[4]),
    .ADR1(DLX_IFinst_IR_latched[20]),
    .ADR2(DLX_EXinst__n0144),
    .ADR3(DLX_IDinst_current_IR[20]),
    .O(DLX_IDinst_Mcompar__n0105_inst_lut4_42)
  );
  X_BUF \DLX_IDinst__n0105/XBUSED  (
    .I(\DLX_IDinst__n0105/CYMUXF ),
    .O(DLX_IDinst__n0105)
  );
  X_BUF \DLX_IDinst__n0105/CYINIT_2872  (
    .I(DLX_IDinst_Mcompar__n0105_inst_cy_263),
    .O(\DLX_IDinst__n0105/CYINIT )
  );
  X_ONE \DLX_IDinst_Mcompar__n0367_inst_cy_263/LOGIC_ONE_2873  (
    .O(\DLX_IDinst_Mcompar__n0367_inst_cy_263/LOGIC_ONE )
  );
  X_ZERO \DLX_IDinst_Mcompar__n0367_inst_cy_263/LOGIC_ZERO_2874  (
    .O(\DLX_IDinst_Mcompar__n0367_inst_cy_263/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mcompar__n0367_inst_cy_262_2875 (
    .IA(\DLX_IDinst_Mcompar__n0367_inst_cy_263/LOGIC_ZERO ),
    .IB(\DLX_IDinst_Mcompar__n0367_inst_cy_263/LOGIC_ONE ),
    .SEL(DLX_IDinst_Mcompar__n0367_inst_lut4_40),
    .O(DLX_IDinst_Mcompar__n0367_inst_cy_262)
  );
  defparam DLX_IDinst_Mcompar__n0367_inst_lut4_401.INIT = 16'h8421;
  X_LUT4 DLX_IDinst_Mcompar__n0367_inst_lut4_401 (
    .ADR0(DLX_MEMinst_reg_dst_out[1]),
    .ADR1(DLX_IDinst_jtarget[21]),
    .ADR2(DLX_IDinst_jtarget[22]),
    .ADR3(DLX_MEMinst_reg_dst_out[0]),
    .O(DLX_IDinst_Mcompar__n0367_inst_lut4_40)
  );
  defparam DLX_IDinst_Mcompar__n0367_inst_lut4_411.INIT = 16'h9009;
  X_LUT4 DLX_IDinst_Mcompar__n0367_inst_lut4_411 (
    .ADR0(DLX_IDinst_jtarget[23]),
    .ADR1(DLX_MEMinst_reg_dst_out[2]),
    .ADR2(DLX_IDinst_jtarget[24]),
    .ADR3(DLX_MEMinst_reg_dst_out[3]),
    .O(DLX_IDinst_Mcompar__n0367_inst_lut4_41)
  );
  X_BUF \DLX_IDinst_Mcompar__n0367_inst_cy_263/COUTUSED  (
    .I(\DLX_IDinst_Mcompar__n0367_inst_cy_263/CYMUXG ),
    .O(DLX_IDinst_Mcompar__n0367_inst_cy_263)
  );
  X_MUX2 DLX_IDinst_Mcompar__n0367_inst_cy_263_2876 (
    .IA(\DLX_IDinst_Mcompar__n0367_inst_cy_263/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mcompar__n0367_inst_cy_262),
    .SEL(DLX_IDinst_Mcompar__n0367_inst_lut4_41),
    .O(\DLX_IDinst_Mcompar__n0367_inst_cy_263/CYMUXG )
  );
  X_ZERO \DLX_IDinst__n0367/LOGIC_ZERO_2877  (
    .O(\DLX_IDinst__n0367/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mcompar__n0367_inst_cy_264 (
    .IA(\DLX_IDinst__n0367/LOGIC_ZERO ),
    .IB(\DLX_IDinst__n0367/CYINIT ),
    .SEL(DLX_IDinst_Mcompar__n0367_inst_lut4_42),
    .O(\DLX_IDinst__n0367/CYMUXF )
  );
  defparam DLX_IDinst_Mcompar__n0367_inst_lut4_421.INIT = 16'hC399;
  X_LUT4 DLX_IDinst_Mcompar__n0367_inst_lut4_421 (
    .ADR0(DLX_IDinst_current_IR[25]),
    .ADR1(DLX_MEMinst_reg_dst_out[4]),
    .ADR2(DLX_IFinst_IR_latched[25]),
    .ADR3(DLX_EXinst__n0144),
    .O(DLX_IDinst_Mcompar__n0367_inst_lut4_42)
  );
  X_BUF \DLX_IDinst__n0367/XBUSED  (
    .I(\DLX_IDinst__n0367/CYMUXF ),
    .O(DLX_IDinst__n0367)
  );
  X_BUF \DLX_IDinst__n0367/CYINIT_2878  (
    .I(DLX_IDinst_Mcompar__n0367_inst_cy_263),
    .O(\DLX_IDinst__n0367/CYINIT )
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<20>1 .INIT = 16'h5C0C;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<20>1  (
    .ADR0(DLX_MEMinst_opcode_of_WB[2]),
    .ADR1(DLX_MEMinst_RF_data_in[20]),
    .ADR2(DLX_IDinst__n0161),
    .ADR3(DLX_IDinst_Mmux__n0162__net105),
    .O(\DLX_IDinst_RegFile_10_20/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_10_20/YUSED  (
    .I(\DLX_IDinst_RegFile_10_20/GROM ),
    .O(DLX_IDinst_WB_data_eff[20])
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<21>1 .INIT = 16'h50D8;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<21>1  (
    .ADR0(DLX_IDinst__n0161),
    .ADR1(DLX_IDinst_Mmux__n0162__net105),
    .ADR2(DLX_MEMinst_RF_data_in[21]),
    .ADR3(DLX_MEMinst_opcode_of_WB[2]),
    .O(\DLX_IDinst_RegFile_10_21/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_10_21/YUSED  (
    .I(\DLX_IDinst_RegFile_10_21/GROM ),
    .O(DLX_IDinst_WB_data_eff[21])
  );
  defparam DLX_IDinst_RegFile_29_29_2879.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_29_29_2879 (
    .I(DLX_IDinst_WB_data_eff[29]),
    .CE(DLX_IDinst__n0608),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_29_29)
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<22>1 .INIT = 16'h44E4;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<22>1  (
    .ADR0(DLX_IDinst__n0161),
    .ADR1(DLX_MEMinst_RF_data_in[22]),
    .ADR2(DLX_IDinst_Mmux__n0162__net105),
    .ADR3(DLX_MEMinst_opcode_of_WB[2]),
    .O(\DLX_IDinst_RegFile_10_22/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_10_22/YUSED  (
    .I(\DLX_IDinst_RegFile_10_22/GROM ),
    .O(DLX_IDinst_WB_data_eff[22])
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<23>1 .INIT = 16'h22E2;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<23>1  (
    .ADR0(DLX_MEMinst_RF_data_in[23]),
    .ADR1(DLX_IDinst__n0161),
    .ADR2(DLX_IDinst_Mmux__n0162__net105),
    .ADR3(DLX_MEMinst_opcode_of_WB[2]),
    .O(\DLX_IDinst_RegFile_10_23/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_10_23/YUSED  (
    .I(\DLX_IDinst_RegFile_10_23/GROM ),
    .O(DLX_IDinst_WB_data_eff[23])
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<31>1 .INIT = 16'h22E2;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<31>1  (
    .ADR0(DLX_MEMinst_RF_data_in[31]),
    .ADR1(DLX_IDinst__n0161),
    .ADR2(DLX_IDinst_Mmux__n0162__net105),
    .ADR3(DLX_MEMinst_opcode_of_WB[2]),
    .O(\DLX_IDinst_RegFile_10_31/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_10_31/YUSED  (
    .I(\DLX_IDinst_RegFile_10_31/GROM ),
    .O(DLX_IDinst_WB_data_eff[31])
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<24>1 .INIT = 16'h7520;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<24>1  (
    .ADR0(DLX_IDinst__n0161),
    .ADR1(DLX_MEMinst_opcode_of_WB[2]),
    .ADR2(DLX_IDinst_Mmux__n0162__net105),
    .ADR3(DLX_MEMinst_RF_data_in[24]),
    .O(\DLX_IDinst_RegFile_10_24/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_10_24/YUSED  (
    .I(\DLX_IDinst_RegFile_10_24/GROM ),
    .O(DLX_IDinst_WB_data_eff[24])
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<16>1 .INIT = 16'h30B8;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<16>1  (
    .ADR0(DLX_IDinst_Mmux__n0162__net105),
    .ADR1(DLX_IDinst__n0161),
    .ADR2(DLX_MEMinst_RF_data_in[16]),
    .ADR3(DLX_MEMinst_opcode_of_WB[2]),
    .O(\DLX_IDinst_RegFile_10_16/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_10_16/YUSED  (
    .I(\DLX_IDinst_RegFile_10_16/GROM ),
    .O(DLX_IDinst_WB_data_eff[16])
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<25>1 .INIT = 16'h7250;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<25>1  (
    .ADR0(DLX_IDinst__n0161),
    .ADR1(DLX_MEMinst_opcode_of_WB[2]),
    .ADR2(DLX_MEMinst_RF_data_in[25]),
    .ADR3(DLX_IDinst_Mmux__n0162__net105),
    .O(\DLX_IDinst_RegFile_10_25/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_10_25/YUSED  (
    .I(\DLX_IDinst_RegFile_10_25/GROM ),
    .O(DLX_IDinst_WB_data_eff[25])
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<17>1 .INIT = 16'h2E22;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<17>1  (
    .ADR0(DLX_MEMinst_RF_data_in[17]),
    .ADR1(DLX_IDinst__n0161),
    .ADR2(DLX_MEMinst_opcode_of_WB[2]),
    .ADR3(DLX_IDinst_Mmux__n0162__net105),
    .O(\DLX_IDinst_RegFile_10_17/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_10_17/YUSED  (
    .I(\DLX_IDinst_RegFile_10_17/GROM ),
    .O(DLX_IDinst_WB_data_eff[17])
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<26>1 .INIT = 16'h0CAA;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<26>1  (
    .ADR0(DLX_MEMinst_RF_data_in[26]),
    .ADR1(DLX_IDinst_Mmux__n0162__net105),
    .ADR2(DLX_MEMinst_opcode_of_WB[2]),
    .ADR3(DLX_IDinst__n0161),
    .O(\DLX_IDinst_RegFile_10_26/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_10_26/YUSED  (
    .I(\DLX_IDinst_RegFile_10_26/GROM ),
    .O(DLX_IDinst_WB_data_eff[26])
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<18>1 .INIT = 16'h44E4;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<18>1  (
    .ADR0(DLX_IDinst__n0161),
    .ADR1(DLX_MEMinst_RF_data_in[18]),
    .ADR2(DLX_IDinst_Mmux__n0162__net105),
    .ADR3(DLX_MEMinst_opcode_of_WB[2]),
    .O(\DLX_IDinst_RegFile_10_18/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_10_18/YUSED  (
    .I(\DLX_IDinst_RegFile_10_18/GROM ),
    .O(DLX_IDinst_WB_data_eff[18])
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<27>1 .INIT = 16'h7430;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<27>1  (
    .ADR0(DLX_MEMinst_opcode_of_WB[2]),
    .ADR1(DLX_IDinst__n0161),
    .ADR2(DLX_MEMinst_RF_data_in[27]),
    .ADR3(DLX_IDinst_Mmux__n0162__net105),
    .O(\DLX_IDinst_RegFile_10_27/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_10_27/YUSED  (
    .I(\DLX_IDinst_RegFile_10_27/GROM ),
    .O(DLX_IDinst_WB_data_eff[27])
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<19>1 .INIT = 16'h7250;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<19>1  (
    .ADR0(DLX_IDinst__n0161),
    .ADR1(DLX_MEMinst_opcode_of_WB[2]),
    .ADR2(DLX_MEMinst_RF_data_in[19]),
    .ADR3(DLX_IDinst_Mmux__n0162__net105),
    .O(\DLX_IDinst_RegFile_10_19/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_10_19/YUSED  (
    .I(\DLX_IDinst_RegFile_10_19/GROM ),
    .O(DLX_IDinst_WB_data_eff[19])
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<28>1 .INIT = 16'h44E4;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<28>1  (
    .ADR0(DLX_IDinst__n0161),
    .ADR1(DLX_MEMinst_RF_data_in[28]),
    .ADR2(DLX_IDinst_Mmux__n0162__net105),
    .ADR3(DLX_MEMinst_opcode_of_WB[2]),
    .O(\DLX_IDinst_RegFile_10_28/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_10_28/YUSED  (
    .I(\DLX_IDinst_RegFile_10_28/GROM ),
    .O(DLX_IDinst_WB_data_eff[28])
  );
  defparam \DLX_IDinst_Mmux_WB_data_eff_Result<29>1 .INIT = 16'h0ACC;
  X_LUT4 \DLX_IDinst_Mmux_WB_data_eff_Result<29>1  (
    .ADR0(DLX_IDinst_Mmux__n0162__net105),
    .ADR1(DLX_MEMinst_RF_data_in[29]),
    .ADR2(DLX_MEMinst_opcode_of_WB[2]),
    .ADR3(DLX_IDinst__n0161),
    .O(\DLX_IDinst_RegFile_10_29/GROM )
  );
  X_BUF \DLX_IDinst_RegFile_10_29/YUSED  (
    .I(\DLX_IDinst_RegFile_10_29/GROM ),
    .O(DLX_IDinst_WB_data_eff[29])
  );
  defparam DLX_IDinst__n0124_2880.INIT = 16'h00C8;
  X_LUT4 DLX_IDinst__n0124_2880 (
    .ADR0(N127400),
    .ADR1(DLX_IDinst_jtarget[10]),
    .ADR2(DLX_IDinst__n0453),
    .ADR3(DLX_IDinst_N108456),
    .O(DLX_IDinst__n0124)
  );
  defparam \DLX_IDinst__n0142<0> .INIT = 16'h00E0;
  X_LUT4 \DLX_IDinst__n0142<0>  (
    .ADR0(N127400),
    .ADR1(DLX_IDinst__n0453),
    .ADR2(DLX_IDinst_IR_latched[26]),
    .ADR3(DLX_IDinst_N108456),
    .O(DLX_IDinst__n0142[0])
  );
  defparam DLX_IDinst__n0125_2881.INIT = 16'h3200;
  X_LUT4 DLX_IDinst__n0125_2881 (
    .ADR0(N127400),
    .ADR1(DLX_IDinst_N108456),
    .ADR2(DLX_IDinst__n0453),
    .ADR3(DLX_IDinst_jtarget[9]),
    .O(DLX_IDinst__n0125)
  );
  defparam \DLX_IDinst__n0142<2> .INIT = 16'h3200;
  X_LUT4 \DLX_IDinst__n0142<2>  (
    .ADR0(N127400),
    .ADR1(DLX_IDinst_N108456),
    .ADR2(DLX_IDinst__n0453),
    .ADR3(DLX_IDinst_IR_latched[28]),
    .O(DLX_IDinst__n0142[2])
  );
  defparam \DLX_IDinst__n0143<4> .INIT = 16'h00E0;
  X_LUT4 \DLX_IDinst__n0143<4>  (
    .ADR0(N127400),
    .ADR1(DLX_IDinst__n0453),
    .ADR2(DLX_IDinst_jtarget[4]),
    .ADR3(DLX_IDinst_Ker1084541_1),
    .O(DLX_IDinst__n0143[4])
  );
  defparam \DLX_IDinst__n0142<5> .INIT = 16'h3200;
  X_LUT4 \DLX_IDinst__n0142<5>  (
    .ADR0(N127652),
    .ADR1(DLX_IDinst_Ker1084541_1),
    .ADR2(DLX_IDinst__n0453),
    .ADR3(DLX_IDinst_IR_latched[31]),
    .O(DLX_IDinst__n0142[5])
  );
  defparam \DLX_EXinst__n0007<10>2491 .INIT = 16'hFCCC;
  X_LUT4 \DLX_EXinst__n0007<10>2491  (
    .ADR0(VCC),
    .ADR1(CHOICE4498),
    .ADR2(DLX_EXinst__n0012[10]),
    .ADR3(DLX_EXinst_N73959),
    .O(\DLX_EXinst_ALU_result_10_1/GROM )
  );
  X_BUF \DLX_EXinst_ALU_result_10_1/YUSED  (
    .I(\DLX_EXinst_ALU_result_10_1/GROM ),
    .O(N162867)
  );
  defparam \DLX_EXinst__n0007<11>2491 .INIT = 16'hFCCC;
  X_LUT4 \DLX_EXinst__n0007<11>2491  (
    .ADR0(VCC),
    .ADR1(CHOICE4438),
    .ADR2(DLX_EXinst_N73959),
    .ADR3(DLX_EXinst__n0012[11]),
    .O(\DLX_EXinst_ALU_result_11_1/GROM )
  );
  X_BUF \DLX_EXinst_ALU_result_11_1/YUSED  (
    .I(\DLX_EXinst_ALU_result_11_1/GROM ),
    .O(N162828)
  );
  defparam \DLX_EXinst__n0007<12>2401 .INIT = 16'hFF88;
  X_LUT4 \DLX_EXinst__n0007<12>2401  (
    .ADR0(DLX_EXinst__n0012[12]),
    .ADR1(DLX_EXinst_N73959),
    .ADR2(VCC),
    .ADR3(CHOICE3813),
    .O(\DLX_EXinst_ALU_result_12_1/GROM )
  );
  X_BUF \DLX_EXinst_ALU_result_12_1/YUSED  (
    .I(\DLX_EXinst_ALU_result_12_1/GROM ),
    .O(N162832)
  );
  defparam \DLX_EXinst__n0007<13>2401 .INIT = 16'hFF88;
  X_LUT4 \DLX_EXinst__n0007<13>2401  (
    .ADR0(DLX_EXinst__n0012[13]),
    .ADR1(DLX_EXinst_N73959),
    .ADR2(VCC),
    .ADR3(CHOICE3758),
    .O(\DLX_EXinst_ALU_result_13_1/GROM )
  );
  X_BUF \DLX_EXinst_ALU_result_13_1/YUSED  (
    .I(\DLX_EXinst_ALU_result_13_1/GROM ),
    .O(N162857)
  );
  defparam \DLX_EXinst__n0007<14>2401 .INIT = 16'hEEAA;
  X_LUT4 \DLX_EXinst__n0007<14>2401  (
    .ADR0(CHOICE3703),
    .ADR1(DLX_EXinst_N73959),
    .ADR2(VCC),
    .ADR3(DLX_EXinst__n0012[14]),
    .O(\DLX_EXinst_ALU_result_14_1/GROM )
  );
  X_BUF \DLX_EXinst_ALU_result_14_1/YUSED  (
    .I(\DLX_EXinst_ALU_result_14_1/GROM ),
    .O(N162813)
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<0>1 .INIT = 16'hF0E2;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<0>1  (
    .ADR0(DLX_IFinst_IR_latched[0]),
    .ADR1(DLX_IDinst_counter[0]),
    .ADR2(DLX_IDinst_current_IR[0]),
    .ADR3(DLX_IDinst_counter[1]),
    .O(\DLX_IDinst_current_IR<0>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<0>/YUSED  (
    .I(\DLX_IDinst_current_IR<0>/GROM ),
    .O(DLX_IDinst_jtarget[0])
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<1>1 .INIT = 16'hCCCA;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<1>1  (
    .ADR0(DLX_IFinst_IR_latched[1]),
    .ADR1(DLX_IDinst_current_IR[1]),
    .ADR2(DLX_IDinst_counter[1]),
    .ADR3(DLX_IDinst_counter[0]),
    .O(\DLX_IDinst_current_IR<1>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<1>/YUSED  (
    .I(\DLX_IDinst_current_IR<1>/GROM ),
    .O(DLX_IDinst_jtarget[1])
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<2>1 .INIT = 16'hF0E2;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<2>1  (
    .ADR0(DLX_IFinst_IR_latched[2]),
    .ADR1(DLX_IDinst_counter[1]),
    .ADR2(DLX_IDinst_current_IR[2]),
    .ADR3(DLX_IDinst_counter[0]),
    .O(\DLX_IDinst_current_IR<2>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<2>/YUSED  (
    .I(\DLX_IDinst_current_IR<2>/GROM ),
    .O(DLX_IDinst_jtarget[2])
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<3>1 .INIT = 16'hCDC8;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<3>1  (
    .ADR0(DLX_IDinst_counter[0]),
    .ADR1(DLX_IDinst_current_IR[3]),
    .ADR2(DLX_IDinst_counter[1]),
    .ADR3(DLX_IFinst_IR_latched[3]),
    .O(\DLX_IDinst_current_IR<3>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<3>/YUSED  (
    .I(\DLX_IDinst_current_IR<3>/GROM ),
    .O(DLX_IDinst_jtarget[3])
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<4>1 .INIT = 16'hFE02;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<4>1  (
    .ADR0(DLX_IFinst_IR_latched[4]),
    .ADR1(DLX_IDinst_counter[0]),
    .ADR2(DLX_IDinst_counter[1]),
    .ADR3(DLX_IDinst_current_IR[4]),
    .O(\DLX_IDinst_current_IR<4>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<4>/YUSED  (
    .I(\DLX_IDinst_current_IR<4>/GROM ),
    .O(DLX_IDinst_jtarget[4])
  );
  defparam \DLX_IDinst__n0145<1>1 .INIT = 16'hC00C;
  X_LUT4 \DLX_IDinst__n0145<1>1  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst__n0387),
    .ADR2(DLX_IDinst_counter[0]),
    .ADR3(DLX_IDinst_counter[1]),
    .O(DLX_IDinst__n0145[1])
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<5>1 .INIT = 16'hFE02;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<5>1  (
    .ADR0(DLX_IFinst_IR_latched[5]),
    .ADR1(DLX_IDinst_counter[0]),
    .ADR2(DLX_IDinst_counter[1]),
    .ADR3(DLX_IDinst_current_IR[5]),
    .O(\DLX_IDinst_current_IR<5>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<5>/YUSED  (
    .I(\DLX_IDinst_current_IR<5>/GROM ),
    .O(DLX_IDinst_jtarget[5])
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<6>1 .INIT = 16'hAAB8;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<6>1  (
    .ADR0(DLX_IDinst_current_IR[6]),
    .ADR1(DLX_IDinst_counter[1]),
    .ADR2(DLX_IFinst_IR_latched[6]),
    .ADR3(DLX_IDinst_counter[0]),
    .O(\DLX_IDinst_current_IR<6>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<6>/YUSED  (
    .I(\DLX_IDinst_current_IR<6>/GROM ),
    .O(DLX_IDinst_jtarget[6])
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<7>1 .INIT = 16'hFE04;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<7>1  (
    .ADR0(DLX_IDinst_counter[1]),
    .ADR1(DLX_IFinst_IR_latched[7]),
    .ADR2(DLX_IDinst_counter[0]),
    .ADR3(DLX_IDinst_current_IR[7]),
    .O(\DLX_IDinst_current_IR<7>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<7>/YUSED  (
    .I(\DLX_IDinst_current_IR<7>/GROM ),
    .O(DLX_IDinst_jtarget[7])
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<8>1 .INIT = 16'hFE04;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<8>1  (
    .ADR0(DLX_IDinst_counter[1]),
    .ADR1(DLX_IFinst_IR_latched[8]),
    .ADR2(DLX_IDinst_counter[0]),
    .ADR3(DLX_IDinst_current_IR[8]),
    .O(\DLX_IDinst_current_IR<8>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<8>/YUSED  (
    .I(\DLX_IDinst_current_IR<8>/GROM ),
    .O(DLX_IDinst_jtarget[8])
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<9>1 .INIT = 16'hF0E4;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<9>1  (
    .ADR0(DLX_IDinst_counter[0]),
    .ADR1(DLX_IFinst_IR_latched[9]),
    .ADR2(DLX_IDinst_current_IR[9]),
    .ADR3(DLX_IDinst_counter[1]),
    .O(\DLX_IDinst_current_IR<9>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<9>/YUSED  (
    .I(\DLX_IDinst_current_IR<9>/GROM ),
    .O(DLX_IDinst_jtarget[9])
  );
  defparam \DLX_EXinst__n0008<9>1 .INIT = 16'hAA00;
  X_LUT4 \DLX_EXinst__n0008<9>1  (
    .ADR0(DLX_IDinst_reg_out_B[9]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N72765),
    .O(DLX_EXinst__n0008[9])
  );
  defparam \DLX_EXinst__n0008<8>1 .INIT = 16'hA0A0;
  X_LUT4 \DLX_EXinst__n0008<8>1  (
    .ADR0(DLX_IDinst_reg_out_B[8]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N72765),
    .ADR3(VCC),
    .O(DLX_EXinst__n0008[8])
  );
  defparam \DLX_EXinst__n0007<8>3011 .INIT = 16'hEECC;
  X_LUT4 \DLX_EXinst__n0007<8>3011  (
    .ADR0(DLX_EXinst_N73959),
    .ADR1(CHOICE5191),
    .ADR2(VCC),
    .ADR3(DLX_EXinst__n0012[8]),
    .O(\DLX_EXinst_ALU_result<8>/GROM )
  );
  X_BUF \DLX_EXinst_ALU_result<8>/YUSED  (
    .I(\DLX_EXinst_ALU_result<8>/GROM ),
    .O(N162844)
  );
  defparam \DLX_EXinst__n0008<11>1 .INIT = 16'h8888;
  X_LUT4 \DLX_EXinst__n0008<11>1  (
    .ADR0(DLX_IDinst_reg_out_B[11]),
    .ADR1(DLX_EXinst_N72765),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst__n0008[11])
  );
  defparam \DLX_EXinst__n0008<10>1 .INIT = 16'h8888;
  X_LUT4 \DLX_EXinst__n0008<10>1  (
    .ADR0(DLX_EXinst_N72765),
    .ADR1(DLX_IDinst_reg_out_B[10]),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst__n0008[10])
  );
  defparam \DLX_EXinst__n0008<13>1 .INIT = 16'hCC00;
  X_LUT4 \DLX_EXinst__n0008<13>1  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N72765),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[13]),
    .O(DLX_EXinst__n0008[13])
  );
  defparam \DLX_EXinst__n0008<12>1 .INIT = 16'hA0A0;
  X_LUT4 \DLX_EXinst__n0008<12>1  (
    .ADR0(DLX_EXinst_N72765),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[12]),
    .ADR3(VCC),
    .O(DLX_EXinst__n0008[12])
  );
  defparam \DLX_EXinst__n0008<16>1 .INIT = 16'hAA00;
  X_LUT4 \DLX_EXinst__n0008<16>1  (
    .ADR0(DLX_EXinst_N72746),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_reg_out_B[16]),
    .O(DLX_EXinst__n0008[16])
  );
  defparam \DLX_EXinst__n0008<20>1 .INIT = 16'hAA00;
  X_LUT4 \DLX_EXinst__n0008<20>1  (
    .ADR0(DLX_IDinst_reg_out_B[20]),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_N72746),
    .O(DLX_EXinst__n0008[20])
  );
  defparam \DLX_EXinst__n0008<17>1 .INIT = 16'hF000;
  X_LUT4 \DLX_EXinst__n0008<17>1  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[17]),
    .ADR3(DLX_EXinst_N72746),
    .O(DLX_EXinst__n0008[17])
  );
  defparam \DLX_EXinst__n0008<21>1 .INIT = 16'hF000;
  X_LUT4 \DLX_EXinst__n0008<21>1  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[21]),
    .ADR3(DLX_EXinst_N72746),
    .O(DLX_EXinst__n0008[21])
  );
  defparam \DLX_EXinst__n0008<14>1 .INIT = 16'hC0C0;
  X_LUT4 \DLX_EXinst__n0008<14>1  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N72765),
    .ADR2(DLX_IDinst_reg_out_B[14]),
    .ADR3(VCC),
    .O(DLX_EXinst__n0008[14])
  );
  defparam \DLX_EXinst__n0008<19>1 .INIT = 16'hA0A0;
  X_LUT4 \DLX_EXinst__n0008<19>1  (
    .ADR0(DLX_IDinst_reg_out_B[19]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N72746),
    .ADR3(VCC),
    .O(DLX_EXinst__n0008[19])
  );
  defparam \DLX_EXinst__n0008<22>1 .INIT = 16'hF000;
  X_LUT4 \DLX_EXinst__n0008<22>1  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N72746),
    .ADR3(DLX_IDinst_reg_out_B[22]),
    .O(DLX_EXinst__n0008[22])
  );
  defparam \DLX_EXinst__n0008<24>1 .INIT = 16'hC0C0;
  X_LUT4 \DLX_EXinst__n0008<24>1  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_N72746),
    .ADR2(DLX_IDinst_reg_out_B[24]),
    .ADR3(VCC),
    .O(DLX_EXinst__n0008[24])
  );
  defparam \DLX_EXinst__n0008<23>1 .INIT = 16'h8888;
  X_LUT4 \DLX_EXinst__n0008<23>1  (
    .ADR0(DLX_IDinst_reg_out_B[23]),
    .ADR1(DLX_EXinst_N72746),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(DLX_EXinst__n0008[23])
  );
  defparam \DLX_EXinst__n0008<27>1 .INIT = 16'hA0A0;
  X_LUT4 \DLX_EXinst__n0008<27>1  (
    .ADR0(DLX_IDinst_reg_out_B[27]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N72746),
    .ADR3(VCC),
    .O(DLX_EXinst__n0008[27])
  );
  defparam \DLX_EXinst__n0008<25>1 .INIT = 16'hF000;
  X_LUT4 \DLX_EXinst__n0008<25>1  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N72746),
    .ADR3(DLX_IDinst_reg_out_B[25]),
    .O(DLX_EXinst__n0008[25])
  );
  defparam \DLX_EXinst__n0008<29>1 .INIT = 16'hA0A0;
  X_LUT4 \DLX_EXinst__n0008<29>1  (
    .ADR0(DLX_EXinst_N72746),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_out_B[29]),
    .ADR3(VCC),
    .O(DLX_EXinst__n0008[29])
  );
  defparam \DLX_EXinst__n0008<28>1 .INIT = 16'hA0A0;
  X_LUT4 \DLX_EXinst__n0008<28>1  (
    .ADR0(DLX_IDinst_reg_out_B[28]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_N72746),
    .ADR3(VCC),
    .O(DLX_EXinst__n0008[28])
  );
  defparam DLX_IDinst__n01551.INIT = 16'h000E;
  X_LUT4 DLX_IDinst__n01551 (
    .ADR0(DLX_IDinst__n0453),
    .ADR1(DLX_IDinst__n0098),
    .ADR2(DLX_IDinst__n0387),
    .ADR3(DLX_IDinst_Ker1084541_1),
    .O(DLX_IDinst__n0155)
  );
  defparam DLX_IDinst__n01191.INIT = 16'h4CCC;
  X_LUT4 DLX_IDinst__n01191 (
    .ADR0(DLX_IDinst_IR_latched[26]),
    .ADR1(DLX_IDinst__n0018[4]),
    .ADR2(DLX_IDinst_IR_latched[27]),
    .ADR3(DLX_IDinst_N108165),
    .O(DLX_IDinst__n0119)
  );
  defparam \DLX_IDinst__n0143<5>1 .INIT = 16'hEAAA;
  X_LUT4 \DLX_IDinst__n0143<5>1  (
    .ADR0(DLX_IDinst__n0025[5]),
    .ADR1(DLX_IDinst_IR_latched[26]),
    .ADR2(DLX_IDinst_IR_latched[27]),
    .ADR3(DLX_IDinst_N108165),
    .O(DLX_IDinst__n0143[5])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<29>1 .INIT = 16'hACAC;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<29>1  (
    .ADR0(DM_read_data[29]),
    .ADR1(DLX_EXinst_ALU_result[29]),
    .ADR2(DLX_EXinst_mem_to_reg_EX),
    .ADR3(VCC),
    .O(DLX_MEMinst__n0000[29])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<10>1 .INIT = 16'hAFA0;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<10>1  (
    .ADR0(DM_read_data[10]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_mem_to_reg_EX),
    .ADR3(DLX_EXinst_ALU_result[10]),
    .O(DLX_MEMinst__n0000[10])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<28>1 .INIT = 16'hDD88;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<28>1  (
    .ADR0(DLX_EXinst_mem_to_reg_EX),
    .ADR1(DM_read_data[28]),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_ALU_result[28]),
    .O(DLX_MEMinst__n0000[28])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<11>1 .INIT = 16'hE4E4;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<11>1  (
    .ADR0(DLX_EXinst_mem_to_reg_EX),
    .ADR1(DLX_EXinst_ALU_result[11]),
    .ADR2(DM_read_data[11]),
    .ADR3(VCC),
    .O(DLX_MEMinst__n0000[11])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<27>1 .INIT = 16'hCCAA;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<27>1  (
    .ADR0(DLX_EXinst_ALU_result[27]),
    .ADR1(DM_read_data[27]),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_mem_to_reg_EX),
    .O(DLX_MEMinst__n0000[27])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<20>1 .INIT = 16'hF0CC;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<20>1  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_ALU_result[20]),
    .ADR2(DM_read_data[20]),
    .ADR3(DLX_EXinst_mem_to_reg_EX),
    .O(DLX_MEMinst__n0000[20])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<26>1 .INIT = 16'hE4E4;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<26>1  (
    .ADR0(DLX_EXinst_mem_to_reg_EX),
    .ADR1(DLX_EXinst_ALU_result[26]),
    .ADR2(DM_read_data[26]),
    .ADR3(VCC),
    .O(DLX_MEMinst__n0000[26])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<12>1 .INIT = 16'hFC30;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<12>1  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_mem_to_reg_EX),
    .ADR2(DLX_EXinst_ALU_result[12]),
    .ADR3(DM_read_data[12]),
    .O(DLX_MEMinst__n0000[12])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<25>1 .INIT = 16'hEE44;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<25>1  (
    .ADR0(DLX_EXinst_mem_to_reg_EX),
    .ADR1(DLX_EXinst_ALU_result[25]),
    .ADR2(VCC),
    .ADR3(DM_read_data[25]),
    .O(DLX_MEMinst__n0000[25])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<21>1 .INIT = 16'hE4E4;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<21>1  (
    .ADR0(DLX_EXinst_mem_to_reg_EX),
    .ADR1(DLX_EXinst_ALU_result[21]),
    .ADR2(DM_read_data[21]),
    .ADR3(VCC),
    .O(DLX_MEMinst__n0000[21])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<23>1 .INIT = 16'hCACA;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<23>1  (
    .ADR0(DLX_EXinst_ALU_result[23]),
    .ADR1(DM_read_data[23]),
    .ADR2(DLX_EXinst_mem_to_reg_EX),
    .ADR3(VCC),
    .O(DLX_MEMinst__n0000[23])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<13>1 .INIT = 16'hCFC0;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<13>1  (
    .ADR0(VCC),
    .ADR1(DM_read_data[13]),
    .ADR2(DLX_EXinst_mem_to_reg_EX),
    .ADR3(DLX_EXinst_ALU_result[13]),
    .O(DLX_MEMinst__n0000[13])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<22>1 .INIT = 16'hF0AA;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<22>1  (
    .ADR0(DLX_EXinst_ALU_result[22]),
    .ADR1(VCC),
    .ADR2(DM_read_data[22]),
    .ADR3(DLX_EXinst_mem_to_reg_EX),
    .O(DLX_MEMinst__n0000[22])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<30>1 .INIT = 16'hBB88;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<30>1  (
    .ADR0(DM_read_data[30]),
    .ADR1(DLX_EXinst_mem_to_reg_EX),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_ALU_result[30]),
    .O(DLX_MEMinst__n0000[30])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<19>1 .INIT = 16'hBB88;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<19>1  (
    .ADR0(DM_read_data[19]),
    .ADR1(DLX_EXinst_mem_to_reg_EX),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_ALU_result[19]),
    .O(DLX_MEMinst__n0000[19])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<14>1 .INIT = 16'hFC30;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<14>1  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_mem_to_reg_EX),
    .ADR2(DLX_EXinst_ALU_result[14]),
    .ADR3(DM_read_data[14]),
    .O(DLX_MEMinst__n0000[14])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<18>1 .INIT = 16'hCACA;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<18>1  (
    .ADR0(DLX_EXinst_ALU_result[18]),
    .ADR1(DM_read_data[18]),
    .ADR2(DLX_EXinst_mem_to_reg_EX),
    .ADR3(VCC),
    .O(DLX_MEMinst__n0000[18])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<15>1 .INIT = 16'hF0AA;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<15>1  (
    .ADR0(DLX_EXinst_ALU_result[15]),
    .ADR1(VCC),
    .ADR2(DM_read_data[15]),
    .ADR3(DLX_EXinst_mem_to_reg_EX),
    .O(DLX_MEMinst__n0000[15])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<17>1 .INIT = 16'hF0AA;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<17>1  (
    .ADR0(DLX_EXinst_ALU_result[17]),
    .ADR1(VCC),
    .ADR2(DM_read_data[17]),
    .ADR3(DLX_EXinst_mem_to_reg_EX),
    .O(DLX_MEMinst__n0000[17])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<31>1 .INIT = 16'hF0AA;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<31>1  (
    .ADR0(DLX_EXinst_ALU_result[31]),
    .ADR1(VCC),
    .ADR2(DM_read_data[31]),
    .ADR3(DLX_EXinst_mem_to_reg_EX),
    .O(DLX_MEMinst__n0000[31])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<9>1 .INIT = 16'hF0CC;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<9>1  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_ALU_result[9]),
    .ADR2(DM_read_data[9]),
    .ADR3(DLX_EXinst_mem_to_reg_EX),
    .O(DLX_MEMinst__n0000[9])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<16>1 .INIT = 16'hCCF0;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<16>1  (
    .ADR0(VCC),
    .ADR1(DM_read_data[16]),
    .ADR2(DLX_EXinst_ALU_result[16]),
    .ADR3(DLX_EXinst_mem_to_reg_EX),
    .O(DLX_MEMinst__n0000[16])
  );
  defparam DLX_IDinst__n0126_2882.INIT = 16'h5400;
  X_LUT4 DLX_IDinst__n0126_2882 (
    .ADR0(DLX_IDinst_N108456),
    .ADR1(N127400),
    .ADR2(DLX_IDinst__n0453),
    .ADR3(DLX_IDinst_jtarget[8]),
    .O(DLX_IDinst__n0126)
  );
  defparam \DLX_IDinst__n0135<0> .INIT = 16'h00C8;
  X_LUT4 \DLX_IDinst__n0135<0>  (
    .ADR0(N127400),
    .ADR1(DLX_IDinst_jtarget[16]),
    .ADR2(DLX_IDinst__n0453),
    .ADR3(DLX_IDinst_N108456),
    .O(DLX_IDinst__n0135[0])
  );
  defparam DLX_IFinst_IR_previous_26.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_26 (
    .I(DLX_IFinst_IR_latched[26]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[26])
  );
  defparam DLX_IDinst__n0127_2883.INIT = 16'h4440;
  X_LUT4 DLX_IDinst__n0127_2883 (
    .ADR0(DLX_IDinst_N108456),
    .ADR1(DLX_IDinst_jtarget[7]),
    .ADR2(DLX_IDinst__n0453),
    .ADR3(N127400),
    .O(DLX_IDinst__n0127)
  );
  defparam \DLX_IDinst__n0135<1> .INIT = 16'h2220;
  X_LUT4 \DLX_IDinst__n0135<1>  (
    .ADR0(DLX_IDinst_jtarget[17]),
    .ADR1(DLX_IDinst_N108456),
    .ADR2(DLX_IDinst__n0453),
    .ADR3(N127400),
    .O(DLX_IDinst__n0135[1])
  );
  defparam DLX_IDinst__n0128_2884.INIT = 16'h5400;
  X_LUT4 DLX_IDinst__n0128_2884 (
    .ADR0(DLX_IDinst_N108456),
    .ADR1(DLX_IDinst__n0453),
    .ADR2(N127400),
    .ADR3(DLX_IDinst_jtarget[6]),
    .O(DLX_IDinst__n0128)
  );
  defparam \DLX_IDinst__n0135<2> .INIT = 16'h3200;
  X_LUT4 \DLX_IDinst__n0135<2>  (
    .ADR0(DLX_IDinst__n0453),
    .ADR1(DLX_IDinst_N108456),
    .ADR2(N127400),
    .ADR3(DLX_IDinst_jtarget[18]),
    .O(DLX_IDinst__n0135[2])
  );
  defparam \DLX_IDinst__n0135<3> .INIT = 16'h3200;
  X_LUT4 \DLX_IDinst__n0135<3>  (
    .ADR0(N127400),
    .ADR1(DLX_IDinst_N108456),
    .ADR2(DLX_IDinst__n0453),
    .ADR3(DLX_IDinst_jtarget[19]),
    .O(DLX_IDinst__n0135[3])
  );
  defparam \DLX_IDinst__n0143<1> .INIT = 16'h00C8;
  X_LUT4 \DLX_IDinst__n0143<1>  (
    .ADR0(N127400),
    .ADR1(DLX_IDinst_jtarget[1]),
    .ADR2(DLX_IDinst__n0453),
    .ADR3(DLX_IDinst_Ker1084541_1),
    .O(\DLX_IDinst_Imm<1>/GROM )
  );
  X_BUF \DLX_IDinst_Imm<1>/YUSED  (
    .I(\DLX_IDinst_Imm<1>/GROM ),
    .O(DLX_IDinst__n0143[1])
  );
  defparam \DLX_IDinst__n0143<2> .INIT = 16'h00A8;
  X_LUT4 \DLX_IDinst__n0143<2>  (
    .ADR0(DLX_IDinst_jtarget[2]),
    .ADR1(N127400),
    .ADR2(DLX_IDinst__n0453),
    .ADR3(DLX_IDinst_Ker1084541_1),
    .O(\DLX_IDinst_Imm<2>/GROM )
  );
  X_BUF \DLX_IDinst_Imm<2>/YUSED  (
    .I(\DLX_IDinst_Imm<2>/GROM ),
    .O(DLX_IDinst__n0143[2])
  );
  defparam \DLX_IDinst__n0143<3> .INIT = 16'h5040;
  X_LUT4 \DLX_IDinst__n0143<3>  (
    .ADR0(DLX_IDinst_Ker1084541_1),
    .ADR1(N127400),
    .ADR2(DLX_IDinst_jtarget[3]),
    .ADR3(DLX_IDinst__n0453),
    .O(\DLX_IDinst_Imm<3>/GROM )
  );
  X_BUF \DLX_IDinst_Imm<3>/YUSED  (
    .I(\DLX_IDinst_Imm<3>/GROM ),
    .O(DLX_IDinst__n0143[3])
  );
  defparam DLX_IDinst__n0140_2885.INIT = 16'h2000;
  X_LUT4 DLX_IDinst__n0140_2885 (
    .ADR0(N139563),
    .ADR1(N127137),
    .ADR2(DLX_IDinst__n0163),
    .ADR3(DLX_IDinst__n0164),
    .O(DLX_IDinst__n0140)
  );
  defparam DLX_IDinst__n01531.INIT = 16'hD8DC;
  X_LUT4 DLX_IDinst__n01531 (
    .ADR0(DLX_IDinst_Ker1084541_1),
    .ADR1(DLX_IDinst_CLI),
    .ADR2(DLX_IDinst__n0453),
    .ADR3(DLX_IDinst__n0098),
    .O(\DLX_IDinst_CLI/GROM )
  );
  X_BUF \DLX_IDinst_CLI/YUSED  (
    .I(\DLX_IDinst_CLI/GROM ),
    .O(DLX_IDinst__n0153)
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<10>1 .INIT = 16'hCCCA;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<10>1  (
    .ADR0(DLX_IFinst_IR_latched[10]),
    .ADR1(DLX_IDinst_current_IR[10]),
    .ADR2(DLX_IDinst_counter[1]),
    .ADR3(DLX_IDinst_counter[0]),
    .O(\DLX_IDinst_current_IR<10>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<10>/YUSED  (
    .I(\DLX_IDinst_current_IR<10>/GROM ),
    .O(DLX_IDinst_jtarget[10])
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<11>1 .INIT = 16'hCCCA;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<11>1  (
    .ADR0(DLX_IFinst_IR_latched[11]),
    .ADR1(DLX_IDinst_current_IR[11]),
    .ADR2(DLX_IDinst_counter[1]),
    .ADR3(DLX_IDinst_counter[0]),
    .O(\DLX_IDinst_current_IR<11>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<11>/YUSED  (
    .I(\DLX_IDinst_current_IR<11>/GROM ),
    .O(DLX_IDinst_jtarget[11])
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<20>1 .INIT = 16'hABA8;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<20>1  (
    .ADR0(DLX_IDinst_current_IR[20]),
    .ADR1(DLX_IDinst_counter[0]),
    .ADR2(DLX_IDinst_counter[1]),
    .ADR3(DLX_IFinst_IR_latched[20]),
    .O(\DLX_IDinst_current_IR<20>/FROM )
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_581.INIT = 16'h8000;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_581 (
    .ADR0(DLX_IDinst_jtarget[18]),
    .ADR1(DLX_IDinst_jtarget[19]),
    .ADR2(DLX_IDinst_jtarget[17]),
    .ADR3(DLX_IDinst_jtarget[20]),
    .O(\DLX_IDinst_current_IR<20>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<20>/XUSED  (
    .I(\DLX_IDinst_current_IR<20>/FROM ),
    .O(DLX_IDinst_jtarget[20])
  );
  X_BUF \DLX_IDinst_current_IR<20>/YUSED  (
    .I(\DLX_IDinst_current_IR<20>/GROM ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_58)
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<12>1 .INIT = 16'hCCD8;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<12>1  (
    .ADR0(DLX_IDinst_counter[0]),
    .ADR1(DLX_IDinst_current_IR[12]),
    .ADR2(DLX_IFinst_IR_latched[12]),
    .ADR3(DLX_IDinst_counter[1]),
    .O(\DLX_IDinst_current_IR<12>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<12>/YUSED  (
    .I(\DLX_IDinst_current_IR<12>/GROM ),
    .O(DLX_IDinst_jtarget[12])
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<13>1 .INIT = 16'hFE02;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<13>1  (
    .ADR0(DLX_IFinst_IR_latched[13]),
    .ADR1(DLX_IDinst_counter[0]),
    .ADR2(DLX_IDinst_counter[1]),
    .ADR3(DLX_IDinst_current_IR[13]),
    .O(\DLX_IDinst_current_IR<13>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<13>/YUSED  (
    .I(\DLX_IDinst_current_IR<13>/GROM ),
    .O(DLX_IDinst_jtarget[13])
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<30>1 .INIT = 16'hF1E0;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<30>1  (
    .ADR0(DLX_IDinst_counter[0]),
    .ADR1(DLX_IDinst_counter[1]),
    .ADR2(DLX_IDinst_current_IR[30]),
    .ADR3(DLX_IFinst_IR_latched[30]),
    .O(\DLX_IDinst_current_IR<30>/FROM )
  );
  defparam DLX_IDinst_Ker107607.INIT = 16'hC0EA;
  X_LUT4 DLX_IDinst_Ker107607 (
    .ADR0(N136696),
    .ADR1(DLX_IDinst_N108574),
    .ADR2(DLX_IDinst_N108221),
    .ADR3(DLX_IDinst_IR_latched[30]),
    .O(\DLX_IDinst_current_IR<30>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<30>/XUSED  (
    .I(\DLX_IDinst_current_IR<30>/FROM ),
    .O(DLX_IDinst_IR_latched[30])
  );
  X_BUF \DLX_IDinst_current_IR<30>/YUSED  (
    .I(\DLX_IDinst_current_IR<30>/GROM ),
    .O(DLX_IDinst_N107609)
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<14>1 .INIT = 16'hF1E0;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<14>1  (
    .ADR0(DLX_IDinst_counter[0]),
    .ADR1(DLX_IDinst_counter[1]),
    .ADR2(DLX_IDinst_current_IR[14]),
    .ADR3(DLX_IFinst_IR_latched[14]),
    .O(\DLX_IDinst_current_IR<14>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<14>/YUSED  (
    .I(\DLX_IDinst_current_IR<14>/GROM ),
    .O(DLX_IDinst_jtarget[14])
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<22>1 .INIT = 16'hCDC8;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<22>1  (
    .ADR0(DLX_IDinst_counter[1]),
    .ADR1(DLX_IDinst_current_IR[22]),
    .ADR2(DLX_IDinst_counter[0]),
    .ADR3(DLX_IFinst_IR_latched[22]),
    .O(\DLX_IDinst_current_IR<22>/FROM )
  );
  defparam \DLX_IDinst__n0146<6>39 .INIT = 16'h3088;
  X_LUT4 \DLX_IDinst__n0146<6>39  (
    .ADR0(\DLX_IDinst_Cause_Reg[6] ),
    .ADR1(DLX_IDinst_jtarget[21]),
    .ADR2(DLX_IDinst_EPC[6]),
    .ADR3(DLX_IDinst_jtarget[22]),
    .O(\DLX_IDinst_current_IR<22>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<22>/XUSED  (
    .I(\DLX_IDinst_current_IR<22>/FROM ),
    .O(DLX_IDinst_jtarget[22])
  );
  X_BUF \DLX_IDinst_current_IR<22>/YUSED  (
    .I(\DLX_IDinst_current_IR<22>/GROM ),
    .O(CHOICE3211)
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<23>1 .INIT = 16'hFE10;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<23>1  (
    .ADR0(DLX_IDinst_counter[1]),
    .ADR1(DLX_IDinst_counter[0]),
    .ADR2(DLX_IFinst_IR_latched[23]),
    .ADR3(DLX_IDinst_current_IR[23]),
    .O(\DLX_IDinst_current_IR<23>/FROM )
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_5831.INIT = 16'h0008;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_5831 (
    .ADR0(DLX_IDinst_jtarget[24]),
    .ADR1(DLX_IDinst_jtarget[25]),
    .ADR2(DLX_IDinst_jtarget[22]),
    .ADR3(DLX_IDinst_jtarget[23]),
    .O(\DLX_IDinst_current_IR<23>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<23>/XUSED  (
    .I(\DLX_IDinst_current_IR<23>/FROM ),
    .O(DLX_IDinst_jtarget[23])
  );
  X_BUF \DLX_IDinst_current_IR<23>/YUSED  (
    .I(\DLX_IDinst_current_IR<23>/GROM ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_583)
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<31>1 .INIT = 16'hCDC8;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<31>1  (
    .ADR0(DLX_IDinst_counter[0]),
    .ADR1(DLX_IDinst_current_IR[31]),
    .ADR2(DLX_IDinst_counter[1]),
    .ADR3(DLX_IFinst_IR_latched[31]),
    .O(\DLX_IDinst_current_IR<31>/FROM )
  );
  defparam DLX_IDinst_Ker1084741.INIT = 16'h5300;
  X_LUT4 DLX_IDinst_Ker1084741 (
    .ADR0(DLX_IFinst_IR_latched[30]),
    .ADR1(DLX_IDinst_current_IR[30]),
    .ADR2(DLX_EXinst__n0144),
    .ADR3(DLX_IDinst_IR_latched[31]),
    .O(\DLX_IDinst_current_IR<31>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<31>/XUSED  (
    .I(\DLX_IDinst_current_IR<31>/FROM ),
    .O(DLX_IDinst_IR_latched[31])
  );
  X_BUF \DLX_IDinst_current_IR<31>/YUSED  (
    .I(\DLX_IDinst_current_IR<31>/GROM ),
    .O(DLX_IDinst_N108476)
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<15>1 .INIT = 16'hF0E2;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<15>1  (
    .ADR0(DLX_IFinst_IR_latched[15]),
    .ADR1(DLX_IDinst_counter[1]),
    .ADR2(DLX_IDinst_current_IR[15]),
    .ADR3(DLX_IDinst_counter[0]),
    .O(\DLX_IDinst_current_IR<15>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<15>/YUSED  (
    .I(\DLX_IDinst_current_IR<15>/GROM ),
    .O(DLX_IDinst_jtarget[15])
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<24>1 .INIT = 16'hF0E2;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<24>1  (
    .ADR0(DLX_IFinst_IR_latched[24]),
    .ADR1(DLX_IDinst_counter[1]),
    .ADR2(DLX_IDinst_current_IR[24]),
    .ADR3(DLX_IDinst_counter[0]),
    .O(\DLX_IDinst_current_IR<24>/FROM )
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_5791.INIT = 16'h0004;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_5791 (
    .ADR0(DLX_IDinst_jtarget[23]),
    .ADR1(DLX_IDinst_jtarget[25]),
    .ADR2(DLX_IDinst_jtarget[22]),
    .ADR3(DLX_IDinst_jtarget[24]),
    .O(\DLX_IDinst_current_IR<24>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<24>/XUSED  (
    .I(\DLX_IDinst_current_IR<24>/FROM ),
    .O(DLX_IDinst_jtarget[24])
  );
  X_BUF \DLX_IDinst_current_IR<24>/YUSED  (
    .I(\DLX_IDinst_current_IR<24>/GROM ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_579)
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<25>1 .INIT = 16'hF0E2;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<25>1  (
    .ADR0(DLX_IFinst_IR_latched[25]),
    .ADR1(DLX_IDinst_counter[1]),
    .ADR2(DLX_IDinst_current_IR[25]),
    .ADR3(DLX_IDinst_counter[0]),
    .O(\DLX_IDinst_current_IR<25>/FROM )
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_5711.INIT = 16'h0001;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_5711 (
    .ADR0(DLX_IDinst_jtarget[23]),
    .ADR1(DLX_IDinst_jtarget[22]),
    .ADR2(DLX_IDinst_jtarget[24]),
    .ADR3(DLX_IDinst_jtarget[25]),
    .O(\DLX_IDinst_current_IR<25>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<25>/XUSED  (
    .I(\DLX_IDinst_current_IR<25>/FROM ),
    .O(DLX_IDinst_jtarget[25])
  );
  X_BUF \DLX_IDinst_current_IR<25>/YUSED  (
    .I(\DLX_IDinst_current_IR<25>/GROM ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_571)
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<17>1 .INIT = 16'hCDC8;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<17>1  (
    .ADR0(DLX_IDinst_counter[0]),
    .ADR1(DLX_IDinst_current_IR[17]),
    .ADR2(DLX_IDinst_counter[1]),
    .ADR3(DLX_IFinst_IR_latched[17]),
    .O(\DLX_IDinst_current_IR<17>/FROM )
  );
  defparam DLX_IDinst__n0381_SW0.INIT = 16'hFFCC;
  X_LUT4 DLX_IDinst__n0381_SW0 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_jtarget[16]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_jtarget[17]),
    .O(\DLX_IDinst_current_IR<17>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<17>/XUSED  (
    .I(\DLX_IDinst_current_IR<17>/FROM ),
    .O(DLX_IDinst_jtarget[17])
  );
  X_BUF \DLX_IDinst_current_IR<17>/YUSED  (
    .I(\DLX_IDinst_current_IR<17>/GROM ),
    .O(N126925)
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<26>1 .INIT = 16'hF0E2;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<26>1  (
    .ADR0(DLX_IFinst_IR_latched[26]),
    .ADR1(DLX_IDinst_counter[0]),
    .ADR2(DLX_IDinst_current_IR[26]),
    .ADR3(DLX_IDinst_counter[1]),
    .O(\DLX_IDinst_current_IR<26>/FROM )
  );
  defparam DLX_IDinst__n00981.INIT = 16'h0020;
  X_LUT4 DLX_IDinst__n00981 (
    .ADR0(DLX_IDinst_N108165),
    .ADR1(DLX_IDinst_IR_latched[27]),
    .ADR2(DLX_IDinst_IR_latched[30]),
    .ADR3(DLX_IDinst_IR_latched[26]),
    .O(\DLX_IDinst_current_IR<26>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<26>/XUSED  (
    .I(\DLX_IDinst_current_IR<26>/FROM ),
    .O(DLX_IDinst_IR_latched[26])
  );
  X_BUF \DLX_IDinst_current_IR<26>/YUSED  (
    .I(\DLX_IDinst_current_IR<26>/GROM ),
    .O(DLX_IDinst__n0098)
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<18>1 .INIT = 16'hAAB8;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<18>1  (
    .ADR0(DLX_IDinst_current_IR[18]),
    .ADR1(DLX_IDinst_counter[1]),
    .ADR2(DLX_IFinst_IR_latched[18]),
    .ADR3(DLX_IDinst_counter[0]),
    .O(\DLX_IDinst_current_IR<18>/FROM )
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5510.INIT = 16'h0020;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5510 (
    .ADR0(DLX_IDinst_jtarget[19]),
    .ADR1(DLX_IDinst_jtarget[17]),
    .ADR2(DLX_IDinst_jtarget[20]),
    .ADR3(DLX_IDinst_jtarget[18]),
    .O(\DLX_IDinst_current_IR<18>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<18>/XUSED  (
    .I(\DLX_IDinst_current_IR<18>/FROM ),
    .O(DLX_IDinst_jtarget[18])
  );
  X_BUF \DLX_IDinst_current_IR<18>/YUSED  (
    .I(\DLX_IDinst_current_IR<18>/GROM ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_55)
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<27>1 .INIT = 16'hAAAC;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<27>1  (
    .ADR0(DLX_IDinst_current_IR[27]),
    .ADR1(DLX_IFinst_IR_latched[27]),
    .ADR2(DLX_IDinst_counter[0]),
    .ADR3(DLX_IDinst_counter[1]),
    .O(\DLX_IDinst_current_IR<27>/FROM )
  );
  defparam DLX_IDinst__n03131.INIT = 16'h0001;
  X_LUT4 DLX_IDinst__n03131 (
    .ADR0(DLX_IDinst_IR_latched[30]),
    .ADR1(DLX_IDinst_IR_latched[28]),
    .ADR2(DLX_IDinst_IR_latched[26]),
    .ADR3(DLX_IDinst_IR_latched[27]),
    .O(\DLX_IDinst_current_IR<27>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<27>/XUSED  (
    .I(\DLX_IDinst_current_IR<27>/FROM ),
    .O(DLX_IDinst_IR_latched[27])
  );
  X_BUF \DLX_IDinst_current_IR<27>/YUSED  (
    .I(\DLX_IDinst_current_IR<27>/GROM ),
    .O(DLX_IDinst__n0313)
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<19>1 .INIT = 16'hF0E2;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<19>1  (
    .ADR0(DLX_IFinst_IR_latched[19]),
    .ADR1(DLX_IDinst_counter[1]),
    .ADR2(DLX_IDinst_current_IR[19]),
    .ADR3(DLX_IDinst_counter[0]),
    .O(\DLX_IDinst_current_IR<19>/FROM )
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5110.INIT = 16'h0004;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5110 (
    .ADR0(DLX_IDinst_jtarget[18]),
    .ADR1(DLX_IDinst_jtarget[20]),
    .ADR2(DLX_IDinst_jtarget[17]),
    .ADR3(DLX_IDinst_jtarget[19]),
    .O(\DLX_IDinst_current_IR<19>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<19>/XUSED  (
    .I(\DLX_IDinst_current_IR<19>/FROM ),
    .O(DLX_IDinst_jtarget[19])
  );
  X_BUF \DLX_IDinst_current_IR<19>/YUSED  (
    .I(\DLX_IDinst_current_IR<19>/GROM ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_51)
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<28>1 .INIT = 16'hCDC8;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<28>1  (
    .ADR0(DLX_IDinst_counter[0]),
    .ADR1(DLX_IDinst_current_IR[28]),
    .ADR2(DLX_IDinst_counter[1]),
    .ADR3(DLX_IFinst_IR_latched[28]),
    .O(\DLX_IDinst_current_IR<28>/FROM )
  );
  defparam DLX_IDinst__n04271.INIT = 16'h00C4;
  X_LUT4 DLX_IDinst__n04271 (
    .ADR0(DLX_IDinst_IR_latched[27]),
    .ADR1(DLX_IDinst_IR_latched[29]),
    .ADR2(DLX_IDinst_IR_latched[26]),
    .ADR3(DLX_IDinst_IR_latched[28]),
    .O(\DLX_IDinst_current_IR<28>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<28>/XUSED  (
    .I(\DLX_IDinst_current_IR<28>/FROM ),
    .O(DLX_IDinst_IR_latched[28])
  );
  X_BUF \DLX_IDinst_current_IR<28>/YUSED  (
    .I(\DLX_IDinst_current_IR<28>/GROM ),
    .O(DLX_IDinst__n0427)
  );
  defparam \DLX_IDinst_Mmux_IR_latched_Result<29>1 .INIT = 16'hFE10;
  X_LUT4 \DLX_IDinst_Mmux_IR_latched_Result<29>1  (
    .ADR0(DLX_IDinst_counter[1]),
    .ADR1(DLX_IDinst_counter[0]),
    .ADR2(DLX_IFinst_IR_latched[29]),
    .ADR3(DLX_IDinst_current_IR[29]),
    .O(\DLX_IDinst_current_IR<29>/FROM )
  );
  defparam DLX_IDinst_Ker1084411.INIT = 16'h0033;
  X_LUT4 DLX_IDinst_Ker1084411 (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_IR_latched[31]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_IR_latched[29]),
    .O(\DLX_IDinst_current_IR<29>/GROM )
  );
  X_BUF \DLX_IDinst_current_IR<29>/XUSED  (
    .I(\DLX_IDinst_current_IR<29>/FROM ),
    .O(DLX_IDinst_IR_latched[29])
  );
  X_BUF \DLX_IDinst_current_IR<29>/YUSED  (
    .I(\DLX_IDinst_current_IR<29>/GROM ),
    .O(DLX_IDinst_N108443)
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<8>1 .INIT = 16'hAFA0;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<8>1  (
    .ADR0(DM_read_data[8]),
    .ADR1(VCC),
    .ADR2(DLX_EXinst_mem_to_reg_EX),
    .ADR3(DLX_EXinst_ALU_result[8]),
    .O(DLX_MEMinst__n0000[8])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<0>1 .INIT = 16'hCFC0;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<0>1  (
    .ADR0(VCC),
    .ADR1(DM_read_data[0]),
    .ADR2(DLX_EXinst_mem_to_reg_EX),
    .ADR3(DLX_EXinst_ALU_result[0]),
    .O(DLX_MEMinst__n0000[0])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<7>1 .INIT = 16'hF3C0;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<7>1  (
    .ADR0(VCC),
    .ADR1(DLX_EXinst_mem_to_reg_EX),
    .ADR2(DM_read_data[7]),
    .ADR3(DLX_EXinst_ALU_result[7]),
    .O(DLX_MEMinst__n0000[7])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<1>1 .INIT = 16'hF5A0;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<1>1  (
    .ADR0(DLX_EXinst_mem_to_reg_EX),
    .ADR1(VCC),
    .ADR2(DM_read_data[1]),
    .ADR3(DLX_EXinst_ALU_result[1]),
    .O(DLX_MEMinst__n0000[1])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<6>1 .INIT = 16'hB8B8;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<6>1  (
    .ADR0(DM_read_data[6]),
    .ADR1(DLX_EXinst_mem_to_reg_EX),
    .ADR2(DLX_EXinst_ALU_result[6]),
    .ADR3(VCC),
    .O(DLX_MEMinst__n0000[6])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<2>1 .INIT = 16'hDD88;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<2>1  (
    .ADR0(DLX_EXinst_mem_to_reg_EX),
    .ADR1(DM_read_data[2]),
    .ADR2(VCC),
    .ADR3(DLX_EXinst_ALU_result[2]),
    .O(DLX_MEMinst__n0000[2])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<5>1 .INIT = 16'hD8D8;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<5>1  (
    .ADR0(DLX_EXinst_mem_to_reg_EX),
    .ADR1(DM_read_data[5]),
    .ADR2(DLX_EXinst_ALU_result[5]),
    .ADR3(VCC),
    .O(DLX_MEMinst__n0000[5])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<3>1 .INIT = 16'hF5A0;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<3>1  (
    .ADR0(DLX_EXinst_mem_to_reg_EX),
    .ADR1(VCC),
    .ADR2(DM_read_data[3]),
    .ADR3(DLX_EXinst_ALU_result[3]),
    .O(DLX_MEMinst__n0000[3])
  );
  defparam \DLX_MEMinst_Mmux__n0000_Result<4>1 .INIT = 16'hCFC0;
  X_LUT4 \DLX_MEMinst_Mmux__n0000_Result<4>1  (
    .ADR0(VCC),
    .ADR1(DM_read_data[4]),
    .ADR2(DLX_EXinst_mem_to_reg_EX),
    .ADR3(DLX_EXinst_ALU_result[4]),
    .O(DLX_MEMinst__n0000[4])
  );
  defparam DLX_IDinst__n01201.INIT = 16'h7F00;
  X_LUT4 DLX_IDinst__n01201 (
    .ADR0(DLX_IDinst_IR_latched[26]),
    .ADR1(DLX_IDinst_N108165),
    .ADR2(DLX_IDinst_IR_latched[27]),
    .ADR3(DLX_IDinst__n0018[3]),
    .O(DLX_IDinst__n0120)
  );
  defparam DLX_IDinst__n01231.INIT = 16'h70F0;
  X_LUT4 DLX_IDinst__n01231 (
    .ADR0(DLX_IDinst_IR_latched[26]),
    .ADR1(DLX_IDinst_N108165),
    .ADR2(DLX_IDinst__n0018[0]),
    .ADR3(DLX_IDinst_IR_latched[27]),
    .O(DLX_IDinst__n0123)
  );
  defparam DLX_IDinst__n01211.INIT = 16'h4CCC;
  X_LUT4 DLX_IDinst__n01211 (
    .ADR0(DLX_IDinst_IR_latched[27]),
    .ADR1(DLX_IDinst__n0018[2]),
    .ADR2(DLX_IDinst_IR_latched[26]),
    .ADR3(DLX_IDinst_N108165),
    .O(DLX_IDinst__n0121)
  );
  defparam DLX_IDinst__n01221.INIT = 16'h4CCC;
  X_LUT4 DLX_IDinst__n01221 (
    .ADR0(DLX_IDinst_N108165),
    .ADR1(DLX_IDinst__n0018[1]),
    .ADR2(DLX_IDinst_IR_latched[26]),
    .ADR3(DLX_IDinst_IR_latched[27]),
    .O(DLX_IDinst__n0122)
  );
  defparam \DLX_IDinst__n0147<2>1 .INIT = 16'hA280;
  X_LUT4 \DLX_IDinst__n0147<2>1  (
    .ADR0(DLX_IDinst_N107173),
    .ADR1(DLX_IDinst__n0176),
    .ADR2(DLX_MEMinst_RF_data_in[2]),
    .ADR3(DLX_IDinst__n0623[2]),
    .O(\DLX_IDinst_reg_out_B<2>/GROM )
  );
  X_BUF \DLX_IDinst_reg_out_B<2>/YUSED  (
    .I(\DLX_IDinst_reg_out_B<2>/GROM ),
    .O(DLX_IDinst__n0147[2])
  );
  defparam \DLX_IDinst__n0147<3>1 .INIT = 16'h88A0;
  X_LUT4 \DLX_IDinst__n0147<3>1  (
    .ADR0(DLX_IDinst_N107173),
    .ADR1(DLX_MEMinst_RF_data_in[3]),
    .ADR2(DLX_IDinst__n0623[3]),
    .ADR3(DLX_IDinst__n0176),
    .O(\DLX_IDinst_reg_out_B<3>/GROM )
  );
  X_BUF \DLX_IDinst_reg_out_B<3>/YUSED  (
    .I(\DLX_IDinst_reg_out_B<3>/GROM ),
    .O(DLX_IDinst__n0147[3])
  );
  defparam DLX_IDinst_reg_out_A_10.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_A_10 (
    .I(N162904),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE2573),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_A[10])
  );
  defparam \DLX_IDinst__n0146<10>491 .INIT = 16'h2000;
  X_LUT4 \DLX_IDinst__n0146<10>491  (
    .ADR0(DLX_IDinst_Ker1084541_1),
    .ADR1(DLX_IDinst__n0387),
    .ADR2(DLX_IDinst__n0116),
    .ADR3(DLX_IFinst_NPC[10]),
    .O(N162904)
  );
  defparam \DLX_IDinst__n0146<11>491 .INIT = 16'h0800;
  X_LUT4 \DLX_IDinst__n0146<11>491  (
    .ADR0(DLX_IFinst_NPC[11]),
    .ADR1(DLX_IDinst__n0116),
    .ADR2(DLX_IDinst__n0387),
    .ADR3(DLX_IDinst_Ker1084541_1),
    .O(N162907)
  );
  defparam \DLX_IDinst__n0146<12>491 .INIT = 16'h0800;
  X_LUT4 \DLX_IDinst__n0146<12>491  (
    .ADR0(DLX_IDinst_Ker1084541_1),
    .ADR1(DLX_IFinst_NPC[12]),
    .ADR2(DLX_IDinst__n0387),
    .ADR3(DLX_IDinst__n0116),
    .O(N162910)
  );
  defparam \DLX_IDinst__n0146<20>491 .INIT = 16'h0080;
  X_LUT4 \DLX_IDinst__n0146<20>491  (
    .ADR0(DLX_IDinst__n0116),
    .ADR1(DLX_IDinst_Ker1084541_1),
    .ADR2(DLX_IFinst_NPC[20]),
    .ADR3(DLX_IDinst__n0387),
    .O(N162934)
  );
  defparam \DLX_IDinst__n0146<13>491 .INIT = 16'h4000;
  X_LUT4 \DLX_IDinst__n0146<13>491  (
    .ADR0(DLX_IDinst__n0387),
    .ADR1(DLX_IDinst_Ker1084541_1),
    .ADR2(DLX_IDinst__n0116),
    .ADR3(DLX_IFinst_NPC[13]),
    .O(N162913)
  );
  defparam \DLX_IDinst__n0146<21>491 .INIT = 16'h2000;
  X_LUT4 \DLX_IDinst__n0146<21>491  (
    .ADR0(DLX_IDinst__n0116),
    .ADR1(DLX_IDinst__n0387),
    .ADR2(DLX_IFinst_NPC[21]),
    .ADR3(DLX_IDinst_Ker1084541_1),
    .O(N162937)
  );
  defparam \DLX_IDinst__n0146<14>491 .INIT = 16'h2000;
  X_LUT4 \DLX_IDinst__n0146<14>491  (
    .ADR0(DLX_IDinst__n0116),
    .ADR1(DLX_IDinst__n0387),
    .ADR2(DLX_IDinst_Ker1084541_1),
    .ADR3(DLX_IFinst_NPC[14]),
    .O(N162916)
  );
  defparam \DLX_IDinst__n0146<22>491 .INIT = 16'h4000;
  X_LUT4 \DLX_IDinst__n0146<22>491  (
    .ADR0(DLX_IDinst__n0387),
    .ADR1(DLX_IFinst_NPC[22]),
    .ADR2(DLX_IDinst_Ker1084541_1),
    .ADR3(DLX_IDinst__n0116),
    .O(N162940)
  );
  defparam \DLX_IDinst__n0146<31>661 .INIT = 16'h4000;
  X_LUT4 \DLX_IDinst__n0146<31>661  (
    .ADR0(DLX_IDinst__n0387),
    .ADR1(DLX_IDinst_Ker1084541_1),
    .ADR2(DLX_IFinst_NPC[31]),
    .ADR3(DLX_IDinst__n0116),
    .O(N162871)
  );
  defparam \DLX_IDinst__n0146<15>491 .INIT = 16'h0800;
  X_LUT4 \DLX_IDinst__n0146<15>491  (
    .ADR0(DLX_IDinst__n0116),
    .ADR1(DLX_IDinst_Ker1084541_1),
    .ADR2(DLX_IDinst__n0387),
    .ADR3(DLX_IFinst_NPC[15]),
    .O(N162919)
  );
  defparam \DLX_IDinst__n0146<23>491 .INIT = 16'h4000;
  X_LUT4 \DLX_IDinst__n0146<23>491  (
    .ADR0(DLX_IDinst__n0387),
    .ADR1(DLX_IFinst_NPC[23]),
    .ADR2(DLX_IDinst__n0116),
    .ADR3(DLX_IDinst_Ker1084541_1),
    .O(N162943)
  );
  defparam \DLX_IDinst__n0146<16>491 .INIT = 16'h0080;
  X_LUT4 \DLX_IDinst__n0146<16>491  (
    .ADR0(DLX_IDinst__n0116),
    .ADR1(DLX_IFinst_NPC[16]),
    .ADR2(DLX_IDinst_Ker1084541_1),
    .ADR3(DLX_IDinst__n0387),
    .O(N162922)
  );
  defparam \DLX_IDinst__n0146<24>491 .INIT = 16'h4000;
  X_LUT4 \DLX_IDinst__n0146<24>491  (
    .ADR0(DLX_IDinst__n0387),
    .ADR1(DLX_IDinst_Ker1084541_1),
    .ADR2(DLX_IFinst_NPC[24]),
    .ADR3(DLX_IDinst__n0116),
    .O(N162946)
  );
  defparam \DLX_IDinst__n0146<17>491 .INIT = 16'h2000;
  X_LUT4 \DLX_IDinst__n0146<17>491  (
    .ADR0(DLX_IDinst__n0116),
    .ADR1(DLX_IDinst__n0387),
    .ADR2(DLX_IFinst_NPC[17]),
    .ADR3(DLX_IDinst_Ker1084541_1),
    .O(N162925)
  );
  defparam \DLX_IDinst__n0146<25>491 .INIT = 16'h4000;
  X_LUT4 \DLX_IDinst__n0146<25>491  (
    .ADR0(DLX_IDinst__n0387),
    .ADR1(DLX_IFinst_NPC[25]),
    .ADR2(DLX_IDinst__n0116),
    .ADR3(DLX_IDinst_Ker1084541_1),
    .O(N162949)
  );
  defparam \DLX_IDinst__n0147<31>1 .INIT = 16'h88C0;
  X_LUT4 \DLX_IDinst__n0147<31>1  (
    .ADR0(DLX_MEMinst_RF_data_in[31]),
    .ADR1(DLX_IDinst_N107173),
    .ADR2(DLX_IDinst__n0623[31]),
    .ADR3(DLX_IDinst__n0176),
    .O(DLX_IDinst__n0147[31])
  );
  defparam \DLX_IDinst__n0147<10>1 .INIT = 16'hAC00;
  X_LUT4 \DLX_IDinst__n0147<10>1  (
    .ADR0(DLX_MEMinst_RF_data_in[10]),
    .ADR1(DLX_IDinst__n0623[10]),
    .ADR2(DLX_IDinst__n0176),
    .ADR3(DLX_IDinst_N107173),
    .O(DLX_IDinst__n0147[10])
  );
  defparam \DLX_IDinst__n0146<18>491 .INIT = 16'h0080;
  X_LUT4 \DLX_IDinst__n0146<18>491  (
    .ADR0(DLX_IFinst_NPC[18]),
    .ADR1(DLX_IDinst__n0116),
    .ADR2(DLX_IDinst_Ker1084541_1),
    .ADR3(DLX_IDinst__n0387),
    .O(N162928)
  );
  defparam \DLX_IDinst__n0146<26>491 .INIT = 16'h0800;
  X_LUT4 \DLX_IDinst__n0146<26>491  (
    .ADR0(DLX_IDinst_Ker1084541_1),
    .ADR1(DLX_IDinst__n0116),
    .ADR2(DLX_IDinst__n0387),
    .ADR3(DLX_IFinst_NPC[26]),
    .O(N162952)
  );
  defparam \DLX_IDinst__n0147<30>1 .INIT = 16'h8C80;
  X_LUT4 \DLX_IDinst__n0147<30>1  (
    .ADR0(DLX_MEMinst_RF_data_in[30]),
    .ADR1(DLX_IDinst_N107173),
    .ADR2(DLX_IDinst__n0176),
    .ADR3(DLX_IDinst__n0623[30]),
    .O(DLX_IDinst__n0147[30])
  );
  defparam \DLX_IDinst__n0147<11>1 .INIT = 16'hA0C0;
  X_LUT4 \DLX_IDinst__n0147<11>1  (
    .ADR0(DLX_MEMinst_RF_data_in[11]),
    .ADR1(DLX_IDinst__n0623[11]),
    .ADR2(DLX_IDinst_N107173),
    .ADR3(DLX_IDinst__n0176),
    .O(DLX_IDinst__n0147[11])
  );
  defparam DLX_IDinst_RegFile_22_20_2886.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_22_20_2886 (
    .I(DLX_IDinst_WB_data_eff[20]),
    .CE(DLX_IDinst__n0594),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_22_20)
  );
  defparam \DLX_IDinst__n0146<19>491 .INIT = 16'h4000;
  X_LUT4 \DLX_IDinst__n0146<19>491  (
    .ADR0(DLX_IDinst__n0387),
    .ADR1(DLX_IFinst_NPC[19]),
    .ADR2(DLX_IDinst__n0116),
    .ADR3(DLX_IDinst_Ker1084541_1),
    .O(N162931)
  );
  defparam \DLX_IDinst__n0146<27>491 .INIT = 16'h2000;
  X_LUT4 \DLX_IDinst__n0146<27>491  (
    .ADR0(DLX_IDinst__n0116),
    .ADR1(DLX_IDinst__n0387),
    .ADR2(DLX_IDinst_Ker1084541_1),
    .ADR3(DLX_IFinst_NPC[27]),
    .O(N162955)
  );
  defparam \DLX_IDinst__n0147<29>1 .INIT = 16'hAC00;
  X_LUT4 \DLX_IDinst__n0147<29>1  (
    .ADR0(DLX_MEMinst_RF_data_in[29]),
    .ADR1(DLX_IDinst__n0623[29]),
    .ADR2(DLX_IDinst__n0176),
    .ADR3(DLX_IDinst_N107173),
    .O(DLX_IDinst__n0147[29])
  );
  defparam \DLX_IDinst__n0147<20>1 .INIT = 16'hE400;
  X_LUT4 \DLX_IDinst__n0147<20>1  (
    .ADR0(DLX_IDinst__n0176),
    .ADR1(DLX_IDinst__n0623[20]),
    .ADR2(DLX_MEMinst_RF_data_in[20]),
    .ADR3(DLX_IDinst_N107173),
    .O(DLX_IDinst__n0147[20])
  );
  defparam \DLX_IDinst__n0147<27>1 .INIT = 16'hC808;
  X_LUT4 \DLX_IDinst__n0147<27>1  (
    .ADR0(DLX_IDinst__n0623[27]),
    .ADR1(DLX_IDinst_N107173),
    .ADR2(DLX_IDinst__n0176),
    .ADR3(DLX_MEMinst_RF_data_in[27]),
    .O(DLX_IDinst__n0147[27])
  );
  defparam \DLX_IDinst__n0147<12>1 .INIT = 16'hCA00;
  X_LUT4 \DLX_IDinst__n0147<12>1  (
    .ADR0(DLX_IDinst__n0623[12]),
    .ADR1(DLX_MEMinst_RF_data_in[12]),
    .ADR2(DLX_IDinst__n0176),
    .ADR3(DLX_IDinst_N107173),
    .O(DLX_IDinst__n0147[12])
  );
  defparam \DLX_IDinst__n0146<28>491 .INIT = 16'h0800;
  X_LUT4 \DLX_IDinst__n0146<28>491  (
    .ADR0(DLX_IDinst_Ker1084541_1),
    .ADR1(DLX_IDinst__n0116),
    .ADR2(DLX_IDinst__n0387),
    .ADR3(DLX_IFinst_NPC[28]),
    .O(N162958)
  );
  defparam \DLX_IDinst__n0147<26>1 .INIT = 16'hC0A0;
  X_LUT4 \DLX_IDinst__n0147<26>1  (
    .ADR0(DLX_IDinst__n0623[26]),
    .ADR1(DLX_MEMinst_RF_data_in[26]),
    .ADR2(DLX_IDinst_N107173),
    .ADR3(DLX_IDinst__n0176),
    .O(DLX_IDinst__n0147[26])
  );
  defparam \DLX_IDinst__n0147<21>1 .INIT = 16'hA088;
  X_LUT4 \DLX_IDinst__n0147<21>1  (
    .ADR0(DLX_IDinst_N107173),
    .ADR1(DLX_IDinst__n0623[21]),
    .ADR2(DLX_MEMinst_RF_data_in[21]),
    .ADR3(DLX_IDinst__n0176),
    .O(DLX_IDinst__n0147[21])
  );
  defparam \DLX_IDinst__n0147<25>1 .INIT = 16'hB800;
  X_LUT4 \DLX_IDinst__n0147<25>1  (
    .ADR0(DLX_MEMinst_RF_data_in[25]),
    .ADR1(DLX_IDinst__n0176),
    .ADR2(DLX_IDinst__n0623[25]),
    .ADR3(DLX_IDinst_N107173),
    .O(DLX_IDinst__n0147[25])
  );
  defparam \DLX_IDinst__n0147<13>1 .INIT = 16'hCA00;
  X_LUT4 \DLX_IDinst__n0147<13>1  (
    .ADR0(DLX_IDinst__n0623[13]),
    .ADR1(DLX_MEMinst_RF_data_in[13]),
    .ADR2(DLX_IDinst__n0176),
    .ADR3(DLX_IDinst_N107173),
    .O(DLX_IDinst__n0147[13])
  );
  defparam \DLX_IDinst__n0146<29>491 .INIT = 16'h0080;
  X_LUT4 \DLX_IDinst__n0146<29>491  (
    .ADR0(DLX_IFinst_NPC[29]),
    .ADR1(DLX_IDinst__n0116),
    .ADR2(DLX_IDinst_Ker1084541_1),
    .ADR3(DLX_IDinst__n0387),
    .O(N162961)
  );
  defparam \DLX_IDinst__n0147<24>1 .INIT = 16'hA280;
  X_LUT4 \DLX_IDinst__n0147<24>1  (
    .ADR0(DLX_IDinst_N107173),
    .ADR1(DLX_IDinst__n0176),
    .ADR2(DLX_MEMinst_RF_data_in[24]),
    .ADR3(DLX_IDinst__n0623[24]),
    .O(DLX_IDinst__n0147[24])
  );
  defparam \DLX_IDinst__n0147<22>1 .INIT = 16'hB080;
  X_LUT4 \DLX_IDinst__n0147<22>1  (
    .ADR0(DLX_MEMinst_RF_data_in[22]),
    .ADR1(DLX_IDinst__n0176),
    .ADR2(DLX_IDinst_N107173),
    .ADR3(DLX_IDinst__n0623[22]),
    .O(DLX_IDinst__n0147[22])
  );
  defparam \DLX_IDinst__n0147<23>1 .INIT = 16'hC840;
  X_LUT4 \DLX_IDinst__n0147<23>1  (
    .ADR0(DLX_IDinst__n0176),
    .ADR1(DLX_IDinst_N107173),
    .ADR2(DLX_IDinst__n0623[23]),
    .ADR3(DLX_MEMinst_RF_data_in[23]),
    .O(DLX_IDinst__n0147[23])
  );
  defparam \DLX_IDinst__n0147<14>1 .INIT = 16'hAC00;
  X_LUT4 \DLX_IDinst__n0147<14>1  (
    .ADR0(DLX_MEMinst_RF_data_in[14]),
    .ADR1(DLX_IDinst__n0623[14]),
    .ADR2(DLX_IDinst__n0176),
    .ADR3(DLX_IDinst_N107173),
    .O(DLX_IDinst__n0147[14])
  );
  defparam \DLX_IDinst__n0147<19>1 .INIT = 16'hA820;
  X_LUT4 \DLX_IDinst__n0147<19>1  (
    .ADR0(DLX_IDinst_N107173),
    .ADR1(DLX_IDinst__n0176),
    .ADR2(DLX_IDinst__n0623[19]),
    .ADR3(DLX_MEMinst_RF_data_in[19]),
    .O(DLX_IDinst__n0147[19])
  );
  defparam \DLX_IDinst__n0147<15>1 .INIT = 16'hC088;
  X_LUT4 \DLX_IDinst__n0147<15>1  (
    .ADR0(DLX_IDinst__n0623[15]),
    .ADR1(DLX_IDinst_N107173),
    .ADR2(DLX_MEMinst_RF_data_in[15]),
    .ADR3(DLX_IDinst__n0176),
    .O(DLX_IDinst__n0147[15])
  );
  defparam \DLX_IDinst__n0147<18>1 .INIT = 16'hD800;
  X_LUT4 \DLX_IDinst__n0147<18>1  (
    .ADR0(DLX_IDinst__n0176),
    .ADR1(DLX_MEMinst_RF_data_in[18]),
    .ADR2(DLX_IDinst__n0623[18]),
    .ADR3(DLX_IDinst_N107173),
    .O(DLX_IDinst__n0147[18])
  );
  defparam \DLX_IDinst__n0147<16>1 .INIT = 16'hE200;
  X_LUT4 \DLX_IDinst__n0147<16>1  (
    .ADR0(DLX_IDinst__n0623[16]),
    .ADR1(DLX_IDinst__n0176),
    .ADR2(DLX_MEMinst_RF_data_in[16]),
    .ADR3(DLX_IDinst_N107173),
    .O(DLX_IDinst__n0147[16])
  );
  defparam \DLX_IDinst__n0147<9>1 .INIT = 16'hC840;
  X_LUT4 \DLX_IDinst__n0147<9>1  (
    .ADR0(DLX_IDinst__n0176),
    .ADR1(DLX_IDinst_N107173),
    .ADR2(DLX_IDinst__n0623[9]),
    .ADR3(DLX_MEMinst_RF_data_in[9]),
    .O(DLX_IDinst__n0147[9])
  );
  defparam \DLX_IDinst__n0147<17>1 .INIT = 16'hA088;
  X_LUT4 \DLX_IDinst__n0147<17>1  (
    .ADR0(DLX_IDinst_N107173),
    .ADR1(DLX_IDinst__n0623[17]),
    .ADR2(DLX_MEMinst_RF_data_in[17]),
    .ADR3(DLX_IDinst__n0176),
    .O(DLX_IDinst__n0147[17])
  );
  defparam \DLX_IDinst__n0146<0>661 .INIT = 16'h0080;
  X_LUT4 \DLX_IDinst__n0146<0>661  (
    .ADR0(DLX_IDinst__n0116),
    .ADR1(DLX_IDinst_Ker1084541_1),
    .ADR2(DLX_IFinst_NPC[0]),
    .ADR3(DLX_IDinst__n0387),
    .O(N162874)
  );
  defparam \DLX_IDinst__n0146<1>491 .INIT = 16'h4000;
  X_LUT4 \DLX_IDinst__n0146<1>491  (
    .ADR0(DLX_IDinst__n0387),
    .ADR1(DLX_IDinst__n0116),
    .ADR2(DLX_IDinst_Ker1084541_1),
    .ADR3(DLX_IFinst_NPC[1]),
    .O(N162877)
  );
  defparam \DLX_IDinst__n0146<2>491 .INIT = 16'h0800;
  X_LUT4 \DLX_IDinst__n0146<2>491  (
    .ADR0(DLX_IDinst_Ker1084541_1),
    .ADR1(DLX_IFinst_NPC[2]),
    .ADR2(DLX_IDinst__n0387),
    .ADR3(DLX_IDinst__n0116),
    .O(N162880)
  );
  defparam \DLX_IDinst__n0146<3>491 .INIT = 16'h0080;
  X_LUT4 \DLX_IDinst__n0146<3>491  (
    .ADR0(DLX_IDinst_Ker1084541_1),
    .ADR1(DLX_IFinst_NPC[3]),
    .ADR2(DLX_IDinst__n0116),
    .ADR3(DLX_IDinst__n0387),
    .O(N162883)
  );
  defparam \DLX_IDinst__n0146<4>491 .INIT = 16'h0800;
  X_LUT4 \DLX_IDinst__n0146<4>491  (
    .ADR0(DLX_IDinst__n0116),
    .ADR1(DLX_IFinst_NPC[4]),
    .ADR2(DLX_IDinst__n0387),
    .ADR3(DLX_IDinst_Ker1084541_1),
    .O(N162886)
  );
  defparam \DLX_IDinst__n0147<8>1 .INIT = 16'h8C80;
  X_LUT4 \DLX_IDinst__n0147<8>1  (
    .ADR0(DLX_MEMinst_RF_data_in[8]),
    .ADR1(DLX_IDinst_N107173),
    .ADR2(DLX_IDinst__n0176),
    .ADR3(DLX_IDinst__n0623[8]),
    .O(DLX_IDinst__n0147[8])
  );
  defparam \DLX_IDinst__n0147<1>1 .INIT = 16'hC088;
  X_LUT4 \DLX_IDinst__n0147<1>1  (
    .ADR0(DLX_IDinst__n0623[1]),
    .ADR1(DLX_IDinst_N107173),
    .ADR2(DLX_MEMinst_RF_data_in[1]),
    .ADR3(DLX_IDinst__n0176),
    .O(DLX_IDinst__n0147[1])
  );
  defparam \DLX_IDinst__n0146<5>491 .INIT = 16'h2000;
  X_LUT4 \DLX_IDinst__n0146<5>491  (
    .ADR0(DLX_IFinst_NPC[5]),
    .ADR1(DLX_IDinst__n0387),
    .ADR2(DLX_IDinst_Ker1084541_1),
    .ADR3(DLX_IDinst__n0116),
    .O(N162889)
  );
  defparam \DLX_IDinst__n0146<6>661 .INIT = 16'h4000;
  X_LUT4 \DLX_IDinst__n0146<6>661  (
    .ADR0(DLX_IDinst__n0387),
    .ADR1(DLX_IFinst_NPC[6]),
    .ADR2(DLX_IDinst__n0116),
    .ADR3(DLX_IDinst_Ker1084541_1),
    .O(N162892)
  );
  defparam \DLX_IDinst__n0146<7>491 .INIT = 16'h2000;
  X_LUT4 \DLX_IDinst__n0146<7>491  (
    .ADR0(DLX_IDinst__n0116),
    .ADR1(DLX_IDinst__n0387),
    .ADR2(DLX_IFinst_NPC[7]),
    .ADR3(DLX_IDinst_Ker1084541_1),
    .O(N162895)
  );
  defparam \DLX_IDinst__n0147<7>1 .INIT = 16'hE400;
  X_LUT4 \DLX_IDinst__n0147<7>1  (
    .ADR0(DLX_IDinst__n0176),
    .ADR1(DLX_IDinst__n0623[7]),
    .ADR2(DLX_MEMinst_RF_data_in[7]),
    .ADR3(DLX_IDinst_N107173),
    .O(DLX_IDinst__n0147[7])
  );
  defparam \DLX_IDinst__n0147<4>1 .INIT = 16'hE400;
  X_LUT4 \DLX_IDinst__n0147<4>1  (
    .ADR0(DLX_IDinst__n0176),
    .ADR1(DLX_IDinst__n0623[4]),
    .ADR2(DLX_MEMinst_RF_data_in[4]),
    .ADR3(DLX_IDinst_N107173),
    .O(DLX_IDinst__n0147[4])
  );
  defparam \DLX_IDinst__n0146<8>491 .INIT = 16'h2000;
  X_LUT4 \DLX_IDinst__n0146<8>491  (
    .ADR0(DLX_IDinst__n0116),
    .ADR1(DLX_IDinst__n0387),
    .ADR2(DLX_IDinst_Ker1084541_1),
    .ADR3(DLX_IFinst_NPC[8]),
    .O(N162898)
  );
  defparam \DLX_IDinst__n0147<6>1 .INIT = 16'hC840;
  X_LUT4 \DLX_IDinst__n0147<6>1  (
    .ADR0(DLX_IDinst__n0176),
    .ADR1(DLX_IDinst_N107173),
    .ADR2(DLX_IDinst__n0623[6]),
    .ADR3(DLX_MEMinst_RF_data_in[6]),
    .O(DLX_IDinst__n0147[6])
  );
  defparam \DLX_IDinst__n0147<5>1 .INIT = 16'h88C0;
  X_LUT4 \DLX_IDinst__n0147<5>1  (
    .ADR0(DLX_MEMinst_RF_data_in[5]),
    .ADR1(DLX_IDinst_N107173),
    .ADR2(DLX_IDinst__n0623[5]),
    .ADR3(DLX_IDinst__n0176),
    .O(DLX_IDinst__n0147[5])
  );
  defparam DLX_IDinst_IR_opcode_field_1.INIT = 1'b0;
  X_SFF DLX_IDinst_IR_opcode_field_1 (
    .I(DLX_IDinst__n0142[1]),
    .CE(DLX_IDinst__n0116),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_IDinst__n0115),
    .O(DLX_IDinst_IR_opcode_field[1])
  );
  defparam \DLX_IDinst__n0146<9>491 .INIT = 16'h0800;
  X_LUT4 \DLX_IDinst__n0146<9>491  (
    .ADR0(DLX_IFinst_NPC[9]),
    .ADR1(DLX_IDinst__n0116),
    .ADR2(DLX_IDinst__n0387),
    .ADR3(DLX_IDinst_Ker1084541_1),
    .O(N162901)
  );
  defparam \DLX_EXinst_Mmux_reg_dst_of_EX_Result<0>1 .INIT = 16'hF0AA;
  X_LUT4 \DLX_EXinst_Mmux_reg_dst_of_EX_Result<0>1  (
    .ADR0(DLX_IDinst_rt_addr[0]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_rd_addr[0]),
    .ADR3(DLX_IDinst_reg_dst),
    .O(\DLX_EXinst_reg_dst_out<0>/GROM )
  );
  X_BUF \DLX_EXinst_reg_dst_out<0>/YUSED  (
    .I(\DLX_EXinst_reg_dst_out<0>/GROM ),
    .O(DLX_reg_dst_of_EX[0])
  );
  defparam \DLX_EXinst_Mmux_reg_dst_of_EX_Result<1>1 .INIT = 16'hDD88;
  X_LUT4 \DLX_EXinst_Mmux_reg_dst_of_EX_Result<1>1  (
    .ADR0(DLX_IDinst_reg_dst),
    .ADR1(DLX_IDinst_rd_addr[1]),
    .ADR2(VCC),
    .ADR3(DLX_IDinst_rt_addr[1]),
    .O(\DLX_EXinst_reg_dst_out<1>/GROM )
  );
  X_BUF \DLX_EXinst_reg_dst_out<1>/YUSED  (
    .I(\DLX_EXinst_reg_dst_out<1>/GROM ),
    .O(DLX_reg_dst_of_EX[1])
  );
  defparam \DLX_EXinst_Mmux_reg_dst_of_EX_Result<2>1 .INIT = 16'hCFC0;
  X_LUT4 \DLX_EXinst_Mmux_reg_dst_of_EX_Result<2>1  (
    .ADR0(VCC),
    .ADR1(DLX_IDinst_rd_addr[2]),
    .ADR2(DLX_IDinst_reg_dst),
    .ADR3(DLX_IDinst_rt_addr[2]),
    .O(\DLX_EXinst_reg_dst_out<2>/GROM )
  );
  X_BUF \DLX_EXinst_reg_dst_out<2>/YUSED  (
    .I(\DLX_EXinst_reg_dst_out<2>/GROM ),
    .O(DLX_reg_dst_of_EX[2])
  );
  defparam \DLX_EXinst_Mmux_reg_dst_of_EX_Result<3>1 .INIT = 16'hF5A0;
  X_LUT4 \DLX_EXinst_Mmux_reg_dst_of_EX_Result<3>1  (
    .ADR0(DLX_IDinst_reg_dst),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_rd_addr[3]),
    .ADR3(DLX_IDinst_rt_addr[3]),
    .O(\DLX_EXinst_reg_dst_out<3>/GROM )
  );
  X_BUF \DLX_EXinst_reg_dst_out<3>/YUSED  (
    .I(\DLX_EXinst_reg_dst_out<3>/GROM ),
    .O(DLX_reg_dst_of_EX[3])
  );
  X_ZERO \DLX_EXinst_reg_dst_out<4>/LOGIC_ZERO_2887  (
    .O(\DLX_EXinst_reg_dst_out<4>/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mcompar__n0100_inst_cy_264 (
    .IA(\DLX_EXinst_reg_dst_out<4>/LOGIC_ZERO ),
    .IB(\DLX_EXinst_reg_dst_out<4>/CYINIT ),
    .SEL(DLX_IDinst_Mcompar__n0100_inst_lut4_42),
    .O(\DLX_EXinst_reg_dst_out<4>/CYMUXF )
  );
  defparam DLX_IDinst_Mcompar__n0100_inst_lut4_421.INIT = 16'hD287;
  X_LUT4 DLX_IDinst_Mcompar__n0100_inst_lut4_421 (
    .ADR0(DLX_EXinst__n0144),
    .ADR1(DLX_IFinst_IR_latched[25]),
    .ADR2(DLX_reg_dst_of_EX[4]),
    .ADR3(DLX_IDinst_current_IR[25]),
    .O(DLX_IDinst_Mcompar__n0100_inst_lut4_42)
  );
  defparam \DLX_EXinst_Mmux_reg_dst_of_EX_Result<4>1 .INIT = 16'hFA0A;
  X_LUT4 \DLX_EXinst_Mmux_reg_dst_of_EX_Result<4>1  (
    .ADR0(DLX_IDinst_rt_addr[4]),
    .ADR1(VCC),
    .ADR2(DLX_IDinst_reg_dst),
    .ADR3(DLX_IDinst_rd_addr[4]),
    .O(\DLX_EXinst_reg_dst_out<4>/GROM )
  );
  X_BUF \DLX_EXinst_reg_dst_out<4>/XBUSED  (
    .I(\DLX_EXinst_reg_dst_out<4>/CYMUXF ),
    .O(DLX_IDinst__n0100)
  );
  X_BUF \DLX_EXinst_reg_dst_out<4>/YUSED  (
    .I(\DLX_EXinst_reg_dst_out<4>/GROM ),
    .O(DLX_reg_dst_of_EX[4])
  );
  X_BUF \DLX_EXinst_reg_dst_out<4>/CYINIT_2888  (
    .I(DLX_IDinst_Mcompar__n0100_inst_cy_263),
    .O(\DLX_EXinst_reg_dst_out<4>/CYINIT )
  );
  defparam \DLX_EXinst_Mshift__n0023_Sh<2> .INIT = 16'h2075;
  X_LUT4 \DLX_EXinst_Mshift__n0023_Sh<2>  (
    .ADR0(DLX_IDinst_reg_out_B[1]),
    .ADR1(DLX_IDinst_reg_out_B[0]),
    .ADR2(DLX_IDinst_reg_out_A[0]),
    .ADR3(N131631),
    .O(\DLX_EXinst_reg_out_B_EX<6>/FROM )
  );
  defparam \DLX_EXinst__n0007<18>367_SW0 .INIT = 16'hF4F0;
  X_LUT4 \DLX_EXinst__n0007<18>367_SW0  (
    .ADR0(DLX_EXinst_N72822),
    .ADR1(DLX_EXinst_N75973),
    .ADR2(CHOICE5266),
    .ADR3(\DLX_EXinst_Mshift__n0023_Sh[2] ),
    .O(\DLX_EXinst_reg_out_B_EX<6>/GROM )
  );
  X_BUF \DLX_EXinst_reg_out_B_EX<6>/XUSED  (
    .I(\DLX_EXinst_reg_out_B_EX<6>/FROM ),
    .O(\DLX_EXinst_Mshift__n0023_Sh[2] )
  );
  X_BUF \DLX_EXinst_reg_out_B_EX<6>/YUSED  (
    .I(\DLX_EXinst_reg_out_B_EX<6>/GROM ),
    .O(N163290)
  );
  defparam DLX_IDinst_Imm_0_1_2889.INIT = 1'b0;
  X_SFF DLX_IDinst_Imm_0_1_2889 (
    .I(\DLX_IDinst_Imm<0>/GROM ),
    .CE(DLX_IDinst__n0116),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_IDinst__n0115),
    .O(DLX_IDinst_Imm_0_1)
  );
  defparam DLX_IDinst_IR_opcode_field_3.INIT = 1'b0;
  X_SFF DLX_IDinst_IR_opcode_field_3 (
    .I(DLX_IDinst__n0142[3]),
    .CE(DLX_IDinst__n0116),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_IDinst__n0115),
    .O(DLX_IDinst_IR_opcode_field[3])
  );
  X_ZERO \DLX_IDinst_RegFile_12_10/LOGIC_ZERO_2890  (
    .O(\DLX_IDinst_RegFile_12_10/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_166_2891 (
    .IA(\DLX_IDinst_RegFile_12_10/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_12_10/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_225),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_166)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2251.INIT = 16'hB8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2251 (
    .ADR0(DLX_IDinst_RegFile_13_10),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR2(DLX_IDinst_RegFile_12_10),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_49),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_225)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2261.INIT = 16'hB8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2261 (
    .ADR0(DLX_IDinst_RegFile_15_10),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR2(DLX_IDinst_RegFile_14_10),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_50),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_226)
  );
  X_BUF \DLX_IDinst_RegFile_12_10/COUTUSED  (
    .I(\DLX_IDinst_RegFile_12_10/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_167)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_167_2892 (
    .IA(\DLX_IDinst_RegFile_12_10/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_166),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_226),
    .O(\DLX_IDinst_RegFile_12_10/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_12_10/CYINIT_2893  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_165),
    .O(\DLX_IDinst_RegFile_12_10/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_20_10/LOGIC_ZERO_2894  (
    .O(\DLX_IDinst_RegFile_20_10/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_170_2895 (
    .IA(\DLX_IDinst_RegFile_20_10/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_20_10/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_229),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_170)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2291.INIT = 16'hF7B3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2291 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_53),
    .ADR2(DLX_IDinst_RegFile_21_10),
    .ADR3(DLX_IDinst_RegFile_20_10),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_229)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2301.INIT = 16'hF7D5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2301 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_54),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR2(DLX_IDinst_RegFile_23_10),
    .ADR3(DLX_IDinst_RegFile_22_10),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_230)
  );
  X_BUF \DLX_IDinst_RegFile_20_10/COUTUSED  (
    .I(\DLX_IDinst_RegFile_20_10/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_171)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_171_2896 (
    .IA(\DLX_IDinst_RegFile_20_10/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_170),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_230),
    .O(\DLX_IDinst_RegFile_20_10/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_20_10/CYINIT_2897  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_169),
    .O(\DLX_IDinst_RegFile_20_10/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_12_11/LOGIC_ZERO_2898  (
    .O(\DLX_IDinst_RegFile_12_11/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_182_2899 (
    .IA(\DLX_IDinst_RegFile_12_11/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_12_11/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_241),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_182)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2411.INIT = 16'hDF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2411 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR1(DLX_IDinst_RegFile_13_11),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_49),
    .ADR3(DLX_IDinst_RegFile_12_11),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_241)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2421.INIT = 16'hAFCF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2421 (
    .ADR0(DLX_IDinst_RegFile_15_11),
    .ADR1(DLX_IDinst_RegFile_14_11),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_50),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_242)
  );
  X_BUF \DLX_IDinst_RegFile_12_11/COUTUSED  (
    .I(\DLX_IDinst_RegFile_12_11/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_183)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_183_2900 (
    .IA(\DLX_IDinst_RegFile_12_11/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_182),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_242),
    .O(\DLX_IDinst_RegFile_12_11/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_12_11/CYINIT_2901  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_181),
    .O(\DLX_IDinst_RegFile_12_11/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_20_11/LOGIC_ZERO_2902  (
    .O(\DLX_IDinst_RegFile_20_11/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_186_2903 (
    .IA(\DLX_IDinst_RegFile_20_11/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_20_11/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_245),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_186)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2451.INIT = 16'hFB3B;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2451 (
    .ADR0(DLX_IDinst_RegFile_20_11),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_53),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR3(DLX_IDinst_RegFile_21_11),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_245)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2461.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2461 (
    .ADR0(DLX_IDinst_RegFile_23_11),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_54),
    .ADR2(DLX_IDinst_RegFile_22_11),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_246)
  );
  X_BUF \DLX_IDinst_RegFile_20_11/COUTUSED  (
    .I(\DLX_IDinst_RegFile_20_11/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_187)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_187_2904 (
    .IA(\DLX_IDinst_RegFile_20_11/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_186),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_246),
    .O(\DLX_IDinst_RegFile_20_11/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_20_11/CYINIT_2905  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_185),
    .O(\DLX_IDinst_RegFile_20_11/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_12_20/LOGIC_ZERO_2906  (
    .O(\DLX_IDinst_RegFile_12_20/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_326_2907 (
    .IA(\DLX_IDinst_RegFile_12_20/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_12_20/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_385),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_326)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3851.INIT = 16'hB8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3851 (
    .ADR0(DLX_IDinst_RegFile_13_20),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR2(DLX_IDinst_RegFile_12_20),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_49),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_385)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3861.INIT = 16'hAFCF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3861 (
    .ADR0(DLX_IDinst_RegFile_15_20),
    .ADR1(DLX_IDinst_RegFile_14_20),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_50),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_386)
  );
  X_BUF \DLX_IDinst_RegFile_12_20/COUTUSED  (
    .I(\DLX_IDinst_RegFile_12_20/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_327)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_327_2908 (
    .IA(\DLX_IDinst_RegFile_12_20/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_326),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_386),
    .O(\DLX_IDinst_RegFile_12_20/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_12_20/CYINIT_2909  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_325),
    .O(\DLX_IDinst_RegFile_12_20/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_12_12/LOGIC_ZERO_2910  (
    .O(\DLX_IDinst_RegFile_12_12/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_198_2911 (
    .IA(\DLX_IDinst_RegFile_12_12/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_12_12/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_257),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_198)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2571.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2571 (
    .ADR0(DLX_IDinst_RegFile_13_12),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_49),
    .ADR2(DLX_IDinst_RegFile_12_12),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_257)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2581.INIT = 16'hE4FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2581 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR1(DLX_IDinst_RegFile_14_12),
    .ADR2(DLX_IDinst_RegFile_15_12),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_50),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_258)
  );
  X_BUF \DLX_IDinst_RegFile_12_12/COUTUSED  (
    .I(\DLX_IDinst_RegFile_12_12/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_199)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_199_2912 (
    .IA(\DLX_IDinst_RegFile_12_12/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_198),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_258),
    .O(\DLX_IDinst_RegFile_12_12/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_12_12/CYINIT_2913  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_197),
    .O(\DLX_IDinst_RegFile_12_12/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_20_20/LOGIC_ZERO_2914  (
    .O(\DLX_IDinst_RegFile_20_20/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_330_2915 (
    .IA(\DLX_IDinst_RegFile_20_20/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_20_20/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_389),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_330)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3891.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3891 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_53),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR2(DLX_IDinst_RegFile_20_20),
    .ADR3(DLX_IDinst_RegFile_21_20),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_389)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3901.INIT = 16'hDFD5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3901 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_54),
    .ADR1(DLX_IDinst_RegFile_23_20),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR3(DLX_IDinst_RegFile_22_20),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_390)
  );
  X_BUF \DLX_IDinst_RegFile_20_20/COUTUSED  (
    .I(\DLX_IDinst_RegFile_20_20/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_331)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_331_2916 (
    .IA(\DLX_IDinst_RegFile_20_20/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_330),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_390),
    .O(\DLX_IDinst_RegFile_20_20/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_20_20/CYINIT_2917  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_329),
    .O(\DLX_IDinst_RegFile_20_20/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_20_12/LOGIC_ZERO_2918  (
    .O(\DLX_IDinst_RegFile_20_12/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_202_2919 (
    .IA(\DLX_IDinst_RegFile_20_12/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_20_12/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_261),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_202)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2611.INIT = 16'hBF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2611 (
    .ADR0(DLX_IDinst_RegFile_21_12),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_53),
    .ADR3(DLX_IDinst_RegFile_20_12),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_261)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2621.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2621 (
    .ADR0(DLX_IDinst_RegFile_22_12),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_54),
    .ADR2(DLX_IDinst_RegFile_23_12),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_5 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_262)
  );
  X_BUF \DLX_IDinst_RegFile_20_12/COUTUSED  (
    .I(\DLX_IDinst_RegFile_20_12/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_203)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_203_2920 (
    .IA(\DLX_IDinst_RegFile_20_12/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_202),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_262),
    .O(\DLX_IDinst_RegFile_20_12/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_20_12/CYINIT_2921  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_201),
    .O(\DLX_IDinst_RegFile_20_12/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_12_21/LOGIC_ZERO_2922  (
    .O(\DLX_IDinst_RegFile_12_21/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_342_2923 (
    .IA(\DLX_IDinst_RegFile_12_21/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_12_21/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_401),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_342)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4011.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4011 (
    .ADR0(DLX_IDinst_RegFile_12_21),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_49),
    .ADR3(DLX_IDinst_RegFile_13_21),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_401)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4021.INIT = 16'hE2FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4021 (
    .ADR0(DLX_IDinst_RegFile_14_21),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR2(DLX_IDinst_RegFile_15_21),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_50),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_402)
  );
  X_BUF \DLX_IDinst_RegFile_12_21/COUTUSED  (
    .I(\DLX_IDinst_RegFile_12_21/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_343)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_343_2924 (
    .IA(\DLX_IDinst_RegFile_12_21/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_342),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_402),
    .O(\DLX_IDinst_RegFile_12_21/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_12_21/CYINIT_2925  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_341),
    .O(\DLX_IDinst_RegFile_12_21/CYINIT )
  );
  defparam DLX_IDinst_IR_opcode_field_4.INIT = 1'b0;
  X_SFF DLX_IDinst_IR_opcode_field_4 (
    .I(DLX_IDinst__n0142[4]),
    .CE(DLX_IDinst__n0116),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_IDinst__n0115),
    .O(DLX_IDinst_IR_opcode_field[4])
  );
  X_ZERO \DLX_IDinst_RegFile_12_13/LOGIC_ZERO_2926  (
    .O(\DLX_IDinst_RegFile_12_13/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_214_2927 (
    .IA(\DLX_IDinst_RegFile_12_13/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_12_13/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_273),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_214)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2731.INIT = 16'hFD5D;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2731 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_49),
    .ADR1(DLX_IDinst_RegFile_12_13),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR3(DLX_IDinst_RegFile_13_13),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_273)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2741.INIT = 16'hCFAF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2741 (
    .ADR0(DLX_IDinst_RegFile_14_13),
    .ADR1(DLX_IDinst_RegFile_15_13),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_50),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_274)
  );
  X_BUF \DLX_IDinst_RegFile_12_13/COUTUSED  (
    .I(\DLX_IDinst_RegFile_12_13/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_215)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_215_2928 (
    .IA(\DLX_IDinst_RegFile_12_13/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_214),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_274),
    .O(\DLX_IDinst_RegFile_12_13/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_12_13/CYINIT_2929  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_213),
    .O(\DLX_IDinst_RegFile_12_13/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_20_21/LOGIC_ZERO_2930  (
    .O(\DLX_IDinst_RegFile_20_21/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_346_2931 (
    .IA(\DLX_IDinst_RegFile_20_21/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_20_21/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_405),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_346)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4051.INIT = 16'hFB3B;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4051 (
    .ADR0(DLX_IDinst_RegFile_20_21),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_53),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR3(DLX_IDinst_RegFile_21_21),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_405)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4061.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4061 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR1(DLX_IDinst_RegFile_22_21),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_54),
    .ADR3(DLX_IDinst_RegFile_23_21),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_406)
  );
  X_BUF \DLX_IDinst_RegFile_20_21/COUTUSED  (
    .I(\DLX_IDinst_RegFile_20_21/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_347)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_347_2932 (
    .IA(\DLX_IDinst_RegFile_20_21/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_346),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_406),
    .O(\DLX_IDinst_RegFile_20_21/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_20_21/CYINIT_2933  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_345),
    .O(\DLX_IDinst_RegFile_20_21/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_20_13/LOGIC_ZERO_2934  (
    .O(\DLX_IDinst_RegFile_20_13/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_218_2935 (
    .IA(\DLX_IDinst_RegFile_20_13/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_20_13/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_277),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_218)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2771.INIT = 16'hFB73;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2771 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_53),
    .ADR2(DLX_IDinst_RegFile_20_13),
    .ADR3(DLX_IDinst_RegFile_21_13),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_277)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2781.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2781 (
    .ADR0(DLX_IDinst_RegFile_22_13),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_54),
    .ADR2(DLX_IDinst_RegFile_23_13),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_278)
  );
  X_BUF \DLX_IDinst_RegFile_20_13/COUTUSED  (
    .I(\DLX_IDinst_RegFile_20_13/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_219)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_219_2936 (
    .IA(\DLX_IDinst_RegFile_20_13/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_218),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_278),
    .O(\DLX_IDinst_RegFile_20_13/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_20_13/CYINIT_2937  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_217),
    .O(\DLX_IDinst_RegFile_20_13/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_12_30/LOGIC_ZERO_2938  (
    .O(\DLX_IDinst_RegFile_12_30/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_998_2939 (
    .IA(\DLX_IDinst_RegFile_12_30/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_12_30/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1073),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_998)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10731.INIT = 16'hFB73;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10731 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_577),
    .ADR2(DLX_IDinst_RegFile_12_30),
    .ADR3(DLX_IDinst_RegFile_13_30),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1073)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10741.INIT = 16'hAFCF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10741 (
    .ADR0(DLX_IDinst_RegFile_15_30),
    .ADR1(DLX_IDinst_RegFile_14_30),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_578),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1074)
  );
  X_BUF \DLX_IDinst_RegFile_12_30/COUTUSED  (
    .I(\DLX_IDinst_RegFile_12_30/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_999)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_999_2940 (
    .IA(\DLX_IDinst_RegFile_12_30/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_998),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1074),
    .O(\DLX_IDinst_RegFile_12_30/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_12_30/CYINIT_2941  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_997),
    .O(\DLX_IDinst_RegFile_12_30/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_12_22/LOGIC_ZERO_2942  (
    .O(\DLX_IDinst_RegFile_12_22/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_358_2943 (
    .IA(\DLX_IDinst_RegFile_12_22/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_12_22/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_417),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_358)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4171.INIT = 16'hFD5D;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4171 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_49),
    .ADR1(DLX_IDinst_RegFile_12_22),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR3(DLX_IDinst_RegFile_13_22),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_417)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4181.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4181 (
    .ADR0(DLX_IDinst_RegFile_14_22),
    .ADR1(DLX_IDinst_RegFile_15_22),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_50),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_418)
  );
  X_BUF \DLX_IDinst_RegFile_12_22/COUTUSED  (
    .I(\DLX_IDinst_RegFile_12_22/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_359)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_359_2944 (
    .IA(\DLX_IDinst_RegFile_12_22/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_358),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_418),
    .O(\DLX_IDinst_RegFile_12_22/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_12_22/CYINIT_2945  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_357),
    .O(\DLX_IDinst_RegFile_12_22/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_12_14/LOGIC_ZERO_2946  (
    .O(\DLX_IDinst_RegFile_12_14/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_230_2947 (
    .IA(\DLX_IDinst_RegFile_12_14/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_12_14/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_289),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_230)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2891.INIT = 16'hDDF5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2891 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_49),
    .ADR1(DLX_IDinst_RegFile_13_14),
    .ADR2(DLX_IDinst_RegFile_12_14),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_289)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2901.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2901 (
    .ADR0(DLX_IDinst_RegFile_15_14),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_50),
    .ADR2(DLX_IDinst_RegFile_14_14),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_290)
  );
  X_BUF \DLX_IDinst_RegFile_12_14/COUTUSED  (
    .I(\DLX_IDinst_RegFile_12_14/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_231)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_231_2948 (
    .IA(\DLX_IDinst_RegFile_12_14/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_230),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_290),
    .O(\DLX_IDinst_RegFile_12_14/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_12_14/CYINIT_2949  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_229),
    .O(\DLX_IDinst_RegFile_12_14/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_20_30/LOGIC_ZERO_2950  (
    .O(\DLX_IDinst_RegFile_20_30/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_1002_2951 (
    .IA(\DLX_IDinst_RegFile_20_30/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_20_30/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1077),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_1002)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10771.INIT = 16'hACFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10771 (
    .ADR0(DLX_IDinst_RegFile_21_30),
    .ADR1(DLX_IDinst_RegFile_20_30),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_581),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1077)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10781.INIT = 16'hCFAF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10781 (
    .ADR0(DLX_IDinst_RegFile_22_30),
    .ADR1(DLX_IDinst_RegFile_23_30),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_582),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1078)
  );
  X_BUF \DLX_IDinst_RegFile_20_30/COUTUSED  (
    .I(\DLX_IDinst_RegFile_20_30/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_1003)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_1003_2952 (
    .IA(\DLX_IDinst_RegFile_20_30/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_1002),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1078),
    .O(\DLX_IDinst_RegFile_20_30/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_20_30/CYINIT_2953  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_1001),
    .O(\DLX_IDinst_RegFile_20_30/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_20_22/LOGIC_ZERO_2954  (
    .O(\DLX_IDinst_RegFile_20_22/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_362_2955 (
    .IA(\DLX_IDinst_RegFile_20_22/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_20_22/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_421),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_362)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4211.INIT = 16'hBF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4211 (
    .ADR0(DLX_IDinst_RegFile_21_22),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_53),
    .ADR3(DLX_IDinst_RegFile_20_22),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_421)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4221.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4221 (
    .ADR0(DLX_IDinst_RegFile_22_22),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_54),
    .ADR3(DLX_IDinst_RegFile_23_22),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_422)
  );
  X_BUF \DLX_IDinst_RegFile_20_22/COUTUSED  (
    .I(\DLX_IDinst_RegFile_20_22/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_363)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_363_2956 (
    .IA(\DLX_IDinst_RegFile_20_22/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_362),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_422),
    .O(\DLX_IDinst_RegFile_20_22/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_20_22/CYINIT_2957  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_361),
    .O(\DLX_IDinst_RegFile_20_22/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_20_14/LOGIC_ZERO_2958  (
    .O(\DLX_IDinst_RegFile_20_14/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_234_2959 (
    .IA(\DLX_IDinst_RegFile_20_14/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_20_14/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_293),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_234)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2931.INIT = 16'hDFD5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2931 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_53),
    .ADR1(DLX_IDinst_RegFile_21_14),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR3(DLX_IDinst_RegFile_20_14),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_293)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_2941.INIT = 16'hBFB3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_2941 (
    .ADR0(DLX_IDinst_RegFile_23_14),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_54),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR3(DLX_IDinst_RegFile_22_14),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_294)
  );
  X_BUF \DLX_IDinst_RegFile_20_14/COUTUSED  (
    .I(\DLX_IDinst_RegFile_20_14/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_235)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_235_2960 (
    .IA(\DLX_IDinst_RegFile_20_14/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_234),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_294),
    .O(\DLX_IDinst_RegFile_20_14/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_20_14/CYINIT_2961  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_233),
    .O(\DLX_IDinst_RegFile_20_14/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_12_23/LOGIC_ZERO_2962  (
    .O(\DLX_IDinst_RegFile_12_23/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_374_2963 (
    .IA(\DLX_IDinst_RegFile_12_23/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_12_23/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_433),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_374)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4331.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4331 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_49),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR2(DLX_IDinst_RegFile_12_23),
    .ADR3(DLX_IDinst_RegFile_13_23),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_433)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4341.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4341 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR1(DLX_IDinst_RegFile_14_23),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_50),
    .ADR3(DLX_IDinst_RegFile_15_23),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_434)
  );
  X_BUF \DLX_IDinst_RegFile_12_23/COUTUSED  (
    .I(\DLX_IDinst_RegFile_12_23/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_375)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_375_2964 (
    .IA(\DLX_IDinst_RegFile_12_23/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_374),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_434),
    .O(\DLX_IDinst_RegFile_12_23/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_12_23/CYINIT_2965  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_373),
    .O(\DLX_IDinst_RegFile_12_23/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_12_15/LOGIC_ZERO_2966  (
    .O(\DLX_IDinst_RegFile_12_15/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_246_2967 (
    .IA(\DLX_IDinst_RegFile_12_15/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_12_15/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_305),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_246)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3051.INIT = 16'hFD5D;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3051 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_49),
    .ADR1(DLX_IDinst_RegFile_12_15),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR3(DLX_IDinst_RegFile_13_15),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_305)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3061.INIT = 16'hF5DD;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3061 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_50),
    .ADR1(DLX_IDinst_RegFile_14_15),
    .ADR2(DLX_IDinst_RegFile_15_15),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_306)
  );
  X_BUF \DLX_IDinst_RegFile_12_15/COUTUSED  (
    .I(\DLX_IDinst_RegFile_12_15/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_247)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_247_2968 (
    .IA(\DLX_IDinst_RegFile_12_15/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_246),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_306),
    .O(\DLX_IDinst_RegFile_12_15/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_12_15/CYINIT_2969  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_245),
    .O(\DLX_IDinst_RegFile_12_15/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_20_23/LOGIC_ZERO_2970  (
    .O(\DLX_IDinst_RegFile_20_23/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_378_2971 (
    .IA(\DLX_IDinst_RegFile_20_23/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_20_23/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_437),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_378)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4371.INIT = 16'hACFF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4371 (
    .ADR0(DLX_IDinst_RegFile_21_23),
    .ADR1(DLX_IDinst_RegFile_20_23),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_53),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_437)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4381.INIT = 16'hDF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4381 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR1(DLX_IDinst_RegFile_23_23),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_54),
    .ADR3(DLX_IDinst_RegFile_22_23),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_438)
  );
  X_BUF \DLX_IDinst_RegFile_20_23/COUTUSED  (
    .I(\DLX_IDinst_RegFile_20_23/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_379)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_379_2972 (
    .IA(\DLX_IDinst_RegFile_20_23/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_378),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_438),
    .O(\DLX_IDinst_RegFile_20_23/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_20_23/CYINIT_2973  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_377),
    .O(\DLX_IDinst_RegFile_20_23/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_20_15/LOGIC_ZERO_2974  (
    .O(\DLX_IDinst_RegFile_20_15/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_250_2975 (
    .IA(\DLX_IDinst_RegFile_20_15/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_20_15/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_309),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_250)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3091.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3091 (
    .ADR0(DLX_IDinst_RegFile_21_15),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_53),
    .ADR2(DLX_IDinst_RegFile_20_15),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_309)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3101.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3101 (
    .ADR0(DLX_IDinst_RegFile_23_15),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_54),
    .ADR2(DLX_IDinst_RegFile_22_15),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_310)
  );
  X_BUF \DLX_IDinst_RegFile_20_15/COUTUSED  (
    .I(\DLX_IDinst_RegFile_20_15/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_251)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_251_2976 (
    .IA(\DLX_IDinst_RegFile_20_15/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_250),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_310),
    .O(\DLX_IDinst_RegFile_20_15/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_20_15/CYINIT_2977  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_249),
    .O(\DLX_IDinst_RegFile_20_15/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_12_31/LOGIC_ZERO_2978  (
    .O(\DLX_IDinst_RegFile_12_31/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_1014_2979 (
    .IA(\DLX_IDinst_RegFile_12_31/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_12_31/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1089),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_1014)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10891.INIT = 16'hCFAF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10891 (
    .ADR0(DLX_IDinst_RegFile_12_31),
    .ADR1(DLX_IDinst_RegFile_13_31),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_577),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1089)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10901.INIT = 16'hAFCF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10901 (
    .ADR0(DLX_IDinst_RegFile_15_31),
    .ADR1(DLX_IDinst_RegFile_14_31),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_578),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1090)
  );
  X_BUF \DLX_IDinst_RegFile_12_31/COUTUSED  (
    .I(\DLX_IDinst_RegFile_12_31/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_1015)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_1015_2980 (
    .IA(\DLX_IDinst_RegFile_12_31/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_1014),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1090),
    .O(\DLX_IDinst_RegFile_12_31/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_12_31/CYINIT_2981  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_1013),
    .O(\DLX_IDinst_RegFile_12_31/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_20_31/LOGIC_ZERO_2982  (
    .O(\DLX_IDinst_RegFile_20_31/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_1018_2983 (
    .IA(\DLX_IDinst_RegFile_20_31/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_20_31/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1093),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_1018)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10931.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10931 (
    .ADR0(DLX_IDinst_RegFile_20_31),
    .ADR1(DLX_IDinst_RegFile_21_31),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_581),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1093)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10941.INIT = 16'hE2FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10941 (
    .ADR0(DLX_IDinst_RegFile_22_31),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR2(DLX_IDinst_RegFile_23_31),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_582),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1094)
  );
  X_BUF \DLX_IDinst_RegFile_20_31/COUTUSED  (
    .I(\DLX_IDinst_RegFile_20_31/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_1019)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_1019_2984 (
    .IA(\DLX_IDinst_RegFile_20_31/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_1018),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1094),
    .O(\DLX_IDinst_RegFile_20_31/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_20_31/CYINIT_2985  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_1017),
    .O(\DLX_IDinst_RegFile_20_31/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_12_24/LOGIC_ZERO_2986  (
    .O(\DLX_IDinst_RegFile_12_24/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_390_2987 (
    .IA(\DLX_IDinst_RegFile_12_24/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_12_24/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_449),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_390)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4491.INIT = 16'hFB73;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4491 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_49),
    .ADR2(DLX_IDinst_RegFile_12_24),
    .ADR3(DLX_IDinst_RegFile_13_24),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_449)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4501.INIT = 16'hD8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4501 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR1(DLX_IDinst_RegFile_15_24),
    .ADR2(DLX_IDinst_RegFile_14_24),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_50),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_450)
  );
  X_BUF \DLX_IDinst_RegFile_12_24/COUTUSED  (
    .I(\DLX_IDinst_RegFile_12_24/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_391)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_391_2988 (
    .IA(\DLX_IDinst_RegFile_12_24/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_390),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_450),
    .O(\DLX_IDinst_RegFile_12_24/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_12_24/CYINIT_2989  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_389),
    .O(\DLX_IDinst_RegFile_12_24/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_12_16/LOGIC_ZERO_2990  (
    .O(\DLX_IDinst_RegFile_12_16/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_262_2991 (
    .IA(\DLX_IDinst_RegFile_12_16/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_12_16/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_321),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_262)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3211.INIT = 16'hFB3B;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3211 (
    .ADR0(DLX_IDinst_RegFile_12_16),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_49),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR3(DLX_IDinst_RegFile_13_16),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_321)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3221.INIT = 16'hBFB3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3221 (
    .ADR0(DLX_IDinst_RegFile_15_16),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_50),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR3(DLX_IDinst_RegFile_14_16),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_322)
  );
  X_BUF \DLX_IDinst_RegFile_12_16/COUTUSED  (
    .I(\DLX_IDinst_RegFile_12_16/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_263)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_263_2992 (
    .IA(\DLX_IDinst_RegFile_12_16/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_262),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_322),
    .O(\DLX_IDinst_RegFile_12_16/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_12_16/CYINIT_2993  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_261),
    .O(\DLX_IDinst_RegFile_12_16/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_20_24/LOGIC_ZERO_2994  (
    .O(\DLX_IDinst_RegFile_20_24/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_394_2995 (
    .IA(\DLX_IDinst_RegFile_20_24/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_20_24/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_453),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_394)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4531.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4531 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_53),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR2(DLX_IDinst_RegFile_20_24),
    .ADR3(DLX_IDinst_RegFile_21_24),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_453)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4541.INIT = 16'hFD5D;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4541 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_54),
    .ADR1(DLX_IDinst_RegFile_22_24),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR3(DLX_IDinst_RegFile_23_24),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_454)
  );
  X_BUF \DLX_IDinst_RegFile_20_24/COUTUSED  (
    .I(\DLX_IDinst_RegFile_20_24/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_395)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_395_2996 (
    .IA(\DLX_IDinst_RegFile_20_24/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_394),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_454),
    .O(\DLX_IDinst_RegFile_20_24/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_20_24/CYINIT_2997  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_393),
    .O(\DLX_IDinst_RegFile_20_24/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_20_16/LOGIC_ZERO_2998  (
    .O(\DLX_IDinst_RegFile_20_16/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_266_2999 (
    .IA(\DLX_IDinst_RegFile_20_16/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_20_16/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_325),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_266)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3251.INIT = 16'hE2FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3251 (
    .ADR0(DLX_IDinst_RegFile_20_16),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR2(DLX_IDinst_RegFile_21_16),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_53),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_325)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3261.INIT = 16'hB8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3261 (
    .ADR0(DLX_IDinst_RegFile_23_16),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR2(DLX_IDinst_RegFile_22_16),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_54),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_326)
  );
  X_BUF \DLX_IDinst_RegFile_20_16/COUTUSED  (
    .I(\DLX_IDinst_RegFile_20_16/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_267)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_267_3000 (
    .IA(\DLX_IDinst_RegFile_20_16/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_266),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_326),
    .O(\DLX_IDinst_RegFile_20_16/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_20_16/CYINIT_3001  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_265),
    .O(\DLX_IDinst_RegFile_20_16/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_12_25/LOGIC_ZERO_3002  (
    .O(\DLX_IDinst_RegFile_12_25/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_406_3003 (
    .IA(\DLX_IDinst_RegFile_12_25/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_12_25/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_465),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_406)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4651.INIT = 16'hAFCF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4651 (
    .ADR0(DLX_IDinst_RegFile_13_25),
    .ADR1(DLX_IDinst_RegFile_12_25),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_49),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_465)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4661.INIT = 16'hDF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4661 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR1(DLX_IDinst_RegFile_15_25),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_50),
    .ADR3(DLX_IDinst_RegFile_14_25),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_466)
  );
  X_BUF \DLX_IDinst_RegFile_12_25/COUTUSED  (
    .I(\DLX_IDinst_RegFile_12_25/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_407)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_407_3004 (
    .IA(\DLX_IDinst_RegFile_12_25/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_406),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_466),
    .O(\DLX_IDinst_RegFile_12_25/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_12_25/CYINIT_3005  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_405),
    .O(\DLX_IDinst_RegFile_12_25/CYINIT )
  );
  defparam DLX_IDinst_RegFile_2_6_3006.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_2_6_3006 (
    .I(DLX_MEMinst_RF_data_in[6]),
    .CE(DLX_IDinst__n0554),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_2_6)
  );
  X_ZERO \DLX_IDinst_RegFile_12_17/LOGIC_ZERO_3007  (
    .O(\DLX_IDinst_RegFile_12_17/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_278_3008 (
    .IA(\DLX_IDinst_RegFile_12_17/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_12_17/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_337),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_278)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3371.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3371 (
    .ADR0(DLX_IDinst_RegFile_13_17),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_49),
    .ADR2(DLX_IDinst_RegFile_12_17),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_337)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3381.INIT = 16'hE4FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3381 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR1(DLX_IDinst_RegFile_14_17),
    .ADR2(DLX_IDinst_RegFile_15_17),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_50),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_338)
  );
  X_BUF \DLX_IDinst_RegFile_12_17/COUTUSED  (
    .I(\DLX_IDinst_RegFile_12_17/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_279)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_279_3009 (
    .IA(\DLX_IDinst_RegFile_12_17/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_278),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_338),
    .O(\DLX_IDinst_RegFile_12_17/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_12_17/CYINIT_3010  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_277),
    .O(\DLX_IDinst_RegFile_12_17/CYINIT )
  );
  defparam DLX_IDinst_Imm_0.INIT = 1'b0;
  X_SFF DLX_IDinst_Imm_0 (
    .I(DLX_IDinst__n0143[0]),
    .CE(DLX_IDinst__n0116),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_IDinst__n0115),
    .O(\DLX_IDinst_Imm[0] )
  );
  X_ZERO \DLX_IDinst_RegFile_20_25/LOGIC_ZERO_3011  (
    .O(\DLX_IDinst_RegFile_20_25/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_410_3012 (
    .IA(\DLX_IDinst_RegFile_20_25/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_20_25/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_469),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_410)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4691.INIT = 16'hD8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4691 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR1(DLX_IDinst_RegFile_21_25),
    .ADR2(DLX_IDinst_RegFile_20_25),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_53),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_469)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4701.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4701 (
    .ADR0(DLX_IDinst_RegFile_22_25),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_54),
    .ADR2(DLX_IDinst_RegFile_23_25),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_470)
  );
  X_BUF \DLX_IDinst_RegFile_20_25/COUTUSED  (
    .I(\DLX_IDinst_RegFile_20_25/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_411)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_411_3013 (
    .IA(\DLX_IDinst_RegFile_20_25/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_410),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_470),
    .O(\DLX_IDinst_RegFile_20_25/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_20_25/CYINIT_3014  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_409),
    .O(\DLX_IDinst_RegFile_20_25/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_20_17/LOGIC_ZERO_3015  (
    .O(\DLX_IDinst_RegFile_20_17/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_282_3016 (
    .IA(\DLX_IDinst_RegFile_20_17/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_20_17/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_341),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_282)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3411.INIT = 16'hDDF5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3411 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_53),
    .ADR1(DLX_IDinst_RegFile_21_17),
    .ADR2(DLX_IDinst_RegFile_20_17),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_341)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3421.INIT = 16'hFD5D;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3421 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_54),
    .ADR1(DLX_IDinst_RegFile_22_17),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_4 ),
    .ADR3(DLX_IDinst_RegFile_23_17),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_342)
  );
  X_BUF \DLX_IDinst_RegFile_20_17/COUTUSED  (
    .I(\DLX_IDinst_RegFile_20_17/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_283)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_283_3017 (
    .IA(\DLX_IDinst_RegFile_20_17/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_282),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_342),
    .O(\DLX_IDinst_RegFile_20_17/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_20_17/CYINIT_3018  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_281),
    .O(\DLX_IDinst_RegFile_20_17/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_12_26/LOGIC_ZERO_3019  (
    .O(\DLX_IDinst_RegFile_12_26/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_422_3020 (
    .IA(\DLX_IDinst_RegFile_12_26/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_12_26/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_481),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_422)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4811.INIT = 16'hF7B3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4811 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_49),
    .ADR2(DLX_IDinst_RegFile_13_26),
    .ADR3(DLX_IDinst_RegFile_12_26),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_481)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4821.INIT = 16'hDFD5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4821 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_50),
    .ADR1(DLX_IDinst_RegFile_15_26),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR3(DLX_IDinst_RegFile_14_26),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_482)
  );
  X_BUF \DLX_IDinst_RegFile_12_26/COUTUSED  (
    .I(\DLX_IDinst_RegFile_12_26/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_423)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_423_3021 (
    .IA(\DLX_IDinst_RegFile_12_26/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_422),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_482),
    .O(\DLX_IDinst_RegFile_12_26/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_12_26/CYINIT_3022  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_421),
    .O(\DLX_IDinst_RegFile_12_26/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_12_18/LOGIC_ZERO_3023  (
    .O(\DLX_IDinst_RegFile_12_18/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_806_3024 (
    .IA(\DLX_IDinst_RegFile_12_18/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_12_18/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_881),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_806)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8811.INIT = 16'hF7B3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8811 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_577),
    .ADR2(DLX_IDinst_RegFile_13_18),
    .ADR3(DLX_IDinst_RegFile_12_18),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_881)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8821.INIT = 16'hDDF5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8821 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_578),
    .ADR1(DLX_IDinst_RegFile_15_18),
    .ADR2(DLX_IDinst_RegFile_14_18),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_882)
  );
  X_BUF \DLX_IDinst_RegFile_12_18/COUTUSED  (
    .I(\DLX_IDinst_RegFile_12_18/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_807)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_807_3025 (
    .IA(\DLX_IDinst_RegFile_12_18/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_806),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_882),
    .O(\DLX_IDinst_RegFile_12_18/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_12_18/CYINIT_3026  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_805),
    .O(\DLX_IDinst_RegFile_12_18/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_13_10/LOGIC_ZERO_3027  (
    .O(\DLX_IDinst_RegFile_13_10/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_678_3028 (
    .IA(\DLX_IDinst_RegFile_13_10/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_13_10/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_753),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_678)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7531.INIT = 16'hB8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7531 (
    .ADR0(DLX_IDinst_RegFile_13_10),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR2(DLX_IDinst_RegFile_12_10),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_577),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_753)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7541.INIT = 16'hDDF5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7541 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_578),
    .ADR1(DLX_IDinst_RegFile_15_10),
    .ADR2(DLX_IDinst_RegFile_14_10),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_754)
  );
  X_BUF \DLX_IDinst_RegFile_13_10/COUTUSED  (
    .I(\DLX_IDinst_RegFile_13_10/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_679)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_679_3029 (
    .IA(\DLX_IDinst_RegFile_13_10/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_678),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_754),
    .O(\DLX_IDinst_RegFile_13_10/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_13_10/CYINIT_3030  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_677),
    .O(\DLX_IDinst_RegFile_13_10/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_20_26/LOGIC_ZERO_3031  (
    .O(\DLX_IDinst_RegFile_20_26/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_426_3032 (
    .IA(\DLX_IDinst_RegFile_20_26/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_20_26/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_485),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_426)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4851.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4851 (
    .ADR0(DLX_IDinst_RegFile_20_26),
    .ADR1(DLX_IDinst_RegFile_21_26),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_53),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_485)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4861.INIT = 16'hAFCF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4861 (
    .ADR0(DLX_IDinst_RegFile_23_26),
    .ADR1(DLX_IDinst_RegFile_22_26),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_54),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_486)
  );
  X_BUF \DLX_IDinst_RegFile_20_26/COUTUSED  (
    .I(\DLX_IDinst_RegFile_20_26/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_427)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_427_3033 (
    .IA(\DLX_IDinst_RegFile_20_26/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_426),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_486),
    .O(\DLX_IDinst_RegFile_20_26/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_20_26/CYINIT_3034  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_425),
    .O(\DLX_IDinst_RegFile_20_26/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_20_18/LOGIC_ZERO_3035  (
    .O(\DLX_IDinst_RegFile_20_18/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_298_3036 (
    .IA(\DLX_IDinst_RegFile_20_18/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_20_18/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_357),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_298)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3571.INIT = 16'hBFB3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3571 (
    .ADR0(DLX_IDinst_RegFile_21_18),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_53),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR3(DLX_IDinst_RegFile_20_18),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_357)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3581.INIT = 16'hFB3B;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3581 (
    .ADR0(DLX_IDinst_RegFile_22_18),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_54),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR3(DLX_IDinst_RegFile_23_18),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_358)
  );
  X_BUF \DLX_IDinst_RegFile_20_18/COUTUSED  (
    .I(\DLX_IDinst_RegFile_20_18/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_299)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_299_3037 (
    .IA(\DLX_IDinst_RegFile_20_18/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_298),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_358),
    .O(\DLX_IDinst_RegFile_20_18/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_20_18/CYINIT_3038  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_297),
    .O(\DLX_IDinst_RegFile_20_18/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_21_10/LOGIC_ZERO_3039  (
    .O(\DLX_IDinst_RegFile_21_10/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_682_3040 (
    .IA(\DLX_IDinst_RegFile_21_10/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_21_10/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_757),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_682)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7571.INIT = 16'hFB3B;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7571 (
    .ADR0(DLX_IDinst_RegFile_20_10),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_581),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR3(DLX_IDinst_RegFile_21_10),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_757)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7581.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7581 (
    .ADR0(DLX_IDinst_RegFile_22_10),
    .ADR1(DLX_IDinst_RegFile_23_10),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_582),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_758)
  );
  X_BUF \DLX_IDinst_RegFile_21_10/COUTUSED  (
    .I(\DLX_IDinst_RegFile_21_10/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_683)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_683_3041 (
    .IA(\DLX_IDinst_RegFile_21_10/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_682),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_758),
    .O(\DLX_IDinst_RegFile_21_10/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_21_10/CYINIT_3042  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_681),
    .O(\DLX_IDinst_RegFile_21_10/CYINIT )
  );
  defparam DLX_IFinst_PC_20.INIT = 1'b0;
  X_SFF DLX_IFinst_PC_20 (
    .I(DLX_IFinst_NPC[20]),
    .CE(DLX_IFinst_PC_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_IFinst_PC[20])
  );
  X_ZERO \DLX_IDinst_RegFile_12_27/LOGIC_ZERO_3043  (
    .O(\DLX_IDinst_RegFile_12_27/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_950_3044 (
    .IA(\DLX_IDinst_RegFile_12_27/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_12_27/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1025),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_950)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10251.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10251 (
    .ADR0(DLX_IDinst_jtarget[21]),
    .ADR1(DLX_IDinst_RegFile_12_27),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_577),
    .ADR3(DLX_IDinst_RegFile_13_27),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1025)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10261.INIT = 16'hBFB3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10261 (
    .ADR0(DLX_IDinst_RegFile_15_27),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_578),
    .ADR2(DLX_IDinst_jtarget[21]),
    .ADR3(DLX_IDinst_RegFile_14_27),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1026)
  );
  X_BUF \DLX_IDinst_RegFile_12_27/COUTUSED  (
    .I(\DLX_IDinst_RegFile_12_27/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_951)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_951_3045 (
    .IA(\DLX_IDinst_RegFile_12_27/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_950),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1026),
    .O(\DLX_IDinst_RegFile_12_27/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_12_27/CYINIT_3046  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_949),
    .O(\DLX_IDinst_RegFile_12_27/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_12_19/LOGIC_ZERO_3047  (
    .O(\DLX_IDinst_RegFile_12_19/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_310_3048 (
    .IA(\DLX_IDinst_RegFile_12_19/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_12_19/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_369),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_310)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3691.INIT = 16'hFB3B;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3691 (
    .ADR0(DLX_IDinst_RegFile_12_19),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_49),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR3(DLX_IDinst_RegFile_13_19),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_369)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3701.INIT = 16'hDFD5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3701 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_50),
    .ADR1(DLX_IDinst_RegFile_15_19),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR3(DLX_IDinst_RegFile_14_19),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_370)
  );
  X_BUF \DLX_IDinst_RegFile_12_19/COUTUSED  (
    .I(\DLX_IDinst_RegFile_12_19/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_311)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_311_3049 (
    .IA(\DLX_IDinst_RegFile_12_19/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_310),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_370),
    .O(\DLX_IDinst_RegFile_12_19/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_12_19/CYINIT_3050  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_309),
    .O(\DLX_IDinst_RegFile_12_19/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_13_11/LOGIC_ZERO_3051  (
    .O(\DLX_IDinst_RegFile_13_11/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_694_3052 (
    .IA(\DLX_IDinst_RegFile_13_11/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_13_11/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_769),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_694)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7691.INIT = 16'hF5DD;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7691 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_577),
    .ADR1(DLX_IDinst_RegFile_12_11),
    .ADR2(DLX_IDinst_RegFile_13_11),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_769)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7701.INIT = 16'hFB3B;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7701 (
    .ADR0(DLX_IDinst_RegFile_14_11),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_578),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR3(DLX_IDinst_RegFile_15_11),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_770)
  );
  X_BUF \DLX_IDinst_RegFile_13_11/COUTUSED  (
    .I(\DLX_IDinst_RegFile_13_11/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_695)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_695_3053 (
    .IA(\DLX_IDinst_RegFile_13_11/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_694),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_770),
    .O(\DLX_IDinst_RegFile_13_11/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_13_11/CYINIT_3054  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_693),
    .O(\DLX_IDinst_RegFile_13_11/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_20_27/LOGIC_ZERO_3055  (
    .O(\DLX_IDinst_RegFile_20_27/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_954_3056 (
    .IA(\DLX_IDinst_RegFile_20_27/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_20_27/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1029),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_954)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10291.INIT = 16'hF7B3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10291 (
    .ADR0(DLX_IDinst_jtarget[21]),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_581),
    .ADR2(DLX_IDinst_RegFile_21_27),
    .ADR3(DLX_IDinst_RegFile_20_27),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1029)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10301.INIT = 16'hCFAF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10301 (
    .ADR0(DLX_IDinst_RegFile_22_27),
    .ADR1(DLX_IDinst_RegFile_23_27),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_582),
    .ADR3(DLX_IDinst_jtarget[21]),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1030)
  );
  X_BUF \DLX_IDinst_RegFile_20_27/COUTUSED  (
    .I(\DLX_IDinst_RegFile_20_27/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_955)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_955_3057 (
    .IA(\DLX_IDinst_RegFile_20_27/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_954),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1030),
    .O(\DLX_IDinst_RegFile_20_27/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_20_27/CYINIT_3058  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_953),
    .O(\DLX_IDinst_RegFile_20_27/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_20_19/LOGIC_ZERO_3059  (
    .O(\DLX_IDinst_RegFile_20_19/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_314_3060 (
    .IA(\DLX_IDinst_RegFile_20_19/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_20_19/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_373),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_314)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3731.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3731 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_53),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR2(DLX_IDinst_RegFile_20_19),
    .ADR3(DLX_IDinst_RegFile_21_19),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_373)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_3741.INIT = 16'hBF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_3741 (
    .ADR0(DLX_IDinst_RegFile_23_19),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_3 ),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_54),
    .ADR3(DLX_IDinst_RegFile_22_19),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_374)
  );
  X_BUF \DLX_IDinst_RegFile_20_19/COUTUSED  (
    .I(\DLX_IDinst_RegFile_20_19/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_315)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_315_3061 (
    .IA(\DLX_IDinst_RegFile_20_19/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_314),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_374),
    .O(\DLX_IDinst_RegFile_20_19/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_20_19/CYINIT_3062  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_313),
    .O(\DLX_IDinst_RegFile_20_19/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_21_11/LOGIC_ZERO_3063  (
    .O(\DLX_IDinst_RegFile_21_11/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_698_3064 (
    .IA(\DLX_IDinst_RegFile_21_11/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_21_11/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_773),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_698)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7731.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7731 (
    .ADR0(DLX_IDinst_RegFile_20_11),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_581),
    .ADR3(DLX_IDinst_RegFile_21_11),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_773)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7741.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7741 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_582),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR2(DLX_IDinst_RegFile_22_11),
    .ADR3(DLX_IDinst_RegFile_23_11),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_774)
  );
  X_BUF \DLX_IDinst_RegFile_21_11/COUTUSED  (
    .I(\DLX_IDinst_RegFile_21_11/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_699)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_699_3065 (
    .IA(\DLX_IDinst_RegFile_21_11/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_698),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_774),
    .O(\DLX_IDinst_RegFile_21_11/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_21_11/CYINIT_3066  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_697),
    .O(\DLX_IDinst_RegFile_21_11/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_12_28/LOGIC_ZERO_3067  (
    .O(\DLX_IDinst_RegFile_12_28/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_966_3068 (
    .IA(\DLX_IDinst_RegFile_12_28/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_12_28/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1041),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_966)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10411.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10411 (
    .ADR0(DLX_IDinst_RegFile_12_28),
    .ADR1(DLX_IDinst_RegFile_13_28),
    .ADR2(DLX_IDinst_jtarget[21]),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_577),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1041)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10421.INIT = 16'hDF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10421 (
    .ADR0(DLX_IDinst_jtarget[21]),
    .ADR1(DLX_IDinst_RegFile_15_28),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_578),
    .ADR3(DLX_IDinst_RegFile_14_28),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1042)
  );
  X_BUF \DLX_IDinst_RegFile_12_28/COUTUSED  (
    .I(\DLX_IDinst_RegFile_12_28/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_967)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_967_3069 (
    .IA(\DLX_IDinst_RegFile_12_28/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_966),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1042),
    .O(\DLX_IDinst_RegFile_12_28/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_12_28/CYINIT_3070  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_965),
    .O(\DLX_IDinst_RegFile_12_28/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_13_20/LOGIC_ZERO_3071  (
    .O(\DLX_IDinst_RegFile_13_20/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_838_3072 (
    .IA(\DLX_IDinst_RegFile_13_20/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_13_20/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_913),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_838)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9131.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9131 (
    .ADR0(DLX_IDinst_RegFile_13_20),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_577),
    .ADR2(DLX_IDinst_RegFile_12_20),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_913)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9141.INIT = 16'hDDF5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9141 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_578),
    .ADR1(DLX_IDinst_RegFile_15_20),
    .ADR2(DLX_IDinst_RegFile_14_20),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_914)
  );
  X_BUF \DLX_IDinst_RegFile_13_20/COUTUSED  (
    .I(\DLX_IDinst_RegFile_13_20/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_839)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_839_3073 (
    .IA(\DLX_IDinst_RegFile_13_20/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_838),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_914),
    .O(\DLX_IDinst_RegFile_13_20/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_13_20/CYINIT_3074  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_837),
    .O(\DLX_IDinst_RegFile_13_20/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_13_12/LOGIC_ZERO_3075  (
    .O(\DLX_IDinst_RegFile_13_12/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_710_3076 (
    .IA(\DLX_IDinst_RegFile_13_12/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_13_12/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_785),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_710)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7851.INIT = 16'hD8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7851 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR1(DLX_IDinst_RegFile_13_12),
    .ADR2(DLX_IDinst_RegFile_12_12),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_577),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_785)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7861.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7861 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR1(DLX_IDinst_RegFile_14_12),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_578),
    .ADR3(DLX_IDinst_RegFile_15_12),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_786)
  );
  X_BUF \DLX_IDinst_RegFile_13_12/COUTUSED  (
    .I(\DLX_IDinst_RegFile_13_12/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_711)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_711_3077 (
    .IA(\DLX_IDinst_RegFile_13_12/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_710),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_786),
    .O(\DLX_IDinst_RegFile_13_12/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_13_12/CYINIT_3078  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_709),
    .O(\DLX_IDinst_RegFile_13_12/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_20_28/LOGIC_ZERO_3079  (
    .O(\DLX_IDinst_RegFile_20_28/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_970_3080 (
    .IA(\DLX_IDinst_RegFile_20_28/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_20_28/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1045),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_970)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10451.INIT = 16'hBF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10451 (
    .ADR0(DLX_IDinst_RegFile_21_28),
    .ADR1(DLX_IDinst_jtarget[21]),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_581),
    .ADR3(DLX_IDinst_RegFile_20_28),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1045)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10461.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10461 (
    .ADR0(DLX_IDinst_RegFile_22_28),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_582),
    .ADR2(DLX_IDinst_RegFile_23_28),
    .ADR3(DLX_IDinst_jtarget[21]),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1046)
  );
  X_BUF \DLX_IDinst_RegFile_20_28/COUTUSED  (
    .I(\DLX_IDinst_RegFile_20_28/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_971)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_971_3081 (
    .IA(\DLX_IDinst_RegFile_20_28/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_970),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1046),
    .O(\DLX_IDinst_RegFile_20_28/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_20_28/CYINIT_3082  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_969),
    .O(\DLX_IDinst_RegFile_20_28/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_21_20/LOGIC_ZERO_3083  (
    .O(\DLX_IDinst_RegFile_21_20/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_842_3084 (
    .IA(\DLX_IDinst_RegFile_21_20/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_21_20/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_917),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_842)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9171.INIT = 16'hF7D5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9171 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_581),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR2(DLX_IDinst_RegFile_21_20),
    .ADR3(DLX_IDinst_RegFile_20_20),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_917)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9181.INIT = 16'hCFAF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9181 (
    .ADR0(DLX_IDinst_RegFile_22_20),
    .ADR1(DLX_IDinst_RegFile_23_20),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_582),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_918)
  );
  X_BUF \DLX_IDinst_RegFile_21_20/COUTUSED  (
    .I(\DLX_IDinst_RegFile_21_20/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_843)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_843_3085 (
    .IA(\DLX_IDinst_RegFile_21_20/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_842),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_918),
    .O(\DLX_IDinst_RegFile_21_20/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_21_20/CYINIT_3086  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_841),
    .O(\DLX_IDinst_RegFile_21_20/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_21_12/LOGIC_ZERO_3087  (
    .O(\DLX_IDinst_RegFile_21_12/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_714_3088 (
    .IA(\DLX_IDinst_RegFile_21_12/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_21_12/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_789),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_714)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7891.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7891 (
    .ADR0(DLX_IDinst_RegFile_21_12),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_581),
    .ADR2(DLX_IDinst_RegFile_20_12),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_789)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7901.INIT = 16'hF5DD;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7901 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_582),
    .ADR1(DLX_IDinst_RegFile_22_12),
    .ADR2(DLX_IDinst_RegFile_23_12),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_790)
  );
  X_BUF \DLX_IDinst_RegFile_21_12/COUTUSED  (
    .I(\DLX_IDinst_RegFile_21_12/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_715)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_715_3089 (
    .IA(\DLX_IDinst_RegFile_21_12/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_714),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_790),
    .O(\DLX_IDinst_RegFile_21_12/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_21_12/CYINIT_3090  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_713),
    .O(\DLX_IDinst_RegFile_21_12/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_12_29/LOGIC_ZERO_3091  (
    .O(\DLX_IDinst_RegFile_12_29/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_982_3092 (
    .IA(\DLX_IDinst_RegFile_12_29/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_12_29/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1057),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_982)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10571.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10571 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR1(DLX_IDinst_RegFile_12_29),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_577),
    .ADR3(DLX_IDinst_RegFile_13_29),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1057)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10581.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10581 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_578),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR2(DLX_IDinst_RegFile_14_29),
    .ADR3(DLX_IDinst_RegFile_15_29),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1058)
  );
  X_BUF \DLX_IDinst_RegFile_12_29/COUTUSED  (
    .I(\DLX_IDinst_RegFile_12_29/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_983)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_983_3093 (
    .IA(\DLX_IDinst_RegFile_12_29/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_982),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1058),
    .O(\DLX_IDinst_RegFile_12_29/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_12_29/CYINIT_3094  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_981),
    .O(\DLX_IDinst_RegFile_12_29/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_13_21/LOGIC_ZERO_3095  (
    .O(\DLX_IDinst_RegFile_13_21/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_854_3096 (
    .IA(\DLX_IDinst_RegFile_13_21/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_13_21/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_929),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_854)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9291.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9291 (
    .ADR0(DLX_IDinst_RegFile_12_21),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_577),
    .ADR3(DLX_IDinst_RegFile_13_21),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_929)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9301.INIT = 16'hACFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9301 (
    .ADR0(DLX_IDinst_RegFile_15_21),
    .ADR1(DLX_IDinst_RegFile_14_21),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_578),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_930)
  );
  X_BUF \DLX_IDinst_RegFile_13_21/COUTUSED  (
    .I(\DLX_IDinst_RegFile_13_21/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_855)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_855_3097 (
    .IA(\DLX_IDinst_RegFile_13_21/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_854),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_930),
    .O(\DLX_IDinst_RegFile_13_21/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_13_21/CYINIT_3098  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_853),
    .O(\DLX_IDinst_RegFile_13_21/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_13_13/LOGIC_ZERO_3099  (
    .O(\DLX_IDinst_RegFile_13_13/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_726_3100 (
    .IA(\DLX_IDinst_RegFile_13_13/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_13_13/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_801),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_726)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8011.INIT = 16'hF7D5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8011 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_577),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR2(DLX_IDinst_RegFile_13_13),
    .ADR3(DLX_IDinst_RegFile_12_13),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_801)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8021.INIT = 16'hE4FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8021 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR1(DLX_IDinst_RegFile_14_13),
    .ADR2(DLX_IDinst_RegFile_15_13),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_578),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_802)
  );
  X_BUF \DLX_IDinst_RegFile_13_13/COUTUSED  (
    .I(\DLX_IDinst_RegFile_13_13/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_727)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_727_3101 (
    .IA(\DLX_IDinst_RegFile_13_13/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_726),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_802),
    .O(\DLX_IDinst_RegFile_13_13/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_13_13/CYINIT_3102  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_725),
    .O(\DLX_IDinst_RegFile_13_13/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_20_29/LOGIC_ZERO_3103  (
    .O(\DLX_IDinst_RegFile_20_29/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_986_3104 (
    .IA(\DLX_IDinst_RegFile_20_29/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_20_29/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1061),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_986)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10611.INIT = 16'hE2FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10611 (
    .ADR0(DLX_IDinst_RegFile_20_29),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR2(DLX_IDinst_RegFile_21_29),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_581),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1061)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10621.INIT = 16'hF7D5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10621 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_582),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_5 ),
    .ADR2(DLX_IDinst_RegFile_23_29),
    .ADR3(DLX_IDinst_RegFile_22_29),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1062)
  );
  X_BUF \DLX_IDinst_RegFile_20_29/COUTUSED  (
    .I(\DLX_IDinst_RegFile_20_29/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_987)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_987_3105 (
    .IA(\DLX_IDinst_RegFile_20_29/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_986),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1062),
    .O(\DLX_IDinst_RegFile_20_29/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_20_29/CYINIT_3106  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_985),
    .O(\DLX_IDinst_RegFile_20_29/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_21_21/LOGIC_ZERO_3107  (
    .O(\DLX_IDinst_RegFile_21_21/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_858_3108 (
    .IA(\DLX_IDinst_RegFile_21_21/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_21_21/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_933),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_858)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9331.INIT = 16'hFB3B;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9331 (
    .ADR0(DLX_IDinst_RegFile_20_21),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_581),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR3(DLX_IDinst_RegFile_21_21),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_933)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9341.INIT = 16'hACFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9341 (
    .ADR0(DLX_IDinst_RegFile_23_21),
    .ADR1(DLX_IDinst_RegFile_22_21),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_582),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_934)
  );
  X_BUF \DLX_IDinst_RegFile_21_21/COUTUSED  (
    .I(\DLX_IDinst_RegFile_21_21/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_859)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_859_3109 (
    .IA(\DLX_IDinst_RegFile_21_21/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_858),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_934),
    .O(\DLX_IDinst_RegFile_21_21/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_21_21/CYINIT_3110  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_857),
    .O(\DLX_IDinst_RegFile_21_21/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_21_13/LOGIC_ZERO_3111  (
    .O(\DLX_IDinst_RegFile_21_13/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_730_3112 (
    .IA(\DLX_IDinst_RegFile_21_13/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_21_13/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_805),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_730)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8051.INIT = 16'hD8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8051 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR1(DLX_IDinst_RegFile_21_13),
    .ADR2(DLX_IDinst_RegFile_20_13),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_581),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_805)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8061.INIT = 16'hFB73;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8061 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_582),
    .ADR2(DLX_IDinst_RegFile_22_13),
    .ADR3(DLX_IDinst_RegFile_23_13),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_806)
  );
  X_BUF \DLX_IDinst_RegFile_21_13/COUTUSED  (
    .I(\DLX_IDinst_RegFile_21_13/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_731)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_731_3113 (
    .IA(\DLX_IDinst_RegFile_21_13/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_730),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_806),
    .O(\DLX_IDinst_RegFile_21_13/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_21_13/CYINIT_3114  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_729),
    .O(\DLX_IDinst_RegFile_21_13/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_13_30/LOGIC_ZERO_3115  (
    .O(\DLX_IDinst_RegFile_13_30/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_486_3116 (
    .IA(\DLX_IDinst_RegFile_13_30/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_13_30/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_545),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_486)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5451.INIT = 16'hF7D5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5451 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_49),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR2(DLX_IDinst_RegFile_13_30),
    .ADR3(DLX_IDinst_RegFile_12_30),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_545)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5461.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5461 (
    .ADR0(DLX_IDinst_RegFile_14_30),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_50),
    .ADR2(DLX_IDinst_RegFile_15_30),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_546)
  );
  X_BUF \DLX_IDinst_RegFile_13_30/COUTUSED  (
    .I(\DLX_IDinst_RegFile_13_30/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_487)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_487_3117 (
    .IA(\DLX_IDinst_RegFile_13_30/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_486),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_546),
    .O(\DLX_IDinst_RegFile_13_30/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_13_30/CYINIT_3118  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_485),
    .O(\DLX_IDinst_RegFile_13_30/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_13_22/LOGIC_ZERO_3119  (
    .O(\DLX_IDinst_RegFile_13_22/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_870_3120 (
    .IA(\DLX_IDinst_RegFile_13_22/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_13_22/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_945),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_870)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9451.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9451 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_577),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR2(DLX_IDinst_RegFile_12_22),
    .ADR3(DLX_IDinst_RegFile_13_22),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_945)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9461.INIT = 16'hBFB3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9461 (
    .ADR0(DLX_IDinst_RegFile_15_22),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_578),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR3(DLX_IDinst_RegFile_14_22),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_946)
  );
  X_BUF \DLX_IDinst_RegFile_13_22/COUTUSED  (
    .I(\DLX_IDinst_RegFile_13_22/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_871)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_871_3121 (
    .IA(\DLX_IDinst_RegFile_13_22/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_870),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_946),
    .O(\DLX_IDinst_RegFile_13_22/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_13_22/CYINIT_3122  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_869),
    .O(\DLX_IDinst_RegFile_13_22/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_13_14/LOGIC_ZERO_3123  (
    .O(\DLX_IDinst_RegFile_13_14/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_742_3124 (
    .IA(\DLX_IDinst_RegFile_13_14/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_13_14/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_817),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_742)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8171.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8171 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_577),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR2(DLX_IDinst_RegFile_12_14),
    .ADR3(DLX_IDinst_RegFile_13_14),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_817)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8181.INIT = 16'hD8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8181 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR1(DLX_IDinst_RegFile_15_14),
    .ADR2(DLX_IDinst_RegFile_14_14),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_578),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_818)
  );
  X_BUF \DLX_IDinst_RegFile_13_14/COUTUSED  (
    .I(\DLX_IDinst_RegFile_13_14/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_743)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_743_3125 (
    .IA(\DLX_IDinst_RegFile_13_14/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_742),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_818),
    .O(\DLX_IDinst_RegFile_13_14/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_13_14/CYINIT_3126  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_741),
    .O(\DLX_IDinst_RegFile_13_14/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_21_30/LOGIC_ZERO_3127  (
    .O(\DLX_IDinst_RegFile_21_30/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_490_3128 (
    .IA(\DLX_IDinst_RegFile_21_30/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_21_30/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_549),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_490)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5491.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5491 (
    .ADR0(DLX_IDinst_RegFile_21_30),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_53),
    .ADR2(DLX_IDinst_RegFile_20_30),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_549)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5501.INIT = 16'hBF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5501 (
    .ADR0(DLX_IDinst_RegFile_23_30),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_54),
    .ADR3(DLX_IDinst_RegFile_22_30),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_550)
  );
  X_BUF \DLX_IDinst_RegFile_21_30/COUTUSED  (
    .I(\DLX_IDinst_RegFile_21_30/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_491)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_491_3129 (
    .IA(\DLX_IDinst_RegFile_21_30/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_490),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_550),
    .O(\DLX_IDinst_RegFile_21_30/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_21_30/CYINIT_3130  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_489),
    .O(\DLX_IDinst_RegFile_21_30/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_21_22/LOGIC_ZERO_3131  (
    .O(\DLX_IDinst_RegFile_21_22/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_874_3132 (
    .IA(\DLX_IDinst_RegFile_21_22/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_21_22/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_949),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_874)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9491.INIT = 16'hFD5D;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9491 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_581),
    .ADR1(DLX_IDinst_RegFile_20_22),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR3(DLX_IDinst_RegFile_21_22),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_949)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9501.INIT = 16'hDFD5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9501 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_582),
    .ADR1(DLX_IDinst_RegFile_23_22),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR3(DLX_IDinst_RegFile_22_22),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_950)
  );
  X_BUF \DLX_IDinst_RegFile_21_22/COUTUSED  (
    .I(\DLX_IDinst_RegFile_21_22/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_875)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_875_3133 (
    .IA(\DLX_IDinst_RegFile_21_22/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_874),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_950),
    .O(\DLX_IDinst_RegFile_21_22/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_21_22/CYINIT_3134  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_873),
    .O(\DLX_IDinst_RegFile_21_22/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_21_14/LOGIC_ZERO_3135  (
    .O(\DLX_IDinst_RegFile_21_14/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_746_3136 (
    .IA(\DLX_IDinst_RegFile_21_14/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_21_14/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_821),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_746)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8211.INIT = 16'hB8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8211 (
    .ADR0(DLX_IDinst_RegFile_21_14),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR2(DLX_IDinst_RegFile_20_14),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_581),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_821)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8221.INIT = 16'hACFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8221 (
    .ADR0(DLX_IDinst_RegFile_23_14),
    .ADR1(DLX_IDinst_RegFile_22_14),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_582),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_822)
  );
  X_BUF \DLX_IDinst_RegFile_21_14/COUTUSED  (
    .I(\DLX_IDinst_RegFile_21_14/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_747)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_747_3137 (
    .IA(\DLX_IDinst_RegFile_21_14/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_746),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_822),
    .O(\DLX_IDinst_RegFile_21_14/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_21_14/CYINIT_3138  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_745),
    .O(\DLX_IDinst_RegFile_21_14/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_13_23/LOGIC_ZERO_3139  (
    .O(\DLX_IDinst_RegFile_13_23/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_886_3140 (
    .IA(\DLX_IDinst_RegFile_13_23/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_13_23/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_961),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_886)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9611.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9611 (
    .ADR0(DLX_IDinst_RegFile_12_23),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_577),
    .ADR3(DLX_IDinst_RegFile_13_23),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_961)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9621.INIT = 16'hDFD5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9621 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_578),
    .ADR1(DLX_IDinst_RegFile_15_23),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR3(DLX_IDinst_RegFile_14_23),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_962)
  );
  X_BUF \DLX_IDinst_RegFile_13_23/COUTUSED  (
    .I(\DLX_IDinst_RegFile_13_23/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_887)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_887_3141 (
    .IA(\DLX_IDinst_RegFile_13_23/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_886),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_962),
    .O(\DLX_IDinst_RegFile_13_23/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_13_23/CYINIT_3142  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_885),
    .O(\DLX_IDinst_RegFile_13_23/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_13_15/LOGIC_ZERO_3143  (
    .O(\DLX_IDinst_RegFile_13_15/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_758_3144 (
    .IA(\DLX_IDinst_RegFile_13_15/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_13_15/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_833),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_758)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8331.INIT = 16'hE2FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8331 (
    .ADR0(DLX_IDinst_RegFile_12_15),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR2(DLX_IDinst_RegFile_13_15),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_577),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_833)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8341.INIT = 16'hAFCF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8341 (
    .ADR0(DLX_IDinst_RegFile_15_15),
    .ADR1(DLX_IDinst_RegFile_14_15),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_578),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_834)
  );
  X_BUF \DLX_IDinst_RegFile_13_15/COUTUSED  (
    .I(\DLX_IDinst_RegFile_13_15/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_759)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_759_3145 (
    .IA(\DLX_IDinst_RegFile_13_15/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_758),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_834),
    .O(\DLX_IDinst_RegFile_13_15/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_13_15/CYINIT_3146  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_757),
    .O(\DLX_IDinst_RegFile_13_15/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_21_23/LOGIC_ZERO_3147  (
    .O(\DLX_IDinst_RegFile_21_23/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_890_3148 (
    .IA(\DLX_IDinst_RegFile_21_23/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_21_23/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_965),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_890)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9651.INIT = 16'hCFAF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9651 (
    .ADR0(DLX_IDinst_RegFile_20_23),
    .ADR1(DLX_IDinst_RegFile_21_23),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_581),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_965)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9661.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9661 (
    .ADR0(DLX_IDinst_RegFile_22_23),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_582),
    .ADR2(DLX_IDinst_RegFile_23_23),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_966)
  );
  X_BUF \DLX_IDinst_RegFile_21_23/COUTUSED  (
    .I(\DLX_IDinst_RegFile_21_23/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_891)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_891_3149 (
    .IA(\DLX_IDinst_RegFile_21_23/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_890),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_966),
    .O(\DLX_IDinst_RegFile_21_23/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_21_23/CYINIT_3150  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_889),
    .O(\DLX_IDinst_RegFile_21_23/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_21_15/LOGIC_ZERO_3151  (
    .O(\DLX_IDinst_RegFile_21_15/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_762_3152 (
    .IA(\DLX_IDinst_RegFile_21_15/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_21_15/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_837),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_762)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8371.INIT = 16'hDF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8371 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR1(DLX_IDinst_RegFile_21_15),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_581),
    .ADR3(DLX_IDinst_RegFile_20_15),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_837)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8381.INIT = 16'hD8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8381 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR1(DLX_IDinst_RegFile_23_15),
    .ADR2(DLX_IDinst_RegFile_22_15),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_582),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_838)
  );
  X_BUF \DLX_IDinst_RegFile_21_15/COUTUSED  (
    .I(\DLX_IDinst_RegFile_21_15/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_763)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_763_3153 (
    .IA(\DLX_IDinst_RegFile_21_15/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_762),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_838),
    .O(\DLX_IDinst_RegFile_21_15/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_21_15/CYINIT_3154  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_761),
    .O(\DLX_IDinst_RegFile_21_15/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_13_31/LOGIC_ZERO_3155  (
    .O(\DLX_IDinst_RegFile_13_31/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_502_3156 (
    .IA(\DLX_IDinst_RegFile_13_31/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_13_31/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_561),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_502)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5611.INIT = 16'hE2FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5611 (
    .ADR0(DLX_IDinst_RegFile_12_31),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR2(DLX_IDinst_RegFile_13_31),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_49),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_561)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5621.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5621 (
    .ADR0(DLX_IDinst_RegFile_14_31),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_50),
    .ADR3(DLX_IDinst_RegFile_15_31),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_562)
  );
  X_BUF \DLX_IDinst_RegFile_13_31/COUTUSED  (
    .I(\DLX_IDinst_RegFile_13_31/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_503)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_503_3157 (
    .IA(\DLX_IDinst_RegFile_13_31/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_502),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_562),
    .O(\DLX_IDinst_RegFile_13_31/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_13_31/CYINIT_3158  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_501),
    .O(\DLX_IDinst_RegFile_13_31/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_21_31/LOGIC_ZERO_3159  (
    .O(\DLX_IDinst_RegFile_21_31/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_506_3160 (
    .IA(\DLX_IDinst_RegFile_21_31/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_21_31/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_565),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_506)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5651.INIT = 16'hD8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5651 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR1(DLX_IDinst_RegFile_21_31),
    .ADR2(DLX_IDinst_RegFile_20_31),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_53),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_565)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5661.INIT = 16'hCFAF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5661 (
    .ADR0(DLX_IDinst_RegFile_22_31),
    .ADR1(DLX_IDinst_RegFile_23_31),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_54),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_566)
  );
  X_BUF \DLX_IDinst_RegFile_21_31/COUTUSED  (
    .I(\DLX_IDinst_RegFile_21_31/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_507)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_507_3161 (
    .IA(\DLX_IDinst_RegFile_21_31/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_506),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_566),
    .O(\DLX_IDinst_RegFile_21_31/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_21_31/CYINIT_3162  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_505),
    .O(\DLX_IDinst_RegFile_21_31/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_13_24/LOGIC_ZERO_3163  (
    .O(\DLX_IDinst_RegFile_13_24/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_902_3164 (
    .IA(\DLX_IDinst_RegFile_13_24/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_13_24/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_977),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_902)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9771.INIT = 16'hE4FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9771 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR1(DLX_IDinst_RegFile_12_24),
    .ADR2(DLX_IDinst_RegFile_13_24),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_577),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_977)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9781.INIT = 16'hF7D5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9781 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_578),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR2(DLX_IDinst_RegFile_15_24),
    .ADR3(DLX_IDinst_RegFile_14_24),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_978)
  );
  X_BUF \DLX_IDinst_RegFile_13_24/COUTUSED  (
    .I(\DLX_IDinst_RegFile_13_24/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_903)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_903_3165 (
    .IA(\DLX_IDinst_RegFile_13_24/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_902),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_978),
    .O(\DLX_IDinst_RegFile_13_24/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_13_24/CYINIT_3166  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_901),
    .O(\DLX_IDinst_RegFile_13_24/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_13_16/LOGIC_ZERO_3167  (
    .O(\DLX_IDinst_RegFile_13_16/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_774_3168 (
    .IA(\DLX_IDinst_RegFile_13_16/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_13_16/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_849),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_774)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8491.INIT = 16'hDFD5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8491 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_577),
    .ADR1(DLX_IDinst_RegFile_13_16),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR3(DLX_IDinst_RegFile_12_16),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_849)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8501.INIT = 16'hFD5D;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8501 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_578),
    .ADR1(DLX_IDinst_RegFile_14_16),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR3(DLX_IDinst_RegFile_15_16),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_850)
  );
  X_BUF \DLX_IDinst_RegFile_13_16/COUTUSED  (
    .I(\DLX_IDinst_RegFile_13_16/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_775)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_775_3169 (
    .IA(\DLX_IDinst_RegFile_13_16/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_774),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_850),
    .O(\DLX_IDinst_RegFile_13_16/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_13_16/CYINIT_3170  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_773),
    .O(\DLX_IDinst_RegFile_13_16/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_21_24/LOGIC_ZERO_3171  (
    .O(\DLX_IDinst_RegFile_21_24/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_906_3172 (
    .IA(\DLX_IDinst_RegFile_21_24/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_21_24/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_981),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_906)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9811.INIT = 16'hFB73;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9811 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_581),
    .ADR2(DLX_IDinst_RegFile_20_24),
    .ADR3(DLX_IDinst_RegFile_21_24),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_981)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9821.INIT = 16'hBFB3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9821 (
    .ADR0(DLX_IDinst_RegFile_23_24),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_582),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR3(DLX_IDinst_RegFile_22_24),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_982)
  );
  X_BUF \DLX_IDinst_RegFile_21_24/COUTUSED  (
    .I(\DLX_IDinst_RegFile_21_24/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_907)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_907_3173 (
    .IA(\DLX_IDinst_RegFile_21_24/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_906),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_982),
    .O(\DLX_IDinst_RegFile_21_24/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_21_24/CYINIT_3174  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_905),
    .O(\DLX_IDinst_RegFile_21_24/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_21_16/LOGIC_ZERO_3175  (
    .O(\DLX_IDinst_RegFile_21_16/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_778_3176 (
    .IA(\DLX_IDinst_RegFile_21_16/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_21_16/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_853),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_778)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8531.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8531 (
    .ADR0(DLX_IDinst_RegFile_20_16),
    .ADR1(DLX_IDinst_RegFile_21_16),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_581),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_853)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8541.INIT = 16'hFB3B;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8541 (
    .ADR0(DLX_IDinst_RegFile_22_16),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_582),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR3(DLX_IDinst_RegFile_23_16),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_854)
  );
  X_BUF \DLX_IDinst_RegFile_21_16/COUTUSED  (
    .I(\DLX_IDinst_RegFile_21_16/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_779)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_779_3177 (
    .IA(\DLX_IDinst_RegFile_21_16/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_778),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_854),
    .O(\DLX_IDinst_RegFile_21_16/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_21_16/CYINIT_3178  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_777),
    .O(\DLX_IDinst_RegFile_21_16/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_13_25/LOGIC_ZERO_3179  (
    .O(\DLX_IDinst_RegFile_13_25/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_918_3180 (
    .IA(\DLX_IDinst_RegFile_13_25/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_13_25/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_993),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_918)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9931.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9931 (
    .ADR0(DLX_IDinst_RegFile_12_25),
    .ADR1(DLX_IDinst_RegFile_13_25),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_577),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_993)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9941.INIT = 16'hCFAF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9941 (
    .ADR0(DLX_IDinst_RegFile_14_25),
    .ADR1(DLX_IDinst_RegFile_15_25),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_578),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_994)
  );
  X_BUF \DLX_IDinst_RegFile_13_25/COUTUSED  (
    .I(\DLX_IDinst_RegFile_13_25/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_919)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_919_3181 (
    .IA(\DLX_IDinst_RegFile_13_25/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_918),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_994),
    .O(\DLX_IDinst_RegFile_13_25/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_13_25/CYINIT_3182  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_917),
    .O(\DLX_IDinst_RegFile_13_25/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_13_17/LOGIC_ZERO_3183  (
    .O(\DLX_IDinst_RegFile_13_17/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_790_3184 (
    .IA(\DLX_IDinst_RegFile_13_17/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_13_17/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_865),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_790)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8651.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8651 (
    .ADR0(DLX_IDinst_RegFile_12_17),
    .ADR1(DLX_IDinst_RegFile_13_17),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_577),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_865)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8661.INIT = 16'hF5DD;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8661 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_578),
    .ADR1(DLX_IDinst_RegFile_14_17),
    .ADR2(DLX_IDinst_RegFile_15_17),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_866)
  );
  X_BUF \DLX_IDinst_RegFile_13_17/COUTUSED  (
    .I(\DLX_IDinst_RegFile_13_17/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_791)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_791_3185 (
    .IA(\DLX_IDinst_RegFile_13_17/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_790),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_866),
    .O(\DLX_IDinst_RegFile_13_17/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_13_17/CYINIT_3186  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_789),
    .O(\DLX_IDinst_RegFile_13_17/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_21_25/LOGIC_ZERO_3187  (
    .O(\DLX_IDinst_RegFile_21_25/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_922_3188 (
    .IA(\DLX_IDinst_RegFile_21_25/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_21_25/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_997),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_922)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9971.INIT = 16'hF5DD;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9971 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_581),
    .ADR1(DLX_IDinst_RegFile_20_25),
    .ADR2(DLX_IDinst_RegFile_21_25),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_997)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9981.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9981 (
    .ADR0(DLX_IDinst_RegFile_22_25),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_582),
    .ADR3(DLX_IDinst_RegFile_23_25),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_998)
  );
  X_BUF \DLX_IDinst_RegFile_21_25/COUTUSED  (
    .I(\DLX_IDinst_RegFile_21_25/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_923)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_923_3189 (
    .IA(\DLX_IDinst_RegFile_21_25/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_922),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_998),
    .O(\DLX_IDinst_RegFile_21_25/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_21_25/CYINIT_3190  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_921),
    .O(\DLX_IDinst_RegFile_21_25/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_21_17/LOGIC_ZERO_3191  (
    .O(\DLX_IDinst_RegFile_21_17/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_794_3192 (
    .IA(\DLX_IDinst_RegFile_21_17/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_21_17/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_869),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_794)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8691.INIT = 16'hFD5D;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8691 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_581),
    .ADR1(DLX_IDinst_RegFile_20_17),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR3(DLX_IDinst_RegFile_21_17),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_869)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8701.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8701 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_582),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR2(DLX_IDinst_RegFile_22_17),
    .ADR3(DLX_IDinst_RegFile_23_17),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_870)
  );
  X_BUF \DLX_IDinst_RegFile_21_17/COUTUSED  (
    .I(\DLX_IDinst_RegFile_21_17/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_795)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_795_3193 (
    .IA(\DLX_IDinst_RegFile_21_17/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_794),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_870),
    .O(\DLX_IDinst_RegFile_21_17/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_21_17/CYINIT_3194  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_793),
    .O(\DLX_IDinst_RegFile_21_17/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_13_26/LOGIC_ZERO_3195  (
    .O(\DLX_IDinst_RegFile_13_26/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_934_3196 (
    .IA(\DLX_IDinst_RegFile_13_26/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_13_26/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1009),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_934)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10091.INIT = 16'hBFB3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10091 (
    .ADR0(DLX_IDinst_RegFile_13_26),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_577),
    .ADR2(DLX_IDinst_jtarget[21]),
    .ADR3(DLX_IDinst_RegFile_12_26),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1009)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10101.INIT = 16'hDFD5;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10101 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_578),
    .ADR1(DLX_IDinst_RegFile_15_26),
    .ADR2(DLX_IDinst_jtarget[21]),
    .ADR3(DLX_IDinst_RegFile_14_26),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1010)
  );
  X_BUF \DLX_IDinst_RegFile_13_26/COUTUSED  (
    .I(\DLX_IDinst_RegFile_13_26/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_935)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_935_3197 (
    .IA(\DLX_IDinst_RegFile_13_26/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_934),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1010),
    .O(\DLX_IDinst_RegFile_13_26/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_13_26/CYINIT_3198  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_933),
    .O(\DLX_IDinst_RegFile_13_26/CYINIT )
  );
  defparam DLX_IFinst_PC_30.INIT = 1'b0;
  X_SFF DLX_IFinst_PC_30 (
    .I(DLX_IFinst_NPC[30]),
    .CE(DLX_IFinst_PC_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_IFinst_PC[30])
  );
  X_ZERO \DLX_IDinst_RegFile_21_26/LOGIC_ZERO_3199  (
    .O(\DLX_IDinst_RegFile_21_26/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_938_3200 (
    .IA(\DLX_IDinst_RegFile_21_26/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_21_26/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1013),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_938)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10131.INIT = 16'hF7B3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10131 (
    .ADR0(DLX_IDinst_jtarget[21]),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_581),
    .ADR2(DLX_IDinst_RegFile_21_26),
    .ADR3(DLX_IDinst_RegFile_20_26),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1013)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_10141.INIT = 16'hF7B3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_10141 (
    .ADR0(DLX_IDinst_jtarget[21]),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_582),
    .ADR2(DLX_IDinst_RegFile_23_26),
    .ADR3(DLX_IDinst_RegFile_22_26),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_1014)
  );
  X_BUF \DLX_IDinst_RegFile_21_26/COUTUSED  (
    .I(\DLX_IDinst_RegFile_21_26/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_939)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_939_3201 (
    .IA(\DLX_IDinst_RegFile_21_26/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_938),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_1014),
    .O(\DLX_IDinst_RegFile_21_26/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_21_26/CYINIT_3202  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_937),
    .O(\DLX_IDinst_RegFile_21_26/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_21_18/LOGIC_ZERO_3203  (
    .O(\DLX_IDinst_RegFile_21_18/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_810_3204 (
    .IA(\DLX_IDinst_RegFile_21_18/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_21_18/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_885),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_810)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8851.INIT = 16'hFD5D;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8851 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_581),
    .ADR1(DLX_IDinst_RegFile_20_18),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR3(DLX_IDinst_RegFile_21_18),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_885)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8861.INIT = 16'hDF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8861 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR1(DLX_IDinst_RegFile_23_18),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_582),
    .ADR3(DLX_IDinst_RegFile_22_18),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_886)
  );
  X_BUF \DLX_IDinst_RegFile_21_18/COUTUSED  (
    .I(\DLX_IDinst_RegFile_21_18/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_811)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_811_3205 (
    .IA(\DLX_IDinst_RegFile_21_18/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_810),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_886),
    .O(\DLX_IDinst_RegFile_21_18/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_21_18/CYINIT_3206  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_809),
    .O(\DLX_IDinst_RegFile_21_18/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_13_27/LOGIC_ZERO_3207  (
    .O(\DLX_IDinst_RegFile_13_27/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_438_3208 (
    .IA(\DLX_IDinst_RegFile_13_27/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_13_27/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_497),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_438)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4971.INIT = 16'hF5DD;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4971 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_49),
    .ADR1(DLX_IDinst_RegFile_12_27),
    .ADR2(DLX_IDinst_RegFile_13_27),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_497)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_4981.INIT = 16'hE4FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_4981 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR1(DLX_IDinst_RegFile_14_27),
    .ADR2(DLX_IDinst_RegFile_15_27),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_50),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_498)
  );
  X_BUF \DLX_IDinst_RegFile_13_27/COUTUSED  (
    .I(\DLX_IDinst_RegFile_13_27/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_439)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_439_3209 (
    .IA(\DLX_IDinst_RegFile_13_27/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_438),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_498),
    .O(\DLX_IDinst_RegFile_13_27/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_13_27/CYINIT_3210  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_437),
    .O(\DLX_IDinst_RegFile_13_27/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_13_19/LOGIC_ZERO_3211  (
    .O(\DLX_IDinst_RegFile_13_19/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_822_3212 (
    .IA(\DLX_IDinst_RegFile_13_19/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_13_19/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_897),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_822)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8971.INIT = 16'hCFAF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8971 (
    .ADR0(DLX_IDinst_RegFile_12_19),
    .ADR1(DLX_IDinst_RegFile_13_19),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_577),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_897)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_8981.INIT = 16'hDF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_8981 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR1(DLX_IDinst_RegFile_15_19),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_578),
    .ADR3(DLX_IDinst_RegFile_14_19),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_898)
  );
  X_BUF \DLX_IDinst_RegFile_13_19/COUTUSED  (
    .I(\DLX_IDinst_RegFile_13_19/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_823)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_823_3213 (
    .IA(\DLX_IDinst_RegFile_13_19/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_822),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_898),
    .O(\DLX_IDinst_RegFile_13_19/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_13_19/CYINIT_3214  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_821),
    .O(\DLX_IDinst_RegFile_13_19/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_21_27/LOGIC_ZERO_3215  (
    .O(\DLX_IDinst_RegFile_21_27/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_442_3216 (
    .IA(\DLX_IDinst_RegFile_21_27/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_21_27/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_501),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_442)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5011.INIT = 16'hE4FF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5011 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR1(DLX_IDinst_RegFile_20_27),
    .ADR2(DLX_IDinst_RegFile_21_27),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_53),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_501)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5021.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5021 (
    .ADR0(DLX_IDinst_RegFile_22_27),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_54),
    .ADR2(DLX_IDinst_RegFile_23_27),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_502)
  );
  X_BUF \DLX_IDinst_RegFile_21_27/COUTUSED  (
    .I(\DLX_IDinst_RegFile_21_27/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_443)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_443_3217 (
    .IA(\DLX_IDinst_RegFile_21_27/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_442),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_502),
    .O(\DLX_IDinst_RegFile_21_27/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_21_27/CYINIT_3218  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_441),
    .O(\DLX_IDinst_RegFile_21_27/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_21_19/LOGIC_ZERO_3219  (
    .O(\DLX_IDinst_RegFile_21_19/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_826_3220 (
    .IA(\DLX_IDinst_RegFile_21_19/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_21_19/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_901),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_826)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9011.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9011 (
    .ADR0(DLX_IDinst_RegFile_21_19),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_581),
    .ADR2(DLX_IDinst_RegFile_20_19),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_901)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9021.INIT = 16'hB8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9021 (
    .ADR0(DLX_IDinst_RegFile_23_19),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_2 ),
    .ADR2(DLX_IDinst_RegFile_22_19),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_582),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_902)
  );
  X_BUF \DLX_IDinst_RegFile_21_19/COUTUSED  (
    .I(\DLX_IDinst_RegFile_21_19/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_827)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_827_3221 (
    .IA(\DLX_IDinst_RegFile_21_19/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_826),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_902),
    .O(\DLX_IDinst_RegFile_21_19/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_21_19/CYINIT_3222  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_825),
    .O(\DLX_IDinst_RegFile_21_19/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_13_28/LOGIC_ZERO_3223  (
    .O(\DLX_IDinst_RegFile_13_28/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_454_3224 (
    .IA(\DLX_IDinst_RegFile_13_28/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_13_28/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_513),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_454)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5131.INIT = 16'hF5DD;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5131 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_49),
    .ADR1(DLX_IDinst_RegFile_12_28),
    .ADR2(DLX_IDinst_RegFile_13_28),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_513)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5141.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5141 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR1(DLX_IDinst_RegFile_14_28),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_50),
    .ADR3(DLX_IDinst_RegFile_15_28),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_514)
  );
  X_BUF \DLX_IDinst_RegFile_13_28/COUTUSED  (
    .I(\DLX_IDinst_RegFile_13_28/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_455)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_455_3225 (
    .IA(\DLX_IDinst_RegFile_13_28/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_454),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_514),
    .O(\DLX_IDinst_RegFile_13_28/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_13_28/CYINIT_3226  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_453),
    .O(\DLX_IDinst_RegFile_13_28/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_21_28/LOGIC_ZERO_3227  (
    .O(\DLX_IDinst_RegFile_21_28/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_458_3228 (
    .IA(\DLX_IDinst_RegFile_21_28/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_21_28/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_517),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_458)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5171.INIT = 16'hEF4F;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5171 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR1(DLX_IDinst_RegFile_20_28),
    .ADR2(DLX_IDinst_Mmux__COND_4_inst_lut4_53),
    .ADR3(DLX_IDinst_RegFile_21_28),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_517)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5181.INIT = 16'hDFD5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5181 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_54),
    .ADR1(DLX_IDinst_RegFile_23_28),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_2 ),
    .ADR3(DLX_IDinst_RegFile_22_28),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_518)
  );
  X_BUF \DLX_IDinst_RegFile_21_28/COUTUSED  (
    .I(\DLX_IDinst_RegFile_21_28/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_459)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_459_3229 (
    .IA(\DLX_IDinst_RegFile_21_28/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_458),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_518),
    .O(\DLX_IDinst_RegFile_21_28/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_21_28/CYINIT_3230  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_457),
    .O(\DLX_IDinst_RegFile_21_28/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_13_29/LOGIC_ZERO_3231  (
    .O(\DLX_IDinst_RegFile_13_29/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_470_3232 (
    .IA(\DLX_IDinst_RegFile_13_29/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_13_29/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_529),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_470)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5291.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5291 (
    .ADR0(DLX_IDinst_RegFile_12_29),
    .ADR1(DLX_IDinst_Mmux__COND_4_inst_lut4_49),
    .ADR2(DLX_IDinst_RegFile_13_29),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_529)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5301.INIT = 16'hACFF;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5301 (
    .ADR0(DLX_IDinst_RegFile_15_29),
    .ADR1(DLX_IDinst_RegFile_14_29),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR3(DLX_IDinst_Mmux__COND_4_inst_lut4_50),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_530)
  );
  X_BUF \DLX_IDinst_RegFile_13_29/COUTUSED  (
    .I(\DLX_IDinst_RegFile_13_29/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_471)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_471_3233 (
    .IA(\DLX_IDinst_RegFile_13_29/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_470),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_530),
    .O(\DLX_IDinst_RegFile_13_29/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_13_29/CYINIT_3234  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_469),
    .O(\DLX_IDinst_RegFile_13_29/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_21_29/LOGIC_ZERO_3235  (
    .O(\DLX_IDinst_RegFile_21_29/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_474_3236 (
    .IA(\DLX_IDinst_RegFile_21_29/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_21_29/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_533),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_474)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5331.INIT = 16'hDFD5;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5331 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_53),
    .ADR1(DLX_IDinst_RegFile_21_29),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .ADR3(DLX_IDinst_RegFile_20_29),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_533)
  );
  defparam DLX_IDinst_Mmux__COND_4_inst_lut4_5341.INIT = 16'hF5DD;
  X_LUT4 DLX_IDinst_Mmux__COND_4_inst_lut4_5341 (
    .ADR0(DLX_IDinst_Mmux__COND_4_inst_lut4_54),
    .ADR1(DLX_IDinst_RegFile_22_29),
    .ADR2(DLX_IDinst_RegFile_23_29),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<16>1_1 ),
    .O(DLX_IDinst_Mmux__COND_4_inst_lut4_534)
  );
  X_BUF \DLX_IDinst_RegFile_21_29/COUTUSED  (
    .I(\DLX_IDinst_RegFile_21_29/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_4_inst_cy_475)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_4_inst_cy_475_3237 (
    .IA(\DLX_IDinst_RegFile_21_29/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_4_inst_cy_474),
    .SEL(DLX_IDinst_Mmux__COND_4_inst_lut4_534),
    .O(\DLX_IDinst_RegFile_21_29/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_21_29/CYINIT_3238  (
    .I(DLX_IDinst_Mmux__COND_4_inst_cy_473),
    .O(\DLX_IDinst_RegFile_21_29/CYINIT )
  );
  defparam DLX_IFinst_PC_27.INIT = 1'b0;
  X_SFF DLX_IFinst_PC_27 (
    .I(DLX_IFinst_NPC[27]),
    .CE(DLX_IFinst_PC_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_IFinst_PC[27])
  );
  X_ZERO \DLX_IDinst_RegFile_16_10/LOGIC_ZERO_3239  (
    .O(\DLX_IDinst_RegFile_16_10/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_680_3240 (
    .IA(\DLX_IDinst_RegFile_16_10/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_16_10/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_755),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_680)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7551.INIT = 16'hE2FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7551 (
    .ADR0(DLX_IDinst_RegFile_16_10),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR2(DLX_IDinst_RegFile_17_10),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_579),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_755)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7561.INIT = 16'hF3BB;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7561 (
    .ADR0(DLX_IDinst_RegFile_18_10),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_580),
    .ADR2(DLX_IDinst_RegFile_19_10),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_756)
  );
  X_BUF \DLX_IDinst_RegFile_16_10/COUTUSED  (
    .I(\DLX_IDinst_RegFile_16_10/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_681)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_681_3241 (
    .IA(\DLX_IDinst_RegFile_16_10/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_680),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_756),
    .O(\DLX_IDinst_RegFile_16_10/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_16_10/CYINIT_3242  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_679),
    .O(\DLX_IDinst_RegFile_16_10/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_24_10/LOGIC_ZERO_3243  (
    .O(\DLX_IDinst_RegFile_24_10/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_684_3244 (
    .IA(\DLX_IDinst_RegFile_24_10/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_24_10/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_759),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_684)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7591.INIT = 16'hBBF3;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7591 (
    .ADR0(DLX_IDinst_RegFile_25_10),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_583),
    .ADR2(DLX_IDinst_RegFile_24_10),
    .ADR3(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_759)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7601.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7601 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_584),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR2(DLX_IDinst_RegFile_26_10),
    .ADR3(DLX_IDinst_RegFile_27_10),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_760)
  );
  X_BUF \DLX_IDinst_RegFile_24_10/COUTUSED  (
    .I(\DLX_IDinst_RegFile_24_10/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_685)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_685_3245 (
    .IA(\DLX_IDinst_RegFile_24_10/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_684),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_760),
    .O(\DLX_IDinst_RegFile_24_10/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_24_10/CYINIT_3246  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_683),
    .O(\DLX_IDinst_RegFile_24_10/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_16_11/LOGIC_ZERO_3247  (
    .O(\DLX_IDinst_RegFile_16_11/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_696_3248 (
    .IA(\DLX_IDinst_RegFile_16_11/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_16_11/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_771),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_696)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7711.INIT = 16'hCAFF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7711 (
    .ADR0(DLX_IDinst_RegFile_16_11),
    .ADR1(DLX_IDinst_RegFile_17_11),
    .ADR2(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_579),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_771)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7721.INIT = 16'hDF8F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7721 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR1(DLX_IDinst_RegFile_19_11),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_580),
    .ADR3(DLX_IDinst_RegFile_18_11),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_772)
  );
  X_BUF \DLX_IDinst_RegFile_16_11/COUTUSED  (
    .I(\DLX_IDinst_RegFile_16_11/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_697)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_697_3249 (
    .IA(\DLX_IDinst_RegFile_16_11/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_696),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_772),
    .O(\DLX_IDinst_RegFile_16_11/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_16_11/CYINIT_3250  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_695),
    .O(\DLX_IDinst_RegFile_16_11/CYINIT )
  );
  defparam DLX_IFinst_IR_previous_20.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_20 (
    .I(DLX_IFinst_IR_latched[20]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[20])
  );
  X_ZERO \DLX_IDinst_RegFile_24_11/LOGIC_ZERO_3251  (
    .O(\DLX_IDinst_RegFile_24_11/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_700_3252 (
    .IA(\DLX_IDinst_RegFile_24_11/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_24_11/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_775),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_700)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7751.INIT = 16'hD8FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7751 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR1(DLX_IDinst_RegFile_25_11),
    .ADR2(DLX_IDinst_RegFile_24_11),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_583),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_775)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7761.INIT = 16'hFD75;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7761 (
    .ADR0(DLX_IDinst_Mmux__COND_5_inst_lut4_584),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR2(DLX_IDinst_RegFile_26_11),
    .ADR3(DLX_IDinst_RegFile_27_11),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_776)
  );
  X_BUF \DLX_IDinst_RegFile_24_11/COUTUSED  (
    .I(\DLX_IDinst_RegFile_24_11/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_701)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_701_3253 (
    .IA(\DLX_IDinst_RegFile_24_11/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_700),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_776),
    .O(\DLX_IDinst_RegFile_24_11/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_24_11/CYINIT_3254  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_699),
    .O(\DLX_IDinst_RegFile_24_11/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_16_20/LOGIC_ZERO_3255  (
    .O(\DLX_IDinst_RegFile_16_20/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_840_3256 (
    .IA(\DLX_IDinst_RegFile_16_20/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_16_20/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_915),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_840)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9151.INIT = 16'hEF2F;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9151 (
    .ADR0(DLX_IDinst_RegFile_16_20),
    .ADR1(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR2(DLX_IDinst_Mmux__COND_5_inst_lut4_579),
    .ADR3(DLX_IDinst_RegFile_17_20),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_915)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_9161.INIT = 16'hFB73;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_9161 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_1 ),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_580),
    .ADR2(DLX_IDinst_RegFile_18_20),
    .ADR3(DLX_IDinst_RegFile_19_20),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_916)
  );
  X_BUF \DLX_IDinst_RegFile_16_20/COUTUSED  (
    .I(\DLX_IDinst_RegFile_16_20/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_841)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_841_3257 (
    .IA(\DLX_IDinst_RegFile_16_20/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_840),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_916),
    .O(\DLX_IDinst_RegFile_16_20/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_16_20/CYINIT_3258  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_839),
    .O(\DLX_IDinst_RegFile_16_20/CYINIT )
  );
  X_ZERO \DLX_IDinst_RegFile_16_12/LOGIC_ZERO_3259  (
    .O(\DLX_IDinst_RegFile_16_12/LOGIC_ZERO )
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_712_3260 (
    .IA(\DLX_IDinst_RegFile_16_12/LOGIC_ZERO ),
    .IB(\DLX_IDinst_RegFile_16_12/CYINIT ),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_787),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_712)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7871.INIT = 16'hFB73;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7871 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR1(DLX_IDinst_Mmux__COND_5_inst_lut4_579),
    .ADR2(DLX_IDinst_RegFile_16_12),
    .ADR3(DLX_IDinst_RegFile_17_12),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_787)
  );
  defparam DLX_IDinst_Mmux__COND_5_inst_lut4_7881.INIT = 16'hE4FF;
  X_LUT4 DLX_IDinst_Mmux__COND_5_inst_lut4_7881 (
    .ADR0(\DLX_IDinst_Mmux_IR_latched_Result<21>1_3 ),
    .ADR1(DLX_IDinst_RegFile_18_12),
    .ADR2(DLX_IDinst_RegFile_19_12),
    .ADR3(DLX_IDinst_Mmux__COND_5_inst_lut4_580),
    .O(DLX_IDinst_Mmux__COND_5_inst_lut4_788)
  );
  X_BUF \DLX_IDinst_RegFile_16_12/COUTUSED  (
    .I(\DLX_IDinst_RegFile_16_12/CYMUXG ),
    .O(DLX_IDinst_Mmux__COND_5_inst_cy_713)
  );
  X_MUX2 DLX_IDinst_Mmux__COND_5_inst_cy_713_3261 (
    .IA(\DLX_IDinst_RegFile_16_12/LOGIC_ZERO ),
    .IB(DLX_IDinst_Mmux__COND_5_inst_cy_712),
    .SEL(DLX_IDinst_Mmux__COND_5_inst_lut4_788),
    .O(\DLX_IDinst_RegFile_16_12/CYMUXG )
  );
  X_BUF \DLX_IDinst_RegFile_16_12/CYINIT_3262  (
    .I(DLX_IDinst_Mmux__COND_5_inst_cy_711),
    .O(\DLX_IDinst_RegFile_16_12/CYINIT )
  );
  defparam DLX_IDinst_RegFile_2_19_3263.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_2_19_3263 (
    .I(DLX_IDinst_WB_data_eff[19]),
    .CE(DLX_IDinst__n0554),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_2_19)
  );
  defparam DLX_IFinst_IR_previous_16.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_16 (
    .I(DLX_IFinst_IR_latched[16]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[16])
  );
  defparam DLX_IDinst_RegFile_2_27_3264.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_2_27_3264 (
    .I(DLX_IDinst_WB_data_eff[27]),
    .CE(DLX_IDinst__n0554),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_2_27)
  );
  defparam DLX_IDinst_slot_num_FFd2_3265.INIT = 1'b0;
  X_SFF DLX_IDinst_slot_num_FFd2_3265 (
    .I(\DLX_IDinst_slot_num_FFd2-In ),
    .CE(DLX_IDinst__n0530),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_slot_num_FFd2)
  );
  defparam vga_top_vga1__n000839.INIT = 16'h8A00;
  X_LUT4 vga_top_vga1__n000839 (
    .ADR0(vga_top_vga1_hcounter[9]),
    .ADR1(CHOICE3146),
    .ADR2(vga_top_vga1_vcounter[9]),
    .ADR3(CHOICE3149),
    .O(\CHOICE3150/FROM )
  );
  defparam vga_top_vga1__n000846.INIT = 16'hAA00;
  X_LUT4 vga_top_vga1__n000846 (
    .ADR0(CHOICE3139),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(CHOICE3150),
    .O(\CHOICE3150/GROM )
  );
  X_BUF \CHOICE3150/XUSED  (
    .I(\CHOICE3150/FROM ),
    .O(CHOICE3150)
  );
  X_BUF \CHOICE3150/YUSED  (
    .I(\CHOICE3150/GROM ),
    .O(N145733)
  );
  defparam DLX_IDinst_slot_num_FFd3_3266.INIT = 1'b0;
  X_SFF DLX_IDinst_slot_num_FFd3_3266 (
    .I(\DLX_IDinst_slot_num_FFd3-In ),
    .CE(DLX_IDinst__n0530),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_slot_num_FFd3)
  );
  defparam DLX_IDinst_RegFile_2_21_3267.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_2_21_3267 (
    .I(DLX_IDinst_WB_data_eff[21]),
    .CE(DLX_IDinst__n0554),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_2_21)
  );
  defparam DLX_EXinst_noop_3268.INIT = 1'b1;
  X_SFF DLX_EXinst_noop_3268 (
    .I(\DLX_EXinst_noop/LOGIC_ZERO ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GSR),
    .RST(GND),
    .SSET(N139488),
    .SRST(GND),
    .O(DLX_EXinst_noop)
  );
  defparam DLX_IDinst_slot_num_FFd4_3269.INIT = 1'b1;
  X_SFF DLX_IDinst_slot_num_FFd4_3269 (
    .I(\DLX_IDinst_slot_num_FFd4-In ),
    .CE(DLX_IDinst__n0530),
    .CLK(clkdiv),
    .SET(GSR),
    .RST(GND),
    .SSET(reset_IBUF_3),
    .SRST(GND),
    .O(DLX_IDinst_slot_num_FFd4)
  );
  defparam DLX_IDinst_RegFile_2_13_3270.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_2_13_3270 (
    .I(DLX_IDinst_WB_data_eff[13]),
    .CE(DLX_IDinst__n0554),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_2_13)
  );
  defparam DLX_IDinst_RegFile_1_1_3271.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_1_1_3271 (
    .I(DLX_MEMinst_RF_data_in[1]),
    .CE(DLX_IDinst__n0552),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_1_1)
  );
  defparam DLX_EXinst_reg_out_B_EX_7.INIT = 1'b0;
  X_SFF DLX_EXinst_reg_out_B_EX_7 (
    .I(DLX_IDinst_reg_out_B[7]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_reg_out_B_EX[7])
  );
  defparam DLX_IDinst_RegFile_15_5_3272.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_15_5_3272 (
    .I(DLX_MEMinst_RF_data_in[5]),
    .CE(DLX_IDinst__n0580),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_15_5)
  );
  defparam DLX_IFinst_IR_previous_13.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_13 (
    .I(DLX_IFinst_IR_latched[13]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[13])
  );
  defparam DLX_IDinst_RegFile_1_23_3273.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_1_23_3273 (
    .I(DLX_IDinst_WB_data_eff[23]),
    .CE(DLX_IDinst__n0552),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_1_23)
  );
  defparam DLX_IDinst_RegFile_22_6_3274.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_22_6_3274 (
    .I(DLX_MEMinst_RF_data_in[6]),
    .CE(DLX_IDinst__n0594),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_22_6)
  );
  defparam DLX_MEMinst_opcode_of_WB_5.INIT = 1'b0;
  X_SFF DLX_MEMinst_opcode_of_WB_5 (
    .I(DLX_EXinst_opcode_of_EX_reg[5]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_MEMinst_opcode_of_WB[5])
  );
  defparam DLX_IDinst_RegFile_6_6_3275.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_6_6_3275 (
    .I(DLX_MEMinst_RF_data_in[6]),
    .CE(DLX_IDinst__n0562),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_6_6)
  );
  defparam DLX_IDinst_RegFile_15_9_3276.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_15_9_3276 (
    .I(DLX_IDinst_WB_data_eff[9]),
    .CE(DLX_IDinst__n0580),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_15_9)
  );
  defparam DLX_IDinst_RegFile_21_6_3277.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_21_6_3277 (
    .I(DLX_MEMinst_RF_data_in[6]),
    .CE(DLX_IDinst__n0592),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_21_6)
  );
  defparam DLX_IDinst_RegFile_22_2_3278.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_22_2_3278 (
    .I(DLX_MEMinst_RF_data_in[2]),
    .CE(DLX_IDinst__n0594),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_22_2)
  );
  defparam DLX_IDinst_RegFile_13_7_3279.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_13_7_3279 (
    .I(DLX_MEMinst_RF_data_in[7]),
    .CE(DLX_IDinst__n0576),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_13_7)
  );
  defparam DLX_IDinst_RegFile_30_2_3280.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_30_2_3280 (
    .I(DLX_MEMinst_RF_data_in[2]),
    .CE(DLX_IDinst__n0610),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_30_2)
  );
  defparam DLX_IDinst_RegFile_30_3_3281.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_30_3_3281 (
    .I(DLX_MEMinst_RF_data_in[3]),
    .CE(DLX_IDinst__n0610),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_30_3)
  );
  defparam DLX_IDinst_RegFile_14_3_3282.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_14_3_3282 (
    .I(DLX_MEMinst_RF_data_in[3]),
    .CE(DLX_IDinst__n0578),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_14_3)
  );
  defparam DLX_IDinst_RegFile_22_3_3283.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_22_3_3283 (
    .I(DLX_MEMinst_RF_data_in[3]),
    .CE(DLX_IDinst__n0594),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_22_3)
  );
  defparam DLX_IDinst_RegFile_21_7_3284.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_21_7_3284 (
    .I(DLX_MEMinst_RF_data_in[7]),
    .CE(DLX_IDinst__n0592),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_21_7)
  );
  defparam DLX_IDinst_reg_out_B_28.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_B_28 (
    .I(DLX_IDinst__n0147[28]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_B[28])
  );
  defparam DLX_IDinst_branch_address_29.INIT = 1'b0;
  X_SFF DLX_IDinst_branch_address_29 (
    .I(N141265),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_branch_address[29])
  );
  defparam DLX_IDinst_branch_address_28.INIT = 1'b0;
  X_SFF DLX_IDinst_branch_address_28 (
    .I(N141328),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_branch_address[28])
  );
  defparam DLX_IFinst_NPC_24.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_24 (
    .I(DLX_IFinst__n0001[24]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC[24])
  );
  defparam DLX_IFinst_NPC_16.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_16 (
    .I(DLX_IFinst__n0001[16]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC[16])
  );
  defparam DLX_IDinst_RegFile_0_7_3285.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_0_7_3285 (
    .I(DLX_MEMinst_RF_data_in[7]),
    .CE(DLX_IDinst__n0550),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_0_7)
  );
  defparam DLX_IFinst_NPC_25.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_25 (
    .I(DLX_IFinst__n0001[25]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC[25])
  );
  defparam DLX_IFinst_NPC_17.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_17 (
    .I(DLX_IFinst__n0001[17]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC[17])
  );
  defparam DLX_IFinst_NPC_26.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_26 (
    .I(DLX_IFinst__n0001[26]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC[26])
  );
  defparam DLX_IDinst_branch_address_23.INIT = 1'b0;
  X_SFF DLX_IDinst_branch_address_23 (
    .I(N141643),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_branch_address[23])
  );
  defparam DLX_IDinst_branch_address_31.INIT = 1'b0;
  X_SFF DLX_IDinst_branch_address_31 (
    .I(N145908),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_branch_address[31])
  );
  defparam DLX_IDinst_RegFile_3_29_3286.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_3_29_3286 (
    .I(DLX_IDinst_WB_data_eff[29]),
    .CE(DLX_IDinst__n0556),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_3_29)
  );
  defparam DLX_EXinst_ALU_result_0_1_3287.INIT = 1'b0;
  X_SFF DLX_EXinst_ALU_result_0_1_3287 (
    .I(\DLX_EXinst_ALU_result<0>/GROM ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE5945),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_ALU_result_0_1)
  );
  defparam DLX_EXinst_ALU_result_0.INIT = 1'b0;
  X_SFF DLX_EXinst_ALU_result_0 (
    .I(CHOICE6016),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE5945),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_ALU_result[0])
  );
  defparam DLX_IDinst_branch_address_17.INIT = 1'b0;
  X_SFF DLX_IDinst_branch_address_17 (
    .I(N140824),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_branch_address[17])
  );
  defparam DLX_IDinst_branch_address_24.INIT = 1'b0;
  X_SFF DLX_IDinst_branch_address_24 (
    .I(N141580),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_branch_address[24])
  );
  defparam DLX_IDinst_branch_address_25.INIT = 1'b0;
  X_SFF DLX_IDinst_branch_address_25 (
    .I(N141517),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_branch_address[25])
  );
  defparam DLX_IFinst_NPC_31.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_31 (
    .I(DLX_IFinst__n0001[31]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC[31])
  );
  defparam DLX_IFinst_NPC_15.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_15 (
    .I(\DLX_IFinst_NPC<15>/GROM ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC[15])
  );
  defparam DLX_IFinst_NPC_23.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_23 (
    .I(DLX_IFinst__n0001[23]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC[23])
  );
  defparam DLX_IDinst_branch_address_26.INIT = 1'b0;
  X_SFF DLX_IDinst_branch_address_26 (
    .I(N141454),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_branch_address[26])
  );
  defparam DLX_IDinst_branch_address_19.INIT = 1'b0;
  X_SFF DLX_IDinst_branch_address_19 (
    .I(N140950),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_branch_address[19])
  );
  defparam DLX_IDinst_branch_address_18.INIT = 1'b0;
  X_SFF DLX_IDinst_branch_address_18 (
    .I(N140887),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_branch_address[18])
  );
  defparam DLX_IDinst_branch_address_27.INIT = 1'b0;
  X_SFF DLX_IDinst_branch_address_27 (
    .I(N141391),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_branch_address[27])
  );
  defparam DLX_IFinst_NPC_18.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_18 (
    .I(DLX_IFinst__n0001[18]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC[18])
  );
  defparam DLX_IFinst_NPC_27.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_27 (
    .I(DLX_IFinst__n0001[27]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC[27])
  );
  defparam DLX_IFinst_NPC_19.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_19 (
    .I(DLX_IFinst__n0001[19]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC[19])
  );
  defparam DLX_MEMinst_opcode_of_WB_2.INIT = 1'b0;
  X_SFF DLX_MEMinst_opcode_of_WB_2 (
    .I(DLX_EXinst_opcode_of_EX_reg[2]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_MEMinst_opcode_of_WB[2])
  );
  defparam DLX_IFinst_NPC_29.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_29 (
    .I(DLX_IFinst__n0001[29]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC[29])
  );
  defparam DLX_IDinst_RegFile_20_2_3288.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_20_2_3288 (
    .I(DLX_MEMinst_RF_data_in[2]),
    .CE(DLX_IDinst__n0590),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_20_2)
  );
  defparam DLX_IDinst_RegFile_11_7_3289.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_11_7_3289 (
    .I(DLX_MEMinst_RF_data_in[7]),
    .CE(DLX_IDinst__n0572),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_11_7)
  );
  defparam DLX_IDinst_RegFile_20_3_3290.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_20_3_3290 (
    .I(DLX_MEMinst_RF_data_in[3]),
    .CE(DLX_IDinst__n0590),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_20_3)
  );
  defparam DLX_IDinst_RegFile_12_3_3291.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_12_3_3291 (
    .I(DLX_MEMinst_RF_data_in[3]),
    .CE(DLX_IDinst__n0574),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_12_3)
  );
  defparam DLX_IDinst_RegFile_20_4_3292.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_20_4_3292 (
    .I(DLX_MEMinst_RF_data_in[4]),
    .CE(DLX_IDinst__n0590),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_20_4)
  );
  defparam DLX_IDinst_RegFile_11_8_3293.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_11_8_3293 (
    .I(DLX_IDinst_WB_data_eff[8]),
    .CE(DLX_IDinst__n0572),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_11_8)
  );
  defparam DLX_IDinst_RegFile_13_0_3294.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_13_0_3294 (
    .I(DLX_MEMinst_RF_data_in[0]),
    .CE(DLX_IDinst__n0576),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_13_0)
  );
  defparam DLX_IDinst_RegFile_12_4_3295.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_12_4_3295 (
    .I(DLX_MEMinst_RF_data_in[4]),
    .CE(DLX_IDinst__n0574),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_12_4)
  );
  defparam DLX_IDinst_RegFile_2_16_3296.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_2_16_3296 (
    .I(DLX_IDinst_WB_data_eff[16]),
    .CE(DLX_IDinst__n0554),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_2_16)
  );
  defparam DLX_IDinst_RegFile_2_15_3297.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_2_15_3297 (
    .I(DLX_IDinst_WB_data_eff[15]),
    .CE(DLX_IDinst__n0554),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_2_15)
  );
  defparam DLX_IDinst_RegFile_0_12_3298.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_0_12_3298 (
    .I(DLX_IDinst_WB_data_eff[12]),
    .CE(DLX_IDinst__n0550),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_0_12)
  );
  defparam DLX_IDinst_RegFile_16_15_3299.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_16_15_3299 (
    .I(DLX_IDinst_WB_data_eff[15]),
    .CE(DLX_IDinst__n0582),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_16_15)
  );
  defparam DLX_IDinst_RegFile_2_17_3300.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_2_17_3300 (
    .I(DLX_IDinst_WB_data_eff[17]),
    .CE(DLX_IDinst__n0554),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_2_17)
  );
  defparam DLX_IFinst_IR_previous_6.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_6 (
    .I(DLX_IFinst_IR_latched[6]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[6])
  );
  defparam DLX_IDinst_RegFile_23_23_3301.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_23_23_3301 (
    .I(DLX_IDinst_WB_data_eff[23]),
    .CE(DLX_IDinst__n0596),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_23_23)
  );
  defparam DLX_IDinst_RegFile_30_23_3302.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_30_23_3302 (
    .I(DLX_IDinst_WB_data_eff[23]),
    .CE(DLX_IDinst__n0610),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_30_23)
  );
  defparam DLX_IDinst_RegFile_3_13_3303.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_3_13_3303 (
    .I(DLX_IDinst_WB_data_eff[13]),
    .CE(DLX_IDinst__n0556),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_3_13)
  );
  defparam DLX_IDinst_RegFile_2_29_3304.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_2_29_3304 (
    .I(DLX_IDinst_WB_data_eff[29]),
    .CE(DLX_IDinst__n0554),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_2_29)
  );
  defparam DLX_IDinst_RegFile_23_17_3305.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_23_17_3305 (
    .I(DLX_IDinst_WB_data_eff[17]),
    .CE(DLX_IDinst__n0596),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_23_17)
  );
  defparam DLX_IDinst_RegFile_3_31_3306.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_3_31_3306 (
    .I(DLX_IDinst_WB_data_eff[31]),
    .CE(DLX_IDinst__n0556),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_3_31)
  );
  defparam DLX_IDinst_RegFile_3_22_3307.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_3_22_3307 (
    .I(DLX_IDinst_WB_data_eff[22]),
    .CE(DLX_IDinst__n0556),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_3_22)
  );
  defparam DLX_IDinst_RegFile_18_4_3308.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_18_4_3308 (
    .I(DLX_MEMinst_RF_data_in[4]),
    .CE(DLX_IDinst__n0586),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_18_4)
  );
  defparam DLX_IDinst_RegFile_17_18_3309.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_17_18_3309 (
    .I(DLX_IDinst_WB_data_eff[18]),
    .CE(DLX_IDinst__n0584),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_17_18)
  );
  defparam DLX_IDinst_RegFile_29_7_3310.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_29_7_3310 (
    .I(DLX_MEMinst_RF_data_in[7]),
    .CE(DLX_IDinst__n0608),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_29_7)
  );
  defparam DLX_IDinst_RegFile_1_0_3311.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_1_0_3311 (
    .I(DLX_MEMinst_RF_data_in[0]),
    .CE(DLX_IDinst__n0552),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_1_0)
  );
  defparam DLX_IDinst_RegFile_3_25_3312.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_3_25_3312 (
    .I(DLX_IDinst_WB_data_eff[25]),
    .CE(DLX_IDinst__n0556),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_3_25)
  );
  defparam DLX_IDinst_RegFile_3_17_3313.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_3_17_3313 (
    .I(DLX_IDinst_WB_data_eff[17]),
    .CE(DLX_IDinst__n0556),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_3_17)
  );
  defparam DLX_IDinst_RegFile_3_20_3314.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_3_20_3314 (
    .I(DLX_IDinst_WB_data_eff[20]),
    .CE(DLX_IDinst__n0556),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_3_20)
  );
  defparam DLX_IDinst_RegFile_18_1_3315.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_18_1_3315 (
    .I(DLX_MEMinst_RF_data_in[1]),
    .CE(DLX_IDinst__n0586),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_18_1)
  );
  defparam DLX_IFinst_IR_previous_19.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_19 (
    .I(DLX_IFinst_IR_latched[19]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[19])
  );
  defparam DLX_MEMinst_reg_write_MEM_3316.INIT = 1'b0;
  X_SFF DLX_MEMinst_reg_write_MEM_3316 (
    .I(DLX_EXinst_reg_write_EX),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_MEMinst_reg_write_MEM)
  );
  defparam DLX_IDinst_branch_sig_3317.INIT = 1'b0;
  X_SFF DLX_IDinst_branch_sig_3317 (
    .I(\DLX_IDinst_branch_sig/GROM ),
    .CE(DLX_IDinst__n0116),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_IDinst__n0115),
    .O(DLX_IDinst_branch_sig)
  );
  defparam DLX_IDinst_RegFile_10_6_3318.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_10_6_3318 (
    .I(DLX_MEMinst_RF_data_in[6]),
    .CE(DLX_IDinst__n0570),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_10_6)
  );
  defparam DLX_IDinst_Imm_31_1_3319.INIT = 1'b0;
  X_SFF DLX_IDinst_Imm_31_1_3319 (
    .I(\DLX_IDinst_Imm<31>/GROM ),
    .CE(DLX_IDinst__n0116),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_IDinst__n0115),
    .O(DLX_IDinst_Imm_31_1)
  );
  defparam DLX_IDinst_Imm_31.INIT = 1'b0;
  X_SFF DLX_IDinst_Imm_31 (
    .I(N140698),
    .CE(DLX_IDinst__n0116),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_IDinst__n0115),
    .O(\DLX_IDinst_Imm[31] )
  );
  defparam DLX_IDinst_RegFile_11_2_3320.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_11_2_3320 (
    .I(DLX_MEMinst_RF_data_in[2]),
    .CE(DLX_IDinst__n0572),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_11_2)
  );
  defparam DLX_IFinst_IR_curr_30.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_30 (
    .I(IR_MSB_6_OBUF),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[30])
  );
  defparam DLX_IFinst_IR_curr_13.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_13 (
    .I(IR[13]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[13])
  );
  defparam DLX_IFinst_IR_curr_22.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_22 (
    .I(IR[22]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[22])
  );
  defparam DLX_IFinst_IR_curr_14.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_14 (
    .I(IR[14]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[14])
  );
  defparam DLX_IDinst_RegFile_1_5_3321.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_1_5_3321 (
    .I(DLX_MEMinst_RF_data_in[5]),
    .CE(DLX_IDinst__n0552),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_1_5)
  );
  defparam DLX_IDinst_RegFile_22_11_3322.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_22_11_3322 (
    .I(DLX_IDinst_WB_data_eff[11]),
    .CE(DLX_IDinst__n0594),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_22_11)
  );
  defparam DLX_IDinst_stall_3323.INIT = 1'b0;
  X_SFF DLX_IDinst_stall_3323 (
    .I(\DLX_IDinst_stall/GROM ),
    .CE(DLX_IDinst__n0614),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_stall)
  );
  defparam DLX_IFinst_IR_curr_28.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_28 (
    .I(IR_MSB_4_OBUF),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[28])
  );
  defparam DLX_IDinst_reg_out_A_30.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_A_30 (
    .I(N162964),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE2873),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_A[30])
  );
  defparam DLX_IFinst_IR_curr_29.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_29 (
    .I(IR_MSB_5_OBUF),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[29])
  );
  defparam DLX_IDinst_reg_out_B_0.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_B_0 (
    .I(DLX_IDinst__n0147[0]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_B[0])
  );
  defparam DLX_IDinst_slot_num_FFd1_3324.INIT = 1'b0;
  X_SFF DLX_IDinst_slot_num_FFd1_3324 (
    .I(\DLX_IDinst_slot_num_FFd1-In ),
    .CE(DLX_IDinst__n0530),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_slot_num_FFd1)
  );
  defparam DLX_IDinst_RegFile_3_19_3325.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_3_19_3325 (
    .I(DLX_IDinst_WB_data_eff[19]),
    .CE(DLX_IDinst__n0556),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_3_19)
  );
  defparam DLX_IDinst_RegFile_2_5_3326.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_2_5_3326 (
    .I(DLX_MEMinst_RF_data_in[5]),
    .CE(DLX_IDinst__n0554),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_2_5)
  );
  defparam DLX_IDinst_RegFile_3_10_3327.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_3_10_3327 (
    .I(DLX_IDinst_WB_data_eff[10]),
    .CE(DLX_IDinst__n0556),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_3_10)
  );
  defparam DLX_IDinst_RegFile_27_25_3328.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_27_25_3328 (
    .I(DLX_IDinst_WB_data_eff[25]),
    .CE(DLX_IDinst__n0604),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_27_25)
  );
  defparam DLX_IDinst_RegFile_3_1_3329.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_3_1_3329 (
    .I(DLX_MEMinst_RF_data_in[1]),
    .CE(DLX_IDinst__n0556),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_3_1)
  );
  defparam DLX_EXinst_ALU_result_20.INIT = 1'b0;
  X_SFF DLX_EXinst_ALU_result_20 (
    .I(N162820),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE4700),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_ALU_result[20])
  );
  defparam DLX_IDinst_RegFile_3_27_3330.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_3_27_3330 (
    .I(DLX_IDinst_WB_data_eff[27]),
    .CE(DLX_IDinst__n0556),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_3_27)
  );
  defparam DLX_EXinst_ALU_result_21.INIT = 1'b0;
  X_SFF DLX_EXinst_ALU_result_21 (
    .I(CHOICE4185),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE4153),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_ALU_result[21])
  );
  defparam DLX_IDinst_RegFile_7_4_3331.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_7_4_3331 (
    .I(DLX_MEMinst_RF_data_in[4]),
    .CE(DLX_IDinst__n0564),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_7_4)
  );
  defparam DLX_IDinst_RegFile_1_9_3332.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_1_9_3332 (
    .I(DLX_IDinst_WB_data_eff[9]),
    .CE(DLX_IDinst__n0552),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_1_9)
  );
  defparam DLX_IDinst_RegFile_3_11_3333.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_3_11_3333 (
    .I(DLX_IDinst_WB_data_eff[11]),
    .CE(DLX_IDinst__n0556),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_3_11)
  );
  defparam DLX_EXinst_ALU_result_23.INIT = 1'b0;
  X_SFF DLX_EXinst_ALU_result_23 (
    .I(CHOICE4055),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE4023),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_ALU_result[23])
  );
  defparam DLX_IDinst_RegFile_22_8_3334.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_22_8_3334 (
    .I(DLX_IDinst_WB_data_eff[8]),
    .CE(DLX_IDinst__n0594),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_22_8)
  );
  defparam DLX_EXinst_ALU_result_30.INIT = 1'b0;
  X_SFF DLX_EXinst_ALU_result_30 (
    .I(N162838),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE4734),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_ALU_result[30])
  );
  defparam DLX_EXinst_ALU_result_22.INIT = 1'b0;
  X_SFF DLX_EXinst_ALU_result_22 (
    .I(CHOICE4120),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE4088),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_ALU_result[22])
  );
  defparam DLX_IDinst_RegFile_15_7_3335.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_15_7_3335 (
    .I(DLX_MEMinst_RF_data_in[7]),
    .CE(DLX_IDinst__n0580),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_15_7)
  );
  defparam DLX_IDinst_RegFile_23_8_3336.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_23_8_3336 (
    .I(DLX_IDinst_WB_data_eff[8]),
    .CE(DLX_IDinst__n0596),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_23_8)
  );
  defparam DLX_EXinst_ALU_result_16.INIT = 1'b0;
  X_SFF DLX_EXinst_ALU_result_16 (
    .I(CHOICE4629),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE4594),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_ALU_result[16])
  );
  defparam DLX_IDinst_RegFile_7_3_3337.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_7_3_3337 (
    .I(DLX_MEMinst_RF_data_in[3]),
    .CE(DLX_IDinst__n0564),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_7_3)
  );
  defparam DLX_IDinst_RegFile_22_16_3338.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_22_16_3338 (
    .I(DLX_IDinst_WB_data_eff[16]),
    .CE(DLX_IDinst__n0594),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_22_16)
  );
  defparam DLX_EXinst_ALU_result_24.INIT = 1'b0;
  X_SFF DLX_EXinst_ALU_result_24 (
    .I(CHOICE5683),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE5634),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_ALU_result[24])
  );
  defparam DLX_IDinst_RegFile_2_7_3339.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_2_7_3339 (
    .I(DLX_MEMinst_RF_data_in[7]),
    .CE(DLX_IDinst__n0554),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_2_7)
  );
  defparam DLX_EXinst_ALU_result_25.INIT = 1'b0;
  X_SFF DLX_EXinst_ALU_result_25 (
    .I(CHOICE5120),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE5087),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_ALU_result[25])
  );
  defparam DLX_EXinst_ALU_result_17.INIT = 1'b0;
  X_SFF DLX_EXinst_ALU_result_17 (
    .I(CHOICE5428),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE5389),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_ALU_result[17])
  );
  defparam DLX_IDinst_RegFile_3_4_3340.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_3_4_3340 (
    .I(DLX_MEMinst_RF_data_in[4]),
    .CE(DLX_IDinst__n0556),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_3_4)
  );
  defparam DLX_EXinst_ALU_result_26.INIT = 1'b0;
  X_SFF DLX_EXinst_ALU_result_26 (
    .I(CHOICE5053),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE5020),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_ALU_result[26])
  );
  defparam DLX_EXinst_ALU_result_18.INIT = 1'b0;
  X_SFF DLX_EXinst_ALU_result_18 (
    .I(CHOICE5270),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE5231),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_ALU_result[18])
  );
  defparam DLX_EXinst_ALU_result_27.INIT = 1'b0;
  X_SFF DLX_EXinst_ALU_result_27 (
    .I(CHOICE4986),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE4953),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_ALU_result[27])
  );
  defparam DLX_EXinst_ALU_result_19.INIT = 1'b0;
  X_SFF DLX_EXinst_ALU_result_19 (
    .I(CHOICE5349),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE5310),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_ALU_result[19])
  );
  defparam DLX_EXinst_ALU_result_28.INIT = 1'b0;
  X_SFF DLX_EXinst_ALU_result_28 (
    .I(N162804),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE4879),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_ALU_result[28])
  );
  defparam DLX_IFinst_IR_previous_30.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_30 (
    .I(DLX_IFinst_IR_latched[30]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[30])
  );
  defparam DLX_IDinst_RegFile_3_9_3341.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_3_9_3341 (
    .I(DLX_IDinst_WB_data_eff[9]),
    .CE(DLX_IDinst__n0556),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_3_9)
  );
  defparam DLX_IDinst_RegFile_5_0_3342.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_5_0_3342 (
    .I(DLX_MEMinst_RF_data_in[0]),
    .CE(DLX_IDinst__n0560),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_5_0)
  );
  defparam DLX_IFinst_NPC_0.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_0 (
    .I(\DLX_IFinst_NPC<0>/GROM ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC[0])
  );
  defparam DLX_IDinst_RegFile_4_5_3343.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_4_5_3343 (
    .I(DLX_MEMinst_RF_data_in[5]),
    .CE(DLX_IDinst__n0558),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_4_5)
  );
  defparam DLX_IDinst_RegFile_5_1_3344.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_5_1_3344 (
    .I(DLX_MEMinst_RF_data_in[1]),
    .CE(DLX_IDinst__n0560),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_5_1)
  );
  defparam DLX_IDinst_EPC_6.INIT = 1'b0;
  X_SFF DLX_IDinst_EPC_6 (
    .I(DLX_IFinst_NPC[6]),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_EPC[6])
  );
  defparam DLX_IDinst_RegFile_0_1_3345.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_0_1_3345 (
    .I(DLX_MEMinst_RF_data_in[1]),
    .CE(DLX_IDinst__n0550),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_0_1)
  );
  defparam DLX_IDinst_RegFile_0_0_3346.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_0_0_3346 (
    .I(DLX_MEMinst_RF_data_in[0]),
    .CE(DLX_IDinst__n0550),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_0_0)
  );
  defparam DLX_IDinst_RegFile_1_17_3347.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_1_17_3347 (
    .I(DLX_IDinst_WB_data_eff[17]),
    .CE(DLX_IDinst__n0552),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_1_17)
  );
  defparam DLX_EXinst_ALU_result_29.INIT = 1'b0;
  X_SFF DLX_EXinst_ALU_result_29 (
    .I(N162835),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE4805),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_ALU_result[29])
  );
  defparam DLX_IDinst_RegFile_27_29_3348.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_27_29_3348 (
    .I(DLX_IDinst_WB_data_eff[29]),
    .CE(DLX_IDinst__n0604),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_27_29)
  );
  defparam DLX_IDinst_RegFile_23_26_3349.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_23_26_3349 (
    .I(DLX_IDinst_WB_data_eff[26]),
    .CE(DLX_IDinst__n0596),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_23_26)
  );
  defparam DLX_IDinst_RegFile_16_13_3350.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_16_13_3350 (
    .I(DLX_IDinst_WB_data_eff[13]),
    .CE(DLX_IDinst__n0582),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_16_13)
  );
  defparam DLX_IDinst_RegFile_0_2_3351.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_0_2_3351 (
    .I(DLX_MEMinst_RF_data_in[2]),
    .CE(DLX_IDinst__n0550),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_0_2)
  );
  defparam DLX_IDinst_RegFile_0_4_3352.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_0_4_3352 (
    .I(DLX_MEMinst_RF_data_in[4]),
    .CE(DLX_IDinst__n0550),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_0_4)
  );
  defparam DLX_IDinst_RegFile_1_2_3353.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_1_2_3353 (
    .I(DLX_MEMinst_RF_data_in[2]),
    .CE(DLX_IDinst__n0552),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_1_2)
  );
  defparam DLX_IDinst_RegFile_1_3_3354.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_1_3_3354 (
    .I(DLX_MEMinst_RF_data_in[3]),
    .CE(DLX_IDinst__n0552),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_1_3)
  );
  defparam DLX_IDinst_RegFile_4_0_3355.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_4_0_3355 (
    .I(DLX_MEMinst_RF_data_in[0]),
    .CE(DLX_IDinst__n0558),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_4_0)
  );
  defparam DLX_IDinst_RegFile_4_1_3356.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_4_1_3356 (
    .I(DLX_MEMinst_RF_data_in[1]),
    .CE(DLX_IDinst__n0558),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_4_1)
  );
  defparam DLX_IDinst_RegFile_4_2_3357.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_4_2_3357 (
    .I(DLX_MEMinst_RF_data_in[2]),
    .CE(DLX_IDinst__n0558),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_4_2)
  );
  defparam DLX_IDinst_RegFile_4_3_3358.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_4_3_3358 (
    .I(DLX_MEMinst_RF_data_in[3]),
    .CE(DLX_IDinst__n0558),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_4_3)
  );
  defparam DLX_IDinst_RegFile_4_4_3359.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_4_4_3359 (
    .I(DLX_MEMinst_RF_data_in[4]),
    .CE(DLX_IDinst__n0558),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_4_4)
  );
  defparam DLX_IDinst_RegFile_3_7_3360.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_3_7_3360 (
    .I(DLX_MEMinst_RF_data_in[7]),
    .CE(DLX_IDinst__n0556),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_3_7)
  );
  defparam DLX_IDinst_RegFile_6_1_3361.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_6_1_3361 (
    .I(DLX_MEMinst_RF_data_in[1]),
    .CE(DLX_IDinst__n0562),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_6_1)
  );
  defparam DLX_IDinst_RegFile_5_5_3362.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_5_5_3362 (
    .I(DLX_MEMinst_RF_data_in[5]),
    .CE(DLX_IDinst__n0560),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_5_5)
  );
  defparam DLX_IDinst_RegFile_4_9_3363.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_4_9_3363 (
    .I(DLX_IDinst_WB_data_eff[9]),
    .CE(DLX_IDinst__n0558),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_4_9)
  );
  defparam DLX_IDinst_RegFile_5_7_3364.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_5_7_3364 (
    .I(DLX_MEMinst_RF_data_in[7]),
    .CE(DLX_IDinst__n0560),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_5_7)
  );
  defparam DLX_IDinst_RegFile_6_2_3365.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_6_2_3365 (
    .I(DLX_MEMinst_RF_data_in[2]),
    .CE(DLX_IDinst__n0562),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_6_2)
  );
  defparam DLX_IDinst_RegFile_6_3_3366.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_6_3_3366 (
    .I(DLX_MEMinst_RF_data_in[3]),
    .CE(DLX_IDinst__n0562),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_6_3)
  );
  defparam DLX_IDinst_RegFile_5_6_3367.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_5_6_3367 (
    .I(DLX_MEMinst_RF_data_in[6]),
    .CE(DLX_IDinst__n0560),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_5_6)
  );
  defparam DLX_IDinst_RegFile_6_7_3368.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_6_7_3368 (
    .I(DLX_MEMinst_RF_data_in[7]),
    .CE(DLX_IDinst__n0562),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_6_7)
  );
  defparam DLX_IDinst_RegFile_6_5_3369.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_6_5_3369 (
    .I(DLX_MEMinst_RF_data_in[5]),
    .CE(DLX_IDinst__n0562),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_6_5)
  );
  defparam DLX_IDinst_RegFile_6_4_3370.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_6_4_3370 (
    .I(DLX_MEMinst_RF_data_in[4]),
    .CE(DLX_IDinst__n0562),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_6_4)
  );
  defparam DLX_IDinst_RegFile_5_8_3371.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_5_8_3371 (
    .I(DLX_IDinst_WB_data_eff[8]),
    .CE(DLX_IDinst__n0560),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_5_8)
  );
  defparam DLX_IDinst_RegFile_7_0_3372.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_7_0_3372 (
    .I(DLX_MEMinst_RF_data_in[0]),
    .CE(DLX_IDinst__n0564),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_7_0)
  );
  defparam DLX_IDinst_RegFile_5_9_3373.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_5_9_3373 (
    .I(DLX_IDinst_WB_data_eff[9]),
    .CE(DLX_IDinst__n0560),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_5_9)
  );
  defparam DLX_IDinst_RegFile_7_1_3374.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_7_1_3374 (
    .I(DLX_MEMinst_RF_data_in[1]),
    .CE(DLX_IDinst__n0564),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_7_1)
  );
  defparam DLX_IDinst_RegFile_7_6_3375.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_7_6_3375 (
    .I(DLX_MEMinst_RF_data_in[6]),
    .CE(DLX_IDinst__n0564),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_7_6)
  );
  defparam DLX_IDinst_RegFile_8_0_3376.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_8_0_3376 (
    .I(DLX_MEMinst_RF_data_in[0]),
    .CE(DLX_IDinst__n0566),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_8_0)
  );
  defparam DLX_IDinst_RegFile_6_8_3377.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_6_8_3377 (
    .I(DLX_IDinst_WB_data_eff[8]),
    .CE(DLX_IDinst__n0562),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_6_8)
  );
  defparam DLX_IDinst_RegFile_8_1_3378.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_8_1_3378 (
    .I(DLX_MEMinst_RF_data_in[1]),
    .CE(DLX_IDinst__n0566),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_8_1)
  );
  defparam DLX_IDinst_RegFile_8_2_3379.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_8_2_3379 (
    .I(DLX_MEMinst_RF_data_in[2]),
    .CE(DLX_IDinst__n0566),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_8_2)
  );
  defparam DLX_IDinst_RegFile_7_7_3380.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_7_7_3380 (
    .I(DLX_MEMinst_RF_data_in[7]),
    .CE(DLX_IDinst__n0564),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_7_7)
  );
  defparam DLX_IDinst_RegFile_7_8_3381.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_7_8_3381 (
    .I(DLX_IDinst_WB_data_eff[8]),
    .CE(DLX_IDinst__n0564),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_7_8)
  );
  defparam DLX_IDinst_RegFile_8_3_3382.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_8_3_3382 (
    .I(DLX_MEMinst_RF_data_in[3]),
    .CE(DLX_IDinst__n0566),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_8_3)
  );
  defparam DLX_IDinst_RegFile_9_0_3383.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_9_0_3383 (
    .I(DLX_MEMinst_RF_data_in[0]),
    .CE(DLX_IDinst__n0568),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_9_0)
  );
  defparam DLX_IDinst_RegFile_7_9_3384.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_7_9_3384 (
    .I(DLX_IDinst_WB_data_eff[9]),
    .CE(DLX_IDinst__n0564),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_7_9)
  );
  defparam DLX_IDinst_RegFile_8_4_3385.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_8_4_3385 (
    .I(DLX_MEMinst_RF_data_in[4]),
    .CE(DLX_IDinst__n0566),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_8_4)
  );
  defparam DLX_IDinst_RegFile_4_6_3386.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_4_6_3386 (
    .I(DLX_MEMinst_RF_data_in[6]),
    .CE(DLX_IDinst__n0558),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_4_6)
  );
  defparam DLX_IDinst_RegFile_5_2_3387.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_5_2_3387 (
    .I(DLX_MEMinst_RF_data_in[2]),
    .CE(DLX_IDinst__n0560),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_5_2)
  );
  defparam DLX_IDinst_RegFile_4_7_3388.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_4_7_3388 (
    .I(DLX_MEMinst_RF_data_in[7]),
    .CE(DLX_IDinst__n0558),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_4_7)
  );
  defparam DLX_IDinst_RegFile_5_3_3389.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_5_3_3389 (
    .I(DLX_MEMinst_RF_data_in[3]),
    .CE(DLX_IDinst__n0560),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_5_3)
  );
  defparam DLX_IDinst_RegFile_4_8_3390.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_4_8_3390 (
    .I(DLX_IDinst_WB_data_eff[8]),
    .CE(DLX_IDinst__n0558),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_4_8)
  );
  defparam DLX_IDinst_RegFile_5_4_3391.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_5_4_3391 (
    .I(DLX_MEMinst_RF_data_in[4]),
    .CE(DLX_IDinst__n0560),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_5_4)
  );
  defparam DLX_IDinst_RegFile_6_0_3392.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_6_0_3392 (
    .I(DLX_MEMinst_RF_data_in[0]),
    .CE(DLX_IDinst__n0562),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_6_0)
  );
  defparam DLX_IDinst_RegFile_8_5_3393.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_8_5_3393 (
    .I(DLX_MEMinst_RF_data_in[5]),
    .CE(DLX_IDinst__n0566),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_8_5)
  );
  defparam DLX_IDinst_RegFile_9_1_3394.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_9_1_3394 (
    .I(DLX_MEMinst_RF_data_in[1]),
    .CE(DLX_IDinst__n0568),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_9_1)
  );
  defparam DLX_IDinst_RegFile_8_6_3395.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_8_6_3395 (
    .I(DLX_MEMinst_RF_data_in[6]),
    .CE(DLX_IDinst__n0566),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_8_6)
  );
  defparam DLX_IDinst_RegFile_9_2_3396.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_9_2_3396 (
    .I(DLX_MEMinst_RF_data_in[2]),
    .CE(DLX_IDinst__n0568),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_9_2)
  );
  defparam DLX_IDinst_RegFile_9_3_3397.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_9_3_3397 (
    .I(DLX_MEMinst_RF_data_in[3]),
    .CE(DLX_IDinst__n0568),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_9_3)
  );
  defparam DLX_IDinst_RegFile_8_7_3398.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_8_7_3398 (
    .I(DLX_MEMinst_RF_data_in[7]),
    .CE(DLX_IDinst__n0566),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_8_7)
  );
  defparam DLX_IDinst_RegFile_8_8_3399.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_8_8_3399 (
    .I(DLX_IDinst_WB_data_eff[8]),
    .CE(DLX_IDinst__n0566),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_8_8)
  );
  defparam DLX_IDinst_RegFile_9_4_3400.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_9_4_3400 (
    .I(DLX_MEMinst_RF_data_in[4]),
    .CE(DLX_IDinst__n0568),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_9_4)
  );
  defparam DLX_IDinst_RegFile_8_9_3401.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_8_9_3401 (
    .I(DLX_IDinst_WB_data_eff[9]),
    .CE(DLX_IDinst__n0566),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_8_9)
  );
  defparam DLX_IDinst_RegFile_9_7_3402.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_9_7_3402 (
    .I(DLX_MEMinst_RF_data_in[7]),
    .CE(DLX_IDinst__n0568),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_9_7)
  );
  defparam DLX_IDinst_RegFile_9_5_3403.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_9_5_3403 (
    .I(DLX_MEMinst_RF_data_in[5]),
    .CE(DLX_IDinst__n0568),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_9_5)
  );
  defparam DLX_IDinst_RegFile_9_6_3404.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_9_6_3404 (
    .I(DLX_MEMinst_RF_data_in[6]),
    .CE(DLX_IDinst__n0568),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_9_6)
  );
  defparam DLX_IDinst_RegFile_9_8_3405.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_9_8_3405 (
    .I(DLX_IDinst_WB_data_eff[8]),
    .CE(DLX_IDinst__n0568),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_9_8)
  );
  defparam DLX_IDinst_RegFile_9_9_3406.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_9_9_3406 (
    .I(DLX_IDinst_WB_data_eff[9]),
    .CE(DLX_IDinst__n0568),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_9_9)
  );
  defparam DLX_IFinst_NPC_1.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_1 (
    .I(\DLX_IFinst_NPC<1>/GROM ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC[1])
  );
  defparam DLX_IFinst_NPC_2.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_2 (
    .I(\DLX_IFinst_NPC<2>/GROM ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC[2])
  );
  defparam DLX_IDinst_RegFile_11_14_3407.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_11_14_3407 (
    .I(DLX_IDinst_WB_data_eff[14]),
    .CE(DLX_IDinst__n0572),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_11_14)
  );
  defparam DLX_IDinst_RegFile_11_26_3408.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_11_26_3408 (
    .I(DLX_IDinst_WB_data_eff[26]),
    .CE(DLX_IDinst__n0572),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_11_26)
  );
  defparam DLX_IDinst_RegFile_11_28_3409.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_11_28_3409 (
    .I(DLX_IDinst_WB_data_eff[28]),
    .CE(DLX_IDinst__n0572),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_11_28)
  );
  defparam DLX_IDinst_RegFile_7_2_3410.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_7_2_3410 (
    .I(DLX_MEMinst_RF_data_in[2]),
    .CE(DLX_IDinst__n0564),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_7_2)
  );
  defparam DLX_IDinst_EPC_2.INIT = 1'b0;
  X_SFF DLX_IDinst_EPC_2 (
    .I(DLX_IFinst_NPC[2]),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_EPC[2])
  );
  defparam DLX_IDinst_RegFile_2_0_3411.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_2_0_3411 (
    .I(DLX_MEMinst_RF_data_in[0]),
    .CE(DLX_IDinst__n0554),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_2_0)
  );
  defparam DLX_IDinst_EPC_3.INIT = 1'b0;
  X_SFF DLX_IDinst_EPC_3 (
    .I(DLX_IFinst_NPC[3]),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_EPC[3])
  );
  defparam DLX_IFinst_NPC_3.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_3 (
    .I(\DLX_IFinst_NPC<3>/GROM ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC[3])
  );
  defparam DLX_IFinst_NPC_4.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_4 (
    .I(\DLX_IFinst_NPC<4>/GROM ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC[4])
  );
  defparam DLX_IFinst_NPC_5.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_5 (
    .I(\DLX_IFinst_NPC<5>/GROM ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC[5])
  );
  defparam DLX_IFinst_NPC_6.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_6 (
    .I(\DLX_IFinst_NPC<6>/GROM ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC[6])
  );
  defparam DLX_IFinst_NPC_7.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_7 (
    .I(\DLX_IFinst_NPC<7>/GROM ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC[7])
  );
  defparam DLX_IFinst_NPC_8.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_8 (
    .I(\DLX_IFinst_NPC<8>/GROM ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC[8])
  );
  defparam DLX_IFinst_NPC_9.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_9 (
    .I(\DLX_IFinst_NPC<9>/GROM ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC[9])
  );
  defparam DLX_IFinst_IR_curr_7.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_7 (
    .I(IR[7]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[7])
  );
  defparam DLX_IDinst_RegFile_6_16_3412.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_6_16_3412 (
    .I(DLX_IDinst_WB_data_eff[16]),
    .CE(DLX_IDinst__n0562),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_6_16)
  );
  defparam DLX_IDinst_EPC_4.INIT = 1'b0;
  X_SFF DLX_IDinst_EPC_4 (
    .I(DLX_IFinst_NPC[4]),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_EPC[4])
  );
  defparam DLX_IDinst_EPC_5.INIT = 1'b0;
  X_SFF DLX_IDinst_EPC_5 (
    .I(DLX_IFinst_NPC[5]),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_EPC[5])
  );
  defparam DLX_IFinst_PC_10.INIT = 1'b0;
  X_SFF DLX_IFinst_PC_10 (
    .I(DLX_IFinst_NPC[10]),
    .CE(DLX_IFinst_PC_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_PC[10])
  );
  defparam DLX_IDinst_RegFile_6_23_3413.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_6_23_3413 (
    .I(DLX_IDinst_WB_data_eff[23]),
    .CE(DLX_IDinst__n0562),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_6_23)
  );
  defparam DLX_IDinst_RegFile_6_19_3414.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_6_19_3414 (
    .I(DLX_IDinst_WB_data_eff[19]),
    .CE(DLX_IDinst__n0562),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_6_19)
  );
  defparam vga_top_vga1_helpme_3415.INIT = 1'b1;
  X_SFF vga_top_vga1_helpme_3415 (
    .I(\vga_top_vga1_helpme/LOGIC_ZERO ),
    .CE(vga_top_vga1__n0052),
    .CLK(clkdiv),
    .SET(GSR),
    .RST(GND),
    .SSET(reset_IBUF_1),
    .SRST(GND),
    .O(vga_top_vga1_helpme)
  );
  defparam DLX_IDinst_Cause_Reg_0.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_0 (
    .I(DLX_IDinst_Imm_0_1),
    .CE(DLX_IDinst__n0617),
    .CLK(clkdiv),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<0>/FFY/RST ),
    .O(\DLX_IDinst_Cause_Reg[0] )
  );
  X_BUF \DLX_IDinst_Cause_Reg<0>/FFY/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<0>/FFY/RST )
  );
  defparam DLX_IDinst_Cause_Reg_1.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_1 (
    .I(DLX_IDinst_Imm_1_1),
    .CE(DLX_IDinst__n0617),
    .CLK(clkdiv),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<1>/FFY/RST ),
    .O(\DLX_IDinst_Cause_Reg[1] )
  );
  X_BUF \DLX_IDinst_Cause_Reg<1>/FFY/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<1>/FFY/RST )
  );
  defparam DLX_IDinst_Cause_Reg_3.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_3 (
    .I(DLX_IDinst_Imm_3_1),
    .CE(DLX_IDinst__n0617),
    .CLK(clkdiv),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<3>/FFY/RST ),
    .O(\DLX_IDinst_Cause_Reg[3] )
  );
  X_BUF \DLX_IDinst_Cause_Reg<3>/FFY/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<3>/FFY/RST )
  );
  defparam DLX_IDinst_Cause_Reg_2.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_2 (
    .I(DLX_IDinst_Imm_2_1),
    .CE(DLX_IDinst__n0617),
    .CLK(clkdiv),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<2>/FFY/RST ),
    .O(\DLX_IDinst_Cause_Reg[2] )
  );
  X_BUF \DLX_IDinst_Cause_Reg<2>/FFY/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<2>/FFY/RST )
  );
  defparam DLX_IDinst_Cause_Reg_4.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_4 (
    .I(\DLX_IDinst_Imm[4] ),
    .CE(DLX_IDinst__n0617),
    .CLK(clkdiv),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<4>/FFY/RST ),
    .O(\DLX_IDinst_Cause_Reg[4] )
  );
  X_BUF \DLX_IDinst_Cause_Reg<4>/FFY/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<4>/FFY/RST )
  );
  defparam DLX_IDinst_Cause_Reg_5.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_5 (
    .I(\DLX_IDinst_Imm[5] ),
    .CE(DLX_IDinst__n0617),
    .CLK(clkdiv),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<5>/FFY/RST ),
    .O(\DLX_IDinst_Cause_Reg[5] )
  );
  X_BUF \DLX_IDinst_Cause_Reg<5>/FFY/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<5>/FFY/RST )
  );
  defparam DLX_IDinst_branch_address_21.INIT = 1'b0;
  X_SFF DLX_IDinst_branch_address_21 (
    .I(N141076),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_branch_address[21])
  );
  defparam DLX_IFinst_NPC_30.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_30 (
    .I(DLX_IFinst__n0001[30]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC[30])
  );
  defparam DLX_IFinst_NPC_14.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_14 (
    .I(\DLX_IFinst_NPC<14>/GROM ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC[14])
  );
  defparam DLX_IFinst_NPC_22.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_22 (
    .I(DLX_IFinst__n0001[22]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC[22])
  );
  defparam DLX_IDinst_branch_address_22.INIT = 1'b0;
  X_SFF DLX_IDinst_branch_address_22 (
    .I(N141139),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_branch_address[22])
  );
  defparam DLX_IDinst_branch_address_30.INIT = 1'b0;
  X_SFF DLX_IDinst_branch_address_30 (
    .I(N141202),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_branch_address[30])
  );
  defparam DLX_IDinst_branch_address_14.INIT = 1'b0;
  X_SFF DLX_IDinst_branch_address_14 (
    .I(N140571),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_branch_address[14])
  );
  defparam DLX_IDinst_branch_address_15.INIT = 1'b0;
  X_SFF DLX_IDinst_branch_address_15 (
    .I(N140634),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_branch_address[15])
  );
  defparam DLX_IDinst_Cause_Reg_7.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_7 (
    .I(\DLX_IDinst_Imm[7] ),
    .CE(DLX_IDinst__n0617),
    .CLK(clkdiv),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<7>/FFY/RST ),
    .O(\DLX_IDinst_Cause_Reg[7] )
  );
  X_BUF \DLX_IDinst_Cause_Reg<7>/FFY/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<7>/FFY/RST )
  );
  defparam DLX_IDinst_Cause_Reg_8.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_8 (
    .I(\DLX_IDinst_Imm[8] ),
    .CE(DLX_IDinst__n0617),
    .CLK(clkdiv),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<8>/FFY/RST ),
    .O(\DLX_IDinst_Cause_Reg[8] )
  );
  X_BUF \DLX_IDinst_Cause_Reg<8>/FFY/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<8>/FFY/RST )
  );
  defparam DLX_IDinst_Cause_Reg_9.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_9 (
    .I(\DLX_IDinst_Imm[9] ),
    .CE(DLX_IDinst__n0617),
    .CLK(clkdiv),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<9>/FFY/RST ),
    .O(\DLX_IDinst_Cause_Reg[9] )
  );
  X_BUF \DLX_IDinst_Cause_Reg<9>/FFY/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<9>/FFY/RST )
  );
  defparam DLX_IDinst_delay_slot_3416.INIT = 1'b0;
  X_SFF DLX_IDinst_delay_slot_3416 (
    .I(N146881),
    .CE(DLX_IDinst__n0615),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_delay_slot)
  );
  defparam DLX_IDinst_reg_dst_3417.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_dst_3417 (
    .I(N147993),
    .CE(DLX_IDinst__n0116),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_IDinst__n0115),
    .O(DLX_IDinst_reg_dst)
  );
  defparam DLX_IDinst_reg_write_3418.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_write_3418 (
    .I(N148197),
    .CE(DLX_IDinst__n0116),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_IDinst__n0115),
    .O(DLX_IDinst_reg_write)
  );
  defparam DLX_IFinst_IR_curr_0.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_0 (
    .I(IR[0]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[0])
  );
  defparam DLX_IFinst_NPC_10.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_10 (
    .I(\DLX_IFinst_NPC<10>/GROM ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC[10])
  );
  defparam DLX_IFinst_stalled_3419.INIT = 1'b0;
  X_SFF DLX_IFinst_stalled_3419 (
    .I(\DLX_IFinst_stalled/FROM ),
    .CE(\DLX_IFinst_stalled/CEMUXNOT ),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_IFinst_stalled)
  );
  defparam DLX_IDinst_RegFile_6_27_3420.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_6_27_3420 (
    .I(DLX_IDinst_WB_data_eff[27]),
    .CE(DLX_IDinst__n0562),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_6_27)
  );
  defparam DLX_IDinst_RegFile_31_18_3421.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_31_18_3421 (
    .I(DLX_IDinst_WB_data_eff[18]),
    .CE(DLX_IDinst__n0612),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_31_18)
  );
  defparam DLX_IDinst_RegFile_7_20_3422.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_7_20_3422 (
    .I(DLX_IDinst_WB_data_eff[20]),
    .CE(DLX_IDinst__n0564),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_7_20)
  );
  defparam DLX_IDinst_RegFile_31_19_3423.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_31_19_3423 (
    .I(DLX_IDinst_WB_data_eff[19]),
    .CE(DLX_IDinst__n0612),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_31_19)
  );
  defparam DLX_IDinst_RegFile_7_12_3424.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_7_12_3424 (
    .I(DLX_IDinst_WB_data_eff[12]),
    .CE(DLX_IDinst__n0564),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_7_12)
  );
  defparam DLX_IDinst_RegFile_23_27_3425.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_23_27_3425 (
    .I(DLX_IDinst_WB_data_eff[27]),
    .CE(DLX_IDinst__n0596),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_23_27)
  );
  defparam DLX_IFinst_NPC_11.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_11 (
    .I(\DLX_IFinst_NPC<11>/GROM ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC[11])
  );
  defparam DLX_IFinst_NPC_20.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_20 (
    .I(DLX_IFinst__n0001[20]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC[20])
  );
  defparam DLX_IFinst_NPC_12.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_12 (
    .I(\DLX_IFinst_NPC<12>/GROM ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC[12])
  );
  defparam DLX_IFinst_NPC_21.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_21 (
    .I(DLX_IFinst__n0001[21]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC[21])
  );
  defparam DLX_IDinst_branch_address_10.INIT = 1'b0;
  X_SFF DLX_IDinst_branch_address_10 (
    .I(N140319),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_branch_address[10])
  );
  defparam DLX_IFinst_NPC_13.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_13 (
    .I(\DLX_IFinst_NPC<13>/GROM ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC[13])
  );
  defparam DLX_IDinst_RegFile_2_12_3426.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_2_12_3426 (
    .I(DLX_IDinst_WB_data_eff[12]),
    .CE(DLX_IDinst__n0554),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_2_12)
  );
  defparam DLX_IDinst_branch_address_11.INIT = 1'b0;
  X_SFF DLX_IDinst_branch_address_11 (
    .I(N140382),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_branch_address[11])
  );
  defparam DLX_IDinst_branch_address_20.INIT = 1'b0;
  X_SFF DLX_IDinst_branch_address_20 (
    .I(N141013),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_branch_address[20])
  );
  defparam DLX_IDinst_branch_address_12.INIT = 1'b0;
  X_SFF DLX_IDinst_branch_address_12 (
    .I(N140445),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_branch_address[12])
  );
  defparam DLX_IDinst_branch_address_13.INIT = 1'b0;
  X_SFF DLX_IDinst_branch_address_13 (
    .I(N140508),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_branch_address[13])
  );
  defparam DLX_IFinst_IR_latched_0.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_latched_0 (
    .I(DLX_IFinst__n0003[0]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_latched[0])
  );
  defparam DLX_IFinst_IR_latched_1.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_latched_1 (
    .I(DLX_IFinst__n0003[1]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_latched[1])
  );
  defparam DLX_IFinst_IR_latched_3.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_latched_3 (
    .I(DLX_IFinst__n0003[3]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_latched[3])
  );
  defparam DLX_IFinst_IR_latched_2.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_latched_2 (
    .I(DLX_IFinst__n0003[2]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_latched[2])
  );
  defparam DLX_IFinst_IR_latched_4.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_latched_4 (
    .I(DLX_IFinst__n0003[4]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_latched[4])
  );
  defparam DLX_IFinst_IR_latched_5.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_latched_5 (
    .I(DLX_IFinst__n0003[5]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_latched[5])
  );
  defparam DLX_IFinst_IR_latched_6.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_latched_6 (
    .I(DLX_IFinst__n0003[6]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_latched[6])
  );
  defparam DLX_IFinst_IR_latched_7.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_latched_7 (
    .I(DLX_IFinst__n0003[7]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_latched[7])
  );
  defparam DLX_IFinst_IR_latched_8.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_latched_8 (
    .I(DLX_IFinst__n0003[8]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_latched[8])
  );
  defparam DLX_IDinst_RegFile_12_0_3427.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_12_0_3427 (
    .I(DLX_MEMinst_RF_data_in[0]),
    .CE(DLX_IDinst__n0574),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_12_0)
  );
  defparam DLX_IDinst_RegFile_20_0_3428.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_20_0_3428 (
    .I(DLX_MEMinst_RF_data_in[0]),
    .CE(DLX_IDinst__n0590),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_20_0)
  );
  defparam DLX_IDinst_RegFile_11_5_3429.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_11_5_3429 (
    .I(DLX_MEMinst_RF_data_in[5]),
    .CE(DLX_IDinst__n0572),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_11_5)
  );
  defparam DLX_IDinst_RegFile_12_1_3430.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_12_1_3430 (
    .I(DLX_MEMinst_RF_data_in[1]),
    .CE(DLX_IDinst__n0574),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_12_1)
  );
  defparam DLX_IDinst_RegFile_20_1_3431.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_20_1_3431 (
    .I(DLX_MEMinst_RF_data_in[1]),
    .CE(DLX_IDinst__n0590),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_20_1)
  );
  defparam DLX_IDinst_RegFile_12_2_3432.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_12_2_3432 (
    .I(DLX_MEMinst_RF_data_in[2]),
    .CE(DLX_IDinst__n0574),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_12_2)
  );
  defparam DLX_IDinst_RegFile_11_6_3433.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_11_6_3433 (
    .I(DLX_MEMinst_RF_data_in[6]),
    .CE(DLX_IDinst__n0572),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_11_6)
  );
  defparam DLX_IDinst_RegFile_12_6_3434.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_12_6_3434 (
    .I(DLX_MEMinst_RF_data_in[6]),
    .CE(DLX_IDinst__n0574),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_12_6)
  );
  defparam DLX_IDinst_RegFile_13_2_3435.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_13_2_3435 (
    .I(DLX_MEMinst_RF_data_in[2]),
    .CE(DLX_IDinst__n0576),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_13_2)
  );
  defparam DLX_IDinst_RegFile_20_6_3436.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_20_6_3436 (
    .I(DLX_MEMinst_RF_data_in[6]),
    .CE(DLX_IDinst__n0590),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_20_6)
  );
  defparam DLX_IDinst_RegFile_12_7_3437.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_12_7_3437 (
    .I(DLX_MEMinst_RF_data_in[7]),
    .CE(DLX_IDinst__n0574),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_12_7)
  );
  defparam DLX_IDinst_RegFile_21_2_3438.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_21_2_3438 (
    .I(DLX_MEMinst_RF_data_in[2]),
    .CE(DLX_IDinst__n0592),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_21_2)
  );
  defparam DLX_IDinst_RegFile_21_0_3439.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_21_0_3439 (
    .I(DLX_MEMinst_RF_data_in[0]),
    .CE(DLX_IDinst__n0592),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_21_0)
  );
  defparam DLX_IDinst_RegFile_11_9_3440.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_11_9_3440 (
    .I(DLX_IDinst_WB_data_eff[9]),
    .CE(DLX_IDinst__n0572),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_11_9)
  );
  defparam DLX_IDinst_RegFile_12_5_3441.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_12_5_3441 (
    .I(DLX_MEMinst_RF_data_in[5]),
    .CE(DLX_IDinst__n0574),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_12_5)
  );
  defparam DLX_IDinst_RegFile_13_1_3442.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_13_1_3442 (
    .I(DLX_MEMinst_RF_data_in[1]),
    .CE(DLX_IDinst__n0576),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_13_1)
  );
  defparam DLX_IDinst_RegFile_21_1_3443.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_21_1_3443 (
    .I(DLX_MEMinst_RF_data_in[1]),
    .CE(DLX_IDinst__n0592),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_21_1)
  );
  defparam DLX_IDinst_RegFile_20_5_3444.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_20_5_3444 (
    .I(DLX_MEMinst_RF_data_in[5]),
    .CE(DLX_IDinst__n0590),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_20_5)
  );
  defparam DLX_IDinst_RegFile_20_8_3445.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_20_8_3445 (
    .I(DLX_IDinst_WB_data_eff[8]),
    .CE(DLX_IDinst__n0590),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_20_8)
  );
  defparam DLX_IDinst_RegFile_21_4_3446.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_21_4_3446 (
    .I(DLX_MEMinst_RF_data_in[4]),
    .CE(DLX_IDinst__n0592),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_21_4)
  );
  defparam DLX_IDinst_RegFile_13_5_3447.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_13_5_3447 (
    .I(DLX_MEMinst_RF_data_in[5]),
    .CE(DLX_IDinst__n0576),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_13_5)
  );
  defparam DLX_IDinst_RegFile_22_0_3448.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_22_0_3448 (
    .I(DLX_MEMinst_RF_data_in[0]),
    .CE(DLX_IDinst__n0594),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_22_0)
  );
  defparam DLX_IDinst_RegFile_12_9_3449.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_12_9_3449 (
    .I(DLX_IDinst_WB_data_eff[9]),
    .CE(DLX_IDinst__n0574),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_12_9)
  );
  defparam DLX_IDinst_RegFile_30_0_3450.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_30_0_3450 (
    .I(DLX_MEMinst_RF_data_in[0]),
    .CE(DLX_IDinst__n0610),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_30_0)
  );
  defparam DLX_IDinst_RegFile_14_1_3451.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_14_1_3451 (
    .I(DLX_MEMinst_RF_data_in[1]),
    .CE(DLX_IDinst__n0578),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_14_1)
  );
  defparam DLX_IDinst_RegFile_21_5_3452.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_21_5_3452 (
    .I(DLX_MEMinst_RF_data_in[5]),
    .CE(DLX_IDinst__n0592),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_21_5)
  );
  defparam DLX_IDinst_RegFile_20_9_3453.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_20_9_3453 (
    .I(DLX_IDinst_WB_data_eff[9]),
    .CE(DLX_IDinst__n0590),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_20_9)
  );
  defparam DLX_IDinst_RegFile_22_1_3454.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_22_1_3454 (
    .I(DLX_MEMinst_RF_data_in[1]),
    .CE(DLX_IDinst__n0594),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_22_1)
  );
  defparam DLX_IDinst_RegFile_13_6_3455.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_13_6_3455 (
    .I(DLX_MEMinst_RF_data_in[6]),
    .CE(DLX_IDinst__n0576),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_13_6)
  );
  defparam DLX_IDinst_RegFile_14_2_3456.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_14_2_3456 (
    .I(DLX_MEMinst_RF_data_in[2]),
    .CE(DLX_IDinst__n0578),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_14_2)
  );
  defparam DLX_IDinst_RegFile_30_1_3457.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_30_1_3457 (
    .I(DLX_MEMinst_RF_data_in[1]),
    .CE(DLX_IDinst__n0610),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_30_1)
  );
  defparam DLX_IDinst_RegFile_13_3_3458.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_13_3_3458 (
    .I(DLX_MEMinst_RF_data_in[3]),
    .CE(DLX_IDinst__n0576),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_13_3)
  );
  defparam DLX_IDinst_RegFile_20_7_3459.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_20_7_3459 (
    .I(DLX_MEMinst_RF_data_in[7]),
    .CE(DLX_IDinst__n0590),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_20_7)
  );
  defparam DLX_IDinst_RegFile_21_3_3460.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_21_3_3460 (
    .I(DLX_MEMinst_RF_data_in[3]),
    .CE(DLX_IDinst__n0592),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_21_3)
  );
  defparam DLX_IDinst_RegFile_14_0_3461.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_14_0_3461 (
    .I(DLX_MEMinst_RF_data_in[0]),
    .CE(DLX_IDinst__n0578),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_14_0)
  );
  defparam DLX_IDinst_RegFile_12_8_3462.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_12_8_3462 (
    .I(DLX_IDinst_WB_data_eff[8]),
    .CE(DLX_IDinst__n0574),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_12_8)
  );
  defparam DLX_IDinst_RegFile_13_4_3463.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_13_4_3463 (
    .I(DLX_MEMinst_RF_data_in[4]),
    .CE(DLX_IDinst__n0576),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_13_4)
  );
  defparam DLX_IDinst_RegFile_22_5_3464.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_22_5_3464 (
    .I(DLX_MEMinst_RF_data_in[5]),
    .CE(DLX_IDinst__n0594),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_22_5)
  );
  defparam DLX_IDinst_RegFile_14_5_3465.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_14_5_3465 (
    .I(DLX_MEMinst_RF_data_in[5]),
    .CE(DLX_IDinst__n0578),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_14_5)
  );
  defparam DLX_IDinst_RegFile_13_9_3466.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_13_9_3466 (
    .I(DLX_IDinst_WB_data_eff[9]),
    .CE(DLX_IDinst__n0576),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_13_9)
  );
  defparam DLX_IDinst_RegFile_21_9_3467.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_21_9_3467 (
    .I(DLX_IDinst_WB_data_eff[9]),
    .CE(DLX_IDinst__n0592),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_21_9)
  );
  defparam DLX_IDinst_RegFile_15_1_3468.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_15_1_3468 (
    .I(DLX_MEMinst_RF_data_in[1]),
    .CE(DLX_IDinst__n0580),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_15_1)
  );
  defparam DLX_IDinst_RegFile_15_2_3469.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_15_2_3469 (
    .I(DLX_MEMinst_RF_data_in[2]),
    .CE(DLX_IDinst__n0580),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_15_2)
  );
  defparam DLX_IDinst_RegFile_31_1_3470.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_31_1_3470 (
    .I(DLX_MEMinst_RF_data_in[1]),
    .CE(DLX_IDinst__n0612),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_31_1)
  );
  defparam DLX_IDinst_RegFile_30_5_3471.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_30_5_3471 (
    .I(DLX_MEMinst_RF_data_in[5]),
    .CE(DLX_IDinst__n0610),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_30_5)
  );
  defparam DLX_IDinst_RegFile_13_8_3472.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_13_8_3472 (
    .I(DLX_IDinst_WB_data_eff[8]),
    .CE(DLX_IDinst__n0576),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_13_8)
  );
  defparam DLX_IDinst_RegFile_31_0_3473.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_31_0_3473 (
    .I(DLX_MEMinst_RF_data_in[0]),
    .CE(DLX_IDinst__n0612),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_31_0)
  );
  defparam DLX_IDinst_RegFile_22_4_3474.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_22_4_3474 (
    .I(DLX_MEMinst_RF_data_in[4]),
    .CE(DLX_IDinst__n0594),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_22_4)
  );
  defparam DLX_IDinst_RegFile_14_4_3475.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_14_4_3475 (
    .I(DLX_MEMinst_RF_data_in[4]),
    .CE(DLX_IDinst__n0578),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_14_4)
  );
  defparam DLX_IDinst_RegFile_21_8_3476.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_21_8_3476 (
    .I(DLX_IDinst_WB_data_eff[8]),
    .CE(DLX_IDinst__n0592),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_21_8)
  );
  defparam DLX_IDinst_RegFile_15_0_3477.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_15_0_3477 (
    .I(DLX_MEMinst_RF_data_in[0]),
    .CE(DLX_IDinst__n0580),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_15_0)
  );
  defparam DLX_IDinst_RegFile_30_4_3478.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_30_4_3478 (
    .I(DLX_MEMinst_RF_data_in[4]),
    .CE(DLX_IDinst__n0610),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_30_4)
  );
  defparam DLX_IDinst_RegFile_23_0_3479.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_23_0_3479 (
    .I(DLX_MEMinst_RF_data_in[0]),
    .CE(DLX_IDinst__n0596),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_23_0)
  );
  defparam DLX_IDinst_RegFile_30_8_3480.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_30_8_3480 (
    .I(DLX_IDinst_WB_data_eff[8]),
    .CE(DLX_IDinst__n0610),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_30_8)
  );
  defparam DLX_IDinst_RegFile_23_4_3481.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_23_4_3481 (
    .I(DLX_MEMinst_RF_data_in[4]),
    .CE(DLX_IDinst__n0596),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_23_4)
  );
  defparam DLX_IDinst_RegFile_24_0_3482.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_24_0_3482 (
    .I(DLX_MEMinst_RF_data_in[0]),
    .CE(DLX_IDinst__n0598),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_24_0)
  );
  defparam DLX_IDinst_RegFile_31_4_3483.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_31_4_3483 (
    .I(DLX_MEMinst_RF_data_in[4]),
    .CE(DLX_IDinst__n0612),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_31_4)
  );
  defparam DLX_IDinst_RegFile_16_1_3484.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_16_1_3484 (
    .I(DLX_MEMinst_RF_data_in[1]),
    .CE(DLX_IDinst__n0582),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_16_1)
  );
  defparam DLX_IDinst_RegFile_14_9_3485.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_14_9_3485 (
    .I(DLX_IDinst_WB_data_eff[9]),
    .CE(DLX_IDinst__n0578),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_14_9)
  );
  defparam DLX_IDinst_RegFile_23_5_3486.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_23_5_3486 (
    .I(DLX_MEMinst_RF_data_in[5]),
    .CE(DLX_IDinst__n0596),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_23_5)
  );
  defparam DLX_IDinst_RegFile_30_6_3487.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_30_6_3487 (
    .I(DLX_MEMinst_RF_data_in[6]),
    .CE(DLX_IDinst__n0610),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_30_6)
  );
  defparam DLX_IDinst_RegFile_31_2_3488.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_31_2_3488 (
    .I(DLX_MEMinst_RF_data_in[2]),
    .CE(DLX_IDinst__n0612),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_31_2)
  );
  defparam DLX_IDinst_RegFile_31_3_3489.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_31_3_3489 (
    .I(DLX_MEMinst_RF_data_in[3]),
    .CE(DLX_IDinst__n0612),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_31_3)
  );
  defparam DLX_IDinst_RegFile_15_3_3490.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_15_3_3490 (
    .I(DLX_MEMinst_RF_data_in[3]),
    .CE(DLX_IDinst__n0580),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_15_3)
  );
  defparam DLX_IDinst_RegFile_30_7_3491.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_30_7_3491 (
    .I(DLX_MEMinst_RF_data_in[7]),
    .CE(DLX_IDinst__n0610),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_30_7)
  );
  defparam DLX_IDinst_RegFile_22_7_3492.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_22_7_3492 (
    .I(DLX_MEMinst_RF_data_in[7]),
    .CE(DLX_IDinst__n0594),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_22_7)
  );
  defparam DLX_IDinst_RegFile_16_0_3493.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_16_0_3493 (
    .I(DLX_MEMinst_RF_data_in[0]),
    .CE(DLX_IDinst__n0582),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_16_0)
  );
  defparam DLX_IDinst_RegFile_15_4_3494.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_15_4_3494 (
    .I(DLX_MEMinst_RF_data_in[4]),
    .CE(DLX_IDinst__n0580),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_15_4)
  );
  defparam DLX_IDinst_RegFile_17_0_3495.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_17_0_3495 (
    .I(DLX_MEMinst_RF_data_in[0]),
    .CE(DLX_IDinst__n0584),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_17_0)
  );
  defparam DLX_IDinst_RegFile_24_4_3496.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_24_4_3496 (
    .I(DLX_MEMinst_RF_data_in[4]),
    .CE(DLX_IDinst__n0598),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_24_4)
  );
  defparam DLX_IDinst_RegFile_25_0_3497.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_25_0_3497 (
    .I(DLX_MEMinst_RF_data_in[0]),
    .CE(DLX_IDinst__n0600),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_25_0)
  );
  defparam DLX_IDinst_RegFile_31_8_3498.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_31_8_3498 (
    .I(DLX_IDinst_WB_data_eff[8]),
    .CE(DLX_IDinst__n0612),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_31_8)
  );
  defparam DLX_IDinst_RegFile_17_1_3499.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_17_1_3499 (
    .I(DLX_MEMinst_RF_data_in[1]),
    .CE(DLX_IDinst__n0584),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_17_1)
  );
  defparam DLX_IDinst_RegFile_16_5_3500.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_16_5_3500 (
    .I(DLX_MEMinst_RF_data_in[5]),
    .CE(DLX_IDinst__n0582),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_16_5)
  );
  defparam DLX_IDinst_RegFile_24_1_3501.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_24_1_3501 (
    .I(DLX_MEMinst_RF_data_in[1]),
    .CE(DLX_IDinst__n0598),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_24_1)
  );
  defparam DLX_IDinst_RegFile_30_9_3502.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_30_9_3502 (
    .I(DLX_IDinst_WB_data_eff[9]),
    .CE(DLX_IDinst__n0610),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_30_9)
  );
  defparam DLX_IDinst_RegFile_31_5_3503.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_31_5_3503 (
    .I(DLX_MEMinst_RF_data_in[5]),
    .CE(DLX_IDinst__n0612),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_31_5)
  );
  defparam DLX_IDinst_RegFile_24_2_3504.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_24_2_3504 (
    .I(DLX_MEMinst_RF_data_in[2]),
    .CE(DLX_IDinst__n0598),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_24_2)
  );
  defparam DLX_IDinst_RegFile_15_6_3505.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_15_6_3505 (
    .I(DLX_MEMinst_RF_data_in[6]),
    .CE(DLX_IDinst__n0580),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_15_6)
  );
  defparam DLX_IDinst_RegFile_23_6_3506.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_23_6_3506 (
    .I(DLX_MEMinst_RF_data_in[6]),
    .CE(DLX_IDinst__n0596),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_23_6)
  );
  defparam DLX_IDinst_RegFile_16_2_3507.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_16_2_3507 (
    .I(DLX_MEMinst_RF_data_in[2]),
    .CE(DLX_IDinst__n0582),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_16_2)
  );
  defparam DLX_IDinst_RegFile_31_6_3508.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_31_6_3508 (
    .I(DLX_MEMinst_RF_data_in[6]),
    .CE(DLX_IDinst__n0612),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_31_6)
  );
  defparam DLX_IDinst_RegFile_16_3_3509.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_16_3_3509 (
    .I(DLX_MEMinst_RF_data_in[3]),
    .CE(DLX_IDinst__n0582),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_16_3)
  );
  defparam DLX_IDinst_RegFile_24_3_3510.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_24_3_3510 (
    .I(DLX_MEMinst_RF_data_in[3]),
    .CE(DLX_IDinst__n0598),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_24_3)
  );
  defparam DLX_IDinst_RegFile_31_7_3511.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_31_7_3511 (
    .I(DLX_MEMinst_RF_data_in[7]),
    .CE(DLX_IDinst__n0612),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_31_7)
  );
  defparam DLX_IDinst_RegFile_16_4_3512.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_16_4_3512 (
    .I(DLX_MEMinst_RF_data_in[4]),
    .CE(DLX_IDinst__n0582),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_16_4)
  );
  defparam DLX_IDinst_RegFile_15_8_3513.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_15_8_3513 (
    .I(DLX_IDinst_WB_data_eff[8]),
    .CE(DLX_IDinst__n0580),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_15_8)
  );
  defparam DLX_IDinst_RegFile_23_9_3514.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_23_9_3514 (
    .I(DLX_IDinst_WB_data_eff[9]),
    .CE(DLX_IDinst__n0596),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_23_9)
  );
  defparam DLX_IDinst_RegFile_25_1_3515.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_25_1_3515 (
    .I(DLX_MEMinst_RF_data_in[1]),
    .CE(DLX_IDinst__n0600),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_25_1)
  );
  defparam DLX_IDinst_RegFile_24_5_3516.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_24_5_3516 (
    .I(DLX_MEMinst_RF_data_in[5]),
    .CE(DLX_IDinst__n0598),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_24_5)
  );
  defparam DLX_IDinst_RegFile_31_9_3517.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_31_9_3517 (
    .I(DLX_IDinst_WB_data_eff[9]),
    .CE(DLX_IDinst__n0612),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_31_9)
  );
  defparam DLX_IDinst_RegFile_16_6_3518.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_16_6_3518 (
    .I(DLX_MEMinst_RF_data_in[6]),
    .CE(DLX_IDinst__n0582),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_16_6)
  );
  defparam DLX_IDinst_RegFile_17_2_3519.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_17_2_3519 (
    .I(DLX_MEMinst_RF_data_in[2]),
    .CE(DLX_IDinst__n0584),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_17_2)
  );
  defparam DLX_IDinst_RegFile_25_2_3520.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_25_2_3520 (
    .I(DLX_MEMinst_RF_data_in[2]),
    .CE(DLX_IDinst__n0600),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_25_2)
  );
  defparam DLX_IDinst_RegFile_24_6_3521.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_24_6_3521 (
    .I(DLX_MEMinst_RF_data_in[6]),
    .CE(DLX_IDinst__n0598),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_24_6)
  );
  defparam DLX_IDinst_RegFile_17_3_3522.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_17_3_3522 (
    .I(DLX_MEMinst_RF_data_in[3]),
    .CE(DLX_IDinst__n0584),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_17_3)
  );
  defparam DLX_IDinst_RegFile_16_7_3523.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_16_7_3523 (
    .I(DLX_MEMinst_RF_data_in[7]),
    .CE(DLX_IDinst__n0582),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_16_7)
  );
  defparam DLX_IDinst_RegFile_24_7_3524.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_24_7_3524 (
    .I(DLX_MEMinst_RF_data_in[7]),
    .CE(DLX_IDinst__n0598),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_24_7)
  );
  defparam DLX_IDinst_RegFile_25_3_3525.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_25_3_3525 (
    .I(DLX_MEMinst_RF_data_in[3]),
    .CE(DLX_IDinst__n0600),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_25_3)
  );
  defparam DLX_IDinst_RegFile_16_8_3526.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_16_8_3526 (
    .I(DLX_IDinst_WB_data_eff[8]),
    .CE(DLX_IDinst__n0582),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_16_8)
  );
  defparam DLX_IDinst_RegFile_17_4_3527.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_17_4_3527 (
    .I(DLX_MEMinst_RF_data_in[4]),
    .CE(DLX_IDinst__n0584),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_17_4)
  );
  defparam DLX_IDinst_RegFile_18_0_3528.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_18_0_3528 (
    .I(DLX_MEMinst_RF_data_in[0]),
    .CE(DLX_IDinst__n0586),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_18_0)
  );
  defparam DLX_IDinst_RegFile_25_4_3529.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_25_4_3529 (
    .I(DLX_MEMinst_RF_data_in[4]),
    .CE(DLX_IDinst__n0600),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_25_4)
  );
  defparam DLX_IDinst_RegFile_24_8_3530.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_24_8_3530 (
    .I(DLX_IDinst_WB_data_eff[8]),
    .CE(DLX_IDinst__n0598),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_24_8)
  );
  defparam DLX_IDinst_RegFile_16_9_3531.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_16_9_3531 (
    .I(DLX_IDinst_WB_data_eff[9]),
    .CE(DLX_IDinst__n0582),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_16_9)
  );
  defparam DLX_IDinst_RegFile_25_6_3532.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_25_6_3532 (
    .I(DLX_MEMinst_RF_data_in[6]),
    .CE(DLX_IDinst__n0600),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_25_6)
  );
  defparam DLX_IDinst_RegFile_25_7_3533.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_25_7_3533 (
    .I(DLX_MEMinst_RF_data_in[7]),
    .CE(DLX_IDinst__n0600),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_25_7)
  );
  defparam vga_top_vga1_helpcounter_2.INIT = 1'b0;
  X_SFF vga_top_vga1_helpcounter_2 (
    .I(vga_top_vga1_helpcounter__n0000[2]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(vga_top_vga1__n0052),
    .SRST(reset_IBUF_1),
    .O(vga_top_vga1_helpcounter[2])
  );
  defparam DLX_IDinst_RegFile_17_8_3534.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_17_8_3534 (
    .I(DLX_IDinst_WB_data_eff[8]),
    .CE(DLX_IDinst__n0584),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_17_8)
  );
  defparam DLX_IDinst_RegFile_26_4_3535.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_26_4_3535 (
    .I(DLX_MEMinst_RF_data_in[4]),
    .CE(DLX_IDinst__n0602),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_26_4)
  );
  defparam DLX_IDinst_RegFile_27_0_3536.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_27_0_3536 (
    .I(DLX_MEMinst_RF_data_in[0]),
    .CE(DLX_IDinst__n0604),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_27_0)
  );
  defparam DLX_IDinst_RegFile_25_8_3537.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_25_8_3537 (
    .I(DLX_IDinst_WB_data_eff[8]),
    .CE(DLX_IDinst__n0600),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_25_8)
  );
  defparam DLX_IFinst_IR_previous_22.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_22 (
    .I(DLX_IFinst_IR_latched[22]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[22])
  );
  defparam DLX_IDinst_RegFile_17_5_3538.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_17_5_3538 (
    .I(DLX_MEMinst_RF_data_in[5]),
    .CE(DLX_IDinst__n0584),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_17_5)
  );
  defparam DLX_IDinst_RegFile_24_9_3539.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_24_9_3539 (
    .I(DLX_IDinst_WB_data_eff[9]),
    .CE(DLX_IDinst__n0598),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_24_9)
  );
  defparam DLX_IDinst_RegFile_25_5_3540.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_25_5_3540 (
    .I(DLX_MEMinst_RF_data_in[5]),
    .CE(DLX_IDinst__n0600),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_25_5)
  );
  defparam DLX_IDinst_RegFile_18_2_3541.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_18_2_3541 (
    .I(DLX_MEMinst_RF_data_in[2]),
    .CE(DLX_IDinst__n0586),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_18_2)
  );
  defparam DLX_IDinst_RegFile_26_1_3542.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_26_1_3542 (
    .I(DLX_MEMinst_RF_data_in[1]),
    .CE(DLX_IDinst__n0602),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_26_1)
  );
  defparam DLX_IDinst_RegFile_17_6_3543.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_17_6_3543 (
    .I(DLX_MEMinst_RF_data_in[6]),
    .CE(DLX_IDinst__n0584),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_17_6)
  );
  defparam DLX_IDinst_RegFile_19_4_3544.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_19_4_3544 (
    .I(DLX_MEMinst_RF_data_in[4]),
    .CE(DLX_IDinst__n0588),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_19_4)
  );
  defparam DLX_IDinst_RegFile_26_8_3545.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_26_8_3545 (
    .I(DLX_IDinst_WB_data_eff[8]),
    .CE(DLX_IDinst__n0602),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_26_8)
  );
  defparam DLX_IDinst_RegFile_27_4_3546.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_27_4_3546 (
    .I(DLX_MEMinst_RF_data_in[4]),
    .CE(DLX_IDinst__n0604),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_27_4)
  );
  defparam DLX_IDinst_RegFile_28_0_3547.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_28_0_3547 (
    .I(DLX_MEMinst_RF_data_in[0]),
    .CE(DLX_IDinst__n0606),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_28_0)
  );
  defparam DLX_IDinst_RegFile_18_9_3548.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_18_9_3548 (
    .I(DLX_IDinst_WB_data_eff[9]),
    .CE(DLX_IDinst__n0586),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_18_9)
  );
  defparam DLX_IDinst_RegFile_19_5_3549.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_19_5_3549 (
    .I(DLX_MEMinst_RF_data_in[5]),
    .CE(DLX_IDinst__n0588),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_19_5)
  );
  defparam DLX_IDinst_RegFile_26_9_3550.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_26_9_3550 (
    .I(DLX_IDinst_WB_data_eff[9]),
    .CE(DLX_IDinst__n0602),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_26_9)
  );
  defparam DLX_IDinst_RegFile_27_5_3551.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_27_5_3551 (
    .I(DLX_MEMinst_RF_data_in[5]),
    .CE(DLX_IDinst__n0604),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_27_5)
  );
  defparam DLX_IDinst_RegFile_28_1_3552.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_28_1_3552 (
    .I(DLX_MEMinst_RF_data_in[1]),
    .CE(DLX_IDinst__n0606),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_28_1)
  );
  defparam DLX_IDinst_RegFile_19_6_3553.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_19_6_3553 (
    .I(DLX_MEMinst_RF_data_in[6]),
    .CE(DLX_IDinst__n0588),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_19_6)
  );
  defparam DLX_IDinst_RegFile_27_6_3554.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_27_6_3554 (
    .I(DLX_MEMinst_RF_data_in[6]),
    .CE(DLX_IDinst__n0604),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_27_6)
  );
  defparam DLX_IDinst_RegFile_28_2_3555.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_28_2_3555 (
    .I(DLX_MEMinst_RF_data_in[2]),
    .CE(DLX_IDinst__n0606),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_28_2)
  );
  defparam DLX_IDinst_RegFile_19_7_3556.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_19_7_3556 (
    .I(DLX_MEMinst_RF_data_in[7]),
    .CE(DLX_IDinst__n0588),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_19_7)
  );
  defparam DLX_IDinst_RegFile_27_7_3557.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_27_7_3557 (
    .I(DLX_MEMinst_RF_data_in[7]),
    .CE(DLX_IDinst__n0604),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_27_7)
  );
  defparam DLX_IDinst_RegFile_28_3_3558.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_28_3_3558 (
    .I(DLX_MEMinst_RF_data_in[3]),
    .CE(DLX_IDinst__n0606),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_28_3)
  );
  defparam DLX_IDinst_RegFile_19_8_3559.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_19_8_3559 (
    .I(DLX_IDinst_WB_data_eff[8]),
    .CE(DLX_IDinst__n0588),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_19_8)
  );
  defparam DLX_IDinst_RegFile_27_8_3560.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_27_8_3560 (
    .I(DLX_IDinst_WB_data_eff[8]),
    .CE(DLX_IDinst__n0604),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_27_8)
  );
  defparam DLX_IDinst_RegFile_28_4_3561.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_28_4_3561 (
    .I(DLX_MEMinst_RF_data_in[4]),
    .CE(DLX_IDinst__n0606),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_28_4)
  );
  defparam DLX_IDinst_RegFile_29_0_3562.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_29_0_3562 (
    .I(DLX_MEMinst_RF_data_in[0]),
    .CE(DLX_IDinst__n0608),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_29_0)
  );
  defparam DLX_IDinst_RegFile_19_9_3563.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_19_9_3563 (
    .I(DLX_IDinst_WB_data_eff[9]),
    .CE(DLX_IDinst__n0588),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_19_9)
  );
  defparam DLX_IDinst_RegFile_27_9_3564.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_27_9_3564 (
    .I(DLX_IDinst_WB_data_eff[9]),
    .CE(DLX_IDinst__n0604),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_27_9)
  );
  defparam DLX_IDinst_RegFile_28_5_3565.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_28_5_3565 (
    .I(DLX_MEMinst_RF_data_in[5]),
    .CE(DLX_IDinst__n0606),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_28_5)
  );
  defparam DLX_IDinst_RegFile_19_1_3566.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_19_1_3566 (
    .I(DLX_MEMinst_RF_data_in[1]),
    .CE(DLX_IDinst__n0588),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_19_1)
  );
  defparam DLX_IDinst_RegFile_27_1_3567.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_27_1_3567 (
    .I(DLX_MEMinst_RF_data_in[1]),
    .CE(DLX_IDinst__n0604),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_27_1)
  );
  defparam DLX_IDinst_RegFile_26_6_3568.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_26_6_3568 (
    .I(DLX_MEMinst_RF_data_in[6]),
    .CE(DLX_IDinst__n0602),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_26_6)
  );
  defparam DLX_IDinst_RegFile_25_9_3569.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_25_9_3569 (
    .I(DLX_IDinst_WB_data_eff[9]),
    .CE(DLX_IDinst__n0600),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_25_9)
  );
  defparam DLX_IDinst_RegFile_19_2_3570.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_19_2_3570 (
    .I(DLX_MEMinst_RF_data_in[2]),
    .CE(DLX_IDinst__n0588),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_19_2)
  );
  defparam DLX_IDinst_RegFile_18_6_3571.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_18_6_3571 (
    .I(DLX_MEMinst_RF_data_in[6]),
    .CE(DLX_IDinst__n0586),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_18_6)
  );
  defparam DLX_IDinst_RegFile_27_2_3572.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_27_2_3572 (
    .I(DLX_MEMinst_RF_data_in[2]),
    .CE(DLX_IDinst__n0604),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_27_2)
  );
  defparam DLX_IDinst_RegFile_18_7_3573.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_18_7_3573 (
    .I(DLX_MEMinst_RF_data_in[7]),
    .CE(DLX_IDinst__n0586),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_18_7)
  );
  defparam DLX_IDinst_RegFile_19_3_3574.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_19_3_3574 (
    .I(DLX_MEMinst_RF_data_in[3]),
    .CE(DLX_IDinst__n0588),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_19_3)
  );
  defparam DLX_IDinst_RegFile_26_7_3575.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_26_7_3575 (
    .I(DLX_MEMinst_RF_data_in[7]),
    .CE(DLX_IDinst__n0602),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_26_7)
  );
  defparam DLX_IDinst_RegFile_18_8_3576.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_18_8_3576 (
    .I(DLX_IDinst_WB_data_eff[8]),
    .CE(DLX_IDinst__n0586),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_18_8)
  );
  defparam DLX_IDinst_RegFile_27_3_3577.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_27_3_3577 (
    .I(DLX_MEMinst_RF_data_in[3]),
    .CE(DLX_IDinst__n0604),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_27_3)
  );
  defparam DLX_IDinst_RegFile_29_1_3578.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_29_1_3578 (
    .I(DLX_MEMinst_RF_data_in[1]),
    .CE(DLX_IDinst__n0608),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_29_1)
  );
  defparam DLX_IDinst_RegFile_28_6_3579.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_28_6_3579 (
    .I(DLX_MEMinst_RF_data_in[6]),
    .CE(DLX_IDinst__n0606),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_28_6)
  );
  defparam DLX_IDinst_RegFile_29_2_3580.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_29_2_3580 (
    .I(DLX_MEMinst_RF_data_in[2]),
    .CE(DLX_IDinst__n0608),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_29_2)
  );
  defparam DLX_IDinst_RegFile_28_7_3581.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_28_7_3581 (
    .I(DLX_MEMinst_RF_data_in[7]),
    .CE(DLX_IDinst__n0606),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_28_7)
  );
  defparam DLX_IDinst_RegFile_29_3_3582.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_29_3_3582 (
    .I(DLX_MEMinst_RF_data_in[3]),
    .CE(DLX_IDinst__n0608),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_29_3)
  );
  defparam DLX_IDinst_RegFile_28_8_3583.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_28_8_3583 (
    .I(DLX_IDinst_WB_data_eff[8]),
    .CE(DLX_IDinst__n0606),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_28_8)
  );
  defparam DLX_IDinst_RegFile_29_4_3584.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_29_4_3584 (
    .I(DLX_MEMinst_RF_data_in[4]),
    .CE(DLX_IDinst__n0608),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_29_4)
  );
  defparam DLX_IDinst_RegFile_28_9_3585.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_28_9_3585 (
    .I(DLX_IDinst_WB_data_eff[9]),
    .CE(DLX_IDinst__n0606),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_28_9)
  );
  defparam DLX_IDinst_RegFile_29_5_3586.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_29_5_3586 (
    .I(DLX_MEMinst_RF_data_in[5]),
    .CE(DLX_IDinst__n0608),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_29_5)
  );
  defparam DLX_IDinst_RegFile_29_6_3587.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_29_6_3587 (
    .I(DLX_MEMinst_RF_data_in[6]),
    .CE(DLX_IDinst__n0608),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_29_6)
  );
  defparam DLX_IDinst_RegFile_29_8_3588.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_29_8_3588 (
    .I(DLX_IDinst_WB_data_eff[8]),
    .CE(DLX_IDinst__n0608),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_29_8)
  );
  defparam DLX_IDinst_RegFile_29_9_3589.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_29_9_3589 (
    .I(DLX_IDinst_WB_data_eff[9]),
    .CE(DLX_IDinst__n0608),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_29_9)
  );
  defparam DLX_IDinst_RegFile_6_9_3590.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_6_9_3590 (
    .I(DLX_IDinst_WB_data_eff[9]),
    .CE(DLX_IDinst__n0562),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_6_9)
  );
  defparam DLX_IDinst_RegFile_2_14_3591.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_2_14_3591 (
    .I(DLX_IDinst_WB_data_eff[14]),
    .CE(DLX_IDinst__n0554),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_2_14)
  );
  defparam DLX_IDinst_RegFile_0_21_3592.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_0_21_3592 (
    .I(DLX_IDinst_WB_data_eff[21]),
    .CE(DLX_IDinst__n0550),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_0_21)
  );
  defparam DLX_IDinst_RegFile_0_11_3593.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_0_11_3593 (
    .I(DLX_IDinst_WB_data_eff[11]),
    .CE(DLX_IDinst__n0550),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_0_11)
  );
  defparam DLX_IDinst_RegFile_0_13_3594.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_0_13_3594 (
    .I(DLX_IDinst_WB_data_eff[13]),
    .CE(DLX_IDinst__n0550),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_0_13)
  );
  defparam DLX_IDinst_RegFile_0_30_3595.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_0_30_3595 (
    .I(DLX_IDinst_WB_data_eff[30]),
    .CE(DLX_IDinst__n0550),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_0_30)
  );
  defparam DLX_IDinst_RegFile_0_22_3596.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_0_22_3596 (
    .I(DLX_IDinst_WB_data_eff[22]),
    .CE(DLX_IDinst__n0550),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_0_22)
  );
  defparam DLX_IDinst_RegFile_0_14_3597.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_0_14_3597 (
    .I(DLX_IDinst_WB_data_eff[14]),
    .CE(DLX_IDinst__n0550),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_0_14)
  );
  defparam DLX_IDinst_RegFile_0_31_3598.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_0_31_3598 (
    .I(DLX_IDinst_WB_data_eff[31]),
    .CE(DLX_IDinst__n0550),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_0_31)
  );
  defparam DLX_IDinst_RegFile_0_23_3599.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_0_23_3599 (
    .I(DLX_IDinst_WB_data_eff[23]),
    .CE(DLX_IDinst__n0550),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_0_23)
  );
  defparam DLX_IDinst_RegFile_0_15_3600.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_0_15_3600 (
    .I(DLX_IDinst_WB_data_eff[15]),
    .CE(DLX_IDinst__n0550),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_0_15)
  );
  defparam DLX_IDinst_RegFile_0_24_3601.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_0_24_3601 (
    .I(DLX_IDinst_WB_data_eff[24]),
    .CE(DLX_IDinst__n0550),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_0_24)
  );
  defparam DLX_IDinst_RegFile_0_16_3602.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_0_16_3602 (
    .I(DLX_IDinst_WB_data_eff[16]),
    .CE(DLX_IDinst__n0550),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_0_16)
  );
  defparam DLX_IDinst_RegFile_0_17_3603.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_0_17_3603 (
    .I(DLX_IDinst_WB_data_eff[17]),
    .CE(DLX_IDinst__n0550),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_0_17)
  );
  defparam DLX_IDinst_RegFile_0_25_3604.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_0_25_3604 (
    .I(DLX_IDinst_WB_data_eff[25]),
    .CE(DLX_IDinst__n0550),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_0_25)
  );
  defparam DLX_IDinst_RegFile_1_10_3605.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_1_10_3605 (
    .I(DLX_IDinst_WB_data_eff[10]),
    .CE(DLX_IDinst__n0552),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_1_10)
  );
  defparam DLX_IDinst_RegFile_0_26_3606.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_0_26_3606 (
    .I(DLX_IDinst_WB_data_eff[26]),
    .CE(DLX_IDinst__n0550),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_0_26)
  );
  defparam DLX_IDinst_RegFile_0_18_3607.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_0_18_3607 (
    .I(DLX_IDinst_WB_data_eff[18]),
    .CE(DLX_IDinst__n0550),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_0_18)
  );
  defparam DLX_IDinst_RegFile_1_11_3608.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_1_11_3608 (
    .I(DLX_IDinst_WB_data_eff[11]),
    .CE(DLX_IDinst__n0552),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_1_11)
  );
  defparam DLX_IDinst_RegFile_0_27_3609.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_0_27_3609 (
    .I(DLX_IDinst_WB_data_eff[27]),
    .CE(DLX_IDinst__n0550),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_0_27)
  );
  defparam DLX_IDinst_RegFile_0_19_3610.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_0_19_3610 (
    .I(DLX_IDinst_WB_data_eff[19]),
    .CE(DLX_IDinst__n0550),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_0_19)
  );
  defparam DLX_IDinst_RegFile_1_12_3611.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_1_12_3611 (
    .I(DLX_IDinst_WB_data_eff[12]),
    .CE(DLX_IDinst__n0552),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_1_12)
  );
  defparam DLX_IDinst_RegFile_0_28_3612.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_0_28_3612 (
    .I(DLX_IDinst_WB_data_eff[28]),
    .CE(DLX_IDinst__n0550),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_0_28)
  );
  defparam DLX_IDinst_RegFile_1_20_3613.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_1_20_3613 (
    .I(DLX_IDinst_WB_data_eff[20]),
    .CE(DLX_IDinst__n0552),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_1_20)
  );
  defparam DLX_IDinst_RegFile_1_13_3614.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_1_13_3614 (
    .I(DLX_IDinst_WB_data_eff[13]),
    .CE(DLX_IDinst__n0552),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_1_13)
  );
  defparam DLX_IDinst_RegFile_0_29_3615.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_0_29_3615 (
    .I(DLX_IDinst_WB_data_eff[29]),
    .CE(DLX_IDinst__n0550),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_0_29)
  );
  defparam DLX_IDinst_RegFile_1_21_3616.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_1_21_3616 (
    .I(DLX_IDinst_WB_data_eff[21]),
    .CE(DLX_IDinst__n0552),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_1_21)
  );
  defparam DLX_IDinst_RegFile_1_14_3617.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_1_14_3617 (
    .I(DLX_IDinst_WB_data_eff[14]),
    .CE(DLX_IDinst__n0552),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_1_14)
  );
  defparam DLX_IDinst_RegFile_1_30_3618.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_1_30_3618 (
    .I(DLX_IDinst_WB_data_eff[30]),
    .CE(DLX_IDinst__n0552),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_1_30)
  );
  defparam DLX_IDinst_RegFile_1_22_3619.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_1_22_3619 (
    .I(DLX_IDinst_WB_data_eff[22]),
    .CE(DLX_IDinst__n0552),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_1_22)
  );
  defparam DLX_IDinst_RegFile_1_31_3620.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_1_31_3620 (
    .I(DLX_IDinst_WB_data_eff[31]),
    .CE(DLX_IDinst__n0552),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_1_31)
  );
  defparam DLX_IDinst_RegFile_1_15_3621.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_1_15_3621 (
    .I(DLX_IDinst_WB_data_eff[15]),
    .CE(DLX_IDinst__n0552),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_1_15)
  );
  defparam DLX_IDinst_RegFile_1_16_3622.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_1_16_3622 (
    .I(DLX_IDinst_WB_data_eff[16]),
    .CE(DLX_IDinst__n0552),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_1_16)
  );
  defparam DLX_IDinst_RegFile_1_25_3623.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_1_25_3623 (
    .I(DLX_IDinst_WB_data_eff[25]),
    .CE(DLX_IDinst__n0552),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_1_25)
  );
  defparam DLX_IDinst_RegFile_2_10_3624.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_2_10_3624 (
    .I(DLX_IDinst_WB_data_eff[10]),
    .CE(DLX_IDinst__n0554),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_2_10)
  );
  defparam DLX_IDinst_RegFile_1_18_3625.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_1_18_3625 (
    .I(DLX_IDinst_WB_data_eff[18]),
    .CE(DLX_IDinst__n0552),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_1_18)
  );
  defparam DLX_IDinst_RegFile_2_11_3626.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_2_11_3626 (
    .I(DLX_IDinst_WB_data_eff[11]),
    .CE(DLX_IDinst__n0554),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_2_11)
  );
  defparam DLX_IDinst_RegFile_1_27_3627.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_1_27_3627 (
    .I(DLX_IDinst_WB_data_eff[27]),
    .CE(DLX_IDinst__n0552),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_1_27)
  );
  defparam DLX_IDinst_RegFile_4_10_3628.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_4_10_3628 (
    .I(DLX_IDinst_WB_data_eff[10]),
    .CE(DLX_IDinst__n0558),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_4_10)
  );
  defparam DLX_IDinst_RegFile_4_11_3629.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_4_11_3629 (
    .I(DLX_IDinst_WB_data_eff[11]),
    .CE(DLX_IDinst__n0558),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_4_11)
  );
  defparam DLX_IDinst_RegFile_4_12_3630.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_4_12_3630 (
    .I(DLX_IDinst_WB_data_eff[12]),
    .CE(DLX_IDinst__n0558),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_4_12)
  );
  defparam DLX_IDinst_RegFile_4_20_3631.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_4_20_3631 (
    .I(DLX_IDinst_WB_data_eff[20]),
    .CE(DLX_IDinst__n0558),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_4_20)
  );
  defparam DLX_IDinst_RegFile_4_13_3632.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_4_13_3632 (
    .I(DLX_IDinst_WB_data_eff[13]),
    .CE(DLX_IDinst__n0558),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_4_13)
  );
  defparam DLX_IDinst_RegFile_4_14_3633.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_4_14_3633 (
    .I(DLX_IDinst_WB_data_eff[14]),
    .CE(DLX_IDinst__n0558),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_4_14)
  );
  defparam DLX_IDinst_RegFile_4_21_3634.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_4_21_3634 (
    .I(DLX_IDinst_WB_data_eff[21]),
    .CE(DLX_IDinst__n0558),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_4_21)
  );
  defparam DLX_IDinst_RegFile_4_22_3635.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_4_22_3635 (
    .I(DLX_IDinst_WB_data_eff[22]),
    .CE(DLX_IDinst__n0558),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_4_22)
  );
  defparam DLX_IDinst_RegFile_4_30_3636.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_4_30_3636 (
    .I(DLX_IDinst_WB_data_eff[30]),
    .CE(DLX_IDinst__n0558),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_4_30)
  );
  defparam DLX_IDinst_RegFile_4_31_3637.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_4_31_3637 (
    .I(DLX_IDinst_WB_data_eff[31]),
    .CE(DLX_IDinst__n0558),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_4_31)
  );
  defparam DLX_IDinst_RegFile_4_23_3638.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_4_23_3638 (
    .I(DLX_IDinst_WB_data_eff[23]),
    .CE(DLX_IDinst__n0558),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_4_23)
  );
  defparam DLX_IDinst_RegFile_4_15_3639.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_4_15_3639 (
    .I(DLX_IDinst_WB_data_eff[15]),
    .CE(DLX_IDinst__n0558),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_4_15)
  );
  defparam DLX_IDinst_RegFile_4_16_3640.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_4_16_3640 (
    .I(DLX_IDinst_WB_data_eff[16]),
    .CE(DLX_IDinst__n0558),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_4_16)
  );
  defparam DLX_IDinst_RegFile_4_24_3641.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_4_24_3641 (
    .I(DLX_IDinst_WB_data_eff[24]),
    .CE(DLX_IDinst__n0558),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_4_24)
  );
  defparam DLX_IDinst_RegFile_4_17_3642.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_4_17_3642 (
    .I(DLX_IDinst_WB_data_eff[17]),
    .CE(DLX_IDinst__n0558),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_4_17)
  );
  defparam DLX_IDinst_RegFile_4_26_3643.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_4_26_3643 (
    .I(DLX_IDinst_WB_data_eff[26]),
    .CE(DLX_IDinst__n0558),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_4_26)
  );
  defparam DLX_IDinst_RegFile_4_25_3644.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_4_25_3644 (
    .I(DLX_IDinst_WB_data_eff[25]),
    .CE(DLX_IDinst__n0558),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_4_25)
  );
  defparam DLX_IDinst_RegFile_4_18_3645.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_4_18_3645 (
    .I(DLX_IDinst_WB_data_eff[18]),
    .CE(DLX_IDinst__n0558),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_4_18)
  );
  defparam DLX_IDinst_RegFile_5_10_3646.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_5_10_3646 (
    .I(DLX_IDinst_WB_data_eff[10]),
    .CE(DLX_IDinst__n0560),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_5_10)
  );
  defparam DLX_IDinst_RegFile_4_19_3647.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_4_19_3647 (
    .I(DLX_IDinst_WB_data_eff[19]),
    .CE(DLX_IDinst__n0558),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_4_19)
  );
  defparam DLX_IDinst_RegFile_4_27_3648.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_4_27_3648 (
    .I(DLX_IDinst_WB_data_eff[27]),
    .CE(DLX_IDinst__n0558),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_4_27)
  );
  defparam DLX_IDinst_RegFile_4_28_3649.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_4_28_3649 (
    .I(DLX_IDinst_WB_data_eff[28]),
    .CE(DLX_IDinst__n0558),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_4_28)
  );
  defparam DLX_IDinst_RegFile_5_11_3650.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_5_11_3650 (
    .I(DLX_IDinst_WB_data_eff[11]),
    .CE(DLX_IDinst__n0560),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_5_11)
  );
  defparam DLX_IDinst_RegFile_5_20_3651.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_5_20_3651 (
    .I(DLX_IDinst_WB_data_eff[20]),
    .CE(DLX_IDinst__n0560),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_5_20)
  );
  defparam DLX_IDinst_RegFile_5_12_3652.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_5_12_3652 (
    .I(DLX_IDinst_WB_data_eff[12]),
    .CE(DLX_IDinst__n0560),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_5_12)
  );
  defparam DLX_IDinst_RegFile_4_29_3653.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_4_29_3653 (
    .I(DLX_IDinst_WB_data_eff[29]),
    .CE(DLX_IDinst__n0558),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_4_29)
  );
  defparam DLX_IDinst_RegFile_5_13_3654.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_5_13_3654 (
    .I(DLX_IDinst_WB_data_eff[13]),
    .CE(DLX_IDinst__n0560),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_5_13)
  );
  defparam DLX_IDinst_RegFile_5_21_3655.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_5_21_3655 (
    .I(DLX_IDinst_WB_data_eff[21]),
    .CE(DLX_IDinst__n0560),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_5_21)
  );
  defparam DLX_IDinst_RegFile_6_29_3656.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_6_29_3656 (
    .I(DLX_IDinst_WB_data_eff[29]),
    .CE(DLX_IDinst__n0562),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_6_29)
  );
  defparam DLX_IDinst_RegFile_7_21_3657.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_7_21_3657 (
    .I(DLX_IDinst_WB_data_eff[21]),
    .CE(DLX_IDinst__n0564),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_7_21)
  );
  defparam DLX_IDinst_RegFile_7_13_3658.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_7_13_3658 (
    .I(DLX_IDinst_WB_data_eff[13]),
    .CE(DLX_IDinst__n0564),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_7_13)
  );
  defparam DLX_IDinst_RegFile_7_30_3659.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_7_30_3659 (
    .I(DLX_IDinst_WB_data_eff[30]),
    .CE(DLX_IDinst__n0564),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_7_30)
  );
  defparam DLX_IDinst_RegFile_7_22_3660.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_7_22_3660 (
    .I(DLX_IDinst_WB_data_eff[22]),
    .CE(DLX_IDinst__n0564),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_7_22)
  );
  defparam DLX_IDinst_RegFile_7_14_3661.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_7_14_3661 (
    .I(DLX_IDinst_WB_data_eff[14]),
    .CE(DLX_IDinst__n0564),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_7_14)
  );
  defparam DLX_IDinst_RegFile_7_23_3662.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_7_23_3662 (
    .I(DLX_IDinst_WB_data_eff[23]),
    .CE(DLX_IDinst__n0564),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_7_23)
  );
  defparam DLX_IDinst_RegFile_7_15_3663.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_7_15_3663 (
    .I(DLX_IDinst_WB_data_eff[15]),
    .CE(DLX_IDinst__n0564),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_7_15)
  );
  defparam DLX_IDinst_RegFile_7_31_3664.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_7_31_3664 (
    .I(DLX_IDinst_WB_data_eff[31]),
    .CE(DLX_IDinst__n0564),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_7_31)
  );
  defparam DLX_IDinst_RegFile_7_24_3665.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_7_24_3665 (
    .I(DLX_IDinst_WB_data_eff[24]),
    .CE(DLX_IDinst__n0564),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_7_24)
  );
  defparam DLX_IDinst_RegFile_7_16_3666.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_7_16_3666 (
    .I(DLX_IDinst_WB_data_eff[16]),
    .CE(DLX_IDinst__n0564),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_7_16)
  );
  defparam DLX_IDinst_RegFile_7_25_3667.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_7_25_3667 (
    .I(DLX_IDinst_WB_data_eff[25]),
    .CE(DLX_IDinst__n0564),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_7_25)
  );
  defparam DLX_IDinst_RegFile_7_17_3668.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_7_17_3668 (
    .I(DLX_IDinst_WB_data_eff[17]),
    .CE(DLX_IDinst__n0564),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_7_17)
  );
  defparam DLX_IDinst_RegFile_7_26_3669.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_7_26_3669 (
    .I(DLX_IDinst_WB_data_eff[26]),
    .CE(DLX_IDinst__n0564),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_7_26)
  );
  defparam DLX_IDinst_RegFile_7_18_3670.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_7_18_3670 (
    .I(DLX_IDinst_WB_data_eff[18]),
    .CE(DLX_IDinst__n0564),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_7_18)
  );
  defparam DLX_IDinst_RegFile_8_10_3671.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_8_10_3671 (
    .I(DLX_IDinst_WB_data_eff[10]),
    .CE(DLX_IDinst__n0566),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_8_10)
  );
  defparam DLX_IDinst_RegFile_7_19_3672.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_7_19_3672 (
    .I(DLX_IDinst_WB_data_eff[19]),
    .CE(DLX_IDinst__n0564),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_7_19)
  );
  defparam DLX_IDinst_RegFile_7_27_3673.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_7_27_3673 (
    .I(DLX_IDinst_WB_data_eff[27]),
    .CE(DLX_IDinst__n0564),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_7_27)
  );
  defparam DLX_IDinst_RegFile_5_18_3674.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_5_18_3674 (
    .I(DLX_IDinst_WB_data_eff[18]),
    .CE(DLX_IDinst__n0560),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_5_18)
  );
  defparam DLX_IDinst_RegFile_5_27_3675.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_5_27_3675 (
    .I(DLX_IDinst_WB_data_eff[27]),
    .CE(DLX_IDinst__n0560),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_5_27)
  );
  defparam DLX_IDinst_RegFile_5_19_3676.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_5_19_3676 (
    .I(DLX_IDinst_WB_data_eff[19]),
    .CE(DLX_IDinst__n0560),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_5_19)
  );
  defparam DLX_IDinst_RegFile_6_28_3677.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_6_28_3677 (
    .I(DLX_IDinst_WB_data_eff[28]),
    .CE(DLX_IDinst__n0562),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_6_28)
  );
  defparam DLX_IDinst_RegFile_5_28_3678.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_5_28_3678 (
    .I(DLX_IDinst_WB_data_eff[28]),
    .CE(DLX_IDinst__n0560),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_5_28)
  );
  defparam DLX_IDinst_RegFile_5_24_3679.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_5_24_3679 (
    .I(DLX_IDinst_WB_data_eff[24]),
    .CE(DLX_IDinst__n0560),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_5_24)
  );
  defparam DLX_IDinst_RegFile_5_16_3680.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_5_16_3680 (
    .I(DLX_IDinst_WB_data_eff[16]),
    .CE(DLX_IDinst__n0560),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_5_16)
  );
  defparam DLX_IDinst_RegFile_5_25_3681.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_5_25_3681 (
    .I(DLX_IDinst_WB_data_eff[25]),
    .CE(DLX_IDinst__n0560),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_5_25)
  );
  defparam DLX_IDinst_RegFile_5_26_3682.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_5_26_3682 (
    .I(DLX_IDinst_WB_data_eff[26]),
    .CE(DLX_IDinst__n0560),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_5_26)
  );
  defparam DLX_IDinst_RegFile_5_17_3683.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_5_17_3683 (
    .I(DLX_IDinst_WB_data_eff[17]),
    .CE(DLX_IDinst__n0560),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_5_17)
  );
  defparam DLX_IDinst_RegFile_5_30_3684.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_5_30_3684 (
    .I(DLX_IDinst_WB_data_eff[30]),
    .CE(DLX_IDinst__n0560),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_5_30)
  );
  defparam DLX_IDinst_RegFile_5_22_3685.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_5_22_3685 (
    .I(DLX_IDinst_WB_data_eff[22]),
    .CE(DLX_IDinst__n0560),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_5_22)
  );
  defparam DLX_IDinst_RegFile_5_14_3686.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_5_14_3686 (
    .I(DLX_IDinst_WB_data_eff[14]),
    .CE(DLX_IDinst__n0560),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_5_14)
  );
  defparam DLX_IDinst_RegFile_5_15_3687.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_5_15_3687 (
    .I(DLX_IDinst_WB_data_eff[15]),
    .CE(DLX_IDinst__n0560),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_5_15)
  );
  defparam DLX_IDinst_RegFile_5_31_3688.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_5_31_3688 (
    .I(DLX_IDinst_WB_data_eff[31]),
    .CE(DLX_IDinst__n0560),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_5_31)
  );
  defparam DLX_IDinst_RegFile_5_23_3689.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_5_23_3689 (
    .I(DLX_IDinst_WB_data_eff[23]),
    .CE(DLX_IDinst__n0560),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_5_23)
  );
  defparam DLX_IDinst_RegFile_7_28_3690.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_7_28_3690 (
    .I(DLX_IDinst_WB_data_eff[28]),
    .CE(DLX_IDinst__n0564),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_7_28)
  );
  defparam DLX_IDinst_RegFile_8_11_3691.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_8_11_3691 (
    .I(DLX_IDinst_WB_data_eff[11]),
    .CE(DLX_IDinst__n0566),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_8_11)
  );
  defparam DLX_IDinst_RegFile_8_12_3692.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_8_12_3692 (
    .I(DLX_IDinst_WB_data_eff[12]),
    .CE(DLX_IDinst__n0566),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_8_12)
  );
  defparam DLX_IDinst_RegFile_8_20_3693.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_8_20_3693 (
    .I(DLX_IDinst_WB_data_eff[20]),
    .CE(DLX_IDinst__n0566),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_8_20)
  );
  defparam DLX_IDinst_RegFile_8_30_3694.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_8_30_3694 (
    .I(DLX_IDinst_WB_data_eff[30]),
    .CE(DLX_IDinst__n0566),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_8_30)
  );
  defparam DLX_IDinst_RegFile_7_29_3695.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_7_29_3695 (
    .I(DLX_IDinst_WB_data_eff[29]),
    .CE(DLX_IDinst__n0564),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_7_29)
  );
  defparam DLX_IDinst_RegFile_8_13_3696.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_8_13_3696 (
    .I(DLX_IDinst_WB_data_eff[13]),
    .CE(DLX_IDinst__n0566),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_8_13)
  );
  defparam DLX_IDinst_RegFile_8_21_3697.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_8_21_3697 (
    .I(DLX_IDinst_WB_data_eff[21]),
    .CE(DLX_IDinst__n0566),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_8_21)
  );
  defparam DLX_IDinst_RegFile_8_22_3698.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_8_22_3698 (
    .I(DLX_IDinst_WB_data_eff[22]),
    .CE(DLX_IDinst__n0566),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_8_22)
  );
  defparam DLX_IDinst_RegFile_8_14_3699.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_8_14_3699 (
    .I(DLX_IDinst_WB_data_eff[14]),
    .CE(DLX_IDinst__n0566),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_8_14)
  );
  defparam DLX_IDinst_RegFile_8_23_3700.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_8_23_3700 (
    .I(DLX_IDinst_WB_data_eff[23]),
    .CE(DLX_IDinst__n0566),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_8_23)
  );
  defparam DLX_IDinst_RegFile_8_31_3701.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_8_31_3701 (
    .I(DLX_IDinst_WB_data_eff[31]),
    .CE(DLX_IDinst__n0566),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_8_31)
  );
  defparam DLX_IDinst_RegFile_8_15_3702.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_8_15_3702 (
    .I(DLX_IDinst_WB_data_eff[15]),
    .CE(DLX_IDinst__n0566),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_8_15)
  );
  defparam DLX_IDinst_RegFile_9_10_3703.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_9_10_3703 (
    .I(DLX_IDinst_WB_data_eff[10]),
    .CE(DLX_IDinst__n0568),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_9_10)
  );
  defparam DLX_IDinst_RegFile_8_19_3704.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_8_19_3704 (
    .I(DLX_IDinst_WB_data_eff[19]),
    .CE(DLX_IDinst__n0566),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_8_19)
  );
  defparam DLX_IDinst_RegFile_8_27_3705.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_8_27_3705 (
    .I(DLX_IDinst_WB_data_eff[27]),
    .CE(DLX_IDinst__n0566),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_8_27)
  );
  defparam DLX_IDinst_RegFile_8_28_3706.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_8_28_3706 (
    .I(DLX_IDinst_WB_data_eff[28]),
    .CE(DLX_IDinst__n0566),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_8_28)
  );
  defparam DLX_IDinst_RegFile_9_11_3707.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_9_11_3707 (
    .I(DLX_IDinst_WB_data_eff[11]),
    .CE(DLX_IDinst__n0568),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_9_11)
  );
  defparam DLX_IDinst_RegFile_9_30_3708.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_9_30_3708 (
    .I(DLX_IDinst_WB_data_eff[30]),
    .CE(DLX_IDinst__n0568),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_9_30)
  );
  defparam DLX_IDinst_RegFile_9_22_3709.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_9_22_3709 (
    .I(DLX_IDinst_WB_data_eff[22]),
    .CE(DLX_IDinst__n0568),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_9_22)
  );
  defparam DLX_IDinst_RegFile_9_31_3710.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_9_31_3710 (
    .I(DLX_IDinst_WB_data_eff[31]),
    .CE(DLX_IDinst__n0568),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_9_31)
  );
  defparam DLX_IDinst_RegFile_9_14_3711.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_9_14_3711 (
    .I(DLX_IDinst_WB_data_eff[14]),
    .CE(DLX_IDinst__n0568),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_9_14)
  );
  defparam DLX_IDinst_RegFile_9_15_3712.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_9_15_3712 (
    .I(DLX_IDinst_WB_data_eff[15]),
    .CE(DLX_IDinst__n0568),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_9_15)
  );
  defparam DLX_IDinst_RegFile_9_23_3713.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_9_23_3713 (
    .I(DLX_IDinst_WB_data_eff[23]),
    .CE(DLX_IDinst__n0568),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_9_23)
  );
  defparam DLX_IDinst_RegFile_9_18_3714.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_9_18_3714 (
    .I(DLX_IDinst_WB_data_eff[18]),
    .CE(DLX_IDinst__n0568),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_9_18)
  );
  defparam DLX_IDinst_RegFile_9_27_3715.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_9_27_3715 (
    .I(DLX_IDinst_WB_data_eff[27]),
    .CE(DLX_IDinst__n0568),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_9_27)
  );
  defparam DLX_IDinst_RegFile_9_19_3716.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_9_19_3716 (
    .I(DLX_IDinst_WB_data_eff[19]),
    .CE(DLX_IDinst__n0568),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_9_19)
  );
  defparam DLX_IDinst_RegFile_9_29_3717.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_9_29_3717 (
    .I(DLX_IDinst_WB_data_eff[29]),
    .CE(DLX_IDinst__n0568),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_9_29)
  );
  defparam DLX_IDinst_RegFile_9_28_3718.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_9_28_3718 (
    .I(DLX_IDinst_WB_data_eff[28]),
    .CE(DLX_IDinst__n0568),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_9_28)
  );
  defparam DLX_IFinst_PC_0.INIT = 1'b0;
  X_SFF DLX_IFinst_PC_0 (
    .I(DLX_IFinst_NPC[0]),
    .CE(DLX_IFinst_PC_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_PC[0])
  );
  defparam DLX_IDinst_RegFile_8_24_3719.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_8_24_3719 (
    .I(DLX_IDinst_WB_data_eff[24]),
    .CE(DLX_IDinst__n0566),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_8_24)
  );
  defparam DLX_IDinst_RegFile_8_16_3720.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_8_16_3720 (
    .I(DLX_IDinst_WB_data_eff[16]),
    .CE(DLX_IDinst__n0566),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_8_16)
  );
  defparam DLX_IDinst_RegFile_8_25_3721.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_8_25_3721 (
    .I(DLX_IDinst_WB_data_eff[25]),
    .CE(DLX_IDinst__n0566),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_8_25)
  );
  defparam DLX_IDinst_RegFile_8_18_3722.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_8_18_3722 (
    .I(DLX_IDinst_WB_data_eff[18]),
    .CE(DLX_IDinst__n0566),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_8_18)
  );
  defparam DLX_IDinst_RegFile_8_17_3723.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_8_17_3723 (
    .I(DLX_IDinst_WB_data_eff[17]),
    .CE(DLX_IDinst__n0566),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_8_17)
  );
  defparam DLX_IDinst_RegFile_8_26_3724.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_8_26_3724 (
    .I(DLX_IDinst_WB_data_eff[26]),
    .CE(DLX_IDinst__n0566),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_8_26)
  );
  defparam DLX_IDinst_RegFile_9_20_3725.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_9_20_3725 (
    .I(DLX_IDinst_WB_data_eff[20]),
    .CE(DLX_IDinst__n0568),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_9_20)
  );
  defparam DLX_IDinst_RegFile_9_12_3726.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_9_12_3726 (
    .I(DLX_IDinst_WB_data_eff[12]),
    .CE(DLX_IDinst__n0568),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_9_12)
  );
  defparam DLX_IDinst_RegFile_8_29_3727.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_8_29_3727 (
    .I(DLX_IDinst_WB_data_eff[29]),
    .CE(DLX_IDinst__n0566),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_8_29)
  );
  defparam DLX_IDinst_RegFile_9_13_3728.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_9_13_3728 (
    .I(DLX_IDinst_WB_data_eff[13]),
    .CE(DLX_IDinst__n0568),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_9_13)
  );
  defparam DLX_IDinst_RegFile_9_21_3729.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_9_21_3729 (
    .I(DLX_IDinst_WB_data_eff[21]),
    .CE(DLX_IDinst__n0568),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_9_21)
  );
  defparam DLX_IFinst_PC_3.INIT = 1'b0;
  X_SFF DLX_IFinst_PC_3 (
    .I(DLX_IFinst_NPC[3]),
    .CE(DLX_IFinst_PC_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_IFinst_PC[3])
  );
  defparam DLX_IFinst_PC_1.INIT = 1'b0;
  X_SFF DLX_IFinst_PC_1 (
    .I(DLX_IFinst_NPC[1]),
    .CE(DLX_IFinst_PC_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_PC[1])
  );
  defparam DLX_IFinst_PC_2.INIT = 1'b0;
  X_SFF DLX_IFinst_PC_2 (
    .I(DLX_IFinst_NPC[2]),
    .CE(DLX_IFinst_PC_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_IFinst_PC[2])
  );
  defparam DLX_IFinst_PC_4.INIT = 1'b0;
  X_SFF DLX_IFinst_PC_4 (
    .I(DLX_IFinst_NPC[4]),
    .CE(DLX_IFinst_PC_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_IFinst_PC[4])
  );
  defparam DLX_IFinst_PC_5.INIT = 1'b0;
  X_SFF DLX_IFinst_PC_5 (
    .I(DLX_IFinst_NPC[5]),
    .CE(DLX_IFinst_PC_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_IFinst_PC[5])
  );
  defparam DLX_IFinst_PC_6.INIT = 1'b0;
  X_SFF DLX_IFinst_PC_6 (
    .I(DLX_IFinst_NPC[6]),
    .CE(DLX_IFinst_PC_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_IFinst_PC[6])
  );
  defparam DLX_IFinst_PC_7.INIT = 1'b0;
  X_SFF DLX_IFinst_PC_7 (
    .I(DLX_IFinst_NPC[7]),
    .CE(DLX_IFinst_PC_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_IFinst_PC[7])
  );
  defparam DLX_IFinst_PC_8.INIT = 1'b0;
  X_SFF DLX_IFinst_PC_8 (
    .I(DLX_IFinst_NPC[8]),
    .CE(DLX_IFinst_PC_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_IFinst_PC[8])
  );
  defparam DLX_IFinst_PC_9.INIT = 1'b0;
  X_SFF DLX_IFinst_PC_9 (
    .I(DLX_IFinst_NPC[9]),
    .CE(DLX_IFinst_PC_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_IFinst_PC[9])
  );
  defparam DLX_MEMinst_opcode_of_WB_1.INIT = 1'b0;
  X_SFF DLX_MEMinst_opcode_of_WB_1 (
    .I(DLX_EXinst_opcode_of_EX_reg[1]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_MEMinst_opcode_of_WB[1])
  );
  defparam DLX_IFinst_IR_previous_3.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_3 (
    .I(DLX_IFinst_IR_latched[3]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[3])
  );
  defparam DLX_IDinst_RegFile_3_28_3730.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_3_28_3730 (
    .I(DLX_IDinst_WB_data_eff[28]),
    .CE(DLX_IDinst__n0556),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_3_28)
  );
  defparam DLX_IDinst_RegFile_9_24_3731.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_9_24_3731 (
    .I(DLX_IDinst_WB_data_eff[24]),
    .CE(DLX_IDinst__n0568),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_9_24)
  );
  defparam DLX_IDinst_RegFile_9_16_3732.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_9_16_3732 (
    .I(DLX_IDinst_WB_data_eff[16]),
    .CE(DLX_IDinst__n0568),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_9_16)
  );
  defparam DLX_IDinst_RegFile_9_25_3733.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_9_25_3733 (
    .I(DLX_IDinst_WB_data_eff[25]),
    .CE(DLX_IDinst__n0568),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_9_25)
  );
  defparam DLX_IDinst_RegFile_9_26_3734.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_9_26_3734 (
    .I(DLX_IDinst_WB_data_eff[26]),
    .CE(DLX_IDinst__n0568),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_9_26)
  );
  defparam DLX_IDinst_RegFile_9_17_3735.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_9_17_3735 (
    .I(DLX_IDinst_WB_data_eff[17]),
    .CE(DLX_IDinst__n0568),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_RegFile_9_17)
  );
  defparam DLX_IDinst_RegFile_2_1_3736.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_2_1_3736 (
    .I(DLX_MEMinst_RF_data_in[1]),
    .CE(DLX_IDinst__n0554),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_2_1)
  );
  defparam DLX_IDinst_EPC_9.INIT = 1'b0;
  X_SFF DLX_IDinst_EPC_9 (
    .I(DLX_IFinst_NPC[9]),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_EPC[9])
  );
  defparam DLX_IDinst_RegFile_0_10_3737.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_0_10_3737 (
    .I(DLX_IDinst_WB_data_eff[10]),
    .CE(DLX_IDinst__n0550),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_0_10)
  );
  defparam DLX_IDinst_RegFile_0_20_3738.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_0_20_3738 (
    .I(DLX_IDinst_WB_data_eff[20]),
    .CE(DLX_IDinst__n0550),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_0_20)
  );
  defparam DLX_IDinst_RegFile_30_31_3739.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_30_31_3739 (
    .I(DLX_IDinst_WB_data_eff[31]),
    .CE(DLX_IDinst__n0610),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_30_31)
  );
  defparam DLX_IDinst_RegFile_2_2_3740.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_2_2_3740 (
    .I(DLX_MEMinst_RF_data_in[2]),
    .CE(DLX_IDinst__n0554),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_2_2)
  );
  defparam DLX_IDinst_RegFile_2_3_3741.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_2_3_3741 (
    .I(DLX_MEMinst_RF_data_in[3]),
    .CE(DLX_IDinst__n0554),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_2_3)
  );
  defparam DLX_IDinst_RegFile_2_4_3742.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_2_4_3742 (
    .I(DLX_MEMinst_RF_data_in[4]),
    .CE(DLX_IDinst__n0554),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_2_4)
  );
  defparam DLX_EXinst_ALU_result_6.INIT = 1'b0;
  X_SFF DLX_EXinst_ALU_result_6 (
    .I(N162801),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(N136886),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_ALU_result[6])
  );
  defparam DLX_IDinst_RegFile_31_13_3743.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_31_13_3743 (
    .I(DLX_IDinst_WB_data_eff[13]),
    .CE(DLX_IDinst__n0612),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_31_13)
  );
  defparam DLX_IDinst_RegFile_31_22_3744.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_31_22_3744 (
    .I(DLX_IDinst_WB_data_eff[22]),
    .CE(DLX_IDinst__n0612),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_31_22)
  );
  defparam DLX_IDinst_RegFile_31_16_3745.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_31_16_3745 (
    .I(DLX_IDinst_WB_data_eff[16]),
    .CE(DLX_IDinst__n0612),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_31_16)
  );
  defparam DLX_IDinst_RegFile_15_31_3746.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_15_31_3746 (
    .I(DLX_IDinst_WB_data_eff[31]),
    .CE(DLX_IDinst__n0580),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_15_31)
  );
  defparam DLX_IDinst_RegFile_15_18_3747.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_15_18_3747 (
    .I(DLX_IDinst_WB_data_eff[18]),
    .CE(DLX_IDinst__n0580),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_15_18)
  );
  defparam DLX_IDinst_RegFile_15_19_3748.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_15_19_3748 (
    .I(DLX_IDinst_WB_data_eff[19]),
    .CE(DLX_IDinst__n0580),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_15_19)
  );
  defparam DLX_IDinst_RegFile_19_0_3749.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_19_0_3749 (
    .I(DLX_MEMinst_RF_data_in[0]),
    .CE(DLX_IDinst__n0588),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_19_0)
  );
  defparam DLX_IDinst_RegFile_0_3_3750.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_0_3_3750 (
    .I(DLX_MEMinst_RF_data_in[3]),
    .CE(DLX_IDinst__n0550),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_0_3)
  );
  defparam DLX_IDinst_RegFile_23_1_3751.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_23_1_3751 (
    .I(DLX_MEMinst_RF_data_in[1]),
    .CE(DLX_IDinst__n0596),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_23_1)
  );
  defparam DLX_EXinst_ALU_result_5.INIT = 1'b0;
  X_SFF DLX_EXinst_ALU_result_5 (
    .I(N162863),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(N136886),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_ALU_result[5])
  );
  defparam DLX_IDinst_RegFile_14_6_3752.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_14_6_3752 (
    .I(DLX_MEMinst_RF_data_in[6]),
    .CE(DLX_IDinst__n0578),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_14_6)
  );
  defparam DLX_IDinst_RegFile_0_5_3753.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_0_5_3753 (
    .I(DLX_MEMinst_RF_data_in[5]),
    .CE(DLX_IDinst__n0550),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_0_5)
  );
  defparam DLX_IFinst_IR_curr_17.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_17 (
    .I(IR[17]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[17])
  );
  defparam DLX_IFinst_IR_curr_26.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_26 (
    .I(IR_MSB_2_OBUF),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[26])
  );
  defparam DLX_IDinst_RegFile_11_20_3754.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_11_20_3754 (
    .I(DLX_IDinst_WB_data_eff[20]),
    .CE(DLX_IDinst__n0572),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_11_20)
  );
  defparam DLX_IDinst_RegFile_11_30_3755.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_11_30_3755 (
    .I(DLX_IDinst_WB_data_eff[30]),
    .CE(DLX_IDinst__n0572),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_11_30)
  );
  defparam DLX_IDinst_RegFile_11_15_3756.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_11_15_3756 (
    .I(DLX_IDinst_WB_data_eff[15]),
    .CE(DLX_IDinst__n0572),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_11_15)
  );
  defparam DLX_IDinst_RegFile_11_25_3757.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_11_25_3757 (
    .I(DLX_IDinst_WB_data_eff[25]),
    .CE(DLX_IDinst__n0572),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_11_25)
  );
  defparam DLX_IDinst_RegFile_1_24_3758.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_1_24_3758 (
    .I(DLX_IDinst_WB_data_eff[24]),
    .CE(DLX_IDinst__n0552),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_1_24)
  );
  defparam DLX_IDinst_RegFile_3_2_3759.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_3_2_3759 (
    .I(DLX_MEMinst_RF_data_in[2]),
    .CE(DLX_IDinst__n0556),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_3_2)
  );
  defparam DLX_IDinst_RegFile_23_3_3760.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_23_3_3760 (
    .I(DLX_MEMinst_RF_data_in[3]),
    .CE(DLX_IDinst__n0596),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_23_3)
  );
  defparam DLX_IDinst_RegFile_14_8_3761.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_14_8_3761 (
    .I(DLX_IDinst_WB_data_eff[8]),
    .CE(DLX_IDinst__n0578),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_14_8)
  );
  defparam DLX_IDinst_RegFile_3_3_3762.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_3_3_3762 (
    .I(DLX_MEMinst_RF_data_in[3]),
    .CE(DLX_IDinst__n0556),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_3_3)
  );
  defparam DLX_IDinst_RegFile_22_9_3763.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_22_9_3763 (
    .I(DLX_IDinst_WB_data_eff[9]),
    .CE(DLX_IDinst__n0594),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_22_9)
  );
  defparam DLX_IDinst_RegFile_2_8_3764.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_2_8_3764 (
    .I(DLX_IDinst_WB_data_eff[8]),
    .CE(DLX_IDinst__n0554),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_2_8)
  );
  defparam DLX_IDinst_RegFile_7_5_3765.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_7_5_3765 (
    .I(DLX_MEMinst_RF_data_in[5]),
    .CE(DLX_IDinst__n0564),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_7_5)
  );
  defparam DLX_MEMinst_RF_data_in_24.INIT = 1'b0;
  X_SFF DLX_MEMinst_RF_data_in_24 (
    .I(DLX_MEMinst__n0000[24]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_MEMinst_RF_data_in[24])
  );
  defparam DLX_IDinst_RegFile_2_9_3766.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_2_9_3766 (
    .I(DLX_IDinst_WB_data_eff[9]),
    .CE(DLX_IDinst__n0554),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_2_9)
  );
  defparam DLX_IFinst_IR_previous_23.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_23 (
    .I(DLX_IFinst_IR_latched[23]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[23])
  );
  defparam DLX_IDinst_RegFile_10_2_3767.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_10_2_3767 (
    .I(DLX_MEMinst_RF_data_in[2]),
    .CE(DLX_IDinst__n0570),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_10_2)
  );
  defparam DLX_IDinst_RegFile_10_4_3768.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_10_4_3768 (
    .I(DLX_MEMinst_RF_data_in[4]),
    .CE(DLX_IDinst__n0570),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_10_4)
  );
  defparam DLX_IDinst_RegFile_10_5_3769.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_10_5_3769 (
    .I(DLX_MEMinst_RF_data_in[5]),
    .CE(DLX_IDinst__n0570),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_10_5)
  );
  defparam DLX_IDinst_RegFile_23_7_3770.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_23_7_3770 (
    .I(DLX_MEMinst_RF_data_in[7]),
    .CE(DLX_IDinst__n0596),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_23_7)
  );
  defparam DLX_IDinst_RegFile_27_23_3771.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_27_23_3771 (
    .I(DLX_IDinst_WB_data_eff[23]),
    .CE(DLX_IDinst__n0604),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_27_23)
  );
  defparam DLX_IDinst_RegFile_3_5_3772.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_3_5_3772 (
    .I(DLX_MEMinst_RF_data_in[5]),
    .CE(DLX_IDinst__n0556),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_3_5)
  );
  defparam DLX_IFinst_IR_previous_11.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_11 (
    .I(DLX_IFinst_IR_latched[11]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[11])
  );
  defparam DLX_MEMinst_noop_3773.INIT = 1'b1;
  X_SFF DLX_MEMinst_noop_3773 (
    .I(DLX_EXinst_noop),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GSR),
    .RST(GND),
    .SSET(reset_IBUF_1),
    .SRST(GND),
    .O(DLX_MEMinst_noop)
  );
  defparam DLX_IDinst_RegFile_11_1_3774.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_11_1_3774 (
    .I(DLX_MEMinst_RF_data_in[1]),
    .CE(DLX_IDinst__n0572),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_11_1)
  );
  defparam DLX_IFinst_IR_previous_28.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_28 (
    .I(DLX_IFinst_IR_latched[28]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[28])
  );
  defparam DLX_IFinst_IR_previous_29.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_29 (
    .I(DLX_IFinst_IR_latched[29]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[29])
  );
  defparam DLX_IDinst_RegFile_10_7_3775.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_10_7_3775 (
    .I(DLX_MEMinst_RF_data_in[7]),
    .CE(DLX_IDinst__n0570),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_10_7)
  );
  defparam DLX_IDinst_RegFile_6_10_3776.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_6_10_3776 (
    .I(DLX_IDinst_WB_data_eff[10]),
    .CE(DLX_IDinst__n0562),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_6_10)
  );
  defparam DLX_IFinst_IR_previous_0.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_0 (
    .I(DLX_IFinst_IR_latched[0]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[0])
  );
  defparam DLX_IFinst_IR_previous_5.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_5 (
    .I(DLX_IFinst_IR_latched[5]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[5])
  );
  defparam DLX_EXinst_ALU_result_4.INIT = 1'b0;
  X_SFF DLX_EXinst_ALU_result_4 (
    .I(N162850),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(N136886),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_ALU_result[4])
  );
  defparam DLX_IFinst_PC_11.INIT = 1'b0;
  X_SFF DLX_IFinst_PC_11 (
    .I(DLX_IFinst_NPC[11]),
    .CE(DLX_IFinst_PC_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_PC[11])
  );
  defparam DLX_IDinst_RegFile_14_31_3777.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_14_31_3777 (
    .I(DLX_IDinst_WB_data_eff[31]),
    .CE(DLX_IDinst__n0578),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_14_31)
  );
  defparam DLX_IDinst_RegFile_6_22_3778.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_6_22_3778 (
    .I(DLX_IDinst_WB_data_eff[22]),
    .CE(DLX_IDinst__n0562),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_6_22)
  );
  defparam DLX_IDinst_RegFile_14_27_3779.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_14_27_3779 (
    .I(DLX_IDinst_WB_data_eff[27]),
    .CE(DLX_IDinst__n0578),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_14_27)
  );
  defparam DLX_IDinst_RegFile_22_19_3780.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_22_19_3780 (
    .I(DLX_IDinst_WB_data_eff[19]),
    .CE(DLX_IDinst__n0594),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_22_19)
  );
  defparam DLX_IDinst_RegFile_6_14_3781.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_6_14_3781 (
    .I(DLX_IDinst_WB_data_eff[14]),
    .CE(DLX_IDinst__n0562),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_6_14)
  );
  defparam DLX_IDinst_RegFile_6_30_3782.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_6_30_3782 (
    .I(DLX_IDinst_WB_data_eff[30]),
    .CE(DLX_IDinst__n0562),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_6_30)
  );
  defparam DLX_IDinst_RegFile_6_31_3783.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_6_31_3783 (
    .I(DLX_IDinst_WB_data_eff[31]),
    .CE(DLX_IDinst__n0562),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_6_31)
  );
  defparam DLX_IDinst_RegFile_6_15_3784.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_6_15_3784 (
    .I(DLX_IDinst_WB_data_eff[15]),
    .CE(DLX_IDinst__n0562),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_6_15)
  );
  defparam DLX_IDinst_RegFile_30_16_3785.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_30_16_3785 (
    .I(DLX_IDinst_WB_data_eff[16]),
    .CE(DLX_IDinst__n0610),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_30_16)
  );
  defparam DLX_IDinst_RegFile_22_17_3786.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_22_17_3786 (
    .I(DLX_IDinst_WB_data_eff[17]),
    .CE(DLX_IDinst__n0594),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_22_17)
  );
  defparam DLX_IDinst_RegFile_14_18_3787.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_14_18_3787 (
    .I(DLX_IDinst_WB_data_eff[18]),
    .CE(DLX_IDinst__n0578),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_14_18)
  );
  defparam DLX_IDinst_RegFile_6_21_3788.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_6_21_3788 (
    .I(DLX_IDinst_WB_data_eff[21]),
    .CE(DLX_IDinst__n0562),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_6_21)
  );
  defparam DLX_IDinst_RegFile_5_29_3789.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_5_29_3789 (
    .I(DLX_IDinst_WB_data_eff[29]),
    .CE(DLX_IDinst__n0560),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_5_29)
  );
  defparam DLX_IDinst_RegFile_23_10_3790.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_23_10_3790 (
    .I(DLX_IDinst_WB_data_eff[10]),
    .CE(DLX_IDinst__n0596),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_23_10)
  );
  defparam DLX_IDinst_RegFile_6_24_3791.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_6_24_3791 (
    .I(DLX_IDinst_WB_data_eff[24]),
    .CE(DLX_IDinst__n0562),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_6_24)
  );
  defparam DLX_IDinst_RegFile_6_17_3792.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_6_17_3792 (
    .I(DLX_IDinst_WB_data_eff[17]),
    .CE(DLX_IDinst__n0562),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_6_17)
  );
  defparam DLX_IDinst_RegFile_6_25_3793.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_6_25_3793 (
    .I(DLX_IDinst_WB_data_eff[25]),
    .CE(DLX_IDinst__n0562),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_6_25)
  );
  defparam DLX_IDinst_RegFile_7_10_3794.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_7_10_3794 (
    .I(DLX_IDinst_WB_data_eff[10]),
    .CE(DLX_IDinst__n0564),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_7_10)
  );
  defparam DLX_IDinst_RegFile_6_18_3795.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_6_18_3795 (
    .I(DLX_IDinst_WB_data_eff[18]),
    .CE(DLX_IDinst__n0562),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_6_18)
  );
  defparam DLX_IDinst_RegFile_15_17_3796.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_15_17_3796 (
    .I(DLX_IDinst_WB_data_eff[17]),
    .CE(DLX_IDinst__n0580),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_15_17)
  );
  defparam DLX_IDinst_EPC_11.INIT = 1'b0;
  X_SFF DLX_IDinst_EPC_11 (
    .I(DLX_IFinst_NPC[11]),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_EPC[11])
  );
  defparam DLX_IDinst_EPC_10.INIT = 1'b0;
  X_SFF DLX_IDinst_EPC_10 (
    .I(DLX_IFinst_NPC[10]),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_EPC[10])
  );
  defparam DLX_IDinst_EPC_20.INIT = 1'b0;
  X_SFF DLX_IDinst_EPC_20 (
    .I(DLX_IFinst_NPC[20]),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_EPC[20])
  );
  defparam DLX_IDinst_EPC_12.INIT = 1'b0;
  X_SFF DLX_IDinst_EPC_12 (
    .I(DLX_IFinst_NPC[12]),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_EPC[12])
  );
  defparam DLX_IDinst_EPC_21.INIT = 1'b0;
  X_SFF DLX_IDinst_EPC_21 (
    .I(DLX_IFinst_NPC[21]),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_EPC[21])
  );
  defparam DLX_IDinst_EPC_13.INIT = 1'b0;
  X_SFF DLX_IDinst_EPC_13 (
    .I(DLX_IFinst_NPC[13]),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_EPC[13])
  );
  defparam DLX_IDinst_EPC_30.INIT = 1'b0;
  X_SFF DLX_IDinst_EPC_30 (
    .I(DLX_IFinst_NPC[30]),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_EPC[30])
  );
  defparam DLX_IDinst_EPC_23.INIT = 1'b0;
  X_SFF DLX_IDinst_EPC_23 (
    .I(DLX_IFinst_NPC[23]),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_EPC[23])
  );
  defparam DLX_IDinst_EPC_22.INIT = 1'b0;
  X_SFF DLX_IDinst_EPC_22 (
    .I(DLX_IFinst_NPC[22]),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_EPC[22])
  );
  defparam DLX_IDinst_EPC_14.INIT = 1'b0;
  X_SFF DLX_IDinst_EPC_14 (
    .I(DLX_IFinst_NPC[14]),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_EPC[14])
  );
  defparam DLX_IDinst_RegFile_10_30_3797.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_10_30_3797 (
    .I(\DLX_IDinst_RegFile_10_30/GROM ),
    .CE(DLX_IDinst__n0570),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_10_30)
  );
  defparam DLX_IDinst_EPC_15.INIT = 1'b0;
  X_SFF DLX_IDinst_EPC_15 (
    .I(DLX_IFinst_NPC[15]),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_EPC[15])
  );
  defparam DLX_IDinst_EPC_31.INIT = 1'b0;
  X_SFF DLX_IDinst_EPC_31 (
    .I(DLX_IFinst_NPC[31]),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_EPC[31])
  );
  defparam DLX_IDinst_EPC_24.INIT = 1'b0;
  X_SFF DLX_IDinst_EPC_24 (
    .I(DLX_IFinst_NPC[24]),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_EPC[24])
  );
  defparam DLX_IDinst_EPC_16.INIT = 1'b0;
  X_SFF DLX_IDinst_EPC_16 (
    .I(DLX_IFinst_NPC[16]),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_EPC[16])
  );
  defparam DLX_IDinst_EPC_25.INIT = 1'b0;
  X_SFF DLX_IDinst_EPC_25 (
    .I(DLX_IFinst_NPC[25]),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_EPC[25])
  );
  defparam DLX_IDinst_EPC_17.INIT = 1'b0;
  X_SFF DLX_IDinst_EPC_17 (
    .I(DLX_IFinst_NPC[17]),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_EPC[17])
  );
  defparam DLX_IDinst_EPC_26.INIT = 1'b0;
  X_SFF DLX_IDinst_EPC_26 (
    .I(DLX_IFinst_NPC[26]),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_EPC[26])
  );
  defparam DLX_IDinst_EPC_18.INIT = 1'b0;
  X_SFF DLX_IDinst_EPC_18 (
    .I(DLX_IFinst_NPC[18]),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_EPC[18])
  );
  defparam DLX_IDinst_EPC_27.INIT = 1'b0;
  X_SFF DLX_IDinst_EPC_27 (
    .I(DLX_IFinst_NPC[27]),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_EPC[27])
  );
  defparam DLX_IDinst_EPC_19.INIT = 1'b0;
  X_SFF DLX_IDinst_EPC_19 (
    .I(DLX_IFinst_NPC[19]),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_EPC[19])
  );
  defparam DLX_IDinst_EPC_28.INIT = 1'b0;
  X_SFF DLX_IDinst_EPC_28 (
    .I(DLX_IFinst_NPC[28]),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_EPC[28])
  );
  defparam DLX_IDinst_branch_address_7.INIT = 1'b0;
  X_SFF DLX_IDinst_branch_address_7 (
    .I(N140126),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_branch_address[7])
  );
  defparam DLX_IDinst_branch_address_5.INIT = 1'b0;
  X_SFF DLX_IDinst_branch_address_5 (
    .I(N140078),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_branch_address[5])
  );
  defparam DLX_IDinst_EPC_0.INIT = 1'b0;
  X_SFF DLX_IDinst_EPC_0 (
    .I(DLX_IFinst_NPC[0]),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_EPC[0])
  );
  defparam DLX_IDinst_branch_address_6.INIT = 1'b0;
  X_SFF DLX_IDinst_branch_address_6 (
    .I(N145997),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_branch_address[6])
  );
  defparam DLX_IDinst_branch_address_8.INIT = 1'b0;
  X_SFF DLX_IDinst_branch_address_8 (
    .I(N140193),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_branch_address[8])
  );
  defparam DLX_IDinst_branch_address_9.INIT = 1'b0;
  X_SFF DLX_IDinst_branch_address_9 (
    .I(N140256),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_branch_address[9])
  );
  defparam DLX_IDinst_branch_address_0.INIT = 1'b0;
  X_SFF DLX_IDinst_branch_address_0 (
    .I(N145826),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_branch_address[0])
  );
  defparam DLX_IDinst_branch_address_2.INIT = 1'b0;
  X_SFF DLX_IDinst_branch_address_2 (
    .I(N139889),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_branch_address[2])
  );
  defparam DLX_IDinst_branch_address_1.INIT = 1'b0;
  X_SFF DLX_IDinst_branch_address_1 (
    .I(N139826),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_branch_address[1])
  );
  defparam DLX_IDinst_branch_address_3.INIT = 1'b0;
  X_SFF DLX_IDinst_branch_address_3 (
    .I(N139952),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_branch_address[3])
  );
  defparam DLX_IDinst_branch_address_4.INIT = 1'b0;
  X_SFF DLX_IDinst_branch_address_4 (
    .I(N140015),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_branch_address[4])
  );
  defparam DLX_IDinst_counter_0.INIT = 1'b0;
  X_SFF DLX_IDinst_counter_0 (
    .I(N144314),
    .CE(DLX_IDinst__n0549),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_counter[0])
  );
  defparam DLX_IDinst_Cause_Reg_10.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_10 (
    .I(\DLX_IDinst_Imm[10] ),
    .CE(DLX_IDinst__n0617),
    .CLK(clkdiv),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<10>/FFY/RST ),
    .O(\DLX_IDinst_Cause_Reg[10] )
  );
  X_BUF \DLX_IDinst_Cause_Reg<10>/FFY/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<10>/FFY/RST )
  );
  defparam DLX_IDinst_Cause_Reg_12.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_12 (
    .I(\DLX_IDinst_Imm[12] ),
    .CE(DLX_IDinst__n0617),
    .CLK(clkdiv),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<12>/FFY/RST ),
    .O(\DLX_IDinst_Cause_Reg[12] )
  );
  X_BUF \DLX_IDinst_Cause_Reg<12>/FFY/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<12>/FFY/RST )
  );
  defparam DLX_IDinst_Cause_Reg_11.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_11 (
    .I(\DLX_IDinst_Imm[11] ),
    .CE(DLX_IDinst__n0617),
    .CLK(clkdiv),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<11>/FFY/RST ),
    .O(\DLX_IDinst_Cause_Reg[11] )
  );
  X_BUF \DLX_IDinst_Cause_Reg<11>/FFY/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<11>/FFY/RST )
  );
  defparam DLX_IDinst_Cause_Reg_13.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_13 (
    .I(\DLX_IDinst_Imm[13] ),
    .CE(DLX_IDinst__n0617),
    .CLK(clkdiv),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<13>/FFY/RST ),
    .O(\DLX_IDinst_Cause_Reg[13] )
  );
  X_BUF \DLX_IDinst_Cause_Reg<13>/FFY/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<13>/FFY/RST )
  );
  defparam DLX_IDinst_Cause_Reg_14.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_14 (
    .I(\DLX_IDinst_Imm[14] ),
    .CE(DLX_IDinst__n0617),
    .CLK(clkdiv),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<14>/FFY/RST ),
    .O(\DLX_IDinst_Cause_Reg[14] )
  );
  X_BUF \DLX_IDinst_Cause_Reg<14>/FFY/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<14>/FFY/RST )
  );
  defparam DLX_IDinst_Cause_Reg_15.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_15 (
    .I(\DLX_IDinst_Imm[15] ),
    .CE(DLX_IDinst__n0617),
    .CLK(clkdiv),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<15>/FFY/RST ),
    .O(\DLX_IDinst_Cause_Reg[15] )
  );
  X_BUF \DLX_IDinst_Cause_Reg<15>/FFY/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<15>/FFY/RST )
  );
  defparam DLX_IDinst_Cause_Reg_31.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_31 (
    .I(DLX_IDinst_Imm_31_1),
    .CE(DLX_IDinst__n0617),
    .CLK(clkdiv),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<31>/FFY/RST ),
    .O(\DLX_IDinst_Cause_Reg[31] )
  );
  X_BUF \DLX_IDinst_Cause_Reg<31>/FFY/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<31>/FFY/RST )
  );
  defparam vga_top_vga1_helpcounter_0.INIT = 1'b0;
  X_SFF vga_top_vga1_helpcounter_0 (
    .I(\vga_top_vga1_helpcounter<0>/BXMUXNOT ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(vga_top_vga1__n0052),
    .SRST(reset_IBUF_1),
    .O(vga_top_vga1_helpcounter[0])
  );
  defparam vga_top_vga1_helpcounter_1.INIT = 1'b0;
  X_SFF vga_top_vga1_helpcounter_1 (
    .I(vga_top_vga1_helpcounter__n0000[1]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(vga_top_vga1__n0052),
    .SRST(reset_IBUF_1),
    .O(vga_top_vga1_helpcounter[1])
  );
  defparam DLX_MEMinst_reg_dst_out_3.INIT = 1'b0;
  X_SFF DLX_MEMinst_reg_dst_out_3 (
    .I(DLX_EXinst_reg_dst_out[3]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_MEMinst_reg_dst_out[3])
  );
  defparam DLX_MEMinst_reg_dst_out_4.INIT = 1'b0;
  X_SFF DLX_MEMinst_reg_dst_out_4 (
    .I(DLX_EXinst_reg_dst_out[4]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_MEMinst_reg_dst_out[4])
  );
  defparam DLX_EXinst_reg_out_B_EX_1.INIT = 1'b0;
  X_SFF DLX_EXinst_reg_out_B_EX_1 (
    .I(DLX_IDinst_reg_out_B[1]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_reg_out_B_EX[1])
  );
  defparam vga_top_vga1_videoon_3798.INIT = 1'b0;
  X_SFF vga_top_vga1_videoon_3798 (
    .I(\vga_top_vga1_videoon/LOGIC_ONE ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(N147636),
    .O(vga_top_vga1_videoon)
  );
  defparam DLX_MEMinst_reg_dst_out_0.INIT = 1'b0;
  X_SFF DLX_MEMinst_reg_dst_out_0 (
    .I(DLX_EXinst_reg_dst_out[0]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_MEMinst_reg_dst_out[0])
  );
  defparam DLX_MEMinst_reg_dst_out_1.INIT = 1'b0;
  X_SFF DLX_MEMinst_reg_dst_out_1 (
    .I(DLX_EXinst_reg_dst_out[1]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_MEMinst_reg_dst_out[1])
  );
  defparam DLX_MEMinst_reg_dst_out_2.INIT = 1'b0;
  X_SFF DLX_MEMinst_reg_dst_out_2 (
    .I(DLX_EXinst_reg_dst_out[2]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_MEMinst_reg_dst_out[2])
  );
  defparam DLX_EXinst_reg_out_B_EX_26.INIT = 1'b0;
  X_SFF DLX_EXinst_reg_out_B_EX_26 (
    .I(DLX_EXinst__n0008[26]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_reg_out_B_EX[26])
  );
  defparam DLX_EXinst_mem_write_EX_3799.INIT = 1'b0;
  X_SFF DLX_EXinst_mem_write_EX_3799 (
    .I(DLX_IDinst_mem_write),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_mem_write_EX)
  );
  defparam DLX_EXinst_reg_out_B_EX_18.INIT = 1'b0;
  X_SFF DLX_EXinst_reg_out_B_EX_18 (
    .I(DLX_EXinst__n0008[18]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_reg_out_B_EX[18])
  );
  defparam DLX_IDinst_rt_addr_4.INIT = 1'b0;
  X_SFF DLX_IDinst_rt_addr_4 (
    .I(DLX_IDinst__n0135[4]),
    .CE(DLX_IDinst__n0116),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_IDinst__n0115),
    .O(DLX_IDinst_rt_addr[4])
  );
  defparam DLX_EXinst_ALU_result_31.INIT = 1'b0;
  X_SFF DLX_EXinst_ALU_result_31 (
    .I(CHOICE5867),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE5811),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_ALU_result[31])
  );
  defparam DLX_IDinst_rd_addr_4.INIT = 1'b0;
  X_SFF DLX_IDinst_rd_addr_4 (
    .I(DLX_IDinst__n0136[4]),
    .CE(DLX_IDinst__n0116),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_IDinst__n0115),
    .O(DLX_IDinst_rd_addr[4])
  );
  defparam DLX_IDinst_rd_addr_3.INIT = 1'b0;
  X_SFF DLX_IDinst_rd_addr_3 (
    .I(DLX_IDinst__n0136[3]),
    .CE(DLX_IDinst__n0116),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_IDinst__n0115),
    .O(DLX_IDinst_rd_addr[3])
  );
  defparam DLX_IDinst_current_IR_21.INIT = 1'b0;
  X_SFF DLX_IDinst_current_IR_21 (
    .I(\DLX_IDinst_current_IR<21>/FROM ),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_current_IR[21])
  );
  defparam DLX_IDinst_EPC_1.INIT = 1'b0;
  X_SFF DLX_IDinst_EPC_1 (
    .I(DLX_IFinst_NPC[1]),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_EPC[1])
  );
  defparam DLX_IDinst_EPC_7.INIT = 1'b0;
  X_SFF DLX_IDinst_EPC_7 (
    .I(DLX_IFinst_NPC[7]),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_EPC[7])
  );
  defparam DLX_EXinst_ALU_result_1_1_3800.INIT = 1'b0;
  X_SFF DLX_EXinst_ALU_result_1_1_3800 (
    .I(\DLX_EXinst_ALU_result<1>/GROM ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE5717),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_ALU_result_1_1)
  );
  defparam DLX_IDinst_EPC_8.INIT = 1'b0;
  X_SFF DLX_IDinst_EPC_8 (
    .I(DLX_IFinst_NPC[8]),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_EPC[8])
  );
  defparam DLX_EXinst_ALU_result_1.INIT = 1'b0;
  X_SFF DLX_EXinst_ALU_result_1 (
    .I(N162854),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE5717),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_ALU_result[1])
  );
  defparam DLX_IDinst_rd_addr_0.INIT = 1'b0;
  X_SFF DLX_IDinst_rd_addr_0 (
    .I(DLX_IDinst__n0136[0]),
    .CE(DLX_IDinst__n0116),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_IDinst__n0115),
    .O(DLX_IDinst_rd_addr[0])
  );
  defparam DLX_IDinst_Imm_5.INIT = 1'b0;
  X_SFF DLX_IDinst_Imm_5 (
    .I(DLX_IDinst__n0129),
    .CE(DLX_IDinst__n0116),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_IDinst__n0115),
    .O(\DLX_IDinst_Imm[5] )
  );
  defparam DLX_IDinst_rd_addr_1.INIT = 1'b0;
  X_SFF DLX_IDinst_rd_addr_1 (
    .I(DLX_IDinst__n0136[1]),
    .CE(DLX_IDinst__n0116),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_IDinst__n0115),
    .O(DLX_IDinst_rd_addr[1])
  );
  defparam DLX_IDinst_rd_addr_2.INIT = 1'b0;
  X_SFF DLX_IDinst_rd_addr_2 (
    .I(DLX_IDinst__n0136[2]),
    .CE(DLX_IDinst__n0116),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_IDinst__n0115),
    .O(DLX_IDinst_rd_addr[2])
  );
  defparam DLX_IDinst_current_IR_16.INIT = 1'b0;
  X_SFF DLX_IDinst_current_IR_16 (
    .I(\DLX_IDinst_current_IR<16>/FROM ),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_current_IR[16])
  );
  defparam DLX_EXinst_reg_out_B_EX_31.INIT = 1'b0;
  X_SFF DLX_EXinst_reg_out_B_EX_31 (
    .I(DLX_EXinst__n0008[31]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_reg_out_B_EX[31])
  );
  defparam DLX_EXinst_reg_out_B_EX_0.INIT = 1'b0;
  X_SFF DLX_EXinst_reg_out_B_EX_0 (
    .I(DLX_IDinst_reg_out_B[0]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_reg_out_B_EX[0])
  );
  defparam DLX_EXinst_word_3801.INIT = 1'b0;
  X_SFF DLX_EXinst_word_3801 (
    .I(DLX_EXinst__n0011),
    .CE(DLX_EXinst__n0144),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_EXinst_word)
  );
  defparam DLX_EXinst_opcode_of_EX_reg_5.INIT = 1'b0;
  X_SFF DLX_EXinst_opcode_of_EX_reg_5 (
    .I(DLX_IDinst_IR_opcode_field[5]),
    .CE(DLX_EXinst__n0144),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_EXinst_opcode_of_EX_reg[5])
  );
  defparam DLX_EXinst_byte_3802.INIT = 1'b0;
  X_SFF DLX_EXinst_byte_3802 (
    .I(DLX_EXinst__n0010),
    .CE(DLX_EXinst__n0144),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_EXinst_byte)
  );
  defparam DLX_EXinst_ALU_result_9_1_3803.INIT = 1'b0;
  X_SFF DLX_EXinst_ALU_result_9_1_3803 (
    .I(\DLX_EXinst_ALU_result<9>/GROM ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(N136886),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_ALU_result_9_1)
  );
  defparam DLX_EXinst_ALU_result_9.INIT = 1'b0;
  X_SFF DLX_EXinst_ALU_result_9 (
    .I(N162810),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(N136886),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_ALU_result[9])
  );
  defparam DLX_EXinst_ALU_result_2_1_3804.INIT = 1'b0;
  X_SFF DLX_EXinst_ALU_result_2_1_3804 (
    .I(\DLX_EXinst_ALU_result<2>/GROM ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE5538),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_ALU_result_2_1)
  );
  defparam DLX_EXinst_ALU_result_2.INIT = 1'b0;
  X_SFF DLX_EXinst_ALU_result_2 (
    .I(N162841),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE5538),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_ALU_result[2])
  );
  defparam DLX_IDinst_mem_to_reg_3805.INIT = 1'b0;
  X_SFF DLX_IDinst_mem_to_reg_3805 (
    .I(DLX_IDinst__n0139),
    .CE(DLX_IDinst__n0116),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_IDinst__n0115),
    .O(DLX_IDinst_mem_to_reg)
  );
  defparam DLX_EXinst_reg_out_B_EX_15.INIT = 1'b0;
  X_SFF DLX_EXinst_reg_out_B_EX_15 (
    .I(DLX_EXinst__n0008[15]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_reg_out_B_EX[15])
  );
  defparam DLX_EXinst_reg_out_B_EX_2.INIT = 1'b0;
  X_SFF DLX_EXinst_reg_out_B_EX_2 (
    .I(DLX_IDinst_reg_out_B_2_1),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_reg_out_B_EX[2])
  );
  defparam DLX_IDinst_RegFile_10_11_3806.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_10_11_3806 (
    .I(\DLX_IDinst_RegFile_10_11/GROM ),
    .CE(DLX_IDinst__n0570),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_10_11)
  );
  defparam DLX_IDinst_RegFile_10_13_3807.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_10_13_3807 (
    .I(\DLX_IDinst_RegFile_10_13/GROM ),
    .CE(DLX_IDinst__n0570),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_10_13)
  );
  defparam DLX_IDinst_RegFile_10_12_3808.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_10_12_3808 (
    .I(\DLX_IDinst_RegFile_10_12/GROM ),
    .CE(DLX_IDinst__n0570),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_10_12)
  );
  defparam DLX_IDinst_RegFile_10_14_3809.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_10_14_3809 (
    .I(\DLX_IDinst_RegFile_10_14/GROM ),
    .CE(DLX_IDinst__n0570),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_10_14)
  );
  defparam DLX_IDinst_RegFile_10_15_3810.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_10_15_3810 (
    .I(\DLX_IDinst_RegFile_10_15/GROM ),
    .CE(DLX_IDinst__n0570),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_10_15)
  );
  defparam DLX_IDinst_RegFile_0_8_3811.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_0_8_3811 (
    .I(\DLX_IDinst_RegFile_0_8/GROM ),
    .CE(DLX_IDinst__n0550),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_0_8)
  );
  defparam DLX_IDinst_RegFile_0_9_3812.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_0_9_3812 (
    .I(\DLX_IDinst_RegFile_0_9/GROM ),
    .CE(DLX_IDinst__n0550),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_0_9)
  );
  defparam DLX_IDinst_RegFile_10_10_3813.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_10_10_3813 (
    .I(\DLX_IDinst_RegFile_10_10/GROM ),
    .CE(DLX_IDinst__n0570),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_10_10)
  );
  defparam DLX_EXinst_ALU_result_3_1_3814.INIT = 1'b0;
  X_SFF DLX_EXinst_ALU_result_3_1_3814 (
    .I(\DLX_EXinst_ALU_result<3>/GROM ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE5462),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_ALU_result_3_1)
  );
  defparam DLX_EXinst_ALU_result_3.INIT = 1'b0;
  X_SFF DLX_EXinst_ALU_result_3 (
    .I(N162860),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE5462),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_ALU_result[3])
  );
  defparam DLX_EXinst_opcode_of_EX_reg_0.INIT = 1'b0;
  X_SFF DLX_EXinst_opcode_of_EX_reg_0 (
    .I(DLX_IDinst_IR_opcode_field[0]),
    .CE(DLX_EXinst__n0144),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_EXinst_opcode_of_EX_reg[0])
  );
  defparam DLX_EXinst_opcode_of_EX_reg_1.INIT = 1'b0;
  X_SFF DLX_EXinst_opcode_of_EX_reg_1 (
    .I(DLX_IDinst_IR_opcode_field[1]),
    .CE(DLX_EXinst__n0144),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_EXinst_opcode_of_EX_reg[1])
  );
  defparam DLX_EXinst_opcode_of_EX_reg_2.INIT = 1'b0;
  X_SFF DLX_EXinst_opcode_of_EX_reg_2 (
    .I(DLX_IDinst_IR_opcode_field[2]),
    .CE(DLX_EXinst__n0144),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_EXinst_opcode_of_EX_reg[2])
  );
  defparam DLX_EXinst_opcode_of_EX_reg_3.INIT = 1'b0;
  X_SFF DLX_EXinst_opcode_of_EX_reg_3 (
    .I(DLX_IDinst_IR_opcode_field[3]),
    .CE(DLX_EXinst__n0144),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_EXinst_opcode_of_EX_reg[3])
  );
  defparam DLX_EXinst_mem_read_EX_3815.INIT = 1'b0;
  X_SFF DLX_EXinst_mem_read_EX_3815 (
    .I(\DM_read/OD ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_mem_read_EX)
  );
  defparam DLX_EXinst_opcode_of_EX_reg_4.INIT = 1'b0;
  X_SFF DLX_EXinst_opcode_of_EX_reg_4 (
    .I(DLX_IDinst_IR_opcode_field[4]),
    .CE(DLX_EXinst__n0144),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_EXinst_opcode_of_EX_reg[4])
  );
  defparam DLX_IDinst_CLI_1_3816.INIT = 1'b0;
  X_SFF DLX_IDinst_CLI_1_3816 (
    .I(\CLI/OD ),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_CLI_1)
  );
  defparam DLX_EXinst_mem_write_EX_1_3817.INIT = 1'b0;
  X_SFF DLX_EXinst_mem_write_EX_1_3817 (
    .I(\DM_write/OD ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_mem_write_EX_1)
  );
  defparam DLX_IFinst_NPC_0_1_3818.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_0_1_3818 (
    .I(\NPC_eff<0>/OD ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC_0_1)
  );
  defparam DLX_IFinst_NPC_1_1_3819.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_1_1_3819 (
    .I(\NPC_eff<1>/OD ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC_1_1)
  );
  defparam vga_top_vga1_hsyncout_3820.INIT = 1'b1;
  X_SFF vga_top_vga1_hsyncout_3820 (
    .I(\hsync/LOGIC_ZERO ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GSR),
    .RST(GND),
    .SSET(vga_top_vga1__n0010),
    .SRST(GND),
    .O(vga_top_vga1_hsyncout)
  );
  defparam DLX_IDinst_stall_1_3821.INIT = 1'b0;
  X_SFF DLX_IDinst_stall_1_3821 (
    .I(\stall/OD ),
    .CE(DLX_IDinst__n0614),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IDinst_stall_1)
  );
  defparam vga_top_vga1_vsyncout_3822.INIT = 1'b1;
  X_SFF vga_top_vga1_vsyncout_3822 (
    .I(\vsync/LOGIC_ZERO ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GSR),
    .RST(GND),
    .SSET(vga_top_vga1__n0011),
    .SRST(GND),
    .O(vga_top_vga1_vsyncout)
  );
  defparam DLX_IFinst_NPC_2_1_3823.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_2_1_3823 (
    .I(\NPC_eff<2>/OD ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC_2_1)
  );
  defparam DLX_IFinst_NPC_3_1_3824.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_3_1_3824 (
    .I(\NPC_eff<3>/OD ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC_3_1)
  );
  defparam DLX_IFinst_NPC_4_1_3825.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_4_1_3825 (
    .I(\NPC_eff<4>/OD ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC_4_1)
  );
  defparam DLX_IFinst_NPC_5_1_3826.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_5_1_3826 (
    .I(\NPC_eff<5>/OD ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC_5_1)
  );
  defparam DLX_IFinst_NPC_6_1_3827.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_6_1_3827 (
    .I(\NPC_eff<6>/OD ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC_6_1)
  );
  defparam DLX_IFinst_NPC_7_1_3828.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_7_1_3828 (
    .I(\NPC_eff<7>/OD ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC_7_1)
  );
  defparam DLX_IFinst_NPC_8_1_3829.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_8_1_3829 (
    .I(\NPC_eff<8>/OD ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC_8_1)
  );
  defparam DLX_IFinst_NPC_9_1_3830.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_9_1_3830 (
    .I(\NPC_eff<9>/OD ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC_9_1)
  );
  defparam DLX_IFinst_NPC_10_1_3831.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_10_1_3831 (
    .I(\NPC_eff<10>/OD ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC_10_1)
  );
  defparam DLX_IFinst_NPC_11_1_3832.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_11_1_3832 (
    .I(\NPC_eff<11>/OD ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC_11_1)
  );
  defparam DLX_IFinst_NPC_12_1_3833.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_12_1_3833 (
    .I(\NPC_eff<12>/OD ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC_12_1)
  );
  defparam DLX_IFinst_NPC_13_1_3834.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_13_1_3834 (
    .I(\NPC_eff<13>/OD ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC_13_1)
  );
  defparam DLX_IFinst_NPC_14_1_3835.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_14_1_3835 (
    .I(\NPC_eff<14>/OD ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC_14_1)
  );
  defparam DLX_IFinst_NPC_15_1_3836.INIT = 1'b0;
  X_SFF DLX_IFinst_NPC_15_1_3836 (
    .I(\NPC_eff<15>/OD ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_NPC_15_1)
  );
  defparam DLX_EXinst_reg_out_B_EX_0_1_3837.INIT = 1'b0;
  X_SFF DLX_EXinst_reg_out_B_EX_0_1_3837 (
    .I(\DM_write_data<0>/OD ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_reg_out_B_EX_0_1)
  );
  defparam DLX_IDinst_branch_sig_1_3838.INIT = 1'b0;
  X_SFF DLX_IDinst_branch_sig_1_3838 (
    .I(\branch_sig/OD ),
    .CE(DLX_IDinst__n0116),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_IDinst__n0115),
    .O(DLX_IDinst_branch_sig_1)
  );
  defparam DLX_IDinst_RegFile_1_4_3839.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_1_4_3839 (
    .I(DLX_MEMinst_RF_data_in[4]),
    .CE(DLX_IDinst__n0552),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_1_4)
  );
  defparam DLX_IDinst_RegFile_10_0_3840.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_10_0_3840 (
    .I(DLX_MEMinst_RF_data_in[0]),
    .CE(DLX_IDinst__n0570),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_10_0)
  );
  defparam DLX_EXinst_ALU_result_5_1_3841.INIT = 1'b0;
  X_SFF DLX_EXinst_ALU_result_5_1_3841 (
    .I(\DLX_EXinst_ALU_result_5_1/F5MUX ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(N136886),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_ALU_result_5_1)
  );
  defparam DLX_IDinst_RegFile_30_10_3842.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_30_10_3842 (
    .I(DLX_IDinst_WB_data_eff[10]),
    .CE(DLX_IDinst__n0610),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_30_10)
  );
  defparam DLX_EXinst_ALU_result_6_1_3843.INIT = 1'b0;
  X_SFF DLX_EXinst_ALU_result_6_1_3843 (
    .I(\DLX_EXinst_ALU_result_6_1/F5MUX ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(N136886),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_ALU_result_6_1)
  );
  defparam DLX_EXinst_ALU_result_7_1_3844.INIT = 1'b0;
  X_SFF DLX_EXinst_ALU_result_7_1_3844 (
    .I(\DLX_EXinst_ALU_result_7_1/F5MUX ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(N136886),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_ALU_result_7_1)
  );
  defparam DLX_IFinst_IR_curr_4.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_4 (
    .I(IR[4]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[4])
  );
  defparam DLX_IDinst_RegFile_2_31_3845.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_2_31_3845 (
    .I(DLX_IDinst_WB_data_eff[31]),
    .CE(DLX_IDinst__n0554),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_2_31)
  );
  defparam DLX_IFinst_IR_previous_21.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_21 (
    .I(DLX_IFinst_IR_latched[21]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[21])
  );
  defparam DLX_IFinst_IR_latched_9.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_latched_9 (
    .I(DLX_IFinst__n0003[9]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_latched[9])
  );
  defparam DLX_IDinst_RegFile_3_12_3846.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_3_12_3846 (
    .I(DLX_IDinst_WB_data_eff[12]),
    .CE(DLX_IDinst__n0556),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_3_12)
  );
  defparam DLX_IDinst_RegFile_10_3_3847.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_10_3_3847 (
    .I(DLX_MEMinst_RF_data_in[3]),
    .CE(DLX_IDinst__n0570),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_10_3)
  );
  defparam DLX_IDinst_RegFile_2_28_3848.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_2_28_3848 (
    .I(DLX_IDinst_WB_data_eff[28]),
    .CE(DLX_IDinst__n0554),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_2_28)
  );
  defparam DLX_IFinst_IR_previous_1.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_1 (
    .I(DLX_IFinst_IR_latched[1]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[1])
  );
  defparam DLX_IDinst_RegFile_14_21_3849.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_14_21_3849 (
    .I(DLX_IDinst_WB_data_eff[21]),
    .CE(DLX_IDinst__n0578),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_14_21)
  );
  defparam DLX_IFinst_IR_previous_24.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_24 (
    .I(DLX_IFinst_IR_latched[24]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[24])
  );
  defparam DLX_IDinst_RegFile_2_20_3850.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_2_20_3850 (
    .I(DLX_IDinst_WB_data_eff[20]),
    .CE(DLX_IDinst__n0554),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_2_20)
  );
  defparam DLX_IDinst_RegFile_26_0_3851.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_26_0_3851 (
    .I(DLX_MEMinst_RF_data_in[0]),
    .CE(DLX_IDinst__n0602),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_26_0)
  );
  defparam DLX_IDinst_RegFile_17_7_3852.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_17_7_3852 (
    .I(DLX_MEMinst_RF_data_in[7]),
    .CE(DLX_IDinst__n0584),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_17_7)
  );
  defparam DLX_IFinst_IR_previous_4.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_previous_4 (
    .I(DLX_IFinst_IR_latched[4]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_previous[4])
  );
  defparam DLX_IDinst_RegFile_14_10_3853.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_14_10_3853 (
    .I(DLX_IDinst_WB_data_eff[10]),
    .CE(DLX_IDinst__n0578),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_14_10)
  );
  defparam DLX_IDinst_RegFile_11_0_3854.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_11_0_3854 (
    .I(DLX_MEMinst_RF_data_in[0]),
    .CE(DLX_IDinst__n0572),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_11_0)
  );
  defparam DLX_IDinst_RegFile_14_22_3855.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_14_22_3855 (
    .I(DLX_IDinst_WB_data_eff[22]),
    .CE(DLX_IDinst__n0578),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_14_22)
  );
  defparam vga_top_vga1_gridvcounter_1.INIT = 1'b0;
  X_SFF vga_top_vga1_gridvcounter_1 (
    .I(vga_top_vga1_gridvcounter__n0000[1]),
    .CE(vga_top_vga1_N112931),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0014),
    .O(vga_top_vga1_gridvcounter[1])
  );
  defparam vga_top_vga1_gridvcounter_3.INIT = 1'b0;
  X_SFF vga_top_vga1_gridvcounter_3 (
    .I(vga_top_vga1_gridvcounter__n0000[3]),
    .CE(vga_top_vga1_N112931),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0014),
    .O(vga_top_vga1_gridvcounter[3])
  );
  defparam vga_top_vga1_gridvcounter_5.INIT = 1'b0;
  X_SFF vga_top_vga1_gridvcounter_5 (
    .I(vga_top_vga1_gridvcounter__n0000[5]),
    .CE(vga_top_vga1_N112931),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0014),
    .O(vga_top_vga1_gridvcounter[5])
  );
  defparam vga_top_vga1_gridvcounter_0.INIT = 1'b0;
  X_SFF vga_top_vga1_gridvcounter_0 (
    .I(vga_top_vga1_gridvcounter_Madd__n0000_inst_lut2_0),
    .CE(vga_top_vga1_N112931),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0014),
    .O(vga_top_vga1_gridvcounter[0])
  );
  defparam DLX_EXinst_ALU_result_15.INIT = 1'b0;
  X_SFF DLX_EXinst_ALU_result_15 (
    .I(N162847),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE4287),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_ALU_result[15])
  );
  defparam DLX_MEMinst_opcode_of_WB_3.INIT = 1'b0;
  X_SFF DLX_MEMinst_opcode_of_WB_3 (
    .I(DLX_EXinst_opcode_of_EX_reg[3]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_MEMinst_opcode_of_WB[3])
  );
  defparam DLX_IFinst_IR_latched_10.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_latched_10 (
    .I(DLX_IFinst__n0003[10]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_latched[10])
  );
  defparam DLX_IFinst_IR_latched_11.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_latched_11 (
    .I(DLX_IFinst__n0003[11]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_latched[11])
  );
  defparam DLX_IFinst_IR_latched_20.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_latched_20 (
    .I(DLX_IFinst__n0003[20]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_latched[20])
  );
  defparam DLX_IFinst_IR_latched_12.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_latched_12 (
    .I(DLX_IFinst__n0003[12]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_latched[12])
  );
  defparam DLX_MEMinst_RF_data_in_13.INIT = 1'b0;
  X_SFF DLX_MEMinst_RF_data_in_13 (
    .I(DLX_MEMinst__n0000[13]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_MEMinst_RF_data_in[13])
  );
  defparam DLX_MEMinst_RF_data_in_25.INIT = 1'b0;
  X_SFF DLX_MEMinst_RF_data_in_25 (
    .I(DLX_MEMinst__n0000[25]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_MEMinst_RF_data_in[25])
  );
  defparam DLX_MEMinst_RF_data_in_23.INIT = 1'b0;
  X_SFF DLX_MEMinst_RF_data_in_23 (
    .I(DLX_MEMinst__n0000[23]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_MEMinst_RF_data_in[23])
  );
  defparam DLX_MEMinst_RF_data_in_30.INIT = 1'b0;
  X_SFF DLX_MEMinst_RF_data_in_30 (
    .I(DLX_MEMinst__n0000[30]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_MEMinst_RF_data_in[30])
  );
  defparam DLX_MEMinst_RF_data_in_22.INIT = 1'b0;
  X_SFF DLX_MEMinst_RF_data_in_22 (
    .I(DLX_MEMinst__n0000[22]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_MEMinst_RF_data_in[22])
  );
  defparam DLX_MEMinst_RF_data_in_14.INIT = 1'b0;
  X_SFF DLX_MEMinst_RF_data_in_14 (
    .I(DLX_MEMinst__n0000[14]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_MEMinst_RF_data_in[14])
  );
  defparam DLX_MEMinst_RF_data_in_19.INIT = 1'b0;
  X_SFF DLX_MEMinst_RF_data_in_19 (
    .I(DLX_MEMinst__n0000[19]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_MEMinst_RF_data_in[19])
  );
  defparam DLX_MEMinst_RF_data_in_15.INIT = 1'b0;
  X_SFF DLX_MEMinst_RF_data_in_15 (
    .I(DLX_MEMinst__n0000[15]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_MEMinst_RF_data_in[15])
  );
  defparam DLX_MEMinst_RF_data_in_18.INIT = 1'b0;
  X_SFF DLX_MEMinst_RF_data_in_18 (
    .I(DLX_MEMinst__n0000[18]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_MEMinst_RF_data_in[18])
  );
  defparam DLX_MEMinst_RF_data_in_31.INIT = 1'b0;
  X_SFF DLX_MEMinst_RF_data_in_31 (
    .I(DLX_MEMinst__n0000[31]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_MEMinst_RF_data_in[31])
  );
  defparam DLX_MEMinst_RF_data_in_17.INIT = 1'b0;
  X_SFF DLX_MEMinst_RF_data_in_17 (
    .I(DLX_MEMinst__n0000[17]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_MEMinst_RF_data_in[17])
  );
  defparam DLX_MEMinst_RF_data_in_16.INIT = 1'b0;
  X_SFF DLX_MEMinst_RF_data_in_16 (
    .I(DLX_MEMinst__n0000[16]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_MEMinst_RF_data_in[16])
  );
  defparam DLX_IDinst_rt_addr_1.INIT = 1'b0;
  X_SFF DLX_IDinst_rt_addr_1 (
    .I(DLX_IDinst__n0135[1]),
    .CE(DLX_IDinst__n0116),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_IDinst__n0115),
    .O(DLX_IDinst_rt_addr[1])
  );
  defparam DLX_MEMinst_RF_data_in_9.INIT = 1'b0;
  X_SFF DLX_MEMinst_RF_data_in_9 (
    .I(DLX_MEMinst__n0000[9]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_MEMinst_RF_data_in[9])
  );
  defparam DLX_IDinst_rt_addr_0.INIT = 1'b0;
  X_SFF DLX_IDinst_rt_addr_0 (
    .I(DLX_IDinst__n0135[0]),
    .CE(DLX_IDinst__n0116),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_IDinst__n0115),
    .O(DLX_IDinst_rt_addr[0])
  );
  defparam DLX_IFinst_IR_latched_24.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_latched_24 (
    .I(DLX_IFinst__n0003[24]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_latched[24])
  );
  defparam DLX_IFinst_IR_latched_16.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_latched_16 (
    .I(DLX_IFinst__n0003[16]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_latched[16])
  );
  defparam DLX_IFinst_IR_latched_17.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_latched_17 (
    .I(DLX_IFinst__n0003[17]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_latched[17])
  );
  defparam DLX_IFinst_IR_latched_25.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_latched_25 (
    .I(DLX_IFinst__n0003[25]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_latched[25])
  );
  defparam DLX_IFinst_IR_latched_18.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_latched_18 (
    .I(DLX_IFinst__n0003[18]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_latched[18])
  );
  defparam DLX_IFinst_IR_latched_26.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_latched_26 (
    .I(DLX_IFinst__n0003[26]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_latched[26])
  );
  defparam DLX_IFinst_IR_latched_19.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_latched_19 (
    .I(DLX_IFinst__n0003[19]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_latched[19])
  );
  defparam DLX_IFinst_IR_latched_27.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_latched_27 (
    .I(DLX_IFinst__n0003[27]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_latched[27])
  );
  defparam DLX_IDinst_RegFile_30_17_3856.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_30_17_3856 (
    .I(DLX_IDinst_WB_data_eff[17]),
    .CE(DLX_IDinst__n0610),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_30_17)
  );
  defparam DLX_IDinst_RegFile_14_17_3857.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_14_17_3857 (
    .I(DLX_IDinst_WB_data_eff[17]),
    .CE(DLX_IDinst__n0578),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_14_17)
  );
  defparam DLX_IDinst_RegFile_11_3_3858.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_11_3_3858 (
    .I(DLX_MEMinst_RF_data_in[3]),
    .CE(DLX_IDinst__n0572),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_11_3)
  );
  defparam DLX_IFinst_IR_latched_13.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_latched_13 (
    .I(DLX_IFinst__n0003[13]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_latched[13])
  );
  defparam DLX_IFinst_IR_latched_21.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_latched_21 (
    .I(DLX_IFinst__n0003[21]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_latched[21])
  );
  defparam DLX_IFinst_IR_latched_30.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_latched_30 (
    .I(DLX_IFinst__n0003[30]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_latched[30])
  );
  defparam DLX_IFinst_IR_latched_14.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_latched_14 (
    .I(DLX_IFinst__n0003[14]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_latched[14])
  );
  defparam DLX_IFinst_IR_latched_22.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_latched_22 (
    .I(DLX_IFinst__n0003[22]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_latched[22])
  );
  defparam DLX_IFinst_IR_latched_23.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_latched_23 (
    .I(DLX_IFinst__n0003[23]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_latched[23])
  );
  defparam DLX_IFinst_IR_latched_15.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_latched_15 (
    .I(DLX_IFinst__n0003[15]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_latched[15])
  );
  defparam DLX_IFinst_IR_latched_31.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_latched_31 (
    .I(DLX_IFinst__n0003[31]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_latched[31])
  );
  defparam DLX_IDinst_RegFile_30_20_3859.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_30_20_3859 (
    .I(DLX_IDinst_WB_data_eff[20]),
    .CE(DLX_IDinst__n0610),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_30_20)
  );
  defparam DLX_IDinst_RegFile_11_27_3860.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_11_27_3860 (
    .I(DLX_IDinst_WB_data_eff[27]),
    .CE(DLX_IDinst__n0572),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_11_27)
  );
  defparam DLX_IFinst_IR_latched_28.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_latched_28 (
    .I(DLX_IFinst__n0003[28]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_latched[28])
  );
  defparam DLX_IFinst_IR_latched_29.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_latched_29 (
    .I(DLX_IFinst__n0003[29]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_2),
    .O(DLX_IFinst_IR_latched[29])
  );
  defparam DLX_IDinst_RegFile_22_14_3861.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_22_14_3861 (
    .I(DLX_IDinst_WB_data_eff[14]),
    .CE(DLX_IDinst__n0594),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_22_14)
  );
  defparam vga_top_vga1_vcounter_1.INIT = 1'b0;
  X_SFF vga_top_vga1_vcounter_1 (
    .I(vga_top_vga1_vcounter__n0000[1]),
    .CE(N145733),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0007),
    .O(vga_top_vga1_vcounter[1])
  );
  defparam vga_top_vga1_vcounter_3.INIT = 1'b0;
  X_SFF vga_top_vga1_vcounter_3 (
    .I(vga_top_vga1_vcounter__n0000[3]),
    .CE(N145733),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0007),
    .O(vga_top_vga1_vcounter[3])
  );
  defparam vga_top_vga1_vcounter_0.INIT = 1'b0;
  X_SFF vga_top_vga1_vcounter_0 (
    .I(vga_top_vga1_vcounter_Madd__n0000_inst_lut2_9),
    .CE(N145733),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0007),
    .O(vga_top_vga1_vcounter[0])
  );
  defparam vga_top_vga1_vcounter_5.INIT = 1'b0;
  X_SFF vga_top_vga1_vcounter_5 (
    .I(vga_top_vga1_vcounter__n0000[5]),
    .CE(N145733),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0007),
    .O(vga_top_vga1_vcounter[5])
  );
  defparam vga_top_vga1_vcounter_7.INIT = 1'b0;
  X_SFF vga_top_vga1_vcounter_7 (
    .I(vga_top_vga1_vcounter__n0000[7]),
    .CE(N145733),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0007),
    .O(vga_top_vga1_vcounter[7])
  );
  defparam vga_top_vga1_vcounter_2.INIT = 1'b0;
  X_SFF vga_top_vga1_vcounter_2 (
    .I(vga_top_vga1_vcounter__n0000[2]),
    .CE(N145733),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0007),
    .O(vga_top_vga1_vcounter[2])
  );
  defparam vga_top_vga1_vcounter_4.INIT = 1'b0;
  X_SFF vga_top_vga1_vcounter_4 (
    .I(vga_top_vga1_vcounter__n0000[4]),
    .CE(N145733),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0007),
    .O(vga_top_vga1_vcounter[4])
  );
  defparam vga_top_vga1_vcounter_6.INIT = 1'b0;
  X_SFF vga_top_vga1_vcounter_6 (
    .I(vga_top_vga1_vcounter__n0000[6]),
    .CE(N145733),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0007),
    .O(vga_top_vga1_vcounter[6])
  );
  defparam vga_top_vga1_vcounter_9.INIT = 1'b0;
  X_SFF vga_top_vga1_vcounter_9 (
    .I(vga_top_vga1_vcounter__n0000[9]),
    .CE(N145733),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0007),
    .O(vga_top_vga1_vcounter[9])
  );
  defparam vga_top_vga1_vcounter_8.INIT = 1'b0;
  X_SFF vga_top_vga1_vcounter_8 (
    .I(vga_top_vga1_vcounter__n0000[8]),
    .CE(N145733),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0007),
    .O(vga_top_vga1_vcounter[8])
  );
  defparam DLX_IDinst_RegFile_14_12_3862.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_14_12_3862 (
    .I(DLX_IDinst_WB_data_eff[12]),
    .CE(DLX_IDinst__n0578),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_14_12)
  );
  defparam DLX_IDinst_RegFile_18_3_3863.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_18_3_3863 (
    .I(DLX_MEMinst_RF_data_in[3]),
    .CE(DLX_IDinst__n0586),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_18_3)
  );
  defparam DLX_IDinst_RegFile_30_13_3864.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_30_13_3864 (
    .I(DLX_IDinst_WB_data_eff[13]),
    .CE(DLX_IDinst__n0610),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_30_13)
  );
  defparam DLX_IDinst_RegFile_22_26_3865.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_22_26_3865 (
    .I(DLX_IDinst_WB_data_eff[26]),
    .CE(DLX_IDinst__n0594),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_22_26)
  );
  defparam DLX_IDinst_RegFile_15_11_3866.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_15_11_3866 (
    .I(DLX_IDinst_WB_data_eff[11]),
    .CE(DLX_IDinst__n0580),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_15_11)
  );
  defparam DLX_IDinst_RegFile_3_6_3867.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_3_6_3867 (
    .I(DLX_MEMinst_RF_data_in[6]),
    .CE(DLX_IDinst__n0556),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_3_6)
  );
  defparam DLX_EXinst_reg_out_B_EX_30.INIT = 1'b0;
  X_SFF DLX_EXinst_reg_out_B_EX_30 (
    .I(DLX_EXinst__n0008[30]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_reg_out_B_EX[30])
  );
  defparam DLX_IDinst_RegFile_23_21_3868.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_23_21_3868 (
    .I(DLX_IDinst_WB_data_eff[21]),
    .CE(DLX_IDinst__n0596),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_23_21)
  );
  defparam vga_top_vga1_gridvcounter_2.INIT = 1'b0;
  X_SFF vga_top_vga1_gridvcounter_2 (
    .I(vga_top_vga1_gridvcounter__n0000[2]),
    .CE(vga_top_vga1_N112931),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0014),
    .O(vga_top_vga1_gridvcounter[2])
  );
  defparam vga_top_vga1_gridvcounter_4.INIT = 1'b0;
  X_SFF vga_top_vga1_gridvcounter_4 (
    .I(vga_top_vga1_gridvcounter__n0000[4]),
    .CE(vga_top_vga1_N112931),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0014),
    .O(vga_top_vga1_gridvcounter[4])
  );
  defparam vga_top_vga1_gridvcounter_7.INIT = 1'b0;
  X_SFF vga_top_vga1_gridvcounter_7 (
    .I(vga_top_vga1_gridvcounter__n0000[7]),
    .CE(vga_top_vga1_N112931),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0014),
    .O(vga_top_vga1_gridvcounter[7])
  );
  defparam DLX_IDinst_RegFile_30_27_3869.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_30_27_3869 (
    .I(DLX_IDinst_WB_data_eff[27]),
    .CE(DLX_IDinst__n0610),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_30_27)
  );
  defparam vga_top_vga1_gridvcounter_6.INIT = 1'b0;
  X_SFF vga_top_vga1_gridvcounter_6 (
    .I(vga_top_vga1_gridvcounter__n0000[6]),
    .CE(vga_top_vga1_N112931),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0014),
    .O(vga_top_vga1_gridvcounter[6])
  );
  defparam vga_top_vga1_gridvcounter_8.INIT = 1'b0;
  X_SFF vga_top_vga1_gridvcounter_8 (
    .I(vga_top_vga1_gridvcounter__n0000[8]),
    .CE(vga_top_vga1_N112931),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0014),
    .O(vga_top_vga1_gridvcounter[8])
  );
  defparam DLX_IDinst_RegFile_22_30_3870.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_22_30_3870 (
    .I(DLX_IDinst_WB_data_eff[30]),
    .CE(DLX_IDinst__n0594),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_22_30)
  );
  defparam DLX_IDinst_RegFile_30_22_3871.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_30_22_3871 (
    .I(DLX_IDinst_WB_data_eff[22]),
    .CE(DLX_IDinst__n0610),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_30_22)
  );
  defparam DLX_IDinst_RegFile_1_6_3872.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_1_6_3872 (
    .I(DLX_MEMinst_RF_data_in[6]),
    .CE(DLX_IDinst__n0552),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_1_6)
  );
  defparam DLX_IDinst_RegFile_30_18_3873.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_30_18_3873 (
    .I(DLX_IDinst_WB_data_eff[18]),
    .CE(DLX_IDinst__n0610),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_30_18)
  );
  defparam DLX_IDinst_RegFile_22_23_3874.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_22_23_3874 (
    .I(DLX_IDinst_WB_data_eff[23]),
    .CE(DLX_IDinst__n0594),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_22_23)
  );
  defparam DLX_IDinst_RegFile_23_12_3875.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_23_12_3875 (
    .I(DLX_IDinst_WB_data_eff[12]),
    .CE(DLX_IDinst__n0596),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_23_12)
  );
  defparam DLX_IDinst_RegFile_15_20_3876.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_15_20_3876 (
    .I(DLX_IDinst_WB_data_eff[20]),
    .CE(DLX_IDinst__n0580),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_15_20)
  );
  defparam DLX_IDinst_RegFile_14_16_3877.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_14_16_3877 (
    .I(DLX_IDinst_WB_data_eff[16]),
    .CE(DLX_IDinst__n0578),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_14_16)
  );
  defparam DLX_EXinst_mem_to_reg_EX_3878.INIT = 1'b0;
  X_SFF DLX_EXinst_mem_to_reg_EX_3878 (
    .I(DLX_IDinst_mem_to_reg),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_mem_to_reg_EX)
  );
  defparam DLX_IDinst_RegFile_6_20_3879.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_6_20_3879 (
    .I(DLX_IDinst_WB_data_eff[20]),
    .CE(DLX_IDinst__n0562),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_6_20)
  );
  defparam DLX_IDinst_RegFile_6_12_3880.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_6_12_3880 (
    .I(DLX_IDinst_WB_data_eff[12]),
    .CE(DLX_IDinst__n0562),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_6_12)
  );
  defparam DLX_IDinst_RegFile_1_7_3881.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_1_7_3881 (
    .I(DLX_MEMinst_RF_data_in[7]),
    .CE(DLX_IDinst__n0552),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_1_7)
  );
  defparam DLX_IDinst_RegFile_10_9_3882.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_10_9_3882 (
    .I(DLX_IDinst_WB_data_eff[9]),
    .CE(DLX_IDinst__n0570),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_10_9)
  );
  defparam vga_top_vga1_gridhcounter_3.INIT = 1'b0;
  X_SFF vga_top_vga1_gridhcounter_3 (
    .I(vga_top_vga1_gridhcounter__n0000[3]),
    .CE(vga_top_vga1__n0013),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0012),
    .O(vga_top_vga1_gridhcounter[3])
  );
  defparam vga_top_vga1_gridhcounter_1.INIT = 1'b0;
  X_SFF vga_top_vga1_gridhcounter_1 (
    .I(vga_top_vga1_gridhcounter__n0000[1]),
    .CE(vga_top_vga1__n0013),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0012),
    .O(vga_top_vga1_gridhcounter[1])
  );
  defparam vga_top_vga1_gridhcounter_5.INIT = 1'b0;
  X_SFF vga_top_vga1_gridhcounter_5 (
    .I(vga_top_vga1_gridhcounter__n0000[5]),
    .CE(vga_top_vga1__n0013),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0012),
    .O(vga_top_vga1_gridhcounter[5])
  );
  defparam vga_top_vga1_gridhcounter_0.INIT = 1'b0;
  X_SFF vga_top_vga1_gridhcounter_0 (
    .I(vga_top_vga1_gridhcounter_Madd__n0000_inst_lut2_0),
    .CE(vga_top_vga1__n0013),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0012),
    .O(vga_top_vga1_gridhcounter[0])
  );
  defparam DLX_IDinst_RegFile_14_29_3883.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_14_29_3883 (
    .I(DLX_IDinst_WB_data_eff[29]),
    .CE(DLX_IDinst__n0578),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_14_29)
  );
  defparam vga_top_vga1_gridhcounter_2.INIT = 1'b0;
  X_SFF vga_top_vga1_gridhcounter_2 (
    .I(vga_top_vga1_gridhcounter__n0000[2]),
    .CE(vga_top_vga1__n0013),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0012),
    .O(vga_top_vga1_gridhcounter[2])
  );
  defparam vga_top_vga1_hcounter_1.INIT = 1'b0;
  X_SFF vga_top_vga1_hcounter_1 (
    .I(vga_top_vga1_hcounter__n0000[1]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0006),
    .O(vga_top_vga1_hcounter[1])
  );
  defparam vga_top_vga1_gridhcounter_4.INIT = 1'b0;
  X_SFF vga_top_vga1_gridhcounter_4 (
    .I(vga_top_vga1_gridhcounter__n0000[4]),
    .CE(vga_top_vga1__n0013),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0012),
    .O(vga_top_vga1_gridhcounter[4])
  );
  defparam vga_top_vga1_gridhcounter_7.INIT = 1'b0;
  X_SFF vga_top_vga1_gridhcounter_7 (
    .I(vga_top_vga1_gridhcounter__n0000[7]),
    .CE(vga_top_vga1__n0013),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0012),
    .O(vga_top_vga1_gridhcounter[7])
  );
  defparam vga_top_vga1_gridhcounter_8.INIT = 1'b0;
  X_SFF vga_top_vga1_gridhcounter_8 (
    .I(vga_top_vga1_gridhcounter__n0000[8]),
    .CE(vga_top_vga1__n0013),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0012),
    .O(vga_top_vga1_gridhcounter[8])
  );
  defparam vga_top_vga1_gridhcounter_6.INIT = 1'b0;
  X_SFF vga_top_vga1_gridhcounter_6 (
    .I(vga_top_vga1_gridhcounter__n0000[6]),
    .CE(vga_top_vga1__n0013),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0012),
    .O(vga_top_vga1_gridhcounter[6])
  );
  defparam DLX_IDinst_RegFile_6_13_3884.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_6_13_3884 (
    .I(DLX_IDinst_WB_data_eff[13]),
    .CE(DLX_IDinst__n0562),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_6_13)
  );
  defparam vga_top_vga1_hcounter_3.INIT = 1'b0;
  X_SFF vga_top_vga1_hcounter_3 (
    .I(vga_top_vga1_hcounter__n0000[3]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0006),
    .O(vga_top_vga1_hcounter[3])
  );
  defparam vga_top_vga1_hcounter_0.INIT = 1'b0;
  X_SFF vga_top_vga1_hcounter_0 (
    .I(vga_top_vga1_hcounter_Madd__n0000_inst_lut2_19),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0006),
    .O(vga_top_vga1_hcounter[0])
  );
  defparam vga_top_vga1_hcounter_7.INIT = 1'b0;
  X_SFF vga_top_vga1_hcounter_7 (
    .I(vga_top_vga1_hcounter__n0000[7]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0006),
    .O(vga_top_vga1_hcounter[7])
  );
  defparam vga_top_vga1_hcounter_2.INIT = 1'b0;
  X_SFF vga_top_vga1_hcounter_2 (
    .I(vga_top_vga1_hcounter__n0000[2]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0006),
    .O(vga_top_vga1_hcounter[2])
  );
  defparam vga_top_vga1_hcounter_5.INIT = 1'b0;
  X_SFF vga_top_vga1_hcounter_5 (
    .I(vga_top_vga1_hcounter__n0000[5]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0006),
    .O(vga_top_vga1_hcounter[5])
  );
  defparam vga_top_vga1_hcounter_4.INIT = 1'b0;
  X_SFF vga_top_vga1_hcounter_4 (
    .I(vga_top_vga1_hcounter__n0000[4]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0006),
    .O(vga_top_vga1_hcounter[4])
  );
  defparam vga_top_vga1_hcounter_9.INIT = 1'b0;
  X_SFF vga_top_vga1_hcounter_9 (
    .I(vga_top_vga1_hcounter__n0000[9]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0006),
    .O(vga_top_vga1_hcounter[9])
  );
  defparam vga_top_vga1_hcounter_6.INIT = 1'b0;
  X_SFF vga_top_vga1_hcounter_6 (
    .I(vga_top_vga1_hcounter__n0000[6]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0006),
    .O(vga_top_vga1_hcounter[6])
  );
  defparam vga_top_vga1_hcounter_13.INIT = 1'b0;
  X_SFF vga_top_vga1_hcounter_13 (
    .I(vga_top_vga1_hcounter__n0000[13]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0006),
    .O(vga_top_vga1_hcounter[13])
  );
  defparam vga_top_vga1_hcounter_8.INIT = 1'b0;
  X_SFF vga_top_vga1_hcounter_8 (
    .I(vga_top_vga1_hcounter__n0000[8]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0006),
    .O(vga_top_vga1_hcounter[8])
  );
  defparam vga_top_vga1_hcounter_11.INIT = 1'b0;
  X_SFF vga_top_vga1_hcounter_11 (
    .I(vga_top_vga1_hcounter__n0000[11]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0006),
    .O(vga_top_vga1_hcounter[11])
  );
  defparam vga_top_vga1_hcounter_10.INIT = 1'b0;
  X_SFF vga_top_vga1_hcounter_10 (
    .I(vga_top_vga1_hcounter__n0000[10]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0006),
    .O(vga_top_vga1_hcounter[10])
  );
  defparam vga_top_vga1_hcounter_15.INIT = 1'b0;
  X_SFF vga_top_vga1_hcounter_15 (
    .I(vga_top_vga1_hcounter__n0000[15]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0006),
    .O(vga_top_vga1_hcounter[15])
  );
  defparam vga_top_vga1_hcounter_12.INIT = 1'b0;
  X_SFF vga_top_vga1_hcounter_12 (
    .I(vga_top_vga1_hcounter__n0000[12]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0006),
    .O(vga_top_vga1_hcounter[12])
  );
  defparam vga_top_vga1_hcounter_14.INIT = 1'b0;
  X_SFF vga_top_vga1_hcounter_14 (
    .I(vga_top_vga1_hcounter__n0000[14]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(vga_top_vga1__n0006),
    .O(vga_top_vga1_hcounter[14])
  );
  defparam DLX_IDinst_RegFile_3_14_3885.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_3_14_3885 (
    .I(DLX_IDinst_WB_data_eff[14]),
    .CE(DLX_IDinst__n0556),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_3_14)
  );
  defparam DLX_IDinst_RegFile_18_5_3886.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_18_5_3886 (
    .I(DLX_MEMinst_RF_data_in[5]),
    .CE(DLX_IDinst__n0586),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_18_5)
  );
  defparam DLX_EXinst_reg_write_EX_3887.INIT = 1'b0;
  X_SFF DLX_EXinst_reg_write_EX_3887 (
    .I(DLX_IDinst_reg_write),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_reg_write_EX)
  );
  defparam DLX_IDinst_Cause_Reg_6.INIT = 1'b0;
  X_FF DLX_IDinst_Cause_Reg_6 (
    .I(\DLX_IDinst_Imm[6] ),
    .CE(DLX_IDinst__n0617),
    .CLK(clkdiv),
    .SET(GND),
    .RST(\DLX_IDinst_Cause_Reg<6>/FFY/RST ),
    .O(\DLX_IDinst_Cause_Reg[6] )
  );
  X_BUF \DLX_IDinst_Cause_Reg<6>/FFY/RSTOR  (
    .I(GSR),
    .O(\DLX_IDinst_Cause_Reg<6>/FFY/RST )
  );
  defparam DLX_IDinst_RegFile_3_0_3888.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_3_0_3888 (
    .I(DLX_MEMinst_RF_data_in[0]),
    .CE(DLX_IDinst__n0556),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_3_0)
  );
  defparam DLX_IDinst_RegFile_31_11_3889.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_31_11_3889 (
    .I(DLX_IDinst_WB_data_eff[11]),
    .CE(DLX_IDinst__n0612),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_31_11)
  );
  defparam DLX_EXinst_reg_out_B_EX_3.INIT = 1'b0;
  X_SFF DLX_EXinst_reg_out_B_EX_3 (
    .I(DLX_IDinst_reg_out_B_3_1),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_reg_out_B_EX[3])
  );
  defparam DLX_IDinst_RegFile_3_30_3890.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_3_30_3890 (
    .I(DLX_IDinst_WB_data_eff[30]),
    .CE(DLX_IDinst__n0556),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_3_30)
  );
  defparam DLX_IDinst_RegFile_22_28_3891.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_22_28_3891 (
    .I(DLX_IDinst_WB_data_eff[28]),
    .CE(DLX_IDinst__n0594),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_22_28)
  );
  defparam DLX_IDinst_RegFile_23_14_3892.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_23_14_3892 (
    .I(DLX_IDinst_WB_data_eff[14]),
    .CE(DLX_IDinst__n0596),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_23_14)
  );
  defparam DLX_IDinst_RegFile_26_3_3893.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_26_3_3893 (
    .I(DLX_MEMinst_RF_data_in[3]),
    .CE(DLX_IDinst__n0602),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_7),
    .O(DLX_IDinst_RegFile_26_3)
  );
  defparam DLX_IDinst_RegFile_15_23_3894.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_15_23_3894 (
    .I(DLX_IDinst_WB_data_eff[23]),
    .CE(DLX_IDinst__n0580),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_15_23)
  );
  defparam DLX_IFinst_IR_curr_20.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_20 (
    .I(IR[20]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[20])
  );
  defparam DLX_IDinst_RegFile_31_29_3895.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_31_29_3895 (
    .I(DLX_IDinst_WB_data_eff[29]),
    .CE(DLX_IDinst__n0612),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_31_29)
  );
  defparam DLX_IDinst_RegFile_31_23_3896.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_31_23_3896 (
    .I(DLX_IDinst_WB_data_eff[23]),
    .CE(DLX_IDinst__n0612),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_31_23)
  );
  defparam DLX_IDinst_RegFile_1_8_3897.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_1_8_3897 (
    .I(DLX_IDinst_WB_data_eff[8]),
    .CE(DLX_IDinst__n0552),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_1_8)
  );
  defparam DLX_IDinst_RegFile_24_12_3898.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_24_12_3898 (
    .I(DLX_IDinst_WB_data_eff[12]),
    .CE(DLX_IDinst__n0598),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_24_12)
  );
  defparam DLX_IDinst_RegFile_31_20_3899.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_31_20_3899 (
    .I(DLX_IDinst_WB_data_eff[20]),
    .CE(DLX_IDinst__n0612),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_31_20)
  );
  defparam DLX_IFinst_IR_curr_10.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_10 (
    .I(IR[10]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[10])
  );
  defparam DLX_IDinst_RegFile_30_29_3900.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_30_29_3900 (
    .I(DLX_IDinst_WB_data_eff[29]),
    .CE(DLX_IDinst__n0610),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_30_29)
  );
  defparam DLX_IDinst_RegFile_15_13_3901.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_15_13_3901 (
    .I(DLX_IDinst_WB_data_eff[13]),
    .CE(DLX_IDinst__n0580),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_15_13)
  );
  defparam DLX_IFinst_IR_curr_12.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_12 (
    .I(IR[12]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[12])
  );
  defparam DLX_IDinst_RegFile_15_22_3902.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_15_22_3902 (
    .I(DLX_IDinst_WB_data_eff[22]),
    .CE(DLX_IDinst__n0580),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_15_22)
  );
  defparam DLX_IFinst_IR_curr_11.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_11 (
    .I(IR[11]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[11])
  );
  defparam DLX_IDinst_RegFile_31_31_3903.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_31_31_3903 (
    .I(DLX_IDinst_WB_data_eff[31]),
    .CE(DLX_IDinst__n0612),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_31_31)
  );
  defparam DLX_IDinst_RegFile_31_17_3904.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_31_17_3904 (
    .I(DLX_IDinst_WB_data_eff[17]),
    .CE(DLX_IDinst__n0612),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_31_17)
  );
  defparam DLX_IFinst_IR_curr_21.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_21 (
    .I(IR[21]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[21])
  );
  defparam DLX_IDinst_RegFile_3_23_3905.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_3_23_3905 (
    .I(DLX_IDinst_WB_data_eff[23]),
    .CE(DLX_IDinst__n0556),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_3_23)
  );
  defparam DLX_IDinst_RegFile_7_11_3906.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_7_11_3906 (
    .I(DLX_IDinst_WB_data_eff[11]),
    .CE(DLX_IDinst__n0564),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_7_11)
  );
  defparam DLX_EXinst_reg_out_B_EX_5.INIT = 1'b0;
  X_SFF DLX_EXinst_reg_out_B_EX_5 (
    .I(DLX_IDinst_reg_out_B[5]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_reg_out_B_EX[5])
  );
  defparam DLX_IDinst_RegFile_23_16_3907.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_23_16_3907 (
    .I(DLX_IDinst_WB_data_eff[16]),
    .CE(DLX_IDinst__n0596),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_23_16)
  );
  defparam vga_top_vga1_clockcounter_FFd1_3908.INIT = 1'b0;
  X_SFF vga_top_vga1_clockcounter_FFd1_3908 (
    .I(vga_top_vga1_clockcounter_FFd2),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(vga_top_vga1_clockcounter_FFd1)
  );
  defparam DLX_IDinst_RegFile_6_26_3909.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_6_26_3909 (
    .I(DLX_IDinst_WB_data_eff[26]),
    .CE(DLX_IDinst__n0562),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_4),
    .O(DLX_IDinst_RegFile_6_26)
  );
  defparam vga_top_vga1_clockcounter_FFd2_3910.INIT = 1'b1;
  X_SFF vga_top_vga1_clockcounter_FFd2_3910 (
    .I(vga_top_vga1_clockcounter_FFd1),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GSR),
    .RST(GND),
    .SSET(reset_IBUF_1),
    .SRST(GND),
    .O(vga_top_vga1_clockcounter_FFd2)
  );
  defparam DLX_MEMinst_opcode_of_WB_0.INIT = 1'b0;
  X_SFF DLX_MEMinst_opcode_of_WB_0 (
    .I(DLX_EXinst_opcode_of_EX_reg[0]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_MEMinst_opcode_of_WB[0])
  );
  defparam DLX_MEMinst_opcode_of_WB_4.INIT = 1'b0;
  X_SFF DLX_MEMinst_opcode_of_WB_4 (
    .I(DLX_EXinst_opcode_of_EX_reg[4]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_MEMinst_opcode_of_WB[4])
  );
  defparam DLX_IDinst_RegFile_3_16_3911.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_3_16_3911 (
    .I(DLX_IDinst_WB_data_eff[16]),
    .CE(DLX_IDinst__n0556),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_3_16)
  );
  defparam DLX_IDinst_EPC_29.INIT = 1'b0;
  X_SFF DLX_IDinst_EPC_29 (
    .I(DLX_IFinst_NPC[29]),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_EPC[29])
  );
  defparam DLX_IDinst_RegFile_26_10_3912.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_26_10_3912 (
    .I(DLX_IDinst_WB_data_eff[10]),
    .CE(DLX_IDinst__n0602),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_26_10)
  );
  defparam DLX_IDinst_RegFile_2_25_3913.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_2_25_3913 (
    .I(DLX_IDinst_WB_data_eff[25]),
    .CE(DLX_IDinst__n0554),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_2_25)
  );
  defparam DLX_IFinst_IR_curr_15.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_15 (
    .I(IR[15]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[15])
  );
  defparam DLX_IFinst_IR_curr_31.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_31 (
    .I(IR_MSB_7_OBUF),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[31])
  );
  defparam DLX_IDinst_RegFile_2_30_3914.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_2_30_3914 (
    .I(DLX_IDinst_WB_data_eff[30]),
    .CE(DLX_IDinst__n0554),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_2_30)
  );
  defparam DLX_IFinst_IR_curr_24.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_24 (
    .I(IR_MSB_0_OBUF),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[24])
  );
  defparam DLX_IFinst_IR_curr_16.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_16 (
    .I(IR[16]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[16])
  );
  defparam DLX_IDinst_RegFile_0_6_3915.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_0_6_3915 (
    .I(DLX_MEMinst_RF_data_in[6]),
    .CE(DLX_IDinst__n0550),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_0_6)
  );
  defparam DLX_IFinst_IR_curr_25.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_25 (
    .I(IR_MSB_1_OBUF),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[25])
  );
  defparam DLX_IDinst_RegFile_2_18_3916.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_2_18_3916 (
    .I(DLX_IDinst_WB_data_eff[18]),
    .CE(DLX_IDinst__n0554),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_2_18)
  );
  defparam DLX_IDinst_RegFile_1_19_3917.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_1_19_3917 (
    .I(DLX_IDinst_WB_data_eff[19]),
    .CE(DLX_IDinst__n0552),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_1_19)
  );
  defparam DLX_IDinst_RegFile_3_18_3918.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_3_18_3918 (
    .I(DLX_IDinst_WB_data_eff[18]),
    .CE(DLX_IDinst__n0556),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_3_18)
  );
  defparam DLX_IFinst_IR_curr_6.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_6 (
    .I(IR[6]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[6])
  );
  defparam DLX_IDinst_RegFile_11_19_3919.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_11_19_3919 (
    .I(DLX_IDinst_WB_data_eff[19]),
    .CE(DLX_IDinst__n0572),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_11_19)
  );
  defparam DLX_IDinst_RegFile_20_11_3920.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_20_11_3920 (
    .I(DLX_IDinst_WB_data_eff[11]),
    .CE(DLX_IDinst__n0590),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_20_11)
  );
  defparam DLX_IDinst_RegFile_12_11_3921.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_12_11_3921 (
    .I(DLX_IDinst_WB_data_eff[11]),
    .CE(DLX_IDinst__n0574),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_12_11)
  );
  defparam DLX_IDinst_RegFile_12_20_3922.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_12_20_3922 (
    .I(DLX_IDinst_WB_data_eff[20]),
    .CE(DLX_IDinst__n0574),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_12_20)
  );
  defparam DLX_IDinst_RegFile_20_20_3923.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_20_20_3923 (
    .I(DLX_IDinst_WB_data_eff[20]),
    .CE(DLX_IDinst__n0590),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_20_20)
  );
  defparam DLX_IDinst_RegFile_12_12_3924.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_12_12_3924 (
    .I(DLX_IDinst_WB_data_eff[12]),
    .CE(DLX_IDinst__n0574),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_12_12)
  );
  defparam DLX_IDinst_RegFile_20_12_3925.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_20_12_3925 (
    .I(DLX_IDinst_WB_data_eff[12]),
    .CE(DLX_IDinst__n0590),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_20_12)
  );
  defparam DLX_IDinst_RegFile_23_2_3926.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_23_2_3926 (
    .I(DLX_MEMinst_RF_data_in[2]),
    .CE(DLX_IDinst__n0596),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_23_2)
  );
  defparam DLX_IFinst_IR_curr_27.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_27 (
    .I(IR_MSB_3_OBUF),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[27])
  );
  defparam DLX_IDinst_RegFile_2_26_3927.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_2_26_3927 (
    .I(DLX_IDinst_WB_data_eff[26]),
    .CE(DLX_IDinst__n0554),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_2_26)
  );
  defparam DLX_IDinst_RegFile_10_20_3928.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_10_20_3928 (
    .I(\DLX_IDinst_RegFile_10_20/GROM ),
    .CE(DLX_IDinst__n0570),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_10_20)
  );
  defparam DLX_IDinst_RegFile_10_21_3929.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_10_21_3929 (
    .I(\DLX_IDinst_RegFile_10_21/GROM ),
    .CE(DLX_IDinst__n0570),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_10_21)
  );
  defparam DLX_IDinst_RegFile_10_22_3930.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_10_22_3930 (
    .I(\DLX_IDinst_RegFile_10_22/GROM ),
    .CE(DLX_IDinst__n0570),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_10_22)
  );
  defparam DLX_IDinst_RegFile_10_23_3931.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_10_23_3931 (
    .I(\DLX_IDinst_RegFile_10_23/GROM ),
    .CE(DLX_IDinst__n0570),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_10_23)
  );
  defparam DLX_IDinst_RegFile_10_31_3932.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_10_31_3932 (
    .I(\DLX_IDinst_RegFile_10_31/GROM ),
    .CE(DLX_IDinst__n0570),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_10_31)
  );
  defparam DLX_IDinst_RegFile_10_16_3933.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_10_16_3933 (
    .I(\DLX_IDinst_RegFile_10_16/GROM ),
    .CE(DLX_IDinst__n0570),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_10_16)
  );
  defparam DLX_IDinst_RegFile_10_24_3934.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_10_24_3934 (
    .I(\DLX_IDinst_RegFile_10_24/GROM ),
    .CE(DLX_IDinst__n0570),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_10_24)
  );
  defparam DLX_IDinst_RegFile_10_25_3935.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_10_25_3935 (
    .I(\DLX_IDinst_RegFile_10_25/GROM ),
    .CE(DLX_IDinst__n0570),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_10_25)
  );
  defparam DLX_IDinst_RegFile_10_17_3936.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_10_17_3936 (
    .I(\DLX_IDinst_RegFile_10_17/GROM ),
    .CE(DLX_IDinst__n0570),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_10_17)
  );
  defparam DLX_IDinst_RegFile_10_26_3937.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_10_26_3937 (
    .I(\DLX_IDinst_RegFile_10_26/GROM ),
    .CE(DLX_IDinst__n0570),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_10_26)
  );
  defparam DLX_IDinst_RegFile_10_18_3938.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_10_18_3938 (
    .I(\DLX_IDinst_RegFile_10_18/GROM ),
    .CE(DLX_IDinst__n0570),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_10_18)
  );
  defparam DLX_IDinst_RegFile_10_27_3939.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_10_27_3939 (
    .I(\DLX_IDinst_RegFile_10_27/GROM ),
    .CE(DLX_IDinst__n0570),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_10_27)
  );
  defparam DLX_IDinst_RegFile_10_19_3940.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_10_19_3940 (
    .I(\DLX_IDinst_RegFile_10_19/GROM ),
    .CE(DLX_IDinst__n0570),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_10_19)
  );
  defparam DLX_IDinst_RegFile_10_28_3941.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_10_28_3941 (
    .I(\DLX_IDinst_RegFile_10_28/GROM ),
    .CE(DLX_IDinst__n0570),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_10_28)
  );
  defparam DLX_IDinst_RegFile_10_29_3942.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_10_29_3942 (
    .I(\DLX_IDinst_RegFile_10_29/GROM ),
    .CE(DLX_IDinst__n0570),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_10_29)
  );
  defparam DLX_IDinst_Imm_10.INIT = 1'b0;
  X_SFF DLX_IDinst_Imm_10 (
    .I(DLX_IDinst__n0124),
    .CE(DLX_IDinst__n0116),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_IDinst__n0115),
    .O(\DLX_IDinst_Imm[10] )
  );
  defparam DLX_IDinst_IR_opcode_field_0.INIT = 1'b0;
  X_SFF DLX_IDinst_IR_opcode_field_0 (
    .I(DLX_IDinst__n0142[0]),
    .CE(DLX_IDinst__n0116),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_IDinst__n0115),
    .O(DLX_IDinst_IR_opcode_field[0])
  );
  defparam DLX_IDinst_IR_opcode_field_2.INIT = 1'b0;
  X_SFF DLX_IDinst_IR_opcode_field_2 (
    .I(DLX_IDinst__n0142[2]),
    .CE(DLX_IDinst__n0116),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_IDinst__n0115),
    .O(DLX_IDinst_IR_opcode_field[2])
  );
  defparam DLX_IDinst_Imm_9.INIT = 1'b0;
  X_SFF DLX_IDinst_Imm_9 (
    .I(DLX_IDinst__n0125),
    .CE(DLX_IDinst__n0116),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_IDinst__n0115),
    .O(\DLX_IDinst_Imm[9] )
  );
  defparam DLX_EXinst_ALU_result_10.INIT = 1'b0;
  X_SFF DLX_EXinst_ALU_result_10 (
    .I(\DLX_EXinst_ALU_result_10_1/GROM ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(N136886),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_ALU_result[10])
  );
  defparam DLX_IDinst_IR_opcode_field_5.INIT = 1'b0;
  X_SFF DLX_IDinst_IR_opcode_field_5 (
    .I(DLX_IDinst__n0142[5]),
    .CE(DLX_IDinst__n0116),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_IDinst__n0115),
    .O(DLX_IDinst_IR_opcode_field[5])
  );
  defparam DLX_IDinst_RegFile_3_26_3943.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_3_26_3943 (
    .I(DLX_IDinst_WB_data_eff[26]),
    .CE(DLX_IDinst__n0556),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_3_26)
  );
  defparam DLX_IFinst_IR_curr_19.INIT = 1'b0;
  X_SFF DLX_IFinst_IR_curr_19 (
    .I(IR[19]),
    .CE(DLX_IFinst_IR_curr_N3087),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_3),
    .O(DLX_IFinst_IR_curr[19])
  );
  defparam DLX_IDinst_counter_1.INIT = 1'b0;
  X_SFF DLX_IDinst_counter_1 (
    .I(DLX_IDinst__n0145[1]),
    .CE(DLX_IDinst__n0549),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_counter[1])
  );
  defparam DLX_IDinst_current_IR_5.INIT = 1'b0;
  X_SFF DLX_IDinst_current_IR_5 (
    .I(\DLX_IDinst_current_IR<5>/GROM ),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_current_IR[5])
  );
  defparam DLX_IDinst_current_IR_6.INIT = 1'b0;
  X_SFF DLX_IDinst_current_IR_6 (
    .I(\DLX_IDinst_current_IR<6>/GROM ),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_current_IR[6])
  );
  defparam DLX_IDinst_current_IR_7.INIT = 1'b0;
  X_SFF DLX_IDinst_current_IR_7 (
    .I(\DLX_IDinst_current_IR<7>/GROM ),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_current_IR[7])
  );
  defparam DLX_IDinst_current_IR_8.INIT = 1'b0;
  X_SFF DLX_IDinst_current_IR_8 (
    .I(\DLX_IDinst_current_IR<8>/GROM ),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_current_IR[8])
  );
  defparam DLX_IDinst_current_IR_9.INIT = 1'b0;
  X_SFF DLX_IDinst_current_IR_9 (
    .I(\DLX_IDinst_current_IR<9>/GROM ),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_current_IR[9])
  );
  defparam DLX_EXinst_reg_out_B_EX_9.INIT = 1'b0;
  X_SFF DLX_EXinst_reg_out_B_EX_9 (
    .I(DLX_EXinst__n0008[9]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_reg_out_B_EX[9])
  );
  defparam DLX_EXinst_reg_out_B_EX_10.INIT = 1'b0;
  X_SFF DLX_EXinst_reg_out_B_EX_10 (
    .I(DLX_EXinst__n0008[10]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_reg_out_B_EX[10])
  );
  defparam DLX_EXinst_reg_out_B_EX_8.INIT = 1'b0;
  X_SFF DLX_EXinst_reg_out_B_EX_8 (
    .I(DLX_EXinst__n0008[8]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_reg_out_B_EX[8])
  );
  defparam DLX_EXinst_ALU_result_8_1_3944.INIT = 1'b0;
  X_SFF DLX_EXinst_ALU_result_8_1_3944 (
    .I(\DLX_EXinst_ALU_result<8>/GROM ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(N136886),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_ALU_result_8_1)
  );
  defparam DLX_EXinst_ALU_result_8.INIT = 1'b0;
  X_SFF DLX_EXinst_ALU_result_8 (
    .I(N162844),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(N136886),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_ALU_result[8])
  );
  defparam DLX_EXinst_reg_out_B_EX_11.INIT = 1'b0;
  X_SFF DLX_EXinst_reg_out_B_EX_11 (
    .I(DLX_EXinst__n0008[11]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_reg_out_B_EX[11])
  );
  defparam DLX_EXinst_reg_out_B_EX_20.INIT = 1'b0;
  X_SFF DLX_EXinst_reg_out_B_EX_20 (
    .I(DLX_EXinst__n0008[20]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_reg_out_B_EX[20])
  );
  defparam DLX_EXinst_reg_out_B_EX_12.INIT = 1'b0;
  X_SFF DLX_EXinst_reg_out_B_EX_12 (
    .I(DLX_EXinst__n0008[12]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_reg_out_B_EX[12])
  );
  defparam DLX_IDinst_Imm_4.INIT = 1'b0;
  X_SFF DLX_IDinst_Imm_4 (
    .I(DLX_IDinst__n0143[4]),
    .CE(DLX_IDinst__n0116),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_IDinst__n0115),
    .O(\DLX_IDinst_Imm[4] )
  );
  defparam DLX_EXinst_ALU_result_11.INIT = 1'b0;
  X_SFF DLX_EXinst_ALU_result_11 (
    .I(\DLX_EXinst_ALU_result_11_1/GROM ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(N136886),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_ALU_result[11])
  );
  defparam DLX_EXinst_ALU_result_10_1_3945.INIT = 1'b0;
  X_SFF DLX_EXinst_ALU_result_10_1_3945 (
    .I(N162867),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(N136886),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_ALU_result_10_1)
  );
  defparam DLX_EXinst_ALU_result_12.INIT = 1'b0;
  X_SFF DLX_EXinst_ALU_result_12 (
    .I(\DLX_EXinst_ALU_result_12_1/GROM ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(N136886),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_ALU_result[12])
  );
  defparam DLX_EXinst_ALU_result_11_1_3946.INIT = 1'b0;
  X_SFF DLX_EXinst_ALU_result_11_1_3946 (
    .I(N162828),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(N136886),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_ALU_result_11_1)
  );
  defparam DLX_EXinst_ALU_result_13.INIT = 1'b0;
  X_SFF DLX_EXinst_ALU_result_13 (
    .I(\DLX_EXinst_ALU_result_13_1/GROM ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(N136886),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_ALU_result[13])
  );
  defparam DLX_EXinst_ALU_result_12_1_3947.INIT = 1'b0;
  X_SFF DLX_EXinst_ALU_result_12_1_3947 (
    .I(N162832),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(N136886),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_ALU_result_12_1)
  );
  defparam DLX_EXinst_ALU_result_14.INIT = 1'b0;
  X_SFF DLX_EXinst_ALU_result_14 (
    .I(\DLX_EXinst_ALU_result_14_1/GROM ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(N136886),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_ALU_result[14])
  );
  defparam DLX_EXinst_ALU_result_13_1_3948.INIT = 1'b0;
  X_SFF DLX_EXinst_ALU_result_13_1_3948 (
    .I(N162857),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(N136886),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_ALU_result_13_1)
  );
  defparam DLX_IDinst_current_IR_0.INIT = 1'b0;
  X_SFF DLX_IDinst_current_IR_0 (
    .I(\DLX_IDinst_current_IR<0>/GROM ),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_current_IR[0])
  );
  defparam DLX_EXinst_ALU_result_14_1_3949.INIT = 1'b0;
  X_SFF DLX_EXinst_ALU_result_14_1_3949 (
    .I(N162813),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(N136886),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_ALU_result_14_1)
  );
  defparam DLX_IDinst_current_IR_1.INIT = 1'b0;
  X_SFF DLX_IDinst_current_IR_1 (
    .I(\DLX_IDinst_current_IR<1>/GROM ),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_current_IR[1])
  );
  defparam DLX_IDinst_current_IR_2.INIT = 1'b0;
  X_SFF DLX_IDinst_current_IR_2 (
    .I(\DLX_IDinst_current_IR<2>/GROM ),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_current_IR[2])
  );
  defparam DLX_IDinst_current_IR_3.INIT = 1'b0;
  X_SFF DLX_IDinst_current_IR_3 (
    .I(\DLX_IDinst_current_IR<3>/GROM ),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_current_IR[3])
  );
  defparam DLX_IDinst_current_IR_4.INIT = 1'b0;
  X_SFF DLX_IDinst_current_IR_4 (
    .I(\DLX_IDinst_current_IR<4>/GROM ),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_current_IR[4])
  );
  defparam DLX_IDinst_reg_out_A_25.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_A_25 (
    .I(N162949),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE2798),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_A[25])
  );
  defparam DLX_IDinst_reg_out_B_10.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_B_10 (
    .I(DLX_IDinst__n0147[10]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_B[10])
  );
  defparam DLX_IDinst_reg_out_B_31.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_B_31 (
    .I(DLX_IDinst__n0147[31]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_B[31])
  );
  defparam DLX_IDinst_reg_out_A_26.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_A_26 (
    .I(N162952),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE2813),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_A[26])
  );
  defparam DLX_IDinst_reg_out_A_18.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_A_18 (
    .I(N162928),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE2708),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_A[18])
  );
  defparam DLX_IDinst_reg_out_B_11.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_B_11 (
    .I(DLX_IDinst__n0147[11]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_B[11])
  );
  defparam DLX_IDinst_reg_out_B_30.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_B_30 (
    .I(DLX_IDinst__n0147[30]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_B[30])
  );
  defparam DLX_IDinst_reg_out_A_27.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_A_27 (
    .I(N162955),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE2828),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_A[27])
  );
  defparam DLX_IDinst_reg_out_A_19.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_A_19 (
    .I(N162931),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE2693),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_A[19])
  );
  defparam DLX_IDinst_reg_out_B_20.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_B_20 (
    .I(DLX_IDinst__n0147[20]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_B[20])
  );
  defparam DLX_IDinst_reg_out_B_29.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_B_29 (
    .I(DLX_IDinst__n0147[29]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_B[29])
  );
  defparam DLX_IDinst_reg_out_B_21.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_B_21 (
    .I(DLX_IDinst__n0147[21]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_B[21])
  );
  defparam DLX_IDinst_reg_out_B_12.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_B_12 (
    .I(DLX_IDinst__n0147[12]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_B[12])
  );
  defparam DLX_IDinst_reg_out_B_27.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_B_27 (
    .I(DLX_IDinst__n0147[27]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_B[27])
  );
  defparam DLX_IDinst_reg_out_A_28.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_A_28 (
    .I(N162958),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE2843),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_A[28])
  );
  defparam DLX_IDinst_reg_out_B_13.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_B_13 (
    .I(DLX_IDinst__n0147[13]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_B[13])
  );
  defparam DLX_EXinst_reg_out_B_EX_13.INIT = 1'b0;
  X_SFF DLX_EXinst_reg_out_B_EX_13 (
    .I(DLX_EXinst__n0008[13]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_reg_out_B_EX[13])
  );
  defparam DLX_EXinst_reg_out_B_EX_16.INIT = 1'b0;
  X_SFF DLX_EXinst_reg_out_B_EX_16 (
    .I(DLX_EXinst__n0008[16]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_reg_out_B_EX[16])
  );
  defparam DLX_EXinst_reg_out_B_EX_17.INIT = 1'b0;
  X_SFF DLX_EXinst_reg_out_B_EX_17 (
    .I(DLX_EXinst__n0008[17]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_reg_out_B_EX[17])
  );
  defparam DLX_EXinst_reg_out_B_EX_21.INIT = 1'b0;
  X_SFF DLX_EXinst_reg_out_B_EX_21 (
    .I(DLX_EXinst__n0008[21]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_reg_out_B_EX[21])
  );
  defparam DLX_EXinst_reg_out_B_EX_14.INIT = 1'b0;
  X_SFF DLX_EXinst_reg_out_B_EX_14 (
    .I(DLX_EXinst__n0008[14]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_reg_out_B_EX[14])
  );
  defparam DLX_EXinst_reg_out_B_EX_22.INIT = 1'b0;
  X_SFF DLX_EXinst_reg_out_B_EX_22 (
    .I(DLX_EXinst__n0008[22]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_reg_out_B_EX[22])
  );
  defparam DLX_EXinst_reg_out_B_EX_19.INIT = 1'b0;
  X_SFF DLX_EXinst_reg_out_B_EX_19 (
    .I(DLX_EXinst__n0008[19]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_reg_out_B_EX[19])
  );
  defparam DLX_EXinst_reg_out_B_EX_24.INIT = 1'b0;
  X_SFF DLX_EXinst_reg_out_B_EX_24 (
    .I(DLX_EXinst__n0008[24]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_reg_out_B_EX[24])
  );
  defparam DLX_EXinst_reg_out_B_EX_23.INIT = 1'b0;
  X_SFF DLX_EXinst_reg_out_B_EX_23 (
    .I(DLX_EXinst__n0008[23]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_reg_out_B_EX[23])
  );
  defparam DLX_EXinst_reg_out_B_EX_27.INIT = 1'b0;
  X_SFF DLX_EXinst_reg_out_B_EX_27 (
    .I(DLX_EXinst__n0008[27]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_reg_out_B_EX[27])
  );
  defparam DLX_EXinst_reg_out_B_EX_25.INIT = 1'b0;
  X_SFF DLX_EXinst_reg_out_B_EX_25 (
    .I(DLX_EXinst__n0008[25]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_reg_out_B_EX[25])
  );
  defparam DLX_EXinst_reg_out_B_EX_28.INIT = 1'b0;
  X_SFF DLX_EXinst_reg_out_B_EX_28 (
    .I(DLX_EXinst__n0008[28]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_reg_out_B_EX[28])
  );
  defparam DLX_EXinst_reg_out_B_EX_29.INIT = 1'b0;
  X_SFF DLX_EXinst_reg_out_B_EX_29 (
    .I(DLX_EXinst__n0008[29]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_reg_out_B_EX[29])
  );
  defparam DLX_IDinst_intr_slot_3950.INIT = 1'b0;
  X_SFF DLX_IDinst_intr_slot_3950 (
    .I(DLX_IDinst__n0155),
    .CE(DLX_IDinst__n0616),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_intr_slot)
  );
  defparam DLX_IDinst_IR_function_field_5.INIT = 1'b0;
  X_SFF DLX_IDinst_IR_function_field_5 (
    .I(DLX_IDinst__n0143[5]),
    .CE(DLX_IDinst__n0116),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_IDinst__n0115),
    .O(DLX_IDinst_IR_function_field[5])
  );
  defparam DLX_IDinst_Imm_15.INIT = 1'b0;
  X_SFF DLX_IDinst_Imm_15 (
    .I(DLX_IDinst__n0119),
    .CE(DLX_IDinst__n0116),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_IDinst__n0115),
    .O(\DLX_IDinst_Imm[15] )
  );
  defparam DLX_MEMinst_RF_data_in_10.INIT = 1'b0;
  X_SFF DLX_MEMinst_RF_data_in_10 (
    .I(DLX_MEMinst__n0000[10]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_MEMinst_RF_data_in[10])
  );
  defparam DLX_MEMinst_RF_data_in_29.INIT = 1'b0;
  X_SFF DLX_MEMinst_RF_data_in_29 (
    .I(DLX_MEMinst__n0000[29]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_MEMinst_RF_data_in[29])
  );
  defparam DLX_MEMinst_RF_data_in_11.INIT = 1'b0;
  X_SFF DLX_MEMinst_RF_data_in_11 (
    .I(DLX_MEMinst__n0000[11]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_MEMinst_RF_data_in[11])
  );
  defparam DLX_MEMinst_RF_data_in_28.INIT = 1'b0;
  X_SFF DLX_MEMinst_RF_data_in_28 (
    .I(DLX_MEMinst__n0000[28]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_MEMinst_RF_data_in[28])
  );
  defparam DLX_MEMinst_RF_data_in_20.INIT = 1'b0;
  X_SFF DLX_MEMinst_RF_data_in_20 (
    .I(DLX_MEMinst__n0000[20]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_MEMinst_RF_data_in[20])
  );
  defparam DLX_MEMinst_RF_data_in_27.INIT = 1'b0;
  X_SFF DLX_MEMinst_RF_data_in_27 (
    .I(DLX_MEMinst__n0000[27]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_MEMinst_RF_data_in[27])
  );
  defparam DLX_MEMinst_RF_data_in_12.INIT = 1'b0;
  X_SFF DLX_MEMinst_RF_data_in_12 (
    .I(DLX_MEMinst__n0000[12]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_MEMinst_RF_data_in[12])
  );
  defparam DLX_MEMinst_RF_data_in_26.INIT = 1'b0;
  X_SFF DLX_MEMinst_RF_data_in_26 (
    .I(DLX_MEMinst__n0000[26]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_MEMinst_RF_data_in[26])
  );
  defparam DLX_MEMinst_RF_data_in_21.INIT = 1'b0;
  X_SFF DLX_MEMinst_RF_data_in_21 (
    .I(DLX_MEMinst__n0000[21]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_MEMinst_RF_data_in[21])
  );
  defparam DLX_IDinst_reg_out_B_2.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_B_2 (
    .I(DLX_IDinst__n0147[2]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_B[2])
  );
  defparam DLX_IDinst_reg_out_B_3.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_B_3 (
    .I(DLX_IDinst__n0147[3]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_B[3])
  );
  defparam DLX_IDinst_reg_out_A_11.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_A_11 (
    .I(N162907),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE2588),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_A[11])
  );
  defparam DLX_IDinst_reg_out_A_12.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_A_12 (
    .I(N162910),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE2603),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_A[12])
  );
  defparam DLX_IDinst_reg_out_A_20.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_A_20 (
    .I(N162934),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE2723),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_A[20])
  );
  defparam DLX_IDinst_reg_out_A_13.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_A_13 (
    .I(N162913),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE2618),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_A[13])
  );
  defparam DLX_IDinst_reg_out_A_21.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_A_21 (
    .I(N162937),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE2738),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_A[21])
  );
  defparam DLX_IDinst_reg_out_A_14.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_A_14 (
    .I(N162916),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE2633),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_A[14])
  );
  defparam DLX_IDinst_reg_out_A_22.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_A_22 (
    .I(N162940),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE2753),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_A[22])
  );
  defparam DLX_IDinst_reg_out_A_31.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_A_31 (
    .I(N162871),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE3232),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_A[31])
  );
  defparam DLX_IDinst_reg_out_A_15.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_A_15 (
    .I(N162919),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE2648),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_A[15])
  );
  defparam DLX_IDinst_reg_out_A_23.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_A_23 (
    .I(N162943),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE2768),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_A[23])
  );
  defparam DLX_IDinst_reg_out_A_16.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_A_16 (
    .I(N162922),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE2663),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_A[16])
  );
  defparam DLX_IDinst_reg_out_A_24.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_A_24 (
    .I(N162946),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE2783),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_A[24])
  );
  defparam DLX_IDinst_reg_out_A_17.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_A_17 (
    .I(N162925),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE2678),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_A[17])
  );
  defparam DLX_IDinst_Imm_8.INIT = 1'b0;
  X_SFF DLX_IDinst_Imm_8 (
    .I(DLX_IDinst__n0126),
    .CE(DLX_IDinst__n0116),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_IDinst__n0115),
    .O(\DLX_IDinst_Imm[8] )
  );
  defparam DLX_IDinst_Imm_7.INIT = 1'b0;
  X_SFF DLX_IDinst_Imm_7 (
    .I(DLX_IDinst__n0127),
    .CE(DLX_IDinst__n0116),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_IDinst__n0115),
    .O(\DLX_IDinst_Imm[7] )
  );
  defparam DLX_IDinst_rt_addr_2.INIT = 1'b0;
  X_SFF DLX_IDinst_rt_addr_2 (
    .I(DLX_IDinst__n0135[2]),
    .CE(DLX_IDinst__n0116),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_IDinst__n0115),
    .O(DLX_IDinst_rt_addr[2])
  );
  defparam DLX_IDinst_Imm_6.INIT = 1'b0;
  X_SFF DLX_IDinst_Imm_6 (
    .I(DLX_IDinst__n0128),
    .CE(DLX_IDinst__n0116),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_IDinst__n0115),
    .O(\DLX_IDinst_Imm[6] )
  );
  defparam DLX_IDinst_Imm_1_1_3951.INIT = 1'b0;
  X_SFF DLX_IDinst_Imm_1_1_3951 (
    .I(\DLX_IDinst_Imm<1>/GROM ),
    .CE(DLX_IDinst__n0116),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_IDinst__n0115),
    .O(DLX_IDinst_Imm_1_1)
  );
  defparam DLX_IDinst_rt_addr_3.INIT = 1'b0;
  X_SFF DLX_IDinst_rt_addr_3 (
    .I(DLX_IDinst__n0135[3]),
    .CE(DLX_IDinst__n0116),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_IDinst__n0115),
    .O(DLX_IDinst_rt_addr[3])
  );
  defparam DLX_IDinst_Imm_2_1_3952.INIT = 1'b0;
  X_SFF DLX_IDinst_Imm_2_1_3952 (
    .I(\DLX_IDinst_Imm<2>/GROM ),
    .CE(DLX_IDinst__n0116),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_IDinst__n0115),
    .O(DLX_IDinst_Imm_2_1)
  );
  defparam DLX_IDinst_Imm_1.INIT = 1'b0;
  X_SFF DLX_IDinst_Imm_1 (
    .I(DLX_IDinst__n0143[1]),
    .CE(DLX_IDinst__n0116),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_IDinst__n0115),
    .O(\DLX_IDinst_Imm[1] )
  );
  defparam DLX_IDinst_Imm_3_1_3953.INIT = 1'b0;
  X_SFF DLX_IDinst_Imm_3_1_3953 (
    .I(\DLX_IDinst_Imm<3>/GROM ),
    .CE(DLX_IDinst__n0116),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_IDinst__n0115),
    .O(DLX_IDinst_Imm_3_1)
  );
  defparam DLX_IDinst_Imm_2.INIT = 1'b0;
  X_SFF DLX_IDinst_Imm_2 (
    .I(DLX_IDinst__n0143[2]),
    .CE(DLX_IDinst__n0116),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_IDinst__n0115),
    .O(\DLX_IDinst_Imm[2] )
  );
  defparam DLX_IDinst_mem_read_3954.INIT = 1'b0;
  X_SFF DLX_IDinst_mem_read_3954 (
    .I(DLX_IDinst__n0140),
    .CE(DLX_IDinst__n0116),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_IDinst__n0115),
    .O(DLX_IDinst_mem_read)
  );
  defparam DLX_IDinst_Imm_3.INIT = 1'b0;
  X_SFF DLX_IDinst_Imm_3 (
    .I(DLX_IDinst__n0143[3]),
    .CE(DLX_IDinst__n0116),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_IDinst__n0115),
    .O(\DLX_IDinst_Imm[3] )
  );
  defparam DLX_IDinst_CLI_3955.INIT = 1'b0;
  X_SFF DLX_IDinst_CLI_3955 (
    .I(\DLX_IDinst_CLI/GROM ),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_CLI)
  );
  defparam DLX_IDinst_current_IR_10.INIT = 1'b0;
  X_SFF DLX_IDinst_current_IR_10 (
    .I(\DLX_IDinst_current_IR<10>/GROM ),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_current_IR[10])
  );
  defparam DLX_IDinst_current_IR_11.INIT = 1'b0;
  X_SFF DLX_IDinst_current_IR_11 (
    .I(\DLX_IDinst_current_IR<11>/GROM ),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_current_IR[11])
  );
  defparam DLX_IDinst_current_IR_20.INIT = 1'b0;
  X_SFF DLX_IDinst_current_IR_20 (
    .I(\DLX_IDinst_current_IR<20>/FROM ),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_current_IR[20])
  );
  defparam DLX_IDinst_current_IR_12.INIT = 1'b0;
  X_SFF DLX_IDinst_current_IR_12 (
    .I(\DLX_IDinst_current_IR<12>/GROM ),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_current_IR[12])
  );
  defparam DLX_IDinst_current_IR_13.INIT = 1'b0;
  X_SFF DLX_IDinst_current_IR_13 (
    .I(\DLX_IDinst_current_IR<13>/GROM ),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_current_IR[13])
  );
  defparam DLX_IDinst_current_IR_30.INIT = 1'b0;
  X_SFF DLX_IDinst_current_IR_30 (
    .I(\DLX_IDinst_current_IR<30>/FROM ),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_current_IR[30])
  );
  defparam DLX_IDinst_current_IR_22.INIT = 1'b0;
  X_SFF DLX_IDinst_current_IR_22 (
    .I(\DLX_IDinst_current_IR<22>/FROM ),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_current_IR[22])
  );
  defparam DLX_IDinst_current_IR_14.INIT = 1'b0;
  X_SFF DLX_IDinst_current_IR_14 (
    .I(\DLX_IDinst_current_IR<14>/GROM ),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_current_IR[14])
  );
  defparam DLX_IDinst_current_IR_23.INIT = 1'b0;
  X_SFF DLX_IDinst_current_IR_23 (
    .I(\DLX_IDinst_current_IR<23>/FROM ),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_current_IR[23])
  );
  defparam DLX_IDinst_current_IR_15.INIT = 1'b0;
  X_SFF DLX_IDinst_current_IR_15 (
    .I(\DLX_IDinst_current_IR<15>/GROM ),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_current_IR[15])
  );
  defparam DLX_IDinst_current_IR_31.INIT = 1'b0;
  X_SFF DLX_IDinst_current_IR_31 (
    .I(\DLX_IDinst_current_IR<31>/FROM ),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_current_IR[31])
  );
  defparam DLX_IDinst_current_IR_24.INIT = 1'b0;
  X_SFF DLX_IDinst_current_IR_24 (
    .I(\DLX_IDinst_current_IR<24>/FROM ),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_current_IR[24])
  );
  defparam DLX_IDinst_current_IR_25.INIT = 1'b0;
  X_SFF DLX_IDinst_current_IR_25 (
    .I(\DLX_IDinst_current_IR<25>/FROM ),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_current_IR[25])
  );
  defparam DLX_IDinst_current_IR_17.INIT = 1'b0;
  X_SFF DLX_IDinst_current_IR_17 (
    .I(\DLX_IDinst_current_IR<17>/FROM ),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_current_IR[17])
  );
  defparam DLX_IDinst_current_IR_26.INIT = 1'b0;
  X_SFF DLX_IDinst_current_IR_26 (
    .I(\DLX_IDinst_current_IR<26>/FROM ),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_current_IR[26])
  );
  defparam DLX_IDinst_current_IR_18.INIT = 1'b0;
  X_SFF DLX_IDinst_current_IR_18 (
    .I(\DLX_IDinst_current_IR<18>/FROM ),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_current_IR[18])
  );
  defparam DLX_IDinst_current_IR_27.INIT = 1'b0;
  X_SFF DLX_IDinst_current_IR_27 (
    .I(\DLX_IDinst_current_IR<27>/FROM ),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_current_IR[27])
  );
  defparam DLX_IDinst_current_IR_19.INIT = 1'b0;
  X_SFF DLX_IDinst_current_IR_19 (
    .I(\DLX_IDinst_current_IR<19>/FROM ),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_current_IR[19])
  );
  defparam DLX_IDinst_current_IR_28.INIT = 1'b0;
  X_SFF DLX_IDinst_current_IR_28 (
    .I(\DLX_IDinst_current_IR<28>/FROM ),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_current_IR[28])
  );
  defparam DLX_MEMinst_RF_data_in_0.INIT = 1'b0;
  X_SFF DLX_MEMinst_RF_data_in_0 (
    .I(DLX_MEMinst__n0000[0]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_MEMinst_RF_data_in[0])
  );
  defparam DLX_IDinst_current_IR_29.INIT = 1'b0;
  X_SFF DLX_IDinst_current_IR_29 (
    .I(\DLX_IDinst_current_IR<29>/FROM ),
    .CE(DLX_IDinst_N108233),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF),
    .O(DLX_IDinst_current_IR[29])
  );
  defparam DLX_MEMinst_RF_data_in_1.INIT = 1'b0;
  X_SFF DLX_MEMinst_RF_data_in_1 (
    .I(DLX_MEMinst__n0000[1]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_MEMinst_RF_data_in[1])
  );
  defparam DLX_MEMinst_RF_data_in_8.INIT = 1'b0;
  X_SFF DLX_MEMinst_RF_data_in_8 (
    .I(DLX_MEMinst__n0000[8]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_MEMinst_RF_data_in[8])
  );
  defparam DLX_MEMinst_RF_data_in_7.INIT = 1'b0;
  X_SFF DLX_MEMinst_RF_data_in_7 (
    .I(DLX_MEMinst__n0000[7]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_MEMinst_RF_data_in[7])
  );
  defparam DLX_MEMinst_RF_data_in_2.INIT = 1'b0;
  X_SFF DLX_MEMinst_RF_data_in_2 (
    .I(DLX_MEMinst__n0000[2]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_MEMinst_RF_data_in[2])
  );
  defparam DLX_MEMinst_RF_data_in_6.INIT = 1'b0;
  X_SFF DLX_MEMinst_RF_data_in_6 (
    .I(DLX_MEMinst__n0000[6]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_MEMinst_RF_data_in[6])
  );
  defparam DLX_MEMinst_RF_data_in_3.INIT = 1'b0;
  X_SFF DLX_MEMinst_RF_data_in_3 (
    .I(DLX_MEMinst__n0000[3]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_MEMinst_RF_data_in[3])
  );
  defparam DLX_MEMinst_RF_data_in_5.INIT = 1'b0;
  X_SFF DLX_MEMinst_RF_data_in_5 (
    .I(DLX_MEMinst__n0000[5]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_MEMinst_RF_data_in[5])
  );
  defparam DLX_IDinst_Imm_11.INIT = 1'b0;
  X_SFF DLX_IDinst_Imm_11 (
    .I(DLX_IDinst__n0123),
    .CE(DLX_IDinst__n0116),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_IDinst__n0115),
    .O(\DLX_IDinst_Imm[11] )
  );
  defparam DLX_MEMinst_RF_data_in_4.INIT = 1'b0;
  X_SFF DLX_MEMinst_RF_data_in_4 (
    .I(DLX_MEMinst__n0000[4]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_1),
    .O(DLX_MEMinst_RF_data_in[4])
  );
  defparam DLX_IDinst_Imm_14.INIT = 1'b0;
  X_SFF DLX_IDinst_Imm_14 (
    .I(DLX_IDinst__n0120),
    .CE(DLX_IDinst__n0116),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_IDinst__n0115),
    .O(\DLX_IDinst_Imm[14] )
  );
  defparam DLX_IDinst_Imm_12.INIT = 1'b0;
  X_SFF DLX_IDinst_Imm_12 (
    .I(DLX_IDinst__n0122),
    .CE(DLX_IDinst__n0116),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_IDinst__n0115),
    .O(\DLX_IDinst_Imm[12] )
  );
  defparam DLX_IDinst_reg_out_B_3_1_3956.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_B_3_1_3956 (
    .I(\DLX_IDinst_reg_out_B<3>/GROM ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_B_3_1)
  );
  defparam DLX_IDinst_Imm_13.INIT = 1'b0;
  X_SFF DLX_IDinst_Imm_13 (
    .I(DLX_IDinst__n0121),
    .CE(DLX_IDinst__n0116),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_IDinst__n0115),
    .O(\DLX_IDinst_Imm[13] )
  );
  defparam DLX_IDinst_reg_out_B_2_1_3957.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_B_2_1_3957 (
    .I(\DLX_IDinst_reg_out_B<2>/GROM ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_B_2_1)
  );
  defparam DLX_IDinst_RegFile_22_22_3958.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_22_22_3958 (
    .I(DLX_IDinst_WB_data_eff[22]),
    .CE(DLX_IDinst__n0594),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_22_22)
  );
  defparam DLX_IDinst_RegFile_30_30_3959.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_30_30_3959 (
    .I(DLX_IDinst_WB_data_eff[30]),
    .CE(DLX_IDinst__n0610),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_30_30)
  );
  defparam DLX_IDinst_RegFile_30_14_3960.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_30_14_3960 (
    .I(DLX_IDinst_WB_data_eff[14]),
    .CE(DLX_IDinst__n0610),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_30_14)
  );
  defparam DLX_IDinst_RegFile_14_15_3961.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_14_15_3961 (
    .I(DLX_IDinst_WB_data_eff[15]),
    .CE(DLX_IDinst__n0578),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_14_15)
  );
  defparam DLX_IDinst_RegFile_22_15_3962.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_22_15_3962 (
    .I(DLX_IDinst_WB_data_eff[15]),
    .CE(DLX_IDinst__n0594),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_22_15)
  );
  defparam DLX_IDinst_RegFile_30_15_3963.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_30_15_3963 (
    .I(DLX_IDinst_WB_data_eff[15]),
    .CE(DLX_IDinst__n0610),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_30_15)
  );
  defparam DLX_IDinst_RegFile_22_31_3964.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_22_31_3964 (
    .I(DLX_IDinst_WB_data_eff[31]),
    .CE(DLX_IDinst__n0594),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_22_31)
  );
  defparam DLX_IDinst_RegFile_14_24_3965.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_14_24_3965 (
    .I(DLX_IDinst_WB_data_eff[24]),
    .CE(DLX_IDinst__n0578),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_14_24)
  );
  defparam DLX_IDinst_RegFile_22_24_3966.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_22_24_3966 (
    .I(DLX_IDinst_WB_data_eff[24]),
    .CE(DLX_IDinst__n0594),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_22_24)
  );
  defparam DLX_IDinst_RegFile_30_24_3967.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_30_24_3967 (
    .I(DLX_IDinst_WB_data_eff[24]),
    .CE(DLX_IDinst__n0610),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_30_24)
  );
  defparam DLX_IDinst_RegFile_14_25_3968.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_14_25_3968 (
    .I(DLX_IDinst_WB_data_eff[25]),
    .CE(DLX_IDinst__n0578),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_14_25)
  );
  defparam DLX_IDinst_RegFile_22_25_3969.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_22_25_3969 (
    .I(DLX_IDinst_WB_data_eff[25]),
    .CE(DLX_IDinst__n0594),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_22_25)
  );
  defparam DLX_IDinst_RegFile_30_25_3970.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_30_25_3970 (
    .I(DLX_IDinst_WB_data_eff[25]),
    .CE(DLX_IDinst__n0610),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_30_25)
  );
  defparam DLX_IDinst_RegFile_14_26_3971.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_14_26_3971 (
    .I(DLX_IDinst_WB_data_eff[26]),
    .CE(DLX_IDinst__n0578),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_14_26)
  );
  defparam DLX_IDinst_RegFile_15_10_3972.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_15_10_3972 (
    .I(DLX_IDinst_WB_data_eff[10]),
    .CE(DLX_IDinst__n0580),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_15_10)
  );
  defparam DLX_IDinst_RegFile_22_18_3973.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_22_18_3973 (
    .I(DLX_IDinst_WB_data_eff[18]),
    .CE(DLX_IDinst__n0594),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_22_18)
  );
  defparam DLX_IDinst_RegFile_30_26_3974.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_30_26_3974 (
    .I(DLX_IDinst_WB_data_eff[26]),
    .CE(DLX_IDinst__n0610),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_30_26)
  );
  defparam DLX_IDinst_RegFile_31_10_3975.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_31_10_3975 (
    .I(DLX_IDinst_WB_data_eff[10]),
    .CE(DLX_IDinst__n0612),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_31_10)
  );
  defparam DLX_IDinst_RegFile_14_19_3976.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_14_19_3976 (
    .I(DLX_IDinst_WB_data_eff[19]),
    .CE(DLX_IDinst__n0578),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_14_19)
  );
  defparam DLX_IDinst_RegFile_22_27_3977.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_22_27_3977 (
    .I(DLX_IDinst_WB_data_eff[27]),
    .CE(DLX_IDinst__n0594),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_22_27)
  );
  defparam DLX_IDinst_RegFile_23_11_3978.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_23_11_3978 (
    .I(DLX_IDinst_WB_data_eff[11]),
    .CE(DLX_IDinst__n0596),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_23_11)
  );
  defparam DLX_IDinst_RegFile_14_28_3979.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_14_28_3979 (
    .I(DLX_IDinst_WB_data_eff[28]),
    .CE(DLX_IDinst__n0578),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_14_28)
  );
  defparam DLX_IDinst_RegFile_30_19_3980.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_30_19_3980 (
    .I(DLX_IDinst_WB_data_eff[19]),
    .CE(DLX_IDinst__n0610),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_30_19)
  );
  defparam DLX_IDinst_RegFile_11_29_3981.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_11_29_3981 (
    .I(DLX_IDinst_WB_data_eff[29]),
    .CE(DLX_IDinst__n0572),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_11_29)
  );
  defparam DLX_IDinst_RegFile_12_13_3982.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_12_13_3982 (
    .I(DLX_IDinst_WB_data_eff[13]),
    .CE(DLX_IDinst__n0574),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_12_13)
  );
  defparam DLX_IDinst_RegFile_12_21_3983.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_12_21_3983 (
    .I(DLX_IDinst_WB_data_eff[21]),
    .CE(DLX_IDinst__n0574),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_12_21)
  );
  defparam DLX_IDinst_RegFile_12_30_3984.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_12_30_3984 (
    .I(DLX_IDinst_WB_data_eff[30]),
    .CE(DLX_IDinst__n0574),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_12_30)
  );
  defparam DLX_IDinst_RegFile_20_21_3985.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_20_21_3985 (
    .I(DLX_IDinst_WB_data_eff[21]),
    .CE(DLX_IDinst__n0590),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_20_21)
  );
  defparam DLX_IDinst_RegFile_20_13_3986.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_20_13_3986 (
    .I(DLX_IDinst_WB_data_eff[13]),
    .CE(DLX_IDinst__n0590),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_20_13)
  );
  defparam DLX_IDinst_reg_out_A_3.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_A_3 (
    .I(N162883),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE2483),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_A[3])
  );
  defparam DLX_IDinst_reg_out_A_4.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_A_4 (
    .I(N162886),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE2498),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_A[4])
  );
  defparam DLX_IDinst_reg_out_B_1.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_B_1 (
    .I(DLX_IDinst__n0147[1]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_B[1])
  );
  defparam DLX_IDinst_reg_out_B_8.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_B_8 (
    .I(DLX_IDinst__n0147[8]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_B[8])
  );
  defparam DLX_IDinst_reg_out_A_6.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_A_6 (
    .I(N162892),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE3213),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_A[6])
  );
  defparam DLX_IDinst_reg_out_A_5.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_A_5 (
    .I(N162889),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE2513),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_A[5])
  );
  defparam DLX_IDinst_reg_out_A_7.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_A_7 (
    .I(N162895),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE2528),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_A[7])
  );
  defparam DLX_IDinst_reg_out_B_4.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_B_4 (
    .I(DLX_IDinst__n0147[4]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_B[4])
  );
  defparam DLX_IDinst_reg_out_B_7.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_B_7 (
    .I(DLX_IDinst__n0147[7]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_B[7])
  );
  defparam DLX_IDinst_reg_out_B_5.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_B_5 (
    .I(DLX_IDinst__n0147[5]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_B[5])
  );
  defparam DLX_IDinst_reg_out_A_8.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_A_8 (
    .I(N162898),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE2543),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_A[8])
  );
  defparam DLX_IDinst_reg_out_B_6.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_B_6 (
    .I(DLX_IDinst__n0147[6]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_B[6])
  );
  defparam DLX_EXinst_reg_dst_out_0.INIT = 1'b0;
  X_SFF DLX_EXinst_reg_dst_out_0 (
    .I(\DLX_EXinst_reg_dst_out<0>/GROM ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_reg_dst_out[0])
  );
  defparam DLX_IDinst_reg_out_A_9.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_A_9 (
    .I(N162901),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE2558),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_A[9])
  );
  defparam DLX_EXinst_reg_dst_out_1.INIT = 1'b0;
  X_SFF DLX_EXinst_reg_dst_out_1 (
    .I(\DLX_EXinst_reg_dst_out<1>/GROM ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_reg_dst_out[1])
  );
  defparam DLX_IDinst_reg_out_B_26.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_B_26 (
    .I(DLX_IDinst__n0147[26]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_B[26])
  );
  defparam DLX_IDinst_reg_out_B_22.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_B_22 (
    .I(DLX_IDinst__n0147[22]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_B[22])
  );
  defparam DLX_IDinst_reg_out_B_25.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_B_25 (
    .I(DLX_IDinst__n0147[25]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_B[25])
  );
  defparam DLX_IDinst_reg_out_A_29.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_A_29 (
    .I(N162961),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE2858),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_A[29])
  );
  defparam DLX_IDinst_reg_out_B_24.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_B_24 (
    .I(DLX_IDinst__n0147[24]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_B[24])
  );
  defparam DLX_IDinst_reg_out_B_14.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_B_14 (
    .I(DLX_IDinst__n0147[14]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_B[14])
  );
  defparam DLX_IDinst_reg_out_B_23.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_B_23 (
    .I(DLX_IDinst__n0147[23]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_B[23])
  );
  defparam DLX_IDinst_reg_out_B_15.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_B_15 (
    .I(DLX_IDinst__n0147[15]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_B[15])
  );
  defparam DLX_IDinst_reg_out_B_19.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_B_19 (
    .I(DLX_IDinst__n0147[19]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_B[19])
  );
  defparam DLX_IDinst_reg_out_B_16.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_B_16 (
    .I(DLX_IDinst__n0147[16]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_B[16])
  );
  defparam DLX_IDinst_reg_out_A_1.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_A_1 (
    .I(N162877),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE2903),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_A[1])
  );
  defparam DLX_IDinst_reg_out_B_18.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_B_18 (
    .I(DLX_IDinst__n0147[18]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_B[18])
  );
  defparam DLX_IDinst_reg_out_B_17.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_B_17 (
    .I(DLX_IDinst__n0147[17]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_B[17])
  );
  defparam DLX_IDinst_reg_out_A_2.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_A_2 (
    .I(N162880),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE2888),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_A[2])
  );
  defparam DLX_IDinst_reg_out_B_9.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_B_9 (
    .I(DLX_IDinst__n0147[9]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_B[9])
  );
  defparam DLX_IDinst_reg_out_A_0.INIT = 1'b0;
  X_SFF DLX_IDinst_reg_out_A_0 (
    .I(N162874),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(CHOICE3251),
    .SRST(reset_IBUF_14),
    .O(DLX_IDinst_reg_out_A[0])
  );
  defparam DLX_EXinst_reg_dst_out_2.INIT = 1'b0;
  X_SFF DLX_EXinst_reg_dst_out_2 (
    .I(\DLX_EXinst_reg_dst_out<2>/GROM ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_reg_dst_out[2])
  );
  defparam DLX_EXinst_reg_dst_out_3.INIT = 1'b0;
  X_SFF DLX_EXinst_reg_dst_out_3 (
    .I(\DLX_EXinst_reg_dst_out<3>/GROM ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_reg_dst_out[3])
  );
  defparam DLX_EXinst_reg_dst_out_4.INIT = 1'b0;
  X_SFF DLX_EXinst_reg_dst_out_4 (
    .I(\DLX_EXinst_reg_dst_out<4>/GROM ),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_reg_dst_out[4])
  );
  defparam DLX_EXinst_reg_out_B_EX_6.INIT = 1'b0;
  X_SFF DLX_EXinst_reg_out_B_EX_6 (
    .I(DLX_IDinst_reg_out_B[6]),
    .CE(VCC),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(DLX_EXinst__n0006),
    .O(DLX_EXinst_reg_out_B_EX[6])
  );
  defparam DLX_IDinst_RegFile_11_11_3987.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_11_11_3987 (
    .I(DLX_IDinst_WB_data_eff[11]),
    .CE(DLX_IDinst__n0572),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_11_11)
  );
  defparam DLX_IDinst_RegFile_11_12_3988.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_11_12_3988 (
    .I(DLX_IDinst_WB_data_eff[12]),
    .CE(DLX_IDinst__n0572),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_11_12)
  );
  defparam DLX_IDinst_RegFile_11_13_3989.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_11_13_3989 (
    .I(DLX_IDinst_WB_data_eff[13]),
    .CE(DLX_IDinst__n0572),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_11_13)
  );
  defparam DLX_IDinst_RegFile_11_22_3990.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_11_22_3990 (
    .I(DLX_IDinst_WB_data_eff[22]),
    .CE(DLX_IDinst__n0572),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_11_22)
  );
  defparam DLX_IDinst_RegFile_11_23_3991.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_11_23_3991 (
    .I(DLX_IDinst_WB_data_eff[23]),
    .CE(DLX_IDinst__n0572),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_11_23)
  );
  defparam DLX_IDinst_RegFile_11_31_3992.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_11_31_3992 (
    .I(DLX_IDinst_WB_data_eff[31]),
    .CE(DLX_IDinst__n0572),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_11_31)
  );
  defparam DLX_IDinst_RegFile_11_16_3993.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_11_16_3993 (
    .I(DLX_IDinst_WB_data_eff[16]),
    .CE(DLX_IDinst__n0572),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_11_16)
  );
  defparam DLX_IDinst_RegFile_11_17_3994.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_11_17_3994 (
    .I(DLX_IDinst_WB_data_eff[17]),
    .CE(DLX_IDinst__n0572),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_11_17)
  );
  defparam DLX_IDinst_RegFile_11_18_3995.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_11_18_3995 (
    .I(DLX_IDinst_WB_data_eff[18]),
    .CE(DLX_IDinst__n0572),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_13),
    .O(DLX_IDinst_RegFile_11_18)
  );
  defparam DLX_IDinst_RegFile_12_10_3996.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_12_10_3996 (
    .I(DLX_IDinst_WB_data_eff[10]),
    .CE(DLX_IDinst__n0574),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_12_10)
  );
  defparam DLX_IDinst_RegFile_20_10_3997.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_20_10_3997 (
    .I(DLX_IDinst_WB_data_eff[10]),
    .CE(DLX_IDinst__n0590),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_20_10)
  );
  defparam DLX_IDinst_RegFile_13_10_3998.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_13_10_3998 (
    .I(DLX_IDinst_WB_data_eff[10]),
    .CE(DLX_IDinst__n0576),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_13_10)
  );
  defparam DLX_IDinst_RegFile_20_26_3999.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_20_26_3999 (
    .I(DLX_IDinst_WB_data_eff[26]),
    .CE(DLX_IDinst__n0590),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_20_26)
  );
  defparam DLX_IDinst_RegFile_20_18_4000.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_20_18_4000 (
    .I(DLX_IDinst_WB_data_eff[18]),
    .CE(DLX_IDinst__n0590),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_20_18)
  );
  defparam DLX_IDinst_RegFile_12_27_4001.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_12_27_4001 (
    .I(DLX_IDinst_WB_data_eff[27]),
    .CE(DLX_IDinst__n0574),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_12_27)
  );
  defparam DLX_IDinst_RegFile_21_10_4002.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_21_10_4002 (
    .I(DLX_IDinst_WB_data_eff[10]),
    .CE(DLX_IDinst__n0592),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_21_10)
  );
  defparam DLX_IDinst_RegFile_12_22_4003.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_12_22_4003 (
    .I(DLX_IDinst_WB_data_eff[22]),
    .CE(DLX_IDinst__n0574),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_12_22)
  );
  defparam DLX_IDinst_RegFile_12_14_4004.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_12_14_4004 (
    .I(DLX_IDinst_WB_data_eff[14]),
    .CE(DLX_IDinst__n0574),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_12_14)
  );
  defparam DLX_IDinst_RegFile_20_30_4005.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_20_30_4005 (
    .I(DLX_IDinst_WB_data_eff[30]),
    .CE(DLX_IDinst__n0590),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_20_30)
  );
  defparam DLX_IDinst_RegFile_20_14_4006.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_20_14_4006 (
    .I(DLX_IDinst_WB_data_eff[14]),
    .CE(DLX_IDinst__n0590),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_20_14)
  );
  defparam DLX_IDinst_RegFile_20_22_4007.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_20_22_4007 (
    .I(DLX_IDinst_WB_data_eff[22]),
    .CE(DLX_IDinst__n0590),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_20_22)
  );
  defparam DLX_IDinst_RegFile_20_31_4008.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_20_31_4008 (
    .I(DLX_IDinst_WB_data_eff[31]),
    .CE(DLX_IDinst__n0590),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_20_31)
  );
  defparam DLX_IDinst_RegFile_12_24_4009.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_12_24_4009 (
    .I(DLX_IDinst_WB_data_eff[24]),
    .CE(DLX_IDinst__n0574),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_12_24)
  );
  defparam DLX_IDinst_RegFile_12_16_4010.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_12_16_4010 (
    .I(DLX_IDinst_WB_data_eff[16]),
    .CE(DLX_IDinst__n0574),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_12_16)
  );
  defparam DLX_IDinst_RegFile_20_16_4011.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_20_16_4011 (
    .I(DLX_IDinst_WB_data_eff[16]),
    .CE(DLX_IDinst__n0590),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_20_16)
  );
  defparam DLX_IDinst_RegFile_20_24_4012.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_20_24_4012 (
    .I(DLX_IDinst_WB_data_eff[24]),
    .CE(DLX_IDinst__n0590),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_20_24)
  );
  defparam DLX_IDinst_RegFile_12_23_4013.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_12_23_4013 (
    .I(DLX_IDinst_WB_data_eff[23]),
    .CE(DLX_IDinst__n0574),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_12_23)
  );
  defparam DLX_IDinst_RegFile_12_15_4014.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_12_15_4014 (
    .I(DLX_IDinst_WB_data_eff[15]),
    .CE(DLX_IDinst__n0574),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_12_15)
  );
  defparam DLX_IDinst_RegFile_20_23_4015.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_20_23_4015 (
    .I(DLX_IDinst_WB_data_eff[23]),
    .CE(DLX_IDinst__n0590),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_20_23)
  );
  defparam DLX_IDinst_RegFile_12_31_4016.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_12_31_4016 (
    .I(DLX_IDinst_WB_data_eff[31]),
    .CE(DLX_IDinst__n0574),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_12_31)
  );
  defparam DLX_IDinst_RegFile_20_15_4017.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_20_15_4017 (
    .I(DLX_IDinst_WB_data_eff[15]),
    .CE(DLX_IDinst__n0590),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_20_15)
  );
  defparam DLX_IDinst_RegFile_12_25_4018.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_12_25_4018 (
    .I(DLX_IDinst_WB_data_eff[25]),
    .CE(DLX_IDinst__n0574),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_12_25)
  );
  defparam DLX_IDinst_RegFile_12_17_4019.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_12_17_4019 (
    .I(DLX_IDinst_WB_data_eff[17]),
    .CE(DLX_IDinst__n0574),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_12_17)
  );
  defparam DLX_IDinst_RegFile_20_25_4020.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_20_25_4020 (
    .I(DLX_IDinst_WB_data_eff[25]),
    .CE(DLX_IDinst__n0590),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_20_25)
  );
  defparam DLX_IDinst_RegFile_12_18_4021.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_12_18_4021 (
    .I(DLX_IDinst_WB_data_eff[18]),
    .CE(DLX_IDinst__n0574),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_12_18)
  );
  defparam DLX_IDinst_RegFile_20_17_4022.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_20_17_4022 (
    .I(DLX_IDinst_WB_data_eff[17]),
    .CE(DLX_IDinst__n0590),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_20_17)
  );
  defparam DLX_IDinst_RegFile_12_26_4023.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_12_26_4023 (
    .I(DLX_IDinst_WB_data_eff[26]),
    .CE(DLX_IDinst__n0574),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_12_26)
  );
  defparam DLX_IDinst_RegFile_12_28_4024.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_12_28_4024 (
    .I(DLX_IDinst_WB_data_eff[28]),
    .CE(DLX_IDinst__n0574),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_12_28)
  );
  defparam DLX_IDinst_RegFile_13_20_4025.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_13_20_4025 (
    .I(DLX_IDinst_WB_data_eff[20]),
    .CE(DLX_IDinst__n0576),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_13_20)
  );
  defparam DLX_IDinst_RegFile_13_12_4026.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_13_12_4026 (
    .I(DLX_IDinst_WB_data_eff[12]),
    .CE(DLX_IDinst__n0576),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_13_12)
  );
  defparam DLX_IDinst_RegFile_21_12_4027.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_21_12_4027 (
    .I(DLX_IDinst_WB_data_eff[12]),
    .CE(DLX_IDinst__n0592),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_21_12)
  );
  defparam DLX_IDinst_RegFile_20_28_4028.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_20_28_4028 (
    .I(DLX_IDinst_WB_data_eff[28]),
    .CE(DLX_IDinst__n0590),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_20_28)
  );
  defparam DLX_IDinst_RegFile_21_20_4029.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_21_20_4029 (
    .I(DLX_IDinst_WB_data_eff[20]),
    .CE(DLX_IDinst__n0592),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_21_20)
  );
  defparam DLX_IDinst_RegFile_12_19_4030.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_12_19_4030 (
    .I(DLX_IDinst_WB_data_eff[19]),
    .CE(DLX_IDinst__n0574),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_12_19)
  );
  defparam DLX_IDinst_RegFile_13_11_4031.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_13_11_4031 (
    .I(DLX_IDinst_WB_data_eff[11]),
    .CE(DLX_IDinst__n0576),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_13_11)
  );
  defparam DLX_IDinst_RegFile_20_27_4032.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_20_27_4032 (
    .I(DLX_IDinst_WB_data_eff[27]),
    .CE(DLX_IDinst__n0590),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_20_27)
  );
  defparam DLX_IDinst_RegFile_21_11_4033.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_21_11_4033 (
    .I(DLX_IDinst_WB_data_eff[11]),
    .CE(DLX_IDinst__n0592),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_21_11)
  );
  defparam DLX_IDinst_RegFile_20_19_4034.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_20_19_4034 (
    .I(DLX_IDinst_WB_data_eff[19]),
    .CE(DLX_IDinst__n0590),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_20_19)
  );
  defparam DLX_IDinst_RegFile_12_29_4035.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_12_29_4035 (
    .I(DLX_IDinst_WB_data_eff[29]),
    .CE(DLX_IDinst__n0574),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_12_29)
  );
  defparam DLX_IDinst_RegFile_13_21_4036.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_13_21_4036 (
    .I(DLX_IDinst_WB_data_eff[21]),
    .CE(DLX_IDinst__n0576),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_13_21)
  );
  defparam DLX_IDinst_RegFile_13_13_4037.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_13_13_4037 (
    .I(DLX_IDinst_WB_data_eff[13]),
    .CE(DLX_IDinst__n0576),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_13_13)
  );
  defparam DLX_IDinst_RegFile_21_21_4038.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_21_21_4038 (
    .I(DLX_IDinst_WB_data_eff[21]),
    .CE(DLX_IDinst__n0592),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_21_21)
  );
  defparam DLX_IDinst_RegFile_20_29_4039.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_20_29_4039 (
    .I(DLX_IDinst_WB_data_eff[29]),
    .CE(DLX_IDinst__n0590),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_20_29)
  );
  defparam DLX_IDinst_RegFile_21_13_4040.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_21_13_4040 (
    .I(DLX_IDinst_WB_data_eff[13]),
    .CE(DLX_IDinst__n0592),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_21_13)
  );
  defparam DLX_IDinst_RegFile_13_30_4041.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_13_30_4041 (
    .I(DLX_IDinst_WB_data_eff[30]),
    .CE(DLX_IDinst__n0576),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_13_30)
  );
  defparam DLX_IDinst_RegFile_13_22_4042.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_13_22_4042 (
    .I(DLX_IDinst_WB_data_eff[22]),
    .CE(DLX_IDinst__n0576),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_13_22)
  );
  defparam DLX_IDinst_RegFile_21_30_4043.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_21_30_4043 (
    .I(DLX_IDinst_WB_data_eff[30]),
    .CE(DLX_IDinst__n0592),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_21_30)
  );
  defparam DLX_IDinst_RegFile_13_14_4044.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_13_14_4044 (
    .I(DLX_IDinst_WB_data_eff[14]),
    .CE(DLX_IDinst__n0576),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_13_14)
  );
  defparam DLX_IDinst_RegFile_13_31_4045.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_13_31_4045 (
    .I(DLX_IDinst_WB_data_eff[31]),
    .CE(DLX_IDinst__n0576),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_13_31)
  );
  defparam DLX_IDinst_RegFile_21_31_4046.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_21_31_4046 (
    .I(DLX_IDinst_WB_data_eff[31]),
    .CE(DLX_IDinst__n0592),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_21_31)
  );
  defparam DLX_IDinst_RegFile_13_24_4047.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_13_24_4047 (
    .I(DLX_IDinst_WB_data_eff[24]),
    .CE(DLX_IDinst__n0576),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_13_24)
  );
  defparam DLX_IDinst_RegFile_21_24_4048.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_21_24_4048 (
    .I(DLX_IDinst_WB_data_eff[24]),
    .CE(DLX_IDinst__n0592),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_21_24)
  );
  defparam DLX_IDinst_RegFile_13_16_4049.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_13_16_4049 (
    .I(DLX_IDinst_WB_data_eff[16]),
    .CE(DLX_IDinst__n0576),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_13_16)
  );
  defparam DLX_IDinst_RegFile_21_22_4050.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_21_22_4050 (
    .I(DLX_IDinst_WB_data_eff[22]),
    .CE(DLX_IDinst__n0592),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_21_22)
  );
  defparam DLX_IDinst_RegFile_21_14_4051.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_21_14_4051 (
    .I(DLX_IDinst_WB_data_eff[14]),
    .CE(DLX_IDinst__n0592),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_21_14)
  );
  defparam DLX_IDinst_RegFile_13_23_4052.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_13_23_4052 (
    .I(DLX_IDinst_WB_data_eff[23]),
    .CE(DLX_IDinst__n0576),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_13_23)
  );
  defparam DLX_IDinst_RegFile_21_23_4053.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_21_23_4053 (
    .I(DLX_IDinst_WB_data_eff[23]),
    .CE(DLX_IDinst__n0592),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_21_23)
  );
  defparam DLX_IDinst_RegFile_13_15_4054.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_13_15_4054 (
    .I(DLX_IDinst_WB_data_eff[15]),
    .CE(DLX_IDinst__n0576),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_13_15)
  );
  defparam DLX_IDinst_RegFile_21_15_4055.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_21_15_4055 (
    .I(DLX_IDinst_WB_data_eff[15]),
    .CE(DLX_IDinst__n0592),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_21_15)
  );
  defparam DLX_IDinst_RegFile_13_26_4056.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_13_26_4056 (
    .I(DLX_IDinst_WB_data_eff[26]),
    .CE(DLX_IDinst__n0576),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_13_26)
  );
  defparam DLX_IDinst_RegFile_13_18_4057.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_13_18_4057 (
    .I(DLX_IDinst_WB_data_eff[18]),
    .CE(DLX_IDinst__n0576),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_13_18)
  );
  defparam DLX_IDinst_RegFile_21_18_4058.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_21_18_4058 (
    .I(DLX_IDinst_WB_data_eff[18]),
    .CE(DLX_IDinst__n0592),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_21_18)
  );
  defparam DLX_IDinst_RegFile_21_26_4059.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_21_26_4059 (
    .I(DLX_IDinst_WB_data_eff[26]),
    .CE(DLX_IDinst__n0592),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_21_26)
  );
  defparam DLX_IDinst_RegFile_13_27_4060.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_13_27_4060 (
    .I(DLX_IDinst_WB_data_eff[27]),
    .CE(DLX_IDinst__n0576),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_13_27)
  );
  defparam DLX_IDinst_RegFile_22_10_4061.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_22_10_4061 (
    .I(DLX_IDinst_WB_data_eff[10]),
    .CE(DLX_IDinst__n0594),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_22_10)
  );
  defparam DLX_IDinst_RegFile_21_16_4062.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_21_16_4062 (
    .I(DLX_IDinst_WB_data_eff[16]),
    .CE(DLX_IDinst__n0592),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_21_16)
  );
  defparam DLX_IDinst_RegFile_13_25_4063.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_13_25_4063 (
    .I(DLX_IDinst_WB_data_eff[25]),
    .CE(DLX_IDinst__n0576),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_13_25)
  );
  defparam DLX_IDinst_RegFile_13_17_4064.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_13_17_4064 (
    .I(DLX_IDinst_WB_data_eff[17]),
    .CE(DLX_IDinst__n0576),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_13_17)
  );
  defparam DLX_IDinst_RegFile_21_17_4065.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_21_17_4065 (
    .I(DLX_IDinst_WB_data_eff[17]),
    .CE(DLX_IDinst__n0592),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_21_17)
  );
  defparam DLX_IDinst_RegFile_21_25_4066.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_21_25_4066 (
    .I(DLX_IDinst_WB_data_eff[25]),
    .CE(DLX_IDinst__n0592),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_21_25)
  );
  defparam DLX_IDinst_RegFile_14_13_4067.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_14_13_4067 (
    .I(DLX_IDinst_WB_data_eff[13]),
    .CE(DLX_IDinst__n0578),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_14_13)
  );
  defparam DLX_IDinst_RegFile_22_12_4068.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_22_12_4068 (
    .I(DLX_IDinst_WB_data_eff[12]),
    .CE(DLX_IDinst__n0594),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_22_12)
  );
  defparam DLX_IDinst_RegFile_13_29_4069.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_13_29_4069 (
    .I(DLX_IDinst_WB_data_eff[29]),
    .CE(DLX_IDinst__n0576),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_13_29)
  );
  defparam DLX_IDinst_RegFile_30_12_4070.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_30_12_4070 (
    .I(DLX_IDinst_WB_data_eff[12]),
    .CE(DLX_IDinst__n0610),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_30_12)
  );
  defparam DLX_IDinst_RegFile_22_21_4071.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_22_21_4071 (
    .I(DLX_IDinst_WB_data_eff[21]),
    .CE(DLX_IDinst__n0594),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_22_21)
  );
  defparam DLX_IDinst_RegFile_14_14_4072.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_14_14_4072 (
    .I(DLX_IDinst_WB_data_eff[14]),
    .CE(DLX_IDinst__n0578),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_14_14)
  );
  defparam DLX_IDinst_RegFile_21_29_4073.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_21_29_4073 (
    .I(DLX_IDinst_WB_data_eff[29]),
    .CE(DLX_IDinst__n0592),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_21_29)
  );
  defparam DLX_IDinst_RegFile_14_30_4074.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_14_30_4074 (
    .I(DLX_IDinst_WB_data_eff[30]),
    .CE(DLX_IDinst__n0578),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_14_30)
  );
  defparam DLX_IDinst_RegFile_30_21_4075.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_30_21_4075 (
    .I(DLX_IDinst_WB_data_eff[21]),
    .CE(DLX_IDinst__n0610),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_30_21)
  );
  defparam DLX_IDinst_RegFile_13_19_4076.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_13_19_4076 (
    .I(DLX_IDinst_WB_data_eff[19]),
    .CE(DLX_IDinst__n0576),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_13_19)
  );
  defparam DLX_IDinst_RegFile_14_11_4077.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_14_11_4077 (
    .I(DLX_IDinst_WB_data_eff[11]),
    .CE(DLX_IDinst__n0578),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_14_11)
  );
  defparam DLX_IDinst_RegFile_21_19_4078.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_21_19_4078 (
    .I(DLX_IDinst_WB_data_eff[19]),
    .CE(DLX_IDinst__n0592),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_21_19)
  );
  defparam DLX_IDinst_RegFile_21_27_4079.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_21_27_4079 (
    .I(DLX_IDinst_WB_data_eff[27]),
    .CE(DLX_IDinst__n0592),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_21_27)
  );
  defparam DLX_IDinst_RegFile_21_28_4080.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_21_28_4080 (
    .I(DLX_IDinst_WB_data_eff[28]),
    .CE(DLX_IDinst__n0592),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_21_28)
  );
  defparam DLX_IDinst_RegFile_30_11_4081.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_30_11_4081 (
    .I(DLX_IDinst_WB_data_eff[11]),
    .CE(DLX_IDinst__n0610),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_30_11)
  );
  defparam DLX_IDinst_RegFile_14_20_4082.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_14_20_4082 (
    .I(DLX_IDinst_WB_data_eff[20]),
    .CE(DLX_IDinst__n0578),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_14_20)
  );
  defparam DLX_IDinst_RegFile_13_28_4083.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_13_28_4083 (
    .I(DLX_IDinst_WB_data_eff[28]),
    .CE(DLX_IDinst__n0576),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_12),
    .O(DLX_IDinst_RegFile_13_28)
  );
  defparam DLX_IDinst_RegFile_15_12_4084.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_15_12_4084 (
    .I(DLX_IDinst_WB_data_eff[12]),
    .CE(DLX_IDinst__n0580),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_15_12)
  );
  defparam DLX_IDinst_RegFile_23_20_4085.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_23_20_4085 (
    .I(DLX_IDinst_WB_data_eff[20]),
    .CE(DLX_IDinst__n0596),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_23_20)
  );
  defparam DLX_IDinst_RegFile_30_28_4086.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_30_28_4086 (
    .I(DLX_IDinst_WB_data_eff[28]),
    .CE(DLX_IDinst__n0610),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_30_28)
  );
  defparam DLX_IDinst_RegFile_31_12_4087.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_31_12_4087 (
    .I(DLX_IDinst_WB_data_eff[12]),
    .CE(DLX_IDinst__n0612),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_31_12)
  );
  defparam DLX_IDinst_RegFile_15_21_4088.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_15_21_4088 (
    .I(DLX_IDinst_WB_data_eff[21]),
    .CE(DLX_IDinst__n0580),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_15_21)
  );
  defparam DLX_IDinst_RegFile_22_29_4089.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_22_29_4089 (
    .I(DLX_IDinst_WB_data_eff[29]),
    .CE(DLX_IDinst__n0594),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_9),
    .O(DLX_IDinst_RegFile_22_29)
  );
  defparam DLX_IDinst_RegFile_23_13_4090.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_23_13_4090 (
    .I(DLX_IDinst_WB_data_eff[13]),
    .CE(DLX_IDinst__n0596),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_23_13)
  );
  defparam DLX_IDinst_RegFile_31_21_4091.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_31_21_4091 (
    .I(DLX_IDinst_WB_data_eff[21]),
    .CE(DLX_IDinst__n0612),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_31_21)
  );
  defparam DLX_IDinst_RegFile_15_30_4092.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_15_30_4092 (
    .I(DLX_IDinst_WB_data_eff[30]),
    .CE(DLX_IDinst__n0580),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_15_30)
  );
  defparam DLX_IDinst_RegFile_15_14_4093.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_15_14_4093 (
    .I(DLX_IDinst_WB_data_eff[14]),
    .CE(DLX_IDinst__n0580),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_15_14)
  );
  defparam DLX_IDinst_RegFile_23_22_4094.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_23_22_4094 (
    .I(DLX_IDinst_WB_data_eff[22]),
    .CE(DLX_IDinst__n0596),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_23_22)
  );
  defparam DLX_IDinst_RegFile_31_30_4095.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_31_30_4095 (
    .I(DLX_IDinst_WB_data_eff[30]),
    .CE(DLX_IDinst__n0612),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_31_30)
  );
  defparam DLX_IDinst_RegFile_31_14_4096.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_31_14_4096 (
    .I(DLX_IDinst_WB_data_eff[14]),
    .CE(DLX_IDinst__n0612),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_31_14)
  );
  defparam DLX_IDinst_RegFile_15_15_4097.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_15_15_4097 (
    .I(DLX_IDinst_WB_data_eff[15]),
    .CE(DLX_IDinst__n0580),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_15_15)
  );
  defparam DLX_IDinst_RegFile_23_15_4098.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_23_15_4098 (
    .I(DLX_IDinst_WB_data_eff[15]),
    .CE(DLX_IDinst__n0596),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_23_15)
  );
  defparam DLX_IDinst_RegFile_31_15_4099.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_31_15_4099 (
    .I(DLX_IDinst_WB_data_eff[15]),
    .CE(DLX_IDinst__n0612),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_6),
    .O(DLX_IDinst_RegFile_31_15)
  );
  defparam DLX_IDinst_RegFile_23_31_4100.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_23_31_4100 (
    .I(DLX_IDinst_WB_data_eff[31]),
    .CE(DLX_IDinst__n0596),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_23_31)
  );
  defparam DLX_IDinst_RegFile_15_24_4101.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_15_24_4101 (
    .I(DLX_IDinst_WB_data_eff[24]),
    .CE(DLX_IDinst__n0580),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_15_24)
  );
  defparam DLX_IDinst_RegFile_23_24_4102.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_23_24_4102 (
    .I(DLX_IDinst_WB_data_eff[24]),
    .CE(DLX_IDinst__n0596),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_23_24)
  );
  defparam DLX_IDinst_RegFile_31_24_4103.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_31_24_4103 (
    .I(DLX_IDinst_WB_data_eff[24]),
    .CE(DLX_IDinst__n0612),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_31_24)
  );
  defparam DLX_IDinst_RegFile_15_25_4104.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_15_25_4104 (
    .I(DLX_IDinst_WB_data_eff[25]),
    .CE(DLX_IDinst__n0580),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_15_25)
  );
  defparam DLX_IDinst_RegFile_23_25_4105.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_23_25_4105 (
    .I(DLX_IDinst_WB_data_eff[25]),
    .CE(DLX_IDinst__n0596),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_23_25)
  );
  defparam DLX_IDinst_RegFile_31_25_4106.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_31_25_4106 (
    .I(DLX_IDinst_WB_data_eff[25]),
    .CE(DLX_IDinst__n0612),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_31_25)
  );
  defparam DLX_IDinst_RegFile_15_26_4107.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_15_26_4107 (
    .I(DLX_IDinst_WB_data_eff[26]),
    .CE(DLX_IDinst__n0580),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_15_26)
  );
  defparam DLX_IDinst_RegFile_16_10_4108.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_16_10_4108 (
    .I(DLX_IDinst_WB_data_eff[10]),
    .CE(DLX_IDinst__n0582),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_16_10)
  );
  defparam DLX_IDinst_RegFile_23_18_4109.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_23_18_4109 (
    .I(DLX_IDinst_WB_data_eff[18]),
    .CE(DLX_IDinst__n0596),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_23_18)
  );
  defparam DLX_IDinst_RegFile_31_26_4110.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_31_26_4110 (
    .I(DLX_IDinst_WB_data_eff[26]),
    .CE(DLX_IDinst__n0612),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_31_26)
  );
  defparam DLX_IDinst_RegFile_23_19_4111.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_23_19_4111 (
    .I(DLX_IDinst_WB_data_eff[19]),
    .CE(DLX_IDinst__n0596),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_23_19)
  );
  defparam DLX_IDinst_RegFile_24_10_4112.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_24_10_4112 (
    .I(DLX_IDinst_WB_data_eff[10]),
    .CE(DLX_IDinst__n0598),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_24_10)
  );
  defparam DLX_IDinst_RegFile_16_11_4113.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_16_11_4113 (
    .I(DLX_IDinst_WB_data_eff[11]),
    .CE(DLX_IDinst__n0582),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_16_11)
  );
  defparam DLX_IDinst_RegFile_15_27_4114.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_15_27_4114 (
    .I(DLX_IDinst_WB_data_eff[27]),
    .CE(DLX_IDinst__n0580),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_15_27)
  );
  defparam DLX_IDinst_RegFile_15_28_4115.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_15_28_4115 (
    .I(DLX_IDinst_WB_data_eff[28]),
    .CE(DLX_IDinst__n0580),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_15_28)
  );
  defparam DLX_IDinst_RegFile_31_27_4116.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_31_27_4116 (
    .I(DLX_IDinst_WB_data_eff[27]),
    .CE(DLX_IDinst__n0612),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_31_27)
  );
  defparam DLX_IDinst_RegFile_24_11_4117.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_24_11_4117 (
    .I(DLX_IDinst_WB_data_eff[11]),
    .CE(DLX_IDinst__n0598),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_24_11)
  );
  defparam DLX_IDinst_RegFile_16_12_4118.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_16_12_4118 (
    .I(DLX_IDinst_WB_data_eff[12]),
    .CE(DLX_IDinst__n0582),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_16_12)
  );
  defparam DLX_IDinst_RegFile_16_20_4119.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_16_20_4119 (
    .I(DLX_IDinst_WB_data_eff[20]),
    .CE(DLX_IDinst__n0582),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_16_20)
  );
  defparam DLX_IDinst_RegFile_15_29_4120.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_15_29_4120 (
    .I(DLX_IDinst_WB_data_eff[29]),
    .CE(DLX_IDinst__n0580),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_15_29)
  );
  defparam DLX_IDinst_RegFile_23_28_4121.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_23_28_4121 (
    .I(DLX_IDinst_WB_data_eff[28]),
    .CE(DLX_IDinst__n0596),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_23_28)
  );
  defparam DLX_IDinst_RegFile_31_28_4122.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_31_28_4122 (
    .I(DLX_IDinst_WB_data_eff[28]),
    .CE(DLX_IDinst__n0612),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_5),
    .O(DLX_IDinst_RegFile_31_28)
  );
  defparam DLX_IDinst_RegFile_24_20_4123.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_24_20_4123 (
    .I(DLX_IDinst_WB_data_eff[20]),
    .CE(DLX_IDinst__n0598),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_24_20)
  );
  defparam DLX_IDinst_RegFile_16_21_4124.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_16_21_4124 (
    .I(DLX_IDinst_WB_data_eff[21]),
    .CE(DLX_IDinst__n0582),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_16_21)
  );
  defparam DLX_IDinst_RegFile_23_29_4125.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_23_29_4125 (
    .I(DLX_IDinst_WB_data_eff[29]),
    .CE(DLX_IDinst__n0596),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_23_29)
  );
  defparam DLX_IDinst_RegFile_24_21_4126.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_24_21_4126 (
    .I(DLX_IDinst_WB_data_eff[21]),
    .CE(DLX_IDinst__n0598),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_24_21)
  );
  defparam DLX_IDinst_RegFile_24_13_4127.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_24_13_4127 (
    .I(DLX_IDinst_WB_data_eff[13]),
    .CE(DLX_IDinst__n0598),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_24_13)
  );
  defparam DLX_IDinst_RegFile_16_30_4128.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_16_30_4128 (
    .I(DLX_IDinst_WB_data_eff[30]),
    .CE(DLX_IDinst__n0582),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_16_30)
  );
  defparam DLX_IDinst_RegFile_16_22_4129.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_16_22_4129 (
    .I(DLX_IDinst_WB_data_eff[22]),
    .CE(DLX_IDinst__n0582),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_16_22)
  );
  defparam DLX_IDinst_RegFile_24_22_4130.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_24_22_4130 (
    .I(DLX_IDinst_WB_data_eff[22]),
    .CE(DLX_IDinst__n0598),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_24_22)
  );
  defparam DLX_IDinst_RegFile_16_14_4131.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_16_14_4131 (
    .I(DLX_IDinst_WB_data_eff[14]),
    .CE(DLX_IDinst__n0582),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_16_14)
  );
  defparam DLX_IDinst_RegFile_24_14_4132.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_24_14_4132 (
    .I(DLX_IDinst_WB_data_eff[14]),
    .CE(DLX_IDinst__n0598),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_24_14)
  );
  defparam DLX_IDinst_RegFile_16_23_4133.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_16_23_4133 (
    .I(DLX_IDinst_WB_data_eff[23]),
    .CE(DLX_IDinst__n0582),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_16_23)
  );
  defparam DLX_IDinst_RegFile_24_23_4134.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_24_23_4134 (
    .I(DLX_IDinst_WB_data_eff[23]),
    .CE(DLX_IDinst__n0598),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_24_23)
  );
  defparam DLX_IDinst_RegFile_24_15_4135.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_24_15_4135 (
    .I(DLX_IDinst_WB_data_eff[15]),
    .CE(DLX_IDinst__n0598),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_24_15)
  );
  defparam DLX_IDinst_RegFile_16_31_4136.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_16_31_4136 (
    .I(DLX_IDinst_WB_data_eff[31]),
    .CE(DLX_IDinst__n0582),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_16_31)
  );
  defparam DLX_IDinst_RegFile_24_31_4137.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_24_31_4137 (
    .I(DLX_IDinst_WB_data_eff[31]),
    .CE(DLX_IDinst__n0598),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_24_31)
  );
  defparam DLX_IDinst_RegFile_16_24_4138.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_16_24_4138 (
    .I(DLX_IDinst_WB_data_eff[24]),
    .CE(DLX_IDinst__n0582),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_16_24)
  );
  defparam DLX_IDinst_RegFile_16_16_4139.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_16_16_4139 (
    .I(DLX_IDinst_WB_data_eff[16]),
    .CE(DLX_IDinst__n0582),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_16_16)
  );
  defparam DLX_IDinst_RegFile_24_24_4140.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_24_24_4140 (
    .I(DLX_IDinst_WB_data_eff[24]),
    .CE(DLX_IDinst__n0598),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_24_24)
  );
  defparam DLX_IDinst_RegFile_24_16_4141.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_24_16_4141 (
    .I(DLX_IDinst_WB_data_eff[16]),
    .CE(DLX_IDinst__n0598),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_24_16)
  );
  defparam DLX_IDinst_RegFile_16_25_4142.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_16_25_4142 (
    .I(DLX_IDinst_WB_data_eff[25]),
    .CE(DLX_IDinst__n0582),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_16_25)
  );
  defparam DLX_IDinst_RegFile_16_17_4143.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_16_17_4143 (
    .I(DLX_IDinst_WB_data_eff[17]),
    .CE(DLX_IDinst__n0582),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_16_17)
  );
  defparam DLX_IDinst_RegFile_24_25_4144.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_24_25_4144 (
    .I(DLX_IDinst_WB_data_eff[25]),
    .CE(DLX_IDinst__n0598),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_24_25)
  );
  defparam DLX_IDinst_RegFile_24_17_4145.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_24_17_4145 (
    .I(DLX_IDinst_WB_data_eff[17]),
    .CE(DLX_IDinst__n0598),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_24_17)
  );
  defparam DLX_IDinst_RegFile_16_26_4146.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_16_26_4146 (
    .I(DLX_IDinst_WB_data_eff[26]),
    .CE(DLX_IDinst__n0582),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_16_26)
  );
  defparam DLX_IDinst_RegFile_16_18_4147.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_16_18_4147 (
    .I(DLX_IDinst_WB_data_eff[18]),
    .CE(DLX_IDinst__n0582),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_16_18)
  );
  defparam DLX_IDinst_RegFile_17_10_4148.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_17_10_4148 (
    .I(DLX_IDinst_WB_data_eff[10]),
    .CE(DLX_IDinst__n0584),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_17_10)
  );
  defparam DLX_IDinst_RegFile_24_26_4149.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_24_26_4149 (
    .I(DLX_IDinst_WB_data_eff[26]),
    .CE(DLX_IDinst__n0598),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_24_26)
  );
  defparam DLX_IDinst_RegFile_24_18_4150.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_24_18_4150 (
    .I(DLX_IDinst_WB_data_eff[18]),
    .CE(DLX_IDinst__n0598),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_24_18)
  );
  defparam DLX_IDinst_RegFile_25_10_4151.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_25_10_4151 (
    .I(DLX_IDinst_WB_data_eff[10]),
    .CE(DLX_IDinst__n0600),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_25_10)
  );
  defparam DLX_IDinst_RegFile_16_27_4152.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_16_27_4152 (
    .I(DLX_IDinst_WB_data_eff[27]),
    .CE(DLX_IDinst__n0582),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_16_27)
  );
  defparam DLX_IDinst_RegFile_16_19_4153.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_16_19_4153 (
    .I(DLX_IDinst_WB_data_eff[19]),
    .CE(DLX_IDinst__n0582),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_16_19)
  );
  defparam DLX_IDinst_RegFile_17_11_4154.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_17_11_4154 (
    .I(DLX_IDinst_WB_data_eff[11]),
    .CE(DLX_IDinst__n0584),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_17_11)
  );
  defparam DLX_IDinst_RegFile_24_27_4155.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_24_27_4155 (
    .I(DLX_IDinst_WB_data_eff[27]),
    .CE(DLX_IDinst__n0598),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_24_27)
  );
  defparam DLX_IDinst_RegFile_24_19_4156.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_24_19_4156 (
    .I(DLX_IDinst_WB_data_eff[19]),
    .CE(DLX_IDinst__n0598),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_24_19)
  );
  defparam DLX_IDinst_RegFile_25_11_4157.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_25_11_4157 (
    .I(DLX_IDinst_WB_data_eff[11]),
    .CE(DLX_IDinst__n0600),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_25_11)
  );
  defparam DLX_IDinst_RegFile_16_28_4158.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_16_28_4158 (
    .I(DLX_IDinst_WB_data_eff[28]),
    .CE(DLX_IDinst__n0582),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_16_28)
  );
  defparam DLX_IDinst_RegFile_17_20_4159.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_17_20_4159 (
    .I(DLX_IDinst_WB_data_eff[20]),
    .CE(DLX_IDinst__n0584),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_17_20)
  );
  defparam DLX_IDinst_RegFile_17_12_4160.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_17_12_4160 (
    .I(DLX_IDinst_WB_data_eff[12]),
    .CE(DLX_IDinst__n0584),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_17_12)
  );
  defparam DLX_IDinst_RegFile_24_28_4161.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_24_28_4161 (
    .I(DLX_IDinst_WB_data_eff[28]),
    .CE(DLX_IDinst__n0598),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_24_28)
  );
  defparam DLX_IDinst_RegFile_25_20_4162.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_25_20_4162 (
    .I(DLX_IDinst_WB_data_eff[20]),
    .CE(DLX_IDinst__n0600),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_25_20)
  );
  defparam DLX_IDinst_RegFile_25_12_4163.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_25_12_4163 (
    .I(DLX_IDinst_WB_data_eff[12]),
    .CE(DLX_IDinst__n0600),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_25_12)
  );
  defparam DLX_IDinst_RegFile_16_29_4164.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_16_29_4164 (
    .I(DLX_IDinst_WB_data_eff[29]),
    .CE(DLX_IDinst__n0582),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_16_29)
  );
  defparam DLX_IDinst_RegFile_17_21_4165.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_17_21_4165 (
    .I(DLX_IDinst_WB_data_eff[21]),
    .CE(DLX_IDinst__n0584),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_17_21)
  );
  defparam DLX_IDinst_RegFile_17_13_4166.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_17_13_4166 (
    .I(DLX_IDinst_WB_data_eff[13]),
    .CE(DLX_IDinst__n0584),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_17_13)
  );
  defparam DLX_IDinst_RegFile_24_29_4167.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_24_29_4167 (
    .I(DLX_IDinst_WB_data_eff[29]),
    .CE(DLX_IDinst__n0598),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_24_29)
  );
  defparam DLX_IDinst_RegFile_25_21_4168.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_25_21_4168 (
    .I(DLX_IDinst_WB_data_eff[21]),
    .CE(DLX_IDinst__n0600),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_25_21)
  );
  defparam DLX_IDinst_RegFile_25_13_4169.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_25_13_4169 (
    .I(DLX_IDinst_WB_data_eff[13]),
    .CE(DLX_IDinst__n0600),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_25_13)
  );
  defparam DLX_IDinst_RegFile_17_30_4170.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_17_30_4170 (
    .I(DLX_IDinst_WB_data_eff[30]),
    .CE(DLX_IDinst__n0584),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_17_30)
  );
  defparam DLX_IDinst_RegFile_17_22_4171.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_17_22_4171 (
    .I(DLX_IDinst_WB_data_eff[22]),
    .CE(DLX_IDinst__n0584),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_17_22)
  );
  defparam DLX_IDinst_RegFile_17_14_4172.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_17_14_4172 (
    .I(DLX_IDinst_WB_data_eff[14]),
    .CE(DLX_IDinst__n0584),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_17_14)
  );
  defparam DLX_IDinst_RegFile_25_30_4173.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_25_30_4173 (
    .I(DLX_IDinst_WB_data_eff[30]),
    .CE(DLX_IDinst__n0600),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_25_30)
  );
  defparam DLX_IDinst_RegFile_25_22_4174.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_25_22_4174 (
    .I(DLX_IDinst_WB_data_eff[22]),
    .CE(DLX_IDinst__n0600),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_25_22)
  );
  defparam DLX_IDinst_RegFile_17_23_4175.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_17_23_4175 (
    .I(DLX_IDinst_WB_data_eff[23]),
    .CE(DLX_IDinst__n0584),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_17_23)
  );
  defparam DLX_IDinst_RegFile_25_14_4176.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_25_14_4176 (
    .I(DLX_IDinst_WB_data_eff[14]),
    .CE(DLX_IDinst__n0600),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_25_14)
  );
  defparam DLX_IDinst_RegFile_17_15_4177.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_17_15_4177 (
    .I(DLX_IDinst_WB_data_eff[15]),
    .CE(DLX_IDinst__n0584),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_17_15)
  );
  defparam DLX_IDinst_RegFile_25_23_4178.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_25_23_4178 (
    .I(DLX_IDinst_WB_data_eff[23]),
    .CE(DLX_IDinst__n0600),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_25_23)
  );
  defparam DLX_IDinst_RegFile_25_15_4179.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_25_15_4179 (
    .I(DLX_IDinst_WB_data_eff[15]),
    .CE(DLX_IDinst__n0600),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_25_15)
  );
  defparam DLX_IDinst_RegFile_17_31_4180.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_17_31_4180 (
    .I(DLX_IDinst_WB_data_eff[31]),
    .CE(DLX_IDinst__n0584),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_17_31)
  );
  defparam DLX_IDinst_RegFile_25_31_4181.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_25_31_4181 (
    .I(DLX_IDinst_WB_data_eff[31]),
    .CE(DLX_IDinst__n0600),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_25_31)
  );
  defparam DLX_IDinst_RegFile_17_24_4182.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_17_24_4182 (
    .I(DLX_IDinst_WB_data_eff[24]),
    .CE(DLX_IDinst__n0584),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_17_24)
  );
  defparam DLX_IDinst_RegFile_17_16_4183.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_17_16_4183 (
    .I(DLX_IDinst_WB_data_eff[16]),
    .CE(DLX_IDinst__n0584),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_17_16)
  );
  defparam DLX_IDinst_RegFile_25_24_4184.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_25_24_4184 (
    .I(DLX_IDinst_WB_data_eff[24]),
    .CE(DLX_IDinst__n0600),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_25_24)
  );
  defparam DLX_IDinst_RegFile_25_16_4185.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_25_16_4185 (
    .I(DLX_IDinst_WB_data_eff[16]),
    .CE(DLX_IDinst__n0600),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_25_16)
  );
  defparam DLX_IDinst_RegFile_17_25_4186.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_17_25_4186 (
    .I(DLX_IDinst_WB_data_eff[25]),
    .CE(DLX_IDinst__n0584),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_17_25)
  );
  defparam DLX_IDinst_RegFile_25_25_4187.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_25_25_4187 (
    .I(DLX_IDinst_WB_data_eff[25]),
    .CE(DLX_IDinst__n0600),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_25_25)
  );
  defparam DLX_IDinst_RegFile_25_17_4188.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_25_17_4188 (
    .I(DLX_IDinst_WB_data_eff[17]),
    .CE(DLX_IDinst__n0600),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_25_17)
  );
  defparam DLX_IDinst_RegFile_17_26_4189.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_17_26_4189 (
    .I(DLX_IDinst_WB_data_eff[26]),
    .CE(DLX_IDinst__n0584),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_17_26)
  );
  defparam DLX_IDinst_RegFile_18_10_4190.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_18_10_4190 (
    .I(DLX_IDinst_WB_data_eff[10]),
    .CE(DLX_IDinst__n0586),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_18_10)
  );
  defparam DLX_IDinst_RegFile_25_26_4191.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_25_26_4191 (
    .I(DLX_IDinst_WB_data_eff[26]),
    .CE(DLX_IDinst__n0600),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_25_26)
  );
  defparam DLX_IDinst_RegFile_25_18_4192.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_25_18_4192 (
    .I(DLX_IDinst_WB_data_eff[18]),
    .CE(DLX_IDinst__n0600),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_25_18)
  );
  defparam DLX_IDinst_RegFile_17_27_4193.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_17_27_4193 (
    .I(DLX_IDinst_WB_data_eff[27]),
    .CE(DLX_IDinst__n0584),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_17_27)
  );
  defparam DLX_IDinst_RegFile_17_19_4194.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_17_19_4194 (
    .I(DLX_IDinst_WB_data_eff[19]),
    .CE(DLX_IDinst__n0584),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_17_19)
  );
  defparam DLX_IDinst_RegFile_25_27_4195.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_25_27_4195 (
    .I(DLX_IDinst_WB_data_eff[27]),
    .CE(DLX_IDinst__n0600),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_25_27)
  );
  defparam DLX_IDinst_RegFile_25_19_4196.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_25_19_4196 (
    .I(DLX_IDinst_WB_data_eff[19]),
    .CE(DLX_IDinst__n0600),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_25_19)
  );
  defparam DLX_IDinst_RegFile_26_11_4197.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_26_11_4197 (
    .I(DLX_IDinst_WB_data_eff[11]),
    .CE(DLX_IDinst__n0602),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_8),
    .O(DLX_IDinst_RegFile_26_11)
  );
  defparam DLX_IDinst_RegFile_17_28_4198.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_17_28_4198 (
    .I(DLX_IDinst_WB_data_eff[28]),
    .CE(DLX_IDinst__n0584),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_11),
    .O(DLX_IDinst_RegFile_17_28)
  );
  defparam DLX_IDinst_RegFile_18_20_4199.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_18_20_4199 (
    .I(DLX_IDinst_WB_data_eff[20]),
    .CE(DLX_IDinst__n0586),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_18_20)
  );
  defparam DLX_IDinst_RegFile_18_12_4200.INIT = 1'b0;
  X_SFF DLX_IDinst_RegFile_18_12_4200 (
    .I(DLX_IDinst_WB_data_eff[12]),
    .CE(DLX_IDinst__n0586),
    .CLK(clkdiv),
    .SET(GND),
    .RST(GSR),
    .SSET(GND),
    .SRST(reset_IBUF_10),
    .O(DLX_IDinst_RegFile_18_12)
  );
  X_IPAD \clk/PAD  (
    .PAD(clk)
  );
  X_CKBUF \clk/BUF  (
    .I(clk),
    .O(\clk/new_buffer )
  );
  X_CKBUF \clkbuf2/BUF  (
    .I(clk0),
    .O(clk0buf)
  );
  X_CKBUF \clkbuf3/BUF  (
    .I(clkdivub),
    .O(clkdiv)
  );
  defparam \PWR_GND_0/F .INIT = 16'hFFFF;
  X_LUT4 \PWR_GND_0/F  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\PWR_GND_0/FROM )
  );
  defparam \PWR_GND_0/G .INIT = 16'h0000;
  X_LUT4 \PWR_GND_0/G  (
    .ADR0(VCC),
    .ADR1(VCC),
    .ADR2(VCC),
    .ADR3(VCC),
    .O(\PWR_GND_0/GROM )
  );
  X_BUF \PWR_GND_0/XUSED  (
    .I(\PWR_GND_0/FROM ),
    .O(GLOBAL_LOGIC1)
  );
  X_BUF \PWR_GND_0/YUSED  (
    .I(\PWR_GND_0/GROM ),
    .O(GLOBAL_LOGIC0)
  );
  X_ZERO NlwBlock_DLX_top_GND (
    .O(GND)
  );
  X_ONE NlwBlock_DLX_top_VCC (
    .O(VCC)
  );
endmodule

